
module matrixMult_N_M_1_N8_M32 ( clk, rst, x, y, o );
  input [255:0] x;
  input [2047:0] y;
  output [255:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
         n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
         n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
         n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
         n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
         n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
         n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125,
         n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
         n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
         n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
         n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
         n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
         n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
         n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
         n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
         n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
         n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269,
         n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277,
         n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
         n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293,
         n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
         n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
         n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
         n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
         n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
         n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341,
         n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
         n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
         n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
         n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
         n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
         n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397,
         n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
         n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413,
         n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
         n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
         n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
         n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
         n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461,
         n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469,
         n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
         n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485,
         n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
         n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
         n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509,
         n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
         n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
         n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533,
         n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541,
         n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
         n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557,
         n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
         n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
         n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581,
         n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
         n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
         n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
         n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613,
         n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
         n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
         n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
         n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
         n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
         n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773,
         n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
         n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
         n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
         n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
         n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
         n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
         n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
         n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
         n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845,
         n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
         n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
         n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
         n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
         n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
         n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
         n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
         n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
         n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917,
         n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
         n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
         n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
         n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
         n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
         n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
         n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
         n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
         n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
         n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
         n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
         n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
         n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
         n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
         n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
         n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101,
         n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109,
         n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
         n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
         n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
         n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181,
         n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
         n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
         n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205,
         n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
         n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
         n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
         n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
         n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
         n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
         n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
         n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
         n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
         n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
         n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
         n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301,
         n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
         n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
         n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
         n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
         n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
         n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
         n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
         n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
         n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373,
         n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
         n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
         n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
         n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
         n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
         n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
         n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
         n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
         n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
         n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
         n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
         n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
         n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
         n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
         n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
         n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
         n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
         n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
         n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
         n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
         n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
         n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
         n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
         n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
         n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
         n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
         n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
         n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
         n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
         n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
         n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
         n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
         n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
         n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
         n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
         n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
         n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
         n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
         n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
         n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
         n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
         n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
         n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
         n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
         n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
         n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
         n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
         n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
         n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
         n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
         n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
         n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
         n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
         n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
         n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
         n24158, n24159, n24160;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oi_reg[3][31]  ( .D(N256), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oi_reg[3][30]  ( .D(N255), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oi_reg[3][29]  ( .D(N254), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oi_reg[3][28]  ( .D(N253), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oi_reg[3][27]  ( .D(N252), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oi_reg[3][26]  ( .D(N251), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oi_reg[3][25]  ( .D(N250), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oi_reg[3][24]  ( .D(N249), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oi_reg[3][23]  ( .D(N248), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oi_reg[3][22]  ( .D(N247), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oi_reg[3][21]  ( .D(N246), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oi_reg[3][20]  ( .D(N245), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oi_reg[3][19]  ( .D(N244), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oi_reg[3][18]  ( .D(N243), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oi_reg[3][17]  ( .D(N242), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oi_reg[3][16]  ( .D(N241), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oi_reg[3][15]  ( .D(N240), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oi_reg[3][14]  ( .D(N239), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oi_reg[3][13]  ( .D(N238), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oi_reg[3][12]  ( .D(N237), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oi_reg[3][11]  ( .D(N236), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oi_reg[3][10]  ( .D(N235), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oi_reg[3][9]  ( .D(N234), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oi_reg[3][8]  ( .D(N233), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oi_reg[3][7]  ( .D(N232), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oi_reg[3][6]  ( .D(N231), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oi_reg[3][5]  ( .D(N230), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oi_reg[3][4]  ( .D(N229), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oi_reg[3][3]  ( .D(N228), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oi_reg[3][2]  ( .D(N227), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oi_reg[3][1]  ( .D(N226), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oi_reg[3][0]  ( .D(N225), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oi_reg[4][31]  ( .D(N320), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oi_reg[4][30]  ( .D(N319), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oi_reg[4][29]  ( .D(N318), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oi_reg[4][28]  ( .D(N317), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oi_reg[4][27]  ( .D(N316), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oi_reg[4][26]  ( .D(N315), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oi_reg[4][25]  ( .D(N314), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oi_reg[4][24]  ( .D(N313), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oi_reg[4][23]  ( .D(N312), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oi_reg[4][22]  ( .D(N311), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oi_reg[4][21]  ( .D(N310), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oi_reg[4][20]  ( .D(N309), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oi_reg[4][19]  ( .D(N308), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oi_reg[4][18]  ( .D(N307), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oi_reg[4][17]  ( .D(N306), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oi_reg[4][16]  ( .D(N305), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oi_reg[4][15]  ( .D(N304), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oi_reg[4][14]  ( .D(N303), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oi_reg[4][13]  ( .D(N302), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oi_reg[4][12]  ( .D(N301), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oi_reg[4][11]  ( .D(N300), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oi_reg[4][10]  ( .D(N299), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oi_reg[4][9]  ( .D(N298), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oi_reg[4][8]  ( .D(N297), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oi_reg[4][7]  ( .D(N296), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oi_reg[4][6]  ( .D(N295), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oi_reg[4][5]  ( .D(N294), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oi_reg[4][4]  ( .D(N293), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oi_reg[4][3]  ( .D(N292), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oi_reg[4][2]  ( .D(N291), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oi_reg[4][1]  ( .D(N290), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oi_reg[4][0]  ( .D(N289), .CLK(clk), .RST(rst), .Q(o[128]) );
  DFF \oi_reg[5][31]  ( .D(N384), .CLK(clk), .RST(rst), .Q(o[191]) );
  DFF \oi_reg[5][30]  ( .D(N383), .CLK(clk), .RST(rst), .Q(o[190]) );
  DFF \oi_reg[5][29]  ( .D(N382), .CLK(clk), .RST(rst), .Q(o[189]) );
  DFF \oi_reg[5][28]  ( .D(N381), .CLK(clk), .RST(rst), .Q(o[188]) );
  DFF \oi_reg[5][27]  ( .D(N380), .CLK(clk), .RST(rst), .Q(o[187]) );
  DFF \oi_reg[5][26]  ( .D(N379), .CLK(clk), .RST(rst), .Q(o[186]) );
  DFF \oi_reg[5][25]  ( .D(N378), .CLK(clk), .RST(rst), .Q(o[185]) );
  DFF \oi_reg[5][24]  ( .D(N377), .CLK(clk), .RST(rst), .Q(o[184]) );
  DFF \oi_reg[5][23]  ( .D(N376), .CLK(clk), .RST(rst), .Q(o[183]) );
  DFF \oi_reg[5][22]  ( .D(N375), .CLK(clk), .RST(rst), .Q(o[182]) );
  DFF \oi_reg[5][21]  ( .D(N374), .CLK(clk), .RST(rst), .Q(o[181]) );
  DFF \oi_reg[5][20]  ( .D(N373), .CLK(clk), .RST(rst), .Q(o[180]) );
  DFF \oi_reg[5][19]  ( .D(N372), .CLK(clk), .RST(rst), .Q(o[179]) );
  DFF \oi_reg[5][18]  ( .D(N371), .CLK(clk), .RST(rst), .Q(o[178]) );
  DFF \oi_reg[5][17]  ( .D(N370), .CLK(clk), .RST(rst), .Q(o[177]) );
  DFF \oi_reg[5][16]  ( .D(N369), .CLK(clk), .RST(rst), .Q(o[176]) );
  DFF \oi_reg[5][15]  ( .D(N368), .CLK(clk), .RST(rst), .Q(o[175]) );
  DFF \oi_reg[5][14]  ( .D(N367), .CLK(clk), .RST(rst), .Q(o[174]) );
  DFF \oi_reg[5][13]  ( .D(N366), .CLK(clk), .RST(rst), .Q(o[173]) );
  DFF \oi_reg[5][12]  ( .D(N365), .CLK(clk), .RST(rst), .Q(o[172]) );
  DFF \oi_reg[5][11]  ( .D(N364), .CLK(clk), .RST(rst), .Q(o[171]) );
  DFF \oi_reg[5][10]  ( .D(N363), .CLK(clk), .RST(rst), .Q(o[170]) );
  DFF \oi_reg[5][9]  ( .D(N362), .CLK(clk), .RST(rst), .Q(o[169]) );
  DFF \oi_reg[5][8]  ( .D(N361), .CLK(clk), .RST(rst), .Q(o[168]) );
  DFF \oi_reg[5][7]  ( .D(N360), .CLK(clk), .RST(rst), .Q(o[167]) );
  DFF \oi_reg[5][6]  ( .D(N359), .CLK(clk), .RST(rst), .Q(o[166]) );
  DFF \oi_reg[5][5]  ( .D(N358), .CLK(clk), .RST(rst), .Q(o[165]) );
  DFF \oi_reg[5][4]  ( .D(N357), .CLK(clk), .RST(rst), .Q(o[164]) );
  DFF \oi_reg[5][3]  ( .D(N356), .CLK(clk), .RST(rst), .Q(o[163]) );
  DFF \oi_reg[5][2]  ( .D(N355), .CLK(clk), .RST(rst), .Q(o[162]) );
  DFF \oi_reg[5][1]  ( .D(N354), .CLK(clk), .RST(rst), .Q(o[161]) );
  DFF \oi_reg[5][0]  ( .D(N353), .CLK(clk), .RST(rst), .Q(o[160]) );
  DFF \oi_reg[6][31]  ( .D(N448), .CLK(clk), .RST(rst), .Q(o[223]) );
  DFF \oi_reg[6][30]  ( .D(N447), .CLK(clk), .RST(rst), .Q(o[222]) );
  DFF \oi_reg[6][29]  ( .D(N446), .CLK(clk), .RST(rst), .Q(o[221]) );
  DFF \oi_reg[6][28]  ( .D(N445), .CLK(clk), .RST(rst), .Q(o[220]) );
  DFF \oi_reg[6][27]  ( .D(N444), .CLK(clk), .RST(rst), .Q(o[219]) );
  DFF \oi_reg[6][26]  ( .D(N443), .CLK(clk), .RST(rst), .Q(o[218]) );
  DFF \oi_reg[6][25]  ( .D(N442), .CLK(clk), .RST(rst), .Q(o[217]) );
  DFF \oi_reg[6][24]  ( .D(N441), .CLK(clk), .RST(rst), .Q(o[216]) );
  DFF \oi_reg[6][23]  ( .D(N440), .CLK(clk), .RST(rst), .Q(o[215]) );
  DFF \oi_reg[6][22]  ( .D(N439), .CLK(clk), .RST(rst), .Q(o[214]) );
  DFF \oi_reg[6][21]  ( .D(N438), .CLK(clk), .RST(rst), .Q(o[213]) );
  DFF \oi_reg[6][20]  ( .D(N437), .CLK(clk), .RST(rst), .Q(o[212]) );
  DFF \oi_reg[6][19]  ( .D(N436), .CLK(clk), .RST(rst), .Q(o[211]) );
  DFF \oi_reg[6][18]  ( .D(N435), .CLK(clk), .RST(rst), .Q(o[210]) );
  DFF \oi_reg[6][17]  ( .D(N434), .CLK(clk), .RST(rst), .Q(o[209]) );
  DFF \oi_reg[6][16]  ( .D(N433), .CLK(clk), .RST(rst), .Q(o[208]) );
  DFF \oi_reg[6][15]  ( .D(N432), .CLK(clk), .RST(rst), .Q(o[207]) );
  DFF \oi_reg[6][14]  ( .D(N431), .CLK(clk), .RST(rst), .Q(o[206]) );
  DFF \oi_reg[6][13]  ( .D(N430), .CLK(clk), .RST(rst), .Q(o[205]) );
  DFF \oi_reg[6][12]  ( .D(N429), .CLK(clk), .RST(rst), .Q(o[204]) );
  DFF \oi_reg[6][11]  ( .D(N428), .CLK(clk), .RST(rst), .Q(o[203]) );
  DFF \oi_reg[6][10]  ( .D(N427), .CLK(clk), .RST(rst), .Q(o[202]) );
  DFF \oi_reg[6][9]  ( .D(N426), .CLK(clk), .RST(rst), .Q(o[201]) );
  DFF \oi_reg[6][8]  ( .D(N425), .CLK(clk), .RST(rst), .Q(o[200]) );
  DFF \oi_reg[6][7]  ( .D(N424), .CLK(clk), .RST(rst), .Q(o[199]) );
  DFF \oi_reg[6][6]  ( .D(N423), .CLK(clk), .RST(rst), .Q(o[198]) );
  DFF \oi_reg[6][5]  ( .D(N422), .CLK(clk), .RST(rst), .Q(o[197]) );
  DFF \oi_reg[6][4]  ( .D(N421), .CLK(clk), .RST(rst), .Q(o[196]) );
  DFF \oi_reg[6][3]  ( .D(N420), .CLK(clk), .RST(rst), .Q(o[195]) );
  DFF \oi_reg[6][2]  ( .D(N419), .CLK(clk), .RST(rst), .Q(o[194]) );
  DFF \oi_reg[6][1]  ( .D(N418), .CLK(clk), .RST(rst), .Q(o[193]) );
  DFF \oi_reg[6][0]  ( .D(N417), .CLK(clk), .RST(rst), .Q(o[192]) );
  DFF \oi_reg[7][31]  ( .D(N512), .CLK(clk), .RST(rst), .Q(o[255]) );
  DFF \oi_reg[7][30]  ( .D(N511), .CLK(clk), .RST(rst), .Q(o[254]) );
  DFF \oi_reg[7][29]  ( .D(N510), .CLK(clk), .RST(rst), .Q(o[253]) );
  DFF \oi_reg[7][28]  ( .D(N509), .CLK(clk), .RST(rst), .Q(o[252]) );
  DFF \oi_reg[7][27]  ( .D(N508), .CLK(clk), .RST(rst), .Q(o[251]) );
  DFF \oi_reg[7][26]  ( .D(N507), .CLK(clk), .RST(rst), .Q(o[250]) );
  DFF \oi_reg[7][25]  ( .D(N506), .CLK(clk), .RST(rst), .Q(o[249]) );
  DFF \oi_reg[7][24]  ( .D(N505), .CLK(clk), .RST(rst), .Q(o[248]) );
  DFF \oi_reg[7][23]  ( .D(N504), .CLK(clk), .RST(rst), .Q(o[247]) );
  DFF \oi_reg[7][22]  ( .D(N503), .CLK(clk), .RST(rst), .Q(o[246]) );
  DFF \oi_reg[7][21]  ( .D(N502), .CLK(clk), .RST(rst), .Q(o[245]) );
  DFF \oi_reg[7][20]  ( .D(N501), .CLK(clk), .RST(rst), .Q(o[244]) );
  DFF \oi_reg[7][19]  ( .D(N500), .CLK(clk), .RST(rst), .Q(o[243]) );
  DFF \oi_reg[7][18]  ( .D(N499), .CLK(clk), .RST(rst), .Q(o[242]) );
  DFF \oi_reg[7][17]  ( .D(N498), .CLK(clk), .RST(rst), .Q(o[241]) );
  DFF \oi_reg[7][16]  ( .D(N497), .CLK(clk), .RST(rst), .Q(o[240]) );
  DFF \oi_reg[7][15]  ( .D(N496), .CLK(clk), .RST(rst), .Q(o[239]) );
  DFF \oi_reg[7][14]  ( .D(N495), .CLK(clk), .RST(rst), .Q(o[238]) );
  DFF \oi_reg[7][13]  ( .D(N494), .CLK(clk), .RST(rst), .Q(o[237]) );
  DFF \oi_reg[7][12]  ( .D(N493), .CLK(clk), .RST(rst), .Q(o[236]) );
  DFF \oi_reg[7][11]  ( .D(N492), .CLK(clk), .RST(rst), .Q(o[235]) );
  DFF \oi_reg[7][10]  ( .D(N491), .CLK(clk), .RST(rst), .Q(o[234]) );
  DFF \oi_reg[7][9]  ( .D(N490), .CLK(clk), .RST(rst), .Q(o[233]) );
  DFF \oi_reg[7][8]  ( .D(N489), .CLK(clk), .RST(rst), .Q(o[232]) );
  DFF \oi_reg[7][7]  ( .D(N488), .CLK(clk), .RST(rst), .Q(o[231]) );
  DFF \oi_reg[7][6]  ( .D(N487), .CLK(clk), .RST(rst), .Q(o[230]) );
  DFF \oi_reg[7][5]  ( .D(N486), .CLK(clk), .RST(rst), .Q(o[229]) );
  DFF \oi_reg[7][4]  ( .D(N485), .CLK(clk), .RST(rst), .Q(o[228]) );
  DFF \oi_reg[7][3]  ( .D(N484), .CLK(clk), .RST(rst), .Q(o[227]) );
  DFF \oi_reg[7][2]  ( .D(N483), .CLK(clk), .RST(rst), .Q(o[226]) );
  DFF \oi_reg[7][1]  ( .D(N482), .CLK(clk), .RST(rst), .Q(o[225]) );
  DFF \oi_reg[7][0]  ( .D(N481), .CLK(clk), .RST(rst), .Q(o[224]) );
  XNOR U3 ( .A(n8892), .B(n8891), .Z(n8896) );
  XNOR U4 ( .A(n5523), .B(n5522), .Z(n5460) );
  XNOR U5 ( .A(n20129), .B(n20128), .Z(n20130) );
  NAND U6 ( .A(n17486), .B(n17485), .Z(n1) );
  NANDN U7 ( .A(n17484), .B(n17483), .Z(n2) );
  NAND U8 ( .A(n1), .B(n2), .Z(n17596) );
  NAND U9 ( .A(n14267), .B(n14266), .Z(n3) );
  NAND U10 ( .A(n14265), .B(n14264), .Z(n4) );
  NAND U11 ( .A(n3), .B(n4), .Z(n14447) );
  XNOR U12 ( .A(n8783), .B(n8782), .Z(n8784) );
  XNOR U13 ( .A(n20330), .B(n20329), .Z(n20331) );
  NAND U14 ( .A(n20592), .B(n20591), .Z(n5) );
  NAND U15 ( .A(n20590), .B(n20589), .Z(n6) );
  NAND U16 ( .A(n5), .B(n6), .Z(n20755) );
  NAND U17 ( .A(n20560), .B(n20559), .Z(n7) );
  NAND U18 ( .A(n20557), .B(n20558), .Z(n8) );
  NAND U19 ( .A(n7), .B(n8), .Z(n20685) );
  NAND U20 ( .A(n17841), .B(n17840), .Z(n9) );
  NAND U21 ( .A(n17839), .B(n17838), .Z(n10) );
  NAND U22 ( .A(n9), .B(n10), .Z(n18078) );
  NAND U23 ( .A(n17708), .B(n17707), .Z(n11) );
  NAND U24 ( .A(n17706), .B(n17705), .Z(n12) );
  NAND U25 ( .A(n11), .B(n12), .Z(n17831) );
  NAND U26 ( .A(n14357), .B(n14356), .Z(n13) );
  NANDN U27 ( .A(n14359), .B(n14358), .Z(n14) );
  NAND U28 ( .A(n13), .B(n14), .Z(n14483) );
  NAND U29 ( .A(n14444), .B(n14443), .Z(n15) );
  NAND U30 ( .A(n14442), .B(n14441), .Z(n16) );
  AND U31 ( .A(n15), .B(n16), .Z(n14594) );
  NAND U32 ( .A(n20996), .B(n21016), .Z(n17) );
  NAND U33 ( .A(n20994), .B(n20995), .Z(n18) );
  AND U34 ( .A(n17), .B(n18), .Z(n21047) );
  NAND U35 ( .A(n20670), .B(n20669), .Z(n19) );
  NAND U36 ( .A(n20668), .B(n20667), .Z(n20) );
  AND U37 ( .A(n19), .B(n20), .Z(n20906) );
  XNOR U38 ( .A(n17776), .B(n17775), .Z(n17653) );
  XNOR U39 ( .A(n17898), .B(n17897), .Z(n17818) );
  NAND U40 ( .A(n18267), .B(n18268), .Z(n18272) );
  XNOR U41 ( .A(n15243), .B(n15242), .Z(n15134) );
  XNOR U42 ( .A(n12344), .B(n12343), .Z(n12235) );
  NAND U43 ( .A(n9284), .B(n9283), .Z(n21) );
  NAND U44 ( .A(n9281), .B(n9282), .Z(n22) );
  NAND U45 ( .A(n21), .B(n22), .Z(n9414) );
  XNOR U46 ( .A(n3502), .B(n3501), .Z(n3470) );
  NAND U47 ( .A(n20716), .B(n20715), .Z(n23) );
  NAND U48 ( .A(n20714), .B(n20713), .Z(n24) );
  NAND U49 ( .A(n23), .B(n24), .Z(n20846) );
  XNOR U50 ( .A(n21155), .B(n21154), .Z(n21152) );
  NAND U51 ( .A(n18290), .B(n18289), .Z(n25) );
  NAND U52 ( .A(n18288), .B(n18287), .Z(n26) );
  NAND U53 ( .A(n25), .B(n26), .Z(n18291) );
  NAND U54 ( .A(n9424), .B(n9423), .Z(n27) );
  NANDN U55 ( .A(n9426), .B(n9425), .Z(n28) );
  AND U56 ( .A(n27), .B(n28), .Z(n9704) );
  XNOR U57 ( .A(n9694), .B(n9693), .Z(n9691) );
  XNOR U58 ( .A(n24126), .B(n24125), .Z(n23866) );
  XOR U59 ( .A(n21180), .B(n21179), .Z(n29) );
  NAND U60 ( .A(n29), .B(n21178), .Z(n30) );
  NAND U61 ( .A(n21180), .B(n21179), .Z(n31) );
  AND U62 ( .A(n30), .B(n31), .Z(n21181) );
  XNOR U63 ( .A(n12383), .B(n12382), .Z(n12380) );
  XNOR U64 ( .A(n9468), .B(n9467), .Z(n9465) );
  XNOR U65 ( .A(n6814), .B(n6813), .Z(n6525) );
  XNOR U66 ( .A(n3868), .B(n3867), .Z(n3590) );
  XNOR U67 ( .A(n8636), .B(n8635), .Z(n8639) );
  XNOR U68 ( .A(n8556), .B(n8557), .Z(n8646) );
  XNOR U69 ( .A(n5378), .B(n5377), .Z(n5341) );
  XNOR U70 ( .A(n23120), .B(n23119), .Z(n23121) );
  XNOR U71 ( .A(n19920), .B(n19919), .Z(n19957) );
  XNOR U72 ( .A(n20263), .B(n20262), .Z(n20264) );
  XNOR U73 ( .A(n20259), .B(n20258), .Z(n20269) );
  XNOR U74 ( .A(n16626), .B(n16625), .Z(n16607) );
  XNOR U75 ( .A(n16621), .B(n16620), .Z(n16667) );
  NAND U76 ( .A(n17305), .B(n17304), .Z(n32) );
  NANDN U77 ( .A(n17303), .B(n17302), .Z(n33) );
  NAND U78 ( .A(n32), .B(n33), .Z(n17479) );
  NAND U79 ( .A(n14141), .B(n14140), .Z(n34) );
  NAND U80 ( .A(n14139), .B(n14138), .Z(n35) );
  NAND U81 ( .A(n34), .B(n35), .Z(n14264) );
  XNOR U82 ( .A(n10800), .B(n10799), .Z(n10781) );
  XNOR U83 ( .A(n7931), .B(n7930), .Z(n7951) );
  XNOR U84 ( .A(n8401), .B(n8400), .Z(n8438) );
  XOR U85 ( .A(n8698), .B(n8697), .Z(n8702) );
  XNOR U86 ( .A(n8624), .B(n8623), .Z(n8611) );
  XNOR U87 ( .A(n8904), .B(n8903), .Z(n8897) );
  XNOR U88 ( .A(n5511), .B(n5510), .Z(n5462) );
  XNOR U89 ( .A(n5770), .B(n5769), .Z(n5779) );
  NAND U90 ( .A(n19709), .B(n18878), .Z(n36) );
  NAND U91 ( .A(n18877), .B(n19043), .Z(n37) );
  NAND U92 ( .A(n36), .B(n37), .Z(n18968) );
  NAND U93 ( .A(n18901), .B(n18900), .Z(n38) );
  NAND U94 ( .A(n19017), .B(n20453), .Z(n39) );
  NAND U95 ( .A(n38), .B(n39), .Z(n18924) );
  XNOR U96 ( .A(n20143), .B(n20142), .Z(n20131) );
  XNOR U97 ( .A(n16817), .B(n16816), .Z(n16767) );
  XOR U98 ( .A(n16756), .B(n16755), .Z(n16760) );
  NAND U99 ( .A(n17360), .B(n17359), .Z(n40) );
  NAND U100 ( .A(n17358), .B(n17357), .Z(n41) );
  NAND U101 ( .A(n40), .B(n41), .Z(n17426) );
  NAND U102 ( .A(n17271), .B(n17270), .Z(n42) );
  NANDN U103 ( .A(n17406), .B(n17269), .Z(n43) );
  NAND U104 ( .A(n42), .B(n43), .Z(n17421) );
  XNOR U105 ( .A(n17604), .B(n17605), .Z(n17607) );
  NAND U106 ( .A(n17416), .B(n17415), .Z(n44) );
  NAND U107 ( .A(n17413), .B(n17414), .Z(n45) );
  AND U108 ( .A(n44), .B(n45), .Z(n17626) );
  XNOR U109 ( .A(n13051), .B(n13050), .Z(n13014) );
  NAND U110 ( .A(n14285), .B(n14284), .Z(n46) );
  NAND U111 ( .A(n14283), .B(n14282), .Z(n47) );
  NAND U112 ( .A(n46), .B(n47), .Z(n14357) );
  NAND U113 ( .A(n14490), .B(n14489), .Z(n48) );
  NAND U114 ( .A(n14488), .B(n14487), .Z(n49) );
  AND U115 ( .A(n48), .B(n49), .Z(n14660) );
  XNOR U116 ( .A(n10157), .B(n10156), .Z(n10150) );
  XNOR U117 ( .A(n10230), .B(n10229), .Z(n10231) );
  XNOR U118 ( .A(n10995), .B(n10994), .Z(n10945) );
  XNOR U119 ( .A(n8083), .B(n8082), .Z(n8037) );
  XNOR U120 ( .A(n8574), .B(n8573), .Z(n8576) );
  XNOR U121 ( .A(n8979), .B(n8978), .Z(n8847) );
  XNOR U122 ( .A(n8933), .B(n8932), .Z(n8934) );
  XNOR U123 ( .A(n4024), .B(o[39]), .Z(n4019) );
  XNOR U124 ( .A(n5312), .B(n5311), .Z(n5387) );
  XOR U125 ( .A(n5324), .B(n5323), .Z(n5393) );
  XNOR U126 ( .A(n5627), .B(n5626), .Z(n5628) );
  XNOR U127 ( .A(n21688), .B(n21687), .Z(n21675) );
  XNOR U128 ( .A(n23502), .B(n23501), .Z(n23503) );
  XNOR U129 ( .A(n23496), .B(n23495), .Z(n23497) );
  XNOR U130 ( .A(n23590), .B(n23589), .Z(n23644) );
  XNOR U131 ( .A(n23567), .B(n23566), .Z(n23650) );
  NAND U132 ( .A(n18967), .B(n18966), .Z(n50) );
  NAND U133 ( .A(n18965), .B(n19341), .Z(n51) );
  AND U134 ( .A(n50), .B(n51), .Z(n19066) );
  XNOR U135 ( .A(n19063), .B(n19062), .Z(n19055) );
  XNOR U136 ( .A(n19309), .B(n19308), .Z(n19380) );
  XNOR U137 ( .A(n20251), .B(n20250), .Z(n20208) );
  XNOR U138 ( .A(n20332), .B(n20331), .Z(n20323) );
  XNOR U139 ( .A(n20429), .B(n20428), .Z(n20431) );
  NAND U140 ( .A(n20547), .B(n20546), .Z(n52) );
  NAND U141 ( .A(n20545), .B(n20544), .Z(n53) );
  NAND U142 ( .A(n52), .B(n53), .Z(n20728) );
  NAND U143 ( .A(n20674), .B(n20673), .Z(n54) );
  NAND U144 ( .A(n20672), .B(n20671), .Z(n55) );
  NAND U145 ( .A(n54), .B(n55), .Z(n20935) );
  NAND U146 ( .A(n20556), .B(n20555), .Z(n56) );
  NAND U147 ( .A(n20554), .B(n20553), .Z(n57) );
  NAND U148 ( .A(n56), .B(n57), .Z(n20684) );
  XNOR U149 ( .A(n15853), .B(n15852), .Z(n15854) );
  XNOR U150 ( .A(n15967), .B(n15966), .Z(n15970) );
  XNOR U151 ( .A(n16293), .B(n16292), .Z(n16284) );
  NAND U152 ( .A(n16331), .B(n16330), .Z(n58) );
  NAND U153 ( .A(n16329), .B(n16328), .Z(n59) );
  NAND U154 ( .A(n58), .B(n59), .Z(n16481) );
  NAND U155 ( .A(n17611), .B(n17610), .Z(n60) );
  NAND U156 ( .A(n17609), .B(n17608), .Z(n61) );
  NAND U157 ( .A(n60), .B(n61), .Z(n17709) );
  XNOR U158 ( .A(n17673), .B(n17672), .Z(n17756) );
  NAND U159 ( .A(n17695), .B(n17694), .Z(n62) );
  NAND U160 ( .A(n17693), .B(n17692), .Z(n63) );
  NAND U161 ( .A(n62), .B(n63), .Z(n17887) );
  NAND U162 ( .A(n17837), .B(n17836), .Z(n64) );
  NAND U163 ( .A(n17835), .B(n17834), .Z(n65) );
  NAND U164 ( .A(n64), .B(n65), .Z(n18077) );
  NAND U165 ( .A(n17704), .B(n17703), .Z(n66) );
  NAND U166 ( .A(n17702), .B(n17701), .Z(n67) );
  NAND U167 ( .A(n66), .B(n67), .Z(n17830) );
  XNOR U168 ( .A(n10297), .B(n10296), .Z(n10298) );
  XNOR U169 ( .A(n8034), .B(n8033), .Z(n8092) );
  NAND U170 ( .A(n9204), .B(n9203), .Z(n68) );
  NAND U171 ( .A(n9202), .B(n9201), .Z(n69) );
  NAND U172 ( .A(n68), .B(n69), .Z(n9438) );
  NAND U173 ( .A(n9181), .B(n9180), .Z(n70) );
  NAND U174 ( .A(n9179), .B(n9178), .Z(n71) );
  NAND U175 ( .A(n70), .B(n71), .Z(n9461) );
  NAND U176 ( .A(n9045), .B(n9044), .Z(n72) );
  NAND U177 ( .A(n9043), .B(n9042), .Z(n73) );
  NAND U178 ( .A(n72), .B(n73), .Z(n9198) );
  XNOR U179 ( .A(n9252), .B(n9251), .Z(n9159) );
  XNOR U180 ( .A(n1845), .B(n1844), .Z(n1895) );
  XNOR U181 ( .A(n23805), .B(n23804), .Z(n23720) );
  XNOR U182 ( .A(n20737), .B(n20736), .Z(n20738) );
  NAND U183 ( .A(n20765), .B(n20764), .Z(n74) );
  NAND U184 ( .A(n20763), .B(n20762), .Z(n75) );
  NAND U185 ( .A(n74), .B(n75), .Z(n20897) );
  XNOR U186 ( .A(n16313), .B(n16312), .Z(n16314) );
  NAND U187 ( .A(n16488), .B(n16487), .Z(n76) );
  NAND U188 ( .A(n16486), .B(n16485), .Z(n77) );
  NAND U189 ( .A(n76), .B(n77), .Z(n16500) );
  NAND U190 ( .A(n16506), .B(n16505), .Z(n78) );
  NANDN U191 ( .A(n16504), .B(n16503), .Z(n79) );
  AND U192 ( .A(n78), .B(n79), .Z(n16719) );
  NAND U193 ( .A(n17878), .B(n17877), .Z(n80) );
  NAND U194 ( .A(n17876), .B(n17875), .Z(n81) );
  NAND U195 ( .A(n80), .B(n81), .Z(n17991) );
  XOR U196 ( .A(n17809), .B(n17808), .Z(n17803) );
  NAND U197 ( .A(n17747), .B(n17746), .Z(n82) );
  NAND U198 ( .A(n17745), .B(n17744), .Z(n83) );
  NAND U199 ( .A(n82), .B(n83), .Z(n17908) );
  NAND U200 ( .A(n18057), .B(n18056), .Z(n84) );
  NANDN U201 ( .A(n18059), .B(n18058), .Z(n85) );
  AND U202 ( .A(n84), .B(n85), .Z(n18289) );
  NAND U203 ( .A(n17850), .B(n17849), .Z(n86) );
  NAND U204 ( .A(n17848), .B(n17847), .Z(n87) );
  AND U205 ( .A(n86), .B(n87), .Z(n18046) );
  NAND U206 ( .A(n14597), .B(n14596), .Z(n88) );
  NAND U207 ( .A(n14595), .B(n14594), .Z(n89) );
  AND U208 ( .A(n88), .B(n89), .Z(n14608) );
  XNOR U209 ( .A(n15132), .B(n15131), .Z(n15133) );
  XOR U210 ( .A(n15138), .B(n15137), .Z(n15140) );
  XNOR U211 ( .A(n12233), .B(n12232), .Z(n12234) );
  XOR U212 ( .A(n12239), .B(n12238), .Z(n12241) );
  XOR U213 ( .A(n12050), .B(n12049), .Z(n12044) );
  XNOR U214 ( .A(n7020), .B(n7019), .Z(n7033) );
  XNOR U215 ( .A(n9264), .B(n9263), .Z(n9164) );
  XNOR U216 ( .A(n9418), .B(n9417), .Z(n9419) );
  NAND U217 ( .A(n9280), .B(n9279), .Z(n90) );
  NAND U218 ( .A(n9277), .B(n9278), .Z(n91) );
  NAND U219 ( .A(n90), .B(n91), .Z(n9413) );
  XNOR U220 ( .A(n9668), .B(n9667), .Z(n9665) );
  XNOR U221 ( .A(n4071), .B(n4070), .Z(n4084) );
  XNOR U222 ( .A(n3470), .B(n3469), .Z(n3471) );
  XNOR U223 ( .A(n18388), .B(n18387), .Z(n18396) );
  NAND U224 ( .A(n20981), .B(n20980), .Z(n92) );
  NAND U225 ( .A(n20982), .B(n20983), .Z(n93) );
  AND U226 ( .A(n92), .B(n93), .Z(n94) );
  XOR U227 ( .A(n21047), .B(n21046), .Z(n95) );
  XNOR U228 ( .A(n20993), .B(n20992), .Z(n96) );
  XNOR U229 ( .A(n95), .B(n96), .Z(n97) );
  XOR U230 ( .A(n21100), .B(n21099), .Z(n98) );
  XNOR U231 ( .A(n21085), .B(n21084), .Z(n99) );
  XNOR U232 ( .A(n98), .B(n99), .Z(n100) );
  XOR U233 ( .A(n21128), .B(n21127), .Z(n101) );
  XNOR U234 ( .A(n21114), .B(n21113), .Z(n102) );
  XNOR U235 ( .A(n101), .B(n102), .Z(n103) );
  XOR U236 ( .A(n100), .B(n103), .Z(n104) );
  XNOR U237 ( .A(n94), .B(n97), .Z(n105) );
  XNOR U238 ( .A(n104), .B(n105), .Z(n106) );
  NAND U239 ( .A(n20976), .B(n20977), .Z(n107) );
  NAND U240 ( .A(n20978), .B(n20979), .Z(n108) );
  NAND U241 ( .A(n107), .B(n108), .Z(n109) );
  XNOR U242 ( .A(n106), .B(n109), .Z(n21129) );
  NAND U243 ( .A(n20699), .B(n20698), .Z(n110) );
  NAND U244 ( .A(n20697), .B(n20696), .Z(n111) );
  NAND U245 ( .A(n110), .B(n111), .Z(n20829) );
  XNOR U246 ( .A(n15598), .B(n15597), .Z(n15606) );
  NAND U247 ( .A(n17651), .B(n17650), .Z(n112) );
  NAND U248 ( .A(n17648), .B(n17649), .Z(n113) );
  NAND U249 ( .A(n112), .B(n113), .Z(n17793) );
  NAND U250 ( .A(n17918), .B(n17917), .Z(n114) );
  NAND U251 ( .A(n17916), .B(n17915), .Z(n115) );
  NAND U252 ( .A(n114), .B(n115), .Z(n18038) );
  NAND U253 ( .A(n18107), .B(n18106), .Z(n116) );
  NANDN U254 ( .A(n18109), .B(n18108), .Z(n117) );
  AND U255 ( .A(n116), .B(n117), .Z(n118) );
  NANDN U256 ( .A(n18113), .B(n18112), .Z(n119) );
  NANDN U257 ( .A(n18111), .B(n18110), .Z(n120) );
  AND U258 ( .A(n119), .B(n120), .Z(n121) );
  NAND U259 ( .A(n18115), .B(n18114), .Z(n122) );
  NAND U260 ( .A(n18116), .B(n18117), .Z(n123) );
  AND U261 ( .A(n122), .B(n123), .Z(n124) );
  ANDN U262 ( .B(n18272), .A(n18271), .Z(n125) );
  OR U263 ( .A(n18277), .B(n18278), .Z(n126) );
  XNOR U264 ( .A(n125), .B(n126), .Z(n127) );
  XOR U265 ( .A(n18266), .B(n18265), .Z(n128) );
  XNOR U266 ( .A(n18196), .B(n18195), .Z(n129) );
  XNOR U267 ( .A(n128), .B(n129), .Z(n130) );
  XOR U268 ( .A(n127), .B(n130), .Z(n131) );
  XNOR U269 ( .A(n121), .B(n124), .Z(n132) );
  XNOR U270 ( .A(n131), .B(n132), .Z(n133) );
  XNOR U271 ( .A(n118), .B(n133), .Z(n18279) );
  NAND U272 ( .A(n14751), .B(n14750), .Z(n134) );
  NANDN U273 ( .A(n14749), .B(n14748), .Z(n135) );
  AND U274 ( .A(n134), .B(n135), .Z(n14920) );
  XNOR U275 ( .A(n9761), .B(o[99]), .Z(n9763) );
  NAND U276 ( .A(n11886), .B(n11885), .Z(n136) );
  NAND U277 ( .A(n11883), .B(n11884), .Z(n137) );
  AND U278 ( .A(n136), .B(n137), .Z(n12034) );
  OR U279 ( .A(n9230), .B(n9229), .Z(n138) );
  NAND U280 ( .A(n9232), .B(n9231), .Z(n139) );
  NAND U281 ( .A(n138), .B(n139), .Z(n9336) );
  XNOR U282 ( .A(n9704), .B(n9703), .Z(n9701) );
  XNOR U283 ( .A(n9474), .B(n9473), .Z(n9698) );
  NAND U284 ( .A(n4356), .B(n4355), .Z(n140) );
  NANDN U285 ( .A(n4354), .B(n4353), .Z(n141) );
  AND U286 ( .A(n140), .B(n141), .Z(n4508) );
  XNOR U287 ( .A(n6396), .B(n6395), .Z(n6397) );
  XNOR U288 ( .A(n3834), .B(n3833), .Z(n3832) );
  XNOR U289 ( .A(n23866), .B(n23865), .Z(n23861) );
  NANDN U290 ( .A(n21171), .B(n21170), .Z(n142) );
  NANDN U291 ( .A(n21173), .B(n21172), .Z(n143) );
  AND U292 ( .A(n142), .B(n143), .Z(n144) );
  NAND U293 ( .A(n21175), .B(n21174), .Z(n145) );
  NANDN U294 ( .A(n21177), .B(n21176), .Z(n146) );
  AND U295 ( .A(n145), .B(n146), .Z(n147) );
  XNOR U296 ( .A(n144), .B(n147), .Z(n21182) );
  XOR U297 ( .A(n18351), .B(n18352), .Z(n18350) );
  XNOR U298 ( .A(n12635), .B(n12634), .Z(n12663) );
  XNOR U299 ( .A(n9730), .B(n9729), .Z(n9727) );
  NAND U300 ( .A(n4922), .B(n4921), .Z(n148) );
  NANDN U301 ( .A(n4924), .B(n4923), .Z(n149) );
  NAND U302 ( .A(n148), .B(n149), .Z(n5146) );
  XNOR U303 ( .A(n6526), .B(n6525), .Z(n6523) );
  XOR U304 ( .A(n3578), .B(n3579), .Z(n150) );
  NANDN U305 ( .A(n3580), .B(n150), .Z(n151) );
  NAND U306 ( .A(n3578), .B(n3579), .Z(n152) );
  AND U307 ( .A(n151), .B(n152), .Z(n3865) );
  XNOR U308 ( .A(n11505), .B(n11504), .Z(n11506) );
  XNOR U309 ( .A(n8567), .B(n8566), .Z(n8568) );
  XNOR U310 ( .A(n5366), .B(n5365), .Z(n5342) );
  XNOR U311 ( .A(n23122), .B(n23121), .Z(n23131) );
  AND U312 ( .A(n18751), .B(o[203]), .Z(n18826) );
  XNOR U313 ( .A(n19909), .B(o[215]), .Z(n19931) );
  XNOR U314 ( .A(n19913), .B(n19912), .Z(n19959) );
  XOR U315 ( .A(n20290), .B(n20289), .Z(n20268) );
  XNOR U316 ( .A(n20265), .B(n20264), .Z(n20305) );
  XNOR U317 ( .A(n16659), .B(n16658), .Z(n16608) );
  XNOR U318 ( .A(n17126), .B(n17125), .Z(n17163) );
  NAND U319 ( .A(n17348), .B(n17347), .Z(n153) );
  NAND U320 ( .A(n17612), .B(n17468), .Z(n154) );
  NAND U321 ( .A(n153), .B(n154), .Z(n17489) );
  NAND U322 ( .A(n17344), .B(n17343), .Z(n155) );
  NAND U323 ( .A(n17342), .B(n18242), .Z(n156) );
  NAND U324 ( .A(n155), .B(n156), .Z(n17485) );
  XNOR U325 ( .A(n10795), .B(n10794), .Z(n10820) );
  XNOR U326 ( .A(n7926), .B(n7925), .Z(n7912) );
  XNOR U327 ( .A(n7904), .B(n7903), .Z(n7952) );
  XNOR U328 ( .A(n7886), .B(n8063), .Z(n7945) );
  XNOR U329 ( .A(n8026), .B(n8025), .Z(n8027) );
  XNOR U330 ( .A(n8394), .B(n8393), .Z(n8440) );
  XNOR U331 ( .A(n8726), .B(n8725), .Z(n8727) );
  XNOR U332 ( .A(n8958), .B(n8957), .Z(n8938) );
  XNOR U333 ( .A(n5177), .B(n5176), .Z(n5194) );
  XNOR U334 ( .A(n5517), .B(n5516), .Z(n5504) );
  XNOR U335 ( .A(n5780), .B(n5779), .Z(n5781) );
  XNOR U336 ( .A(n2831), .B(n2830), .Z(n2836) );
  NAND U337 ( .A(n18828), .B(n18827), .Z(n157) );
  NAND U338 ( .A(n19017), .B(n20072), .Z(n158) );
  NAND U339 ( .A(n157), .B(n158), .Z(n18873) );
  XNOR U340 ( .A(n19486), .B(n19485), .Z(n19487) );
  XNOR U341 ( .A(n19599), .B(n19598), .Z(n19553) );
  XNOR U342 ( .A(n20387), .B(n20386), .Z(n20423) );
  AND U343 ( .A(n20469), .B(o[218]), .Z(n20560) );
  XNOR U344 ( .A(n16766), .B(n16765), .Z(n16768) );
  XNOR U345 ( .A(n17307), .B(n17306), .Z(n17309) );
  NAND U346 ( .A(n17352), .B(n17351), .Z(n159) );
  NAND U347 ( .A(n17350), .B(n17349), .Z(n160) );
  AND U348 ( .A(n159), .B(n160), .Z(n17419) );
  NAND U349 ( .A(n17412), .B(n17411), .Z(n161) );
  NANDN U350 ( .A(n17410), .B(n17409), .Z(n162) );
  AND U351 ( .A(n161), .B(n162), .Z(n17624) );
  NAND U352 ( .A(n14125), .B(n14124), .Z(n163) );
  NANDN U353 ( .A(n14127), .B(n14126), .Z(n164) );
  NAND U354 ( .A(n163), .B(n164), .Z(n14311) );
  NAND U355 ( .A(n14387), .B(n14386), .Z(n165) );
  NANDN U356 ( .A(n14389), .B(n14388), .Z(n166) );
  NAND U357 ( .A(n165), .B(n166), .Z(n14515) );
  NAND U358 ( .A(n14281), .B(n14280), .Z(n167) );
  NAND U359 ( .A(n14279), .B(n14278), .Z(n168) );
  NAND U360 ( .A(n167), .B(n168), .Z(n14356) );
  NAND U361 ( .A(n14271), .B(n14270), .Z(n169) );
  NAND U362 ( .A(n14269), .B(n14268), .Z(n170) );
  NAND U363 ( .A(n169), .B(n170), .Z(n14445) );
  NAND U364 ( .A(n14247), .B(n14246), .Z(n171) );
  NAND U365 ( .A(n14245), .B(n14244), .Z(n172) );
  NAND U366 ( .A(n171), .B(n172), .Z(n14396) );
  XNOR U367 ( .A(n10182), .B(n10181), .Z(n10151) );
  XNOR U368 ( .A(n10808), .B(n10807), .Z(n10814) );
  XNOR U369 ( .A(n10904), .B(n10903), .Z(n10906) );
  XOR U370 ( .A(n10934), .B(n10933), .Z(n10938) );
  XNOR U371 ( .A(n11124), .B(n11123), .Z(n11126) );
  XNOR U372 ( .A(n7939), .B(n7938), .Z(n7918) );
  XNOR U373 ( .A(n8089), .B(n8088), .Z(n8039) );
  XNOR U374 ( .A(n8222), .B(n8221), .Z(n8224) );
  XNOR U375 ( .A(n8618), .B(n8617), .Z(n8591) );
  XNOR U376 ( .A(n8612), .B(n8611), .Z(n8597) );
  XNOR U377 ( .A(n8848), .B(n8847), .Z(n8849) );
  XNOR U378 ( .A(n8973), .B(n8972), .Z(n8935) );
  XOR U379 ( .A(n9099), .B(n9098), .Z(n9109) );
  XNOR U380 ( .A(n5015), .B(n5014), .Z(n5016) );
  XNOR U381 ( .A(n5349), .B(n5348), .Z(n5321) );
  XOR U382 ( .A(n5931), .B(n5930), .Z(n5933) );
  XNOR U383 ( .A(n5921), .B(n5920), .Z(n5925) );
  XNOR U384 ( .A(n1851), .B(n1850), .Z(n1856) );
  XNOR U385 ( .A(n21674), .B(n21673), .Z(n21676) );
  XNOR U386 ( .A(n22411), .B(n22410), .Z(n22413) );
  NAND U387 ( .A(n23296), .B(n23295), .Z(n173) );
  XOR U388 ( .A(n23296), .B(n23295), .Z(n174) );
  NAND U389 ( .A(n174), .B(n23297), .Z(n175) );
  NAND U390 ( .A(n173), .B(n175), .Z(n23498) );
  XNOR U391 ( .A(n23490), .B(n23489), .Z(n23491) );
  XNOR U392 ( .A(n23609), .B(n23608), .Z(n23610) );
  XNOR U393 ( .A(n23570), .B(n23571), .Z(n23651) );
  XNOR U394 ( .A(n23536), .B(n23535), .Z(n23537) );
  NAND U395 ( .A(n18899), .B(n18898), .Z(n176) );
  NAND U396 ( .A(n19030), .B(n19697), .Z(n177) );
  NAND U397 ( .A(n176), .B(n177), .Z(n18925) );
  NAND U398 ( .A(n18888), .B(n18887), .Z(n178) );
  NAND U399 ( .A(n18886), .B(n18885), .Z(n179) );
  AND U400 ( .A(n178), .B(n179), .Z(n18917) );
  NAND U401 ( .A(n18971), .B(n18970), .Z(n180) );
  NAND U402 ( .A(n18969), .B(n18968), .Z(n181) );
  AND U403 ( .A(n180), .B(n181), .Z(n19068) );
  NAND U404 ( .A(n18930), .B(n18929), .Z(n182) );
  NAND U405 ( .A(n18928), .B(n18927), .Z(n183) );
  NAND U406 ( .A(n182), .B(n183), .Z(n19054) );
  XNOR U407 ( .A(n19353), .B(n19352), .Z(n19376) );
  XNOR U408 ( .A(n19381), .B(n19380), .Z(n19383) );
  XNOR U409 ( .A(n20207), .B(n20206), .Z(n20209) );
  XNOR U410 ( .A(n20525), .B(n20524), .Z(n20607) );
  NAND U411 ( .A(n20588), .B(n20587), .Z(n184) );
  NAND U412 ( .A(n20586), .B(n20585), .Z(n185) );
  NAND U413 ( .A(n184), .B(n185), .Z(n20754) );
  NAND U414 ( .A(n20543), .B(n20542), .Z(n186) );
  NANDN U415 ( .A(n20541), .B(n20540), .Z(n187) );
  NAND U416 ( .A(n186), .B(n187), .Z(n20711) );
  NAND U417 ( .A(n20692), .B(n20693), .Z(n188) );
  NAND U418 ( .A(n20694), .B(n20695), .Z(n189) );
  NAND U419 ( .A(n188), .B(n189), .Z(n20916) );
  NAND U420 ( .A(n20599), .B(n20598), .Z(n190) );
  NAND U421 ( .A(n20597), .B(n20596), .Z(n191) );
  NAND U422 ( .A(n190), .B(n191), .Z(n20669) );
  XNOR U423 ( .A(n15719), .B(o[167]), .Z(n15714) );
  XNOR U424 ( .A(n15971), .B(n15970), .Z(n15972) );
  XNOR U425 ( .A(n16285), .B(n16284), .Z(n16286) );
  XNOR U426 ( .A(n16592), .B(n16591), .Z(n16594) );
  XNOR U427 ( .A(n16762), .B(n16761), .Z(n16820) );
  NAND U428 ( .A(n17424), .B(n17423), .Z(n192) );
  NAND U429 ( .A(n17422), .B(n17421), .Z(n193) );
  AND U430 ( .A(n192), .B(n193), .Z(n17628) );
  NAND U431 ( .A(n17532), .B(n17531), .Z(n194) );
  NAND U432 ( .A(n17530), .B(n17529), .Z(n195) );
  NAND U433 ( .A(n194), .B(n195), .Z(n17755) );
  NAND U434 ( .A(n17554), .B(n17553), .Z(n196) );
  NANDN U435 ( .A(n17556), .B(n17555), .Z(n197) );
  AND U436 ( .A(n196), .B(n197), .Z(n17773) );
  XNOR U437 ( .A(n17712), .B(n17711), .Z(n17767) );
  XOR U438 ( .A(n17752), .B(n17751), .Z(n17762) );
  NAND U439 ( .A(n17855), .B(n17856), .Z(n198) );
  NAND U440 ( .A(n17857), .B(n17858), .Z(n199) );
  NAND U441 ( .A(n198), .B(n199), .Z(n18057) );
  AND U442 ( .A(n18035), .B(o[189]), .Z(n18214) );
  NAND U443 ( .A(n17736), .B(n17735), .Z(n200) );
  NAND U444 ( .A(n17734), .B(n17733), .Z(n201) );
  NAND U445 ( .A(n200), .B(n201), .Z(n17849) );
  XNOR U446 ( .A(n13014), .B(n13013), .Z(n13044) );
  XNOR U447 ( .A(n14793), .B(n14792), .Z(n14894) );
  XOR U448 ( .A(n14890), .B(n14889), .Z(n14900) );
  XNOR U449 ( .A(n10248), .B(n10247), .Z(n10218) );
  XNOR U450 ( .A(n12119), .B(n12118), .Z(n12121) );
  XNOR U451 ( .A(n11902), .B(n11901), .Z(n12001) );
  XNOR U452 ( .A(n7864), .B(n7863), .Z(n7866) );
  XNOR U453 ( .A(n8803), .B(n8802), .Z(n8807) );
  XNOR U454 ( .A(n9123), .B(n9122), .Z(n8984) );
  XNOR U455 ( .A(n9020), .B(n9019), .Z(n9021) );
  NAND U456 ( .A(n9041), .B(n9040), .Z(n202) );
  NAND U457 ( .A(n9039), .B(n9038), .Z(n203) );
  NAND U458 ( .A(n202), .B(n203), .Z(n9197) );
  XNOR U459 ( .A(n9159), .B(n9158), .Z(n9160) );
  XOR U460 ( .A(n4142), .B(n4141), .Z(n4130) );
  XNOR U461 ( .A(n4153), .B(n4152), .Z(n4154) );
  XOR U462 ( .A(n4295), .B(n4294), .Z(n4289) );
  XNOR U463 ( .A(n5695), .B(n5694), .Z(n5701) );
  XOR U464 ( .A(n5714), .B(n5713), .Z(n5707) );
  XNOR U465 ( .A(n6247), .B(n6246), .Z(n6248) );
  XOR U466 ( .A(n6285), .B(n6284), .Z(n6328) );
  NAND U467 ( .A(n2496), .B(n2495), .Z(n204) );
  NANDN U468 ( .A(n2498), .B(n2497), .Z(n205) );
  AND U469 ( .A(n204), .B(n205), .Z(n2623) );
  NAND U470 ( .A(n3179), .B(n3178), .Z(n206) );
  NAND U471 ( .A(n3177), .B(n3176), .Z(n207) );
  NAND U472 ( .A(n206), .B(n207), .Z(n3359) );
  XNOR U473 ( .A(n21418), .B(n21417), .Z(n21420) );
  XNOR U474 ( .A(n23504), .B(n23503), .Z(n23363) );
  XNOR U475 ( .A(n23635), .B(n23634), .Z(n23529) );
  XOR U476 ( .A(n23647), .B(n23646), .Z(n23627) );
  XNOR U477 ( .A(n23617), .B(n23616), .Z(n23657) );
  XNOR U478 ( .A(n23856), .B(n23855), .Z(n23815) );
  XNOR U479 ( .A(n20337), .B(n20336), .Z(n20338) );
  XNOR U480 ( .A(n20739), .B(n20738), .Z(n20766) );
  NAND U481 ( .A(n20761), .B(n20760), .Z(n208) );
  NAND U482 ( .A(n20759), .B(n20758), .Z(n209) );
  NAND U483 ( .A(n208), .B(n209), .Z(n20896) );
  NAND U484 ( .A(n20936), .B(n20935), .Z(n210) );
  NANDN U485 ( .A(n20938), .B(n20937), .Z(n211) );
  AND U486 ( .A(n210), .B(n211), .Z(n21133) );
  NAND U487 ( .A(n20986), .B(n21017), .Z(n212) );
  NAND U488 ( .A(n20984), .B(n20985), .Z(n213) );
  AND U489 ( .A(n212), .B(n213), .Z(n20993) );
  XNOR U490 ( .A(n15677), .B(n15676), .Z(n15669) );
  XOR U491 ( .A(n15823), .B(n15822), .Z(n15797) );
  XNOR U492 ( .A(n15855), .B(n15854), .Z(n15902) );
  NAND U493 ( .A(n16484), .B(n16483), .Z(n214) );
  NAND U494 ( .A(n16482), .B(n16481), .Z(n215) );
  NAND U495 ( .A(n214), .B(n215), .Z(n16499) );
  XOR U496 ( .A(n16858), .B(n16857), .Z(n16851) );
  XNOR U497 ( .A(n16986), .B(n16985), .Z(n16974) );
  NAND U498 ( .A(n17595), .B(n17594), .Z(n216) );
  NAND U499 ( .A(n17593), .B(n17592), .Z(n217) );
  NAND U500 ( .A(n216), .B(n217), .Z(n17654) );
  XNOR U501 ( .A(n17920), .B(n17919), .Z(n17922) );
  XNOR U502 ( .A(n17819), .B(n17818), .Z(n17820) );
  NAND U503 ( .A(n17865), .B(n17864), .Z(n218) );
  NAND U504 ( .A(n17863), .B(n18005), .Z(n219) );
  AND U505 ( .A(n218), .B(n219), .Z(n18063) );
  NAND U506 ( .A(n17743), .B(n17742), .Z(n220) );
  NAND U507 ( .A(n17741), .B(n17740), .Z(n221) );
  NAND U508 ( .A(n220), .B(n221), .Z(n17907) );
  NAND U509 ( .A(n18078), .B(n18077), .Z(n222) );
  NANDN U510 ( .A(n18080), .B(n18079), .Z(n223) );
  AND U511 ( .A(n222), .B(n223), .Z(n18282) );
  NAND U512 ( .A(n18026), .B(n18025), .Z(n224) );
  NAND U513 ( .A(n18236), .B(n18024), .Z(n225) );
  NAND U514 ( .A(n224), .B(n225), .Z(n18117) );
  NAND U515 ( .A(n17833), .B(n17832), .Z(n226) );
  NAND U516 ( .A(n17831), .B(n17830), .Z(n227) );
  AND U517 ( .A(n226), .B(n227), .Z(n18048) );
  NAND U518 ( .A(n17862), .B(n17861), .Z(n228) );
  NAND U519 ( .A(n17860), .B(n17859), .Z(n229) );
  NAND U520 ( .A(n228), .B(n229), .Z(n17972) );
  XNOR U521 ( .A(n13833), .B(n13832), .Z(n13836) );
  XNOR U522 ( .A(n14474), .B(n14473), .Z(n14602) );
  XNOR U523 ( .A(n15051), .B(n15050), .Z(n14945) );
  XNOR U524 ( .A(n10226), .B(n10225), .Z(n10213) );
  XOR U525 ( .A(n11132), .B(n11131), .Z(n11027) );
  XNOR U526 ( .A(n11167), .B(n11166), .Z(n11155) );
  XNOR U527 ( .A(n12153), .B(n12152), .Z(n12186) );
  XNOR U528 ( .A(n7024), .B(n7023), .Z(n7025) );
  XNOR U529 ( .A(n8261), .B(n8260), .Z(n8249) );
  XNOR U530 ( .A(n9165), .B(n9164), .Z(n9167) );
  XNOR U531 ( .A(n4075), .B(n4074), .Z(n4076) );
  XOR U532 ( .A(n5541), .B(n5540), .Z(n5419) );
  XNOR U533 ( .A(n6272), .B(n6271), .Z(n6303) );
  XNOR U534 ( .A(n6520), .B(n6519), .Z(n6482) );
  NAND U535 ( .A(n6505), .B(n6608), .Z(n230) );
  XOR U536 ( .A(n6505), .B(n6608), .Z(n231) );
  NAND U537 ( .A(n231), .B(n6506), .Z(n232) );
  NAND U538 ( .A(n230), .B(n232), .Z(n6755) );
  XNOR U539 ( .A(n1600), .B(n1599), .Z(n1602) );
  XNOR U540 ( .A(n1911), .B(n1910), .Z(n1912) );
  NAND U541 ( .A(n3445), .B(n3700), .Z(n233) );
  XOR U542 ( .A(n3445), .B(n3700), .Z(n234) );
  NAND U543 ( .A(n234), .B(n3446), .Z(n235) );
  NAND U544 ( .A(n233), .B(n235), .Z(n3815) );
  XNOR U545 ( .A(n3622), .B(n3621), .Z(n3619) );
  XNOR U546 ( .A(n3557), .B(n3556), .Z(n3472) );
  XNOR U547 ( .A(n21248), .B(n21247), .Z(n21252) );
  XNOR U548 ( .A(n23809), .B(n23808), .Z(n23810) );
  XNOR U549 ( .A(n23688), .B(n23687), .Z(n23689) );
  XNOR U550 ( .A(n24096), .B(n24095), .Z(n24116) );
  XNOR U551 ( .A(n18393), .B(o[195]), .Z(n18395) );
  XNOR U552 ( .A(n20507), .B(n20506), .Z(n20630) );
  XNOR U553 ( .A(n20996), .B(n20926), .Z(n236) );
  XNOR U554 ( .A(n20925), .B(n236), .Z(n20850) );
  NAND U555 ( .A(n20902), .B(n20901), .Z(n237) );
  NANDN U556 ( .A(n20904), .B(n20903), .Z(n238) );
  NAND U557 ( .A(n237), .B(n238), .Z(n21175) );
  NAND U558 ( .A(n20833), .B(n20832), .Z(n239) );
  NAND U559 ( .A(n20830), .B(n20831), .Z(n240) );
  NAND U560 ( .A(n239), .B(n240), .Z(n20950) );
  XNOR U561 ( .A(n15603), .B(o[163]), .Z(n15605) );
  NAND U562 ( .A(n17914), .B(n17913), .Z(n241) );
  NAND U563 ( .A(n17912), .B(n17911), .Z(n242) );
  NAND U564 ( .A(n241), .B(n242), .Z(n18037) );
  XOR U565 ( .A(n18324), .B(n18323), .Z(n18322) );
  NAND U566 ( .A(n17989), .B(n17988), .Z(n243) );
  NAND U567 ( .A(n17986), .B(n17987), .Z(n244) );
  AND U568 ( .A(n243), .B(n244), .Z(n18094) );
  NAND U569 ( .A(n14611), .B(n14610), .Z(n245) );
  NAND U570 ( .A(n14608), .B(n14609), .Z(n246) );
  AND U571 ( .A(n245), .B(n246), .Z(n14923) );
  XNOR U572 ( .A(n15225), .B(n15224), .Z(n15126) );
  XOR U573 ( .A(n15548), .B(n15547), .Z(n247) );
  XNOR U574 ( .A(n15549), .B(n247), .Z(n15534) );
  XNOR U575 ( .A(n9756), .B(n9755), .Z(n9764) );
  XOR U576 ( .A(n10009), .B(n10010), .Z(n248) );
  NANDN U577 ( .A(n10011), .B(n248), .Z(n249) );
  NAND U578 ( .A(n10009), .B(n10010), .Z(n250) );
  AND U579 ( .A(n249), .B(n250), .Z(n10071) );
  XNOR U580 ( .A(n10293), .B(n10292), .Z(n10366) );
  XNOR U581 ( .A(n12326), .B(n12325), .Z(n12221) );
  XOR U582 ( .A(n12643), .B(n12642), .Z(n12641) );
  NAND U583 ( .A(n6872), .B(n6871), .Z(n251) );
  NANDN U584 ( .A(n6975), .B(n6966), .Z(n252) );
  AND U585 ( .A(n251), .B(n252), .Z(n6904) );
  XNOR U586 ( .A(n7033), .B(n7032), .Z(n7034) );
  XOR U587 ( .A(n8127), .B(n8126), .Z(n8244) );
  XOR U588 ( .A(n9708), .B(n9707), .Z(n9702) );
  NAND U589 ( .A(n9236), .B(n9235), .Z(n253) );
  NAND U590 ( .A(n9234), .B(n9233), .Z(n254) );
  NAND U591 ( .A(n253), .B(n254), .Z(n9367) );
  XNOR U592 ( .A(n3899), .B(o[35]), .Z(n3901) );
  XNOR U593 ( .A(n4084), .B(n4083), .Z(n4085) );
  XNOR U594 ( .A(n5029), .B(n5028), .Z(n4921) );
  XNOR U595 ( .A(n6392), .B(n6391), .Z(n6398) );
  XNOR U596 ( .A(n1089), .B(n1088), .Z(n1091) );
  XOR U597 ( .A(n1201), .B(n1200), .Z(n1191) );
  NAND U598 ( .A(n2401), .B(n2400), .Z(n255) );
  NANDN U599 ( .A(n2399), .B(n2398), .Z(n256) );
  AND U600 ( .A(n255), .B(n256), .Z(n2637) );
  XNOR U601 ( .A(n3083), .B(n3082), .Z(n3085) );
  XNOR U602 ( .A(n3610), .B(n3609), .Z(n3607) );
  XOR U603 ( .A(n3858), .B(n3857), .Z(n3856) );
  NAND U604 ( .A(n21591), .B(n21592), .Z(n257) );
  XOR U605 ( .A(n21591), .B(n21592), .Z(n258) );
  NANDN U606 ( .A(n21590), .B(n258), .Z(n259) );
  NAND U607 ( .A(n257), .B(n259), .Z(n21607) );
  XOR U608 ( .A(n23674), .B(n23675), .Z(n260) );
  NANDN U609 ( .A(n23676), .B(n260), .Z(n261) );
  NAND U610 ( .A(n23674), .B(n23675), .Z(n262) );
  AND U611 ( .A(n261), .B(n262), .Z(n23685) );
  XNOR U612 ( .A(n23862), .B(n23861), .Z(n23859) );
  XOR U613 ( .A(n19187), .B(n19186), .Z(n263) );
  NANDN U614 ( .A(n19188), .B(n263), .Z(n264) );
  NAND U615 ( .A(n19187), .B(n19186), .Z(n265) );
  AND U616 ( .A(n264), .B(n265), .Z(n19393) );
  NAND U617 ( .A(n20829), .B(n20828), .Z(n266) );
  NAND U618 ( .A(n20826), .B(n20827), .Z(n267) );
  AND U619 ( .A(n266), .B(n267), .Z(n20943) );
  NAND U620 ( .A(n15791), .B(n15792), .Z(n268) );
  XOR U621 ( .A(n15791), .B(n15792), .Z(n269) );
  NANDN U622 ( .A(n15790), .B(n269), .Z(n270) );
  NAND U623 ( .A(n268), .B(n270), .Z(n15843) );
  NAND U624 ( .A(n16142), .B(n16143), .Z(n271) );
  XOR U625 ( .A(n16142), .B(n16143), .Z(n272) );
  NANDN U626 ( .A(n16141), .B(n272), .Z(n273) );
  NAND U627 ( .A(n271), .B(n273), .Z(n16309) );
  XOR U628 ( .A(n16497), .B(n16496), .Z(n274) );
  NANDN U629 ( .A(n16495), .B(n274), .Z(n275) );
  NAND U630 ( .A(n16497), .B(n16496), .Z(n276) );
  AND U631 ( .A(n275), .B(n276), .Z(n16598) );
  NAND U632 ( .A(n16841), .B(n16838), .Z(n277) );
  NANDN U633 ( .A(n16841), .B(n16840), .Z(n278) );
  NANDN U634 ( .A(n16839), .B(n278), .Z(n279) );
  NAND U635 ( .A(n277), .B(n279), .Z(n16964) );
  XOR U636 ( .A(n17927), .B(n17926), .Z(n280) );
  NANDN U637 ( .A(n17928), .B(n280), .Z(n281) );
  NAND U638 ( .A(n17927), .B(n17926), .Z(n282) );
  AND U639 ( .A(n281), .B(n282), .Z(n18344) );
  NAND U640 ( .A(n13527), .B(n13528), .Z(n283) );
  XOR U641 ( .A(n13527), .B(n13528), .Z(n284) );
  NANDN U642 ( .A(n13526), .B(n284), .Z(n285) );
  NAND U643 ( .A(n283), .B(n285), .Z(n13733) );
  NAND U644 ( .A(n14341), .B(n14342), .Z(n286) );
  XOR U645 ( .A(n14341), .B(n14342), .Z(n287) );
  NANDN U646 ( .A(n14340), .B(n287), .Z(n288) );
  NAND U647 ( .A(n286), .B(n288), .Z(n14467) );
  XOR U648 ( .A(n15282), .B(n15281), .Z(n15280) );
  XOR U649 ( .A(n12026), .B(n12025), .Z(n289) );
  NANDN U650 ( .A(n12024), .B(n289), .Z(n290) );
  NAND U651 ( .A(n12026), .B(n12025), .Z(n291) );
  AND U652 ( .A(n290), .B(n291), .Z(n12039) );
  NAND U653 ( .A(n12037), .B(n12036), .Z(n292) );
  NAND U654 ( .A(n12034), .B(n12035), .Z(n293) );
  AND U655 ( .A(n292), .B(n293), .Z(n12200) );
  NANDN U656 ( .A(n12649), .B(n12648), .Z(n12653) );
  XOR U657 ( .A(n6883), .B(n6884), .Z(n294) );
  NANDN U658 ( .A(n6885), .B(n294), .Z(n295) );
  NAND U659 ( .A(n6883), .B(n6884), .Z(n296) );
  AND U660 ( .A(n295), .B(n296), .Z(n6909) );
  NAND U661 ( .A(n7672), .B(n7673), .Z(n297) );
  XOR U662 ( .A(n7672), .B(n7673), .Z(n298) );
  NANDN U663 ( .A(n7671), .B(n298), .Z(n299) );
  NAND U664 ( .A(n297), .B(n299), .Z(n7876) );
  NAND U665 ( .A(n9480), .B(n9479), .Z(n300) );
  NAND U666 ( .A(n9481), .B(n9482), .Z(n301) );
  AND U667 ( .A(n300), .B(n301), .Z(n302) );
  AND U668 ( .A(n9690), .B(n9689), .Z(n303) );
  NAND U669 ( .A(n9684), .B(n9683), .Z(n304) );
  XNOR U670 ( .A(n303), .B(n304), .Z(n305) );
  AND U671 ( .A(n9488), .B(n9487), .Z(n306) );
  XNOR U672 ( .A(n9678), .B(n9677), .Z(n307) );
  XNOR U673 ( .A(n306), .B(n307), .Z(n308) );
  NAND U674 ( .A(n9692), .B(n9691), .Z(n309) );
  NANDN U675 ( .A(n9694), .B(n9693), .Z(n310) );
  AND U676 ( .A(n309), .B(n310), .Z(n311) );
  NAND U677 ( .A(n9696), .B(n9695), .Z(n312) );
  NAND U678 ( .A(n9697), .B(n9698), .Z(n313) );
  AND U679 ( .A(n312), .B(n313), .Z(n314) );
  XOR U680 ( .A(n311), .B(n314), .Z(n315) );
  XNOR U681 ( .A(n305), .B(n308), .Z(n316) );
  XNOR U682 ( .A(n315), .B(n316), .Z(n317) );
  XNOR U683 ( .A(n302), .B(n317), .Z(n9699) );
  NAND U684 ( .A(n4510), .B(n4509), .Z(n318) );
  NANDN U685 ( .A(n4508), .B(n4507), .Z(n319) );
  NAND U686 ( .A(n318), .B(n319), .Z(n4598) );
  XOR U687 ( .A(n4914), .B(n4915), .Z(n320) );
  NANDN U688 ( .A(n4916), .B(n320), .Z(n321) );
  NAND U689 ( .A(n4914), .B(n4915), .Z(n322) );
  AND U690 ( .A(n321), .B(n322), .Z(n4918) );
  XNOR U691 ( .A(n5152), .B(n5151), .Z(n5148) );
  NAND U692 ( .A(n6364), .B(n6363), .Z(n323) );
  NANDN U693 ( .A(n6362), .B(n6361), .Z(n324) );
  AND U694 ( .A(n323), .B(n324), .Z(n6524) );
  XOR U695 ( .A(n1055), .B(n1054), .Z(n325) );
  NANDN U696 ( .A(n1056), .B(n325), .Z(n326) );
  NAND U697 ( .A(n1055), .B(n1054), .Z(n327) );
  AND U698 ( .A(n326), .B(n327), .Z(n1095) );
  NAND U699 ( .A(n2396), .B(n2397), .Z(n328) );
  XOR U700 ( .A(n2396), .B(n2397), .Z(n329) );
  NAND U701 ( .A(n329), .B(n2395), .Z(n330) );
  NAND U702 ( .A(n328), .B(n330), .Z(n2642) );
  XOR U703 ( .A(n2931), .B(n2932), .Z(n331) );
  NANDN U704 ( .A(n2933), .B(n331), .Z(n332) );
  NAND U705 ( .A(n2931), .B(n2932), .Z(n333) );
  AND U706 ( .A(n332), .B(n333), .Z(n3089) );
  XNOR U707 ( .A(n3866), .B(n3865), .Z(n3863) );
  XNOR U708 ( .A(n19802), .B(n19801), .Z(n19803) );
  XNOR U709 ( .A(n19911), .B(n19910), .Z(n19912) );
  XNOR U710 ( .A(n8392), .B(n8391), .Z(n8393) );
  XNOR U711 ( .A(n8572), .B(o[88]), .Z(n8587) );
  XNOR U712 ( .A(n8629), .B(n8628), .Z(n8640) );
  XNOR U713 ( .A(n8746), .B(n8745), .Z(n8748) );
  XNOR U714 ( .A(n2686), .B(n2685), .Z(n2687) );
  XNOR U715 ( .A(n23126), .B(n23125), .Z(n23127) );
  XNOR U716 ( .A(n23132), .B(n23131), .Z(n23133) );
  XNOR U717 ( .A(n19152), .B(o[208]), .Z(n19167) );
  XNOR U718 ( .A(n19421), .B(n19420), .Z(n19402) );
  XNOR U719 ( .A(n19849), .B(o[214]), .Z(n19828) );
  XNOR U720 ( .A(n19930), .B(n19929), .Z(n19932) );
  XNOR U721 ( .A(n20068), .B(n20067), .Z(n20062) );
  XNOR U722 ( .A(n20227), .B(n20226), .Z(n20232) );
  XOR U723 ( .A(n20318), .B(n20317), .Z(n20320) );
  XNOR U724 ( .A(n20312), .B(n20311), .Z(n20314) );
  XNOR U725 ( .A(n16754), .B(n16753), .Z(n16755) );
  XNOR U726 ( .A(n17136), .B(n17135), .Z(n17137) );
  XNOR U727 ( .A(n13987), .B(n13986), .Z(n14059) );
  NAND U728 ( .A(n14368), .B(n14367), .Z(n334) );
  NANDN U729 ( .A(n14370), .B(n14369), .Z(n335) );
  AND U730 ( .A(n334), .B(n335), .Z(n14506) );
  XNOR U731 ( .A(n10845), .B(n10844), .Z(n10782) );
  XNOR U732 ( .A(n10932), .B(n10931), .Z(n10933) );
  XNOR U733 ( .A(n11507), .B(n11506), .Z(n11451) );
  XNOR U734 ( .A(n8390), .B(o[87]), .Z(n8412) );
  XNOR U735 ( .A(n8551), .B(n8550), .Z(n8545) );
  XNOR U736 ( .A(n8704), .B(n8703), .Z(n8709) );
  XOR U737 ( .A(n8760), .B(n8759), .Z(n8788) );
  XOR U738 ( .A(n8779), .B(n8778), .Z(n8795) );
  XNOR U739 ( .A(n8879), .B(n8880), .Z(n8860) );
  XNOR U740 ( .A(n8946), .B(n8947), .Z(n8884) );
  XNOR U741 ( .A(n8922), .B(n8923), .Z(n8941) );
  XNOR U742 ( .A(n4950), .B(n4949), .Z(n4931) );
  XNOR U743 ( .A(n5194), .B(n5193), .Z(n5250) );
  XNOR U744 ( .A(n5227), .B(n5226), .Z(n5253) );
  XNOR U745 ( .A(n5441), .B(n5440), .Z(n5478) );
  XNOR U746 ( .A(n5304), .B(n5303), .Z(n5306) );
  XNOR U747 ( .A(n5461), .B(n5460), .Z(n5463) );
  XNOR U748 ( .A(n5503), .B(n5502), .Z(n5505) );
  XNOR U749 ( .A(n2482), .B(n2481), .Z(n2448) );
  XNOR U750 ( .A(n2835), .B(n2834), .Z(n2837) );
  XNOR U751 ( .A(n21499), .B(o[234]), .Z(n21510) );
  XNOR U752 ( .A(n21643), .B(n21642), .Z(n21644) );
  XNOR U753 ( .A(n21659), .B(n22273), .Z(n21638) );
  XNOR U754 ( .A(n22288), .B(n22287), .Z(n22326) );
  XNOR U755 ( .A(n22854), .B(n22853), .Z(n22859) );
  XNOR U756 ( .A(n22866), .B(n22865), .Z(n22803) );
  XNOR U757 ( .A(n23229), .B(n23230), .Z(n23212) );
  XNOR U758 ( .A(n23416), .B(n23415), .Z(n23417) );
  XNOR U759 ( .A(n23422), .B(n23421), .Z(n23424) );
  NAND U760 ( .A(n18881), .B(n18880), .Z(n336) );
  NANDN U761 ( .A(n19429), .B(n18879), .Z(n337) );
  NAND U762 ( .A(n336), .B(n337), .Z(n18969) );
  XNOR U763 ( .A(n19474), .B(n19473), .Z(n19476) );
  XNOR U764 ( .A(n19605), .B(n19604), .Z(n19555) );
  XNOR U765 ( .A(n20135), .B(n20134), .Z(n20136) );
  XNOR U766 ( .A(n20306), .B(n20305), .Z(n20307) );
  XNOR U767 ( .A(n20094), .B(n20095), .Z(n20104) );
  XNOR U768 ( .A(n20117), .B(n20116), .Z(n20118) );
  XNOR U769 ( .A(n20271), .B(n20270), .Z(n20242) );
  XNOR U770 ( .A(n20249), .B(n20248), .Z(n20250) );
  XNOR U771 ( .A(n20452), .B(n20453), .Z(n20455) );
  XNOR U772 ( .A(n20423), .B(n20422), .Z(n20424) );
  XNOR U773 ( .A(n20441), .B(n20440), .Z(n20443) );
  XNOR U774 ( .A(n16184), .B(n16183), .Z(n16156) );
  XNOR U775 ( .A(n16432), .B(n16431), .Z(n16443) );
  XNOR U776 ( .A(n16416), .B(n16415), .Z(n16439) );
  XNOR U777 ( .A(n16668), .B(n16667), .Z(n16669) );
  OR U778 ( .A(n16464), .B(n17406), .Z(n338) );
  NANDN U779 ( .A(n16466), .B(n16465), .Z(n339) );
  AND U780 ( .A(n338), .B(n339), .Z(n16564) );
  XNOR U781 ( .A(n16803), .B(n16802), .Z(n16805) );
  XNOR U782 ( .A(n16726), .B(n16725), .Z(n16728) );
  XNOR U783 ( .A(n16929), .B(n16928), .Z(n16931) );
  XNOR U784 ( .A(n17166), .B(n17165), .Z(n17159) );
  XNOR U785 ( .A(n17319), .B(n17318), .Z(n17320) );
  NAND U786 ( .A(n17356), .B(n17355), .Z(n340) );
  NAND U787 ( .A(n17354), .B(n17353), .Z(n341) );
  NAND U788 ( .A(n340), .B(n341), .Z(n17425) );
  NAND U789 ( .A(n17482), .B(n17481), .Z(n342) );
  NAND U790 ( .A(n17480), .B(n17479), .Z(n343) );
  NAND U791 ( .A(n342), .B(n343), .Z(n17598) );
  XNOR U792 ( .A(n14289), .B(n14288), .Z(n14259) );
  NAND U793 ( .A(n14123), .B(n14122), .Z(n344) );
  NANDN U794 ( .A(n14121), .B(n14120), .Z(n345) );
  NAND U795 ( .A(n344), .B(n345), .Z(n14312) );
  NAND U796 ( .A(n14383), .B(n14382), .Z(n346) );
  NANDN U797 ( .A(n14385), .B(n14384), .Z(n347) );
  AND U798 ( .A(n346), .B(n347), .Z(n14516) );
  NAND U799 ( .A(n14243), .B(n14242), .Z(n348) );
  NAND U800 ( .A(n14241), .B(n14240), .Z(n349) );
  NAND U801 ( .A(n348), .B(n349), .Z(n14361) );
  OR U802 ( .A(n14496), .B(n14495), .Z(n350) );
  NAND U803 ( .A(n14497), .B(n14498), .Z(n351) );
  AND U804 ( .A(n350), .B(n351), .Z(n14698) );
  XOR U805 ( .A(n10167), .B(n10168), .Z(n10152) );
  XNOR U806 ( .A(n10246), .B(n10245), .Z(n10247) );
  XNOR U807 ( .A(n10821), .B(n10820), .Z(n10822) );
  XNOR U808 ( .A(n10981), .B(n10980), .Z(n10983) );
  XNOR U809 ( .A(n10944), .B(n10943), .Z(n10946) );
  NAND U810 ( .A(n11604), .B(n11603), .Z(n352) );
  NANDN U811 ( .A(n11606), .B(n11605), .Z(n353) );
  NAND U812 ( .A(n352), .B(n353), .Z(n11832) );
  XNOR U813 ( .A(n7703), .B(n7702), .Z(n7716) );
  XNOR U814 ( .A(n7913), .B(n7912), .Z(n7914) );
  XNOR U815 ( .A(n8075), .B(n8074), .Z(n8077) );
  XOR U816 ( .A(n8028), .B(n8027), .Z(n8032) );
  XNOR U817 ( .A(n8598), .B(n8597), .Z(n8599) );
  XNOR U818 ( .A(n8581), .B(n8582), .Z(n8573) );
  XNOR U819 ( .A(n8971), .B(n8970), .Z(n8972) );
  XOR U820 ( .A(n8728), .B(n8727), .Z(n8686) );
  XNOR U821 ( .A(n8951), .B(n8950), .Z(n8952) );
  XNOR U822 ( .A(n8872), .B(n8871), .Z(n8874) );
  XOR U823 ( .A(n9055), .B(n9054), .Z(n9115) );
  NAND U824 ( .A(n4747), .B(n4746), .Z(n354) );
  NANDN U825 ( .A(n4749), .B(n4748), .Z(n355) );
  AND U826 ( .A(n354), .B(n355), .Z(n4884) );
  XNOR U827 ( .A(n5003), .B(n5002), .Z(n5005) );
  XNOR U828 ( .A(n5372), .B(n5371), .Z(n5322) );
  XNOR U829 ( .A(n5344), .B(n5343), .Z(n5388) );
  XNOR U830 ( .A(n5382), .B(n5381), .Z(n5384) );
  XNOR U831 ( .A(n5675), .B(n5674), .Z(n5677) );
  XNOR U832 ( .A(n5782), .B(n5781), .Z(n5753) );
  XNOR U833 ( .A(n5908), .B(n5909), .Z(n5890) );
  XNOR U834 ( .A(n6092), .B(n6091), .Z(n6093) );
  XNOR U835 ( .A(n6098), .B(n6097), .Z(n6100) );
  XNOR U836 ( .A(n1394), .B(n1393), .Z(n1387) );
  XNOR U837 ( .A(n1855), .B(n1854), .Z(n1857) );
  XNOR U838 ( .A(n1750), .B(n1749), .Z(n1724) );
  XNOR U839 ( .A(n2555), .B(n2554), .Z(n2611) );
  XNOR U840 ( .A(n3039), .B(n3038), .Z(n3040) );
  XNOR U841 ( .A(n3077), .B(n3076), .Z(n3078) );
  XNOR U842 ( .A(n23595), .B(n23594), .Z(n23596) );
  XNOR U843 ( .A(n23369), .B(n23368), .Z(n23370) );
  XNOR U844 ( .A(n23639), .B(n23638), .Z(n23640) );
  XNOR U845 ( .A(n23588), .B(n23587), .Z(n23589) );
  XNOR U846 ( .A(n23582), .B(n23783), .Z(n23583) );
  NAND U847 ( .A(n18876), .B(n18875), .Z(n356) );
  NAND U848 ( .A(n18874), .B(n18873), .Z(n357) );
  AND U849 ( .A(n356), .B(n357), .Z(n18919) );
  XNOR U850 ( .A(n19067), .B(n19066), .Z(n19069) );
  NAND U851 ( .A(n18924), .B(n18923), .Z(n358) );
  NANDN U852 ( .A(n18926), .B(n18925), .Z(n359) );
  NAND U853 ( .A(n358), .B(n359), .Z(n19056) );
  XOR U854 ( .A(n19488), .B(n19487), .Z(n19397) );
  XNOR U855 ( .A(n19720), .B(n19719), .Z(n19722) );
  XNOR U856 ( .A(n20123), .B(n20122), .Z(n20125) );
  XNOR U857 ( .A(n20056), .B(n20055), .Z(n20057) );
  XNOR U858 ( .A(n20324), .B(n20323), .Z(n20325) );
  XOR U859 ( .A(n20603), .B(n20602), .Z(n20613) );
  XNOR U860 ( .A(n20841), .B(n20840), .Z(n20842) );
  NAND U861 ( .A(n20691), .B(n20690), .Z(n360) );
  NAND U862 ( .A(n20689), .B(n20688), .Z(n361) );
  NAND U863 ( .A(n360), .B(n361), .Z(n20915) );
  XNOR U864 ( .A(n20889), .B(n20888), .Z(n20909) );
  NAND U865 ( .A(n20702), .B(n20701), .Z(n362) );
  NAND U866 ( .A(n20700), .B(n20865), .Z(n363) );
  AND U867 ( .A(n362), .B(n363), .Z(n20922) );
  NAND U868 ( .A(n20930), .B(n20929), .Z(n364) );
  NAND U869 ( .A(n20927), .B(n20928), .Z(n365) );
  NAND U870 ( .A(n364), .B(n365), .Z(n21086) );
  XNOR U871 ( .A(n15827), .B(n15826), .Z(n15828) );
  XOR U872 ( .A(n15973), .B(n15972), .Z(n15955) );
  XNOR U873 ( .A(n16006), .B(n16007), .Z(n15992) );
  XNOR U874 ( .A(n16291), .B(n16290), .Z(n16292) );
  XOR U875 ( .A(n16676), .B(n16675), .Z(n16686) );
  XNOR U876 ( .A(n16821), .B(n16820), .Z(n16822) );
  XNOR U877 ( .A(n17496), .B(n17495), .Z(n17500) );
  NAND U878 ( .A(n17420), .B(n17419), .Z(n366) );
  NANDN U879 ( .A(n17418), .B(n17417), .Z(n367) );
  NAND U880 ( .A(n366), .B(n367), .Z(n17629) );
  NAND U881 ( .A(n17528), .B(n17527), .Z(n368) );
  NAND U882 ( .A(n17526), .B(n17525), .Z(n369) );
  NAND U883 ( .A(n368), .B(n369), .Z(n17757) );
  NAND U884 ( .A(n17552), .B(n17551), .Z(n370) );
  NAND U885 ( .A(n17550), .B(n17549), .Z(n371) );
  AND U886 ( .A(n370), .B(n371), .Z(n17774) );
  XNOR U887 ( .A(n17768), .B(n17767), .Z(n17770) );
  NAND U888 ( .A(n17589), .B(n17588), .Z(n372) );
  NANDN U889 ( .A(n17591), .B(n17590), .Z(n373) );
  AND U890 ( .A(n372), .B(n373), .Z(n17763) );
  NAND U891 ( .A(n17627), .B(n17626), .Z(n374) );
  NANDN U892 ( .A(n17625), .B(n17624), .Z(n375) );
  AND U893 ( .A(n374), .B(n375), .Z(n17658) );
  NAND U894 ( .A(n17691), .B(n17690), .Z(n376) );
  NAND U895 ( .A(n17689), .B(n17688), .Z(n377) );
  NAND U896 ( .A(n376), .B(n377), .Z(n17883) );
  NAND U897 ( .A(n18072), .B(n18071), .Z(n378) );
  NAND U898 ( .A(n18069), .B(n18070), .Z(n379) );
  NAND U899 ( .A(n378), .B(n379), .Z(n18267) );
  XNOR U900 ( .A(n18200), .B(n18199), .Z(n18198) );
  XNOR U901 ( .A(n12915), .B(o[137]), .Z(n12907) );
  XNOR U902 ( .A(n13005), .B(n13004), .Z(n13006) );
  XNOR U903 ( .A(n13154), .B(n13153), .Z(n13156) );
  XNOR U904 ( .A(n13401), .B(n13400), .Z(n13403) );
  XNOR U905 ( .A(n13397), .B(n13396), .Z(n13389) );
  XNOR U906 ( .A(n13703), .B(n13702), .Z(n13704) );
  NAND U907 ( .A(n13937), .B(n13936), .Z(n380) );
  NANDN U908 ( .A(n13939), .B(n13938), .Z(n381) );
  NAND U909 ( .A(n380), .B(n381), .Z(n14077) );
  NAND U910 ( .A(n14135), .B(n14134), .Z(n382) );
  NANDN U911 ( .A(n14137), .B(n14136), .Z(n383) );
  NAND U912 ( .A(n382), .B(n383), .Z(n14328) );
  XNOR U913 ( .A(n14450), .B(n14449), .Z(n14452) );
  NAND U914 ( .A(n14448), .B(n14447), .Z(n384) );
  NAND U915 ( .A(n14446), .B(n14445), .Z(n385) );
  AND U916 ( .A(n384), .B(n385), .Z(n14596) );
  NAND U917 ( .A(n14399), .B(n14398), .Z(n386) );
  NAND U918 ( .A(n14396), .B(n14397), .Z(n387) );
  AND U919 ( .A(n386), .B(n387), .Z(n14591) );
  XNOR U920 ( .A(n15031), .B(n15030), .Z(n15033) );
  XNOR U921 ( .A(n15205), .B(n15204), .Z(n15206) );
  XNOR U922 ( .A(n14914), .B(n14913), .Z(n14773) );
  XOR U923 ( .A(n9933), .B(n10717), .Z(n9935) );
  XNOR U924 ( .A(n10273), .B(n10272), .Z(n10223) );
  XOR U925 ( .A(n10817), .B(n10816), .Z(n10860) );
  XNOR U926 ( .A(n11171), .B(n11170), .Z(n11172) );
  NAND U927 ( .A(n11920), .B(n11919), .Z(n388) );
  NANDN U928 ( .A(n11918), .B(n11917), .Z(n389) );
  NAND U929 ( .A(n388), .B(n389), .Z(n12120) );
  XNOR U930 ( .A(n12452), .B(n12285), .Z(n12286) );
  XNOR U931 ( .A(n12263), .B(n12262), .Z(n12264) );
  XNOR U932 ( .A(n6936), .B(o[70]), .Z(n6928) );
  XNOR U933 ( .A(n7018), .B(n7017), .Z(n7019) );
  XNOR U934 ( .A(n7155), .B(n7154), .Z(n7156) );
  XNOR U935 ( .A(n7249), .B(n7248), .Z(n7242) );
  XNOR U936 ( .A(n7551), .B(n7550), .Z(n7553) );
  XNOR U937 ( .A(n7547), .B(n7546), .Z(n7539) );
  XOR U938 ( .A(n7921), .B(n7920), .Z(n7964) );
  XNOR U939 ( .A(n8000), .B(n7999), .Z(n8094) );
  XNOR U940 ( .A(n8265), .B(n8264), .Z(n8266) );
  XNOR U941 ( .A(n8604), .B(n8603), .Z(n8606) );
  XNOR U942 ( .A(n8539), .B(n8538), .Z(n8540) );
  XNOR U943 ( .A(n8785), .B(n8784), .Z(n8801) );
  XNOR U944 ( .A(n8850), .B(n8849), .Z(n8841) );
  XOR U945 ( .A(n8984), .B(n8983), .Z(n8986) );
  XNOR U946 ( .A(n8990), .B(n8989), .Z(n8992) );
  XNOR U947 ( .A(n9002), .B(n9001), .Z(n9003) );
  XNOR U948 ( .A(n9022), .B(n9021), .Z(n9009) );
  NAND U949 ( .A(n9032), .B(n9031), .Z(n390) );
  NAND U950 ( .A(n9030), .B(n9029), .Z(n391) );
  NAND U951 ( .A(n390), .B(n391), .Z(n9247) );
  XNOR U952 ( .A(n4069), .B(n4068), .Z(n4070) );
  XOR U953 ( .A(n4305), .B(n4306), .Z(n4291) );
  NAND U954 ( .A(n4237), .B(n4236), .Z(n392) );
  NAND U955 ( .A(n4235), .B(n4532), .Z(n393) );
  NAND U956 ( .A(n392), .B(n393), .Z(n4284) );
  XOR U957 ( .A(n5017), .B(n5016), .Z(n4926) );
  XOR U958 ( .A(n5023), .B(n5022), .Z(n5027) );
  XNOR U959 ( .A(n5141), .B(n5140), .Z(n5142) );
  XOR U960 ( .A(n5396), .B(n5395), .Z(n5399) );
  XNOR U961 ( .A(n5706), .B(n5705), .Z(n5708) );
  XNOR U962 ( .A(n5712), .B(n5711), .Z(n5713) );
  XNOR U963 ( .A(n5963), .B(n5962), .Z(n5965) );
  XOR U964 ( .A(n6342), .B(n6341), .Z(n6316) );
  NAND U965 ( .A(n6108), .B(n6107), .Z(n394) );
  NANDN U966 ( .A(n6110), .B(n6109), .Z(n395) );
  AND U967 ( .A(n394), .B(n395), .Z(n6310) );
  XNOR U968 ( .A(n6306), .B(n6305), .Z(n6327) );
  XNOR U969 ( .A(n6265), .B(n6264), .Z(n6267) );
  XNOR U970 ( .A(n6281), .B(o[60]), .Z(n6295) );
  XNOR U971 ( .A(n6684), .B(n6442), .Z(n6443) );
  XOR U972 ( .A(n1154), .B(n1958), .Z(n1156) );
  XNOR U973 ( .A(n1288), .B(n1287), .Z(n1289) );
  NAND U974 ( .A(n2229), .B(n2228), .Z(n396) );
  NANDN U975 ( .A(n2231), .B(n2230), .Z(n397) );
  NAND U976 ( .A(n396), .B(n397), .Z(n2369) );
  NAND U977 ( .A(n2419), .B(n2418), .Z(n398) );
  NANDN U978 ( .A(n2421), .B(n2420), .Z(n399) );
  NAND U979 ( .A(n398), .B(n399), .Z(n2565) );
  NAND U980 ( .A(n3173), .B(n3172), .Z(n400) );
  NANDN U981 ( .A(n3175), .B(n3174), .Z(n401) );
  NAND U982 ( .A(n400), .B(n401), .Z(n3360) );
  XOR U983 ( .A(n21446), .B(n21445), .Z(n21419) );
  XNOR U984 ( .A(n22506), .B(n22505), .Z(n22508) );
  XOR U985 ( .A(n22500), .B(n22499), .Z(n22502) );
  XNOR U986 ( .A(n23492), .B(n23491), .Z(n23362) );
  XNOR U987 ( .A(n23530), .B(n23529), .Z(n23532) );
  XNOR U988 ( .A(n23621), .B(n23620), .Z(n23622) );
  XOR U989 ( .A(n23653), .B(n23652), .Z(n23628) );
  XOR U990 ( .A(n23611), .B(n23610), .Z(n23656) );
  XNOR U991 ( .A(n23524), .B(n23523), .Z(n23525) );
  XNOR U992 ( .A(n23829), .B(n23828), .Z(n23805) );
  XNOR U993 ( .A(n23797), .B(n23796), .Z(n23798) );
  XNOR U994 ( .A(n23766), .B(n23765), .Z(n23820) );
  XOR U995 ( .A(n23833), .B(n23832), .Z(n23835) );
  XNOR U996 ( .A(n24092), .B(n24091), .Z(n24090) );
  XNOR U997 ( .A(n23912), .B(n23911), .Z(n23909) );
  XNOR U998 ( .A(n18527), .B(n18526), .Z(n18534) );
  XNOR U999 ( .A(n19494), .B(n19493), .Z(n19497) );
  XNOR U1000 ( .A(n20345), .B(n20344), .Z(n20339) );
  XNOR U1001 ( .A(n20627), .B(n20626), .Z(n20499) );
  XNOR U1002 ( .A(n20749), .B(n20748), .Z(n20751) );
  XNOR U1003 ( .A(n20767), .B(n20766), .Z(n20768) );
  XOR U1004 ( .A(n20996), .B(n20926), .Z(n402) );
  NANDN U1005 ( .A(n20925), .B(n402), .Z(n403) );
  NAND U1006 ( .A(n20996), .B(n20926), .Z(n404) );
  AND U1007 ( .A(n403), .B(n404), .Z(n21135) );
  NAND U1008 ( .A(n20886), .B(n20885), .Z(n405) );
  NAND U1009 ( .A(n20884), .B(n20986), .Z(n406) );
  NAND U1010 ( .A(n405), .B(n406), .Z(n20979) );
  XNOR U1011 ( .A(n20965), .B(n20964), .Z(n20962) );
  XNOR U1012 ( .A(n15670), .B(n15669), .Z(n15672) );
  XNOR U1013 ( .A(n15978), .B(n15977), .Z(n15979) );
  XOR U1014 ( .A(n16037), .B(n16036), .Z(n16048) );
  XNOR U1015 ( .A(n16706), .B(n16705), .Z(n16709) );
  XOR U1016 ( .A(n16955), .B(n16954), .Z(n16850) );
  NAND U1017 ( .A(n17874), .B(n17873), .Z(n407) );
  NAND U1018 ( .A(n17872), .B(n17871), .Z(n408) );
  NAND U1019 ( .A(n407), .B(n408), .Z(n17990) );
  XNOR U1020 ( .A(n17821), .B(n17820), .Z(n17815) );
  AND U1021 ( .A(n17728), .B(n17727), .Z(n409) );
  AND U1022 ( .A(n18157), .B(y[1955]), .Z(n410) );
  NAND U1023 ( .A(x[244]), .B(n410), .Z(n411) );
  NANDN U1024 ( .A(n409), .B(n411), .Z(n17917) );
  NAND U1025 ( .A(n17732), .B(n17731), .Z(n412) );
  NAND U1026 ( .A(n17730), .B(n17729), .Z(n413) );
  NAND U1027 ( .A(n412), .B(n413), .Z(n17913) );
  NAND U1028 ( .A(n18023), .B(n18022), .Z(n414) );
  NAND U1029 ( .A(n18020), .B(n18021), .Z(n415) );
  NAND U1030 ( .A(n414), .B(n415), .Z(n18114) );
  XNOR U1031 ( .A(n13831), .B(n13830), .Z(n13832) );
  XNOR U1032 ( .A(n14478), .B(n14477), .Z(n14480) );
  XNOR U1033 ( .A(n15134), .B(n15133), .Z(n15139) );
  XNOR U1034 ( .A(n15385), .B(n15384), .Z(n15382) );
  XNOR U1035 ( .A(n15316), .B(n15154), .Z(n15155) );
  XOR U1036 ( .A(n15306), .B(n15305), .Z(n15304) );
  XNOR U1037 ( .A(n14946), .B(n14945), .Z(n14947) );
  NAND U1038 ( .A(n9982), .B(n9981), .Z(n416) );
  NANDN U1039 ( .A(n9984), .B(n9983), .Z(n417) );
  AND U1040 ( .A(n416), .B(n417), .Z(n10020) );
  XNOR U1041 ( .A(n10291), .B(n10290), .Z(n10292) );
  NAND U1042 ( .A(n10520), .B(n10519), .Z(n418) );
  NANDN U1043 ( .A(n10518), .B(n10517), .Z(n419) );
  AND U1044 ( .A(n418), .B(n419), .Z(n10568) );
  XOR U1045 ( .A(n11035), .B(n11034), .Z(n11028) );
  XNOR U1046 ( .A(n12151), .B(n12150), .Z(n12152) );
  XNOR U1047 ( .A(n12235), .B(n12234), .Z(n12240) );
  XOR U1048 ( .A(n12195), .B(n12194), .Z(n12042) );
  XNOR U1049 ( .A(n7978), .B(n7977), .Z(n7981) );
  XOR U1050 ( .A(n8230), .B(n8229), .Z(n8125) );
  XOR U1051 ( .A(n9155), .B(n9154), .Z(n9141) );
  NAND U1052 ( .A(n9380), .B(n9379), .Z(n420) );
  NAND U1053 ( .A(n9378), .B(n9646), .Z(n421) );
  NAND U1054 ( .A(n420), .B(n421), .Z(n9506) );
  XNOR U1055 ( .A(n4147), .B(n4146), .Z(n4148) );
  XNOR U1056 ( .A(n4155), .B(n4154), .Z(n4206) );
  XOR U1057 ( .A(n5535), .B(n5534), .Z(n5421) );
  XNOR U1058 ( .A(n6033), .B(n6032), .Z(n6035) );
  XNOR U1059 ( .A(n6478), .B(n6477), .Z(n6371) );
  XNOR U1060 ( .A(n6386), .B(n6385), .Z(n6378) );
  XNOR U1061 ( .A(n6756), .B(n6755), .Z(n6754) );
  XNOR U1062 ( .A(n6644), .B(n6643), .Z(n6641) );
  XOR U1063 ( .A(n6500), .B(n6499), .Z(n6501) );
  NAND U1064 ( .A(n1238), .B(n1237), .Z(n422) );
  NANDN U1065 ( .A(n1869), .B(n1578), .Z(n423) );
  AND U1066 ( .A(n422), .B(n423), .Z(n1241) );
  NAND U1067 ( .A(n2500), .B(n2499), .Z(n424) );
  NANDN U1068 ( .A(n2502), .B(n2501), .Z(n425) );
  AND U1069 ( .A(n424), .B(n425), .Z(n2505) );
  XOR U1070 ( .A(n3252), .B(n3251), .Z(n3246) );
  XNOR U1071 ( .A(n21281), .B(n21280), .Z(n21282) );
  XNOR U1072 ( .A(n21744), .B(n21743), .Z(n21746) );
  XNOR U1073 ( .A(n21753), .B(n21752), .Z(n21834) );
  XNOR U1074 ( .A(n22359), .B(n22358), .Z(n22362) );
  XNOR U1075 ( .A(n23038), .B(n23037), .Z(n23039) );
  XNOR U1076 ( .A(n23874), .B(n23873), .Z(n23872) );
  XNOR U1077 ( .A(n23811), .B(n23810), .Z(n23705) );
  XNOR U1078 ( .A(n23886), .B(n23885), .Z(n23883) );
  XOR U1079 ( .A(n18698), .B(n18697), .Z(n18700) );
  XNOR U1080 ( .A(n19181), .B(n19180), .Z(n19183) );
  XNOR U1081 ( .A(n19759), .B(n19758), .Z(n19761) );
  XNOR U1082 ( .A(n20030), .B(n20029), .Z(n20032) );
  NAND U1083 ( .A(n20899), .B(n20898), .Z(n426) );
  NAND U1084 ( .A(n20897), .B(n20896), .Z(n427) );
  NAND U1085 ( .A(n426), .B(n427), .Z(n21179) );
  NAND U1086 ( .A(n20823), .B(n20822), .Z(n428) );
  NANDN U1087 ( .A(n20825), .B(n20824), .Z(n429) );
  AND U1088 ( .A(n428), .B(n429), .Z(n21170) );
  NAND U1089 ( .A(n20908), .B(n20907), .Z(n430) );
  NAND U1090 ( .A(n20906), .B(n20905), .Z(n431) );
  AND U1091 ( .A(n430), .B(n431), .Z(n21153) );
  XOR U1092 ( .A(n15721), .B(n15643), .Z(n432) );
  NANDN U1093 ( .A(n15644), .B(n432), .Z(n433) );
  NAND U1094 ( .A(n15721), .B(n15643), .Z(n434) );
  AND U1095 ( .A(n433), .B(n434), .Z(n15701) );
  XNOR U1096 ( .A(n15735), .B(n15734), .Z(n15739) );
  XOR U1097 ( .A(n15902), .B(n15901), .Z(n15904) );
  XNOR U1098 ( .A(n16315), .B(n16314), .Z(n16398) );
  OR U1099 ( .A(n16501), .B(n16502), .Z(n435) );
  NAND U1100 ( .A(n16499), .B(n16500), .Z(n436) );
  NAND U1101 ( .A(n435), .B(n436), .Z(n16720) );
  XNOR U1102 ( .A(n16975), .B(n16974), .Z(n16976) );
  XNOR U1103 ( .A(n17787), .B(n17786), .Z(n17788) );
  NAND U1104 ( .A(n17910), .B(n17909), .Z(n437) );
  NAND U1105 ( .A(n17908), .B(n17907), .Z(n438) );
  NAND U1106 ( .A(n437), .B(n438), .Z(n18039) );
  NAND U1107 ( .A(n18045), .B(n18044), .Z(n439) );
  NAND U1108 ( .A(n18043), .B(n18042), .Z(n440) );
  NAND U1109 ( .A(n439), .B(n440), .Z(n18317) );
  XOR U1110 ( .A(n18300), .B(n18299), .Z(n18298) );
  XNOR U1111 ( .A(n13147), .B(n13146), .Z(n13149) );
  XNOR U1112 ( .A(n13421), .B(n13420), .Z(n13422) );
  XOR U1113 ( .A(n14602), .B(n14601), .Z(n14604) );
  XNOR U1114 ( .A(n14930), .B(n14929), .Z(n15089) );
  XOR U1115 ( .A(n15219), .B(n15218), .Z(n15114) );
  XNOR U1116 ( .A(n15270), .B(n15269), .Z(n15229) );
  XNOR U1117 ( .A(n15294), .B(n15293), .Z(n15291) );
  XNOR U1118 ( .A(n10365), .B(n10364), .Z(n10367) );
  XNOR U1119 ( .A(n11156), .B(n11155), .Z(n11157) );
  XNOR U1120 ( .A(n12371), .B(n12370), .Z(n12330) );
  XNOR U1121 ( .A(n12387), .B(n12386), .Z(n12619) );
  XNOR U1122 ( .A(n7297), .B(n7296), .Z(n7299) );
  XNOR U1123 ( .A(n7567), .B(n7566), .Z(n7568) );
  XNOR U1124 ( .A(n8250), .B(n8249), .Z(n8251) );
  XNOR U1125 ( .A(n8827), .B(n8826), .Z(n8829) );
  XNOR U1126 ( .A(n9420), .B(n9419), .Z(n9338) );
  XNOR U1127 ( .A(n9331), .B(n9330), .Z(n9333) );
  XNOR U1128 ( .A(n9325), .B(n9324), .Z(n9327) );
  NAND U1129 ( .A(n9416), .B(n9415), .Z(n441) );
  NAND U1130 ( .A(n9414), .B(n9413), .Z(n442) );
  AND U1131 ( .A(n441), .B(n442), .Z(n9710) );
  NAND U1132 ( .A(n9430), .B(n9429), .Z(n443) );
  NAND U1133 ( .A(n9428), .B(n9427), .Z(n444) );
  AND U1134 ( .A(n443), .B(n444), .Z(n9692) );
  XOR U1135 ( .A(n9564), .B(n9449), .Z(n445) );
  XNOR U1136 ( .A(n9450), .B(n445), .Z(n9369) );
  XOR U1137 ( .A(n9724), .B(n9723), .Z(n9722) );
  XOR U1138 ( .A(n4106), .B(n4105), .Z(n4092) );
  XNOR U1139 ( .A(n4609), .B(n4608), .Z(n4610) );
  XOR U1140 ( .A(n4715), .B(n4714), .Z(n4797) );
  XNOR U1141 ( .A(n5565), .B(n5564), .Z(n5566) );
  XNOR U1142 ( .A(n6760), .B(n6759), .Z(n6774) );
  XOR U1143 ( .A(n1166), .B(n1165), .Z(n1183) );
  XNOR U1144 ( .A(n1190), .B(n1189), .Z(n1192) );
  XNOR U1145 ( .A(n1616), .B(n1615), .Z(n1618) );
  XNOR U1146 ( .A(n1913), .B(n1912), .Z(n2012) );
  XOR U1147 ( .A(n3840), .B(n3839), .Z(n3838) );
  XNOR U1148 ( .A(n3602), .B(n3601), .Z(n3598) );
  XNOR U1149 ( .A(n3555), .B(n3554), .Z(n3556) );
  NAND U1150 ( .A(n21258), .B(n21257), .Z(n446) );
  XOR U1151 ( .A(n21258), .B(n21257), .Z(n447) );
  NANDN U1152 ( .A(n21259), .B(n447), .Z(n448) );
  NAND U1153 ( .A(n446), .B(n448), .Z(n21278) );
  NAND U1154 ( .A(n21408), .B(n21409), .Z(n449) );
  XOR U1155 ( .A(n21408), .B(n21409), .Z(n450) );
  NANDN U1156 ( .A(n21407), .B(n450), .Z(n451) );
  NAND U1157 ( .A(n449), .B(n451), .Z(n21459) );
  NAND U1158 ( .A(n21607), .B(n21608), .Z(n452) );
  XOR U1159 ( .A(n21607), .B(n21608), .Z(n453) );
  NANDN U1160 ( .A(n21606), .B(n453), .Z(n454) );
  NAND U1161 ( .A(n452), .B(n454), .Z(n21740) );
  XOR U1162 ( .A(n22245), .B(n22246), .Z(n455) );
  NANDN U1163 ( .A(n22247), .B(n455), .Z(n456) );
  NAND U1164 ( .A(n22245), .B(n22246), .Z(n457) );
  AND U1165 ( .A(n456), .B(n457), .Z(n22369) );
  XNOR U1166 ( .A(n22495), .B(n22494), .Z(n22491) );
  NAND U1167 ( .A(n22894), .B(n22895), .Z(n458) );
  XOR U1168 ( .A(n22894), .B(n22895), .Z(n459) );
  NANDN U1169 ( .A(n22893), .B(n459), .Z(n460) );
  NAND U1170 ( .A(n458), .B(n460), .Z(n23034) );
  XOR U1171 ( .A(n23686), .B(n23685), .Z(n461) );
  NANDN U1172 ( .A(n23684), .B(n461), .Z(n462) );
  NAND U1173 ( .A(n23686), .B(n23685), .Z(n463) );
  AND U1174 ( .A(n462), .B(n463), .Z(n24146) );
  NAND U1175 ( .A(n18397), .B(n18396), .Z(n464) );
  NAND U1176 ( .A(n18505), .B(n18395), .Z(n465) );
  NAND U1177 ( .A(n464), .B(n465), .Z(n18418) );
  NAND U1178 ( .A(n18639), .B(n18640), .Z(n466) );
  XOR U1179 ( .A(n18639), .B(n18640), .Z(n467) );
  NANDN U1180 ( .A(n18638), .B(n467), .Z(n468) );
  NAND U1181 ( .A(n466), .B(n468), .Z(n18694) );
  XOR U1182 ( .A(n18852), .B(n18853), .Z(n469) );
  NANDN U1183 ( .A(n18854), .B(n469), .Z(n470) );
  NAND U1184 ( .A(n18852), .B(n18853), .Z(n471) );
  AND U1185 ( .A(n470), .B(n471), .Z(n18985) );
  NAND U1186 ( .A(n19089), .B(n19090), .Z(n472) );
  XOR U1187 ( .A(n19089), .B(n19090), .Z(n473) );
  NANDN U1188 ( .A(n19088), .B(n473), .Z(n474) );
  NAND U1189 ( .A(n472), .B(n474), .Z(n19186) );
  XOR U1190 ( .A(n19503), .B(n19504), .Z(n475) );
  NANDN U1191 ( .A(n19505), .B(n475), .Z(n476) );
  NAND U1192 ( .A(n19503), .B(n19504), .Z(n477) );
  AND U1193 ( .A(n476), .B(n477), .Z(n19627) );
  XOR U1194 ( .A(n20191), .B(n20192), .Z(n478) );
  NANDN U1195 ( .A(n20193), .B(n478), .Z(n479) );
  NAND U1196 ( .A(n20191), .B(n20192), .Z(n480) );
  AND U1197 ( .A(n479), .B(n480), .Z(n20485) );
  NAND U1198 ( .A(n20647), .B(n20648), .Z(n481) );
  XOR U1199 ( .A(n20647), .B(n20648), .Z(n482) );
  NANDN U1200 ( .A(n20646), .B(n482), .Z(n483) );
  NAND U1201 ( .A(n481), .B(n483), .Z(n20781) );
  XNOR U1202 ( .A(n20942), .B(n20943), .Z(n20941) );
  NAND U1203 ( .A(n15607), .B(n15606), .Z(n484) );
  NAND U1204 ( .A(n15713), .B(n15605), .Z(n485) );
  NAND U1205 ( .A(n484), .B(n485), .Z(n15629) );
  NAND U1206 ( .A(n15843), .B(n15844), .Z(n486) );
  XOR U1207 ( .A(n15843), .B(n15844), .Z(n487) );
  NANDN U1208 ( .A(n15842), .B(n487), .Z(n488) );
  NAND U1209 ( .A(n486), .B(n488), .Z(n15898) );
  NAND U1210 ( .A(n16309), .B(n16310), .Z(n489) );
  XOR U1211 ( .A(n16309), .B(n16310), .Z(n490) );
  NANDN U1212 ( .A(n16308), .B(n490), .Z(n491) );
  NAND U1213 ( .A(n489), .B(n491), .Z(n16393) );
  XOR U1214 ( .A(n16598), .B(n16597), .Z(n492) );
  NANDN U1215 ( .A(n16599), .B(n492), .Z(n493) );
  NAND U1216 ( .A(n16598), .B(n16597), .Z(n494) );
  AND U1217 ( .A(n493), .B(n494), .Z(n16716) );
  XOR U1218 ( .A(n16964), .B(n16965), .Z(n495) );
  NANDN U1219 ( .A(n16966), .B(n495), .Z(n496) );
  NAND U1220 ( .A(n16964), .B(n16965), .Z(n497) );
  AND U1221 ( .A(n496), .B(n497), .Z(n16981) );
  XOR U1222 ( .A(n17638), .B(n17639), .Z(n498) );
  NANDN U1223 ( .A(n17640), .B(n498), .Z(n499) );
  NAND U1224 ( .A(n17638), .B(n17639), .Z(n500) );
  AND U1225 ( .A(n499), .B(n500), .Z(n17780) );
  NAND U1226 ( .A(n17796), .B(n17795), .Z(n501) );
  NAND U1227 ( .A(n17793), .B(n17794), .Z(n502) );
  AND U1228 ( .A(n501), .B(n502), .Z(n17927) );
  NAND U1229 ( .A(n17962), .B(n17961), .Z(n503) );
  NANDN U1230 ( .A(n17960), .B(n17959), .Z(n504) );
  AND U1231 ( .A(n503), .B(n504), .Z(n18334) );
  NANDN U1232 ( .A(n12738), .B(n12740), .Z(n505) );
  OR U1233 ( .A(n12740), .B(n12741), .Z(n506) );
  NAND U1234 ( .A(n12739), .B(n506), .Z(n507) );
  NAND U1235 ( .A(n505), .B(n507), .Z(n12759) );
  NAND U1236 ( .A(n12814), .B(n12815), .Z(n508) );
  XOR U1237 ( .A(n12814), .B(n12815), .Z(n509) );
  NANDN U1238 ( .A(n12813), .B(n509), .Z(n510) );
  NAND U1239 ( .A(n508), .B(n510), .Z(n12855) );
  XOR U1240 ( .A(n12955), .B(n12956), .Z(n511) );
  NANDN U1241 ( .A(n12957), .B(n511), .Z(n512) );
  NAND U1242 ( .A(n12955), .B(n12956), .Z(n513) );
  AND U1243 ( .A(n512), .B(n513), .Z(n13073) );
  NAND U1244 ( .A(n13733), .B(n13734), .Z(n514) );
  XOR U1245 ( .A(n13733), .B(n13734), .Z(n515) );
  NANDN U1246 ( .A(n13732), .B(n515), .Z(n516) );
  NAND U1247 ( .A(n514), .B(n516), .Z(n13842) );
  NAND U1248 ( .A(n14090), .B(n14091), .Z(n517) );
  XOR U1249 ( .A(n14090), .B(n14091), .Z(n518) );
  NANDN U1250 ( .A(n14089), .B(n518), .Z(n519) );
  NAND U1251 ( .A(n517), .B(n519), .Z(n14099) );
  NAND U1252 ( .A(n14468), .B(n14469), .Z(n520) );
  XOR U1253 ( .A(n14468), .B(n14469), .Z(n521) );
  NANDN U1254 ( .A(n14467), .B(n521), .Z(n522) );
  NAND U1255 ( .A(n520), .B(n522), .Z(n14598) );
  XOR U1256 ( .A(n14917), .B(n14918), .Z(n523) );
  NANDN U1257 ( .A(n14919), .B(n523), .Z(n524) );
  NAND U1258 ( .A(n14917), .B(n14918), .Z(n525) );
  AND U1259 ( .A(n524), .B(n525), .Z(n15084) );
  NANDN U1260 ( .A(n15548), .B(n15547), .Z(n15552) );
  NAND U1261 ( .A(n9769), .B(n9768), .Z(n526) );
  XOR U1262 ( .A(n9769), .B(n9768), .Z(n527) );
  NANDN U1263 ( .A(n9770), .B(n527), .Z(n528) );
  NAND U1264 ( .A(n526), .B(n528), .Z(n9787) );
  XOR U1265 ( .A(n10201), .B(n10202), .Z(n529) );
  NANDN U1266 ( .A(n10203), .B(n529), .Z(n530) );
  NAND U1267 ( .A(n10201), .B(n10202), .Z(n531) );
  AND U1268 ( .A(n530), .B(n531), .Z(n10277) );
  XOR U1269 ( .A(n10665), .B(n10666), .Z(n532) );
  NANDN U1270 ( .A(n10667), .B(n532), .Z(n533) );
  NAND U1271 ( .A(n10665), .B(n10666), .Z(n534) );
  AND U1272 ( .A(n533), .B(n534), .Z(n10772) );
  XOR U1273 ( .A(n11016), .B(n11017), .Z(n535) );
  NANDN U1274 ( .A(n11018), .B(n535), .Z(n536) );
  NAND U1275 ( .A(n11016), .B(n11017), .Z(n537) );
  AND U1276 ( .A(n536), .B(n537), .Z(n11143) );
  XOR U1277 ( .A(n12038), .B(n12039), .Z(n538) );
  NANDN U1278 ( .A(n12040), .B(n538), .Z(n539) );
  NAND U1279 ( .A(n12038), .B(n12039), .Z(n540) );
  AND U1280 ( .A(n539), .B(n540), .Z(n12199) );
  XNOR U1281 ( .A(n12662), .B(n12663), .Z(n12660) );
  NAND U1282 ( .A(n6857), .B(n6856), .Z(n541) );
  NAND U1283 ( .A(n6966), .B(n6855), .Z(n542) );
  NAND U1284 ( .A(n541), .B(n542), .Z(n6883) );
  XOR U1285 ( .A(n6937), .B(n6938), .Z(n543) );
  NANDN U1286 ( .A(n6939), .B(n543), .Z(n544) );
  NAND U1287 ( .A(n6937), .B(n6938), .Z(n545) );
  AND U1288 ( .A(n544), .B(n545), .Z(n6954) );
  XNOR U1289 ( .A(n7035), .B(n7034), .Z(n7031) );
  NAND U1290 ( .A(n7876), .B(n7877), .Z(n546) );
  XOR U1291 ( .A(n7876), .B(n7877), .Z(n547) );
  NANDN U1292 ( .A(n7875), .B(n547), .Z(n548) );
  NAND U1293 ( .A(n546), .B(n548), .Z(n7987) );
  XOR U1294 ( .A(n8239), .B(n8240), .Z(n549) );
  NANDN U1295 ( .A(n8241), .B(n549), .Z(n550) );
  NAND U1296 ( .A(n8239), .B(n8240), .Z(n551) );
  AND U1297 ( .A(n550), .B(n551), .Z(n8256) );
  XNOR U1298 ( .A(n9718), .B(n9717), .Z(n9716) );
  XNOR U1299 ( .A(n9471), .B(n9472), .Z(n9470) );
  NAND U1300 ( .A(n3903), .B(n3902), .Z(n552) );
  NAND U1301 ( .A(n4018), .B(n3901), .Z(n553) );
  NAND U1302 ( .A(n552), .B(n553), .Z(n3925) );
  XOR U1303 ( .A(n3989), .B(n3990), .Z(n554) );
  NANDN U1304 ( .A(n3991), .B(n554), .Z(n555) );
  NAND U1305 ( .A(n3989), .B(n3990), .Z(n556) );
  AND U1306 ( .A(n555), .B(n556), .Z(n4006) );
  XNOR U1307 ( .A(n4086), .B(n4085), .Z(n4082) );
  XOR U1308 ( .A(n4598), .B(n4599), .Z(n557) );
  NANDN U1309 ( .A(n4600), .B(n557), .Z(n558) );
  NAND U1310 ( .A(n4598), .B(n4599), .Z(n559) );
  AND U1311 ( .A(n558), .B(n559), .Z(n4615) );
  XOR U1312 ( .A(n4918), .B(n4919), .Z(n560) );
  NANDN U1313 ( .A(n4920), .B(n560), .Z(n561) );
  NAND U1314 ( .A(n4918), .B(n4919), .Z(n562) );
  AND U1315 ( .A(n561), .B(n562), .Z(n5147) );
  XNOR U1316 ( .A(n6790), .B(n6789), .Z(n6814) );
  XNOR U1317 ( .A(n1060), .B(n1059), .Z(n1056) );
  XOR U1318 ( .A(n1131), .B(n1130), .Z(n563) );
  NANDN U1319 ( .A(n1132), .B(n563), .Z(n564) );
  NAND U1320 ( .A(n1131), .B(n1130), .Z(n565) );
  AND U1321 ( .A(n564), .B(n565), .Z(n1176) );
  XOR U1322 ( .A(n1605), .B(n1606), .Z(n566) );
  NANDN U1323 ( .A(n1607), .B(n566), .Z(n567) );
  NAND U1324 ( .A(n1605), .B(n1606), .Z(n568) );
  AND U1325 ( .A(n567), .B(n568), .Z(n1622) );
  XOR U1326 ( .A(n1900), .B(n1901), .Z(n569) );
  NANDN U1327 ( .A(n1902), .B(n569), .Z(n570) );
  NAND U1328 ( .A(n1900), .B(n1901), .Z(n571) );
  AND U1329 ( .A(n570), .B(n571), .Z(n2019) );
  NAND U1330 ( .A(n2642), .B(n2643), .Z(n572) );
  XOR U1331 ( .A(n2642), .B(n2643), .Z(n573) );
  NANDN U1332 ( .A(n2641), .B(n573), .Z(n574) );
  NAND U1333 ( .A(n572), .B(n574), .Z(n2782) );
  XOR U1334 ( .A(n3090), .B(n3089), .Z(n575) );
  NANDN U1335 ( .A(n3088), .B(n575), .Z(n576) );
  NAND U1336 ( .A(n3090), .B(n3089), .Z(n577) );
  AND U1337 ( .A(n576), .B(n577), .Z(n3099) );
  XNOR U1338 ( .A(n3594), .B(n3593), .Z(n3592) );
  XNOR U1339 ( .A(n23156), .B(n23318), .Z(n23006) );
  XNOR U1340 ( .A(n16645), .B(n16644), .Z(n16647) );
  XNOR U1341 ( .A(n17295), .B(o[184]), .Z(n17304) );
  XNOR U1342 ( .A(n10831), .B(n10830), .Z(n10833) );
  XNOR U1343 ( .A(n7890), .B(n7889), .Z(n7892) );
  XNOR U1344 ( .A(n8586), .B(n8585), .Z(n8588) );
  XNOR U1345 ( .A(n8405), .B(n8404), .Z(n8407) );
  XNOR U1346 ( .A(n8569), .B(n8568), .Z(n8621) );
  XNOR U1347 ( .A(n8763), .B(o[89]), .Z(n8734) );
  XNOR U1348 ( .A(n5220), .B(n5219), .Z(n5222) );
  XNOR U1349 ( .A(n5353), .B(n5352), .Z(n5355) );
  XNOR U1350 ( .A(n22721), .B(n22720), .Z(n22684) );
  XNOR U1351 ( .A(n22702), .B(n22701), .Z(n22658) );
  XNOR U1352 ( .A(n22784), .B(n22783), .Z(n22821) );
  XNOR U1353 ( .A(n22922), .B(n22921), .Z(n22916) );
  XNOR U1354 ( .A(n23158), .B(n23157), .Z(n23173) );
  XNOR U1355 ( .A(n23128), .B(n23127), .Z(n23167) );
  XNOR U1356 ( .A(n19416), .B(n19415), .Z(n19441) );
  XNOR U1357 ( .A(n19465), .B(n19464), .Z(n19403) );
  XNOR U1358 ( .A(n19827), .B(n19826), .Z(n19829) );
  XNOR U1359 ( .A(n19852), .B(n19851), .Z(n19815) );
  XNOR U1360 ( .A(n19833), .B(n19832), .Z(n19789) );
  XNOR U1361 ( .A(n19804), .B(n19803), .Z(n19783) );
  XNOR U1362 ( .A(n19924), .B(n19923), .Z(n19926) );
  XNOR U1363 ( .A(n19958), .B(n19957), .Z(n19960) );
  XNOR U1364 ( .A(n20213), .B(n20212), .Z(n20214) );
  XNOR U1365 ( .A(n20257), .B(n20256), .Z(n20258) );
  XOR U1366 ( .A(n20221), .B(n20220), .Z(n20225) );
  XNOR U1367 ( .A(n20231), .B(n20230), .Z(n20233) );
  XNOR U1368 ( .A(n16641), .B(n16791), .Z(n16613) );
  XNOR U1369 ( .A(n17076), .B(n17075), .Z(n17039) );
  XNOR U1370 ( .A(n17164), .B(n17163), .Z(n17165) );
  XNOR U1371 ( .A(n17138), .B(n17137), .Z(n17200) );
  XNOR U1372 ( .A(n17444), .B(n17443), .Z(n17446) );
  XNOR U1373 ( .A(n14042), .B(n14041), .Z(n13987) );
  NAND U1374 ( .A(n13923), .B(n13922), .Z(n578) );
  NANDN U1375 ( .A(n13921), .B(n13920), .Z(n579) );
  NAND U1376 ( .A(n578), .B(n579), .Z(n14057) );
  XNOR U1377 ( .A(n10827), .B(n10975), .Z(n10787) );
  XNOR U1378 ( .A(n11255), .B(n11254), .Z(n11218) );
  NAND U1379 ( .A(n11212), .B(n11213), .Z(n580) );
  NAND U1380 ( .A(n11214), .B(n11215), .Z(n581) );
  NAND U1381 ( .A(n580), .B(n581), .Z(n11335) );
  XNOR U1382 ( .A(n8348), .B(o[86]), .Z(n8327) );
  XNOR U1383 ( .A(n8351), .B(n8350), .Z(n8314) );
  XNOR U1384 ( .A(n8439), .B(n8438), .Z(n8441) );
  XNOR U1385 ( .A(n8411), .B(n8410), .Z(n8413) );
  XNOR U1386 ( .A(n8387), .B(n8386), .Z(n8474) );
  XNOR U1387 ( .A(n8708), .B(n8707), .Z(n8710) );
  XNOR U1388 ( .A(n8642), .B(n8641), .Z(n8617) );
  XOR U1389 ( .A(n8791), .B(n8790), .Z(n8714) );
  XNOR U1390 ( .A(n8953), .B(n8952), .Z(n8914) );
  XNOR U1391 ( .A(n8867), .B(n8868), .Z(n8908) );
  XNOR U1392 ( .A(n8902), .B(n8901), .Z(n8903) );
  XNOR U1393 ( .A(n8896), .B(n8895), .Z(n8898) );
  XNOR U1394 ( .A(n4982), .B(n4981), .Z(n4932) );
  XNOR U1395 ( .A(n5370), .B(n5369), .Z(n5371) );
  XNOR U1396 ( .A(n5230), .B(n5439), .Z(n5177) );
  XNOR U1397 ( .A(n5181), .B(n5180), .Z(n5192) );
  XNOR U1398 ( .A(n5639), .B(n5638), .Z(n5633) );
  XNOR U1399 ( .A(n5768), .B(n5767), .Z(n5769) );
  XNOR U1400 ( .A(n1748), .B(n1747), .Z(n1749) );
  XNOR U1401 ( .A(n1849), .B(n1848), .Z(n1850) );
  NAND U1402 ( .A(n2215), .B(n2214), .Z(n582) );
  NANDN U1403 ( .A(n2213), .B(n2212), .Z(n583) );
  NAND U1404 ( .A(n582), .B(n583), .Z(n2355) );
  XNOR U1405 ( .A(n2688), .B(n2687), .Z(n2741) );
  XNOR U1406 ( .A(n2675), .B(n2676), .Z(n2765) );
  XNOR U1407 ( .A(n21616), .B(n21615), .Z(n21618) );
  XOR U1408 ( .A(n21638), .B(n21639), .Z(n21623) );
  XNOR U1409 ( .A(n22858), .B(n22857), .Z(n22860) );
  XNOR U1410 ( .A(n22848), .B(n22847), .Z(n22805) );
  XNOR U1411 ( .A(n23134), .B(n23133), .Z(n23104) );
  NAND U1412 ( .A(n18826), .B(n18825), .Z(n584) );
  NANDN U1413 ( .A(n19245), .B(n18879), .Z(n585) );
  NAND U1414 ( .A(n584), .B(n585), .Z(n18875) );
  XNOR U1415 ( .A(n19254), .B(n19253), .Z(n19231) );
  XNOR U1416 ( .A(n19202), .B(n19201), .Z(n19225) );
  XNOR U1417 ( .A(n19216), .B(n19215), .Z(n19218) );
  XNOR U1418 ( .A(n19429), .B(n19428), .Z(n19435) );
  XNOR U1419 ( .A(n19554), .B(n19553), .Z(n19556) );
  XNOR U1420 ( .A(n19591), .B(n19590), .Z(n19593) );
  XNOR U1421 ( .A(n19906), .B(n19905), .Z(n19993) );
  XNOR U1422 ( .A(n20166), .B(n20165), .Z(n20137) );
  XNOR U1423 ( .A(n20105), .B(n20104), .Z(n20107) );
  XNOR U1424 ( .A(n20160), .B(n20159), .Z(n20111) );
  XNOR U1425 ( .A(n20243), .B(n20242), .Z(n20245) );
  XNOR U1426 ( .A(n20237), .B(n20236), .Z(n20238) );
  XOR U1427 ( .A(n20391), .B(n20390), .Z(n20393) );
  XNOR U1428 ( .A(n16430), .B(n16429), .Z(n16431) );
  XOR U1429 ( .A(n16555), .B(n16554), .Z(n16516) );
  XNOR U1430 ( .A(n16634), .B(n16633), .Z(n16673) );
  XOR U1431 ( .A(n16750), .B(n16749), .Z(n16804) );
  XNOR U1432 ( .A(n16811), .B(n16810), .Z(n16765) );
  XNOR U1433 ( .A(n17057), .B(n17056), .Z(n17013) );
  AND U1434 ( .A(n17461), .B(o[185]), .Z(n17609) );
  NAND U1435 ( .A(n17408), .B(n17407), .Z(n586) );
  NAND U1436 ( .A(n17405), .B(n17406), .Z(n587) );
  AND U1437 ( .A(n586), .B(n587), .Z(n17565) );
  AND U1438 ( .A(n17617), .B(o[186]), .Z(n17708) );
  XNOR U1439 ( .A(n13087), .B(n13086), .Z(n13089) );
  XOR U1440 ( .A(n13109), .B(n13110), .Z(n13094) );
  NAND U1441 ( .A(n13783), .B(n13782), .Z(n588) );
  NANDN U1442 ( .A(n13781), .B(n13780), .Z(n589) );
  AND U1443 ( .A(n588), .B(n589), .Z(n13878) );
  AND U1444 ( .A(n13870), .B(n13869), .Z(n590) );
  AND U1445 ( .A(n15313), .B(y[1929]), .Z(n591) );
  NAND U1446 ( .A(x[225]), .B(n591), .Z(n592) );
  NANDN U1447 ( .A(n590), .B(n592), .Z(n14051) );
  NAND U1448 ( .A(n14064), .B(n14063), .Z(n593) );
  NANDN U1449 ( .A(n14066), .B(n14065), .Z(n594) );
  NAND U1450 ( .A(n593), .B(n594), .Z(n14114) );
  NAND U1451 ( .A(n14153), .B(n14152), .Z(n595) );
  NANDN U1452 ( .A(n14155), .B(n14154), .Z(n596) );
  NAND U1453 ( .A(n595), .B(n596), .Z(n14258) );
  NAND U1454 ( .A(n14494), .B(n14493), .Z(n597) );
  NAND U1455 ( .A(n14492), .B(n14491), .Z(n598) );
  AND U1456 ( .A(n597), .B(n598), .Z(n14662) );
  NAND U1457 ( .A(n14500), .B(n14499), .Z(n599) );
  NANDN U1458 ( .A(n14502), .B(n14501), .Z(n600) );
  AND U1459 ( .A(n599), .B(n600), .Z(n14700) );
  XNOR U1460 ( .A(n10113), .B(o[107]), .Z(n10093) );
  XNOR U1461 ( .A(n10188), .B(n10793), .Z(n10167) );
  XNOR U1462 ( .A(n10271), .B(n10270), .Z(n10272) );
  NAND U1463 ( .A(n10241), .B(n10240), .Z(n601) );
  NANDN U1464 ( .A(n10808), .B(n10239), .Z(n602) );
  NAND U1465 ( .A(n601), .B(n602), .Z(n10349) );
  NAND U1466 ( .A(n10334), .B(n10333), .Z(n603) );
  NAND U1467 ( .A(n10376), .B(n12097), .Z(n604) );
  AND U1468 ( .A(n603), .B(n604), .Z(n10404) );
  XNOR U1469 ( .A(n10729), .B(n10728), .Z(n10689) );
  XOR U1470 ( .A(n10928), .B(n10927), .Z(n10982) );
  XNOR U1471 ( .A(n10989), .B(n10988), .Z(n10943) );
  XNOR U1472 ( .A(n11236), .B(n11235), .Z(n11194) );
  NAND U1473 ( .A(n11473), .B(n11472), .Z(n605) );
  NANDN U1474 ( .A(n11475), .B(n11474), .Z(n606) );
  NAND U1475 ( .A(n605), .B(n606), .Z(n11631) );
  NAND U1476 ( .A(n11452), .B(n11451), .Z(n607) );
  NANDN U1477 ( .A(n11454), .B(n11453), .Z(n608) );
  AND U1478 ( .A(n607), .B(n608), .Z(n11622) );
  XNOR U1479 ( .A(n7687), .B(n7686), .Z(n7710) );
  XNOR U1480 ( .A(n7701), .B(n7700), .Z(n7702) );
  XOR U1481 ( .A(n7827), .B(n7826), .Z(n7788) );
  OR U1482 ( .A(n7737), .B(n8695), .Z(n609) );
  NANDN U1483 ( .A(n7739), .B(n7738), .Z(n610) );
  AND U1484 ( .A(n609), .B(n610), .Z(n7836) );
  XOR U1485 ( .A(n8022), .B(n8021), .Z(n8076) );
  XNOR U1486 ( .A(n8038), .B(n8037), .Z(n8040) );
  XNOR U1487 ( .A(n7998), .B(n7997), .Z(n7999) );
  XNOR U1488 ( .A(n8332), .B(n8331), .Z(n8288) );
  XNOR U1489 ( .A(n8648), .B(n8647), .Z(n8592) );
  XNOR U1490 ( .A(n8720), .B(n8719), .Z(n8722) );
  XNOR U1491 ( .A(n8977), .B(n8976), .Z(n8978) );
  XNOR U1492 ( .A(n8927), .B(n8926), .Z(n8929) );
  XNOR U1493 ( .A(n8963), .B(n8962), .Z(n8965) );
  XNOR U1494 ( .A(n4571), .B(n4570), .Z(n4550) );
  NAND U1495 ( .A(n4654), .B(n4653), .Z(n611) );
  NANDN U1496 ( .A(n5441), .B(n4842), .Z(n612) );
  NAND U1497 ( .A(n611), .B(n612), .Z(n4750) );
  XNOR U1498 ( .A(n4958), .B(n4957), .Z(n4996) );
  NAND U1499 ( .A(n4743), .B(n4742), .Z(n613) );
  NANDN U1500 ( .A(n4745), .B(n4744), .Z(n614) );
  AND U1501 ( .A(n613), .B(n614), .Z(n4885) );
  XNOR U1502 ( .A(n4875), .B(n4874), .Z(n4898) );
  XNOR U1503 ( .A(n5242), .B(n5241), .Z(n5243) );
  XNOR U1504 ( .A(n5467), .B(n5466), .Z(n5469) );
  XNOR U1505 ( .A(n5693), .B(n5692), .Z(n5694) );
  XNOR U1506 ( .A(n5580), .B(n5579), .Z(n5582) );
  XNOR U1507 ( .A(n5925), .B(n5924), .Z(n5926) );
  XOR U1508 ( .A(n6094), .B(n6093), .Z(n6112) );
  XOR U1509 ( .A(n1404), .B(n1405), .Z(n1389) );
  XNOR U1510 ( .A(n1768), .B(n1767), .Z(n1770) );
  XNOR U1511 ( .A(n2077), .B(n2076), .Z(n2126) );
  AND U1512 ( .A(n2156), .B(n2155), .Z(n615) );
  AND U1513 ( .A(n3781), .B(y[1801]), .Z(n616) );
  NAND U1514 ( .A(x[225]), .B(n616), .Z(n617) );
  NANDN U1515 ( .A(n615), .B(n617), .Z(n2349) );
  NAND U1516 ( .A(n2362), .B(n2361), .Z(n618) );
  NANDN U1517 ( .A(n2364), .B(n2363), .Z(n619) );
  NAND U1518 ( .A(n618), .B(n619), .Z(n2408) );
  NAND U1519 ( .A(n2449), .B(n2448), .Z(n620) );
  NANDN U1520 ( .A(n2451), .B(n2450), .Z(n621) );
  NAND U1521 ( .A(n620), .B(n621), .Z(n2612) );
  XNOR U1522 ( .A(n2977), .B(n2978), .Z(n2959) );
  XNOR U1523 ( .A(n3045), .B(n3044), .Z(n3046) );
  XNOR U1524 ( .A(n21337), .B(o[231]), .Z(n21332) );
  XNOR U1525 ( .A(n21450), .B(n21449), .Z(n21451) );
  XOR U1526 ( .A(n21547), .B(n21546), .Z(n21549) );
  XNOR U1527 ( .A(n21737), .B(n21736), .Z(n21685) );
  XNOR U1528 ( .A(n21645), .B(n21644), .Z(n21666) );
  XOR U1529 ( .A(n22353), .B(n22352), .Z(n22357) );
  XNOR U1530 ( .A(n22484), .B(n22483), .Z(n22485) );
  XOR U1531 ( .A(n22474), .B(n22473), .Z(n22478) );
  NAND U1532 ( .A(n23214), .B(n23213), .Z(n622) );
  NAND U1533 ( .A(n23211), .B(n23212), .Z(n623) );
  AND U1534 ( .A(n622), .B(n623), .Z(n23484) );
  XNOR U1535 ( .A(n23601), .B(n23600), .Z(n23603) );
  XNOR U1536 ( .A(n23418), .B(n23417), .Z(n23439) );
  XNOR U1537 ( .A(n23395), .B(n23394), .Z(n23382) );
  XNOR U1538 ( .A(n23597), .B(n23596), .Z(n23645) );
  XNOR U1539 ( .A(n23565), .B(n23564), .Z(n23566) );
  XNOR U1540 ( .A(n23990), .B(n23759), .Z(n23760) );
  XOR U1541 ( .A(n18815), .B(n18816), .Z(n18800) );
  XNOR U1542 ( .A(n19359), .B(n19358), .Z(n19368) );
  XNOR U1543 ( .A(n19621), .B(n19620), .Z(n19622) );
  XOR U1544 ( .A(n20119), .B(n20118), .Z(n20124) );
  XNOR U1545 ( .A(n20308), .B(n20307), .Z(n20330) );
  XNOR U1546 ( .A(n20576), .B(n20575), .Z(n20519) );
  XNOR U1547 ( .A(n20564), .B(n20563), .Z(n20619) );
  AND U1548 ( .A(n20580), .B(n20579), .Z(n624) );
  AND U1549 ( .A(n20999), .B(y[1987]), .Z(n625) );
  NAND U1550 ( .A(x[244]), .B(n625), .Z(n626) );
  NANDN U1551 ( .A(n624), .B(n626), .Z(n20764) );
  NAND U1552 ( .A(n20584), .B(n20583), .Z(n627) );
  NAND U1553 ( .A(n20581), .B(n20582), .Z(n628) );
  NAND U1554 ( .A(n627), .B(n628), .Z(n20760) );
  NAND U1555 ( .A(n20678), .B(n20677), .Z(n629) );
  NAND U1556 ( .A(n20675), .B(n20676), .Z(n630) );
  NAND U1557 ( .A(n629), .B(n630), .Z(n20936) );
  AND U1558 ( .A(n20894), .B(o[221]), .Z(n21116) );
  XNOR U1559 ( .A(n20989), .B(n20887), .Z(n20888) );
  XNOR U1560 ( .A(n15619), .B(o[164]), .Z(n15621) );
  XOR U1561 ( .A(n15752), .B(n16543), .Z(n15754) );
  XOR U1562 ( .A(n15833), .B(n15832), .Z(n15821) );
  XOR U1563 ( .A(n15992), .B(n15991), .Z(n15986) );
  XNOR U1564 ( .A(n16297), .B(n16296), .Z(n16299) );
  NAND U1565 ( .A(n16325), .B(n16324), .Z(n631) );
  NANDN U1566 ( .A(n16327), .B(n16326), .Z(n632) );
  NAND U1567 ( .A(n631), .B(n632), .Z(n16483) );
  NAND U1568 ( .A(n16440), .B(n16439), .Z(n633) );
  NANDN U1569 ( .A(n16442), .B(n16441), .Z(n634) );
  AND U1570 ( .A(n633), .B(n634), .Z(n16573) );
  XNOR U1571 ( .A(n16610), .B(n16609), .Z(n16691) );
  XOR U1572 ( .A(n16670), .B(n16669), .Z(n16687) );
  XNOR U1573 ( .A(n16856), .B(n16855), .Z(n16857) );
  XOR U1574 ( .A(n17321), .B(n17320), .Z(n17326) );
  XNOR U1575 ( .A(n17494), .B(n17493), .Z(n17495) );
  OR U1576 ( .A(n17427), .B(n17428), .Z(n635) );
  NAND U1577 ( .A(n17425), .B(n17426), .Z(n636) );
  NAND U1578 ( .A(n635), .B(n636), .Z(n17594) );
  XNOR U1579 ( .A(n17724), .B(n17723), .Z(n17667) );
  NAND U1580 ( .A(n17621), .B(n17620), .Z(n637) );
  NAND U1581 ( .A(n17619), .B(n17618), .Z(n638) );
  NAND U1582 ( .A(n637), .B(n638), .Z(n17717) );
  NAND U1583 ( .A(n17607), .B(n17606), .Z(n639) );
  NANDN U1584 ( .A(n17604), .B(n17605), .Z(n640) );
  NAND U1585 ( .A(n639), .B(n640), .Z(n17710) );
  NAND U1586 ( .A(n17542), .B(n17541), .Z(n641) );
  NAND U1587 ( .A(n17540), .B(n17539), .Z(n642) );
  NAND U1588 ( .A(n641), .B(n642), .Z(n17670) );
  NAND U1589 ( .A(n17603), .B(n17602), .Z(n643) );
  NAND U1590 ( .A(n17600), .B(n17601), .Z(n644) );
  NAND U1591 ( .A(n643), .B(n644), .Z(n17769) );
  NAND U1592 ( .A(n17599), .B(n17598), .Z(n645) );
  NAND U1593 ( .A(n17597), .B(n17596), .Z(n646) );
  NAND U1594 ( .A(n645), .B(n646), .Z(n17660) );
  XNOR U1595 ( .A(n17980), .B(n17979), .Z(n17981) );
  NAND U1596 ( .A(n17854), .B(n17853), .Z(n647) );
  NAND U1597 ( .A(n17852), .B(n17851), .Z(n648) );
  NAND U1598 ( .A(n647), .B(n648), .Z(n18056) );
  XNOR U1599 ( .A(n18030), .B(n18029), .Z(n18050) );
  XNOR U1600 ( .A(n18234), .B(n18233), .Z(n18171) );
  XNOR U1601 ( .A(n13721), .B(n13720), .Z(n13723) );
  XNOR U1602 ( .A(n13709), .B(n13708), .Z(n13711) );
  XNOR U1603 ( .A(n13705), .B(n13704), .Z(n13630) );
  XNOR U1604 ( .A(n14331), .B(n14330), .Z(n14317) );
  XNOR U1605 ( .A(n14353), .B(n14352), .Z(n14456) );
  XOR U1606 ( .A(n14822), .B(n14821), .Z(n14852) );
  XOR U1607 ( .A(n15379), .B(n15378), .Z(n15377) );
  XOR U1608 ( .A(n14906), .B(n14905), .Z(n14908) );
  XNOR U1609 ( .A(n14773), .B(n14772), .Z(n14775) );
  XNOR U1610 ( .A(n10232), .B(n10231), .Z(n10224) );
  XNOR U1611 ( .A(n10356), .B(n10355), .Z(n10358) );
  NAND U1612 ( .A(n10348), .B(n10347), .Z(n649) );
  NANDN U1613 ( .A(n10346), .B(n10727), .Z(n650) );
  AND U1614 ( .A(n649), .B(n650), .Z(n10447) );
  XOR U1615 ( .A(n10880), .B(n10879), .Z(n10884) );
  XNOR U1616 ( .A(n10784), .B(n10783), .Z(n10865) );
  XOR U1617 ( .A(n10823), .B(n10822), .Z(n10861) );
  XNOR U1618 ( .A(n11033), .B(n11032), .Z(n11034) );
  XOR U1619 ( .A(n11929), .B(n11928), .Z(n11959) );
  XNOR U1620 ( .A(n11947), .B(n11946), .Z(n12013) );
  XOR U1621 ( .A(n11997), .B(n11996), .Z(n12007) );
  XOR U1622 ( .A(n7259), .B(n7260), .Z(n7244) );
  XNOR U1623 ( .A(n7954), .B(n7953), .Z(n7969) );
  XOR U1624 ( .A(n7915), .B(n7914), .Z(n7965) );
  XNOR U1625 ( .A(n8093), .B(n8092), .Z(n8095) );
  XNOR U1626 ( .A(n8131), .B(n8130), .Z(n8132) );
  XOR U1627 ( .A(n8600), .B(n8599), .Z(n8605) );
  XNOR U1628 ( .A(n8801), .B(n8800), .Z(n8802) );
  XNOR U1629 ( .A(n8678), .B(n8677), .Z(n8680) );
  XNOR U1630 ( .A(n8996), .B(n8995), .Z(n8998) );
  XNOR U1631 ( .A(n8842), .B(n8841), .Z(n8844) );
  XNOR U1632 ( .A(n9061), .B(n9060), .Z(n9004) );
  XNOR U1633 ( .A(n9047), .B(n9046), .Z(n9049) );
  XNOR U1634 ( .A(n9008), .B(n9007), .Z(n9010) );
  XOR U1635 ( .A(n9444), .B(n9443), .Z(n9445) );
  XNOR U1636 ( .A(n3988), .B(o[38]), .Z(n3980) );
  XOR U1637 ( .A(n4059), .B(n4854), .Z(n4061) );
  XNOR U1638 ( .A(n4136), .B(n4135), .Z(n4137) );
  NAND U1639 ( .A(n4245), .B(n4244), .Z(n651) );
  NAND U1640 ( .A(n4520), .B(n5336), .Z(n652) );
  AND U1641 ( .A(n651), .B(n652), .Z(n4312) );
  XNOR U1642 ( .A(n5298), .B(n5297), .Z(n5299) );
  XNOR U1643 ( .A(n5539), .B(n5538), .Z(n5540) );
  XNOR U1644 ( .A(n5547), .B(n5546), .Z(n5533) );
  XNOR U1645 ( .A(n5836), .B(n5835), .Z(n5839) );
  NAND U1646 ( .A(n5891), .B(n5890), .Z(n653) );
  NANDN U1647 ( .A(n5893), .B(n5892), .Z(n654) );
  AND U1648 ( .A(n653), .B(n654), .Z(n6156) );
  XOR U1649 ( .A(n6348), .B(n6347), .Z(n6318) );
  NAND U1650 ( .A(n6106), .B(n6105), .Z(n655) );
  NANDN U1651 ( .A(n6104), .B(n6103), .Z(n656) );
  AND U1652 ( .A(n655), .B(n656), .Z(n6311) );
  XOR U1653 ( .A(n6249), .B(n6248), .Z(n6330) );
  XNOR U1654 ( .A(n6334), .B(n6333), .Z(n6335) );
  XNOR U1655 ( .A(n6270), .B(n6461), .Z(n6271) );
  XNOR U1656 ( .A(n1453), .B(n1452), .Z(n1455) );
  XNOR U1657 ( .A(n1917), .B(n1916), .Z(n1919) );
  XOR U1658 ( .A(n2134), .B(n2133), .Z(n2138) );
  XOR U1659 ( .A(n2048), .B(n2047), .Z(n2050) );
  NAND U1660 ( .A(n2417), .B(n2416), .Z(n657) );
  NANDN U1661 ( .A(n2415), .B(n2414), .Z(n658) );
  NAND U1662 ( .A(n657), .B(n658), .Z(n2566) );
  NAND U1663 ( .A(n2488), .B(n2487), .Z(n659) );
  NANDN U1664 ( .A(n2486), .B(n2485), .Z(n660) );
  NAND U1665 ( .A(n659), .B(n660), .Z(n2626) );
  XNOR U1666 ( .A(n3041), .B(n3040), .Z(n3035) );
  XNOR U1667 ( .A(n3079), .B(n3078), .Z(n2947) );
  NAND U1668 ( .A(n3171), .B(n3170), .Z(n661) );
  NANDN U1669 ( .A(n3169), .B(n3168), .Z(n662) );
  NAND U1670 ( .A(n661), .B(n662), .Z(n3362) );
  NAND U1671 ( .A(n3128), .B(n3127), .Z(n663) );
  NANDN U1672 ( .A(n3126), .B(n3125), .Z(n664) );
  NAND U1673 ( .A(n663), .B(n664), .Z(n3374) );
  NAND U1674 ( .A(n3142), .B(n3141), .Z(n665) );
  NANDN U1675 ( .A(n3144), .B(n3143), .Z(n666) );
  NAND U1676 ( .A(n665), .B(n666), .Z(n3350) );
  XNOR U1677 ( .A(n21288), .B(n21287), .Z(n21290) );
  XOR U1678 ( .A(n21340), .B(n21265), .Z(n667) );
  NANDN U1679 ( .A(n21266), .B(n667), .Z(n668) );
  NAND U1680 ( .A(n21340), .B(n21265), .Z(n669) );
  AND U1681 ( .A(n668), .B(n669), .Z(n21318) );
  XNOR U1682 ( .A(n21751), .B(n21750), .Z(n21752) );
  XNOR U1683 ( .A(n22745), .B(n22744), .Z(n22637) );
  XNOR U1684 ( .A(n23051), .B(n23050), .Z(n23053) );
  XNOR U1685 ( .A(n23363), .B(n23362), .Z(n23365) );
  XOR U1686 ( .A(n23371), .B(n23370), .Z(n23357) );
  XNOR U1687 ( .A(n23584), .B(n23583), .Z(n23614) );
  XNOR U1688 ( .A(n23538), .B(n23537), .Z(n23658) );
  XNOR U1689 ( .A(n23633), .B(n23632), .Z(n23634) );
  XNOR U1690 ( .A(n23526), .B(n23525), .Z(n23519) );
  XNOR U1691 ( .A(n23718), .B(n23717), .Z(n23719) );
  XNOR U1692 ( .A(n23803), .B(n23802), .Z(n23804) );
  XNOR U1693 ( .A(n23764), .B(n23917), .Z(n23765) );
  XNOR U1694 ( .A(n23815), .B(n23814), .Z(n23816) );
  XOR U1695 ( .A(n23906), .B(n23905), .Z(n23904) );
  XOR U1696 ( .A(n23898), .B(n23897), .Z(n23896) );
  XNOR U1697 ( .A(n18525), .B(n18524), .Z(n18526) );
  XOR U1698 ( .A(n19399), .B(n19398), .Z(n19499) );
  XNOR U1699 ( .A(n19492), .B(n19491), .Z(n19493) );
  XNOR U1700 ( .A(n19766), .B(n19765), .Z(n19768) );
  XNOR U1701 ( .A(n19880), .B(n19879), .Z(n19882) );
  XNOR U1702 ( .A(n20058), .B(n20057), .Z(n20052) );
  XOR U1703 ( .A(n20201), .B(n20200), .Z(n20203) );
  XNOR U1704 ( .A(n20326), .B(n20325), .Z(n20195) );
  XNOR U1705 ( .A(n20343), .B(n20342), .Z(n20344) );
  XNOR U1706 ( .A(n20499), .B(n20498), .Z(n20501) );
  XOR U1707 ( .A(n20775), .B(n20774), .Z(n20650) );
  NAND U1708 ( .A(n20757), .B(n20756), .Z(n670) );
  NAND U1709 ( .A(n20755), .B(n20754), .Z(n671) );
  NAND U1710 ( .A(n670), .B(n671), .Z(n20898) );
  NAND U1711 ( .A(n20712), .B(n20711), .Z(n672) );
  NANDN U1712 ( .A(n20710), .B(n20709), .Z(n673) );
  NAND U1713 ( .A(n672), .B(n673), .Z(n20822) );
  NAND U1714 ( .A(n20729), .B(n20728), .Z(n674) );
  NAND U1715 ( .A(n20727), .B(n20726), .Z(n675) );
  NAND U1716 ( .A(n674), .B(n675), .Z(n20902) );
  NAND U1717 ( .A(n20706), .B(n20705), .Z(n676) );
  NAND U1718 ( .A(n20704), .B(n20703), .Z(n677) );
  NAND U1719 ( .A(n676), .B(n677), .Z(n20875) );
  NAND U1720 ( .A(n20916), .B(n20915), .Z(n678) );
  NANDN U1721 ( .A(n20918), .B(n20917), .Z(n679) );
  AND U1722 ( .A(n678), .B(n679), .Z(n21142) );
  XNOR U1723 ( .A(n21136), .B(n21135), .Z(n21134) );
  NAND U1724 ( .A(n20883), .B(n20882), .Z(n680) );
  NAND U1725 ( .A(n20880), .B(n20881), .Z(n681) );
  NAND U1726 ( .A(n680), .B(n681), .Z(n20976) );
  XOR U1727 ( .A(n21093), .B(n21094), .Z(n21095) );
  NAND U1728 ( .A(n20687), .B(n20686), .Z(n682) );
  NAND U1729 ( .A(n20685), .B(n20684), .Z(n683) );
  AND U1730 ( .A(n682), .B(n683), .Z(n20907) );
  XOR U1731 ( .A(n20971), .B(n20970), .Z(n20969) );
  XNOR U1732 ( .A(n15733), .B(n15732), .Z(n15734) );
  XNOR U1733 ( .A(n15847), .B(n15846), .Z(n15848) );
  XOR U1734 ( .A(n16287), .B(n16286), .Z(n16279) );
  XNOR U1735 ( .A(n16704), .B(n16703), .Z(n16705) );
  XOR U1736 ( .A(n16823), .B(n16822), .Z(n16827) );
  XNOR U1737 ( .A(n16992), .B(n16991), .Z(n16986) );
  XNOR U1738 ( .A(n17653), .B(n17652), .Z(n17655) );
  NAND U1739 ( .A(n17629), .B(n17628), .Z(n684) );
  NANDN U1740 ( .A(n17631), .B(n17630), .Z(n685) );
  AND U1741 ( .A(n684), .B(n685), .Z(n17648) );
  XNOR U1742 ( .A(n17815), .B(n17814), .Z(n17801) );
  NAND U1743 ( .A(n17884), .B(n17883), .Z(n686) );
  NANDN U1744 ( .A(n17882), .B(n17881), .Z(n687) );
  NAND U1745 ( .A(n686), .B(n687), .Z(n17963) );
  NAND U1746 ( .A(n17888), .B(n17887), .Z(n688) );
  NAND U1747 ( .A(n17886), .B(n17885), .Z(n689) );
  NAND U1748 ( .A(n688), .B(n689), .Z(n18043) );
  XNOR U1749 ( .A(n18103), .B(n18102), .Z(n18100) );
  NAND U1750 ( .A(n17869), .B(n17868), .Z(n690) );
  NAND U1751 ( .A(n17867), .B(n17866), .Z(n691) );
  NAND U1752 ( .A(n690), .B(n691), .Z(n18015) );
  OR U1753 ( .A(n18061), .B(n18060), .Z(n692) );
  NAND U1754 ( .A(n18063), .B(n18062), .Z(n693) );
  NAND U1755 ( .A(n692), .B(n693), .Z(n18287) );
  XNOR U1756 ( .A(n18284), .B(n18283), .Z(n18281) );
  XOR U1757 ( .A(n18113), .B(n18112), .Z(n18111) );
  NAND U1758 ( .A(n12862), .B(n13672), .Z(n694) );
  NANDN U1759 ( .A(n12864), .B(n12863), .Z(n695) );
  AND U1760 ( .A(n694), .B(n695), .Z(n12893) );
  XOR U1761 ( .A(n13044), .B(n13043), .Z(n13046) );
  XOR U1762 ( .A(n13383), .B(n13382), .Z(n13385) );
  XNOR U1763 ( .A(n13953), .B(n13952), .Z(n13955) );
  NAND U1764 ( .A(n14074), .B(n14073), .Z(n696) );
  NANDN U1765 ( .A(n14076), .B(n14075), .Z(n697) );
  AND U1766 ( .A(n696), .B(n697), .Z(n14103) );
  XNOR U1767 ( .A(n14472), .B(n14471), .Z(n14473) );
  NAND U1768 ( .A(n14486), .B(n14485), .Z(n698) );
  NAND U1769 ( .A(n14484), .B(n14483), .Z(n699) );
  NAND U1770 ( .A(n698), .B(n699), .Z(n14750) );
  NAND U1771 ( .A(n14593), .B(n14592), .Z(n700) );
  NAND U1772 ( .A(n14591), .B(n14590), .Z(n701) );
  AND U1773 ( .A(n700), .B(n701), .Z(n14609) );
  XNOR U1774 ( .A(n15049), .B(n15048), .Z(n15050) );
  XNOR U1775 ( .A(n15061), .B(n15060), .Z(n15063) );
  XNOR U1776 ( .A(n15223), .B(n15222), .Z(n15224) );
  XNOR U1777 ( .A(n15156), .B(n15155), .Z(n15234) );
  XOR U1778 ( .A(n15247), .B(n15246), .Z(n15248) );
  XOR U1779 ( .A(n14942), .B(n14941), .Z(n14928) );
  XOR U1780 ( .A(n9891), .B(n9800), .Z(n702) );
  NANDN U1781 ( .A(n9801), .B(n702), .Z(n703) );
  NAND U1782 ( .A(n9891), .B(n9800), .Z(n704) );
  AND U1783 ( .A(n703), .B(n704), .Z(n9857) );
  XNOR U1784 ( .A(n10212), .B(n10211), .Z(n10214) );
  XOR U1785 ( .A(n10432), .B(n10431), .Z(n10460) );
  XOR U1786 ( .A(n11001), .B(n11000), .Z(n11005) );
  XNOR U1787 ( .A(n11173), .B(n11172), .Z(n11167) );
  XNOR U1788 ( .A(n12021), .B(n12020), .Z(n11878) );
  XNOR U1789 ( .A(n12163), .B(n12162), .Z(n12165) );
  XNOR U1790 ( .A(n12324), .B(n12323), .Z(n12325) );
  XNOR U1791 ( .A(n12287), .B(n12286), .Z(n12335) );
  XOR U1792 ( .A(n12348), .B(n12347), .Z(n12349) );
  XNOR U1793 ( .A(n12569), .B(n12568), .Z(n12570) );
  XOR U1794 ( .A(n12556), .B(n12557), .Z(n12558) );
  XNOR U1795 ( .A(n12399), .B(n12398), .Z(n12400) );
  XOR U1796 ( .A(n12393), .B(n12392), .Z(n12394) );
  XNOR U1797 ( .A(n12187), .B(n12186), .Z(n12188) );
  XNOR U1798 ( .A(n6961), .B(n6960), .Z(n6962) );
  XNOR U1799 ( .A(n6987), .B(n6986), .Z(n6989) );
  XOR U1800 ( .A(n6975), .B(n6891), .Z(n705) );
  NANDN U1801 ( .A(n6892), .B(n705), .Z(n706) );
  NAND U1802 ( .A(n6975), .B(n6891), .Z(n707) );
  AND U1803 ( .A(n706), .B(n707), .Z(n6940) );
  XOR U1804 ( .A(n7194), .B(n7193), .Z(n7196) );
  XOR U1805 ( .A(n7533), .B(n7532), .Z(n7535) );
  XNOR U1806 ( .A(n7976), .B(n7975), .Z(n7977) );
  XNOR U1807 ( .A(n8267), .B(n8266), .Z(n8261) );
  XNOR U1808 ( .A(n8672), .B(n8671), .Z(n8674) );
  XNOR U1809 ( .A(n8541), .B(n8540), .Z(n8535) );
  XOR U1810 ( .A(n9149), .B(n9148), .Z(n9143) );
  NAND U1811 ( .A(n9028), .B(n9027), .Z(n708) );
  NAND U1812 ( .A(n9026), .B(n9025), .Z(n709) );
  NAND U1813 ( .A(n708), .B(n709), .Z(n9232) );
  XNOR U1814 ( .A(n9250), .B(n9249), .Z(n9251) );
  XNOR U1815 ( .A(n9262), .B(n9261), .Z(n9263) );
  XNOR U1816 ( .A(n9440), .B(n9439), .Z(n9420) );
  NAND U1817 ( .A(n9276), .B(n9275), .Z(n710) );
  NAND U1818 ( .A(n9274), .B(n9273), .Z(n711) );
  NAND U1819 ( .A(n710), .B(n711), .Z(n9415) );
  NAND U1820 ( .A(n9248), .B(n9247), .Z(n712) );
  NAND U1821 ( .A(n9246), .B(n9245), .Z(n713) );
  NAND U1822 ( .A(n712), .B(n713), .Z(n9424) );
  XOR U1823 ( .A(n9564), .B(n9450), .Z(n714) );
  NANDN U1824 ( .A(n9449), .B(n714), .Z(n715) );
  NAND U1825 ( .A(n9564), .B(n9450), .Z(n716) );
  AND U1826 ( .A(n715), .B(n716), .Z(n9682) );
  XOR U1827 ( .A(n9486), .B(n9485), .Z(n9484) );
  NAND U1828 ( .A(n9227), .B(n9226), .Z(n717) );
  NAND U1829 ( .A(n9225), .B(n9224), .Z(n718) );
  NAND U1830 ( .A(n717), .B(n718), .Z(n9409) );
  NAND U1831 ( .A(n9462), .B(n9461), .Z(n719) );
  NANDN U1832 ( .A(n9464), .B(n9463), .Z(n720) );
  AND U1833 ( .A(n719), .B(n720), .Z(n9679) );
  XNOR U1834 ( .A(n9688), .B(n9687), .Z(n9686) );
  NAND U1835 ( .A(n9200), .B(n9199), .Z(n721) );
  NAND U1836 ( .A(n9198), .B(n9197), .Z(n722) );
  AND U1837 ( .A(n721), .B(n722), .Z(n9429) );
  XNOR U1838 ( .A(n9662), .B(n9661), .Z(n9659) );
  XOR U1839 ( .A(n9498), .B(n9497), .Z(n9496) );
  XNOR U1840 ( .A(n4013), .B(n4012), .Z(n4014) );
  XNOR U1841 ( .A(n4038), .B(n4037), .Z(n4040) );
  XOR U1842 ( .A(n4026), .B(n3939), .Z(n723) );
  NANDN U1843 ( .A(n3940), .B(n723), .Z(n724) );
  NAND U1844 ( .A(n4026), .B(n3939), .Z(n725) );
  AND U1845 ( .A(n724), .B(n725), .Z(n3992) );
  NAND U1846 ( .A(n4287), .B(n4286), .Z(n726) );
  NANDN U1847 ( .A(n4285), .B(n4284), .Z(n727) );
  AND U1848 ( .A(n726), .B(n727), .Z(n4354) );
  XOR U1849 ( .A(n4575), .B(n4574), .Z(n4577) );
  XNOR U1850 ( .A(n4928), .B(n4927), .Z(n5029) );
  XOR U1851 ( .A(n5402), .B(n5401), .Z(n5293) );
  XNOR U1852 ( .A(n6041), .B(n6040), .Z(n6019) );
  XNOR U1853 ( .A(n6283), .B(n6282), .Z(n6284) );
  XNOR U1854 ( .A(n6482), .B(n6481), .Z(n6484) );
  XNOR U1855 ( .A(n6384), .B(n6383), .Z(n6385) );
  XOR U1856 ( .A(n6636), .B(n6635), .Z(n6634) );
  XNOR U1857 ( .A(n6547), .B(n6548), .Z(n6549) );
  XNOR U1858 ( .A(n6444), .B(n6443), .Z(n6487) );
  XOR U1859 ( .A(n6656), .B(n6655), .Z(n6654) );
  XNOR U1860 ( .A(n1164), .B(n1163), .Z(n1165) );
  XNOR U1861 ( .A(n1170), .B(n1169), .Z(n1171) );
  XNOR U1862 ( .A(n1530), .B(n1529), .Z(n1532) );
  XOR U1863 ( .A(n1897), .B(n1896), .Z(n1812) );
  NAND U1864 ( .A(n2366), .B(n2365), .Z(n728) );
  NANDN U1865 ( .A(n2368), .B(n2367), .Z(n729) );
  AND U1866 ( .A(n728), .B(n729), .Z(n2399) );
  XNOR U1867 ( .A(n2793), .B(n2792), .Z(n2795) );
  XNOR U1868 ( .A(n2787), .B(n2786), .Z(n2789) );
  XNOR U1869 ( .A(n3329), .B(n3328), .Z(n3353) );
  XNOR U1870 ( .A(n3244), .B(n3243), .Z(n3245) );
  XNOR U1871 ( .A(n3816), .B(n3815), .Z(n3814) );
  XOR U1872 ( .A(n3636), .B(n3635), .Z(n3634) );
  XOR U1873 ( .A(n3616), .B(n3615), .Z(n3614) );
  XNOR U1874 ( .A(n21833), .B(n21832), .Z(n21835) );
  XNOR U1875 ( .A(n23706), .B(n23705), .Z(n23708) );
  XNOR U1876 ( .A(n23700), .B(n23699), .Z(n23702) );
  XNOR U1877 ( .A(n23799), .B(n23798), .Z(n23712) );
  XOR U1878 ( .A(n24134), .B(n24133), .Z(n24132) );
  XOR U1879 ( .A(n24110), .B(n24109), .Z(n24108) );
  NAND U1880 ( .A(n19053), .B(n19052), .Z(n730) );
  NANDN U1881 ( .A(n19051), .B(n19050), .Z(n731) );
  AND U1882 ( .A(n730), .B(n731), .Z(n19082) );
  XNOR U1883 ( .A(n15909), .B(n15908), .Z(n15910) );
  XNOR U1884 ( .A(n15980), .B(n15979), .Z(n16049) );
  XNOR U1885 ( .A(n16122), .B(n16121), .Z(n16123) );
  XOR U1886 ( .A(n17244), .B(n17243), .Z(n17246) );
  XNOR U1887 ( .A(n17944), .B(n17943), .Z(n17949) );
  NAND U1888 ( .A(n17993), .B(n17992), .Z(n732) );
  NAND U1889 ( .A(n17991), .B(n17990), .Z(n733) );
  AND U1890 ( .A(n732), .B(n733), .Z(n18081) );
  NAND U1891 ( .A(n18047), .B(n18046), .Z(n734) );
  NANDN U1892 ( .A(n18049), .B(n18048), .Z(n735) );
  AND U1893 ( .A(n734), .B(n735), .Z(n18297) );
  NAND U1894 ( .A(n17972), .B(n17971), .Z(n736) );
  NAND U1895 ( .A(n17969), .B(n17970), .Z(n737) );
  AND U1896 ( .A(n736), .B(n737), .Z(n18085) );
  NAND U1897 ( .A(n12748), .B(n12831), .Z(n738) );
  XOR U1898 ( .A(n12748), .B(n12831), .Z(n739) );
  NANDN U1899 ( .A(n12747), .B(n739), .Z(n740) );
  NAND U1900 ( .A(n738), .B(n740), .Z(n12801) );
  XNOR U1901 ( .A(n13229), .B(n13228), .Z(n13231) );
  XNOR U1902 ( .A(n13318), .B(n13317), .Z(n13320) );
  XOR U1903 ( .A(n13436), .B(n13435), .Z(n13423) );
  XNOR U1904 ( .A(n13521), .B(n13520), .Z(n13523) );
  XNOR U1905 ( .A(n13959), .B(n13958), .Z(n13960) );
  XOR U1906 ( .A(n15229), .B(n15228), .Z(n15231) );
  XNOR U1907 ( .A(n15286), .B(n15285), .Z(n15524) );
  XNOR U1908 ( .A(n15500), .B(n15499), .Z(n15498) );
  XNOR U1909 ( .A(n9820), .B(n9819), .Z(n9821) );
  XOR U1910 ( .A(n9958), .B(n9957), .Z(n9997) );
  XNOR U1911 ( .A(n10552), .B(n10551), .Z(n10554) );
  XOR U1912 ( .A(n11421), .B(n11420), .Z(n11423) );
  XNOR U1913 ( .A(n12330), .B(n12329), .Z(n12332) );
  XOR U1914 ( .A(n12649), .B(n12648), .Z(n741) );
  XNOR U1915 ( .A(n12650), .B(n741), .Z(n12634) );
  XNOR U1916 ( .A(n12625), .B(n12624), .Z(n12623) );
  XNOR U1917 ( .A(n12601), .B(n12600), .Z(n12599) );
  XNOR U1918 ( .A(n6853), .B(o[67]), .Z(n6855) );
  XNOR U1919 ( .A(n7040), .B(n7039), .Z(n7042) );
  XOR U1920 ( .A(n7582), .B(n7581), .Z(n7569) );
  XNOR U1921 ( .A(n7666), .B(n7665), .Z(n7668) );
  XOR U1922 ( .A(n8519), .B(n8518), .Z(n8521) );
  XNOR U1923 ( .A(n9293), .B(n9292), .Z(n9295) );
  XNOR U1924 ( .A(n4091), .B(n4090), .Z(n4093) );
  XNOR U1925 ( .A(n4206), .B(n4205), .Z(n4208) );
  XNOR U1926 ( .A(n4213), .B(n4212), .Z(n4214) );
  XNOR U1927 ( .A(n5279), .B(n5278), .Z(n5281) );
  XOR U1928 ( .A(n5853), .B(n5852), .Z(n5855) );
  XNOR U1929 ( .A(n5860), .B(n5859), .Z(n5862) );
  XNOR U1930 ( .A(n6476), .B(n6475), .Z(n6477) );
  XOR U1931 ( .A(n6538), .B(n6537), .Z(n6536) );
  XNOR U1932 ( .A(n6780), .B(n6779), .Z(n6778) );
  XOR U1933 ( .A(n994), .B(n993), .Z(n742) );
  NANDN U1934 ( .A(n995), .B(n742), .Z(n743) );
  NAND U1935 ( .A(n994), .B(n993), .Z(n744) );
  AND U1936 ( .A(n743), .B(n744), .Z(n1016) );
  XNOR U1937 ( .A(n1301), .B(n1300), .Z(n1303) );
  XOR U1938 ( .A(n21278), .B(n21277), .Z(n745) );
  NANDN U1939 ( .A(n21279), .B(n745), .Z(n746) );
  NAND U1940 ( .A(n21278), .B(n21277), .Z(n747) );
  AND U1941 ( .A(n746), .B(n747), .Z(n21313) );
  XOR U1942 ( .A(n21459), .B(n21460), .Z(n748) );
  NANDN U1943 ( .A(n21461), .B(n748), .Z(n749) );
  NAND U1944 ( .A(n21459), .B(n21460), .Z(n750) );
  AND U1945 ( .A(n749), .B(n750), .Z(n21528) );
  XOR U1946 ( .A(n21740), .B(n21741), .Z(n751) );
  NANDN U1947 ( .A(n21742), .B(n751), .Z(n752) );
  NAND U1948 ( .A(n21740), .B(n21741), .Z(n753) );
  AND U1949 ( .A(n752), .B(n753), .Z(n21827) );
  XOR U1950 ( .A(n22489), .B(n22490), .Z(n754) );
  NANDN U1951 ( .A(n22491), .B(n754), .Z(n755) );
  NAND U1952 ( .A(n22489), .B(n22490), .Z(n756) );
  AND U1953 ( .A(n755), .B(n756), .Z(n22616) );
  XNOR U1954 ( .A(n22758), .B(n22757), .Z(n22751) );
  XOR U1955 ( .A(n23034), .B(n23035), .Z(n757) );
  NANDN U1956 ( .A(n23036), .B(n757), .Z(n758) );
  NAND U1957 ( .A(n23034), .B(n23035), .Z(n759) );
  AND U1958 ( .A(n758), .B(n759), .Z(n23187) );
  NAND U1959 ( .A(n23508), .B(n23509), .Z(n760) );
  XOR U1960 ( .A(n23508), .B(n23509), .Z(n761) );
  NANDN U1961 ( .A(n23507), .B(n761), .Z(n762) );
  NAND U1962 ( .A(n760), .B(n762), .Z(n23674) );
  XNOR U1963 ( .A(n24146), .B(n24145), .Z(n24144) );
  XOR U1964 ( .A(n18418), .B(n18419), .Z(n763) );
  NANDN U1965 ( .A(n18420), .B(n763), .Z(n764) );
  NAND U1966 ( .A(n18418), .B(n18419), .Z(n765) );
  AND U1967 ( .A(n764), .B(n765), .Z(n18449) );
  XOR U1968 ( .A(n18530), .B(n18531), .Z(n766) );
  NANDN U1969 ( .A(n18532), .B(n766), .Z(n767) );
  NAND U1970 ( .A(n18530), .B(n18531), .Z(n768) );
  AND U1971 ( .A(n767), .B(n768), .Z(n18583) );
  XOR U1972 ( .A(n18694), .B(n18695), .Z(n769) );
  NANDN U1973 ( .A(n18696), .B(n769), .Z(n770) );
  NAND U1974 ( .A(n18694), .B(n18695), .Z(n771) );
  AND U1975 ( .A(n770), .B(n771), .Z(n18761) );
  XOR U1976 ( .A(n19072), .B(n19073), .Z(n772) );
  NANDN U1977 ( .A(n19074), .B(n772), .Z(n773) );
  NAND U1978 ( .A(n19072), .B(n19073), .Z(n774) );
  AND U1979 ( .A(n773), .B(n774), .Z(n19089) );
  NAND U1980 ( .A(n19393), .B(n19394), .Z(n775) );
  XOR U1981 ( .A(n19393), .B(n19394), .Z(n776) );
  NANDN U1982 ( .A(n19392), .B(n776), .Z(n777) );
  NAND U1983 ( .A(n775), .B(n777), .Z(n19503) );
  XOR U1984 ( .A(n19755), .B(n19756), .Z(n778) );
  NANDN U1985 ( .A(n19757), .B(n778), .Z(n779) );
  NAND U1986 ( .A(n19755), .B(n19756), .Z(n780) );
  AND U1987 ( .A(n779), .B(n780), .Z(n19887) );
  NAND U1988 ( .A(n20182), .B(n20183), .Z(n781) );
  XOR U1989 ( .A(n20182), .B(n20183), .Z(n782) );
  NANDN U1990 ( .A(n20181), .B(n782), .Z(n783) );
  NAND U1991 ( .A(n781), .B(n783), .Z(n20191) );
  NAND U1992 ( .A(n20637), .B(n20638), .Z(n784) );
  XOR U1993 ( .A(n20637), .B(n20638), .Z(n785) );
  NANDN U1994 ( .A(n20636), .B(n785), .Z(n786) );
  NAND U1995 ( .A(n784), .B(n786), .Z(n20647) );
  XOR U1996 ( .A(n15629), .B(n15630), .Z(n787) );
  NANDN U1997 ( .A(n15631), .B(n787), .Z(n788) );
  NAND U1998 ( .A(n15629), .B(n15630), .Z(n789) );
  AND U1999 ( .A(n788), .B(n789), .Z(n15657) );
  NAND U2000 ( .A(n15745), .B(n15746), .Z(n790) );
  XOR U2001 ( .A(n15745), .B(n15746), .Z(n791) );
  NANDN U2002 ( .A(n15744), .B(n791), .Z(n792) );
  NAND U2003 ( .A(n790), .B(n792), .Z(n15791) );
  XOR U2004 ( .A(n15898), .B(n15899), .Z(n793) );
  NANDN U2005 ( .A(n15900), .B(n793), .Z(n794) );
  NAND U2006 ( .A(n15898), .B(n15899), .Z(n795) );
  AND U2007 ( .A(n794), .B(n795), .Z(n15916) );
  XOR U2008 ( .A(n16393), .B(n16394), .Z(n796) );
  NANDN U2009 ( .A(n16395), .B(n796), .Z(n797) );
  NAND U2010 ( .A(n16393), .B(n16394), .Z(n798) );
  AND U2011 ( .A(n797), .B(n798), .Z(n16496) );
  NAND U2012 ( .A(n16716), .B(n16717), .Z(n799) );
  XOR U2013 ( .A(n16716), .B(n16717), .Z(n800) );
  NANDN U2014 ( .A(n16715), .B(n800), .Z(n801) );
  NAND U2015 ( .A(n799), .B(n801), .Z(n16839) );
  NAND U2016 ( .A(n16981), .B(n16982), .Z(n802) );
  XOR U2017 ( .A(n16981), .B(n16982), .Z(n803) );
  NAND U2018 ( .A(n803), .B(n16980), .Z(n804) );
  NAND U2019 ( .A(n802), .B(n804), .Z(n17238) );
  XOR U2020 ( .A(n17798), .B(n17797), .Z(n805) );
  NANDN U2021 ( .A(n17799), .B(n805), .Z(n806) );
  NAND U2022 ( .A(n17798), .B(n17797), .Z(n807) );
  AND U2023 ( .A(n806), .B(n807), .Z(n17926) );
  NAND U2024 ( .A(n18040), .B(n18039), .Z(n808) );
  NAND U2025 ( .A(n18038), .B(n18037), .Z(n809) );
  NAND U2026 ( .A(n808), .B(n809), .Z(n18333) );
  XOR U2027 ( .A(n12759), .B(n12760), .Z(n810) );
  NANDN U2028 ( .A(n12761), .B(n810), .Z(n811) );
  NAND U2029 ( .A(n12759), .B(n12760), .Z(n812) );
  AND U2030 ( .A(n811), .B(n812), .Z(n12794) );
  XOR U2031 ( .A(n12855), .B(n12856), .Z(n813) );
  NANDN U2032 ( .A(n12857), .B(n813), .Z(n814) );
  NAND U2033 ( .A(n12855), .B(n12856), .Z(n815) );
  AND U2034 ( .A(n814), .B(n815), .Z(n12942) );
  XOR U2035 ( .A(n13143), .B(n13144), .Z(n816) );
  NANDN U2036 ( .A(n13145), .B(n816), .Z(n817) );
  NAND U2037 ( .A(n13143), .B(n13144), .Z(n818) );
  AND U2038 ( .A(n817), .B(n818), .Z(n13223) );
  XOR U2039 ( .A(n13842), .B(n13843), .Z(n819) );
  NANDN U2040 ( .A(n13844), .B(n819), .Z(n820) );
  NAND U2041 ( .A(n13842), .B(n13843), .Z(n821) );
  AND U2042 ( .A(n820), .B(n821), .Z(n13965) );
  XOR U2043 ( .A(n14099), .B(n14100), .Z(n822) );
  NANDN U2044 ( .A(n14101), .B(n822), .Z(n823) );
  NAND U2045 ( .A(n14099), .B(n14100), .Z(n824) );
  AND U2046 ( .A(n823), .B(n824), .Z(n14341) );
  XOR U2047 ( .A(n14598), .B(n14599), .Z(n825) );
  NANDN U2048 ( .A(n14600), .B(n825), .Z(n826) );
  NAND U2049 ( .A(n14598), .B(n14599), .Z(n827) );
  AND U2050 ( .A(n826), .B(n827), .Z(n14760) );
  XOR U2051 ( .A(n15085), .B(n15084), .Z(n828) );
  NANDN U2052 ( .A(n15086), .B(n828), .Z(n829) );
  NAND U2053 ( .A(n15085), .B(n15084), .Z(n830) );
  AND U2054 ( .A(n829), .B(n830), .Z(n15095) );
  XOR U2055 ( .A(n15559), .B(n15560), .Z(n15561) );
  XOR U2056 ( .A(n9787), .B(n9786), .Z(n831) );
  NANDN U2057 ( .A(n9788), .B(n831), .Z(n832) );
  NAND U2058 ( .A(n9787), .B(n9786), .Z(n833) );
  AND U2059 ( .A(n832), .B(n833), .Z(n9814) );
  XOR U2060 ( .A(n9915), .B(n9916), .Z(n834) );
  NANDN U2061 ( .A(n9917), .B(n834), .Z(n835) );
  NAND U2062 ( .A(n9915), .B(n9916), .Z(n836) );
  AND U2063 ( .A(n835), .B(n836), .Z(n10002) );
  XOR U2064 ( .A(n10361), .B(n10362), .Z(n837) );
  NANDN U2065 ( .A(n10363), .B(n837), .Z(n838) );
  NAND U2066 ( .A(n10361), .B(n10362), .Z(n839) );
  AND U2067 ( .A(n838), .B(n839), .Z(n10455) );
  XOR U2068 ( .A(n10771), .B(n10772), .Z(n840) );
  NANDN U2069 ( .A(n10773), .B(n840), .Z(n841) );
  NAND U2070 ( .A(n10771), .B(n10772), .Z(n842) );
  AND U2071 ( .A(n841), .B(n842), .Z(n10896) );
  NAND U2072 ( .A(n11162), .B(n11163), .Z(n843) );
  XOR U2073 ( .A(n11162), .B(n11163), .Z(n844) );
  NAND U2074 ( .A(n844), .B(n11161), .Z(n845) );
  NAND U2075 ( .A(n843), .B(n845), .Z(n11415) );
  XOR U2076 ( .A(n11867), .B(n11868), .Z(n846) );
  NANDN U2077 ( .A(n11869), .B(n846), .Z(n847) );
  NAND U2078 ( .A(n11867), .B(n11868), .Z(n848) );
  AND U2079 ( .A(n847), .B(n848), .Z(n12025) );
  XOR U2080 ( .A(n12200), .B(n12199), .Z(n849) );
  NANDN U2081 ( .A(n12201), .B(n849), .Z(n850) );
  NAND U2082 ( .A(n12200), .B(n12199), .Z(n851) );
  AND U2083 ( .A(n850), .B(n851), .Z(n12377) );
  XOR U2084 ( .A(n6909), .B(n6910), .Z(n852) );
  NANDN U2085 ( .A(n6911), .B(n852), .Z(n853) );
  NAND U2086 ( .A(n6909), .B(n6910), .Z(n854) );
  AND U2087 ( .A(n853), .B(n854), .Z(n6938) );
  XOR U2088 ( .A(n7029), .B(n7030), .Z(n855) );
  NANDN U2089 ( .A(n7031), .B(n855), .Z(n856) );
  NAND U2090 ( .A(n7029), .B(n7030), .Z(n857) );
  AND U2091 ( .A(n856), .B(n857), .Z(n7047) );
  XOR U2092 ( .A(n7293), .B(n7294), .Z(n858) );
  NANDN U2093 ( .A(n7295), .B(n858), .Z(n859) );
  NAND U2094 ( .A(n7293), .B(n7294), .Z(n860) );
  AND U2095 ( .A(n859), .B(n860), .Z(n7311) );
  XOR U2096 ( .A(n7556), .B(n7557), .Z(n861) );
  NANDN U2097 ( .A(n7558), .B(n861), .Z(n862) );
  NAND U2098 ( .A(n7556), .B(n7557), .Z(n863) );
  AND U2099 ( .A(n862), .B(n863), .Z(n7573) );
  XOR U2100 ( .A(n7987), .B(n7988), .Z(n864) );
  NANDN U2101 ( .A(n7989), .B(n864), .Z(n865) );
  NAND U2102 ( .A(n7987), .B(n7988), .Z(n866) );
  AND U2103 ( .A(n865), .B(n866), .Z(n8111) );
  NAND U2104 ( .A(n8256), .B(n8257), .Z(n867) );
  XOR U2105 ( .A(n8256), .B(n8257), .Z(n868) );
  NAND U2106 ( .A(n868), .B(n8255), .Z(n869) );
  NAND U2107 ( .A(n867), .B(n869), .Z(n8513) );
  XOR U2108 ( .A(n8832), .B(n8833), .Z(n870) );
  NANDN U2109 ( .A(n8834), .B(n870), .Z(n871) );
  NAND U2110 ( .A(n8832), .B(n8833), .Z(n872) );
  AND U2111 ( .A(n871), .B(n872), .Z(n9128) );
  XOR U2112 ( .A(n3925), .B(n3926), .Z(n873) );
  NANDN U2113 ( .A(n3927), .B(n873), .Z(n874) );
  NAND U2114 ( .A(n3925), .B(n3926), .Z(n875) );
  AND U2115 ( .A(n874), .B(n875), .Z(n3958) );
  XOR U2116 ( .A(n4080), .B(n4081), .Z(n876) );
  NANDN U2117 ( .A(n4082), .B(n876), .Z(n877) );
  NAND U2118 ( .A(n4080), .B(n4081), .Z(n878) );
  AND U2119 ( .A(n877), .B(n878), .Z(n4098) );
  NAND U2120 ( .A(n4512), .B(n4513), .Z(n879) );
  XOR U2121 ( .A(n4512), .B(n4513), .Z(n880) );
  NANDN U2122 ( .A(n4511), .B(n880), .Z(n881) );
  NAND U2123 ( .A(n879), .B(n881), .Z(n4599) );
  NAND U2124 ( .A(n4803), .B(n4804), .Z(n882) );
  XOR U2125 ( .A(n4803), .B(n4804), .Z(n883) );
  NANDN U2126 ( .A(n4802), .B(n883), .Z(n884) );
  NAND U2127 ( .A(n882), .B(n884), .Z(n4914) );
  XOR U2128 ( .A(n5146), .B(n5147), .Z(n885) );
  NANDN U2129 ( .A(n5148), .B(n885), .Z(n886) );
  NAND U2130 ( .A(n5146), .B(n5147), .Z(n887) );
  AND U2131 ( .A(n886), .B(n887), .Z(n5273) );
  XOR U2132 ( .A(n5570), .B(n5571), .Z(n888) );
  NANDN U2133 ( .A(n5572), .B(n888), .Z(n889) );
  NAND U2134 ( .A(n5570), .B(n5571), .Z(n890) );
  AND U2135 ( .A(n889), .B(n890), .Z(n5847) );
  NAND U2136 ( .A(n6353), .B(n6354), .Z(n891) );
  XOR U2137 ( .A(n6353), .B(n6354), .Z(n892) );
  NANDN U2138 ( .A(n6352), .B(n892), .Z(n893) );
  NAND U2139 ( .A(n891), .B(n893), .Z(n6810) );
  NAND U2140 ( .A(n1095), .B(n1094), .Z(n894) );
  XOR U2141 ( .A(n1095), .B(n1094), .Z(n895) );
  NANDN U2142 ( .A(n1096), .B(n895), .Z(n896) );
  NAND U2143 ( .A(n894), .B(n896), .Z(n1131) );
  XOR U2144 ( .A(n1195), .B(n1196), .Z(n897) );
  NANDN U2145 ( .A(n1197), .B(n897), .Z(n898) );
  NAND U2146 ( .A(n1195), .B(n1196), .Z(n899) );
  AND U2147 ( .A(n898), .B(n899), .Z(n1295) );
  NAND U2148 ( .A(n1520), .B(n1521), .Z(n900) );
  XOR U2149 ( .A(n1520), .B(n1521), .Z(n901) );
  NANDN U2150 ( .A(n1519), .B(n901), .Z(n902) );
  NAND U2151 ( .A(n900), .B(n902), .Z(n1605) );
  NAND U2152 ( .A(n1803), .B(n1804), .Z(n903) );
  XOR U2153 ( .A(n1803), .B(n1804), .Z(n904) );
  NANDN U2154 ( .A(n1802), .B(n904), .Z(n905) );
  NAND U2155 ( .A(n903), .B(n905), .Z(n1900) );
  XOR U2156 ( .A(n2032), .B(n2033), .Z(n906) );
  NANDN U2157 ( .A(n2034), .B(n906), .Z(n907) );
  NAND U2158 ( .A(n2032), .B(n2033), .Z(n908) );
  AND U2159 ( .A(n907), .B(n908), .Z(n2252) );
  NAND U2160 ( .A(n2783), .B(n2784), .Z(n909) );
  XOR U2161 ( .A(n2783), .B(n2784), .Z(n910) );
  NANDN U2162 ( .A(n2782), .B(n910), .Z(n911) );
  NAND U2163 ( .A(n909), .B(n911), .Z(n2931) );
  XOR U2164 ( .A(n3099), .B(n3098), .Z(n912) );
  NANDN U2165 ( .A(n3100), .B(n912), .Z(n913) );
  NAND U2166 ( .A(n3099), .B(n3098), .Z(n914) );
  AND U2167 ( .A(n913), .B(n914), .Z(n3408) );
  NAND U2168 ( .A(n21184), .B(n21183), .Z(n915) );
  NANDN U2169 ( .A(n21186), .B(n21185), .Z(n916) );
  AND U2170 ( .A(n915), .B(n916), .Z(n917) );
  NAND U2171 ( .A(n20941), .B(n20940), .Z(n918) );
  NANDN U2172 ( .A(n20942), .B(n20943), .Z(n919) );
  AND U2173 ( .A(n918), .B(n919), .Z(n920) );
  XOR U2174 ( .A(n21182), .B(n21181), .Z(n921) );
  XNOR U2175 ( .A(n21169), .B(n21168), .Z(n922) );
  XNOR U2176 ( .A(n921), .B(n922), .Z(n923) );
  NAND U2177 ( .A(n21187), .B(n21188), .Z(n924) );
  NANDN U2178 ( .A(n21189), .B(n21190), .Z(n925) );
  AND U2179 ( .A(n924), .B(n925), .Z(n926) );
  NAND U2180 ( .A(n21193), .B(n21194), .Z(n927) );
  NAND U2181 ( .A(n21191), .B(n21192), .Z(n928) );
  AND U2182 ( .A(n927), .B(n928), .Z(n929) );
  XOR U2183 ( .A(n926), .B(n929), .Z(n930) );
  XNOR U2184 ( .A(n920), .B(n923), .Z(n931) );
  XNOR U2185 ( .A(n930), .B(n931), .Z(n932) );
  XNOR U2186 ( .A(n917), .B(n932), .Z(N448) );
  NAND U2187 ( .A(n9465), .B(n9466), .Z(n933) );
  NANDN U2188 ( .A(n9468), .B(n9467), .Z(n934) );
  AND U2189 ( .A(n933), .B(n934), .Z(n935) );
  NAND U2190 ( .A(n9469), .B(n9470), .Z(n936) );
  NANDN U2191 ( .A(n9471), .B(n9472), .Z(n937) );
  AND U2192 ( .A(n936), .B(n937), .Z(n938) );
  XOR U2193 ( .A(n9714), .B(n9713), .Z(n939) );
  XNOR U2194 ( .A(n9700), .B(n9699), .Z(n940) );
  XNOR U2195 ( .A(n939), .B(n940), .Z(n941) );
  AND U2196 ( .A(n9726), .B(n9725), .Z(n942) );
  NAND U2197 ( .A(n9720), .B(n9719), .Z(n943) );
  XNOR U2198 ( .A(n942), .B(n943), .Z(n944) );
  XOR U2199 ( .A(n941), .B(n944), .Z(n945) );
  XNOR U2200 ( .A(n935), .B(n938), .Z(n946) );
  XNOR U2201 ( .A(n945), .B(n946), .Z(n947) );
  NAND U2202 ( .A(n9727), .B(n9728), .Z(n948) );
  NANDN U2203 ( .A(n9730), .B(n9729), .Z(n949) );
  NAND U2204 ( .A(n948), .B(n949), .Z(n950) );
  XNOR U2205 ( .A(n947), .B(n950), .Z(N192) );
  NAND U2206 ( .A(n3592), .B(n3591), .Z(n951) );
  NANDN U2207 ( .A(n3594), .B(n3593), .Z(n952) );
  AND U2208 ( .A(n951), .B(n952), .Z(n953) );
  XOR U2209 ( .A(n3862), .B(n3861), .Z(n954) );
  XNOR U2210 ( .A(n3848), .B(n3847), .Z(n955) );
  XNOR U2211 ( .A(n954), .B(n955), .Z(n956) );
  NAND U2212 ( .A(n3864), .B(n3863), .Z(n957) );
  NANDN U2213 ( .A(n3866), .B(n3865), .Z(n958) );
  AND U2214 ( .A(n957), .B(n958), .Z(n959) );
  NAND U2215 ( .A(n3870), .B(n3869), .Z(n960) );
  NANDN U2216 ( .A(n3868), .B(n3867), .Z(n961) );
  AND U2217 ( .A(n960), .B(n961), .Z(n962) );
  XOR U2218 ( .A(n959), .B(n962), .Z(n963) );
  XNOR U2219 ( .A(n953), .B(n956), .Z(n964) );
  XNOR U2220 ( .A(n963), .B(n964), .Z(n965) );
  NAND U2221 ( .A(n3589), .B(n3590), .Z(n966) );
  NAND U2222 ( .A(n3587), .B(n3588), .Z(n967) );
  NAND U2223 ( .A(n966), .B(n967), .Z(n968) );
  XNOR U2224 ( .A(n965), .B(n968), .Z(N64) );
  AND U2225 ( .A(x[224]), .B(y[1792]), .Z(n1633) );
  XOR U2226 ( .A(n1633), .B(o[0]), .Z(N33) );
  AND U2227 ( .A(y[1792]), .B(x[225]), .Z(n970) );
  IV U2228 ( .A(n970), .Z(n978) );
  AND U2229 ( .A(x[224]), .B(y[1793]), .Z(n975) );
  XNOR U2230 ( .A(n975), .B(o[1]), .Z(n969) );
  XOR U2231 ( .A(n978), .B(n969), .Z(n972) );
  NAND U2232 ( .A(n1633), .B(o[0]), .Z(n971) );
  XNOR U2233 ( .A(n972), .B(n971), .Z(N34) );
  NANDN U2234 ( .A(n970), .B(n969), .Z(n974) );
  NAND U2235 ( .A(n972), .B(n971), .Z(n973) );
  AND U2236 ( .A(n974), .B(n973), .Z(n984) );
  AND U2237 ( .A(x[224]), .B(y[1794]), .Z(n989) );
  XNOR U2238 ( .A(n989), .B(o[2]), .Z(n983) );
  XNOR U2239 ( .A(n984), .B(n983), .Z(n986) );
  AND U2240 ( .A(n975), .B(o[1]), .Z(n980) );
  AND U2241 ( .A(x[225]), .B(y[1793]), .Z(n977) );
  NAND U2242 ( .A(x[226]), .B(y[1792]), .Z(n976) );
  XNOR U2243 ( .A(n977), .B(n976), .Z(n979) );
  XNOR U2244 ( .A(n980), .B(n979), .Z(n985) );
  XNOR U2245 ( .A(n986), .B(n985), .Z(N35) );
  AND U2246 ( .A(y[1793]), .B(x[226]), .Z(n1005) );
  NANDN U2247 ( .A(n978), .B(n1005), .Z(n982) );
  NAND U2248 ( .A(n980), .B(n979), .Z(n981) );
  AND U2249 ( .A(n982), .B(n981), .Z(n994) );
  NANDN U2250 ( .A(n984), .B(n983), .Z(n988) );
  NAND U2251 ( .A(n986), .B(n985), .Z(n987) );
  NAND U2252 ( .A(n988), .B(n987), .Z(n993) );
  AND U2253 ( .A(x[225]), .B(y[1794]), .Z(n1104) );
  XOR U2254 ( .A(n1005), .B(o[3]), .Z(n996) );
  XOR U2255 ( .A(n1104), .B(n996), .Z(n998) );
  AND U2256 ( .A(n989), .B(o[2]), .Z(n1002) );
  AND U2257 ( .A(x[227]), .B(y[1792]), .Z(n991) );
  NAND U2258 ( .A(y[1795]), .B(x[224]), .Z(n990) );
  XNOR U2259 ( .A(n991), .B(n990), .Z(n1001) );
  XOR U2260 ( .A(n1002), .B(n1001), .Z(n997) );
  XOR U2261 ( .A(n998), .B(n997), .Z(n995) );
  XOR U2262 ( .A(n993), .B(n995), .Z(n992) );
  XOR U2263 ( .A(n994), .B(n992), .Z(N36) );
  NAND U2264 ( .A(n1104), .B(n996), .Z(n1000) );
  NAND U2265 ( .A(n998), .B(n997), .Z(n999) );
  AND U2266 ( .A(n1000), .B(n999), .Z(n1015) );
  XNOR U2267 ( .A(n1016), .B(n1015), .Z(n1018) );
  AND U2268 ( .A(x[227]), .B(y[1795]), .Z(n1052) );
  NAND U2269 ( .A(n1633), .B(n1052), .Z(n1004) );
  NAND U2270 ( .A(n1002), .B(n1001), .Z(n1003) );
  NAND U2271 ( .A(n1004), .B(n1003), .Z(n1011) );
  AND U2272 ( .A(n1005), .B(o[3]), .Z(n1031) );
  AND U2273 ( .A(y[1796]), .B(x[224]), .Z(n1007) );
  AND U2274 ( .A(y[1792]), .B(x[228]), .Z(n1006) );
  XOR U2275 ( .A(n1007), .B(n1006), .Z(n1030) );
  XOR U2276 ( .A(n1031), .B(n1030), .Z(n1010) );
  AND U2277 ( .A(x[226]), .B(y[1794]), .Z(n1159) );
  NAND U2278 ( .A(y[1795]), .B(x[225]), .Z(n1008) );
  XNOR U2279 ( .A(n1159), .B(n1008), .Z(n1027) );
  AND U2280 ( .A(y[1793]), .B(x[227]), .Z(n1025) );
  XOR U2281 ( .A(n1025), .B(o[4]), .Z(n1026) );
  XOR U2282 ( .A(n1027), .B(n1026), .Z(n1009) );
  XNOR U2283 ( .A(n1010), .B(n1009), .Z(n1012) );
  XOR U2284 ( .A(n1011), .B(n1012), .Z(n1017) );
  XNOR U2285 ( .A(n1018), .B(n1017), .Z(N37) );
  NAND U2286 ( .A(n1010), .B(n1009), .Z(n1014) );
  NANDN U2287 ( .A(n1012), .B(n1011), .Z(n1013) );
  AND U2288 ( .A(n1014), .B(n1013), .Z(n1055) );
  NANDN U2289 ( .A(n1016), .B(n1015), .Z(n1020) );
  NAND U2290 ( .A(n1018), .B(n1017), .Z(n1019) );
  NAND U2291 ( .A(n1020), .B(n1019), .Z(n1054) );
  AND U2292 ( .A(x[226]), .B(y[1795]), .Z(n1113) );
  AND U2293 ( .A(y[1794]), .B(x[227]), .Z(n1022) );
  NAND U2294 ( .A(y[1796]), .B(x[225]), .Z(n1021) );
  XNOR U2295 ( .A(n1022), .B(n1021), .Z(n1036) );
  AND U2296 ( .A(x[228]), .B(y[1793]), .Z(n1050) );
  XOR U2297 ( .A(o[5]), .B(n1050), .Z(n1035) );
  XOR U2298 ( .A(n1036), .B(n1035), .Z(n1039) );
  XOR U2299 ( .A(n1113), .B(n1039), .Z(n1041) );
  AND U2300 ( .A(x[229]), .B(y[1792]), .Z(n1024) );
  NAND U2301 ( .A(y[1797]), .B(x[224]), .Z(n1023) );
  XNOR U2302 ( .A(n1024), .B(n1023), .Z(n1044) );
  AND U2303 ( .A(n1025), .B(o[4]), .Z(n1045) );
  XOR U2304 ( .A(n1044), .B(n1045), .Z(n1040) );
  XOR U2305 ( .A(n1041), .B(n1040), .Z(n1059) );
  NAND U2306 ( .A(n1113), .B(n1104), .Z(n1029) );
  NAND U2307 ( .A(n1027), .B(n1026), .Z(n1028) );
  NAND U2308 ( .A(n1029), .B(n1028), .Z(n1058) );
  AND U2309 ( .A(x[228]), .B(y[1796]), .Z(n1822) );
  NAND U2310 ( .A(n1822), .B(n1633), .Z(n1033) );
  NAND U2311 ( .A(n1031), .B(n1030), .Z(n1032) );
  NAND U2312 ( .A(n1033), .B(n1032), .Z(n1057) );
  XNOR U2313 ( .A(n1058), .B(n1057), .Z(n1060) );
  XOR U2314 ( .A(n1054), .B(n1056), .Z(n1034) );
  XOR U2315 ( .A(n1055), .B(n1034), .Z(N38) );
  AND U2316 ( .A(x[227]), .B(y[1796]), .Z(n1114) );
  NAND U2317 ( .A(n1114), .B(n1104), .Z(n1038) );
  NAND U2318 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U2319 ( .A(n1038), .B(n1037), .Z(n1089) );
  NAND U2320 ( .A(n1113), .B(n1039), .Z(n1043) );
  NAND U2321 ( .A(n1041), .B(n1040), .Z(n1042) );
  NAND U2322 ( .A(n1043), .B(n1042), .Z(n1088) );
  AND U2323 ( .A(y[1797]), .B(x[229]), .Z(n1283) );
  NAND U2324 ( .A(n1633), .B(n1283), .Z(n1047) );
  NAND U2325 ( .A(n1045), .B(n1044), .Z(n1046) );
  NAND U2326 ( .A(n1047), .B(n1046), .Z(n1065) );
  AND U2327 ( .A(x[230]), .B(y[1792]), .Z(n1049) );
  NAND U2328 ( .A(x[224]), .B(y[1798]), .Z(n1048) );
  XNOR U2329 ( .A(n1049), .B(n1048), .Z(n1072) );
  AND U2330 ( .A(o[5]), .B(n1050), .Z(n1071) );
  XOR U2331 ( .A(n1072), .B(n1071), .Z(n1064) );
  XOR U2332 ( .A(n1065), .B(n1064), .Z(n1067) );
  NAND U2333 ( .A(y[1796]), .B(x[226]), .Z(n1051) );
  XNOR U2334 ( .A(n1052), .B(n1051), .Z(n1076) );
  AND U2335 ( .A(y[1797]), .B(x[225]), .Z(n1317) );
  NAND U2336 ( .A(y[1794]), .B(x[228]), .Z(n1053) );
  XNOR U2337 ( .A(n1317), .B(n1053), .Z(n1080) );
  AND U2338 ( .A(y[1793]), .B(x[229]), .Z(n1087) );
  XOR U2339 ( .A(o[6]), .B(n1087), .Z(n1079) );
  XOR U2340 ( .A(n1080), .B(n1079), .Z(n1075) );
  XOR U2341 ( .A(n1076), .B(n1075), .Z(n1066) );
  XOR U2342 ( .A(n1067), .B(n1066), .Z(n1090) );
  XNOR U2343 ( .A(n1091), .B(n1090), .Z(n1096) );
  NAND U2344 ( .A(n1058), .B(n1057), .Z(n1062) );
  NANDN U2345 ( .A(n1060), .B(n1059), .Z(n1061) );
  NAND U2346 ( .A(n1062), .B(n1061), .Z(n1094) );
  XOR U2347 ( .A(n1095), .B(n1094), .Z(n1063) );
  XNOR U2348 ( .A(n1096), .B(n1063), .Z(N39) );
  NAND U2349 ( .A(n1065), .B(n1064), .Z(n1069) );
  NAND U2350 ( .A(n1067), .B(n1066), .Z(n1068) );
  AND U2351 ( .A(n1069), .B(n1068), .Z(n1136) );
  AND U2352 ( .A(y[1794]), .B(x[229]), .Z(n1204) );
  NAND U2353 ( .A(x[225]), .B(y[1798]), .Z(n1070) );
  XNOR U2354 ( .A(n1204), .B(n1070), .Z(n1107) );
  AND U2355 ( .A(y[1793]), .B(x[230]), .Z(n1110) );
  XOR U2356 ( .A(o[7]), .B(n1110), .Z(n1106) );
  XNOR U2357 ( .A(n1107), .B(n1106), .Z(n1125) );
  AND U2358 ( .A(y[1798]), .B(x[230]), .Z(n1336) );
  NAND U2359 ( .A(n1633), .B(n1336), .Z(n1074) );
  NAND U2360 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U2361 ( .A(n1074), .B(n1073), .Z(n1124) );
  XOR U2362 ( .A(n1125), .B(n1124), .Z(n1126) );
  NAND U2363 ( .A(n1113), .B(n1114), .Z(n1078) );
  NAND U2364 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U2365 ( .A(n1078), .B(n1077), .Z(n1127) );
  XOR U2366 ( .A(n1126), .B(n1127), .Z(n1134) );
  AND U2367 ( .A(x[228]), .B(y[1797]), .Z(n1638) );
  NAND U2368 ( .A(n1638), .B(n1104), .Z(n1082) );
  NAND U2369 ( .A(n1080), .B(n1079), .Z(n1081) );
  AND U2370 ( .A(n1082), .B(n1081), .Z(n1101) );
  AND U2371 ( .A(y[1797]), .B(x[226]), .Z(n1084) );
  NAND U2372 ( .A(y[1795]), .B(x[228]), .Z(n1083) );
  XNOR U2373 ( .A(n1084), .B(n1083), .Z(n1115) );
  XNOR U2374 ( .A(n1115), .B(n1114), .Z(n1099) );
  AND U2375 ( .A(x[231]), .B(y[1792]), .Z(n1086) );
  NAND U2376 ( .A(y[1799]), .B(x[224]), .Z(n1085) );
  XNOR U2377 ( .A(n1086), .B(n1085), .Z(n1119) );
  AND U2378 ( .A(o[6]), .B(n1087), .Z(n1118) );
  XNOR U2379 ( .A(n1119), .B(n1118), .Z(n1098) );
  XOR U2380 ( .A(n1099), .B(n1098), .Z(n1100) );
  XOR U2381 ( .A(n1101), .B(n1100), .Z(n1133) );
  XOR U2382 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U2383 ( .A(n1136), .B(n1135), .Z(n1132) );
  NANDN U2384 ( .A(n1089), .B(n1088), .Z(n1093) );
  NAND U2385 ( .A(n1091), .B(n1090), .Z(n1092) );
  NAND U2386 ( .A(n1093), .B(n1092), .Z(n1130) );
  XOR U2387 ( .A(n1130), .B(n1131), .Z(n1097) );
  XNOR U2388 ( .A(n1132), .B(n1097), .Z(N40) );
  NAND U2389 ( .A(n1099), .B(n1098), .Z(n1103) );
  NAND U2390 ( .A(n1101), .B(n1100), .Z(n1102) );
  AND U2391 ( .A(n1103), .B(n1102), .Z(n1172) );
  AND U2392 ( .A(y[1798]), .B(x[229]), .Z(n1105) );
  NAND U2393 ( .A(n1105), .B(n1104), .Z(n1109) );
  NAND U2394 ( .A(n1107), .B(n1106), .Z(n1108) );
  AND U2395 ( .A(n1109), .B(n1108), .Z(n1170) );
  AND U2396 ( .A(o[7]), .B(n1110), .Z(n1150) );
  AND U2397 ( .A(x[229]), .B(y[1795]), .Z(n1729) );
  NAND U2398 ( .A(y[1799]), .B(x[225]), .Z(n1111) );
  XNOR U2399 ( .A(n1729), .B(n1111), .Z(n1151) );
  XNOR U2400 ( .A(n1150), .B(n1151), .Z(n1155) );
  NAND U2401 ( .A(x[227]), .B(y[1797]), .Z(n1958) );
  AND U2402 ( .A(y[1794]), .B(x[230]), .Z(n1112) );
  AND U2403 ( .A(x[226]), .B(y[1798]), .Z(n2102) );
  XOR U2404 ( .A(n1112), .B(n2102), .Z(n1160) );
  XOR U2405 ( .A(n1822), .B(n1160), .Z(n1154) );
  XOR U2406 ( .A(n1155), .B(n1156), .Z(n1169) );
  XOR U2407 ( .A(n1172), .B(n1171), .Z(n1185) );
  NAND U2408 ( .A(n1638), .B(n1113), .Z(n1117) );
  NAND U2409 ( .A(n1115), .B(n1114), .Z(n1116) );
  AND U2410 ( .A(n1117), .B(n1116), .Z(n1166) );
  AND U2411 ( .A(y[1799]), .B(x[231]), .Z(n1490) );
  NAND U2412 ( .A(n1633), .B(n1490), .Z(n1121) );
  NAND U2413 ( .A(n1119), .B(n1118), .Z(n1120) );
  AND U2414 ( .A(n1121), .B(n1120), .Z(n1164) );
  AND U2415 ( .A(x[232]), .B(y[1792]), .Z(n1123) );
  NAND U2416 ( .A(y[1800]), .B(x[224]), .Z(n1122) );
  XNOR U2417 ( .A(n1123), .B(n1122), .Z(n1142) );
  AND U2418 ( .A(y[1793]), .B(x[231]), .Z(n1146) );
  XOR U2419 ( .A(o[8]), .B(n1146), .Z(n1141) );
  XOR U2420 ( .A(n1142), .B(n1141), .Z(n1163) );
  NAND U2421 ( .A(n1125), .B(n1124), .Z(n1129) );
  NAND U2422 ( .A(n1127), .B(n1126), .Z(n1128) );
  NAND U2423 ( .A(n1129), .B(n1128), .Z(n1182) );
  XOR U2424 ( .A(n1183), .B(n1182), .Z(n1184) );
  XOR U2425 ( .A(n1185), .B(n1184), .Z(n1178) );
  NAND U2426 ( .A(n1134), .B(n1133), .Z(n1138) );
  NAND U2427 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U2428 ( .A(n1138), .B(n1137), .Z(n1177) );
  IV U2429 ( .A(n1177), .Z(n1175) );
  XOR U2430 ( .A(n1176), .B(n1175), .Z(n1139) );
  XNOR U2431 ( .A(n1178), .B(n1139), .Z(N41) );
  AND U2432 ( .A(x[232]), .B(y[1800]), .Z(n1140) );
  NAND U2433 ( .A(n1140), .B(n1633), .Z(n1144) );
  NAND U2434 ( .A(n1142), .B(n1141), .Z(n1143) );
  AND U2435 ( .A(n1144), .B(n1143), .Z(n1234) );
  AND U2436 ( .A(y[1794]), .B(x[231]), .Z(n1553) );
  NAND U2437 ( .A(x[229]), .B(y[1796]), .Z(n1145) );
  XNOR U2438 ( .A(n1553), .B(n1145), .Z(n1206) );
  AND U2439 ( .A(o[8]), .B(n1146), .Z(n1205) );
  XNOR U2440 ( .A(n1206), .B(n1205), .Z(n1232) );
  AND U2441 ( .A(x[233]), .B(y[1792]), .Z(n1148) );
  NAND U2442 ( .A(y[1801]), .B(x[224]), .Z(n1147) );
  XNOR U2443 ( .A(n1148), .B(n1147), .Z(n1213) );
  AND U2444 ( .A(y[1793]), .B(x[232]), .Z(n1223) );
  XOR U2445 ( .A(o[9]), .B(n1223), .Z(n1212) );
  XNOR U2446 ( .A(n1213), .B(n1212), .Z(n1231) );
  XOR U2447 ( .A(n1232), .B(n1231), .Z(n1233) );
  XNOR U2448 ( .A(n1234), .B(n1233), .Z(n1228) );
  AND U2449 ( .A(x[230]), .B(y[1795]), .Z(n1567) );
  NAND U2450 ( .A(y[1800]), .B(x[225]), .Z(n1149) );
  XNOR U2451 ( .A(n1567), .B(n1149), .Z(n1218) );
  XNOR U2452 ( .A(n1638), .B(n1218), .Z(n1238) );
  AND U2453 ( .A(y[1799]), .B(x[226]), .Z(n1869) );
  NAND U2454 ( .A(y[1798]), .B(x[227]), .Z(n1578) );
  XNOR U2455 ( .A(n1869), .B(n1578), .Z(n1237) );
  XNOR U2456 ( .A(n1238), .B(n1237), .Z(n1226) );
  NAND U2457 ( .A(y[1799]), .B(x[229]), .Z(n1403) );
  AND U2458 ( .A(x[225]), .B(y[1795]), .Z(n1216) );
  NANDN U2459 ( .A(n1403), .B(n1216), .Z(n1153) );
  NAND U2460 ( .A(n1151), .B(n1150), .Z(n1152) );
  NAND U2461 ( .A(n1153), .B(n1152), .Z(n1225) );
  XOR U2462 ( .A(n1226), .B(n1225), .Z(n1227) );
  XNOR U2463 ( .A(n1228), .B(n1227), .Z(n1200) );
  NANDN U2464 ( .A(n1154), .B(n1958), .Z(n1158) );
  NANDN U2465 ( .A(n1156), .B(n1155), .Z(n1157) );
  NAND U2466 ( .A(n1158), .B(n1157), .Z(n1198) );
  NAND U2467 ( .A(n1336), .B(n1159), .Z(n1162) );
  NAND U2468 ( .A(n1822), .B(n1160), .Z(n1161) );
  AND U2469 ( .A(n1162), .B(n1161), .Z(n1199) );
  XNOR U2470 ( .A(n1198), .B(n1199), .Z(n1201) );
  NANDN U2471 ( .A(n1164), .B(n1163), .Z(n1168) );
  NANDN U2472 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U2473 ( .A(n1168), .B(n1167), .Z(n1190) );
  NANDN U2474 ( .A(n1170), .B(n1169), .Z(n1174) );
  NAND U2475 ( .A(n1172), .B(n1171), .Z(n1173) );
  NAND U2476 ( .A(n1174), .B(n1173), .Z(n1189) );
  XNOR U2477 ( .A(n1191), .B(n1192), .Z(n1197) );
  NANDN U2478 ( .A(n1175), .B(n1176), .Z(n1181) );
  NOR U2479 ( .A(n1177), .B(n1176), .Z(n1179) );
  OR U2480 ( .A(n1179), .B(n1178), .Z(n1180) );
  AND U2481 ( .A(n1181), .B(n1180), .Z(n1195) );
  NAND U2482 ( .A(n1183), .B(n1182), .Z(n1187) );
  NANDN U2483 ( .A(n1185), .B(n1184), .Z(n1186) );
  AND U2484 ( .A(n1187), .B(n1186), .Z(n1196) );
  XOR U2485 ( .A(n1195), .B(n1196), .Z(n1188) );
  XNOR U2486 ( .A(n1197), .B(n1188), .Z(N42) );
  NANDN U2487 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U2488 ( .A(n1192), .B(n1191), .Z(n1193) );
  NAND U2489 ( .A(n1194), .B(n1193), .Z(n1294) );
  IV U2490 ( .A(n1294), .Z(n1293) );
  NAND U2491 ( .A(n1199), .B(n1198), .Z(n1203) );
  NANDN U2492 ( .A(n1201), .B(n1200), .Z(n1202) );
  NAND U2493 ( .A(n1203), .B(n1202), .Z(n1302) );
  AND U2494 ( .A(y[1796]), .B(x[231]), .Z(n1277) );
  NAND U2495 ( .A(n1277), .B(n1204), .Z(n1208) );
  NAND U2496 ( .A(n1206), .B(n1205), .Z(n1207) );
  AND U2497 ( .A(n1208), .B(n1207), .Z(n1290) );
  AND U2498 ( .A(x[231]), .B(y[1795]), .Z(n1210) );
  NAND U2499 ( .A(x[228]), .B(y[1798]), .Z(n1209) );
  XNOR U2500 ( .A(n1210), .B(n1209), .Z(n1261) );
  AND U2501 ( .A(y[1796]), .B(x[230]), .Z(n1260) );
  XOR U2502 ( .A(n1261), .B(n1260), .Z(n1288) );
  AND U2503 ( .A(x[232]), .B(y[1794]), .Z(n1464) );
  AND U2504 ( .A(y[1793]), .B(x[233]), .Z(n1269) );
  XOR U2505 ( .A(o[10]), .B(n1269), .Z(n1282) );
  XOR U2506 ( .A(n1464), .B(n1282), .Z(n1284) );
  XNOR U2507 ( .A(n1284), .B(n1283), .Z(n1287) );
  XNOR U2508 ( .A(n1290), .B(n1289), .Z(n1249) );
  AND U2509 ( .A(x[233]), .B(y[1801]), .Z(n1211) );
  NAND U2510 ( .A(n1211), .B(n1633), .Z(n1215) );
  NAND U2511 ( .A(n1213), .B(n1212), .Z(n1214) );
  NAND U2512 ( .A(n1215), .B(n1214), .Z(n1247) );
  AND U2513 ( .A(y[1800]), .B(x[230]), .Z(n1217) );
  NAND U2514 ( .A(n1217), .B(n1216), .Z(n1220) );
  NAND U2515 ( .A(n1638), .B(n1218), .Z(n1219) );
  NAND U2516 ( .A(n1220), .B(n1219), .Z(n1255) );
  AND U2517 ( .A(x[234]), .B(y[1792]), .Z(n1222) );
  NAND U2518 ( .A(y[1802]), .B(x[224]), .Z(n1221) );
  XNOR U2519 ( .A(n1222), .B(n1221), .Z(n1266) );
  AND U2520 ( .A(o[9]), .B(n1223), .Z(n1265) );
  XOR U2521 ( .A(n1266), .B(n1265), .Z(n1253) );
  AND U2522 ( .A(x[227]), .B(y[1799]), .Z(n2192) );
  NAND U2523 ( .A(y[1801]), .B(x[225]), .Z(n1224) );
  XNOR U2524 ( .A(n2192), .B(n1224), .Z(n1278) );
  AND U2525 ( .A(y[1800]), .B(x[226]), .Z(n1279) );
  XOR U2526 ( .A(n1278), .B(n1279), .Z(n1252) );
  XOR U2527 ( .A(n1253), .B(n1252), .Z(n1254) );
  XOR U2528 ( .A(n1255), .B(n1254), .Z(n1246) );
  XOR U2529 ( .A(n1247), .B(n1246), .Z(n1248) );
  XOR U2530 ( .A(n1249), .B(n1248), .Z(n1301) );
  NAND U2531 ( .A(n1226), .B(n1225), .Z(n1230) );
  NAND U2532 ( .A(n1228), .B(n1227), .Z(n1229) );
  AND U2533 ( .A(n1230), .B(n1229), .Z(n1243) );
  NAND U2534 ( .A(n1232), .B(n1231), .Z(n1236) );
  NAND U2535 ( .A(n1234), .B(n1233), .Z(n1235) );
  AND U2536 ( .A(n1236), .B(n1235), .Z(n1240) );
  XOR U2537 ( .A(n1240), .B(n1241), .Z(n1242) );
  XOR U2538 ( .A(n1243), .B(n1242), .Z(n1300) );
  XOR U2539 ( .A(n1302), .B(n1303), .Z(n1296) );
  XNOR U2540 ( .A(n1295), .B(n1296), .Z(n1239) );
  XOR U2541 ( .A(n1293), .B(n1239), .Z(N43) );
  NAND U2542 ( .A(n1241), .B(n1240), .Z(n1245) );
  NANDN U2543 ( .A(n1243), .B(n1242), .Z(n1244) );
  AND U2544 ( .A(n1245), .B(n1244), .Z(n1371) );
  NAND U2545 ( .A(n1247), .B(n1246), .Z(n1251) );
  NAND U2546 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U2547 ( .A(n1251), .B(n1250), .Z(n1369) );
  NAND U2548 ( .A(n1253), .B(n1252), .Z(n1257) );
  NAND U2549 ( .A(n1255), .B(n1254), .Z(n1256) );
  NAND U2550 ( .A(n1257), .B(n1256), .Z(n1358) );
  AND U2551 ( .A(y[1798]), .B(x[231]), .Z(n1259) );
  AND U2552 ( .A(x[228]), .B(y[1795]), .Z(n1258) );
  NAND U2553 ( .A(n1259), .B(n1258), .Z(n1263) );
  NAND U2554 ( .A(n1261), .B(n1260), .Z(n1262) );
  NAND U2555 ( .A(n1263), .B(n1262), .Z(n1356) );
  AND U2556 ( .A(x[234]), .B(y[1802]), .Z(n1264) );
  NAND U2557 ( .A(n1264), .B(n1633), .Z(n1268) );
  NAND U2558 ( .A(n1266), .B(n1265), .Z(n1267) );
  NAND U2559 ( .A(n1268), .B(n1267), .Z(n1352) );
  AND U2560 ( .A(o[10]), .B(n1269), .Z(n1327) );
  AND U2561 ( .A(x[235]), .B(y[1792]), .Z(n1271) );
  NAND U2562 ( .A(x[224]), .B(y[1803]), .Z(n1270) );
  XNOR U2563 ( .A(n1271), .B(n1270), .Z(n1328) );
  XOR U2564 ( .A(n1327), .B(n1328), .Z(n1350) );
  AND U2565 ( .A(x[230]), .B(y[1797]), .Z(n1273) );
  NAND U2566 ( .A(y[1802]), .B(x[225]), .Z(n1272) );
  XNOR U2567 ( .A(n1273), .B(n1272), .Z(n1319) );
  AND U2568 ( .A(y[1793]), .B(x[234]), .Z(n1337) );
  XOR U2569 ( .A(o[11]), .B(n1337), .Z(n1318) );
  XOR U2570 ( .A(n1319), .B(n1318), .Z(n1349) );
  XOR U2571 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U2572 ( .A(n1352), .B(n1351), .Z(n1355) );
  XOR U2573 ( .A(n1356), .B(n1355), .Z(n1357) );
  XNOR U2574 ( .A(n1358), .B(n1357), .Z(n1340) );
  NAND U2575 ( .A(y[1800]), .B(x[227]), .Z(n2321) );
  AND U2576 ( .A(x[226]), .B(y[1801]), .Z(n1275) );
  NAND U2577 ( .A(x[229]), .B(y[1798]), .Z(n1274) );
  XNOR U2578 ( .A(n1275), .B(n1274), .Z(n1314) );
  AND U2579 ( .A(x[228]), .B(y[1799]), .Z(n1313) );
  XNOR U2580 ( .A(n1314), .B(n1313), .Z(n1344) );
  XOR U2581 ( .A(n2321), .B(n1344), .Z(n1346) );
  NAND U2582 ( .A(y[1794]), .B(x[233]), .Z(n1276) );
  XNOR U2583 ( .A(n1277), .B(n1276), .Z(n1332) );
  AND U2584 ( .A(x[232]), .B(y[1795]), .Z(n1331) );
  XNOR U2585 ( .A(n1332), .B(n1331), .Z(n1345) );
  XNOR U2586 ( .A(n1346), .B(n1345), .Z(n1310) );
  NAND U2587 ( .A(y[1801]), .B(x[227]), .Z(n1394) );
  AND U2588 ( .A(x[225]), .B(y[1799]), .Z(n1628) );
  NANDN U2589 ( .A(n1394), .B(n1628), .Z(n1281) );
  NAND U2590 ( .A(n1279), .B(n1278), .Z(n1280) );
  NAND U2591 ( .A(n1281), .B(n1280), .Z(n1308) );
  NAND U2592 ( .A(n1464), .B(n1282), .Z(n1286) );
  NAND U2593 ( .A(n1284), .B(n1283), .Z(n1285) );
  NAND U2594 ( .A(n1286), .B(n1285), .Z(n1307) );
  XOR U2595 ( .A(n1308), .B(n1307), .Z(n1309) );
  XNOR U2596 ( .A(n1310), .B(n1309), .Z(n1339) );
  NANDN U2597 ( .A(n1288), .B(n1287), .Z(n1292) );
  NAND U2598 ( .A(n1290), .B(n1289), .Z(n1291) );
  NAND U2599 ( .A(n1292), .B(n1291), .Z(n1338) );
  XOR U2600 ( .A(n1339), .B(n1338), .Z(n1341) );
  XNOR U2601 ( .A(n1340), .B(n1341), .Z(n1368) );
  XOR U2602 ( .A(n1369), .B(n1368), .Z(n1370) );
  XOR U2603 ( .A(n1371), .B(n1370), .Z(n1364) );
  OR U2604 ( .A(n1295), .B(n1293), .Z(n1299) );
  ANDN U2605 ( .B(n1295), .A(n1294), .Z(n1297) );
  OR U2606 ( .A(n1297), .B(n1296), .Z(n1298) );
  AND U2607 ( .A(n1299), .B(n1298), .Z(n1363) );
  NANDN U2608 ( .A(n1301), .B(n1300), .Z(n1305) );
  NAND U2609 ( .A(n1303), .B(n1302), .Z(n1304) );
  AND U2610 ( .A(n1305), .B(n1304), .Z(n1362) );
  IV U2611 ( .A(n1362), .Z(n1361) );
  XOR U2612 ( .A(n1363), .B(n1361), .Z(n1306) );
  XNOR U2613 ( .A(n1364), .B(n1306), .Z(N44) );
  NAND U2614 ( .A(n1308), .B(n1307), .Z(n1312) );
  NAND U2615 ( .A(n1310), .B(n1309), .Z(n1311) );
  NAND U2616 ( .A(n1312), .B(n1311), .Z(n1435) );
  AND U2617 ( .A(y[1801]), .B(x[229]), .Z(n1860) );
  NAND U2618 ( .A(n2102), .B(n1860), .Z(n1316) );
  NAND U2619 ( .A(n1314), .B(n1313), .Z(n1315) );
  NAND U2620 ( .A(n1316), .B(n1315), .Z(n1382) );
  AND U2621 ( .A(x[230]), .B(y[1802]), .Z(n1645) );
  NAND U2622 ( .A(n1645), .B(n1317), .Z(n1321) );
  NAND U2623 ( .A(n1319), .B(n1318), .Z(n1320) );
  NAND U2624 ( .A(n1321), .B(n1320), .Z(n1381) );
  XOR U2625 ( .A(n1382), .B(n1381), .Z(n1384) );
  AND U2626 ( .A(x[233]), .B(y[1795]), .Z(n2097) );
  AND U2627 ( .A(y[1794]), .B(x[234]), .Z(n2080) );
  AND U2628 ( .A(y[1800]), .B(x[228]), .Z(n1322) );
  XOR U2629 ( .A(n2080), .B(n1322), .Z(n1425) );
  XOR U2630 ( .A(n2097), .B(n1425), .Z(n1404) );
  NAND U2631 ( .A(x[231]), .B(y[1797]), .Z(n1402) );
  XOR U2632 ( .A(n1403), .B(n1402), .Z(n1405) );
  AND U2633 ( .A(x[236]), .B(y[1792]), .Z(n1324) );
  NAND U2634 ( .A(y[1804]), .B(x[224]), .Z(n1323) );
  XNOR U2635 ( .A(n1324), .B(n1323), .Z(n1419) );
  AND U2636 ( .A(y[1793]), .B(x[235]), .Z(n1399) );
  XOR U2637 ( .A(o[12]), .B(n1399), .Z(n1418) );
  XOR U2638 ( .A(n1419), .B(n1418), .Z(n1388) );
  AND U2639 ( .A(y[1802]), .B(x[226]), .Z(n1326) );
  NAND U2640 ( .A(y[1796]), .B(x[232]), .Z(n1325) );
  XNOR U2641 ( .A(n1326), .B(n1325), .Z(n1393) );
  XOR U2642 ( .A(n1388), .B(n1387), .Z(n1390) );
  XOR U2643 ( .A(n1389), .B(n1390), .Z(n1383) );
  XOR U2644 ( .A(n1384), .B(n1383), .Z(n1433) );
  AND U2645 ( .A(y[1803]), .B(x[235]), .Z(n2443) );
  NAND U2646 ( .A(n2443), .B(n1633), .Z(n1330) );
  NAND U2647 ( .A(n1328), .B(n1327), .Z(n1329) );
  NAND U2648 ( .A(n1330), .B(n1329), .Z(n1411) );
  AND U2649 ( .A(x[233]), .B(y[1796]), .Z(n1401) );
  NAND U2650 ( .A(n1553), .B(n1401), .Z(n1334) );
  NAND U2651 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U2652 ( .A(n1334), .B(n1333), .Z(n1409) );
  NAND U2653 ( .A(x[225]), .B(y[1803]), .Z(n1335) );
  XNOR U2654 ( .A(n1336), .B(n1335), .Z(n1415) );
  AND U2655 ( .A(o[11]), .B(n1337), .Z(n1414) );
  XOR U2656 ( .A(n1415), .B(n1414), .Z(n1408) );
  XOR U2657 ( .A(n1409), .B(n1408), .Z(n1410) );
  XOR U2658 ( .A(n1411), .B(n1410), .Z(n1432) );
  XOR U2659 ( .A(n1433), .B(n1432), .Z(n1434) );
  XNOR U2660 ( .A(n1435), .B(n1434), .Z(n1439) );
  NAND U2661 ( .A(n1339), .B(n1338), .Z(n1343) );
  NAND U2662 ( .A(n1341), .B(n1340), .Z(n1342) );
  NAND U2663 ( .A(n1343), .B(n1342), .Z(n1438) );
  XOR U2664 ( .A(n1439), .B(n1438), .Z(n1441) );
  IV U2665 ( .A(n2321), .Z(n2111) );
  NANDN U2666 ( .A(n2111), .B(n1344), .Z(n1348) );
  NAND U2667 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U2668 ( .A(n1348), .B(n1347), .Z(n1376) );
  NAND U2669 ( .A(n1350), .B(n1349), .Z(n1354) );
  NAND U2670 ( .A(n1352), .B(n1351), .Z(n1353) );
  AND U2671 ( .A(n1354), .B(n1353), .Z(n1375) );
  XOR U2672 ( .A(n1376), .B(n1375), .Z(n1377) );
  NAND U2673 ( .A(n1356), .B(n1355), .Z(n1360) );
  NAND U2674 ( .A(n1358), .B(n1357), .Z(n1359) );
  AND U2675 ( .A(n1360), .B(n1359), .Z(n1378) );
  XOR U2676 ( .A(n1377), .B(n1378), .Z(n1440) );
  XNOR U2677 ( .A(n1441), .B(n1440), .Z(n1447) );
  OR U2678 ( .A(n1363), .B(n1361), .Z(n1367) );
  ANDN U2679 ( .B(n1363), .A(n1362), .Z(n1365) );
  OR U2680 ( .A(n1365), .B(n1364), .Z(n1366) );
  AND U2681 ( .A(n1367), .B(n1366), .Z(n1445) );
  NAND U2682 ( .A(n1369), .B(n1368), .Z(n1373) );
  NANDN U2683 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U2684 ( .A(n1373), .B(n1372), .Z(n1446) );
  IV U2685 ( .A(n1446), .Z(n1444) );
  XOR U2686 ( .A(n1445), .B(n1444), .Z(n1374) );
  XNOR U2687 ( .A(n1447), .B(n1374), .Z(N45) );
  NAND U2688 ( .A(n1376), .B(n1375), .Z(n1380) );
  NAND U2689 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U2690 ( .A(n1380), .B(n1379), .Z(n1525) );
  NAND U2691 ( .A(n1382), .B(n1381), .Z(n1386) );
  NAND U2692 ( .A(n1384), .B(n1383), .Z(n1385) );
  NAND U2693 ( .A(n1386), .B(n1385), .Z(n1508) );
  NAND U2694 ( .A(n1388), .B(n1387), .Z(n1392) );
  NAND U2695 ( .A(n1390), .B(n1389), .Z(n1391) );
  NAND U2696 ( .A(n1392), .B(n1391), .Z(n1515) );
  AND U2697 ( .A(y[1802]), .B(x[232]), .Z(n2668) );
  AND U2698 ( .A(x[226]), .B(y[1796]), .Z(n1563) );
  NAND U2699 ( .A(n2668), .B(n1563), .Z(n1396) );
  NANDN U2700 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U2701 ( .A(n1396), .B(n1395), .Z(n1479) );
  AND U2702 ( .A(y[1804]), .B(x[225]), .Z(n1398) );
  NAND U2703 ( .A(x[231]), .B(y[1798]), .Z(n1397) );
  XNOR U2704 ( .A(n1398), .B(n1397), .Z(n1470) );
  AND U2705 ( .A(o[12]), .B(n1399), .Z(n1469) );
  XOR U2706 ( .A(n1470), .B(n1469), .Z(n1477) );
  AND U2707 ( .A(y[1799]), .B(x[230]), .Z(n2480) );
  NAND U2708 ( .A(x[226]), .B(y[1803]), .Z(n1400) );
  XNOR U2709 ( .A(n1401), .B(n1400), .Z(n1483) );
  XOR U2710 ( .A(n2480), .B(n1483), .Z(n1476) );
  XOR U2711 ( .A(n1477), .B(n1476), .Z(n1478) );
  XOR U2712 ( .A(n1479), .B(n1478), .Z(n1514) );
  NAND U2713 ( .A(n1403), .B(n1402), .Z(n1407) );
  ANDN U2714 ( .B(n1405), .A(n1404), .Z(n1406) );
  ANDN U2715 ( .B(n1407), .A(n1406), .Z(n1513) );
  XOR U2716 ( .A(n1514), .B(n1513), .Z(n1516) );
  XOR U2717 ( .A(n1515), .B(n1516), .Z(n1507) );
  XOR U2718 ( .A(n1508), .B(n1507), .Z(n1510) );
  NAND U2719 ( .A(n1409), .B(n1408), .Z(n1413) );
  NAND U2720 ( .A(n1411), .B(n1410), .Z(n1412) );
  NAND U2721 ( .A(n1413), .B(n1412), .Z(n1454) );
  AND U2722 ( .A(y[1803]), .B(x[230]), .Z(n1861) );
  AND U2723 ( .A(y[1798]), .B(x[225]), .Z(n1468) );
  NAND U2724 ( .A(n1861), .B(n1468), .Z(n1417) );
  NAND U2725 ( .A(n1415), .B(n1414), .Z(n1416) );
  NAND U2726 ( .A(n1417), .B(n1416), .Z(n1461) );
  AND U2727 ( .A(x[236]), .B(y[1804]), .Z(n2674) );
  NAND U2728 ( .A(n2674), .B(n1633), .Z(n1421) );
  NAND U2729 ( .A(n1419), .B(n1418), .Z(n1420) );
  NAND U2730 ( .A(n1421), .B(n1420), .Z(n1459) );
  AND U2731 ( .A(x[234]), .B(y[1795]), .Z(n2333) );
  AND U2732 ( .A(y[1794]), .B(x[235]), .Z(n2294) );
  NAND U2733 ( .A(y[1797]), .B(x[232]), .Z(n1422) );
  XNOR U2734 ( .A(n2294), .B(n1422), .Z(n1465) );
  XOR U2735 ( .A(n2333), .B(n1465), .Z(n1458) );
  XOR U2736 ( .A(n1459), .B(n1458), .Z(n1460) );
  XOR U2737 ( .A(n1461), .B(n1460), .Z(n1452) );
  AND U2738 ( .A(x[234]), .B(y[1800]), .Z(n1424) );
  AND U2739 ( .A(x[228]), .B(y[1794]), .Z(n1423) );
  NAND U2740 ( .A(n1424), .B(n1423), .Z(n1427) );
  NAND U2741 ( .A(n2097), .B(n1425), .Z(n1426) );
  NAND U2742 ( .A(n1427), .B(n1426), .Z(n1503) );
  AND U2743 ( .A(x[237]), .B(y[1792]), .Z(n1429) );
  NAND U2744 ( .A(y[1805]), .B(x[224]), .Z(n1428) );
  XNOR U2745 ( .A(n1429), .B(n1428), .Z(n1496) );
  AND U2746 ( .A(y[1793]), .B(x[236]), .Z(n1488) );
  XOR U2747 ( .A(o[13]), .B(n1488), .Z(n1495) );
  XOR U2748 ( .A(n1496), .B(n1495), .Z(n1502) );
  AND U2749 ( .A(y[1802]), .B(x[227]), .Z(n1431) );
  NAND U2750 ( .A(x[229]), .B(y[1800]), .Z(n1430) );
  XNOR U2751 ( .A(n1431), .B(n1430), .Z(n1491) );
  AND U2752 ( .A(x[228]), .B(y[1801]), .Z(n1492) );
  XOR U2753 ( .A(n1491), .B(n1492), .Z(n1501) );
  XOR U2754 ( .A(n1502), .B(n1501), .Z(n1504) );
  XNOR U2755 ( .A(n1503), .B(n1504), .Z(n1453) );
  XOR U2756 ( .A(n1454), .B(n1455), .Z(n1509) );
  XNOR U2757 ( .A(n1510), .B(n1509), .Z(n1523) );
  NAND U2758 ( .A(n1433), .B(n1432), .Z(n1437) );
  NAND U2759 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U2760 ( .A(n1437), .B(n1436), .Z(n1522) );
  XOR U2761 ( .A(n1523), .B(n1522), .Z(n1524) );
  XOR U2762 ( .A(n1525), .B(n1524), .Z(n1521) );
  NAND U2763 ( .A(n1439), .B(n1438), .Z(n1443) );
  NAND U2764 ( .A(n1441), .B(n1440), .Z(n1442) );
  NAND U2765 ( .A(n1443), .B(n1442), .Z(n1519) );
  NANDN U2766 ( .A(n1444), .B(n1445), .Z(n1450) );
  NOR U2767 ( .A(n1446), .B(n1445), .Z(n1448) );
  OR U2768 ( .A(n1448), .B(n1447), .Z(n1449) );
  AND U2769 ( .A(n1450), .B(n1449), .Z(n1520) );
  XOR U2770 ( .A(n1519), .B(n1520), .Z(n1451) );
  XNOR U2771 ( .A(n1521), .B(n1451), .Z(N46) );
  NANDN U2772 ( .A(n1453), .B(n1452), .Z(n1457) );
  NAND U2773 ( .A(n1455), .B(n1454), .Z(n1456) );
  NAND U2774 ( .A(n1457), .B(n1456), .Z(n1531) );
  NAND U2775 ( .A(n1459), .B(n1458), .Z(n1463) );
  NAND U2776 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U2777 ( .A(n1463), .B(n1462), .Z(n1538) );
  AND U2778 ( .A(x[235]), .B(y[1797]), .Z(n1659) );
  NAND U2779 ( .A(n1659), .B(n1464), .Z(n1467) );
  NAND U2780 ( .A(n1465), .B(n2333), .Z(n1466) );
  NAND U2781 ( .A(n1467), .B(n1466), .Z(n1594) );
  AND U2782 ( .A(y[1804]), .B(x[231]), .Z(n2112) );
  NAND U2783 ( .A(n2112), .B(n1468), .Z(n1472) );
  NAND U2784 ( .A(n1470), .B(n1469), .Z(n1471) );
  NAND U2785 ( .A(n1472), .B(n1471), .Z(n1593) );
  XOR U2786 ( .A(n1594), .B(n1593), .Z(n1596) );
  AND U2787 ( .A(x[228]), .B(y[1802]), .Z(n1967) );
  AND U2788 ( .A(x[232]), .B(y[1798]), .Z(n1474) );
  NAND U2789 ( .A(x[227]), .B(y[1803]), .Z(n1473) );
  XNOR U2790 ( .A(n1474), .B(n1473), .Z(n1579) );
  XOR U2791 ( .A(n1860), .B(n1579), .Z(n1588) );
  XOR U2792 ( .A(n1967), .B(n1588), .Z(n1590) );
  AND U2793 ( .A(x[233]), .B(y[1797]), .Z(n2157) );
  AND U2794 ( .A(y[1804]), .B(x[226]), .Z(n1475) );
  AND U2795 ( .A(y[1796]), .B(x[234]), .Z(n2187) );
  XOR U2796 ( .A(n1475), .B(n2187), .Z(n1564) );
  XOR U2797 ( .A(n2157), .B(n1564), .Z(n1589) );
  XOR U2798 ( .A(n1590), .B(n1589), .Z(n1595) );
  XNOR U2799 ( .A(n1596), .B(n1595), .Z(n1536) );
  NAND U2800 ( .A(n1477), .B(n1476), .Z(n1481) );
  NAND U2801 ( .A(n1479), .B(n1478), .Z(n1480) );
  AND U2802 ( .A(n1481), .B(n1480), .Z(n1535) );
  XOR U2803 ( .A(n1536), .B(n1535), .Z(n1537) );
  XOR U2804 ( .A(n1538), .B(n1537), .Z(n1530) );
  AND U2805 ( .A(y[1803]), .B(x[233]), .Z(n1482) );
  NAND U2806 ( .A(n1482), .B(n1563), .Z(n1485) );
  NAND U2807 ( .A(n1483), .B(n2480), .Z(n1484) );
  NAND U2808 ( .A(n1485), .B(n1484), .Z(n1550) );
  AND U2809 ( .A(x[238]), .B(y[1792]), .Z(n1487) );
  NAND U2810 ( .A(y[1806]), .B(x[224]), .Z(n1486) );
  XNOR U2811 ( .A(n1487), .B(n1486), .Z(n1574) );
  AND U2812 ( .A(o[13]), .B(n1488), .Z(n1573) );
  XOR U2813 ( .A(n1574), .B(n1573), .Z(n1548) );
  NAND U2814 ( .A(y[1794]), .B(x[236]), .Z(n1489) );
  XNOR U2815 ( .A(n1490), .B(n1489), .Z(n1555) );
  AND U2816 ( .A(y[1793]), .B(x[237]), .Z(n1562) );
  XOR U2817 ( .A(o[14]), .B(n1562), .Z(n1554) );
  XOR U2818 ( .A(n1555), .B(n1554), .Z(n1547) );
  XOR U2819 ( .A(n1548), .B(n1547), .Z(n1549) );
  XOR U2820 ( .A(n1550), .B(n1549), .Z(n1600) );
  AND U2821 ( .A(y[1802]), .B(x[229]), .Z(n1646) );
  NANDN U2822 ( .A(n2321), .B(n1646), .Z(n1494) );
  NAND U2823 ( .A(n1492), .B(n1491), .Z(n1493) );
  AND U2824 ( .A(n1494), .B(n1493), .Z(n1544) );
  AND U2825 ( .A(y[1805]), .B(x[237]), .Z(n3051) );
  NAND U2826 ( .A(n3051), .B(n1633), .Z(n1498) );
  NAND U2827 ( .A(n1496), .B(n1495), .Z(n1497) );
  NAND U2828 ( .A(n1498), .B(n1497), .Z(n1542) );
  AND U2829 ( .A(y[1795]), .B(x[235]), .Z(n1500) );
  NAND U2830 ( .A(x[230]), .B(y[1800]), .Z(n1499) );
  XNOR U2831 ( .A(n1500), .B(n1499), .Z(n1569) );
  AND U2832 ( .A(x[225]), .B(y[1805]), .Z(n1570) );
  XOR U2833 ( .A(n1569), .B(n1570), .Z(n1541) );
  XOR U2834 ( .A(n1542), .B(n1541), .Z(n1543) );
  XOR U2835 ( .A(n1544), .B(n1543), .Z(n1599) );
  NAND U2836 ( .A(n1502), .B(n1501), .Z(n1506) );
  NAND U2837 ( .A(n1504), .B(n1503), .Z(n1505) );
  AND U2838 ( .A(n1506), .B(n1505), .Z(n1601) );
  XNOR U2839 ( .A(n1602), .B(n1601), .Z(n1529) );
  XOR U2840 ( .A(n1531), .B(n1532), .Z(n1611) );
  NAND U2841 ( .A(n1508), .B(n1507), .Z(n1512) );
  NAND U2842 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U2843 ( .A(n1512), .B(n1511), .Z(n1609) );
  NAND U2844 ( .A(n1514), .B(n1513), .Z(n1518) );
  NAND U2845 ( .A(n1516), .B(n1515), .Z(n1517) );
  NAND U2846 ( .A(n1518), .B(n1517), .Z(n1608) );
  XOR U2847 ( .A(n1609), .B(n1608), .Z(n1610) );
  XNOR U2848 ( .A(n1611), .B(n1610), .Z(n1607) );
  NAND U2849 ( .A(n1523), .B(n1522), .Z(n1527) );
  NANDN U2850 ( .A(n1525), .B(n1524), .Z(n1526) );
  AND U2851 ( .A(n1527), .B(n1526), .Z(n1606) );
  XOR U2852 ( .A(n1605), .B(n1606), .Z(n1528) );
  XNOR U2853 ( .A(n1607), .B(n1528), .Z(N47) );
  NANDN U2854 ( .A(n1530), .B(n1529), .Z(n1534) );
  NAND U2855 ( .A(n1532), .B(n1531), .Z(n1533) );
  NAND U2856 ( .A(n1534), .B(n1533), .Z(n1617) );
  NAND U2857 ( .A(n1536), .B(n1535), .Z(n1540) );
  NAND U2858 ( .A(n1538), .B(n1537), .Z(n1539) );
  NAND U2859 ( .A(n1540), .B(n1539), .Z(n1689) );
  NAND U2860 ( .A(n1542), .B(n1541), .Z(n1546) );
  NANDN U2861 ( .A(n1544), .B(n1543), .Z(n1545) );
  NAND U2862 ( .A(n1546), .B(n1545), .Z(n1695) );
  NAND U2863 ( .A(n1548), .B(n1547), .Z(n1552) );
  NAND U2864 ( .A(n1550), .B(n1549), .Z(n1551) );
  NAND U2865 ( .A(n1552), .B(n1551), .Z(n1693) );
  AND U2866 ( .A(x[236]), .B(y[1799]), .Z(n2103) );
  NAND U2867 ( .A(n2103), .B(n1553), .Z(n1557) );
  NAND U2868 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U2869 ( .A(n1557), .B(n1556), .Z(n1669) );
  AND U2870 ( .A(y[1796]), .B(x[235]), .Z(n1559) );
  NAND U2871 ( .A(y[1794]), .B(x[237]), .Z(n1558) );
  XNOR U2872 ( .A(n1559), .B(n1558), .Z(n1673) );
  AND U2873 ( .A(x[236]), .B(y[1795]), .Z(n1672) );
  XNOR U2874 ( .A(n1673), .B(n1672), .Z(n1667) );
  AND U2875 ( .A(x[239]), .B(y[1792]), .Z(n1561) );
  NAND U2876 ( .A(y[1807]), .B(x[224]), .Z(n1560) );
  XNOR U2877 ( .A(n1561), .B(n1560), .Z(n1635) );
  AND U2878 ( .A(o[14]), .B(n1562), .Z(n1634) );
  XNOR U2879 ( .A(n1635), .B(n1634), .Z(n1666) );
  XOR U2880 ( .A(n1667), .B(n1666), .Z(n1668) );
  XNOR U2881 ( .A(n1669), .B(n1668), .Z(n1701) );
  NAND U2882 ( .A(x[234]), .B(y[1804]), .Z(n2482) );
  NANDN U2883 ( .A(n2482), .B(n1563), .Z(n1566) );
  NAND U2884 ( .A(n2157), .B(n1564), .Z(n1565) );
  NAND U2885 ( .A(n1566), .B(n1565), .Z(n1699) );
  AND U2886 ( .A(y[1800]), .B(x[235]), .Z(n1568) );
  NAND U2887 ( .A(n1568), .B(n1567), .Z(n1572) );
  NAND U2888 ( .A(n1570), .B(n1569), .Z(n1571) );
  NAND U2889 ( .A(n1572), .B(n1571), .Z(n1698) );
  XOR U2890 ( .A(n1699), .B(n1698), .Z(n1700) );
  XOR U2891 ( .A(n1701), .B(n1700), .Z(n1692) );
  XOR U2892 ( .A(n1693), .B(n1692), .Z(n1694) );
  XNOR U2893 ( .A(n1695), .B(n1694), .Z(n1686) );
  AND U2894 ( .A(y[1806]), .B(x[238]), .Z(n3311) );
  NAND U2895 ( .A(n3311), .B(n1633), .Z(n1576) );
  NAND U2896 ( .A(n1574), .B(n1573), .Z(n1575) );
  NAND U2897 ( .A(n1576), .B(n1575), .Z(n1661) );
  AND U2898 ( .A(y[1803]), .B(x[232]), .Z(n1577) );
  NANDN U2899 ( .A(n1578), .B(n1577), .Z(n1581) );
  NAND U2900 ( .A(n1579), .B(n1860), .Z(n1580) );
  NAND U2901 ( .A(n1581), .B(n1580), .Z(n1660) );
  XOR U2902 ( .A(n1661), .B(n1660), .Z(n1663) );
  AND U2903 ( .A(y[1797]), .B(x[234]), .Z(n1583) );
  NAND U2904 ( .A(x[228]), .B(y[1803]), .Z(n1582) );
  XNOR U2905 ( .A(n1583), .B(n1582), .Z(n1641) );
  AND U2906 ( .A(y[1800]), .B(x[231]), .Z(n1640) );
  XNOR U2907 ( .A(n1641), .B(n1640), .Z(n1648) );
  NAND U2908 ( .A(y[1801]), .B(x[230]), .Z(n1738) );
  XNOR U2909 ( .A(n1738), .B(n1646), .Z(n1647) );
  XNOR U2910 ( .A(n1648), .B(n1647), .Z(n1682) );
  AND U2911 ( .A(y[1805]), .B(x[226]), .Z(n1585) );
  NAND U2912 ( .A(x[233]), .B(y[1798]), .Z(n1584) );
  XNOR U2913 ( .A(n1585), .B(n1584), .Z(n1651) );
  AND U2914 ( .A(y[1804]), .B(x[227]), .Z(n1652) );
  XOR U2915 ( .A(n1651), .B(n1652), .Z(n1681) );
  AND U2916 ( .A(y[1806]), .B(x[225]), .Z(n1587) );
  NAND U2917 ( .A(y[1799]), .B(x[232]), .Z(n1586) );
  XNOR U2918 ( .A(n1587), .B(n1586), .Z(n1630) );
  AND U2919 ( .A(y[1793]), .B(x[238]), .Z(n1657) );
  XOR U2920 ( .A(o[15]), .B(n1657), .Z(n1629) );
  XOR U2921 ( .A(n1630), .B(n1629), .Z(n1680) );
  XOR U2922 ( .A(n1681), .B(n1680), .Z(n1683) );
  XOR U2923 ( .A(n1682), .B(n1683), .Z(n1662) );
  XNOR U2924 ( .A(n1663), .B(n1662), .Z(n1705) );
  NAND U2925 ( .A(n1967), .B(n1588), .Z(n1592) );
  NAND U2926 ( .A(n1590), .B(n1589), .Z(n1591) );
  AND U2927 ( .A(n1592), .B(n1591), .Z(n1704) );
  XOR U2928 ( .A(n1705), .B(n1704), .Z(n1706) );
  NAND U2929 ( .A(n1594), .B(n1593), .Z(n1598) );
  NAND U2930 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U2931 ( .A(n1598), .B(n1597), .Z(n1707) );
  XOR U2932 ( .A(n1706), .B(n1707), .Z(n1687) );
  XOR U2933 ( .A(n1686), .B(n1687), .Z(n1688) );
  XOR U2934 ( .A(n1689), .B(n1688), .Z(n1616) );
  NANDN U2935 ( .A(n1600), .B(n1599), .Z(n1604) );
  NAND U2936 ( .A(n1602), .B(n1601), .Z(n1603) );
  AND U2937 ( .A(n1604), .B(n1603), .Z(n1615) );
  XOR U2938 ( .A(n1617), .B(n1618), .Z(n1624) );
  NAND U2939 ( .A(n1609), .B(n1608), .Z(n1613) );
  NAND U2940 ( .A(n1611), .B(n1610), .Z(n1612) );
  AND U2941 ( .A(n1613), .B(n1612), .Z(n1623) );
  IV U2942 ( .A(n1623), .Z(n1621) );
  XOR U2943 ( .A(n1622), .B(n1621), .Z(n1614) );
  XNOR U2944 ( .A(n1624), .B(n1614), .Z(N48) );
  NANDN U2945 ( .A(n1616), .B(n1615), .Z(n1620) );
  NAND U2946 ( .A(n1618), .B(n1617), .Z(n1619) );
  AND U2947 ( .A(n1620), .B(n1619), .Z(n1802) );
  NANDN U2948 ( .A(n1621), .B(n1622), .Z(n1627) );
  NOR U2949 ( .A(n1623), .B(n1622), .Z(n1625) );
  OR U2950 ( .A(n1625), .B(n1624), .Z(n1626) );
  AND U2951 ( .A(n1627), .B(n1626), .Z(n1803) );
  AND U2952 ( .A(x[232]), .B(y[1806]), .Z(n1968) );
  NAND U2953 ( .A(n1968), .B(n1628), .Z(n1632) );
  NAND U2954 ( .A(n1630), .B(n1629), .Z(n1631) );
  AND U2955 ( .A(n1632), .B(n1631), .Z(n1768) );
  AND U2956 ( .A(x[239]), .B(y[1807]), .Z(n3761) );
  NAND U2957 ( .A(n3761), .B(n1633), .Z(n1637) );
  NAND U2958 ( .A(n1635), .B(n1634), .Z(n1636) );
  NAND U2959 ( .A(n1637), .B(n1636), .Z(n1767) );
  AND U2960 ( .A(y[1803]), .B(x[234]), .Z(n1639) );
  NAND U2961 ( .A(n1639), .B(n1638), .Z(n1643) );
  NAND U2962 ( .A(n1641), .B(n1640), .Z(n1642) );
  NAND U2963 ( .A(n1643), .B(n1642), .Z(n1725) );
  AND U2964 ( .A(x[224]), .B(y[1808]), .Z(n1747) );
  NAND U2965 ( .A(y[1792]), .B(x[240]), .Z(n1748) );
  NAND U2966 ( .A(y[1793]), .B(x[239]), .Z(n1735) );
  XOR U2967 ( .A(o[16]), .B(n1735), .Z(n1750) );
  NAND U2968 ( .A(x[231]), .B(y[1801]), .Z(n1644) );
  XNOR U2969 ( .A(n1645), .B(n1644), .Z(n1740) );
  AND U2970 ( .A(y[1798]), .B(x[234]), .Z(n1739) );
  XOR U2971 ( .A(n1740), .B(n1739), .Z(n1723) );
  XOR U2972 ( .A(n1724), .B(n1723), .Z(n1726) );
  XOR U2973 ( .A(n1725), .B(n1726), .Z(n1769) );
  XNOR U2974 ( .A(n1770), .B(n1769), .Z(n1720) );
  NANDN U2975 ( .A(n1646), .B(n1738), .Z(n1650) );
  NAND U2976 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U2977 ( .A(n1650), .B(n1649), .Z(n1718) );
  AND U2978 ( .A(x[233]), .B(y[1805]), .Z(n2463) );
  NAND U2979 ( .A(n2463), .B(n2102), .Z(n1654) );
  NAND U2980 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U2981 ( .A(n1654), .B(n1653), .Z(n1758) );
  AND U2982 ( .A(y[1807]), .B(x[225]), .Z(n1656) );
  NAND U2983 ( .A(y[1800]), .B(x[232]), .Z(n1655) );
  XNOR U2984 ( .A(n1656), .B(n1655), .Z(n1744) );
  AND U2985 ( .A(o[15]), .B(n1657), .Z(n1743) );
  XOR U2986 ( .A(n1744), .B(n1743), .Z(n1755) );
  NAND U2987 ( .A(y[1794]), .B(x[238]), .Z(n1658) );
  XNOR U2988 ( .A(n1659), .B(n1658), .Z(n1779) );
  NAND U2989 ( .A(x[228]), .B(y[1804]), .Z(n1780) );
  XNOR U2990 ( .A(n1779), .B(n1780), .Z(n1756) );
  XOR U2991 ( .A(n1755), .B(n1756), .Z(n1757) );
  XOR U2992 ( .A(n1758), .B(n1757), .Z(n1717) );
  XOR U2993 ( .A(n1718), .B(n1717), .Z(n1719) );
  XOR U2994 ( .A(n1720), .B(n1719), .Z(n1761) );
  NAND U2995 ( .A(n1661), .B(n1660), .Z(n1665) );
  NAND U2996 ( .A(n1663), .B(n1662), .Z(n1664) );
  AND U2997 ( .A(n1665), .B(n1664), .Z(n1762) );
  XOR U2998 ( .A(n1761), .B(n1762), .Z(n1764) );
  NAND U2999 ( .A(n1667), .B(n1666), .Z(n1671) );
  NAND U3000 ( .A(n1669), .B(n1668), .Z(n1670) );
  NAND U3001 ( .A(n1671), .B(n1670), .Z(n1793) );
  AND U3002 ( .A(x[237]), .B(y[1796]), .Z(n1789) );
  NAND U3003 ( .A(n2294), .B(n1789), .Z(n1675) );
  NAND U3004 ( .A(n1673), .B(n1672), .Z(n1674) );
  NAND U3005 ( .A(n1675), .B(n1674), .Z(n1776) );
  AND U3006 ( .A(x[226]), .B(y[1806]), .Z(n1677) );
  NAND U3007 ( .A(y[1799]), .B(x[233]), .Z(n1676) );
  XNOR U3008 ( .A(n1677), .B(n1676), .Z(n1783) );
  NAND U3009 ( .A(x[227]), .B(y[1805]), .Z(n1784) );
  XNOR U3010 ( .A(n1783), .B(n1784), .Z(n1774) );
  AND U3011 ( .A(x[236]), .B(y[1796]), .Z(n2452) );
  AND U3012 ( .A(y[1795]), .B(x[237]), .Z(n1679) );
  NAND U3013 ( .A(x[229]), .B(y[1803]), .Z(n1678) );
  XNOR U3014 ( .A(n1679), .B(n1678), .Z(n1730) );
  XOR U3015 ( .A(n2452), .B(n1730), .Z(n1773) );
  XOR U3016 ( .A(n1774), .B(n1773), .Z(n1775) );
  XNOR U3017 ( .A(n1776), .B(n1775), .Z(n1790) );
  NAND U3018 ( .A(n1681), .B(n1680), .Z(n1685) );
  NAND U3019 ( .A(n1683), .B(n1682), .Z(n1684) );
  AND U3020 ( .A(n1685), .B(n1684), .Z(n1791) );
  XOR U3021 ( .A(n1790), .B(n1791), .Z(n1792) );
  XOR U3022 ( .A(n1793), .B(n1792), .Z(n1763) );
  XNOR U3023 ( .A(n1764), .B(n1763), .Z(n1797) );
  NAND U3024 ( .A(n1687), .B(n1686), .Z(n1691) );
  NAND U3025 ( .A(n1689), .B(n1688), .Z(n1690) );
  AND U3026 ( .A(n1691), .B(n1690), .Z(n1796) );
  XOR U3027 ( .A(n1797), .B(n1796), .Z(n1799) );
  NAND U3028 ( .A(n1693), .B(n1692), .Z(n1697) );
  NAND U3029 ( .A(n1695), .B(n1694), .Z(n1696) );
  NAND U3030 ( .A(n1697), .B(n1696), .Z(n1714) );
  NAND U3031 ( .A(n1699), .B(n1698), .Z(n1703) );
  NAND U3032 ( .A(n1701), .B(n1700), .Z(n1702) );
  NAND U3033 ( .A(n1703), .B(n1702), .Z(n1712) );
  NAND U3034 ( .A(n1705), .B(n1704), .Z(n1709) );
  NAND U3035 ( .A(n1707), .B(n1706), .Z(n1708) );
  AND U3036 ( .A(n1709), .B(n1708), .Z(n1711) );
  XOR U3037 ( .A(n1712), .B(n1711), .Z(n1713) );
  XOR U3038 ( .A(n1714), .B(n1713), .Z(n1798) );
  XOR U3039 ( .A(n1799), .B(n1798), .Z(n1804) );
  XNOR U3040 ( .A(n1803), .B(n1804), .Z(n1710) );
  XOR U3041 ( .A(n1802), .B(n1710), .Z(N49) );
  NAND U3042 ( .A(n1712), .B(n1711), .Z(n1716) );
  NAND U3043 ( .A(n1714), .B(n1713), .Z(n1715) );
  AND U3044 ( .A(n1716), .B(n1715), .Z(n1906) );
  NAND U3045 ( .A(n1718), .B(n1717), .Z(n1722) );
  NAND U3046 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U3047 ( .A(n1722), .B(n1721), .Z(n1815) );
  NAND U3048 ( .A(n1724), .B(n1723), .Z(n1728) );
  NAND U3049 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U3050 ( .A(n1728), .B(n1727), .Z(n1897) );
  AND U3051 ( .A(y[1803]), .B(x[237]), .Z(n2682) );
  NAND U3052 ( .A(n2682), .B(n1729), .Z(n1732) );
  NAND U3053 ( .A(n1730), .B(n2452), .Z(n1731) );
  AND U3054 ( .A(n1732), .B(n1731), .Z(n1845) );
  AND U3055 ( .A(y[1808]), .B(x[225]), .Z(n1734) );
  NAND U3056 ( .A(y[1800]), .B(x[233]), .Z(n1733) );
  XNOR U3057 ( .A(n1734), .B(n1733), .Z(n1865) );
  NANDN U3058 ( .A(n1735), .B(o[16]), .Z(n1866) );
  XNOR U3059 ( .A(n1865), .B(n1866), .Z(n1843) );
  AND U3060 ( .A(y[1794]), .B(x[239]), .Z(n1737) );
  NAND U3061 ( .A(y[1797]), .B(x[236]), .Z(n1736) );
  XNOR U3062 ( .A(n1737), .B(n1736), .Z(n1819) );
  AND U3063 ( .A(x[238]), .B(y[1795]), .Z(n1818) );
  XOR U3064 ( .A(n1819), .B(n1818), .Z(n1842) );
  XOR U3065 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U3066 ( .A(x[231]), .B(y[1802]), .Z(n1877) );
  NANDN U3067 ( .A(n1738), .B(n1877), .Z(n1742) );
  NAND U3068 ( .A(n1740), .B(n1739), .Z(n1741) );
  AND U3069 ( .A(n1742), .B(n1741), .Z(n1855) );
  AND U3070 ( .A(x[232]), .B(y[1807]), .Z(n2585) );
  AND U3071 ( .A(x[225]), .B(y[1800]), .Z(n1946) );
  NAND U3072 ( .A(n2585), .B(n1946), .Z(n1746) );
  NAND U3073 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U3074 ( .A(n1746), .B(n1745), .Z(n1854) );
  NANDN U3075 ( .A(n1748), .B(n1747), .Z(n1752) );
  NANDN U3076 ( .A(n1750), .B(n1749), .Z(n1751) );
  AND U3077 ( .A(n1752), .B(n1751), .Z(n1851) );
  AND U3078 ( .A(x[224]), .B(y[1809]), .Z(n1833) );
  AND U3079 ( .A(x[241]), .B(y[1792]), .Z(n1832) );
  XOR U3080 ( .A(n1833), .B(n1832), .Z(n1835) );
  AND U3081 ( .A(y[1793]), .B(x[240]), .Z(n1829) );
  XOR U3082 ( .A(n1829), .B(o[17]), .Z(n1834) );
  XOR U3083 ( .A(n1835), .B(n1834), .Z(n1848) );
  AND U3084 ( .A(y[1807]), .B(x[226]), .Z(n1754) );
  NAND U3085 ( .A(y[1799]), .B(x[234]), .Z(n1753) );
  XNOR U3086 ( .A(n1754), .B(n1753), .Z(n1870) );
  NAND U3087 ( .A(y[1806]), .B(x[227]), .Z(n1871) );
  XOR U3088 ( .A(n1870), .B(n1871), .Z(n1849) );
  XOR U3089 ( .A(n1857), .B(n1856), .Z(n1894) );
  XOR U3090 ( .A(n1895), .B(n1894), .Z(n1896) );
  NAND U3091 ( .A(n1756), .B(n1755), .Z(n1760) );
  NANDN U3092 ( .A(n1758), .B(n1757), .Z(n1759) );
  AND U3093 ( .A(n1760), .B(n1759), .Z(n1813) );
  XOR U3094 ( .A(n1812), .B(n1813), .Z(n1814) );
  XNOR U3095 ( .A(n1815), .B(n1814), .Z(n1904) );
  NAND U3096 ( .A(n1762), .B(n1761), .Z(n1766) );
  NAND U3097 ( .A(n1764), .B(n1763), .Z(n1765) );
  AND U3098 ( .A(n1766), .B(n1765), .Z(n1809) );
  NANDN U3099 ( .A(n1768), .B(n1767), .Z(n1772) );
  NAND U3100 ( .A(n1770), .B(n1769), .Z(n1771) );
  NAND U3101 ( .A(n1772), .B(n1771), .Z(n1891) );
  NAND U3102 ( .A(n1774), .B(n1773), .Z(n1778) );
  NAND U3103 ( .A(n1776), .B(n1775), .Z(n1777) );
  NAND U3104 ( .A(n1778), .B(n1777), .Z(n1889) );
  NAND U3105 ( .A(x[238]), .B(y[1797]), .Z(n2077) );
  NANDN U3106 ( .A(n2077), .B(n2294), .Z(n1782) );
  NANDN U3107 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U3108 ( .A(n1782), .B(n1781), .Z(n1883) );
  AND U3109 ( .A(x[233]), .B(y[1806]), .Z(n2663) );
  NAND U3110 ( .A(n1869), .B(n2663), .Z(n1786) );
  NANDN U3111 ( .A(n1784), .B(n1783), .Z(n1785) );
  NAND U3112 ( .A(n1786), .B(n1785), .Z(n1882) );
  XNOR U3113 ( .A(n1883), .B(n1882), .Z(n1884) );
  AND U3114 ( .A(y[1804]), .B(x[229]), .Z(n1928) );
  NAND U3115 ( .A(y[1801]), .B(x[232]), .Z(n1787) );
  XNOR U3116 ( .A(n1928), .B(n1787), .Z(n1862) );
  XOR U3117 ( .A(n1862), .B(n1861), .Z(n1876) );
  XOR U3118 ( .A(n1876), .B(n1877), .Z(n1878) );
  NAND U3119 ( .A(y[1805]), .B(x[228]), .Z(n1788) );
  XNOR U3120 ( .A(n1789), .B(n1788), .Z(n1823) );
  NAND U3121 ( .A(y[1798]), .B(x[235]), .Z(n1824) );
  XOR U3122 ( .A(n1823), .B(n1824), .Z(n1879) );
  XOR U3123 ( .A(n1878), .B(n1879), .Z(n1885) );
  XNOR U3124 ( .A(n1884), .B(n1885), .Z(n1888) );
  XOR U3125 ( .A(n1889), .B(n1888), .Z(n1890) );
  XNOR U3126 ( .A(n1891), .B(n1890), .Z(n1807) );
  NAND U3127 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U3128 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U3129 ( .A(n1795), .B(n1794), .Z(n1806) );
  XOR U3130 ( .A(n1807), .B(n1806), .Z(n1808) );
  XOR U3131 ( .A(n1809), .B(n1808), .Z(n1903) );
  XOR U3132 ( .A(n1904), .B(n1903), .Z(n1905) );
  XOR U3133 ( .A(n1906), .B(n1905), .Z(n1902) );
  NAND U3134 ( .A(n1797), .B(n1796), .Z(n1801) );
  NAND U3135 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U3136 ( .A(n1801), .B(n1800), .Z(n1901) );
  XOR U3137 ( .A(n1901), .B(n1900), .Z(n1805) );
  XNOR U3138 ( .A(n1902), .B(n1805), .Z(N50) );
  NAND U3139 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U3140 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U3141 ( .A(n1811), .B(n1810), .Z(n2015) );
  NAND U3142 ( .A(n1813), .B(n1812), .Z(n1817) );
  NAND U3143 ( .A(n1815), .B(n1814), .Z(n1816) );
  AND U3144 ( .A(n1817), .B(n1816), .Z(n2013) );
  AND U3145 ( .A(x[239]), .B(y[1797]), .Z(n2110) );
  AND U3146 ( .A(x[236]), .B(y[1794]), .Z(n2150) );
  NAND U3147 ( .A(n2110), .B(n2150), .Z(n1821) );
  NAND U3148 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U3149 ( .A(n1821), .B(n1820), .Z(n1994) );
  NAND U3150 ( .A(n3051), .B(n1822), .Z(n1826) );
  NANDN U3151 ( .A(n1824), .B(n1823), .Z(n1825) );
  AND U3152 ( .A(n1826), .B(n1825), .Z(n1985) );
  AND U3153 ( .A(x[225]), .B(y[1809]), .Z(n1828) );
  NAND U3154 ( .A(y[1800]), .B(x[234]), .Z(n1827) );
  XNOR U3155 ( .A(n1828), .B(n1827), .Z(n1948) );
  AND U3156 ( .A(n1829), .B(o[17]), .Z(n1947) );
  XOR U3157 ( .A(n1948), .B(n1947), .Z(n1982) );
  AND U3158 ( .A(y[1795]), .B(x[239]), .Z(n1831) );
  NAND U3159 ( .A(y[1801]), .B(x[233]), .Z(n1830) );
  XNOR U3160 ( .A(n1831), .B(n1830), .Z(n1939) );
  AND U3161 ( .A(x[238]), .B(y[1796]), .Z(n1938) );
  XNOR U3162 ( .A(n1939), .B(n1938), .Z(n1983) );
  XNOR U3163 ( .A(n1982), .B(n1983), .Z(n1984) );
  XNOR U3164 ( .A(n1985), .B(n1984), .Z(n1995) );
  XOR U3165 ( .A(n1994), .B(n1995), .Z(n1997) );
  NAND U3166 ( .A(n1833), .B(n1832), .Z(n1837) );
  NAND U3167 ( .A(n1835), .B(n1834), .Z(n1836) );
  NAND U3168 ( .A(n1837), .B(n1836), .Z(n2006) );
  AND U3169 ( .A(y[1794]), .B(x[240]), .Z(n1839) );
  NAND U3170 ( .A(x[235]), .B(y[1799]), .Z(n1838) );
  XNOR U3171 ( .A(n1839), .B(n1838), .Z(n1934) );
  NAND U3172 ( .A(x[226]), .B(y[1808]), .Z(n1935) );
  XNOR U3173 ( .A(n1934), .B(n1935), .Z(n2007) );
  XOR U3174 ( .A(n2006), .B(n2007), .Z(n2009) );
  AND U3175 ( .A(x[229]), .B(y[1805]), .Z(n2059) );
  NAND U3176 ( .A(x[230]), .B(y[1804]), .Z(n1840) );
  XNOR U3177 ( .A(n2059), .B(n1840), .Z(n1930) );
  NAND U3178 ( .A(y[1806]), .B(x[228]), .Z(n1841) );
  XNOR U3179 ( .A(n2668), .B(n1841), .Z(n1969) );
  NAND U3180 ( .A(y[1803]), .B(x[231]), .Z(n1970) );
  XNOR U3181 ( .A(n1969), .B(n1970), .Z(n1929) );
  XOR U3182 ( .A(n1930), .B(n1929), .Z(n2008) );
  XOR U3183 ( .A(n2009), .B(n2008), .Z(n1996) );
  XOR U3184 ( .A(n1997), .B(n1996), .Z(n1917) );
  NAND U3185 ( .A(n1843), .B(n1842), .Z(n1847) );
  NANDN U3186 ( .A(n1845), .B(n1844), .Z(n1846) );
  AND U3187 ( .A(n1847), .B(n1846), .Z(n1989) );
  NANDN U3188 ( .A(n1849), .B(n1848), .Z(n1853) );
  NANDN U3189 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U3190 ( .A(n1853), .B(n1852), .Z(n1988) );
  XOR U3191 ( .A(n1989), .B(n1988), .Z(n1991) );
  NANDN U3192 ( .A(n1855), .B(n1854), .Z(n1859) );
  NAND U3193 ( .A(n1857), .B(n1856), .Z(n1858) );
  AND U3194 ( .A(n1859), .B(n1858), .Z(n1990) );
  XOR U3195 ( .A(n1991), .B(n1990), .Z(n1916) );
  AND U3196 ( .A(x[232]), .B(y[1804]), .Z(n2193) );
  NAND U3197 ( .A(n2193), .B(n1860), .Z(n1864) );
  NAND U3198 ( .A(n1862), .B(n1861), .Z(n1863) );
  NAND U3199 ( .A(n1864), .B(n1863), .Z(n2001) );
  AND U3200 ( .A(x[233]), .B(y[1808]), .Z(n2823) );
  NAND U3201 ( .A(n2823), .B(n1946), .Z(n1868) );
  NANDN U3202 ( .A(n1866), .B(n1865), .Z(n1867) );
  NAND U3203 ( .A(n1868), .B(n1867), .Z(n2000) );
  XOR U3204 ( .A(n2001), .B(n2000), .Z(n2003) );
  AND U3205 ( .A(x[234]), .B(y[1807]), .Z(n2691) );
  IV U3206 ( .A(n2691), .Z(n2822) );
  NANDN U3207 ( .A(n2822), .B(n1869), .Z(n1873) );
  NANDN U3208 ( .A(n1871), .B(n1870), .Z(n1872) );
  AND U3209 ( .A(n1873), .B(n1872), .Z(n1979) );
  AND U3210 ( .A(x[224]), .B(y[1810]), .Z(n1952) );
  AND U3211 ( .A(y[1792]), .B(x[242]), .Z(n1951) );
  XOR U3212 ( .A(n1952), .B(n1951), .Z(n1954) );
  AND U3213 ( .A(x[241]), .B(y[1793]), .Z(n1973) );
  XOR U3214 ( .A(n1973), .B(o[18]), .Z(n1953) );
  XOR U3215 ( .A(n1954), .B(n1953), .Z(n1976) );
  AND U3216 ( .A(y[1797]), .B(x[237]), .Z(n1875) );
  NAND U3217 ( .A(y[1807]), .B(x[227]), .Z(n1874) );
  XNOR U3218 ( .A(n1875), .B(n1874), .Z(n1960) );
  AND U3219 ( .A(y[1798]), .B(x[236]), .Z(n1959) );
  XNOR U3220 ( .A(n1960), .B(n1959), .Z(n1977) );
  XNOR U3221 ( .A(n1976), .B(n1977), .Z(n1978) );
  XNOR U3222 ( .A(n1979), .B(n1978), .Z(n2002) );
  XOR U3223 ( .A(n2003), .B(n2002), .Z(n1923) );
  NAND U3224 ( .A(n1877), .B(n1876), .Z(n1881) );
  NANDN U3225 ( .A(n1879), .B(n1878), .Z(n1880) );
  AND U3226 ( .A(n1881), .B(n1880), .Z(n1922) );
  XNOR U3227 ( .A(n1923), .B(n1922), .Z(n1924) );
  NANDN U3228 ( .A(n1883), .B(n1882), .Z(n1887) );
  NANDN U3229 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U3230 ( .A(n1887), .B(n1886), .Z(n1925) );
  XNOR U3231 ( .A(n1924), .B(n1925), .Z(n1918) );
  XOR U3232 ( .A(n1919), .B(n1918), .Z(n1913) );
  NAND U3233 ( .A(n1889), .B(n1888), .Z(n1893) );
  NAND U3234 ( .A(n1891), .B(n1890), .Z(n1892) );
  AND U3235 ( .A(n1893), .B(n1892), .Z(n1911) );
  NAND U3236 ( .A(n1895), .B(n1894), .Z(n1899) );
  NANDN U3237 ( .A(n1897), .B(n1896), .Z(n1898) );
  NAND U3238 ( .A(n1899), .B(n1898), .Z(n1910) );
  XOR U3239 ( .A(n2013), .B(n2012), .Z(n2014) );
  XOR U3240 ( .A(n2015), .B(n2014), .Z(n2021) );
  NAND U3241 ( .A(n1904), .B(n1903), .Z(n1908) );
  NANDN U3242 ( .A(n1906), .B(n1905), .Z(n1907) );
  AND U3243 ( .A(n1908), .B(n1907), .Z(n2020) );
  IV U3244 ( .A(n2020), .Z(n2018) );
  XOR U3245 ( .A(n2019), .B(n2018), .Z(n1909) );
  XNOR U3246 ( .A(n2021), .B(n1909), .Z(N51) );
  NANDN U3247 ( .A(n1911), .B(n1910), .Z(n1915) );
  NANDN U3248 ( .A(n1913), .B(n1912), .Z(n1914) );
  AND U3249 ( .A(n1915), .B(n1914), .Z(n2029) );
  NANDN U3250 ( .A(n1917), .B(n1916), .Z(n1921) );
  NAND U3251 ( .A(n1919), .B(n1918), .Z(n1920) );
  AND U3252 ( .A(n1921), .B(n1920), .Z(n2027) );
  NANDN U3253 ( .A(n1923), .B(n1922), .Z(n1927) );
  NANDN U3254 ( .A(n1925), .B(n1924), .Z(n1926) );
  AND U3255 ( .A(n1927), .B(n1926), .Z(n2038) );
  AND U3256 ( .A(y[1805]), .B(x[230]), .Z(n1975) );
  NAND U3257 ( .A(n1975), .B(n1928), .Z(n1932) );
  NAND U3258 ( .A(n1930), .B(n1929), .Z(n1931) );
  AND U3259 ( .A(n1932), .B(n1931), .Z(n2043) );
  AND U3260 ( .A(y[1799]), .B(x[240]), .Z(n1933) );
  NAND U3261 ( .A(n1933), .B(n2294), .Z(n1937) );
  NANDN U3262 ( .A(n1935), .B(n1934), .Z(n1936) );
  AND U3263 ( .A(n1937), .B(n1936), .Z(n2042) );
  AND U3264 ( .A(x[239]), .B(y[1801]), .Z(n2696) );
  NAND U3265 ( .A(n2696), .B(n2097), .Z(n1941) );
  NAND U3266 ( .A(n1939), .B(n1938), .Z(n1940) );
  NAND U3267 ( .A(n1941), .B(n1940), .Z(n2127) );
  AND U3268 ( .A(x[225]), .B(y[1810]), .Z(n1943) );
  NAND U3269 ( .A(x[232]), .B(y[1803]), .Z(n1942) );
  XNOR U3270 ( .A(n1943), .B(n1942), .Z(n2076) );
  AND U3271 ( .A(x[226]), .B(y[1809]), .Z(n1945) );
  NAND U3272 ( .A(x[237]), .B(y[1798]), .Z(n1944) );
  XNOR U3273 ( .A(n1945), .B(n1944), .Z(n2104) );
  XOR U3274 ( .A(n2104), .B(n2103), .Z(n2125) );
  XOR U3275 ( .A(n2126), .B(n2125), .Z(n2128) );
  XOR U3276 ( .A(n2127), .B(n2128), .Z(n2041) );
  XOR U3277 ( .A(n2042), .B(n2041), .Z(n2044) );
  XOR U3278 ( .A(n2043), .B(n2044), .Z(n2036) );
  NAND U3279 ( .A(x[234]), .B(y[1809]), .Z(n3141) );
  NANDN U3280 ( .A(n3141), .B(n1946), .Z(n1950) );
  NAND U3281 ( .A(n1948), .B(n1947), .Z(n1949) );
  NAND U3282 ( .A(n1950), .B(n1949), .Z(n2087) );
  NAND U3283 ( .A(n1952), .B(n1951), .Z(n1956) );
  NAND U3284 ( .A(n1954), .B(n1953), .Z(n1955) );
  NAND U3285 ( .A(n1956), .B(n1955), .Z(n2085) );
  AND U3286 ( .A(y[1795]), .B(x[240]), .Z(n2747) );
  NAND U3287 ( .A(y[1802]), .B(x[233]), .Z(n1957) );
  XNOR U3288 ( .A(n2747), .B(n1957), .Z(n2098) );
  NAND U3289 ( .A(x[239]), .B(y[1796]), .Z(n2099) );
  XNOR U3290 ( .A(n2098), .B(n2099), .Z(n2086) );
  XOR U3291 ( .A(n2085), .B(n2086), .Z(n2088) );
  XNOR U3292 ( .A(n2087), .B(n2088), .Z(n2049) );
  AND U3293 ( .A(x[237]), .B(y[1807]), .Z(n3341) );
  NANDN U3294 ( .A(n1958), .B(n3341), .Z(n1962) );
  NAND U3295 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U3296 ( .A(n1962), .B(n1961), .Z(n2093) );
  AND U3297 ( .A(y[1801]), .B(x[234]), .Z(n1964) );
  NAND U3298 ( .A(y[1794]), .B(x[241]), .Z(n1963) );
  XNOR U3299 ( .A(n1964), .B(n1963), .Z(n2081) );
  NAND U3300 ( .A(y[1793]), .B(x[242]), .Z(n2118) );
  XOR U3301 ( .A(o[19]), .B(n2118), .Z(n2082) );
  XNOR U3302 ( .A(n2081), .B(n2082), .Z(n2092) );
  AND U3303 ( .A(y[1808]), .B(x[227]), .Z(n1966) );
  NAND U3304 ( .A(x[235]), .B(y[1800]), .Z(n1965) );
  XNOR U3305 ( .A(n1966), .B(n1965), .Z(n2113) );
  XOR U3306 ( .A(n2113), .B(n2112), .Z(n2091) );
  XOR U3307 ( .A(n2092), .B(n2091), .Z(n2094) );
  XOR U3308 ( .A(n2093), .B(n2094), .Z(n2048) );
  NAND U3309 ( .A(n1968), .B(n1967), .Z(n1972) );
  NANDN U3310 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U3311 ( .A(n1972), .B(n1971), .Z(n2121) );
  AND U3312 ( .A(x[224]), .B(y[1811]), .Z(n2063) );
  NAND U3313 ( .A(y[1792]), .B(x[243]), .Z(n2064) );
  XNOR U3314 ( .A(n2063), .B(n2064), .Z(n2065) );
  NAND U3315 ( .A(n1973), .B(o[18]), .Z(n2066) );
  XNOR U3316 ( .A(n2065), .B(n2066), .Z(n2120) );
  AND U3317 ( .A(x[228]), .B(y[1807]), .Z(n2207) );
  NAND U3318 ( .A(x[229]), .B(y[1806]), .Z(n1974) );
  XNOR U3319 ( .A(n1975), .B(n1974), .Z(n2060) );
  XOR U3320 ( .A(n2207), .B(n2060), .Z(n2119) );
  XOR U3321 ( .A(n2120), .B(n2119), .Z(n2122) );
  XNOR U3322 ( .A(n2121), .B(n2122), .Z(n2047) );
  XOR U3323 ( .A(n2049), .B(n2050), .Z(n2055) );
  NANDN U3324 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U3325 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U3326 ( .A(n1981), .B(n1980), .Z(n2054) );
  NANDN U3327 ( .A(n1983), .B(n1982), .Z(n1987) );
  NANDN U3328 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U3329 ( .A(n1987), .B(n1986), .Z(n2053) );
  XOR U3330 ( .A(n2054), .B(n2053), .Z(n2056) );
  XOR U3331 ( .A(n2055), .B(n2056), .Z(n2035) );
  XNOR U3332 ( .A(n2036), .B(n2035), .Z(n2037) );
  XOR U3333 ( .A(n2038), .B(n2037), .Z(n2139) );
  NAND U3334 ( .A(n1989), .B(n1988), .Z(n1993) );
  NAND U3335 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U3336 ( .A(n1993), .B(n1992), .Z(n2137) );
  NAND U3337 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U3338 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U3339 ( .A(n1999), .B(n1998), .Z(n2133) );
  NAND U3340 ( .A(n2001), .B(n2000), .Z(n2005) );
  NAND U3341 ( .A(n2003), .B(n2002), .Z(n2004) );
  NAND U3342 ( .A(n2005), .B(n2004), .Z(n2132) );
  NAND U3343 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U3344 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U3345 ( .A(n2011), .B(n2010), .Z(n2131) );
  XNOR U3346 ( .A(n2132), .B(n2131), .Z(n2134) );
  XNOR U3347 ( .A(n2137), .B(n2138), .Z(n2140) );
  XOR U3348 ( .A(n2139), .B(n2140), .Z(n2026) );
  XOR U3349 ( .A(n2027), .B(n2026), .Z(n2028) );
  XOR U3350 ( .A(n2029), .B(n2028), .Z(n2034) );
  NAND U3351 ( .A(n2013), .B(n2012), .Z(n2017) );
  NAND U3352 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U3353 ( .A(n2017), .B(n2016), .Z(n2033) );
  NANDN U3354 ( .A(n2018), .B(n2019), .Z(n2024) );
  NOR U3355 ( .A(n2020), .B(n2019), .Z(n2022) );
  OR U3356 ( .A(n2022), .B(n2021), .Z(n2023) );
  AND U3357 ( .A(n2024), .B(n2023), .Z(n2032) );
  XOR U3358 ( .A(n2033), .B(n2032), .Z(n2025) );
  XNOR U3359 ( .A(n2034), .B(n2025), .Z(N52) );
  NAND U3360 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U3361 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U3362 ( .A(n2031), .B(n2030), .Z(n2251) );
  IV U3363 ( .A(n2251), .Z(n2250) );
  NANDN U3364 ( .A(n2036), .B(n2035), .Z(n2040) );
  NANDN U3365 ( .A(n2038), .B(n2037), .Z(n2039) );
  AND U3366 ( .A(n2040), .B(n2039), .Z(n2240) );
  NANDN U3367 ( .A(n2042), .B(n2041), .Z(n2046) );
  OR U3368 ( .A(n2044), .B(n2043), .Z(n2045) );
  AND U3369 ( .A(n2046), .B(n2045), .Z(n2247) );
  NANDN U3370 ( .A(n2048), .B(n2047), .Z(n2052) );
  NANDN U3371 ( .A(n2050), .B(n2049), .Z(n2051) );
  AND U3372 ( .A(n2052), .B(n2051), .Z(n2245) );
  NANDN U3373 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U3374 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U3375 ( .A(n2058), .B(n2057), .Z(n2244) );
  XNOR U3376 ( .A(n2245), .B(n2244), .Z(n2246) );
  XOR U3377 ( .A(n2247), .B(n2246), .Z(n2239) );
  AND U3378 ( .A(y[1806]), .B(x[230]), .Z(n2164) );
  NAND U3379 ( .A(n2164), .B(n2059), .Z(n2062) );
  NAND U3380 ( .A(n2207), .B(n2060), .Z(n2061) );
  AND U3381 ( .A(n2062), .B(n2061), .Z(n2172) );
  NANDN U3382 ( .A(n2064), .B(n2063), .Z(n2068) );
  NANDN U3383 ( .A(n2066), .B(n2065), .Z(n2067) );
  AND U3384 ( .A(n2068), .B(n2067), .Z(n2170) );
  AND U3385 ( .A(y[1794]), .B(x[242]), .Z(n2070) );
  NAND U3386 ( .A(y[1800]), .B(x[236]), .Z(n2069) );
  XNOR U3387 ( .A(n2070), .B(n2069), .Z(n2151) );
  NAND U3388 ( .A(x[241]), .B(y[1795]), .Z(n2152) );
  XNOR U3389 ( .A(n2151), .B(n2152), .Z(n2169) );
  XNOR U3390 ( .A(n2170), .B(n2169), .Z(n2171) );
  XOR U3391 ( .A(n2172), .B(n2171), .Z(n2176) );
  AND U3392 ( .A(x[237]), .B(y[1799]), .Z(n2072) );
  NAND U3393 ( .A(x[227]), .B(y[1809]), .Z(n2071) );
  XNOR U3394 ( .A(n2072), .B(n2071), .Z(n2194) );
  XOR U3395 ( .A(n2194), .B(n2193), .Z(n2165) );
  AND U3396 ( .A(x[229]), .B(y[1807]), .Z(n2074) );
  NAND U3397 ( .A(y[1808]), .B(x[228]), .Z(n2073) );
  XNOR U3398 ( .A(n2074), .B(n2073), .Z(n2209) );
  AND U3399 ( .A(y[1805]), .B(x[231]), .Z(n2208) );
  XNOR U3400 ( .A(n2209), .B(n2208), .Z(n2163) );
  XOR U3401 ( .A(n2164), .B(n2163), .Z(n2166) );
  XOR U3402 ( .A(n2165), .B(n2166), .Z(n2218) );
  AND U3403 ( .A(y[1810]), .B(x[232]), .Z(n3291) );
  AND U3404 ( .A(y[1803]), .B(x[225]), .Z(n2075) );
  NAND U3405 ( .A(n3291), .B(n2075), .Z(n2079) );
  NANDN U3406 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U3407 ( .A(n2079), .B(n2078), .Z(n2217) );
  NAND U3408 ( .A(x[241]), .B(y[1801]), .Z(n2977) );
  NANDN U3409 ( .A(n2977), .B(n2080), .Z(n2084) );
  NANDN U3410 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U3411 ( .A(n2084), .B(n2083), .Z(n2216) );
  XOR U3412 ( .A(n2217), .B(n2216), .Z(n2219) );
  XNOR U3413 ( .A(n2218), .B(n2219), .Z(n2175) );
  XOR U3414 ( .A(n2176), .B(n2175), .Z(n2178) );
  NAND U3415 ( .A(n2086), .B(n2085), .Z(n2090) );
  NAND U3416 ( .A(n2088), .B(n2087), .Z(n2089) );
  AND U3417 ( .A(n2090), .B(n2089), .Z(n2177) );
  XOR U3418 ( .A(n2178), .B(n2177), .Z(n2233) );
  NAND U3419 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U3420 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U3421 ( .A(n2096), .B(n2095), .Z(n2232) );
  XOR U3422 ( .A(n2233), .B(n2232), .Z(n2235) );
  AND U3423 ( .A(x[240]), .B(y[1802]), .Z(n2971) );
  NAND U3424 ( .A(n2971), .B(n2097), .Z(n2101) );
  NANDN U3425 ( .A(n2099), .B(n2098), .Z(n2100) );
  AND U3426 ( .A(n2101), .B(n2100), .Z(n2182) );
  AND U3427 ( .A(y[1809]), .B(x[237]), .Z(n3454) );
  NAND U3428 ( .A(n3454), .B(n2102), .Z(n2106) );
  NAND U3429 ( .A(n2104), .B(n2103), .Z(n2105) );
  AND U3430 ( .A(n2106), .B(n2105), .Z(n2225) );
  AND U3431 ( .A(y[1796]), .B(x[240]), .Z(n2108) );
  NAND U3432 ( .A(y[1802]), .B(x[234]), .Z(n2107) );
  XNOR U3433 ( .A(n2108), .B(n2107), .Z(n2188) );
  NAND U3434 ( .A(y[1810]), .B(x[226]), .Z(n2189) );
  XNOR U3435 ( .A(n2188), .B(n2189), .Z(n2222) );
  NAND U3436 ( .A(x[233]), .B(y[1803]), .Z(n2109) );
  XNOR U3437 ( .A(n2110), .B(n2109), .Z(n2158) );
  NAND U3438 ( .A(y[1798]), .B(x[238]), .Z(n2159) );
  XOR U3439 ( .A(n2158), .B(n2159), .Z(n2223) );
  XNOR U3440 ( .A(n2222), .B(n2223), .Z(n2224) );
  XNOR U3441 ( .A(n2225), .B(n2224), .Z(n2181) );
  XNOR U3442 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U3443 ( .A(x[235]), .B(y[1808]), .Z(n3143) );
  NANDN U3444 ( .A(n3143), .B(n2111), .Z(n2115) );
  NAND U3445 ( .A(n2113), .B(n2112), .Z(n2114) );
  AND U3446 ( .A(n2115), .B(n2114), .Z(n2231) );
  AND U3447 ( .A(x[235]), .B(y[1801]), .Z(n2117) );
  NAND U3448 ( .A(x[225]), .B(y[1811]), .Z(n2116) );
  XNOR U3449 ( .A(n2117), .B(n2116), .Z(n2156) );
  AND U3450 ( .A(y[1793]), .B(x[243]), .Z(n2162) );
  XOR U3451 ( .A(o[20]), .B(n2162), .Z(n2155) );
  XOR U3452 ( .A(n2156), .B(n2155), .Z(n2229) );
  AND U3453 ( .A(x[224]), .B(y[1812]), .Z(n2212) );
  NAND U3454 ( .A(y[1792]), .B(x[244]), .Z(n2213) );
  XNOR U3455 ( .A(n2212), .B(n2213), .Z(n2215) );
  ANDN U3456 ( .B(o[19]), .A(n2118), .Z(n2214) );
  XOR U3457 ( .A(n2215), .B(n2214), .Z(n2228) );
  XOR U3458 ( .A(n2229), .B(n2228), .Z(n2230) );
  XOR U3459 ( .A(n2231), .B(n2230), .Z(n2184) );
  XOR U3460 ( .A(n2183), .B(n2184), .Z(n2146) );
  NAND U3461 ( .A(n2120), .B(n2119), .Z(n2124) );
  NAND U3462 ( .A(n2122), .B(n2121), .Z(n2123) );
  AND U3463 ( .A(n2124), .B(n2123), .Z(n2145) );
  NAND U3464 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U3465 ( .A(n2128), .B(n2127), .Z(n2129) );
  AND U3466 ( .A(n2130), .B(n2129), .Z(n2144) );
  XOR U3467 ( .A(n2145), .B(n2144), .Z(n2147) );
  XOR U3468 ( .A(n2146), .B(n2147), .Z(n2234) );
  XNOR U3469 ( .A(n2235), .B(n2234), .Z(n2238) );
  XOR U3470 ( .A(n2239), .B(n2238), .Z(n2241) );
  XOR U3471 ( .A(n2240), .B(n2241), .Z(n2259) );
  NAND U3472 ( .A(n2132), .B(n2131), .Z(n2136) );
  NANDN U3473 ( .A(n2134), .B(n2133), .Z(n2135) );
  AND U3474 ( .A(n2136), .B(n2135), .Z(n2258) );
  NANDN U3475 ( .A(n2138), .B(n2137), .Z(n2142) );
  NAND U3476 ( .A(n2140), .B(n2139), .Z(n2141) );
  AND U3477 ( .A(n2142), .B(n2141), .Z(n2257) );
  XOR U3478 ( .A(n2258), .B(n2257), .Z(n2260) );
  XOR U3479 ( .A(n2259), .B(n2260), .Z(n2253) );
  XNOR U3480 ( .A(n2252), .B(n2253), .Z(n2143) );
  XOR U3481 ( .A(n2250), .B(n2143), .Z(N53) );
  NAND U3482 ( .A(n2145), .B(n2144), .Z(n2149) );
  NAND U3483 ( .A(n2147), .B(n2146), .Z(n2148) );
  AND U3484 ( .A(n2149), .B(n2148), .Z(n2272) );
  AND U3485 ( .A(y[1800]), .B(x[242]), .Z(n2980) );
  NAND U3486 ( .A(n2980), .B(n2150), .Z(n2154) );
  NANDN U3487 ( .A(n2152), .B(n2151), .Z(n2153) );
  AND U3488 ( .A(n2154), .B(n2153), .Z(n2350) );
  AND U3489 ( .A(y[1811]), .B(x[235]), .Z(n3781) );
  XNOR U3490 ( .A(n2350), .B(n2349), .Z(n2352) );
  AND U3491 ( .A(y[1803]), .B(x[239]), .Z(n2966) );
  NAND U3492 ( .A(n2966), .B(n2157), .Z(n2161) );
  NANDN U3493 ( .A(n2159), .B(n2158), .Z(n2160) );
  NAND U3494 ( .A(n2161), .B(n2160), .Z(n2307) );
  AND U3495 ( .A(x[224]), .B(y[1813]), .Z(n2327) );
  AND U3496 ( .A(y[1792]), .B(x[245]), .Z(n2328) );
  XOR U3497 ( .A(n2327), .B(n2328), .Z(n2330) );
  AND U3498 ( .A(o[20]), .B(n2162), .Z(n2329) );
  XOR U3499 ( .A(n2330), .B(n2329), .Z(n2306) );
  AND U3500 ( .A(y[1808]), .B(x[229]), .Z(n2312) );
  AND U3501 ( .A(x[240]), .B(y[1797]), .Z(n2311) );
  XOR U3502 ( .A(n2312), .B(n2311), .Z(n2314) );
  AND U3503 ( .A(y[1798]), .B(x[239]), .Z(n2313) );
  XOR U3504 ( .A(n2314), .B(n2313), .Z(n2305) );
  XOR U3505 ( .A(n2306), .B(n2305), .Z(n2308) );
  XOR U3506 ( .A(n2307), .B(n2308), .Z(n2351) );
  XOR U3507 ( .A(n2352), .B(n2351), .Z(n2344) );
  NANDN U3508 ( .A(n2164), .B(n2163), .Z(n2168) );
  OR U3509 ( .A(n2166), .B(n2165), .Z(n2167) );
  NAND U3510 ( .A(n2168), .B(n2167), .Z(n2343) );
  XNOR U3511 ( .A(n2344), .B(n2343), .Z(n2345) );
  NANDN U3512 ( .A(n2170), .B(n2169), .Z(n2174) );
  NANDN U3513 ( .A(n2172), .B(n2171), .Z(n2173) );
  NAND U3514 ( .A(n2174), .B(n2173), .Z(n2346) );
  XOR U3515 ( .A(n2345), .B(n2346), .Z(n2270) );
  NAND U3516 ( .A(n2176), .B(n2175), .Z(n2180) );
  NAND U3517 ( .A(n2178), .B(n2177), .Z(n2179) );
  AND U3518 ( .A(n2180), .B(n2179), .Z(n2271) );
  XOR U3519 ( .A(n2270), .B(n2271), .Z(n2273) );
  XNOR U3520 ( .A(n2272), .B(n2273), .Z(n2266) );
  NANDN U3521 ( .A(n2182), .B(n2181), .Z(n2186) );
  NANDN U3522 ( .A(n2184), .B(n2183), .Z(n2185) );
  AND U3523 ( .A(n2186), .B(n2185), .Z(n2368) );
  NAND U3524 ( .A(n2971), .B(n2187), .Z(n2191) );
  NANDN U3525 ( .A(n2189), .B(n2188), .Z(n2190) );
  AND U3526 ( .A(n2191), .B(n2190), .Z(n2277) );
  NAND U3527 ( .A(n3454), .B(n2192), .Z(n2196) );
  NAND U3528 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U3529 ( .A(n2196), .B(n2195), .Z(n2364) );
  AND U3530 ( .A(y[1794]), .B(x[243]), .Z(n2198) );
  NAND U3531 ( .A(y[1802]), .B(x[235]), .Z(n2197) );
  XNOR U3532 ( .A(n2198), .B(n2197), .Z(n2296) );
  AND U3533 ( .A(y[1793]), .B(x[244]), .Z(n2326) );
  XOR U3534 ( .A(n2326), .B(o[21]), .Z(n2295) );
  XOR U3535 ( .A(n2296), .B(n2295), .Z(n2362) );
  AND U3536 ( .A(y[1795]), .B(x[242]), .Z(n2200) );
  NAND U3537 ( .A(x[234]), .B(y[1803]), .Z(n2199) );
  XNOR U3538 ( .A(n2200), .B(n2199), .Z(n2334) );
  AND U3539 ( .A(y[1812]), .B(x[225]), .Z(n2335) );
  XOR U3540 ( .A(n2334), .B(n2335), .Z(n2361) );
  XOR U3541 ( .A(n2362), .B(n2361), .Z(n2363) );
  XNOR U3542 ( .A(n2364), .B(n2363), .Z(n2276) );
  XNOR U3543 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U3544 ( .A(y[1806]), .B(x[231]), .Z(n2584) );
  AND U3545 ( .A(x[230]), .B(y[1807]), .Z(n2202) );
  NAND U3546 ( .A(x[238]), .B(y[1799]), .Z(n2201) );
  XNOR U3547 ( .A(n2202), .B(n2201), .Z(n2338) );
  XNOR U3548 ( .A(n2584), .B(n2338), .Z(n2285) );
  NAND U3549 ( .A(x[233]), .B(y[1804]), .Z(n2283) );
  NAND U3550 ( .A(x[232]), .B(y[1805]), .Z(n2282) );
  XOR U3551 ( .A(n2283), .B(n2282), .Z(n2284) );
  XNOR U3552 ( .A(n2285), .B(n2284), .Z(n2302) );
  AND U3553 ( .A(y[1801]), .B(x[236]), .Z(n2204) );
  NAND U3554 ( .A(y[1796]), .B(x[241]), .Z(n2203) );
  XNOR U3555 ( .A(n2204), .B(n2203), .Z(n2288) );
  AND U3556 ( .A(y[1811]), .B(x[226]), .Z(n2289) );
  XOR U3557 ( .A(n2288), .B(n2289), .Z(n2300) );
  AND U3558 ( .A(x[237]), .B(y[1800]), .Z(n2206) );
  NAND U3559 ( .A(x[227]), .B(y[1810]), .Z(n2205) );
  XNOR U3560 ( .A(n2206), .B(n2205), .Z(n2323) );
  AND U3561 ( .A(x[228]), .B(y[1809]), .Z(n2322) );
  XOR U3562 ( .A(n2323), .B(n2322), .Z(n2299) );
  XOR U3563 ( .A(n2300), .B(n2299), .Z(n2301) );
  XOR U3564 ( .A(n2302), .B(n2301), .Z(n2357) );
  NAND U3565 ( .A(n2312), .B(n2207), .Z(n2211) );
  NAND U3566 ( .A(n2209), .B(n2208), .Z(n2210) );
  AND U3567 ( .A(n2211), .B(n2210), .Z(n2356) );
  XOR U3568 ( .A(n2356), .B(n2355), .Z(n2358) );
  XOR U3569 ( .A(n2357), .B(n2358), .Z(n2279) );
  XNOR U3570 ( .A(n2278), .B(n2279), .Z(n2366) );
  NANDN U3571 ( .A(n2217), .B(n2216), .Z(n2221) );
  OR U3572 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U3573 ( .A(n2221), .B(n2220), .Z(n2371) );
  NANDN U3574 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U3575 ( .A(n2225), .B(n2224), .Z(n2226) );
  NAND U3576 ( .A(n2227), .B(n2226), .Z(n2370) );
  XOR U3577 ( .A(n2370), .B(n2369), .Z(n2372) );
  XOR U3578 ( .A(n2371), .B(n2372), .Z(n2365) );
  XOR U3579 ( .A(n2366), .B(n2365), .Z(n2367) );
  XOR U3580 ( .A(n2368), .B(n2367), .Z(n2265) );
  NAND U3581 ( .A(n2233), .B(n2232), .Z(n2237) );
  NAND U3582 ( .A(n2235), .B(n2234), .Z(n2236) );
  NAND U3583 ( .A(n2237), .B(n2236), .Z(n2264) );
  XOR U3584 ( .A(n2265), .B(n2264), .Z(n2267) );
  XNOR U3585 ( .A(n2266), .B(n2267), .Z(n2384) );
  NANDN U3586 ( .A(n2239), .B(n2238), .Z(n2243) );
  NANDN U3587 ( .A(n2241), .B(n2240), .Z(n2242) );
  AND U3588 ( .A(n2243), .B(n2242), .Z(n2383) );
  NANDN U3589 ( .A(n2245), .B(n2244), .Z(n2249) );
  NAND U3590 ( .A(n2247), .B(n2246), .Z(n2248) );
  AND U3591 ( .A(n2249), .B(n2248), .Z(n2382) );
  XOR U3592 ( .A(n2383), .B(n2382), .Z(n2385) );
  XOR U3593 ( .A(n2384), .B(n2385), .Z(n2378) );
  OR U3594 ( .A(n2252), .B(n2250), .Z(n2256) );
  ANDN U3595 ( .B(n2252), .A(n2251), .Z(n2254) );
  OR U3596 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U3597 ( .A(n2256), .B(n2255), .Z(n2377) );
  NAND U3598 ( .A(n2258), .B(n2257), .Z(n2262) );
  NAND U3599 ( .A(n2260), .B(n2259), .Z(n2261) );
  AND U3600 ( .A(n2262), .B(n2261), .Z(n2376) );
  IV U3601 ( .A(n2376), .Z(n2375) );
  XOR U3602 ( .A(n2377), .B(n2375), .Z(n2263) );
  XNOR U3603 ( .A(n2378), .B(n2263), .Z(N54) );
  NAND U3604 ( .A(n2265), .B(n2264), .Z(n2269) );
  NAND U3605 ( .A(n2267), .B(n2266), .Z(n2268) );
  AND U3606 ( .A(n2269), .B(n2268), .Z(n2392) );
  NAND U3607 ( .A(n2271), .B(n2270), .Z(n2275) );
  NAND U3608 ( .A(n2273), .B(n2272), .Z(n2274) );
  NAND U3609 ( .A(n2275), .B(n2274), .Z(n2389) );
  NANDN U3610 ( .A(n2277), .B(n2276), .Z(n2281) );
  NANDN U3611 ( .A(n2279), .B(n2278), .Z(n2280) );
  AND U3612 ( .A(n2281), .B(n2280), .Z(n2502) );
  NAND U3613 ( .A(n2283), .B(n2282), .Z(n2287) );
  NAND U3614 ( .A(n2285), .B(n2284), .Z(n2286) );
  AND U3615 ( .A(n2287), .B(n2286), .Z(n2498) );
  NANDN U3616 ( .A(n2977), .B(n2452), .Z(n2291) );
  NAND U3617 ( .A(n2289), .B(n2288), .Z(n2290) );
  AND U3618 ( .A(n2291), .B(n2290), .Z(n2431) );
  AND U3619 ( .A(y[1809]), .B(x[229]), .Z(n2473) );
  AND U3620 ( .A(x[241]), .B(y[1797]), .Z(n2474) );
  XOR U3621 ( .A(n2473), .B(n2474), .Z(n2475) );
  AND U3622 ( .A(y[1798]), .B(x[240]), .Z(n2476) );
  XOR U3623 ( .A(n2475), .B(n2476), .Z(n2428) );
  AND U3624 ( .A(y[1796]), .B(x[242]), .Z(n2293) );
  NAND U3625 ( .A(y[1802]), .B(x[236]), .Z(n2292) );
  XNOR U3626 ( .A(n2293), .B(n2292), .Z(n2453) );
  AND U3627 ( .A(x[228]), .B(y[1810]), .Z(n2454) );
  XNOR U3628 ( .A(n2453), .B(n2454), .Z(n2429) );
  XNOR U3629 ( .A(n2428), .B(n2429), .Z(n2430) );
  XOR U3630 ( .A(n2431), .B(n2430), .Z(n2495) );
  AND U3631 ( .A(x[243]), .B(y[1802]), .Z(n3493) );
  NAND U3632 ( .A(n3493), .B(n2294), .Z(n2298) );
  NAND U3633 ( .A(n2296), .B(n2295), .Z(n2297) );
  AND U3634 ( .A(n2298), .B(n2297), .Z(n2496) );
  XOR U3635 ( .A(n2495), .B(n2496), .Z(n2497) );
  XOR U3636 ( .A(n2498), .B(n2497), .Z(n2499) );
  NAND U3637 ( .A(n2300), .B(n2299), .Z(n2304) );
  NAND U3638 ( .A(n2302), .B(n2301), .Z(n2303) );
  AND U3639 ( .A(n2304), .B(n2303), .Z(n2486) );
  NAND U3640 ( .A(n2306), .B(n2305), .Z(n2310) );
  NAND U3641 ( .A(n2308), .B(n2307), .Z(n2309) );
  NAND U3642 ( .A(n2310), .B(n2309), .Z(n2485) );
  XNOR U3643 ( .A(n2486), .B(n2485), .Z(n2488) );
  NAND U3644 ( .A(n2312), .B(n2311), .Z(n2316) );
  AND U3645 ( .A(n2314), .B(n2313), .Z(n2315) );
  ANDN U3646 ( .B(n2316), .A(n2315), .Z(n2451) );
  AND U3647 ( .A(x[237]), .B(y[1801]), .Z(n2318) );
  NAND U3648 ( .A(y[1794]), .B(x[244]), .Z(n2317) );
  XNOR U3649 ( .A(n2318), .B(n2317), .Z(n2469) );
  AND U3650 ( .A(y[1812]), .B(x[226]), .Z(n2470) );
  XOR U3651 ( .A(n2469), .B(n2470), .Z(n2449) );
  AND U3652 ( .A(x[230]), .B(y[1808]), .Z(n2320) );
  NAND U3653 ( .A(x[239]), .B(y[1799]), .Z(n2319) );
  XNOR U3654 ( .A(n2320), .B(n2319), .Z(n2481) );
  XOR U3655 ( .A(n2449), .B(n2448), .Z(n2450) );
  XNOR U3656 ( .A(n2451), .B(n2450), .Z(n2489) );
  AND U3657 ( .A(y[1810]), .B(x[237]), .Z(n3779) );
  NANDN U3658 ( .A(n2321), .B(n3779), .Z(n2325) );
  NAND U3659 ( .A(n2323), .B(n2322), .Z(n2324) );
  AND U3660 ( .A(n2325), .B(n2324), .Z(n2421) );
  AND U3661 ( .A(x[225]), .B(y[1813]), .Z(n2442) );
  XOR U3662 ( .A(n2443), .B(n2442), .Z(n2441) );
  AND U3663 ( .A(n2326), .B(o[21]), .Z(n2440) );
  XOR U3664 ( .A(n2441), .B(n2440), .Z(n2419) );
  AND U3665 ( .A(y[1800]), .B(x[238]), .Z(n2434) );
  AND U3666 ( .A(y[1811]), .B(x[227]), .Z(n2435) );
  XOR U3667 ( .A(n2434), .B(n2435), .Z(n2436) );
  AND U3668 ( .A(y[1795]), .B(x[243]), .Z(n2437) );
  XOR U3669 ( .A(n2436), .B(n2437), .Z(n2418) );
  XOR U3670 ( .A(n2419), .B(n2418), .Z(n2420) );
  XNOR U3671 ( .A(n2421), .B(n2420), .Z(n2490) );
  XOR U3672 ( .A(n2489), .B(n2490), .Z(n2492) );
  NAND U3673 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U3674 ( .A(n2330), .B(n2329), .Z(n2331) );
  AND U3675 ( .A(n2332), .B(n2331), .Z(n2415) );
  AND U3676 ( .A(y[1803]), .B(x[242]), .Z(n3495) );
  NAND U3677 ( .A(n3495), .B(n2333), .Z(n2337) );
  NAND U3678 ( .A(n2335), .B(n2334), .Z(n2336) );
  NAND U3679 ( .A(n2337), .B(n2336), .Z(n2414) );
  XNOR U3680 ( .A(n2415), .B(n2414), .Z(n2417) );
  AND U3681 ( .A(x[238]), .B(y[1807]), .Z(n3506) );
  NAND U3682 ( .A(n3506), .B(n2480), .Z(n2340) );
  NAND U3683 ( .A(n2338), .B(n2584), .Z(n2339) );
  NAND U3684 ( .A(n2340), .B(n2339), .Z(n2424) );
  AND U3685 ( .A(x[224]), .B(y[1814]), .Z(n2457) );
  AND U3686 ( .A(x[246]), .B(y[1792]), .Z(n2458) );
  XOR U3687 ( .A(n2457), .B(n2458), .Z(n2460) );
  AND U3688 ( .A(y[1793]), .B(x[245]), .Z(n2479) );
  XOR U3689 ( .A(o[22]), .B(n2479), .Z(n2459) );
  XOR U3690 ( .A(n2460), .B(n2459), .Z(n2423) );
  AND U3691 ( .A(x[231]), .B(y[1807]), .Z(n2342) );
  NAND U3692 ( .A(y[1806]), .B(x[232]), .Z(n2341) );
  XNOR U3693 ( .A(n2342), .B(n2341), .Z(n2464) );
  XOR U3694 ( .A(n2464), .B(n2463), .Z(n2422) );
  XOR U3695 ( .A(n2423), .B(n2422), .Z(n2425) );
  XOR U3696 ( .A(n2424), .B(n2425), .Z(n2416) );
  XOR U3697 ( .A(n2417), .B(n2416), .Z(n2491) );
  XOR U3698 ( .A(n2492), .B(n2491), .Z(n2487) );
  XOR U3699 ( .A(n2488), .B(n2487), .Z(n2500) );
  XOR U3700 ( .A(n2499), .B(n2500), .Z(n2501) );
  XOR U3701 ( .A(n2502), .B(n2501), .Z(n2404) );
  NANDN U3702 ( .A(n2344), .B(n2343), .Z(n2348) );
  NANDN U3703 ( .A(n2346), .B(n2345), .Z(n2347) );
  AND U3704 ( .A(n2348), .B(n2347), .Z(n2403) );
  NANDN U3705 ( .A(n2350), .B(n2349), .Z(n2354) );
  NAND U3706 ( .A(n2352), .B(n2351), .Z(n2353) );
  AND U3707 ( .A(n2354), .B(n2353), .Z(n2410) );
  NANDN U3708 ( .A(n2356), .B(n2355), .Z(n2360) );
  NANDN U3709 ( .A(n2358), .B(n2357), .Z(n2359) );
  AND U3710 ( .A(n2360), .B(n2359), .Z(n2409) );
  XOR U3711 ( .A(n2409), .B(n2408), .Z(n2411) );
  XNOR U3712 ( .A(n2410), .B(n2411), .Z(n2402) );
  XOR U3713 ( .A(n2403), .B(n2402), .Z(n2405) );
  XOR U3714 ( .A(n2404), .B(n2405), .Z(n2400) );
  NAND U3715 ( .A(n2370), .B(n2369), .Z(n2374) );
  NAND U3716 ( .A(n2372), .B(n2371), .Z(n2373) );
  NAND U3717 ( .A(n2374), .B(n2373), .Z(n2398) );
  XNOR U3718 ( .A(n2399), .B(n2398), .Z(n2401) );
  XOR U3719 ( .A(n2400), .B(n2401), .Z(n2390) );
  XOR U3720 ( .A(n2389), .B(n2390), .Z(n2391) );
  XNOR U3721 ( .A(n2392), .B(n2391), .Z(n2395) );
  OR U3722 ( .A(n2377), .B(n2375), .Z(n2381) );
  ANDN U3723 ( .B(n2377), .A(n2376), .Z(n2379) );
  OR U3724 ( .A(n2379), .B(n2378), .Z(n2380) );
  AND U3725 ( .A(n2381), .B(n2380), .Z(n2396) );
  NANDN U3726 ( .A(n2383), .B(n2382), .Z(n2387) );
  NANDN U3727 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U3728 ( .A(n2387), .B(n2386), .Z(n2397) );
  XOR U3729 ( .A(n2396), .B(n2397), .Z(n2388) );
  XNOR U3730 ( .A(n2395), .B(n2388), .Z(N55) );
  NAND U3731 ( .A(n2390), .B(n2389), .Z(n2394) );
  NAND U3732 ( .A(n2392), .B(n2391), .Z(n2393) );
  NAND U3733 ( .A(n2394), .B(n2393), .Z(n2641) );
  NANDN U3734 ( .A(n2403), .B(n2402), .Z(n2407) );
  NANDN U3735 ( .A(n2405), .B(n2404), .Z(n2406) );
  AND U3736 ( .A(n2407), .B(n2406), .Z(n2636) );
  NANDN U3737 ( .A(n2409), .B(n2408), .Z(n2413) );
  OR U3738 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U3739 ( .A(n2413), .B(n2412), .Z(n2620) );
  NAND U3740 ( .A(n2423), .B(n2422), .Z(n2427) );
  NAND U3741 ( .A(n2425), .B(n2424), .Z(n2426) );
  NAND U3742 ( .A(n2427), .B(n2426), .Z(n2564) );
  XOR U3743 ( .A(n2565), .B(n2564), .Z(n2567) );
  XOR U3744 ( .A(n2566), .B(n2567), .Z(n2631) );
  NANDN U3745 ( .A(n2429), .B(n2428), .Z(n2433) );
  NANDN U3746 ( .A(n2431), .B(n2430), .Z(n2432) );
  NAND U3747 ( .A(n2433), .B(n2432), .Z(n2629) );
  NAND U3748 ( .A(n2435), .B(n2434), .Z(n2439) );
  NAND U3749 ( .A(n2437), .B(n2436), .Z(n2438) );
  NAND U3750 ( .A(n2439), .B(n2438), .Z(n2511) );
  AND U3751 ( .A(n2441), .B(n2440), .Z(n2445) );
  NAND U3752 ( .A(n2443), .B(n2442), .Z(n2444) );
  NANDN U3753 ( .A(n2445), .B(n2444), .Z(n2510) );
  XOR U3754 ( .A(n2511), .B(n2510), .Z(n2513) );
  AND U3755 ( .A(x[231]), .B(y[1808]), .Z(n2447) );
  NAND U3756 ( .A(y[1806]), .B(x[233]), .Z(n2446) );
  XNOR U3757 ( .A(n2447), .B(n2446), .Z(n2586) );
  XOR U3758 ( .A(n2585), .B(n2586), .Z(n2516) );
  AND U3759 ( .A(x[234]), .B(y[1805]), .Z(n2517) );
  XOR U3760 ( .A(n2516), .B(n2517), .Z(n2519) );
  AND U3761 ( .A(y[1809]), .B(x[230]), .Z(n2576) );
  AND U3762 ( .A(x[239]), .B(y[1800]), .Z(n2577) );
  XOR U3763 ( .A(n2576), .B(n2577), .Z(n2578) );
  AND U3764 ( .A(y[1804]), .B(x[235]), .Z(n2579) );
  XOR U3765 ( .A(n2578), .B(n2579), .Z(n2518) );
  XOR U3766 ( .A(n2519), .B(n2518), .Z(n2512) );
  XOR U3767 ( .A(n2513), .B(n2512), .Z(n2630) );
  XOR U3768 ( .A(n2629), .B(n2630), .Z(n2632) );
  XOR U3769 ( .A(n2631), .B(n2632), .Z(n2618) );
  NAND U3770 ( .A(x[242]), .B(y[1802]), .Z(n3329) );
  NANDN U3771 ( .A(n3329), .B(n2452), .Z(n2456) );
  NAND U3772 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U3773 ( .A(n2456), .B(n2455), .Z(n2553) );
  NAND U3774 ( .A(n2458), .B(n2457), .Z(n2462) );
  NAND U3775 ( .A(n2460), .B(n2459), .Z(n2461) );
  NAND U3776 ( .A(n2462), .B(n2461), .Z(n2552) );
  XOR U3777 ( .A(n2553), .B(n2552), .Z(n2554) );
  NAND U3778 ( .A(n2584), .B(n2585), .Z(n2466) );
  NAND U3779 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U3780 ( .A(n2466), .B(n2465), .Z(n2548) );
  AND U3781 ( .A(x[224]), .B(y[1815]), .Z(n2595) );
  AND U3782 ( .A(y[1792]), .B(x[247]), .Z(n2596) );
  XOR U3783 ( .A(n2595), .B(n2596), .Z(n2598) );
  AND U3784 ( .A(x[246]), .B(y[1793]), .Z(n2575) );
  XOR U3785 ( .A(o[23]), .B(n2575), .Z(n2597) );
  XOR U3786 ( .A(n2598), .B(n2597), .Z(n2547) );
  AND U3787 ( .A(y[1795]), .B(x[244]), .Z(n3180) );
  NAND U3788 ( .A(x[240]), .B(y[1799]), .Z(n2467) );
  XNOR U3789 ( .A(n3180), .B(n2467), .Z(n2571) );
  AND U3790 ( .A(y[1796]), .B(x[243]), .Z(n2572) );
  XOR U3791 ( .A(n2571), .B(n2572), .Z(n2546) );
  XOR U3792 ( .A(n2547), .B(n2546), .Z(n2549) );
  XNOR U3793 ( .A(n2548), .B(n2549), .Z(n2555) );
  XOR U3794 ( .A(n2612), .B(n2611), .Z(n2614) );
  AND U3795 ( .A(x[244]), .B(y[1801]), .Z(n3517) );
  AND U3796 ( .A(x[237]), .B(y[1794]), .Z(n2468) );
  NAND U3797 ( .A(n3517), .B(n2468), .Z(n2472) );
  NAND U3798 ( .A(n2470), .B(n2469), .Z(n2471) );
  NAND U3799 ( .A(n2472), .B(n2471), .Z(n2606) );
  NAND U3800 ( .A(n2474), .B(n2473), .Z(n2478) );
  NAND U3801 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U3802 ( .A(n2478), .B(n2477), .Z(n2560) );
  AND U3803 ( .A(x[237]), .B(y[1802]), .Z(n2534) );
  AND U3804 ( .A(x[226]), .B(y[1813]), .Z(n2535) );
  XOR U3805 ( .A(n2534), .B(n2535), .Z(n2536) );
  AND U3806 ( .A(x[245]), .B(y[1794]), .Z(n2537) );
  XOR U3807 ( .A(n2536), .B(n2537), .Z(n2559) );
  AND U3808 ( .A(y[1803]), .B(x[236]), .Z(n2589) );
  AND U3809 ( .A(x[225]), .B(y[1814]), .Z(n2590) );
  XOR U3810 ( .A(n2589), .B(n2590), .Z(n2592) );
  AND U3811 ( .A(o[22]), .B(n2479), .Z(n2591) );
  XOR U3812 ( .A(n2592), .B(n2591), .Z(n2558) );
  XOR U3813 ( .A(n2559), .B(n2558), .Z(n2561) );
  XOR U3814 ( .A(n2560), .B(n2561), .Z(n2605) );
  XOR U3815 ( .A(n2606), .B(n2605), .Z(n2608) );
  AND U3816 ( .A(x[239]), .B(y[1808]), .Z(n3732) );
  NAND U3817 ( .A(n3732), .B(n2480), .Z(n2484) );
  NANDN U3818 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U3819 ( .A(n2484), .B(n2483), .Z(n2542) );
  AND U3820 ( .A(y[1801]), .B(x[238]), .Z(n2528) );
  AND U3821 ( .A(y[1812]), .B(x[227]), .Z(n2529) );
  XOR U3822 ( .A(n2528), .B(n2529), .Z(n2530) );
  AND U3823 ( .A(x[228]), .B(y[1811]), .Z(n2531) );
  XOR U3824 ( .A(n2530), .B(n2531), .Z(n2541) );
  AND U3825 ( .A(y[1810]), .B(x[229]), .Z(n2522) );
  AND U3826 ( .A(x[242]), .B(y[1797]), .Z(n2523) );
  XOR U3827 ( .A(n2522), .B(n2523), .Z(n2525) );
  AND U3828 ( .A(x[241]), .B(y[1798]), .Z(n2524) );
  XOR U3829 ( .A(n2525), .B(n2524), .Z(n2540) );
  XOR U3830 ( .A(n2541), .B(n2540), .Z(n2543) );
  XOR U3831 ( .A(n2542), .B(n2543), .Z(n2607) );
  XOR U3832 ( .A(n2608), .B(n2607), .Z(n2613) );
  XOR U3833 ( .A(n2614), .B(n2613), .Z(n2617) );
  XOR U3834 ( .A(n2618), .B(n2617), .Z(n2619) );
  XNOR U3835 ( .A(n2620), .B(n2619), .Z(n2506) );
  NAND U3836 ( .A(n2490), .B(n2489), .Z(n2494) );
  NAND U3837 ( .A(n2492), .B(n2491), .Z(n2493) );
  NAND U3838 ( .A(n2494), .B(n2493), .Z(n2624) );
  XOR U3839 ( .A(n2624), .B(n2623), .Z(n2625) );
  XNOR U3840 ( .A(n2626), .B(n2625), .Z(n2504) );
  XOR U3841 ( .A(n2504), .B(n2505), .Z(n2507) );
  XOR U3842 ( .A(n2506), .B(n2507), .Z(n2635) );
  XOR U3843 ( .A(n2636), .B(n2635), .Z(n2638) );
  XNOR U3844 ( .A(n2637), .B(n2638), .Z(n2643) );
  XNOR U3845 ( .A(n2642), .B(n2643), .Z(n2503) );
  XNOR U3846 ( .A(n2641), .B(n2503), .Z(N56) );
  NAND U3847 ( .A(n2505), .B(n2504), .Z(n2509) );
  NAND U3848 ( .A(n2507), .B(n2506), .Z(n2508) );
  AND U3849 ( .A(n2509), .B(n2508), .Z(n2779) );
  NAND U3850 ( .A(n2511), .B(n2510), .Z(n2515) );
  NAND U3851 ( .A(n2513), .B(n2512), .Z(n2514) );
  NAND U3852 ( .A(n2515), .B(n2514), .Z(n2720) );
  NAND U3853 ( .A(n2517), .B(n2516), .Z(n2521) );
  NAND U3854 ( .A(n2519), .B(n2518), .Z(n2520) );
  NAND U3855 ( .A(n2521), .B(n2520), .Z(n2718) );
  NAND U3856 ( .A(n2523), .B(n2522), .Z(n2527) );
  NAND U3857 ( .A(n2525), .B(n2524), .Z(n2526) );
  NAND U3858 ( .A(n2527), .B(n2526), .Z(n2744) );
  AND U3859 ( .A(y[1816]), .B(x[224]), .Z(n2699) );
  AND U3860 ( .A(y[1792]), .B(x[248]), .Z(n2700) );
  XOR U3861 ( .A(n2699), .B(n2700), .Z(n2701) );
  NAND U3862 ( .A(y[1793]), .B(x[247]), .Z(n2692) );
  XNOR U3863 ( .A(o[24]), .B(n2692), .Z(n2702) );
  XOR U3864 ( .A(n2701), .B(n2702), .Z(n2742) );
  AND U3865 ( .A(y[1809]), .B(x[231]), .Z(n2685) );
  NAND U3866 ( .A(y[1798]), .B(x[242]), .Z(n2686) );
  NAND U3867 ( .A(x[241]), .B(y[1799]), .Z(n2688) );
  XOR U3868 ( .A(n2742), .B(n2741), .Z(n2743) );
  XOR U3869 ( .A(n2744), .B(n2743), .Z(n2732) );
  NAND U3870 ( .A(n2529), .B(n2528), .Z(n2533) );
  NAND U3871 ( .A(n2531), .B(n2530), .Z(n2532) );
  NAND U3872 ( .A(n2533), .B(n2532), .Z(n2730) );
  NAND U3873 ( .A(n2535), .B(n2534), .Z(n2539) );
  NAND U3874 ( .A(n2537), .B(n2536), .Z(n2538) );
  NAND U3875 ( .A(n2539), .B(n2538), .Z(n2729) );
  XOR U3876 ( .A(n2730), .B(n2729), .Z(n2731) );
  XOR U3877 ( .A(n2732), .B(n2731), .Z(n2717) );
  XOR U3878 ( .A(n2718), .B(n2717), .Z(n2719) );
  XNOR U3879 ( .A(n2720), .B(n2719), .Z(n2725) );
  NAND U3880 ( .A(n2541), .B(n2540), .Z(n2545) );
  NAND U3881 ( .A(n2543), .B(n2542), .Z(n2544) );
  AND U3882 ( .A(n2545), .B(n2544), .Z(n2771) );
  NAND U3883 ( .A(n2547), .B(n2546), .Z(n2551) );
  NAND U3884 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U3885 ( .A(n2551), .B(n2550), .Z(n2770) );
  XOR U3886 ( .A(n2771), .B(n2770), .Z(n2773) );
  NAND U3887 ( .A(n2553), .B(n2552), .Z(n2557) );
  NANDN U3888 ( .A(n2555), .B(n2554), .Z(n2556) );
  AND U3889 ( .A(n2557), .B(n2556), .Z(n2772) );
  XOR U3890 ( .A(n2773), .B(n2772), .Z(n2723) );
  NAND U3891 ( .A(n2559), .B(n2558), .Z(n2563) );
  NAND U3892 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U3893 ( .A(n2563), .B(n2562), .Z(n2724) );
  XOR U3894 ( .A(n2723), .B(n2724), .Z(n2726) );
  XOR U3895 ( .A(n2725), .B(n2726), .Z(n2652) );
  NAND U3896 ( .A(n2565), .B(n2564), .Z(n2569) );
  NAND U3897 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U3898 ( .A(n2569), .B(n2568), .Z(n2651) );
  XOR U3899 ( .A(n2652), .B(n2651), .Z(n2654) );
  AND U3900 ( .A(y[1799]), .B(x[244]), .Z(n2570) );
  NAND U3901 ( .A(n2570), .B(n2747), .Z(n2574) );
  NAND U3902 ( .A(n2572), .B(n2571), .Z(n2573) );
  NAND U3903 ( .A(n2574), .B(n2573), .Z(n2767) );
  AND U3904 ( .A(x[246]), .B(y[1794]), .Z(n2673) );
  XOR U3905 ( .A(n2674), .B(n2673), .Z(n2676) );
  NAND U3906 ( .A(x[226]), .B(y[1814]), .Z(n2675) );
  AND U3907 ( .A(x[225]), .B(y[1815]), .Z(n2681) );
  XOR U3908 ( .A(n2682), .B(n2681), .Z(n2680) );
  AND U3909 ( .A(o[23]), .B(n2575), .Z(n2679) );
  XOR U3910 ( .A(n2680), .B(n2679), .Z(n2764) );
  XOR U3911 ( .A(n2765), .B(n2764), .Z(n2766) );
  XOR U3912 ( .A(n2767), .B(n2766), .Z(n2712) );
  NAND U3913 ( .A(n2577), .B(n2576), .Z(n2581) );
  NAND U3914 ( .A(n2579), .B(n2578), .Z(n2580) );
  NAND U3915 ( .A(n2581), .B(n2580), .Z(n2761) );
  AND U3916 ( .A(x[240]), .B(y[1800]), .Z(n2583) );
  NAND U3917 ( .A(y[1795]), .B(x[245]), .Z(n2582) );
  XNOR U3918 ( .A(n2583), .B(n2582), .Z(n2748) );
  AND U3919 ( .A(y[1811]), .B(x[229]), .Z(n2749) );
  XOR U3920 ( .A(n2748), .B(n2749), .Z(n2759) );
  AND U3921 ( .A(y[1810]), .B(x[230]), .Z(n3062) );
  AND U3922 ( .A(x[244]), .B(y[1796]), .Z(n2896) );
  XOR U3923 ( .A(n3062), .B(n2896), .Z(n2754) );
  AND U3924 ( .A(y[1797]), .B(x[243]), .Z(n2755) );
  XOR U3925 ( .A(n2754), .B(n2755), .Z(n2758) );
  XOR U3926 ( .A(n2759), .B(n2758), .Z(n2760) );
  XOR U3927 ( .A(n2761), .B(n2760), .Z(n2738) );
  NAND U3928 ( .A(n2823), .B(n2584), .Z(n2588) );
  NAND U3929 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U3930 ( .A(n2588), .B(n2587), .Z(n2736) );
  NAND U3931 ( .A(n2590), .B(n2589), .Z(n2594) );
  NAND U3932 ( .A(n2592), .B(n2591), .Z(n2593) );
  NAND U3933 ( .A(n2594), .B(n2593), .Z(n2735) );
  XOR U3934 ( .A(n2736), .B(n2735), .Z(n2737) );
  XOR U3935 ( .A(n2738), .B(n2737), .Z(n2711) );
  XOR U3936 ( .A(n2712), .B(n2711), .Z(n2714) );
  NAND U3937 ( .A(n2596), .B(n2595), .Z(n2600) );
  NAND U3938 ( .A(n2598), .B(n2597), .Z(n2599) );
  NAND U3939 ( .A(n2600), .B(n2599), .Z(n2706) );
  AND U3940 ( .A(x[227]), .B(y[1813]), .Z(n2695) );
  XOR U3941 ( .A(n2696), .B(n2695), .Z(n2694) );
  AND U3942 ( .A(x[228]), .B(y[1812]), .Z(n2693) );
  XOR U3943 ( .A(n2694), .B(n2693), .Z(n2705) );
  XOR U3944 ( .A(n2706), .B(n2705), .Z(n2708) );
  AND U3945 ( .A(y[1807]), .B(x[233]), .Z(n2602) );
  NAND U3946 ( .A(y[1806]), .B(x[234]), .Z(n2601) );
  XNOR U3947 ( .A(n2602), .B(n2601), .Z(n2665) );
  AND U3948 ( .A(y[1802]), .B(x[238]), .Z(n2604) );
  NAND U3949 ( .A(y[1808]), .B(x[232]), .Z(n2603) );
  XNOR U3950 ( .A(n2604), .B(n2603), .Z(n2669) );
  AND U3951 ( .A(y[1805]), .B(x[235]), .Z(n2670) );
  XOR U3952 ( .A(n2669), .B(n2670), .Z(n2664) );
  XOR U3953 ( .A(n2665), .B(n2664), .Z(n2707) );
  XOR U3954 ( .A(n2708), .B(n2707), .Z(n2713) );
  XNOR U3955 ( .A(n2714), .B(n2713), .Z(n2658) );
  NAND U3956 ( .A(n2606), .B(n2605), .Z(n2610) );
  NAND U3957 ( .A(n2608), .B(n2607), .Z(n2609) );
  AND U3958 ( .A(n2610), .B(n2609), .Z(n2657) );
  XOR U3959 ( .A(n2658), .B(n2657), .Z(n2659) );
  NAND U3960 ( .A(n2612), .B(n2611), .Z(n2616) );
  NAND U3961 ( .A(n2614), .B(n2613), .Z(n2615) );
  AND U3962 ( .A(n2616), .B(n2615), .Z(n2660) );
  XOR U3963 ( .A(n2659), .B(n2660), .Z(n2653) );
  XNOR U3964 ( .A(n2654), .B(n2653), .Z(n2777) );
  NAND U3965 ( .A(n2618), .B(n2617), .Z(n2622) );
  NAND U3966 ( .A(n2620), .B(n2619), .Z(n2621) );
  NAND U3967 ( .A(n2622), .B(n2621), .Z(n2647) );
  NAND U3968 ( .A(n2624), .B(n2623), .Z(n2628) );
  NAND U3969 ( .A(n2626), .B(n2625), .Z(n2627) );
  NAND U3970 ( .A(n2628), .B(n2627), .Z(n2646) );
  NAND U3971 ( .A(n2630), .B(n2629), .Z(n2634) );
  NAND U3972 ( .A(n2632), .B(n2631), .Z(n2633) );
  NAND U3973 ( .A(n2634), .B(n2633), .Z(n2645) );
  XOR U3974 ( .A(n2646), .B(n2645), .Z(n2648) );
  XOR U3975 ( .A(n2647), .B(n2648), .Z(n2776) );
  XOR U3976 ( .A(n2777), .B(n2776), .Z(n2778) );
  XOR U3977 ( .A(n2779), .B(n2778), .Z(n2784) );
  NANDN U3978 ( .A(n2636), .B(n2635), .Z(n2640) );
  NANDN U3979 ( .A(n2638), .B(n2637), .Z(n2639) );
  AND U3980 ( .A(n2640), .B(n2639), .Z(n2783) );
  XOR U3981 ( .A(n2783), .B(n2782), .Z(n2644) );
  XNOR U3982 ( .A(n2784), .B(n2644), .Z(N57) );
  NAND U3983 ( .A(n2646), .B(n2645), .Z(n2650) );
  NAND U3984 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U3985 ( .A(n2650), .B(n2649), .Z(n2927) );
  NAND U3986 ( .A(n2652), .B(n2651), .Z(n2656) );
  NAND U3987 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U3988 ( .A(n2656), .B(n2655), .Z(n2925) );
  NAND U3989 ( .A(n2658), .B(n2657), .Z(n2662) );
  NAND U3990 ( .A(n2660), .B(n2659), .Z(n2661) );
  AND U3991 ( .A(n2662), .B(n2661), .Z(n2787) );
  NANDN U3992 ( .A(n2822), .B(n2663), .Z(n2667) );
  NAND U3993 ( .A(n2665), .B(n2664), .Z(n2666) );
  NAND U3994 ( .A(n2667), .B(n2666), .Z(n2847) );
  AND U3995 ( .A(x[238]), .B(y[1808]), .Z(n3647) );
  NAND U3996 ( .A(n3647), .B(n2668), .Z(n2672) );
  NAND U3997 ( .A(n2670), .B(n2669), .Z(n2671) );
  NAND U3998 ( .A(n2672), .B(n2671), .Z(n2873) );
  AND U3999 ( .A(y[1806]), .B(x[235]), .Z(n2893) );
  AND U4000 ( .A(x[236]), .B(y[1805]), .Z(n2891) );
  NAND U4001 ( .A(y[1810]), .B(x[231]), .Z(n2890) );
  XNOR U4002 ( .A(n2891), .B(n2890), .Z(n2892) );
  XOR U4003 ( .A(n2893), .B(n2892), .Z(n2871) );
  NAND U4004 ( .A(y[1793]), .B(x[248]), .Z(n2889) );
  XNOR U4005 ( .A(o[25]), .B(n2889), .Z(n2860) );
  AND U4006 ( .A(y[1816]), .B(x[225]), .Z(n2859) );
  XOR U4007 ( .A(n2860), .B(n2859), .Z(n2862) );
  AND U4008 ( .A(y[1804]), .B(x[237]), .Z(n2861) );
  XOR U4009 ( .A(n2862), .B(n2861), .Z(n2872) );
  XOR U4010 ( .A(n2871), .B(n2872), .Z(n2874) );
  XOR U4011 ( .A(n2873), .B(n2874), .Z(n2846) );
  XOR U4012 ( .A(n2847), .B(n2846), .Z(n2849) );
  NAND U4013 ( .A(n2674), .B(n2673), .Z(n2678) );
  ANDN U4014 ( .B(n2676), .A(n2675), .Z(n2677) );
  ANDN U4015 ( .B(n2678), .A(n2677), .Z(n2835) );
  AND U4016 ( .A(n2680), .B(n2679), .Z(n2684) );
  NAND U4017 ( .A(n2682), .B(n2681), .Z(n2683) );
  NANDN U4018 ( .A(n2684), .B(n2683), .Z(n2834) );
  NANDN U4019 ( .A(n2686), .B(n2685), .Z(n2690) );
  NANDN U4020 ( .A(n2688), .B(n2687), .Z(n2689) );
  AND U4021 ( .A(n2690), .B(n2689), .Z(n2831) );
  AND U4022 ( .A(x[232]), .B(y[1809]), .Z(n2825) );
  XOR U4023 ( .A(n2823), .B(n2691), .Z(n2824) );
  XOR U4024 ( .A(n2825), .B(n2824), .Z(n2829) );
  ANDN U4025 ( .B(o[24]), .A(n2692), .Z(n2818) );
  AND U4026 ( .A(y[1792]), .B(x[249]), .Z(n2817) );
  NAND U4027 ( .A(x[224]), .B(y[1817]), .Z(n2816) );
  XOR U4028 ( .A(n2817), .B(n2816), .Z(n2819) );
  XNOR U4029 ( .A(n2818), .B(n2819), .Z(n2828) );
  XOR U4030 ( .A(n2829), .B(n2828), .Z(n2830) );
  XOR U4031 ( .A(n2837), .B(n2836), .Z(n2848) );
  XNOR U4032 ( .A(n2849), .B(n2848), .Z(n2807) );
  AND U4033 ( .A(n2694), .B(n2693), .Z(n2698) );
  NAND U4034 ( .A(n2696), .B(n2695), .Z(n2697) );
  NANDN U4035 ( .A(n2698), .B(n2697), .Z(n2910) );
  NAND U4036 ( .A(n2700), .B(n2699), .Z(n2704) );
  NAND U4037 ( .A(n2702), .B(n2701), .Z(n2703) );
  NAND U4038 ( .A(n2704), .B(n2703), .Z(n2908) );
  AND U4039 ( .A(y[1803]), .B(x[238]), .Z(n2866) );
  AND U4040 ( .A(x[226]), .B(y[1815]), .Z(n2865) );
  XOR U4041 ( .A(n2866), .B(n2865), .Z(n2868) );
  AND U4042 ( .A(x[227]), .B(y[1814]), .Z(n2867) );
  XOR U4043 ( .A(n2868), .B(n2867), .Z(n2907) );
  XOR U4044 ( .A(n2908), .B(n2907), .Z(n2909) );
  XNOR U4045 ( .A(n2910), .B(n2909), .Z(n2805) );
  NAND U4046 ( .A(n2706), .B(n2705), .Z(n2710) );
  NAND U4047 ( .A(n2708), .B(n2707), .Z(n2709) );
  AND U4048 ( .A(n2710), .B(n2709), .Z(n2804) );
  XOR U4049 ( .A(n2805), .B(n2804), .Z(n2806) );
  XOR U4050 ( .A(n2807), .B(n2806), .Z(n2798) );
  NAND U4051 ( .A(n2712), .B(n2711), .Z(n2716) );
  NAND U4052 ( .A(n2714), .B(n2713), .Z(n2715) );
  AND U4053 ( .A(n2716), .B(n2715), .Z(n2799) );
  XOR U4054 ( .A(n2798), .B(n2799), .Z(n2800) );
  NAND U4055 ( .A(n2718), .B(n2717), .Z(n2722) );
  NAND U4056 ( .A(n2720), .B(n2719), .Z(n2721) );
  AND U4057 ( .A(n2722), .B(n2721), .Z(n2801) );
  XOR U4058 ( .A(n2800), .B(n2801), .Z(n2786) );
  NAND U4059 ( .A(n2724), .B(n2723), .Z(n2728) );
  NAND U4060 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U4061 ( .A(n2728), .B(n2727), .Z(n2794) );
  NAND U4062 ( .A(n2730), .B(n2729), .Z(n2734) );
  NAND U4063 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U4064 ( .A(n2734), .B(n2733), .Z(n2811) );
  NAND U4065 ( .A(n2736), .B(n2735), .Z(n2740) );
  NAND U4066 ( .A(n2738), .B(n2737), .Z(n2739) );
  NAND U4067 ( .A(n2740), .B(n2739), .Z(n2810) );
  XOR U4068 ( .A(n2811), .B(n2810), .Z(n2813) );
  NAND U4069 ( .A(n2742), .B(n2741), .Z(n2746) );
  NAND U4070 ( .A(n2744), .B(n2743), .Z(n2745) );
  AND U4071 ( .A(n2746), .B(n2745), .Z(n2843) );
  AND U4072 ( .A(x[245]), .B(y[1800]), .Z(n3774) );
  NAND U4073 ( .A(n3774), .B(n2747), .Z(n2751) );
  NAND U4074 ( .A(n2749), .B(n2748), .Z(n2750) );
  NAND U4075 ( .A(n2751), .B(n2750), .Z(n2916) );
  AND U4076 ( .A(x[246]), .B(y[1795]), .Z(n2885) );
  AND U4077 ( .A(y[1812]), .B(x[229]), .Z(n2884) );
  NAND U4078 ( .A(x[241]), .B(y[1800]), .Z(n2883) );
  XOR U4079 ( .A(n2884), .B(n2883), .Z(n2886) );
  XNOR U4080 ( .A(n2885), .B(n2886), .Z(n2914) );
  AND U4081 ( .A(y[1797]), .B(x[244]), .Z(n2753) );
  NAND U4082 ( .A(y[1796]), .B(x[245]), .Z(n2752) );
  XNOR U4083 ( .A(n2753), .B(n2752), .Z(n2898) );
  AND U4084 ( .A(y[1798]), .B(x[243]), .Z(n2897) );
  XOR U4085 ( .A(n2898), .B(n2897), .Z(n2913) );
  XOR U4086 ( .A(n2914), .B(n2913), .Z(n2915) );
  XNOR U4087 ( .A(n2916), .B(n2915), .Z(n2841) );
  NAND U4088 ( .A(n2896), .B(n3062), .Z(n2757) );
  NAND U4089 ( .A(n2755), .B(n2754), .Z(n2756) );
  AND U4090 ( .A(n2757), .B(n2756), .Z(n2922) );
  AND U4091 ( .A(x[239]), .B(y[1802]), .Z(n2903) );
  AND U4092 ( .A(y[1799]), .B(x[242]), .Z(n2902) );
  NAND U4093 ( .A(y[1811]), .B(x[230]), .Z(n2901) );
  XOR U4094 ( .A(n2902), .B(n2901), .Z(n2904) );
  XNOR U4095 ( .A(n2903), .B(n2904), .Z(n2920) );
  AND U4096 ( .A(x[247]), .B(y[1794]), .Z(n2879) );
  AND U4097 ( .A(x[228]), .B(y[1813]), .Z(n2878) );
  NAND U4098 ( .A(y[1801]), .B(x[240]), .Z(n2877) );
  XOR U4099 ( .A(n2878), .B(n2877), .Z(n2880) );
  XNOR U4100 ( .A(n2879), .B(n2880), .Z(n2919) );
  XOR U4101 ( .A(n2920), .B(n2919), .Z(n2921) );
  XOR U4102 ( .A(n2922), .B(n2921), .Z(n2840) );
  XOR U4103 ( .A(n2841), .B(n2840), .Z(n2842) );
  XNOR U4104 ( .A(n2843), .B(n2842), .Z(n2855) );
  NAND U4105 ( .A(n2759), .B(n2758), .Z(n2763) );
  NAND U4106 ( .A(n2761), .B(n2760), .Z(n2762) );
  NAND U4107 ( .A(n2763), .B(n2762), .Z(n2853) );
  NAND U4108 ( .A(n2765), .B(n2764), .Z(n2769) );
  NAND U4109 ( .A(n2767), .B(n2766), .Z(n2768) );
  NAND U4110 ( .A(n2769), .B(n2768), .Z(n2852) );
  XOR U4111 ( .A(n2853), .B(n2852), .Z(n2854) );
  XOR U4112 ( .A(n2855), .B(n2854), .Z(n2812) );
  XOR U4113 ( .A(n2813), .B(n2812), .Z(n2793) );
  NAND U4114 ( .A(n2771), .B(n2770), .Z(n2775) );
  NAND U4115 ( .A(n2773), .B(n2772), .Z(n2774) );
  NAND U4116 ( .A(n2775), .B(n2774), .Z(n2792) );
  XOR U4117 ( .A(n2794), .B(n2795), .Z(n2788) );
  XOR U4118 ( .A(n2789), .B(n2788), .Z(n2926) );
  XOR U4119 ( .A(n2925), .B(n2926), .Z(n2928) );
  XOR U4120 ( .A(n2927), .B(n2928), .Z(n2933) );
  NAND U4121 ( .A(n2777), .B(n2776), .Z(n2781) );
  NAND U4122 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U4123 ( .A(n2781), .B(n2780), .Z(n2932) );
  XOR U4124 ( .A(n2932), .B(n2931), .Z(n2785) );
  XNOR U4125 ( .A(n2933), .B(n2785), .Z(N58) );
  NANDN U4126 ( .A(n2787), .B(n2786), .Z(n2791) );
  NAND U4127 ( .A(n2789), .B(n2788), .Z(n2790) );
  AND U4128 ( .A(n2791), .B(n2790), .Z(n3082) );
  NANDN U4129 ( .A(n2793), .B(n2792), .Z(n2797) );
  NAND U4130 ( .A(n2795), .B(n2794), .Z(n2796) );
  NAND U4131 ( .A(n2797), .B(n2796), .Z(n3083) );
  NAND U4132 ( .A(n2799), .B(n2798), .Z(n2803) );
  NAND U4133 ( .A(n2801), .B(n2800), .Z(n2802) );
  AND U4134 ( .A(n2803), .B(n2802), .Z(n2935) );
  NAND U4135 ( .A(n2805), .B(n2804), .Z(n2809) );
  NAND U4136 ( .A(n2807), .B(n2806), .Z(n2808) );
  AND U4137 ( .A(n2809), .B(n2808), .Z(n2936) );
  XOR U4138 ( .A(n2935), .B(n2936), .Z(n2938) );
  NAND U4139 ( .A(n2811), .B(n2810), .Z(n2815) );
  NAND U4140 ( .A(n2813), .B(n2812), .Z(n2814) );
  NAND U4141 ( .A(n2815), .B(n2814), .Z(n2944) );
  AND U4142 ( .A(y[1816]), .B(x[226]), .Z(n2965) );
  XOR U4143 ( .A(n2966), .B(n2965), .Z(n2968) );
  NAND U4144 ( .A(x[248]), .B(y[1794]), .Z(n2967) );
  XNOR U4145 ( .A(n2968), .B(n2967), .Z(n3001) );
  NANDN U4146 ( .A(n2817), .B(n2816), .Z(n2821) );
  OR U4147 ( .A(n2819), .B(n2818), .Z(n2820) );
  NAND U4148 ( .A(n2821), .B(n2820), .Z(n3002) );
  XNOR U4149 ( .A(n3001), .B(n3002), .Z(n3004) );
  NANDN U4150 ( .A(n2823), .B(n2822), .Z(n2827) );
  NANDN U4151 ( .A(n2825), .B(n2824), .Z(n2826) );
  AND U4152 ( .A(n2827), .B(n2826), .Z(n3003) );
  XOR U4153 ( .A(n3004), .B(n3003), .Z(n3039) );
  NAND U4154 ( .A(n2829), .B(n2828), .Z(n2833) );
  NANDN U4155 ( .A(n2831), .B(n2830), .Z(n2832) );
  AND U4156 ( .A(n2833), .B(n2832), .Z(n3038) );
  NANDN U4157 ( .A(n2835), .B(n2834), .Z(n2839) );
  NAND U4158 ( .A(n2837), .B(n2836), .Z(n2838) );
  NAND U4159 ( .A(n2839), .B(n2838), .Z(n3041) );
  NAND U4160 ( .A(n2841), .B(n2840), .Z(n2845) );
  NAND U4161 ( .A(n2843), .B(n2842), .Z(n2844) );
  NAND U4162 ( .A(n2845), .B(n2844), .Z(n3033) );
  NAND U4163 ( .A(n2847), .B(n2846), .Z(n2851) );
  NAND U4164 ( .A(n2849), .B(n2848), .Z(n2850) );
  AND U4165 ( .A(n2851), .B(n2850), .Z(n3032) );
  XOR U4166 ( .A(n3033), .B(n3032), .Z(n3034) );
  XNOR U4167 ( .A(n3035), .B(n3034), .Z(n2942) );
  NAND U4168 ( .A(n2853), .B(n2852), .Z(n2857) );
  NAND U4169 ( .A(n2855), .B(n2854), .Z(n2856) );
  NAND U4170 ( .A(n2857), .B(n2856), .Z(n2950) );
  AND U4171 ( .A(x[236]), .B(y[1806]), .Z(n3151) );
  AND U4172 ( .A(y[1813]), .B(x[229]), .Z(n3015) );
  XOR U4173 ( .A(n3151), .B(n3015), .Z(n3017) );
  NAND U4174 ( .A(x[234]), .B(y[1808]), .Z(n3016) );
  XNOR U4175 ( .A(n3017), .B(n3016), .Z(n3047) );
  AND U4176 ( .A(y[1811]), .B(x[231]), .Z(n3044) );
  NAND U4177 ( .A(x[230]), .B(y[1812]), .Z(n2858) );
  XNOR U4178 ( .A(n3291), .B(n2858), .Z(n3063) );
  NAND U4179 ( .A(x[233]), .B(y[1809]), .Z(n3064) );
  XOR U4180 ( .A(n3063), .B(n3064), .Z(n3045) );
  XOR U4181 ( .A(n3047), .B(n3046), .Z(n2991) );
  NAND U4182 ( .A(n2860), .B(n2859), .Z(n2864) );
  NAND U4183 ( .A(n2862), .B(n2861), .Z(n2863) );
  NAND U4184 ( .A(n2864), .B(n2863), .Z(n2990) );
  NAND U4185 ( .A(n2866), .B(n2865), .Z(n2870) );
  NAND U4186 ( .A(n2868), .B(n2867), .Z(n2869) );
  NAND U4187 ( .A(n2870), .B(n2869), .Z(n2989) );
  XOR U4188 ( .A(n2990), .B(n2989), .Z(n2992) );
  XNOR U4189 ( .A(n2991), .B(n2992), .Z(n3027) );
  NAND U4190 ( .A(n2872), .B(n2871), .Z(n2876) );
  NAND U4191 ( .A(n2874), .B(n2873), .Z(n2875) );
  AND U4192 ( .A(n2876), .B(n2875), .Z(n3026) );
  XOR U4193 ( .A(n3027), .B(n3026), .Z(n3029) );
  NANDN U4194 ( .A(n2878), .B(n2877), .Z(n2882) );
  OR U4195 ( .A(n2880), .B(n2879), .Z(n2881) );
  AND U4196 ( .A(n2882), .B(n2881), .Z(n2953) );
  NANDN U4197 ( .A(n2884), .B(n2883), .Z(n2888) );
  OR U4198 ( .A(n2886), .B(n2885), .Z(n2887) );
  NAND U4199 ( .A(n2888), .B(n2887), .Z(n2954) );
  XNOR U4200 ( .A(n2953), .B(n2954), .Z(n2955) );
  ANDN U4201 ( .B(o[25]), .A(n2889), .Z(n3056) );
  NAND U4202 ( .A(y[1804]), .B(x[238]), .Z(n3057) );
  XNOR U4203 ( .A(n3056), .B(n3057), .Z(n3058) );
  NAND U4204 ( .A(x[225]), .B(y[1817]), .Z(n3059) );
  XNOR U4205 ( .A(n3058), .B(n3059), .Z(n3007) );
  NAND U4206 ( .A(y[1793]), .B(x[249]), .Z(n3067) );
  XNOR U4207 ( .A(o[26]), .B(n3067), .Z(n3020) );
  NAND U4208 ( .A(y[1792]), .B(x[250]), .Z(n3021) );
  XNOR U4209 ( .A(n3020), .B(n3021), .Z(n3022) );
  NAND U4210 ( .A(x[224]), .B(y[1818]), .Z(n3023) );
  XOR U4211 ( .A(n3022), .B(n3023), .Z(n3008) );
  XNOR U4212 ( .A(n3007), .B(n3008), .Z(n3009) );
  NANDN U4213 ( .A(n2891), .B(n2890), .Z(n2895) );
  NANDN U4214 ( .A(n2893), .B(n2892), .Z(n2894) );
  NAND U4215 ( .A(n2895), .B(n2894), .Z(n3010) );
  XOR U4216 ( .A(n3009), .B(n3010), .Z(n2956) );
  XOR U4217 ( .A(n2955), .B(n2956), .Z(n2997) );
  AND U4218 ( .A(x[245]), .B(y[1797]), .Z(n3050) );
  NAND U4219 ( .A(n2896), .B(n3050), .Z(n2900) );
  NAND U4220 ( .A(n2898), .B(n2897), .Z(n2899) );
  NAND U4221 ( .A(n2900), .B(n2899), .Z(n2985) );
  XOR U4222 ( .A(n3051), .B(n3050), .Z(n3053) );
  NAND U4223 ( .A(y[1798]), .B(x[244]), .Z(n3052) );
  XNOR U4224 ( .A(n3053), .B(n3052), .Z(n2984) );
  NAND U4225 ( .A(y[1795]), .B(x[247]), .Z(n2972) );
  XNOR U4226 ( .A(n2971), .B(n2972), .Z(n2974) );
  AND U4227 ( .A(x[246]), .B(y[1796]), .Z(n2973) );
  XOR U4228 ( .A(n2974), .B(n2973), .Z(n2983) );
  XOR U4229 ( .A(n2984), .B(n2983), .Z(n2986) );
  XNOR U4230 ( .A(n2985), .B(n2986), .Z(n2996) );
  AND U4231 ( .A(x[228]), .B(y[1814]), .Z(n2979) );
  XOR U4232 ( .A(n2980), .B(n2979), .Z(n2978) );
  AND U4233 ( .A(y[1799]), .B(x[243]), .Z(n3068) );
  NAND U4234 ( .A(y[1807]), .B(x[235]), .Z(n3069) );
  XNOR U4235 ( .A(n3068), .B(n3069), .Z(n3070) );
  NAND U4236 ( .A(x[227]), .B(y[1815]), .Z(n3071) );
  XOR U4237 ( .A(n3070), .B(n3071), .Z(n2960) );
  XNOR U4238 ( .A(n2959), .B(n2960), .Z(n2962) );
  NANDN U4239 ( .A(n2902), .B(n2901), .Z(n2906) );
  OR U4240 ( .A(n2904), .B(n2903), .Z(n2905) );
  AND U4241 ( .A(n2906), .B(n2905), .Z(n2961) );
  XNOR U4242 ( .A(n2962), .B(n2961), .Z(n2995) );
  XOR U4243 ( .A(n2996), .B(n2995), .Z(n2998) );
  XOR U4244 ( .A(n2997), .B(n2998), .Z(n3028) );
  XNOR U4245 ( .A(n3029), .B(n3028), .Z(n2948) );
  NAND U4246 ( .A(n2908), .B(n2907), .Z(n2912) );
  NAND U4247 ( .A(n2910), .B(n2909), .Z(n2911) );
  AND U4248 ( .A(n2912), .B(n2911), .Z(n3079) );
  NAND U4249 ( .A(n2914), .B(n2913), .Z(n2918) );
  NAND U4250 ( .A(n2916), .B(n2915), .Z(n2917) );
  AND U4251 ( .A(n2918), .B(n2917), .Z(n3077) );
  NAND U4252 ( .A(n2920), .B(n2919), .Z(n2924) );
  NANDN U4253 ( .A(n2922), .B(n2921), .Z(n2923) );
  NAND U4254 ( .A(n2924), .B(n2923), .Z(n3076) );
  XOR U4255 ( .A(n2948), .B(n2947), .Z(n2949) );
  XOR U4256 ( .A(n2950), .B(n2949), .Z(n2941) );
  XOR U4257 ( .A(n2942), .B(n2941), .Z(n2943) );
  XOR U4258 ( .A(n2944), .B(n2943), .Z(n2937) );
  XOR U4259 ( .A(n2938), .B(n2937), .Z(n3084) );
  XNOR U4260 ( .A(n3085), .B(n3084), .Z(n3090) );
  NAND U4261 ( .A(n2926), .B(n2925), .Z(n2930) );
  NAND U4262 ( .A(n2928), .B(n2927), .Z(n2929) );
  AND U4263 ( .A(n2930), .B(n2929), .Z(n3088) );
  XNOR U4264 ( .A(n3088), .B(n3089), .Z(n2934) );
  XNOR U4265 ( .A(n3090), .B(n2934), .Z(N59) );
  NAND U4266 ( .A(n2936), .B(n2935), .Z(n2940) );
  NAND U4267 ( .A(n2938), .B(n2937), .Z(n2939) );
  AND U4268 ( .A(n2940), .B(n2939), .Z(n3095) );
  NAND U4269 ( .A(n2942), .B(n2941), .Z(n2946) );
  NAND U4270 ( .A(n2944), .B(n2943), .Z(n2945) );
  AND U4271 ( .A(n2946), .B(n2945), .Z(n3093) );
  NAND U4272 ( .A(n2948), .B(n2947), .Z(n2952) );
  NAND U4273 ( .A(n2950), .B(n2949), .Z(n2951) );
  NAND U4274 ( .A(n2952), .B(n2951), .Z(n3103) );
  NANDN U4275 ( .A(n2954), .B(n2953), .Z(n2958) );
  NANDN U4276 ( .A(n2956), .B(n2955), .Z(n2957) );
  AND U4277 ( .A(n2958), .B(n2957), .Z(n3221) );
  NANDN U4278 ( .A(n2960), .B(n2959), .Z(n2964) );
  NAND U4279 ( .A(n2962), .B(n2961), .Z(n2963) );
  AND U4280 ( .A(n2964), .B(n2963), .Z(n3219) );
  NAND U4281 ( .A(n2966), .B(n2965), .Z(n2970) );
  ANDN U4282 ( .B(n2968), .A(n2967), .Z(n2969) );
  ANDN U4283 ( .B(n2970), .A(n2969), .Z(n3126) );
  NANDN U4284 ( .A(n2972), .B(n2971), .Z(n2976) );
  NAND U4285 ( .A(n2974), .B(n2973), .Z(n2975) );
  NAND U4286 ( .A(n2976), .B(n2975), .Z(n3125) );
  XNOR U4287 ( .A(n3126), .B(n3125), .Z(n3128) );
  ANDN U4288 ( .B(n2978), .A(n2977), .Z(n2982) );
  NAND U4289 ( .A(n2980), .B(n2979), .Z(n2981) );
  NANDN U4290 ( .A(n2982), .B(n2981), .Z(n3138) );
  AND U4291 ( .A(x[224]), .B(y[1819]), .Z(n3206) );
  NAND U4292 ( .A(y[1792]), .B(x[251]), .Z(n3207) );
  XNOR U4293 ( .A(n3206), .B(n3207), .Z(n3208) );
  NAND U4294 ( .A(x[250]), .B(y[1793]), .Z(n3197) );
  XOR U4295 ( .A(o[27]), .B(n3197), .Z(n3209) );
  XNOR U4296 ( .A(n3208), .B(n3209), .Z(n3135) );
  AND U4297 ( .A(y[1810]), .B(x[233]), .Z(n3191) );
  NAND U4298 ( .A(y[1798]), .B(x[245]), .Z(n3192) );
  XNOR U4299 ( .A(n3191), .B(n3192), .Z(n3193) );
  NAND U4300 ( .A(y[1801]), .B(x[242]), .Z(n3194) );
  XNOR U4301 ( .A(n3193), .B(n3194), .Z(n3136) );
  XOR U4302 ( .A(n3135), .B(n3136), .Z(n3137) );
  XOR U4303 ( .A(n3138), .B(n3137), .Z(n3127) );
  XOR U4304 ( .A(n3128), .B(n3127), .Z(n3218) );
  XNOR U4305 ( .A(n3219), .B(n3218), .Z(n3220) );
  XOR U4306 ( .A(n3221), .B(n3220), .Z(n3238) );
  NAND U4307 ( .A(n2984), .B(n2983), .Z(n2988) );
  NAND U4308 ( .A(n2986), .B(n2985), .Z(n2987) );
  AND U4309 ( .A(n2988), .B(n2987), .Z(n3237) );
  NAND U4310 ( .A(n2990), .B(n2989), .Z(n2994) );
  NAND U4311 ( .A(n2992), .B(n2991), .Z(n2993) );
  AND U4312 ( .A(n2994), .B(n2993), .Z(n3236) );
  XOR U4313 ( .A(n3237), .B(n3236), .Z(n3239) );
  XNOR U4314 ( .A(n3238), .B(n3239), .Z(n3102) );
  NAND U4315 ( .A(n2996), .B(n2995), .Z(n3000) );
  NAND U4316 ( .A(n2998), .B(n2997), .Z(n2999) );
  AND U4317 ( .A(n3000), .B(n2999), .Z(n3225) );
  NANDN U4318 ( .A(n3002), .B(n3001), .Z(n3006) );
  NAND U4319 ( .A(n3004), .B(n3003), .Z(n3005) );
  AND U4320 ( .A(n3006), .B(n3005), .Z(n3214) );
  NANDN U4321 ( .A(n3008), .B(n3007), .Z(n3012) );
  NANDN U4322 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U4323 ( .A(n3012), .B(n3011), .Z(n3213) );
  AND U4324 ( .A(y[1800]), .B(x[243]), .Z(n3185) );
  NAND U4325 ( .A(x[249]), .B(y[1794]), .Z(n3186) );
  XNOR U4326 ( .A(n3185), .B(n3186), .Z(n3187) );
  NAND U4327 ( .A(y[1813]), .B(x[230]), .Z(n3188) );
  XNOR U4328 ( .A(n3187), .B(n3188), .Z(n3177) );
  AND U4329 ( .A(x[239]), .B(y[1804]), .Z(n3156) );
  AND U4330 ( .A(x[226]), .B(y[1817]), .Z(n3157) );
  XOR U4331 ( .A(n3156), .B(n3157), .Z(n3158) );
  AND U4332 ( .A(y[1816]), .B(x[227]), .Z(n3159) );
  XOR U4333 ( .A(n3158), .B(n3159), .Z(n3176) );
  XOR U4334 ( .A(n3177), .B(n3176), .Z(n3179) );
  NAND U4335 ( .A(y[1803]), .B(x[240]), .Z(n3142) );
  XNOR U4336 ( .A(n3142), .B(n3141), .Z(n3144) );
  XOR U4337 ( .A(n3143), .B(n3144), .Z(n3152) );
  AND U4338 ( .A(x[237]), .B(y[1806]), .Z(n3014) );
  NAND U4339 ( .A(y[1807]), .B(x[236]), .Z(n3013) );
  XNOR U4340 ( .A(n3014), .B(n3013), .Z(n3153) );
  XOR U4341 ( .A(n3152), .B(n3153), .Z(n3178) );
  XOR U4342 ( .A(n3179), .B(n3178), .Z(n3121) );
  NAND U4343 ( .A(n3151), .B(n3015), .Z(n3019) );
  ANDN U4344 ( .B(n3017), .A(n3016), .Z(n3018) );
  ANDN U4345 ( .B(n3019), .A(n3018), .Z(n3120) );
  NANDN U4346 ( .A(n3021), .B(n3020), .Z(n3025) );
  NANDN U4347 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U4348 ( .A(n3025), .B(n3024), .Z(n3119) );
  XOR U4349 ( .A(n3120), .B(n3119), .Z(n3122) );
  XNOR U4350 ( .A(n3121), .B(n3122), .Z(n3212) );
  XOR U4351 ( .A(n3213), .B(n3212), .Z(n3215) );
  XOR U4352 ( .A(n3214), .B(n3215), .Z(n3224) );
  XOR U4353 ( .A(n3225), .B(n3224), .Z(n3227) );
  NAND U4354 ( .A(n3027), .B(n3026), .Z(n3031) );
  NAND U4355 ( .A(n3029), .B(n3028), .Z(n3030) );
  AND U4356 ( .A(n3031), .B(n3030), .Z(n3226) );
  XOR U4357 ( .A(n3227), .B(n3226), .Z(n3101) );
  XNOR U4358 ( .A(n3102), .B(n3101), .Z(n3104) );
  XOR U4359 ( .A(n3103), .B(n3104), .Z(n3109) );
  NAND U4360 ( .A(n3033), .B(n3032), .Z(n3037) );
  NAND U4361 ( .A(n3035), .B(n3034), .Z(n3036) );
  NAND U4362 ( .A(n3037), .B(n3036), .Z(n3108) );
  NANDN U4363 ( .A(n3039), .B(n3038), .Z(n3043) );
  NANDN U4364 ( .A(n3041), .B(n3040), .Z(n3042) );
  NAND U4365 ( .A(n3043), .B(n3042), .Z(n3114) );
  NANDN U4366 ( .A(n3045), .B(n3044), .Z(n3049) );
  NAND U4367 ( .A(n3047), .B(n3046), .Z(n3048) );
  NAND U4368 ( .A(n3049), .B(n3048), .Z(n3232) );
  NAND U4369 ( .A(n3051), .B(n3050), .Z(n3055) );
  ANDN U4370 ( .B(n3053), .A(n3052), .Z(n3054) );
  ANDN U4371 ( .B(n3055), .A(n3054), .Z(n3169) );
  NANDN U4372 ( .A(n3057), .B(n3056), .Z(n3061) );
  NANDN U4373 ( .A(n3059), .B(n3058), .Z(n3060) );
  NAND U4374 ( .A(n3061), .B(n3060), .Z(n3168) );
  XNOR U4375 ( .A(n3169), .B(n3168), .Z(n3171) );
  AND U4376 ( .A(y[1812]), .B(x[232]), .Z(n3199) );
  NAND U4377 ( .A(n3199), .B(n3062), .Z(n3066) );
  NANDN U4378 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U4379 ( .A(n3066), .B(n3065), .Z(n3131) );
  AND U4380 ( .A(x[238]), .B(y[1805]), .Z(n3162) );
  AND U4381 ( .A(x[225]), .B(y[1818]), .Z(n3163) );
  XOR U4382 ( .A(n3162), .B(n3163), .Z(n3165) );
  ANDN U4383 ( .B(o[26]), .A(n3067), .Z(n3164) );
  XOR U4384 ( .A(n3165), .B(n3164), .Z(n3130) );
  AND U4385 ( .A(x[241]), .B(y[1802]), .Z(n3200) );
  NAND U4386 ( .A(x[228]), .B(y[1815]), .Z(n3201) );
  XNOR U4387 ( .A(n3200), .B(n3201), .Z(n3203) );
  AND U4388 ( .A(y[1814]), .B(x[229]), .Z(n3202) );
  XOR U4389 ( .A(n3203), .B(n3202), .Z(n3129) );
  XOR U4390 ( .A(n3130), .B(n3129), .Z(n3132) );
  XOR U4391 ( .A(n3131), .B(n3132), .Z(n3170) );
  XOR U4392 ( .A(n3171), .B(n3170), .Z(n3231) );
  NANDN U4393 ( .A(n3069), .B(n3068), .Z(n3073) );
  NANDN U4394 ( .A(n3071), .B(n3070), .Z(n3072) );
  AND U4395 ( .A(n3073), .B(n3072), .Z(n3175) );
  AND U4396 ( .A(y[1795]), .B(x[248]), .Z(n3075) );
  NAND U4397 ( .A(x[244]), .B(y[1799]), .Z(n3074) );
  XNOR U4398 ( .A(n3075), .B(n3074), .Z(n3181) );
  NAND U4399 ( .A(y[1812]), .B(x[231]), .Z(n3182) );
  XNOR U4400 ( .A(n3181), .B(n3182), .Z(n3173) );
  AND U4401 ( .A(x[232]), .B(y[1811]), .Z(n3145) );
  AND U4402 ( .A(y[1796]), .B(x[247]), .Z(n3146) );
  XOR U4403 ( .A(n3145), .B(n3146), .Z(n3147) );
  AND U4404 ( .A(x[246]), .B(y[1797]), .Z(n3148) );
  XOR U4405 ( .A(n3147), .B(n3148), .Z(n3172) );
  XOR U4406 ( .A(n3173), .B(n3172), .Z(n3174) );
  XNOR U4407 ( .A(n3175), .B(n3174), .Z(n3230) );
  XOR U4408 ( .A(n3231), .B(n3230), .Z(n3233) );
  XNOR U4409 ( .A(n3232), .B(n3233), .Z(n3113) );
  XOR U4410 ( .A(n3114), .B(n3113), .Z(n3116) );
  NANDN U4411 ( .A(n3077), .B(n3076), .Z(n3081) );
  NANDN U4412 ( .A(n3079), .B(n3078), .Z(n3080) );
  AND U4413 ( .A(n3081), .B(n3080), .Z(n3115) );
  XOR U4414 ( .A(n3116), .B(n3115), .Z(n3107) );
  XOR U4415 ( .A(n3108), .B(n3107), .Z(n3110) );
  XOR U4416 ( .A(n3109), .B(n3110), .Z(n3092) );
  XOR U4417 ( .A(n3093), .B(n3092), .Z(n3094) );
  XOR U4418 ( .A(n3095), .B(n3094), .Z(n3100) );
  NANDN U4419 ( .A(n3083), .B(n3082), .Z(n3087) );
  NAND U4420 ( .A(n3085), .B(n3084), .Z(n3086) );
  NAND U4421 ( .A(n3087), .B(n3086), .Z(n3098) );
  XOR U4422 ( .A(n3098), .B(n3099), .Z(n3091) );
  XNOR U4423 ( .A(n3100), .B(n3091), .Z(N60) );
  NAND U4424 ( .A(n3093), .B(n3092), .Z(n3097) );
  NAND U4425 ( .A(n3095), .B(n3094), .Z(n3096) );
  NAND U4426 ( .A(n3097), .B(n3096), .Z(n3409) );
  IV U4427 ( .A(n3409), .Z(n3407) );
  NAND U4428 ( .A(n3102), .B(n3101), .Z(n3106) );
  NANDN U4429 ( .A(n3104), .B(n3103), .Z(n3105) );
  NAND U4430 ( .A(n3106), .B(n3105), .Z(n3402) );
  NAND U4431 ( .A(n3108), .B(n3107), .Z(n3112) );
  NAND U4432 ( .A(n3110), .B(n3109), .Z(n3111) );
  AND U4433 ( .A(n3112), .B(n3111), .Z(n3401) );
  XOR U4434 ( .A(n3402), .B(n3401), .Z(n3404) );
  NAND U4435 ( .A(n3114), .B(n3113), .Z(n3118) );
  NAND U4436 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U4437 ( .A(n3118), .B(n3117), .Z(n3243) );
  NANDN U4438 ( .A(n3120), .B(n3119), .Z(n3124) );
  NANDN U4439 ( .A(n3122), .B(n3121), .Z(n3123) );
  NAND U4440 ( .A(n3124), .B(n3123), .Z(n3268) );
  NAND U4441 ( .A(n3130), .B(n3129), .Z(n3134) );
  NAND U4442 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U4443 ( .A(n3134), .B(n3133), .Z(n3372) );
  NAND U4444 ( .A(n3136), .B(n3135), .Z(n3140) );
  NAND U4445 ( .A(n3138), .B(n3137), .Z(n3139) );
  NAND U4446 ( .A(n3140), .B(n3139), .Z(n3371) );
  XOR U4447 ( .A(n3372), .B(n3371), .Z(n3373) );
  XOR U4448 ( .A(n3374), .B(n3373), .Z(n3267) );
  XOR U4449 ( .A(n3268), .B(n3267), .Z(n3270) );
  AND U4450 ( .A(x[231]), .B(y[1813]), .Z(n3314) );
  AND U4451 ( .A(x[236]), .B(y[1808]), .Z(n3315) );
  XOR U4452 ( .A(n3314), .B(n3315), .Z(n3317) );
  AND U4453 ( .A(y[1809]), .B(x[235]), .Z(n3316) );
  XNOR U4454 ( .A(n3317), .B(n3316), .Z(n3348) );
  AND U4455 ( .A(y[1793]), .B(x[251]), .Z(n3326) );
  XOR U4456 ( .A(o[28]), .B(n3326), .Z(n3335) );
  AND U4457 ( .A(x[250]), .B(y[1794]), .Z(n3336) );
  XOR U4458 ( .A(n3335), .B(n3336), .Z(n3338) );
  AND U4459 ( .A(x[239]), .B(y[1805]), .Z(n3337) );
  XNOR U4460 ( .A(n3338), .B(n3337), .Z(n3347) );
  XOR U4461 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4462 ( .A(n3350), .B(n3349), .Z(n3377) );
  NAND U4463 ( .A(n3146), .B(n3145), .Z(n3150) );
  NAND U4464 ( .A(n3148), .B(n3147), .Z(n3149) );
  NAND U4465 ( .A(n3150), .B(n3149), .Z(n3356) );
  AND U4466 ( .A(x[241]), .B(y[1803]), .Z(n3279) );
  AND U4467 ( .A(x[246]), .B(y[1798]), .Z(n3280) );
  XOR U4468 ( .A(n3279), .B(n3280), .Z(n3281) );
  AND U4469 ( .A(x[228]), .B(y[1816]), .Z(n3282) );
  XOR U4470 ( .A(n3281), .B(n3282), .Z(n3354) );
  AND U4471 ( .A(x[230]), .B(y[1814]), .Z(n3535) );
  AND U4472 ( .A(y[1801]), .B(x[243]), .Z(n3327) );
  XOR U4473 ( .A(n3535), .B(n3327), .Z(n3328) );
  XOR U4474 ( .A(n3354), .B(n3353), .Z(n3355) );
  XOR U4475 ( .A(n3356), .B(n3355), .Z(n3378) );
  XOR U4476 ( .A(n3377), .B(n3378), .Z(n3380) );
  NAND U4477 ( .A(n3341), .B(n3151), .Z(n3155) );
  NAND U4478 ( .A(n3153), .B(n3152), .Z(n3154) );
  NAND U4479 ( .A(n3155), .B(n3154), .Z(n3276) );
  NAND U4480 ( .A(n3157), .B(n3156), .Z(n3161) );
  NAND U4481 ( .A(n3159), .B(n3158), .Z(n3160) );
  NAND U4482 ( .A(n3161), .B(n3160), .Z(n3274) );
  NAND U4483 ( .A(n3163), .B(n3162), .Z(n3167) );
  NAND U4484 ( .A(n3165), .B(n3164), .Z(n3166) );
  NAND U4485 ( .A(n3167), .B(n3166), .Z(n3273) );
  XOR U4486 ( .A(n3274), .B(n3273), .Z(n3275) );
  XOR U4487 ( .A(n3276), .B(n3275), .Z(n3379) );
  XOR U4488 ( .A(n3380), .B(n3379), .Z(n3269) );
  XOR U4489 ( .A(n3270), .B(n3269), .Z(n3264) );
  XOR U4490 ( .A(n3360), .B(n3359), .Z(n3361) );
  XNOR U4491 ( .A(n3362), .B(n3361), .Z(n3262) );
  AND U4492 ( .A(y[1799]), .B(x[248]), .Z(n3659) );
  NAND U4493 ( .A(n3659), .B(n3180), .Z(n3184) );
  NANDN U4494 ( .A(n3182), .B(n3181), .Z(n3183) );
  NAND U4495 ( .A(n3184), .B(n3183), .Z(n3398) );
  AND U4496 ( .A(x[249]), .B(y[1795]), .Z(n3310) );
  XOR U4497 ( .A(n3311), .B(n3310), .Z(n3309) );
  AND U4498 ( .A(x[225]), .B(y[1819]), .Z(n3308) );
  XOR U4499 ( .A(n3309), .B(n3308), .Z(n3396) );
  AND U4500 ( .A(y[1804]), .B(x[240]), .Z(n3302) );
  AND U4501 ( .A(x[248]), .B(y[1796]), .Z(n3303) );
  XOR U4502 ( .A(n3302), .B(n3303), .Z(n3304) );
  AND U4503 ( .A(x[226]), .B(y[1818]), .Z(n3305) );
  XOR U4504 ( .A(n3304), .B(n3305), .Z(n3395) );
  XOR U4505 ( .A(n3396), .B(n3395), .Z(n3397) );
  XNOR U4506 ( .A(n3398), .B(n3397), .Z(n3367) );
  NANDN U4507 ( .A(n3186), .B(n3185), .Z(n3190) );
  NANDN U4508 ( .A(n3188), .B(n3187), .Z(n3189) );
  NAND U4509 ( .A(n3190), .B(n3189), .Z(n3392) );
  AND U4510 ( .A(y[1817]), .B(x[227]), .Z(n3342) );
  XOR U4511 ( .A(n3341), .B(n3342), .Z(n3343) );
  AND U4512 ( .A(x[247]), .B(y[1797]), .Z(n3344) );
  XOR U4513 ( .A(n3343), .B(n3344), .Z(n3390) );
  AND U4514 ( .A(y[1815]), .B(x[229]), .Z(n3320) );
  AND U4515 ( .A(y[1799]), .B(x[245]), .Z(n3321) );
  XOR U4516 ( .A(n3320), .B(n3321), .Z(n3322) );
  AND U4517 ( .A(y[1800]), .B(x[244]), .Z(n3323) );
  XOR U4518 ( .A(n3322), .B(n3323), .Z(n3389) );
  XOR U4519 ( .A(n3390), .B(n3389), .Z(n3391) );
  XNOR U4520 ( .A(n3392), .B(n3391), .Z(n3366) );
  NANDN U4521 ( .A(n3192), .B(n3191), .Z(n3196) );
  NANDN U4522 ( .A(n3194), .B(n3193), .Z(n3195) );
  NAND U4523 ( .A(n3196), .B(n3195), .Z(n3299) );
  AND U4524 ( .A(x[224]), .B(y[1820]), .Z(n3286) );
  AND U4525 ( .A(x[252]), .B(y[1792]), .Z(n3285) );
  XOR U4526 ( .A(n3286), .B(n3285), .Z(n3288) );
  ANDN U4527 ( .B(o[27]), .A(n3197), .Z(n3287) );
  XOR U4528 ( .A(n3288), .B(n3287), .Z(n3297) );
  NAND U4529 ( .A(y[1810]), .B(x[234]), .Z(n3198) );
  XNOR U4530 ( .A(n3199), .B(n3198), .Z(n3293) );
  AND U4531 ( .A(x[233]), .B(y[1811]), .Z(n3292) );
  XOR U4532 ( .A(n3293), .B(n3292), .Z(n3296) );
  XOR U4533 ( .A(n3297), .B(n3296), .Z(n3298) );
  XOR U4534 ( .A(n3299), .B(n3298), .Z(n3386) );
  NANDN U4535 ( .A(n3201), .B(n3200), .Z(n3205) );
  NAND U4536 ( .A(n3203), .B(n3202), .Z(n3204) );
  NAND U4537 ( .A(n3205), .B(n3204), .Z(n3384) );
  NANDN U4538 ( .A(n3207), .B(n3206), .Z(n3211) );
  NANDN U4539 ( .A(n3209), .B(n3208), .Z(n3210) );
  NAND U4540 ( .A(n3211), .B(n3210), .Z(n3383) );
  XOR U4541 ( .A(n3384), .B(n3383), .Z(n3385) );
  XNOR U4542 ( .A(n3386), .B(n3385), .Z(n3365) );
  XOR U4543 ( .A(n3366), .B(n3365), .Z(n3368) );
  XOR U4544 ( .A(n3367), .B(n3368), .Z(n3261) );
  XOR U4545 ( .A(n3262), .B(n3261), .Z(n3263) );
  XOR U4546 ( .A(n3264), .B(n3263), .Z(n3257) );
  NANDN U4547 ( .A(n3213), .B(n3212), .Z(n3217) );
  OR U4548 ( .A(n3215), .B(n3214), .Z(n3216) );
  AND U4549 ( .A(n3217), .B(n3216), .Z(n3256) );
  NANDN U4550 ( .A(n3219), .B(n3218), .Z(n3223) );
  NANDN U4551 ( .A(n3221), .B(n3220), .Z(n3222) );
  NAND U4552 ( .A(n3223), .B(n3222), .Z(n3255) );
  XOR U4553 ( .A(n3256), .B(n3255), .Z(n3258) );
  XOR U4554 ( .A(n3257), .B(n3258), .Z(n3244) );
  NAND U4555 ( .A(n3225), .B(n3224), .Z(n3229) );
  NAND U4556 ( .A(n3227), .B(n3226), .Z(n3228) );
  NAND U4557 ( .A(n3229), .B(n3228), .Z(n3251) );
  NAND U4558 ( .A(n3231), .B(n3230), .Z(n3235) );
  NAND U4559 ( .A(n3233), .B(n3232), .Z(n3234) );
  NAND U4560 ( .A(n3235), .B(n3234), .Z(n3249) );
  NAND U4561 ( .A(n3237), .B(n3236), .Z(n3241) );
  NAND U4562 ( .A(n3239), .B(n3238), .Z(n3240) );
  AND U4563 ( .A(n3241), .B(n3240), .Z(n3250) );
  XNOR U4564 ( .A(n3249), .B(n3250), .Z(n3252) );
  XNOR U4565 ( .A(n3245), .B(n3246), .Z(n3403) );
  XOR U4566 ( .A(n3404), .B(n3403), .Z(n3410) );
  XNOR U4567 ( .A(n3408), .B(n3410), .Z(n3242) );
  XOR U4568 ( .A(n3407), .B(n3242), .Z(N61) );
  NANDN U4569 ( .A(n3244), .B(n3243), .Z(n3248) );
  NANDN U4570 ( .A(n3246), .B(n3245), .Z(n3247) );
  NAND U4571 ( .A(n3248), .B(n3247), .Z(n3583) );
  NAND U4572 ( .A(n3250), .B(n3249), .Z(n3254) );
  NANDN U4573 ( .A(n3252), .B(n3251), .Z(n3253) );
  NAND U4574 ( .A(n3254), .B(n3253), .Z(n3581) );
  NANDN U4575 ( .A(n3256), .B(n3255), .Z(n3260) );
  NANDN U4576 ( .A(n3258), .B(n3257), .Z(n3259) );
  AND U4577 ( .A(n3260), .B(n3259), .Z(n3416) );
  NAND U4578 ( .A(n3262), .B(n3261), .Z(n3266) );
  NANDN U4579 ( .A(n3264), .B(n3263), .Z(n3265) );
  AND U4580 ( .A(n3266), .B(n3265), .Z(n3415) );
  XNOR U4581 ( .A(n3416), .B(n3415), .Z(n3418) );
  NAND U4582 ( .A(n3268), .B(n3267), .Z(n3272) );
  NAND U4583 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U4584 ( .A(n3272), .B(n3271), .Z(n3567) );
  NAND U4585 ( .A(n3274), .B(n3273), .Z(n3278) );
  NAND U4586 ( .A(n3276), .B(n3275), .Z(n3277) );
  AND U4587 ( .A(n3278), .B(n3277), .Z(n3424) );
  NAND U4588 ( .A(n3280), .B(n3279), .Z(n3284) );
  NAND U4589 ( .A(n3282), .B(n3281), .Z(n3283) );
  NAND U4590 ( .A(n3284), .B(n3283), .Z(n3458) );
  NAND U4591 ( .A(n3286), .B(n3285), .Z(n3290) );
  NAND U4592 ( .A(n3288), .B(n3287), .Z(n3289) );
  NAND U4593 ( .A(n3290), .B(n3289), .Z(n3457) );
  XOR U4594 ( .A(n3458), .B(n3457), .Z(n3460) );
  AND U4595 ( .A(y[1812]), .B(x[234]), .Z(n3455) );
  NAND U4596 ( .A(n3455), .B(n3291), .Z(n3295) );
  NAND U4597 ( .A(n3293), .B(n3292), .Z(n3294) );
  NAND U4598 ( .A(n3295), .B(n3294), .Z(n3429) );
  AND U4599 ( .A(x[236]), .B(y[1809]), .Z(n3780) );
  AND U4600 ( .A(y[1820]), .B(x[225]), .Z(n3511) );
  XOR U4601 ( .A(n3780), .B(n3511), .Z(n3513) );
  AND U4602 ( .A(x[246]), .B(y[1799]), .Z(n3512) );
  XOR U4603 ( .A(n3513), .B(n3512), .Z(n3428) );
  AND U4604 ( .A(x[239]), .B(y[1806]), .Z(n3516) );
  XOR U4605 ( .A(n3516), .B(n3774), .Z(n3518) );
  XOR U4606 ( .A(n3518), .B(n3517), .Z(n3427) );
  XOR U4607 ( .A(n3428), .B(n3427), .Z(n3430) );
  XOR U4608 ( .A(n3429), .B(n3430), .Z(n3459) );
  XNOR U4609 ( .A(n3460), .B(n3459), .Z(n3422) );
  NAND U4610 ( .A(n3297), .B(n3296), .Z(n3301) );
  NAND U4611 ( .A(n3299), .B(n3298), .Z(n3300) );
  AND U4612 ( .A(n3301), .B(n3300), .Z(n3421) );
  XOR U4613 ( .A(n3422), .B(n3421), .Z(n3423) );
  XNOR U4614 ( .A(n3424), .B(n3423), .Z(n3466) );
  NAND U4615 ( .A(n3303), .B(n3302), .Z(n3307) );
  NAND U4616 ( .A(n3305), .B(n3304), .Z(n3306) );
  NAND U4617 ( .A(n3307), .B(n3306), .Z(n3434) );
  AND U4618 ( .A(n3309), .B(n3308), .Z(n3313) );
  NAND U4619 ( .A(n3311), .B(n3310), .Z(n3312) );
  NANDN U4620 ( .A(n3313), .B(n3312), .Z(n3433) );
  XOR U4621 ( .A(n3434), .B(n3433), .Z(n3436) );
  NAND U4622 ( .A(n3315), .B(n3314), .Z(n3319) );
  NAND U4623 ( .A(n3317), .B(n3316), .Z(n3318) );
  NAND U4624 ( .A(n3319), .B(n3318), .Z(n3477) );
  AND U4625 ( .A(y[1798]), .B(x[247]), .Z(n3526) );
  AND U4626 ( .A(x[237]), .B(y[1808]), .Z(n3524) );
  AND U4627 ( .A(x[248]), .B(y[1797]), .Z(n3744) );
  XOR U4628 ( .A(n3524), .B(n3744), .Z(n3525) );
  XOR U4629 ( .A(n3526), .B(n3525), .Z(n3476) );
  AND U4630 ( .A(y[1810]), .B(x[235]), .Z(n3532) );
  AND U4631 ( .A(x[227]), .B(y[1818]), .Z(n3530) );
  AND U4632 ( .A(x[241]), .B(y[1804]), .Z(n3529) );
  XOR U4633 ( .A(n3530), .B(n3529), .Z(n3531) );
  XOR U4634 ( .A(n3532), .B(n3531), .Z(n3475) );
  XOR U4635 ( .A(n3476), .B(n3475), .Z(n3478) );
  XOR U4636 ( .A(n3477), .B(n3478), .Z(n3435) );
  XOR U4637 ( .A(n3436), .B(n3435), .Z(n3557) );
  NAND U4638 ( .A(n3321), .B(n3320), .Z(n3325) );
  NAND U4639 ( .A(n3323), .B(n3322), .Z(n3324) );
  NAND U4640 ( .A(n3325), .B(n3324), .Z(n3544) );
  AND U4641 ( .A(x[226]), .B(y[1819]), .Z(n3494) );
  XOR U4642 ( .A(n3494), .B(n3493), .Z(n3496) );
  XOR U4643 ( .A(n3496), .B(n3495), .Z(n3543) );
  AND U4644 ( .A(y[1805]), .B(x[240]), .Z(n3482) );
  AND U4645 ( .A(x[251]), .B(y[1794]), .Z(n3481) );
  XOR U4646 ( .A(n3482), .B(n3481), .Z(n3484) );
  AND U4647 ( .A(o[28]), .B(n3326), .Z(n3483) );
  XOR U4648 ( .A(n3484), .B(n3483), .Z(n3542) );
  XOR U4649 ( .A(n3543), .B(n3542), .Z(n3545) );
  XOR U4650 ( .A(n3544), .B(n3545), .Z(n3555) );
  NAND U4651 ( .A(n3327), .B(n3535), .Z(n3331) );
  NANDN U4652 ( .A(n3329), .B(n3328), .Z(n3330) );
  AND U4653 ( .A(n3331), .B(n3330), .Z(n3442) );
  AND U4654 ( .A(x[250]), .B(y[1795]), .Z(n3505) );
  XOR U4655 ( .A(n3506), .B(n3505), .Z(n3508) );
  AND U4656 ( .A(x[249]), .B(y[1796]), .Z(n3507) );
  XNOR U4657 ( .A(n3508), .B(n3507), .Z(n3440) );
  AND U4658 ( .A(x[252]), .B(y[1793]), .Z(n3523) );
  XOR U4659 ( .A(o[29]), .B(n3523), .Z(n3450) );
  AND U4660 ( .A(x[224]), .B(y[1821]), .Z(n3448) );
  AND U4661 ( .A(y[1792]), .B(x[253]), .Z(n3447) );
  XOR U4662 ( .A(n3448), .B(n3447), .Z(n3449) );
  XNOR U4663 ( .A(n3450), .B(n3449), .Z(n3439) );
  XOR U4664 ( .A(n3440), .B(n3439), .Z(n3441) );
  XOR U4665 ( .A(n3442), .B(n3441), .Z(n3554) );
  AND U4666 ( .A(x[228]), .B(y[1817]), .Z(n3488) );
  AND U4667 ( .A(x[234]), .B(y[1811]), .Z(n3487) );
  XOR U4668 ( .A(n3488), .B(n3487), .Z(n3490) );
  AND U4669 ( .A(y[1816]), .B(x[229]), .Z(n3489) );
  XNOR U4670 ( .A(n3490), .B(n3489), .Z(n3446) );
  NAND U4671 ( .A(y[1812]), .B(x[233]), .Z(n3700) );
  AND U4672 ( .A(y[1815]), .B(x[230]), .Z(n3333) );
  NAND U4673 ( .A(y[1814]), .B(x[231]), .Z(n3332) );
  XNOR U4674 ( .A(n3333), .B(n3332), .Z(n3537) );
  AND U4675 ( .A(x[232]), .B(y[1813]), .Z(n3536) );
  XNOR U4676 ( .A(n3537), .B(n3536), .Z(n3445) );
  XOR U4677 ( .A(n3700), .B(n3445), .Z(n3334) );
  XNOR U4678 ( .A(n3446), .B(n3334), .Z(n3501) );
  NAND U4679 ( .A(n3336), .B(n3335), .Z(n3340) );
  NAND U4680 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U4681 ( .A(n3340), .B(n3339), .Z(n3500) );
  NAND U4682 ( .A(n3342), .B(n3341), .Z(n3346) );
  NAND U4683 ( .A(n3344), .B(n3343), .Z(n3345) );
  NAND U4684 ( .A(n3346), .B(n3345), .Z(n3499) );
  XNOR U4685 ( .A(n3500), .B(n3499), .Z(n3502) );
  NAND U4686 ( .A(n3348), .B(n3347), .Z(n3352) );
  NAND U4687 ( .A(n3350), .B(n3349), .Z(n3351) );
  NAND U4688 ( .A(n3352), .B(n3351), .Z(n3469) );
  XNOR U4689 ( .A(n3472), .B(n3471), .Z(n3464) );
  NAND U4690 ( .A(n3354), .B(n3353), .Z(n3358) );
  NAND U4691 ( .A(n3356), .B(n3355), .Z(n3357) );
  NAND U4692 ( .A(n3358), .B(n3357), .Z(n3463) );
  XOR U4693 ( .A(n3464), .B(n3463), .Z(n3465) );
  XOR U4694 ( .A(n3466), .B(n3465), .Z(n3566) );
  XOR U4695 ( .A(n3567), .B(n3566), .Z(n3569) );
  NAND U4696 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U4697 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U4698 ( .A(n3364), .B(n3363), .Z(n3561) );
  NAND U4699 ( .A(n3366), .B(n3365), .Z(n3370) );
  NAND U4700 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U4701 ( .A(n3370), .B(n3369), .Z(n3560) );
  XOR U4702 ( .A(n3561), .B(n3560), .Z(n3563) );
  NAND U4703 ( .A(n3372), .B(n3371), .Z(n3376) );
  NAND U4704 ( .A(n3374), .B(n3373), .Z(n3375) );
  NAND U4705 ( .A(n3376), .B(n3375), .Z(n3574) );
  NAND U4706 ( .A(n3378), .B(n3377), .Z(n3382) );
  NAND U4707 ( .A(n3380), .B(n3379), .Z(n3381) );
  NAND U4708 ( .A(n3382), .B(n3381), .Z(n3572) );
  NAND U4709 ( .A(n3384), .B(n3383), .Z(n3388) );
  NAND U4710 ( .A(n3386), .B(n3385), .Z(n3387) );
  NAND U4711 ( .A(n3388), .B(n3387), .Z(n3551) );
  NAND U4712 ( .A(n3390), .B(n3389), .Z(n3394) );
  NAND U4713 ( .A(n3392), .B(n3391), .Z(n3393) );
  NAND U4714 ( .A(n3394), .B(n3393), .Z(n3549) );
  NAND U4715 ( .A(n3396), .B(n3395), .Z(n3400) );
  NAND U4716 ( .A(n3398), .B(n3397), .Z(n3399) );
  NAND U4717 ( .A(n3400), .B(n3399), .Z(n3548) );
  XOR U4718 ( .A(n3549), .B(n3548), .Z(n3550) );
  XOR U4719 ( .A(n3551), .B(n3550), .Z(n3573) );
  XOR U4720 ( .A(n3572), .B(n3573), .Z(n3575) );
  XOR U4721 ( .A(n3574), .B(n3575), .Z(n3562) );
  XOR U4722 ( .A(n3563), .B(n3562), .Z(n3568) );
  XOR U4723 ( .A(n3569), .B(n3568), .Z(n3417) );
  XOR U4724 ( .A(n3418), .B(n3417), .Z(n3582) );
  XNOR U4725 ( .A(n3581), .B(n3582), .Z(n3584) );
  XOR U4726 ( .A(n3583), .B(n3584), .Z(n3580) );
  NAND U4727 ( .A(n3402), .B(n3401), .Z(n3406) );
  NAND U4728 ( .A(n3404), .B(n3403), .Z(n3405) );
  NAND U4729 ( .A(n3406), .B(n3405), .Z(n3579) );
  NANDN U4730 ( .A(n3407), .B(n3408), .Z(n3413) );
  NOR U4731 ( .A(n3409), .B(n3408), .Z(n3411) );
  OR U4732 ( .A(n3411), .B(n3410), .Z(n3412) );
  AND U4733 ( .A(n3413), .B(n3412), .Z(n3578) );
  XOR U4734 ( .A(n3579), .B(n3578), .Z(n3414) );
  XNOR U4735 ( .A(n3580), .B(n3414), .Z(N62) );
  NANDN U4736 ( .A(n3416), .B(n3415), .Z(n3420) );
  NAND U4737 ( .A(n3418), .B(n3417), .Z(n3419) );
  AND U4738 ( .A(n3420), .B(n3419), .Z(n3588) );
  NAND U4739 ( .A(n3422), .B(n3421), .Z(n3426) );
  NAND U4740 ( .A(n3424), .B(n3423), .Z(n3425) );
  AND U4741 ( .A(n3426), .B(n3425), .Z(n3837) );
  NAND U4742 ( .A(n3428), .B(n3427), .Z(n3432) );
  NAND U4743 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U4744 ( .A(n3432), .B(n3431), .Z(n3822) );
  NAND U4745 ( .A(n3434), .B(n3433), .Z(n3438) );
  NAND U4746 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U4747 ( .A(n3438), .B(n3437), .Z(n3821) );
  XOR U4748 ( .A(n3822), .B(n3821), .Z(n3820) );
  NAND U4749 ( .A(n3440), .B(n3439), .Z(n3444) );
  NAND U4750 ( .A(n3442), .B(n3441), .Z(n3443) );
  NAND U4751 ( .A(n3444), .B(n3443), .Z(n3819) );
  XOR U4752 ( .A(n3820), .B(n3819), .Z(n3840) );
  NAND U4753 ( .A(n3448), .B(n3447), .Z(n3452) );
  NAND U4754 ( .A(n3450), .B(n3449), .Z(n3451) );
  NAND U4755 ( .A(n3452), .B(n3451), .Z(n3627) );
  NAND U4756 ( .A(x[236]), .B(y[1810]), .Z(n3453) );
  XNOR U4757 ( .A(n3454), .B(n3453), .Z(n3782) );
  XOR U4758 ( .A(n3782), .B(n3781), .Z(n3698) );
  AND U4759 ( .A(y[1813]), .B(x[233]), .Z(n3456) );
  XOR U4760 ( .A(n3456), .B(n3455), .Z(n3697) );
  XOR U4761 ( .A(n3698), .B(n3697), .Z(n3630) );
  AND U4762 ( .A(y[1795]), .B(x[251]), .Z(n3764) );
  AND U4763 ( .A(x[225]), .B(y[1821]), .Z(n3763) );
  XOR U4764 ( .A(n3764), .B(n3763), .Z(n3762) );
  XOR U4765 ( .A(n3762), .B(n3761), .Z(n3629) );
  XOR U4766 ( .A(n3630), .B(n3629), .Z(n3628) );
  XOR U4767 ( .A(n3627), .B(n3628), .Z(n3816) );
  NAND U4768 ( .A(n3458), .B(n3457), .Z(n3462) );
  NAND U4769 ( .A(n3460), .B(n3459), .Z(n3461) );
  AND U4770 ( .A(n3462), .B(n3461), .Z(n3813) );
  XNOR U4771 ( .A(n3814), .B(n3813), .Z(n3839) );
  XNOR U4772 ( .A(n3837), .B(n3838), .Z(n3868) );
  NAND U4773 ( .A(n3464), .B(n3463), .Z(n3468) );
  NAND U4774 ( .A(n3466), .B(n3465), .Z(n3467) );
  AND U4775 ( .A(n3468), .B(n3467), .Z(n3870) );
  NANDN U4776 ( .A(n3470), .B(n3469), .Z(n3474) );
  NAND U4777 ( .A(n3472), .B(n3471), .Z(n3473) );
  AND U4778 ( .A(n3474), .B(n3473), .Z(n3855) );
  NAND U4779 ( .A(n3476), .B(n3475), .Z(n3480) );
  NAND U4780 ( .A(n3478), .B(n3477), .Z(n3479) );
  AND U4781 ( .A(n3480), .B(n3479), .Z(n3833) );
  NAND U4782 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U4783 ( .A(n3484), .B(n3483), .Z(n3485) );
  NAND U4784 ( .A(n3486), .B(n3485), .Z(n3797) );
  NAND U4785 ( .A(n3488), .B(n3487), .Z(n3492) );
  NAND U4786 ( .A(n3490), .B(n3489), .Z(n3491) );
  NAND U4787 ( .A(n3492), .B(n3491), .Z(n3800) );
  AND U4788 ( .A(y[1816]), .B(x[230]), .Z(n3756) );
  AND U4789 ( .A(y[1817]), .B(x[229]), .Z(n3758) );
  AND U4790 ( .A(y[1803]), .B(x[243]), .Z(n3757) );
  XOR U4791 ( .A(n3758), .B(n3757), .Z(n3755) );
  XNOR U4792 ( .A(n3756), .B(n3755), .Z(n3633) );
  AND U4793 ( .A(x[228]), .B(y[1818]), .Z(n3748) );
  AND U4794 ( .A(x[227]), .B(y[1819]), .Z(n3750) );
  AND U4795 ( .A(x[242]), .B(y[1804]), .Z(n3749) );
  XOR U4796 ( .A(n3750), .B(n3749), .Z(n3747) );
  XOR U4797 ( .A(n3748), .B(n3747), .Z(n3636) );
  NAND U4798 ( .A(n3494), .B(n3493), .Z(n3498) );
  NAND U4799 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U4800 ( .A(n3498), .B(n3497), .Z(n3635) );
  XOR U4801 ( .A(n3633), .B(n3634), .Z(n3799) );
  XOR U4802 ( .A(n3800), .B(n3799), .Z(n3798) );
  XOR U4803 ( .A(n3797), .B(n3798), .Z(n3834) );
  NAND U4804 ( .A(n3500), .B(n3499), .Z(n3504) );
  NANDN U4805 ( .A(n3502), .B(n3501), .Z(n3503) );
  AND U4806 ( .A(n3504), .B(n3503), .Z(n3831) );
  XOR U4807 ( .A(n3832), .B(n3831), .Z(n3858) );
  AND U4808 ( .A(n3506), .B(n3505), .Z(n3510) );
  NAND U4809 ( .A(n3508), .B(n3507), .Z(n3509) );
  NANDN U4810 ( .A(n3510), .B(n3509), .Z(n3791) );
  AND U4811 ( .A(n3780), .B(n3511), .Z(n3515) );
  NAND U4812 ( .A(n3513), .B(n3512), .Z(n3514) );
  NANDN U4813 ( .A(n3515), .B(n3514), .Z(n3794) );
  NAND U4814 ( .A(n3516), .B(n3774), .Z(n3520) );
  NAND U4815 ( .A(n3518), .B(n3517), .Z(n3519) );
  AND U4816 ( .A(n3520), .B(n3519), .Z(n3608) );
  AND U4817 ( .A(y[1799]), .B(x[247]), .Z(n3742) );
  AND U4818 ( .A(y[1797]), .B(x[249]), .Z(n3522) );
  AND U4819 ( .A(x[248]), .B(y[1798]), .Z(n3521) );
  XOR U4820 ( .A(n3522), .B(n3521), .Z(n3741) );
  XOR U4821 ( .A(n3742), .B(n3741), .Z(n3610) );
  AND U4822 ( .A(n3523), .B(o[29]), .Z(n3722) );
  AND U4823 ( .A(x[252]), .B(y[1794]), .Z(n3724) );
  AND U4824 ( .A(y[1806]), .B(x[240]), .Z(n3723) );
  XOR U4825 ( .A(n3724), .B(n3723), .Z(n3721) );
  XNOR U4826 ( .A(n3722), .B(n3721), .Z(n3609) );
  XNOR U4827 ( .A(n3608), .B(n3607), .Z(n3793) );
  XOR U4828 ( .A(n3794), .B(n3793), .Z(n3792) );
  XOR U4829 ( .A(n3791), .B(n3792), .Z(n3596) );
  NAND U4830 ( .A(n3524), .B(n3744), .Z(n3528) );
  NAND U4831 ( .A(n3526), .B(n3525), .Z(n3527) );
  NAND U4832 ( .A(n3528), .B(n3527), .Z(n3604) );
  NAND U4833 ( .A(n3530), .B(n3529), .Z(n3534) );
  NAND U4834 ( .A(n3532), .B(n3531), .Z(n3533) );
  AND U4835 ( .A(n3534), .B(n3533), .Z(n3620) );
  AND U4836 ( .A(x[224]), .B(y[1822]), .Z(n3692) );
  AND U4837 ( .A(y[1793]), .B(x[253]), .Z(n3678) );
  XOR U4838 ( .A(o[30]), .B(n3678), .Z(n3694) );
  AND U4839 ( .A(y[1792]), .B(x[254]), .Z(n3693) );
  XOR U4840 ( .A(n3694), .B(n3693), .Z(n3691) );
  XOR U4841 ( .A(n3692), .B(n3691), .Z(n3622) );
  AND U4842 ( .A(x[244]), .B(y[1802]), .Z(n3648) );
  XOR U4843 ( .A(n3648), .B(n3647), .Z(n3646) );
  AND U4844 ( .A(x[232]), .B(y[1814]), .Z(n3645) );
  XNOR U4845 ( .A(n3646), .B(n3645), .Z(n3621) );
  XNOR U4846 ( .A(n3620), .B(n3619), .Z(n3603) );
  XOR U4847 ( .A(n3604), .B(n3603), .Z(n3601) );
  AND U4848 ( .A(x[231]), .B(y[1815]), .Z(n3776) );
  NAND U4849 ( .A(n3535), .B(n3776), .Z(n3539) );
  NAND U4850 ( .A(n3537), .B(n3536), .Z(n3538) );
  AND U4851 ( .A(n3539), .B(n3538), .Z(n3613) );
  AND U4852 ( .A(y[1801]), .B(x[245]), .Z(n3541) );
  AND U4853 ( .A(y[1800]), .B(x[246]), .Z(n3540) );
  XOR U4854 ( .A(n3541), .B(n3540), .Z(n3775) );
  XOR U4855 ( .A(n3776), .B(n3775), .Z(n3616) );
  AND U4856 ( .A(x[241]), .B(y[1805]), .Z(n3640) );
  AND U4857 ( .A(y[1820]), .B(x[226]), .Z(n3642) );
  AND U4858 ( .A(x[250]), .B(y[1796]), .Z(n3641) );
  XOR U4859 ( .A(n3642), .B(n3641), .Z(n3639) );
  XNOR U4860 ( .A(n3640), .B(n3639), .Z(n3615) );
  XNOR U4861 ( .A(n3613), .B(n3614), .Z(n3602) );
  NAND U4862 ( .A(n3543), .B(n3542), .Z(n3547) );
  NAND U4863 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U4864 ( .A(n3547), .B(n3546), .Z(n3597) );
  XOR U4865 ( .A(n3598), .B(n3597), .Z(n3595) );
  XOR U4866 ( .A(n3596), .B(n3595), .Z(n3857) );
  XNOR U4867 ( .A(n3855), .B(n3856), .Z(n3594) );
  NAND U4868 ( .A(n3549), .B(n3548), .Z(n3553) );
  NAND U4869 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U4870 ( .A(n3553), .B(n3552), .Z(n3593) );
  NANDN U4871 ( .A(n3555), .B(n3554), .Z(n3559) );
  NANDN U4872 ( .A(n3557), .B(n3556), .Z(n3558) );
  NAND U4873 ( .A(n3559), .B(n3558), .Z(n3591) );
  XOR U4874 ( .A(n3592), .B(n3591), .Z(n3869) );
  XOR U4875 ( .A(n3870), .B(n3869), .Z(n3867) );
  NAND U4876 ( .A(n3561), .B(n3560), .Z(n3565) );
  NAND U4877 ( .A(n3563), .B(n3562), .Z(n3564) );
  AND U4878 ( .A(n3565), .B(n3564), .Z(n3852) );
  NAND U4879 ( .A(n3567), .B(n3566), .Z(n3571) );
  NAND U4880 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U4881 ( .A(n3571), .B(n3570), .Z(n3851) );
  XOR U4882 ( .A(n3852), .B(n3851), .Z(n3850) );
  NAND U4883 ( .A(n3573), .B(n3572), .Z(n3577) );
  NAND U4884 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U4885 ( .A(n3577), .B(n3576), .Z(n3849) );
  XOR U4886 ( .A(n3850), .B(n3849), .Z(n3589) );
  XOR U4887 ( .A(n3590), .B(n3589), .Z(n3587) );
  XOR U4888 ( .A(n3588), .B(n3587), .Z(n3864) );
  NAND U4889 ( .A(n3582), .B(n3581), .Z(n3586) );
  NANDN U4890 ( .A(n3584), .B(n3583), .Z(n3585) );
  NAND U4891 ( .A(n3586), .B(n3585), .Z(n3866) );
  XNOR U4892 ( .A(n3864), .B(n3863), .Z(N63) );
  NAND U4893 ( .A(n3596), .B(n3595), .Z(n3600) );
  NAND U4894 ( .A(n3598), .B(n3597), .Z(n3599) );
  AND U4895 ( .A(n3600), .B(n3599), .Z(n3848) );
  NANDN U4896 ( .A(n3602), .B(n3601), .Z(n3606) );
  NAND U4897 ( .A(n3604), .B(n3603), .Z(n3605) );
  AND U4898 ( .A(n3606), .B(n3605), .Z(n3830) );
  NAND U4899 ( .A(n3608), .B(n3607), .Z(n3612) );
  NANDN U4900 ( .A(n3610), .B(n3609), .Z(n3611) );
  AND U4901 ( .A(n3612), .B(n3611), .Z(n3812) );
  NANDN U4902 ( .A(n3614), .B(n3613), .Z(n3618) );
  NANDN U4903 ( .A(n3616), .B(n3615), .Z(n3617) );
  AND U4904 ( .A(n3618), .B(n3617), .Z(n3626) );
  NAND U4905 ( .A(n3620), .B(n3619), .Z(n3624) );
  NANDN U4906 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U4907 ( .A(n3624), .B(n3623), .Z(n3625) );
  XNOR U4908 ( .A(n3626), .B(n3625), .Z(n3810) );
  NAND U4909 ( .A(n3628), .B(n3627), .Z(n3632) );
  NAND U4910 ( .A(n3630), .B(n3629), .Z(n3631) );
  AND U4911 ( .A(n3632), .B(n3631), .Z(n3808) );
  NANDN U4912 ( .A(n3634), .B(n3633), .Z(n3638) );
  NANDN U4913 ( .A(n3636), .B(n3635), .Z(n3637) );
  AND U4914 ( .A(n3638), .B(n3637), .Z(n3718) );
  NAND U4915 ( .A(n3640), .B(n3639), .Z(n3644) );
  NAND U4916 ( .A(n3642), .B(n3641), .Z(n3643) );
  AND U4917 ( .A(n3644), .B(n3643), .Z(n3652) );
  NAND U4918 ( .A(n3646), .B(n3645), .Z(n3650) );
  NAND U4919 ( .A(n3648), .B(n3647), .Z(n3649) );
  NAND U4920 ( .A(n3650), .B(n3649), .Z(n3651) );
  XNOR U4921 ( .A(n3652), .B(n3651), .Z(n3716) );
  AND U4922 ( .A(x[229]), .B(y[1818]), .Z(n3654) );
  NAND U4923 ( .A(x[231]), .B(y[1816]), .Z(n3653) );
  XNOR U4924 ( .A(n3654), .B(n3653), .Z(n3658) );
  AND U4925 ( .A(y[1805]), .B(x[242]), .Z(n3656) );
  NAND U4926 ( .A(x[227]), .B(y[1820]), .Z(n3655) );
  XNOR U4927 ( .A(n3656), .B(n3655), .Z(n3657) );
  XOR U4928 ( .A(n3658), .B(n3657), .Z(n3661) );
  AND U4929 ( .A(x[246]), .B(y[1801]), .Z(n3773) );
  XNOR U4930 ( .A(n3773), .B(n3659), .Z(n3660) );
  XNOR U4931 ( .A(n3661), .B(n3660), .Z(n3677) );
  AND U4932 ( .A(y[1794]), .B(x[253]), .Z(n3663) );
  NAND U4933 ( .A(x[244]), .B(y[1803]), .Z(n3662) );
  XNOR U4934 ( .A(n3663), .B(n3662), .Z(n3667) );
  AND U4935 ( .A(x[238]), .B(y[1809]), .Z(n3665) );
  NAND U4936 ( .A(x[254]), .B(y[1793]), .Z(n3664) );
  XNOR U4937 ( .A(n3665), .B(n3664), .Z(n3666) );
  XOR U4938 ( .A(n3667), .B(n3666), .Z(n3675) );
  AND U4939 ( .A(x[255]), .B(y[1792]), .Z(n3669) );
  NAND U4940 ( .A(y[1819]), .B(x[228]), .Z(n3668) );
  XNOR U4941 ( .A(n3669), .B(n3668), .Z(n3673) );
  AND U4942 ( .A(x[240]), .B(y[1807]), .Z(n3671) );
  NAND U4943 ( .A(y[1806]), .B(x[241]), .Z(n3670) );
  XNOR U4944 ( .A(n3671), .B(n3670), .Z(n3672) );
  XNOR U4945 ( .A(n3673), .B(n3672), .Z(n3674) );
  XNOR U4946 ( .A(n3675), .B(n3674), .Z(n3676) );
  XOR U4947 ( .A(n3677), .B(n3676), .Z(n3690) );
  AND U4948 ( .A(y[1802]), .B(x[245]), .Z(n3684) );
  AND U4949 ( .A(n3678), .B(o[30]), .Z(n3682) );
  AND U4950 ( .A(y[1798]), .B(x[249]), .Z(n3743) );
  XOR U4951 ( .A(n3743), .B(o[31]), .Z(n3680) );
  AND U4952 ( .A(x[234]), .B(y[1813]), .Z(n3699) );
  XNOR U4953 ( .A(n3779), .B(n3699), .Z(n3679) );
  XNOR U4954 ( .A(n3680), .B(n3679), .Z(n3681) );
  XNOR U4955 ( .A(n3682), .B(n3681), .Z(n3683) );
  XNOR U4956 ( .A(n3684), .B(n3683), .Z(n3688) );
  AND U4957 ( .A(x[230]), .B(y[1817]), .Z(n3686) );
  NAND U4958 ( .A(x[243]), .B(y[1804]), .Z(n3685) );
  XNOR U4959 ( .A(n3686), .B(n3685), .Z(n3687) );
  XNOR U4960 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U4961 ( .A(n3690), .B(n3689), .Z(n3706) );
  NAND U4962 ( .A(n3692), .B(n3691), .Z(n3696) );
  NAND U4963 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U4964 ( .A(n3696), .B(n3695), .Z(n3704) );
  NAND U4965 ( .A(n3698), .B(n3697), .Z(n3702) );
  NANDN U4966 ( .A(n3700), .B(n3699), .Z(n3701) );
  NAND U4967 ( .A(n3702), .B(n3701), .Z(n3703) );
  XNOR U4968 ( .A(n3704), .B(n3703), .Z(n3705) );
  XOR U4969 ( .A(n3706), .B(n3705), .Z(n3714) );
  AND U4970 ( .A(x[247]), .B(y[1800]), .Z(n3708) );
  NAND U4971 ( .A(y[1815]), .B(x[232]), .Z(n3707) );
  XNOR U4972 ( .A(n3708), .B(n3707), .Z(n3712) );
  AND U4973 ( .A(x[251]), .B(y[1796]), .Z(n3710) );
  NAND U4974 ( .A(y[1821]), .B(x[226]), .Z(n3709) );
  XNOR U4975 ( .A(n3710), .B(n3709), .Z(n3711) );
  XNOR U4976 ( .A(n3712), .B(n3711), .Z(n3713) );
  XNOR U4977 ( .A(n3714), .B(n3713), .Z(n3715) );
  XNOR U4978 ( .A(n3716), .B(n3715), .Z(n3717) );
  XNOR U4979 ( .A(n3718), .B(n3717), .Z(n3790) );
  AND U4980 ( .A(x[236]), .B(y[1811]), .Z(n3720) );
  NAND U4981 ( .A(y[1795]), .B(x[252]), .Z(n3719) );
  XNOR U4982 ( .A(n3720), .B(n3719), .Z(n3740) );
  NAND U4983 ( .A(n3722), .B(n3721), .Z(n3726) );
  NAND U4984 ( .A(n3724), .B(n3723), .Z(n3725) );
  AND U4985 ( .A(n3726), .B(n3725), .Z(n3738) );
  AND U4986 ( .A(y[1822]), .B(x[225]), .Z(n3728) );
  NAND U4987 ( .A(y[1823]), .B(x[224]), .Z(n3727) );
  XNOR U4988 ( .A(n3728), .B(n3727), .Z(n3736) );
  AND U4989 ( .A(y[1797]), .B(x[250]), .Z(n3734) );
  AND U4990 ( .A(y[1814]), .B(x[233]), .Z(n3730) );
  NAND U4991 ( .A(x[235]), .B(y[1812]), .Z(n3729) );
  XNOR U4992 ( .A(n3730), .B(n3729), .Z(n3731) );
  XNOR U4993 ( .A(n3732), .B(n3731), .Z(n3733) );
  XNOR U4994 ( .A(n3734), .B(n3733), .Z(n3735) );
  XNOR U4995 ( .A(n3736), .B(n3735), .Z(n3737) );
  XNOR U4996 ( .A(n3738), .B(n3737), .Z(n3739) );
  XOR U4997 ( .A(n3740), .B(n3739), .Z(n3772) );
  NAND U4998 ( .A(n3742), .B(n3741), .Z(n3746) );
  NAND U4999 ( .A(n3744), .B(n3743), .Z(n3745) );
  AND U5000 ( .A(n3746), .B(n3745), .Z(n3754) );
  NAND U5001 ( .A(n3748), .B(n3747), .Z(n3752) );
  NAND U5002 ( .A(n3750), .B(n3749), .Z(n3751) );
  NAND U5003 ( .A(n3752), .B(n3751), .Z(n3753) );
  XNOR U5004 ( .A(n3754), .B(n3753), .Z(n3770) );
  NAND U5005 ( .A(n3756), .B(n3755), .Z(n3760) );
  NAND U5006 ( .A(n3758), .B(n3757), .Z(n3759) );
  AND U5007 ( .A(n3760), .B(n3759), .Z(n3768) );
  NAND U5008 ( .A(n3762), .B(n3761), .Z(n3766) );
  NAND U5009 ( .A(n3764), .B(n3763), .Z(n3765) );
  NAND U5010 ( .A(n3766), .B(n3765), .Z(n3767) );
  XNOR U5011 ( .A(n3768), .B(n3767), .Z(n3769) );
  XNOR U5012 ( .A(n3770), .B(n3769), .Z(n3771) );
  XNOR U5013 ( .A(n3772), .B(n3771), .Z(n3788) );
  AND U5014 ( .A(n3774), .B(n3773), .Z(n3778) );
  AND U5015 ( .A(n3776), .B(n3775), .Z(n3777) );
  NOR U5016 ( .A(n3778), .B(n3777), .Z(n3786) );
  NAND U5017 ( .A(n3780), .B(n3779), .Z(n3784) );
  NAND U5018 ( .A(n3782), .B(n3781), .Z(n3783) );
  AND U5019 ( .A(n3784), .B(n3783), .Z(n3785) );
  XNOR U5020 ( .A(n3786), .B(n3785), .Z(n3787) );
  XOR U5021 ( .A(n3788), .B(n3787), .Z(n3789) );
  XNOR U5022 ( .A(n3790), .B(n3789), .Z(n3806) );
  NAND U5023 ( .A(n3792), .B(n3791), .Z(n3796) );
  NAND U5024 ( .A(n3794), .B(n3793), .Z(n3795) );
  AND U5025 ( .A(n3796), .B(n3795), .Z(n3804) );
  NAND U5026 ( .A(n3798), .B(n3797), .Z(n3802) );
  NAND U5027 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U5028 ( .A(n3802), .B(n3801), .Z(n3803) );
  XNOR U5029 ( .A(n3804), .B(n3803), .Z(n3805) );
  XNOR U5030 ( .A(n3806), .B(n3805), .Z(n3807) );
  XNOR U5031 ( .A(n3808), .B(n3807), .Z(n3809) );
  XNOR U5032 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR U5033 ( .A(n3812), .B(n3811), .Z(n3828) );
  NAND U5034 ( .A(n3814), .B(n3813), .Z(n3818) );
  NANDN U5035 ( .A(n3816), .B(n3815), .Z(n3817) );
  AND U5036 ( .A(n3818), .B(n3817), .Z(n3826) );
  NAND U5037 ( .A(n3820), .B(n3819), .Z(n3824) );
  NAND U5038 ( .A(n3822), .B(n3821), .Z(n3823) );
  NAND U5039 ( .A(n3824), .B(n3823), .Z(n3825) );
  XNOR U5040 ( .A(n3826), .B(n3825), .Z(n3827) );
  XNOR U5041 ( .A(n3828), .B(n3827), .Z(n3829) );
  XNOR U5042 ( .A(n3830), .B(n3829), .Z(n3846) );
  NAND U5043 ( .A(n3832), .B(n3831), .Z(n3836) );
  NANDN U5044 ( .A(n3834), .B(n3833), .Z(n3835) );
  AND U5045 ( .A(n3836), .B(n3835), .Z(n3844) );
  NANDN U5046 ( .A(n3838), .B(n3837), .Z(n3842) );
  NANDN U5047 ( .A(n3840), .B(n3839), .Z(n3841) );
  NAND U5048 ( .A(n3842), .B(n3841), .Z(n3843) );
  XNOR U5049 ( .A(n3844), .B(n3843), .Z(n3845) );
  XNOR U5050 ( .A(n3846), .B(n3845), .Z(n3847) );
  NAND U5051 ( .A(n3850), .B(n3849), .Z(n3854) );
  NAND U5052 ( .A(n3852), .B(n3851), .Z(n3853) );
  AND U5053 ( .A(n3854), .B(n3853), .Z(n3862) );
  NANDN U5054 ( .A(n3856), .B(n3855), .Z(n3860) );
  NANDN U5055 ( .A(n3858), .B(n3857), .Z(n3859) );
  NAND U5056 ( .A(n3860), .B(n3859), .Z(n3861) );
  AND U5057 ( .A(x[224]), .B(y[1824]), .Z(n4520) );
  XOR U5058 ( .A(n4520), .B(o[32]), .Z(N97) );
  AND U5059 ( .A(x[225]), .B(y[1824]), .Z(n3879) );
  AND U5060 ( .A(x[224]), .B(y[1825]), .Z(n3878) );
  XNOR U5061 ( .A(n3878), .B(o[33]), .Z(n3871) );
  XNOR U5062 ( .A(n3879), .B(n3871), .Z(n3873) );
  NAND U5063 ( .A(n4520), .B(o[32]), .Z(n3872) );
  XNOR U5064 ( .A(n3873), .B(n3872), .Z(N98) );
  NANDN U5065 ( .A(n3879), .B(n3871), .Z(n3875) );
  NAND U5066 ( .A(n3873), .B(n3872), .Z(n3874) );
  AND U5067 ( .A(n3875), .B(n3874), .Z(n3885) );
  AND U5068 ( .A(x[224]), .B(y[1826]), .Z(n3892) );
  XNOR U5069 ( .A(n3892), .B(o[34]), .Z(n3884) );
  XNOR U5070 ( .A(n3885), .B(n3884), .Z(n3887) );
  AND U5071 ( .A(y[1824]), .B(x[226]), .Z(n3877) );
  NAND U5072 ( .A(y[1825]), .B(x[225]), .Z(n3876) );
  XNOR U5073 ( .A(n3877), .B(n3876), .Z(n3881) );
  AND U5074 ( .A(n3878), .B(o[33]), .Z(n3880) );
  XNOR U5075 ( .A(n3881), .B(n3880), .Z(n3886) );
  XNOR U5076 ( .A(n3887), .B(n3886), .Z(N99) );
  NAND U5077 ( .A(x[226]), .B(y[1825]), .Z(n3899) );
  NANDN U5078 ( .A(n3899), .B(n3879), .Z(n3883) );
  NAND U5079 ( .A(n3881), .B(n3880), .Z(n3882) );
  AND U5080 ( .A(n3883), .B(n3882), .Z(n3905) );
  NANDN U5081 ( .A(n3885), .B(n3884), .Z(n3889) );
  NAND U5082 ( .A(n3887), .B(n3886), .Z(n3888) );
  AND U5083 ( .A(n3889), .B(n3888), .Z(n3904) );
  XNOR U5084 ( .A(n3905), .B(n3904), .Z(n3907) );
  AND U5085 ( .A(x[225]), .B(y[1826]), .Z(n4018) );
  XOR U5086 ( .A(n4018), .B(n3901), .Z(n3903) );
  AND U5087 ( .A(y[1824]), .B(x[227]), .Z(n3891) );
  NAND U5088 ( .A(y[1827]), .B(x[224]), .Z(n3890) );
  XNOR U5089 ( .A(n3891), .B(n3890), .Z(n3893) );
  AND U5090 ( .A(n3892), .B(o[34]), .Z(n3894) );
  XOR U5091 ( .A(n3893), .B(n3894), .Z(n3902) );
  XOR U5092 ( .A(n3903), .B(n3902), .Z(n3906) );
  XOR U5093 ( .A(n3907), .B(n3906), .Z(N100) );
  AND U5094 ( .A(x[227]), .B(y[1827]), .Z(n3949) );
  NAND U5095 ( .A(n4520), .B(n3949), .Z(n3896) );
  NAND U5096 ( .A(n3894), .B(n3893), .Z(n3895) );
  AND U5097 ( .A(n3896), .B(n3895), .Z(n3931) );
  AND U5098 ( .A(y[1828]), .B(x[224]), .Z(n3898) );
  NAND U5099 ( .A(y[1824]), .B(x[228]), .Z(n3897) );
  XNOR U5100 ( .A(n3898), .B(n3897), .Z(n3922) );
  ANDN U5101 ( .B(o[35]), .A(n3899), .Z(n3921) );
  XOR U5102 ( .A(n3922), .B(n3921), .Z(n3929) );
  AND U5103 ( .A(x[226]), .B(y[1826]), .Z(n4064) );
  NAND U5104 ( .A(y[1827]), .B(x[225]), .Z(n3900) );
  XNOR U5105 ( .A(n4064), .B(n3900), .Z(n3918) );
  AND U5106 ( .A(x[227]), .B(y[1825]), .Z(n3913) );
  XOR U5107 ( .A(o[36]), .B(n3913), .Z(n3917) );
  XOR U5108 ( .A(n3918), .B(n3917), .Z(n3928) );
  XOR U5109 ( .A(n3929), .B(n3928), .Z(n3930) );
  XOR U5110 ( .A(n3931), .B(n3930), .Z(n3927) );
  NANDN U5111 ( .A(n3905), .B(n3904), .Z(n3909) );
  NAND U5112 ( .A(n3907), .B(n3906), .Z(n3908) );
  NAND U5113 ( .A(n3909), .B(n3908), .Z(n3926) );
  XOR U5114 ( .A(n3925), .B(n3926), .Z(n3910) );
  XNOR U5115 ( .A(n3927), .B(n3910), .Z(N101) );
  AND U5116 ( .A(y[1826]), .B(x[227]), .Z(n3912) );
  NAND U5117 ( .A(y[1828]), .B(x[225]), .Z(n3911) );
  XNOR U5118 ( .A(n3912), .B(n3911), .Z(n3936) );
  AND U5119 ( .A(x[228]), .B(y[1825]), .Z(n3945) );
  XOR U5120 ( .A(n3945), .B(o[37]), .Z(n3935) );
  XNOR U5121 ( .A(n3936), .B(n3935), .Z(n3939) );
  NAND U5122 ( .A(x[226]), .B(y[1827]), .Z(n4026) );
  AND U5123 ( .A(o[36]), .B(n3913), .Z(n3941) );
  AND U5124 ( .A(y[1824]), .B(x[229]), .Z(n3915) );
  NAND U5125 ( .A(y[1829]), .B(x[224]), .Z(n3914) );
  XNOR U5126 ( .A(n3915), .B(n3914), .Z(n3942) );
  XOR U5127 ( .A(n3941), .B(n3942), .Z(n3940) );
  XOR U5128 ( .A(n4026), .B(n3940), .Z(n3916) );
  XOR U5129 ( .A(n3939), .B(n3916), .Z(n3954) );
  NANDN U5130 ( .A(n4026), .B(n4018), .Z(n3920) );
  NAND U5131 ( .A(n3918), .B(n3917), .Z(n3919) );
  NAND U5132 ( .A(n3920), .B(n3919), .Z(n3952) );
  AND U5133 ( .A(x[228]), .B(y[1828]), .Z(n4722) );
  NAND U5134 ( .A(n4722), .B(n4520), .Z(n3924) );
  NAND U5135 ( .A(n3922), .B(n3921), .Z(n3923) );
  NAND U5136 ( .A(n3924), .B(n3923), .Z(n3951) );
  XOR U5137 ( .A(n3952), .B(n3951), .Z(n3953) );
  XOR U5138 ( .A(n3954), .B(n3953), .Z(n3960) );
  NAND U5139 ( .A(n3929), .B(n3928), .Z(n3933) );
  NANDN U5140 ( .A(n3931), .B(n3930), .Z(n3932) );
  AND U5141 ( .A(n3933), .B(n3932), .Z(n3959) );
  IV U5142 ( .A(n3959), .Z(n3957) );
  XOR U5143 ( .A(n3958), .B(n3957), .Z(n3934) );
  XNOR U5144 ( .A(n3960), .B(n3934), .Z(N102) );
  AND U5145 ( .A(x[227]), .B(y[1828]), .Z(n4027) );
  NAND U5146 ( .A(n4027), .B(n4018), .Z(n3938) );
  NAND U5147 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U5148 ( .A(n3938), .B(n3937), .Z(n3993) );
  XOR U5149 ( .A(n3993), .B(n3992), .Z(n3995) );
  AND U5150 ( .A(x[229]), .B(y[1829]), .Z(n4188) );
  NAND U5151 ( .A(n4520), .B(n4188), .Z(n3944) );
  NAND U5152 ( .A(n3942), .B(n3941), .Z(n3943) );
  NAND U5153 ( .A(n3944), .B(n3943), .Z(n3966) );
  AND U5154 ( .A(n3945), .B(o[37]), .Z(n3972) );
  AND U5155 ( .A(y[1824]), .B(x[230]), .Z(n3947) );
  NAND U5156 ( .A(y[1830]), .B(x[224]), .Z(n3946) );
  XNOR U5157 ( .A(n3947), .B(n3946), .Z(n3973) );
  XOR U5158 ( .A(n3972), .B(n3973), .Z(n3965) );
  XOR U5159 ( .A(n3966), .B(n3965), .Z(n3968) );
  NAND U5160 ( .A(y[1828]), .B(x[226]), .Z(n3948) );
  XNOR U5161 ( .A(n3949), .B(n3948), .Z(n3977) );
  AND U5162 ( .A(y[1829]), .B(x[225]), .Z(n4235) );
  NAND U5163 ( .A(y[1826]), .B(x[228]), .Z(n3950) );
  XNOR U5164 ( .A(n4235), .B(n3950), .Z(n3981) );
  NAND U5165 ( .A(x[229]), .B(y[1825]), .Z(n3988) );
  XOR U5166 ( .A(n3981), .B(n3980), .Z(n3976) );
  XOR U5167 ( .A(n3977), .B(n3976), .Z(n3967) );
  XOR U5168 ( .A(n3968), .B(n3967), .Z(n3994) );
  XNOR U5169 ( .A(n3995), .B(n3994), .Z(n3991) );
  NAND U5170 ( .A(n3952), .B(n3951), .Z(n3956) );
  NAND U5171 ( .A(n3954), .B(n3953), .Z(n3955) );
  NAND U5172 ( .A(n3956), .B(n3955), .Z(n3990) );
  NANDN U5173 ( .A(n3957), .B(n3958), .Z(n3963) );
  NOR U5174 ( .A(n3959), .B(n3958), .Z(n3961) );
  OR U5175 ( .A(n3961), .B(n3960), .Z(n3962) );
  AND U5176 ( .A(n3963), .B(n3962), .Z(n3989) );
  XOR U5177 ( .A(n3990), .B(n3989), .Z(n3964) );
  XNOR U5178 ( .A(n3991), .B(n3964), .Z(N103) );
  NAND U5179 ( .A(n3966), .B(n3965), .Z(n3970) );
  NAND U5180 ( .A(n3968), .B(n3967), .Z(n3969) );
  AND U5181 ( .A(n3970), .B(n3969), .Z(n4002) );
  AND U5182 ( .A(y[1826]), .B(x[229]), .Z(n4109) );
  NAND U5183 ( .A(y[1830]), .B(x[225]), .Z(n3971) );
  XNOR U5184 ( .A(n4109), .B(n3971), .Z(n4020) );
  NAND U5185 ( .A(x[230]), .B(y[1825]), .Z(n4024) );
  XOR U5186 ( .A(n4020), .B(n4019), .Z(n4038) );
  AND U5187 ( .A(x[230]), .B(y[1830]), .Z(n4253) );
  NAND U5188 ( .A(n4520), .B(n4253), .Z(n3975) );
  NAND U5189 ( .A(n3973), .B(n3972), .Z(n3974) );
  AND U5190 ( .A(n3975), .B(n3974), .Z(n4037) );
  NANDN U5191 ( .A(n4026), .B(n4027), .Z(n3979) );
  NAND U5192 ( .A(n3977), .B(n3976), .Z(n3978) );
  AND U5193 ( .A(n3979), .B(n3978), .Z(n4039) );
  XOR U5194 ( .A(n4040), .B(n4039), .Z(n4000) );
  AND U5195 ( .A(x[228]), .B(y[1829]), .Z(n4525) );
  NAND U5196 ( .A(n4525), .B(n4018), .Z(n3983) );
  NAND U5197 ( .A(n3981), .B(n3980), .Z(n3982) );
  AND U5198 ( .A(n3983), .B(n3982), .Z(n4015) );
  AND U5199 ( .A(y[1829]), .B(x[226]), .Z(n3985) );
  NAND U5200 ( .A(y[1827]), .B(x[228]), .Z(n3984) );
  XNOR U5201 ( .A(n3985), .B(n3984), .Z(n4028) );
  XOR U5202 ( .A(n4028), .B(n4027), .Z(n4013) );
  AND U5203 ( .A(y[1824]), .B(x[231]), .Z(n3987) );
  NAND U5204 ( .A(y[1831]), .B(x[224]), .Z(n3986) );
  XNOR U5205 ( .A(n3987), .B(n3986), .Z(n4032) );
  ANDN U5206 ( .B(o[38]), .A(n3988), .Z(n4031) );
  XNOR U5207 ( .A(n4032), .B(n4031), .Z(n4012) );
  XOR U5208 ( .A(n4015), .B(n4014), .Z(n3999) );
  XOR U5209 ( .A(n4000), .B(n3999), .Z(n4001) );
  XNOR U5210 ( .A(n4002), .B(n4001), .Z(n4008) );
  NAND U5211 ( .A(n3993), .B(n3992), .Z(n3997) );
  NAND U5212 ( .A(n3995), .B(n3994), .Z(n3996) );
  AND U5213 ( .A(n3997), .B(n3996), .Z(n4007) );
  IV U5214 ( .A(n4007), .Z(n4005) );
  XOR U5215 ( .A(n4006), .B(n4005), .Z(n3998) );
  XNOR U5216 ( .A(n4008), .B(n3998), .Z(N104) );
  NAND U5217 ( .A(n4000), .B(n3999), .Z(n4004) );
  NAND U5218 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U5219 ( .A(n4004), .B(n4003), .Z(n4081) );
  NANDN U5220 ( .A(n4005), .B(n4006), .Z(n4011) );
  NOR U5221 ( .A(n4007), .B(n4006), .Z(n4009) );
  OR U5222 ( .A(n4009), .B(n4008), .Z(n4010) );
  AND U5223 ( .A(n4011), .B(n4010), .Z(n4080) );
  NANDN U5224 ( .A(n4013), .B(n4012), .Z(n4017) );
  NAND U5225 ( .A(n4015), .B(n4014), .Z(n4016) );
  AND U5226 ( .A(n4017), .B(n4016), .Z(n4077) );
  AND U5227 ( .A(x[229]), .B(y[1830]), .Z(n4180) );
  NAND U5228 ( .A(n4180), .B(n4018), .Z(n4022) );
  NAND U5229 ( .A(n4020), .B(n4019), .Z(n4021) );
  AND U5230 ( .A(n4022), .B(n4021), .Z(n4075) );
  AND U5231 ( .A(y[1827]), .B(x[229]), .Z(n4639) );
  NAND U5232 ( .A(y[1831]), .B(x[225]), .Z(n4023) );
  XNOR U5233 ( .A(n4639), .B(n4023), .Z(n4056) );
  ANDN U5234 ( .B(o[39]), .A(n4024), .Z(n4055) );
  XNOR U5235 ( .A(n4056), .B(n4055), .Z(n4060) );
  NAND U5236 ( .A(x[227]), .B(y[1829]), .Z(n4854) );
  AND U5237 ( .A(x[230]), .B(y[1826]), .Z(n4025) );
  AND U5238 ( .A(y[1830]), .B(x[226]), .Z(n4948) );
  XOR U5239 ( .A(n4025), .B(n4948), .Z(n4065) );
  XOR U5240 ( .A(n4722), .B(n4065), .Z(n4059) );
  XOR U5241 ( .A(n4060), .B(n4061), .Z(n4074) );
  XOR U5242 ( .A(n4077), .B(n4076), .Z(n4086) );
  NANDN U5243 ( .A(n4026), .B(n4525), .Z(n4030) );
  NAND U5244 ( .A(n4028), .B(n4027), .Z(n4029) );
  AND U5245 ( .A(n4030), .B(n4029), .Z(n4071) );
  AND U5246 ( .A(x[231]), .B(y[1831]), .Z(n4411) );
  NAND U5247 ( .A(n4520), .B(n4411), .Z(n4034) );
  NAND U5248 ( .A(n4032), .B(n4031), .Z(n4033) );
  AND U5249 ( .A(n4034), .B(n4033), .Z(n4069) );
  AND U5250 ( .A(y[1824]), .B(x[232]), .Z(n4036) );
  NAND U5251 ( .A(y[1832]), .B(x[224]), .Z(n4035) );
  XNOR U5252 ( .A(n4036), .B(n4035), .Z(n4046) );
  AND U5253 ( .A(x[231]), .B(y[1825]), .Z(n4051) );
  XOR U5254 ( .A(o[40]), .B(n4051), .Z(n4045) );
  XOR U5255 ( .A(n4046), .B(n4045), .Z(n4068) );
  NANDN U5256 ( .A(n4038), .B(n4037), .Z(n4042) );
  NAND U5257 ( .A(n4040), .B(n4039), .Z(n4041) );
  NAND U5258 ( .A(n4042), .B(n4041), .Z(n4083) );
  XNOR U5259 ( .A(n4080), .B(n4082), .Z(n4043) );
  XOR U5260 ( .A(n4081), .B(n4043), .Z(N105) );
  AND U5261 ( .A(x[232]), .B(y[1832]), .Z(n4044) );
  NAND U5262 ( .A(n4044), .B(n4520), .Z(n4048) );
  NAND U5263 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U5264 ( .A(n4048), .B(n4047), .Z(n4138) );
  AND U5265 ( .A(y[1828]), .B(x[229]), .Z(n4050) );
  NAND U5266 ( .A(y[1826]), .B(x[231]), .Z(n4049) );
  XNOR U5267 ( .A(n4050), .B(n4049), .Z(n4111) );
  AND U5268 ( .A(o[40]), .B(n4051), .Z(n4110) );
  XOR U5269 ( .A(n4111), .B(n4110), .Z(n4136) );
  AND U5270 ( .A(y[1824]), .B(x[233]), .Z(n4053) );
  NAND U5271 ( .A(y[1833]), .B(x[224]), .Z(n4052) );
  XNOR U5272 ( .A(n4053), .B(n4052), .Z(n4118) );
  AND U5273 ( .A(x[232]), .B(y[1825]), .Z(n4127) );
  XOR U5274 ( .A(o[41]), .B(n4127), .Z(n4117) );
  XNOR U5275 ( .A(n4118), .B(n4117), .Z(n4135) );
  XNOR U5276 ( .A(n4138), .B(n4137), .Z(n4132) );
  AND U5277 ( .A(y[1827]), .B(x[230]), .Z(n4470) );
  NAND U5278 ( .A(y[1832]), .B(x[225]), .Z(n4054) );
  XNOR U5279 ( .A(n4470), .B(n4054), .Z(n4122) );
  XOR U5280 ( .A(n4525), .B(n4122), .Z(n4142) );
  AND U5281 ( .A(x[226]), .B(y[1831]), .Z(n4765) );
  AND U5282 ( .A(x[227]), .B(y[1830]), .Z(n4480) );
  XOR U5283 ( .A(n4765), .B(n4480), .Z(n4141) );
  NAND U5284 ( .A(x[229]), .B(y[1831]), .Z(n4239) );
  AND U5285 ( .A(x[225]), .B(y[1827]), .Z(n4121) );
  NANDN U5286 ( .A(n4239), .B(n4121), .Z(n4058) );
  NAND U5287 ( .A(n4056), .B(n4055), .Z(n4057) );
  NAND U5288 ( .A(n4058), .B(n4057), .Z(n4129) );
  XOR U5289 ( .A(n4130), .B(n4129), .Z(n4131) );
  XNOR U5290 ( .A(n4132), .B(n4131), .Z(n4105) );
  NANDN U5291 ( .A(n4059), .B(n4854), .Z(n4063) );
  NANDN U5292 ( .A(n4061), .B(n4060), .Z(n4062) );
  NAND U5293 ( .A(n4063), .B(n4062), .Z(n4103) );
  NAND U5294 ( .A(n4253), .B(n4064), .Z(n4067) );
  NAND U5295 ( .A(n4722), .B(n4065), .Z(n4066) );
  AND U5296 ( .A(n4067), .B(n4066), .Z(n4104) );
  XNOR U5297 ( .A(n4103), .B(n4104), .Z(n4106) );
  NANDN U5298 ( .A(n4069), .B(n4068), .Z(n4073) );
  NANDN U5299 ( .A(n4071), .B(n4070), .Z(n4072) );
  AND U5300 ( .A(n4073), .B(n4072), .Z(n4091) );
  NANDN U5301 ( .A(n4075), .B(n4074), .Z(n4079) );
  NAND U5302 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U5303 ( .A(n4079), .B(n4078), .Z(n4090) );
  XNOR U5304 ( .A(n4092), .B(n4093), .Z(n4099) );
  NANDN U5305 ( .A(n4084), .B(n4083), .Z(n4088) );
  NANDN U5306 ( .A(n4086), .B(n4085), .Z(n4087) );
  AND U5307 ( .A(n4088), .B(n4087), .Z(n4097) );
  IV U5308 ( .A(n4097), .Z(n4096) );
  XOR U5309 ( .A(n4098), .B(n4096), .Z(n4089) );
  XNOR U5310 ( .A(n4099), .B(n4089), .Z(N106) );
  NANDN U5311 ( .A(n4091), .B(n4090), .Z(n4095) );
  NAND U5312 ( .A(n4093), .B(n4092), .Z(n4094) );
  NAND U5313 ( .A(n4095), .B(n4094), .Z(n4199) );
  IV U5314 ( .A(n4199), .Z(n4198) );
  OR U5315 ( .A(n4098), .B(n4096), .Z(n4102) );
  ANDN U5316 ( .B(n4098), .A(n4097), .Z(n4100) );
  OR U5317 ( .A(n4100), .B(n4099), .Z(n4101) );
  AND U5318 ( .A(n4102), .B(n4101), .Z(n4200) );
  NAND U5319 ( .A(n4104), .B(n4103), .Z(n4108) );
  NANDN U5320 ( .A(n4106), .B(n4105), .Z(n4107) );
  NAND U5321 ( .A(n4108), .B(n4107), .Z(n4207) );
  AND U5322 ( .A(x[231]), .B(y[1828]), .Z(n4182) );
  NAND U5323 ( .A(n4182), .B(n4109), .Z(n4113) );
  NAND U5324 ( .A(n4111), .B(n4110), .Z(n4112) );
  AND U5325 ( .A(n4113), .B(n4112), .Z(n4195) );
  AND U5326 ( .A(y[1827]), .B(x[231]), .Z(n4115) );
  NAND U5327 ( .A(y[1830]), .B(x[228]), .Z(n4114) );
  XNOR U5328 ( .A(n4115), .B(n4114), .Z(n4166) );
  AND U5329 ( .A(x[230]), .B(y[1828]), .Z(n4165) );
  XNOR U5330 ( .A(n4166), .B(n4165), .Z(n4193) );
  AND U5331 ( .A(x[232]), .B(y[1826]), .Z(n4375) );
  NAND U5332 ( .A(x[233]), .B(y[1825]), .Z(n4176) );
  XNOR U5333 ( .A(o[42]), .B(n4176), .Z(n4187) );
  XOR U5334 ( .A(n4375), .B(n4187), .Z(n4189) );
  XNOR U5335 ( .A(n4189), .B(n4188), .Z(n4192) );
  XOR U5336 ( .A(n4193), .B(n4192), .Z(n4194) );
  XOR U5337 ( .A(n4195), .B(n4194), .Z(n4155) );
  AND U5338 ( .A(x[233]), .B(y[1833]), .Z(n4116) );
  NAND U5339 ( .A(n4116), .B(n4520), .Z(n4120) );
  NAND U5340 ( .A(n4118), .B(n4117), .Z(n4119) );
  AND U5341 ( .A(n4120), .B(n4119), .Z(n4153) );
  AND U5342 ( .A(x[230]), .B(y[1832]), .Z(n4402) );
  NAND U5343 ( .A(n4402), .B(n4121), .Z(n4124) );
  NAND U5344 ( .A(n4525), .B(n4122), .Z(n4123) );
  NAND U5345 ( .A(n4124), .B(n4123), .Z(n4161) );
  AND U5346 ( .A(y[1824]), .B(x[234]), .Z(n4126) );
  NAND U5347 ( .A(y[1834]), .B(x[224]), .Z(n4125) );
  XNOR U5348 ( .A(n4126), .B(n4125), .Z(n4171) );
  AND U5349 ( .A(o[41]), .B(n4127), .Z(n4170) );
  XOR U5350 ( .A(n4171), .B(n4170), .Z(n4159) );
  AND U5351 ( .A(y[1831]), .B(x[227]), .Z(n5084) );
  NAND U5352 ( .A(y[1833]), .B(x[225]), .Z(n4128) );
  XNOR U5353 ( .A(n5084), .B(n4128), .Z(n4183) );
  AND U5354 ( .A(x[226]), .B(y[1832]), .Z(n4184) );
  XOR U5355 ( .A(n4183), .B(n4184), .Z(n4158) );
  XOR U5356 ( .A(n4159), .B(n4158), .Z(n4160) );
  XOR U5357 ( .A(n4161), .B(n4160), .Z(n4152) );
  NAND U5358 ( .A(n4130), .B(n4129), .Z(n4134) );
  NAND U5359 ( .A(n4132), .B(n4131), .Z(n4133) );
  AND U5360 ( .A(n4134), .B(n4133), .Z(n4149) );
  NANDN U5361 ( .A(n4136), .B(n4135), .Z(n4140) );
  NAND U5362 ( .A(n4138), .B(n4137), .Z(n4139) );
  AND U5363 ( .A(n4140), .B(n4139), .Z(n4146) );
  NOR U5364 ( .A(n4480), .B(n4765), .Z(n4144) );
  NANDN U5365 ( .A(n4142), .B(n4141), .Z(n4143) );
  NANDN U5366 ( .A(n4144), .B(n4143), .Z(n4147) );
  XOR U5367 ( .A(n4149), .B(n4148), .Z(n4205) );
  XOR U5368 ( .A(n4207), .B(n4208), .Z(n4201) );
  XNOR U5369 ( .A(n4200), .B(n4201), .Z(n4145) );
  XOR U5370 ( .A(n4198), .B(n4145), .Z(N107) );
  NANDN U5371 ( .A(n4147), .B(n4146), .Z(n4151) );
  NANDN U5372 ( .A(n4149), .B(n4148), .Z(n4150) );
  AND U5373 ( .A(n4151), .B(n4150), .Z(n4215) );
  NANDN U5374 ( .A(n4153), .B(n4152), .Z(n4157) );
  NANDN U5375 ( .A(n4155), .B(n4154), .Z(n4156) );
  AND U5376 ( .A(n4157), .B(n4156), .Z(n4213) );
  NAND U5377 ( .A(n4159), .B(n4158), .Z(n4163) );
  NAND U5378 ( .A(n4161), .B(n4160), .Z(n4162) );
  NAND U5379 ( .A(n4163), .B(n4162), .Z(n4273) );
  AND U5380 ( .A(x[231]), .B(y[1830]), .Z(n4299) );
  AND U5381 ( .A(x[228]), .B(y[1827]), .Z(n4164) );
  NAND U5382 ( .A(n4299), .B(n4164), .Z(n4168) );
  NAND U5383 ( .A(n4166), .B(n4165), .Z(n4167) );
  NAND U5384 ( .A(n4168), .B(n4167), .Z(n4271) );
  AND U5385 ( .A(x[234]), .B(y[1834]), .Z(n4169) );
  NAND U5386 ( .A(n4169), .B(n4520), .Z(n4173) );
  NAND U5387 ( .A(n4171), .B(n4170), .Z(n4172) );
  NAND U5388 ( .A(n4173), .B(n4172), .Z(n4267) );
  AND U5389 ( .A(y[1824]), .B(x[235]), .Z(n4175) );
  NAND U5390 ( .A(y[1835]), .B(x[224]), .Z(n4174) );
  XNOR U5391 ( .A(n4175), .B(n4174), .Z(n4245) );
  ANDN U5392 ( .B(o[42]), .A(n4176), .Z(n4244) );
  XOR U5393 ( .A(n4245), .B(n4244), .Z(n4266) );
  AND U5394 ( .A(y[1829]), .B(x[230]), .Z(n4178) );
  NAND U5395 ( .A(y[1834]), .B(x[225]), .Z(n4177) );
  XNOR U5396 ( .A(n4178), .B(n4177), .Z(n4237) );
  AND U5397 ( .A(x[234]), .B(y[1825]), .Z(n4251) );
  XOR U5398 ( .A(o[43]), .B(n4251), .Z(n4236) );
  XOR U5399 ( .A(n4237), .B(n4236), .Z(n4265) );
  XOR U5400 ( .A(n4266), .B(n4265), .Z(n4268) );
  XOR U5401 ( .A(n4267), .B(n4268), .Z(n4272) );
  XNOR U5402 ( .A(n4271), .B(n4272), .Z(n4274) );
  XOR U5403 ( .A(n4273), .B(n4274), .Z(n4256) );
  AND U5404 ( .A(x[227]), .B(y[1832]), .Z(n5213) );
  NAND U5405 ( .A(y[1833]), .B(x[226]), .Z(n4179) );
  XNOR U5406 ( .A(n4180), .B(n4179), .Z(n4232) );
  AND U5407 ( .A(x[228]), .B(y[1831]), .Z(n4231) );
  XNOR U5408 ( .A(n4232), .B(n4231), .Z(n4260) );
  XNOR U5409 ( .A(n5213), .B(n4260), .Z(n4262) );
  NAND U5410 ( .A(y[1826]), .B(x[233]), .Z(n4181) );
  XNOR U5411 ( .A(n4182), .B(n4181), .Z(n4248) );
  AND U5412 ( .A(x[232]), .B(y[1827]), .Z(n4247) );
  XNOR U5413 ( .A(n4248), .B(n4247), .Z(n4261) );
  XNOR U5414 ( .A(n4262), .B(n4261), .Z(n4228) );
  NAND U5415 ( .A(x[227]), .B(y[1833]), .Z(n4295) );
  AND U5416 ( .A(x[225]), .B(y[1831]), .Z(n4515) );
  NANDN U5417 ( .A(n4295), .B(n4515), .Z(n4186) );
  NAND U5418 ( .A(n4184), .B(n4183), .Z(n4185) );
  NAND U5419 ( .A(n4186), .B(n4185), .Z(n4226) );
  NAND U5420 ( .A(n4187), .B(n4375), .Z(n4191) );
  NAND U5421 ( .A(n4189), .B(n4188), .Z(n4190) );
  NAND U5422 ( .A(n4191), .B(n4190), .Z(n4225) );
  XOR U5423 ( .A(n4226), .B(n4225), .Z(n4227) );
  XNOR U5424 ( .A(n4228), .B(n4227), .Z(n4255) );
  NAND U5425 ( .A(n4193), .B(n4192), .Z(n4197) );
  NAND U5426 ( .A(n4195), .B(n4194), .Z(n4196) );
  NAND U5427 ( .A(n4197), .B(n4196), .Z(n4254) );
  XOR U5428 ( .A(n4255), .B(n4254), .Z(n4257) );
  XNOR U5429 ( .A(n4256), .B(n4257), .Z(n4212) );
  XOR U5430 ( .A(n4215), .B(n4214), .Z(n4221) );
  OR U5431 ( .A(n4200), .B(n4198), .Z(n4204) );
  ANDN U5432 ( .B(n4200), .A(n4199), .Z(n4202) );
  OR U5433 ( .A(n4202), .B(n4201), .Z(n4203) );
  AND U5434 ( .A(n4204), .B(n4203), .Z(n4220) );
  NANDN U5435 ( .A(n4206), .B(n4205), .Z(n4210) );
  NAND U5436 ( .A(n4208), .B(n4207), .Z(n4209) );
  AND U5437 ( .A(n4210), .B(n4209), .Z(n4219) );
  IV U5438 ( .A(n4219), .Z(n4218) );
  XOR U5439 ( .A(n4220), .B(n4218), .Z(n4211) );
  XNOR U5440 ( .A(n4221), .B(n4211), .Z(N108) );
  NANDN U5441 ( .A(n4213), .B(n4212), .Z(n4217) );
  NANDN U5442 ( .A(n4215), .B(n4214), .Z(n4216) );
  NAND U5443 ( .A(n4217), .B(n4216), .Z(n4340) );
  IV U5444 ( .A(n4340), .Z(n4339) );
  OR U5445 ( .A(n4220), .B(n4218), .Z(n4224) );
  ANDN U5446 ( .B(n4220), .A(n4219), .Z(n4222) );
  OR U5447 ( .A(n4222), .B(n4221), .Z(n4223) );
  AND U5448 ( .A(n4224), .B(n4223), .Z(n4341) );
  NAND U5449 ( .A(n4226), .B(n4225), .Z(n4230) );
  NAND U5450 ( .A(n4228), .B(n4227), .Z(n4229) );
  NAND U5451 ( .A(n4230), .B(n4229), .Z(n4335) );
  AND U5452 ( .A(x[229]), .B(y[1833]), .Z(n4756) );
  NAND U5453 ( .A(n4948), .B(n4756), .Z(n4234) );
  NAND U5454 ( .A(n4232), .B(n4231), .Z(n4233) );
  AND U5455 ( .A(n4234), .B(n4233), .Z(n4285) );
  AND U5456 ( .A(x[230]), .B(y[1834]), .Z(n4532) );
  XNOR U5457 ( .A(n4285), .B(n4284), .Z(n4287) );
  AND U5458 ( .A(x[233]), .B(y[1827]), .Z(n4943) );
  AND U5459 ( .A(y[1826]), .B(x[234]), .Z(n4985) );
  NAND U5460 ( .A(y[1832]), .B(x[228]), .Z(n4238) );
  XNOR U5461 ( .A(n4985), .B(n4238), .Z(n4326) );
  XOR U5462 ( .A(n4943), .B(n4326), .Z(n4305) );
  IV U5463 ( .A(n4239), .Z(n4304) );
  NAND U5464 ( .A(x[231]), .B(y[1829]), .Z(n4303) );
  XNOR U5465 ( .A(n4304), .B(n4303), .Z(n4306) );
  AND U5466 ( .A(y[1824]), .B(x[236]), .Z(n4241) );
  NAND U5467 ( .A(y[1836]), .B(x[224]), .Z(n4240) );
  XNOR U5468 ( .A(n4241), .B(n4240), .Z(n4320) );
  AND U5469 ( .A(x[235]), .B(y[1825]), .Z(n4300) );
  XOR U5470 ( .A(o[44]), .B(n4300), .Z(n4319) );
  XOR U5471 ( .A(n4320), .B(n4319), .Z(n4288) );
  AND U5472 ( .A(y[1834]), .B(x[226]), .Z(n4243) );
  NAND U5473 ( .A(y[1828]), .B(x[232]), .Z(n4242) );
  XNOR U5474 ( .A(n4243), .B(n4242), .Z(n4294) );
  XNOR U5475 ( .A(n4288), .B(n4289), .Z(n4290) );
  XOR U5476 ( .A(n4291), .B(n4290), .Z(n4286) );
  XOR U5477 ( .A(n4287), .B(n4286), .Z(n4334) );
  AND U5478 ( .A(x[235]), .B(y[1835]), .Z(n5336) );
  AND U5479 ( .A(x[231]), .B(y[1826]), .Z(n4456) );
  AND U5480 ( .A(x[233]), .B(y[1828]), .Z(n4246) );
  NAND U5481 ( .A(n4456), .B(n4246), .Z(n4250) );
  NAND U5482 ( .A(n4248), .B(n4247), .Z(n4249) );
  AND U5483 ( .A(n4250), .B(n4249), .Z(n4310) );
  AND U5484 ( .A(o[43]), .B(n4251), .Z(n4315) );
  NAND U5485 ( .A(y[1835]), .B(x[225]), .Z(n4252) );
  XNOR U5486 ( .A(n4253), .B(n4252), .Z(n4316) );
  XOR U5487 ( .A(n4315), .B(n4316), .Z(n4309) );
  XNOR U5488 ( .A(n4310), .B(n4309), .Z(n4311) );
  XNOR U5489 ( .A(n4312), .B(n4311), .Z(n4333) );
  XOR U5490 ( .A(n4334), .B(n4333), .Z(n4336) );
  XNOR U5491 ( .A(n4335), .B(n4336), .Z(n4347) );
  NAND U5492 ( .A(n4255), .B(n4254), .Z(n4259) );
  NAND U5493 ( .A(n4257), .B(n4256), .Z(n4258) );
  NAND U5494 ( .A(n4259), .B(n4258), .Z(n4346) );
  XOR U5495 ( .A(n4347), .B(n4346), .Z(n4349) );
  NANDN U5496 ( .A(n5213), .B(n4260), .Z(n4264) );
  NAND U5497 ( .A(n4262), .B(n4261), .Z(n4263) );
  NAND U5498 ( .A(n4264), .B(n4263), .Z(n4278) );
  NAND U5499 ( .A(n4266), .B(n4265), .Z(n4270) );
  NAND U5500 ( .A(n4268), .B(n4267), .Z(n4269) );
  AND U5501 ( .A(n4270), .B(n4269), .Z(n4279) );
  XOR U5502 ( .A(n4278), .B(n4279), .Z(n4281) );
  NAND U5503 ( .A(n4272), .B(n4271), .Z(n4276) );
  NANDN U5504 ( .A(n4274), .B(n4273), .Z(n4275) );
  AND U5505 ( .A(n4276), .B(n4275), .Z(n4280) );
  XOR U5506 ( .A(n4281), .B(n4280), .Z(n4348) );
  XOR U5507 ( .A(n4349), .B(n4348), .Z(n4342) );
  XNOR U5508 ( .A(n4341), .B(n4342), .Z(n4277) );
  XOR U5509 ( .A(n4339), .B(n4277), .Z(N109) );
  NAND U5510 ( .A(n4279), .B(n4278), .Z(n4283) );
  NAND U5511 ( .A(n4281), .B(n4280), .Z(n4282) );
  NAND U5512 ( .A(n4283), .B(n4282), .Z(n4427) );
  NANDN U5513 ( .A(n4289), .B(n4288), .Z(n4293) );
  NAND U5514 ( .A(n4291), .B(n4290), .Z(n4292) );
  NAND U5515 ( .A(n4293), .B(n4292), .Z(n4359) );
  AND U5516 ( .A(y[1834]), .B(x[232]), .Z(n5637) );
  AND U5517 ( .A(x[226]), .B(y[1828]), .Z(n4466) );
  NAND U5518 ( .A(n5637), .B(n4466), .Z(n4297) );
  NANDN U5519 ( .A(n4295), .B(n4294), .Z(n4296) );
  NAND U5520 ( .A(n4297), .B(n4296), .Z(n4390) );
  NAND U5521 ( .A(y[1836]), .B(x[225]), .Z(n4298) );
  XNOR U5522 ( .A(n4299), .B(n4298), .Z(n4381) );
  AND U5523 ( .A(o[44]), .B(n4300), .Z(n4380) );
  XOR U5524 ( .A(n4381), .B(n4380), .Z(n4388) );
  AND U5525 ( .A(x[230]), .B(y[1831]), .Z(n5376) );
  AND U5526 ( .A(y[1835]), .B(x[226]), .Z(n4302) );
  NAND U5527 ( .A(y[1828]), .B(x[233]), .Z(n4301) );
  XNOR U5528 ( .A(n4302), .B(n4301), .Z(n4404) );
  XOR U5529 ( .A(n5376), .B(n4404), .Z(n4387) );
  XOR U5530 ( .A(n4388), .B(n4387), .Z(n4389) );
  XOR U5531 ( .A(n4390), .B(n4389), .Z(n4358) );
  NANDN U5532 ( .A(n4304), .B(n4303), .Z(n4308) );
  ANDN U5533 ( .B(n4306), .A(n4305), .Z(n4307) );
  ANDN U5534 ( .B(n4308), .A(n4307), .Z(n4357) );
  XOR U5535 ( .A(n4358), .B(n4357), .Z(n4360) );
  XOR U5536 ( .A(n4359), .B(n4360), .Z(n4353) );
  XNOR U5537 ( .A(n4354), .B(n4353), .Z(n4356) );
  NANDN U5538 ( .A(n4310), .B(n4309), .Z(n4314) );
  NANDN U5539 ( .A(n4312), .B(n4311), .Z(n4313) );
  NAND U5540 ( .A(n4314), .B(n4313), .Z(n4366) );
  AND U5541 ( .A(x[230]), .B(y[1835]), .Z(n4696) );
  IV U5542 ( .A(n4696), .Z(n4758) );
  AND U5543 ( .A(x[225]), .B(y[1830]), .Z(n4379) );
  NANDN U5544 ( .A(n4758), .B(n4379), .Z(n4318) );
  NAND U5545 ( .A(n4316), .B(n4315), .Z(n4317) );
  NAND U5546 ( .A(n4318), .B(n4317), .Z(n4372) );
  AND U5547 ( .A(x[236]), .B(y[1836]), .Z(n5645) );
  NAND U5548 ( .A(n5645), .B(n4520), .Z(n4322) );
  NAND U5549 ( .A(n4320), .B(n4319), .Z(n4321) );
  NAND U5550 ( .A(n4322), .B(n4321), .Z(n4370) );
  AND U5551 ( .A(x[234]), .B(y[1827]), .Z(n5225) );
  AND U5552 ( .A(y[1826]), .B(x[235]), .Z(n5186) );
  NAND U5553 ( .A(y[1829]), .B(x[232]), .Z(n4323) );
  XNOR U5554 ( .A(n5186), .B(n4323), .Z(n4376) );
  XOR U5555 ( .A(n5225), .B(n4376), .Z(n4369) );
  XOR U5556 ( .A(n4370), .B(n4369), .Z(n4371) );
  XOR U5557 ( .A(n4372), .B(n4371), .Z(n4364) );
  AND U5558 ( .A(x[234]), .B(y[1832]), .Z(n4325) );
  AND U5559 ( .A(x[228]), .B(y[1826]), .Z(n4324) );
  NAND U5560 ( .A(n4325), .B(n4324), .Z(n4328) );
  NAND U5561 ( .A(n4326), .B(n4943), .Z(n4327) );
  NAND U5562 ( .A(n4328), .B(n4327), .Z(n4415) );
  AND U5563 ( .A(y[1824]), .B(x[237]), .Z(n4330) );
  NAND U5564 ( .A(y[1837]), .B(x[224]), .Z(n4329) );
  XNOR U5565 ( .A(n4330), .B(n4329), .Z(n4398) );
  AND U5566 ( .A(x[236]), .B(y[1825]), .Z(n4409) );
  XOR U5567 ( .A(o[45]), .B(n4409), .Z(n4397) );
  XOR U5568 ( .A(n4398), .B(n4397), .Z(n4413) );
  AND U5569 ( .A(y[1832]), .B(x[229]), .Z(n4332) );
  NAND U5570 ( .A(y[1834]), .B(x[227]), .Z(n4331) );
  XNOR U5571 ( .A(n4332), .B(n4331), .Z(n4393) );
  AND U5572 ( .A(x[228]), .B(y[1833]), .Z(n4394) );
  XOR U5573 ( .A(n4393), .B(n4394), .Z(n4412) );
  XOR U5574 ( .A(n4413), .B(n4412), .Z(n4414) );
  XOR U5575 ( .A(n4415), .B(n4414), .Z(n4363) );
  XOR U5576 ( .A(n4364), .B(n4363), .Z(n4365) );
  XOR U5577 ( .A(n4366), .B(n4365), .Z(n4355) );
  XNOR U5578 ( .A(n4356), .B(n4355), .Z(n4426) );
  NAND U5579 ( .A(n4334), .B(n4333), .Z(n4338) );
  NAND U5580 ( .A(n4336), .B(n4335), .Z(n4337) );
  AND U5581 ( .A(n4338), .B(n4337), .Z(n4425) );
  XNOR U5582 ( .A(n4426), .B(n4425), .Z(n4428) );
  XOR U5583 ( .A(n4427), .B(n4428), .Z(n4421) );
  OR U5584 ( .A(n4341), .B(n4339), .Z(n4345) );
  ANDN U5585 ( .B(n4341), .A(n4340), .Z(n4343) );
  OR U5586 ( .A(n4343), .B(n4342), .Z(n4344) );
  AND U5587 ( .A(n4345), .B(n4344), .Z(n4419) );
  NAND U5588 ( .A(n4347), .B(n4346), .Z(n4351) );
  NAND U5589 ( .A(n4349), .B(n4348), .Z(n4350) );
  NAND U5590 ( .A(n4351), .B(n4350), .Z(n4420) );
  IV U5591 ( .A(n4420), .Z(n4418) );
  XOR U5592 ( .A(n4419), .B(n4418), .Z(n4352) );
  XNOR U5593 ( .A(n4421), .B(n4352), .Z(N110) );
  NAND U5594 ( .A(n4358), .B(n4357), .Z(n4362) );
  NAND U5595 ( .A(n4360), .B(n4359), .Z(n4361) );
  NAND U5596 ( .A(n4362), .B(n4361), .Z(n4507) );
  XNOR U5597 ( .A(n4508), .B(n4507), .Z(n4510) );
  NAND U5598 ( .A(n4364), .B(n4363), .Z(n4368) );
  NAND U5599 ( .A(n4366), .B(n4365), .Z(n4367) );
  NAND U5600 ( .A(n4368), .B(n4367), .Z(n4435) );
  NAND U5601 ( .A(n4370), .B(n4369), .Z(n4374) );
  NAND U5602 ( .A(n4372), .B(n4371), .Z(n4373) );
  AND U5603 ( .A(n4374), .B(n4373), .Z(n4441) );
  AND U5604 ( .A(x[235]), .B(y[1829]), .Z(n4547) );
  NAND U5605 ( .A(n4547), .B(n4375), .Z(n4378) );
  NAND U5606 ( .A(n4376), .B(n5225), .Z(n4377) );
  NAND U5607 ( .A(n4378), .B(n4377), .Z(n4496) );
  NAND U5608 ( .A(x[231]), .B(y[1836]), .Z(n4958) );
  NANDN U5609 ( .A(n4958), .B(n4379), .Z(n4383) );
  NAND U5610 ( .A(n4381), .B(n4380), .Z(n4382) );
  NAND U5611 ( .A(n4383), .B(n4382), .Z(n4495) );
  XOR U5612 ( .A(n4496), .B(n4495), .Z(n4498) );
  AND U5613 ( .A(x[228]), .B(y[1834]), .Z(n4863) );
  AND U5614 ( .A(y[1835]), .B(x[227]), .Z(n4385) );
  NAND U5615 ( .A(y[1830]), .B(x[232]), .Z(n4384) );
  XNOR U5616 ( .A(n4385), .B(n4384), .Z(n4481) );
  XOR U5617 ( .A(n4756), .B(n4481), .Z(n4490) );
  XOR U5618 ( .A(n4863), .B(n4490), .Z(n4492) );
  AND U5619 ( .A(x[233]), .B(y[1829]), .Z(n5039) );
  AND U5620 ( .A(y[1836]), .B(x[226]), .Z(n4386) );
  AND U5621 ( .A(y[1828]), .B(x[234]), .Z(n5079) );
  XOR U5622 ( .A(n4386), .B(n5079), .Z(n4467) );
  XOR U5623 ( .A(n5039), .B(n4467), .Z(n4491) );
  XOR U5624 ( .A(n4492), .B(n4491), .Z(n4497) );
  XNOR U5625 ( .A(n4498), .B(n4497), .Z(n4439) );
  NAND U5626 ( .A(n4388), .B(n4387), .Z(n4392) );
  NAND U5627 ( .A(n4390), .B(n4389), .Z(n4391) );
  AND U5628 ( .A(n4392), .B(n4391), .Z(n4438) );
  XOR U5629 ( .A(n4439), .B(n4438), .Z(n4440) );
  XNOR U5630 ( .A(n4441), .B(n4440), .Z(n4433) );
  NAND U5631 ( .A(x[229]), .B(y[1834]), .Z(n4534) );
  NANDN U5632 ( .A(n4534), .B(n5213), .Z(n4396) );
  NAND U5633 ( .A(n4394), .B(n4393), .Z(n4395) );
  NAND U5634 ( .A(n4396), .B(n4395), .Z(n4447) );
  AND U5635 ( .A(x[237]), .B(y[1837]), .Z(n5987) );
  NAND U5636 ( .A(n5987), .B(n4520), .Z(n4400) );
  NAND U5637 ( .A(n4398), .B(n4397), .Z(n4399) );
  NAND U5638 ( .A(n4400), .B(n4399), .Z(n4445) );
  NAND U5639 ( .A(y[1827]), .B(x[235]), .Z(n4401) );
  XNOR U5640 ( .A(n4402), .B(n4401), .Z(n4471) );
  AND U5641 ( .A(x[225]), .B(y[1837]), .Z(n4472) );
  XOR U5642 ( .A(n4471), .B(n4472), .Z(n4444) );
  XOR U5643 ( .A(n4445), .B(n4444), .Z(n4446) );
  XNOR U5644 ( .A(n4447), .B(n4446), .Z(n4502) );
  AND U5645 ( .A(x[233]), .B(y[1835]), .Z(n4403) );
  NAND U5646 ( .A(n4403), .B(n4466), .Z(n4406) );
  NAND U5647 ( .A(n4404), .B(n5376), .Z(n4405) );
  AND U5648 ( .A(n4406), .B(n4405), .Z(n4453) );
  AND U5649 ( .A(y[1824]), .B(x[238]), .Z(n4408) );
  NAND U5650 ( .A(y[1838]), .B(x[224]), .Z(n4407) );
  XNOR U5651 ( .A(n4408), .B(n4407), .Z(n4476) );
  AND U5652 ( .A(o[45]), .B(n4409), .Z(n4475) );
  XOR U5653 ( .A(n4476), .B(n4475), .Z(n4451) );
  NAND U5654 ( .A(y[1826]), .B(x[236]), .Z(n4410) );
  XNOR U5655 ( .A(n4411), .B(n4410), .Z(n4457) );
  NAND U5656 ( .A(x[237]), .B(y[1825]), .Z(n4465) );
  XNOR U5657 ( .A(o[46]), .B(n4465), .Z(n4458) );
  XOR U5658 ( .A(n4457), .B(n4458), .Z(n4450) );
  XOR U5659 ( .A(n4451), .B(n4450), .Z(n4452) );
  XOR U5660 ( .A(n4453), .B(n4452), .Z(n4501) );
  XOR U5661 ( .A(n4502), .B(n4501), .Z(n4504) );
  NAND U5662 ( .A(n4413), .B(n4412), .Z(n4417) );
  NAND U5663 ( .A(n4415), .B(n4414), .Z(n4416) );
  AND U5664 ( .A(n4417), .B(n4416), .Z(n4503) );
  XNOR U5665 ( .A(n4504), .B(n4503), .Z(n4432) );
  XOR U5666 ( .A(n4433), .B(n4432), .Z(n4434) );
  XOR U5667 ( .A(n4435), .B(n4434), .Z(n4509) );
  XOR U5668 ( .A(n4510), .B(n4509), .Z(n4513) );
  NANDN U5669 ( .A(n4418), .B(n4419), .Z(n4424) );
  NOR U5670 ( .A(n4420), .B(n4419), .Z(n4422) );
  OR U5671 ( .A(n4422), .B(n4421), .Z(n4423) );
  AND U5672 ( .A(n4424), .B(n4423), .Z(n4512) );
  NAND U5673 ( .A(n4426), .B(n4425), .Z(n4430) );
  NANDN U5674 ( .A(n4428), .B(n4427), .Z(n4429) );
  NAND U5675 ( .A(n4430), .B(n4429), .Z(n4511) );
  XOR U5676 ( .A(n4512), .B(n4511), .Z(n4431) );
  XNOR U5677 ( .A(n4513), .B(n4431), .Z(N111) );
  NAND U5678 ( .A(n4433), .B(n4432), .Z(n4437) );
  NAND U5679 ( .A(n4435), .B(n4434), .Z(n4436) );
  AND U5680 ( .A(n4437), .B(n4436), .Z(n4604) );
  NAND U5681 ( .A(n4439), .B(n4438), .Z(n4443) );
  NAND U5682 ( .A(n4441), .B(n4440), .Z(n4442) );
  NAND U5683 ( .A(n4443), .B(n4442), .Z(n4576) );
  NAND U5684 ( .A(n4445), .B(n4444), .Z(n4449) );
  NAND U5685 ( .A(n4447), .B(n4446), .Z(n4448) );
  NAND U5686 ( .A(n4449), .B(n4448), .Z(n4583) );
  NAND U5687 ( .A(n4451), .B(n4450), .Z(n4455) );
  NANDN U5688 ( .A(n4453), .B(n4452), .Z(n4454) );
  NAND U5689 ( .A(n4455), .B(n4454), .Z(n4581) );
  NAND U5690 ( .A(x[236]), .B(y[1831]), .Z(n4950) );
  NANDN U5691 ( .A(n4950), .B(n4456), .Z(n4460) );
  NAND U5692 ( .A(n4458), .B(n4457), .Z(n4459) );
  AND U5693 ( .A(n4460), .B(n4459), .Z(n4557) );
  AND U5694 ( .A(y[1828]), .B(x[235]), .Z(n4462) );
  NAND U5695 ( .A(y[1826]), .B(x[237]), .Z(n4461) );
  XNOR U5696 ( .A(n4462), .B(n4461), .Z(n4561) );
  AND U5697 ( .A(x[236]), .B(y[1827]), .Z(n4560) );
  XNOR U5698 ( .A(n4561), .B(n4560), .Z(n4555) );
  AND U5699 ( .A(y[1824]), .B(x[239]), .Z(n4464) );
  NAND U5700 ( .A(y[1839]), .B(x[224]), .Z(n4463) );
  XNOR U5701 ( .A(n4464), .B(n4463), .Z(n4522) );
  ANDN U5702 ( .B(o[46]), .A(n4465), .Z(n4521) );
  XNOR U5703 ( .A(n4522), .B(n4521), .Z(n4554) );
  XOR U5704 ( .A(n4555), .B(n4554), .Z(n4556) );
  XNOR U5705 ( .A(n4557), .B(n4556), .Z(n4589) );
  NAND U5706 ( .A(x[234]), .B(y[1836]), .Z(n5378) );
  NANDN U5707 ( .A(n5378), .B(n4466), .Z(n4469) );
  NAND U5708 ( .A(n5039), .B(n4467), .Z(n4468) );
  NAND U5709 ( .A(n4469), .B(n4468), .Z(n4587) );
  AND U5710 ( .A(x[235]), .B(y[1832]), .Z(n4862) );
  NAND U5711 ( .A(n4862), .B(n4470), .Z(n4474) );
  NAND U5712 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U5713 ( .A(n4474), .B(n4473), .Z(n4586) );
  XOR U5714 ( .A(n4587), .B(n4586), .Z(n4588) );
  XOR U5715 ( .A(n4589), .B(n4588), .Z(n4580) );
  XOR U5716 ( .A(n4581), .B(n4580), .Z(n4582) );
  XOR U5717 ( .A(n4583), .B(n4582), .Z(n4575) );
  AND U5718 ( .A(x[238]), .B(y[1838]), .Z(n6261) );
  NAND U5719 ( .A(n6261), .B(n4520), .Z(n4478) );
  NAND U5720 ( .A(n4476), .B(n4475), .Z(n4477) );
  NAND U5721 ( .A(n4478), .B(n4477), .Z(n4549) );
  AND U5722 ( .A(x[232]), .B(y[1835]), .Z(n4479) );
  NAND U5723 ( .A(n4480), .B(n4479), .Z(n4483) );
  NAND U5724 ( .A(n4481), .B(n4756), .Z(n4482) );
  NAND U5725 ( .A(n4483), .B(n4482), .Z(n4548) );
  XOR U5726 ( .A(n4549), .B(n4548), .Z(n4551) );
  AND U5727 ( .A(y[1829]), .B(x[234]), .Z(n4485) );
  NAND U5728 ( .A(y[1835]), .B(x[228]), .Z(n4484) );
  XNOR U5729 ( .A(n4485), .B(n4484), .Z(n4528) );
  AND U5730 ( .A(x[231]), .B(y[1832]), .Z(n4527) );
  XNOR U5731 ( .A(n4528), .B(n4527), .Z(n4536) );
  NAND U5732 ( .A(x[230]), .B(y[1833]), .Z(n4533) );
  XOR U5733 ( .A(n4533), .B(n4534), .Z(n4535) );
  XOR U5734 ( .A(n4536), .B(n4535), .Z(n4571) );
  AND U5735 ( .A(y[1837]), .B(x[226]), .Z(n4487) );
  NAND U5736 ( .A(y[1830]), .B(x[233]), .Z(n4486) );
  XNOR U5737 ( .A(n4487), .B(n4486), .Z(n4539) );
  AND U5738 ( .A(x[227]), .B(y[1836]), .Z(n4540) );
  XOR U5739 ( .A(n4539), .B(n4540), .Z(n4569) );
  AND U5740 ( .A(y[1838]), .B(x[225]), .Z(n4489) );
  NAND U5741 ( .A(y[1831]), .B(x[232]), .Z(n4488) );
  XNOR U5742 ( .A(n4489), .B(n4488), .Z(n4517) );
  NAND U5743 ( .A(x[238]), .B(y[1825]), .Z(n4545) );
  XNOR U5744 ( .A(o[47]), .B(n4545), .Z(n4516) );
  XOR U5745 ( .A(n4517), .B(n4516), .Z(n4568) );
  XOR U5746 ( .A(n4569), .B(n4568), .Z(n4570) );
  XNOR U5747 ( .A(n4551), .B(n4550), .Z(n4593) );
  NAND U5748 ( .A(n4863), .B(n4490), .Z(n4494) );
  NAND U5749 ( .A(n4492), .B(n4491), .Z(n4493) );
  AND U5750 ( .A(n4494), .B(n4493), .Z(n4592) );
  XOR U5751 ( .A(n4593), .B(n4592), .Z(n4595) );
  NAND U5752 ( .A(n4496), .B(n4495), .Z(n4500) );
  NAND U5753 ( .A(n4498), .B(n4497), .Z(n4499) );
  AND U5754 ( .A(n4500), .B(n4499), .Z(n4594) );
  XOR U5755 ( .A(n4595), .B(n4594), .Z(n4574) );
  XOR U5756 ( .A(n4576), .B(n4577), .Z(n4601) );
  NAND U5757 ( .A(n4502), .B(n4501), .Z(n4506) );
  NAND U5758 ( .A(n4504), .B(n4503), .Z(n4505) );
  AND U5759 ( .A(n4506), .B(n4505), .Z(n4602) );
  XOR U5760 ( .A(n4601), .B(n4602), .Z(n4603) );
  XOR U5761 ( .A(n4604), .B(n4603), .Z(n4600) );
  XOR U5762 ( .A(n4598), .B(n4599), .Z(n4514) );
  XNOR U5763 ( .A(n4600), .B(n4514), .Z(N112) );
  AND U5764 ( .A(x[232]), .B(y[1838]), .Z(n4864) );
  NAND U5765 ( .A(n4864), .B(n4515), .Z(n4519) );
  NAND U5766 ( .A(n4517), .B(n4516), .Z(n4518) );
  AND U5767 ( .A(n4519), .B(n4518), .Z(n4676) );
  AND U5768 ( .A(x[239]), .B(y[1839]), .Z(n6698) );
  NAND U5769 ( .A(n6698), .B(n4520), .Z(n4524) );
  NAND U5770 ( .A(n4522), .B(n4521), .Z(n4523) );
  NAND U5771 ( .A(n4524), .B(n4523), .Z(n4675) );
  XNOR U5772 ( .A(n4676), .B(n4675), .Z(n4678) );
  AND U5773 ( .A(x[234]), .B(y[1835]), .Z(n4526) );
  NAND U5774 ( .A(n4526), .B(n4525), .Z(n4530) );
  NAND U5775 ( .A(n4528), .B(n4527), .Z(n4529) );
  NAND U5776 ( .A(n4530), .B(n4529), .Z(n4635) );
  AND U5777 ( .A(x[224]), .B(y[1840]), .Z(n4655) );
  NAND U5778 ( .A(x[240]), .B(y[1824]), .Z(n4656) );
  XNOR U5779 ( .A(n4655), .B(n4656), .Z(n4657) );
  NAND U5780 ( .A(x[239]), .B(y[1825]), .Z(n4645) );
  XOR U5781 ( .A(o[48]), .B(n4645), .Z(n4658) );
  XNOR U5782 ( .A(n4657), .B(n4658), .Z(n4634) );
  NAND U5783 ( .A(y[1833]), .B(x[231]), .Z(n4531) );
  XNOR U5784 ( .A(n4532), .B(n4531), .Z(n4650) );
  AND U5785 ( .A(x[234]), .B(y[1830]), .Z(n4649) );
  XOR U5786 ( .A(n4650), .B(n4649), .Z(n4633) );
  XOR U5787 ( .A(n4634), .B(n4633), .Z(n4636) );
  XOR U5788 ( .A(n4635), .B(n4636), .Z(n4677) );
  XNOR U5789 ( .A(n4678), .B(n4677), .Z(n4630) );
  IV U5790 ( .A(n4533), .Z(n4648) );
  NANDN U5791 ( .A(n4648), .B(n4534), .Z(n4538) );
  NAND U5792 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U5793 ( .A(n4538), .B(n4537), .Z(n4628) );
  AND U5794 ( .A(x[233]), .B(y[1837]), .Z(n5358) );
  NAND U5795 ( .A(n5358), .B(n4948), .Z(n4542) );
  NAND U5796 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U5797 ( .A(n4542), .B(n4541), .Z(n4665) );
  AND U5798 ( .A(y[1839]), .B(x[225]), .Z(n4544) );
  NAND U5799 ( .A(y[1832]), .B(x[232]), .Z(n4543) );
  XNOR U5800 ( .A(n4544), .B(n4543), .Z(n4654) );
  ANDN U5801 ( .B(o[47]), .A(n4545), .Z(n4653) );
  XOR U5802 ( .A(n4654), .B(n4653), .Z(n4664) );
  NAND U5803 ( .A(y[1826]), .B(x[238]), .Z(n4546) );
  XNOR U5804 ( .A(n4547), .B(n4546), .Z(n4687) );
  NAND U5805 ( .A(x[228]), .B(y[1836]), .Z(n4688) );
  XNOR U5806 ( .A(n4687), .B(n4688), .Z(n4663) );
  XOR U5807 ( .A(n4664), .B(n4663), .Z(n4666) );
  XNOR U5808 ( .A(n4665), .B(n4666), .Z(n4627) );
  XOR U5809 ( .A(n4628), .B(n4627), .Z(n4629) );
  XOR U5810 ( .A(n4630), .B(n4629), .Z(n4669) );
  NAND U5811 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U5812 ( .A(n4551), .B(n4550), .Z(n4552) );
  AND U5813 ( .A(n4553), .B(n4552), .Z(n4670) );
  XOR U5814 ( .A(n4669), .B(n4670), .Z(n4672) );
  NAND U5815 ( .A(n4555), .B(n4554), .Z(n4559) );
  NAND U5816 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U5817 ( .A(n4559), .B(n4558), .Z(n4701) );
  AND U5818 ( .A(x[237]), .B(y[1828]), .Z(n4698) );
  NAND U5819 ( .A(n5186), .B(n4698), .Z(n4563) );
  NAND U5820 ( .A(n4561), .B(n4560), .Z(n4562) );
  AND U5821 ( .A(n4563), .B(n4562), .Z(n4684) );
  AND U5822 ( .A(y[1838]), .B(x[226]), .Z(n4565) );
  NAND U5823 ( .A(y[1831]), .B(x[233]), .Z(n4564) );
  XNOR U5824 ( .A(n4565), .B(n4564), .Z(n4691) );
  NAND U5825 ( .A(x[227]), .B(y[1837]), .Z(n4692) );
  XNOR U5826 ( .A(n4691), .B(n4692), .Z(n4681) );
  AND U5827 ( .A(x[236]), .B(y[1828]), .Z(n5347) );
  AND U5828 ( .A(y[1835]), .B(x[229]), .Z(n4567) );
  NAND U5829 ( .A(y[1827]), .B(x[237]), .Z(n4566) );
  XOR U5830 ( .A(n4567), .B(n4566), .Z(n4640) );
  XOR U5831 ( .A(n5347), .B(n4640), .Z(n4682) );
  XNOR U5832 ( .A(n4681), .B(n4682), .Z(n4683) );
  XOR U5833 ( .A(n4684), .B(n4683), .Z(n4699) );
  NAND U5834 ( .A(n4569), .B(n4568), .Z(n4573) );
  NANDN U5835 ( .A(n4571), .B(n4570), .Z(n4572) );
  AND U5836 ( .A(n4573), .B(n4572), .Z(n4700) );
  XOR U5837 ( .A(n4699), .B(n4700), .Z(n4702) );
  XOR U5838 ( .A(n4701), .B(n4702), .Z(n4671) );
  XOR U5839 ( .A(n4672), .B(n4671), .Z(n4609) );
  NANDN U5840 ( .A(n4575), .B(n4574), .Z(n4579) );
  NANDN U5841 ( .A(n4577), .B(n4576), .Z(n4578) );
  AND U5842 ( .A(n4579), .B(n4578), .Z(n4608) );
  NAND U5843 ( .A(n4581), .B(n4580), .Z(n4585) );
  NAND U5844 ( .A(n4583), .B(n4582), .Z(n4584) );
  NAND U5845 ( .A(n4585), .B(n4584), .Z(n4624) );
  NAND U5846 ( .A(n4587), .B(n4586), .Z(n4591) );
  NAND U5847 ( .A(n4589), .B(n4588), .Z(n4590) );
  NAND U5848 ( .A(n4591), .B(n4590), .Z(n4622) );
  NAND U5849 ( .A(n4593), .B(n4592), .Z(n4597) );
  NAND U5850 ( .A(n4595), .B(n4594), .Z(n4596) );
  AND U5851 ( .A(n4597), .B(n4596), .Z(n4621) );
  XOR U5852 ( .A(n4622), .B(n4621), .Z(n4623) );
  XNOR U5853 ( .A(n4624), .B(n4623), .Z(n4611) );
  XNOR U5854 ( .A(n4610), .B(n4611), .Z(n4617) );
  NAND U5855 ( .A(n4602), .B(n4601), .Z(n4606) );
  NANDN U5856 ( .A(n4604), .B(n4603), .Z(n4605) );
  AND U5857 ( .A(n4606), .B(n4605), .Z(n4616) );
  IV U5858 ( .A(n4616), .Z(n4614) );
  XOR U5859 ( .A(n4615), .B(n4614), .Z(n4607) );
  XNOR U5860 ( .A(n4617), .B(n4607), .Z(N113) );
  NANDN U5861 ( .A(n4609), .B(n4608), .Z(n4613) );
  NANDN U5862 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5863 ( .A(n4613), .B(n4612), .Z(n4802) );
  NANDN U5864 ( .A(n4614), .B(n4615), .Z(n4620) );
  NOR U5865 ( .A(n4616), .B(n4615), .Z(n4618) );
  OR U5866 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U5867 ( .A(n4620), .B(n4619), .Z(n4803) );
  NAND U5868 ( .A(n4622), .B(n4621), .Z(n4626) );
  NAND U5869 ( .A(n4624), .B(n4623), .Z(n4625) );
  NAND U5870 ( .A(n4626), .B(n4625), .Z(n4799) );
  NAND U5871 ( .A(n4628), .B(n4627), .Z(n4632) );
  NAND U5872 ( .A(n4630), .B(n4629), .Z(n4631) );
  NAND U5873 ( .A(n4632), .B(n4631), .Z(n4714) );
  NAND U5874 ( .A(n4634), .B(n4633), .Z(n4638) );
  NAND U5875 ( .A(n4636), .B(n4635), .Z(n4637) );
  AND U5876 ( .A(n4638), .B(n4637), .Z(n4793) );
  AND U5877 ( .A(x[237]), .B(y[1835]), .Z(n5651) );
  NAND U5878 ( .A(n5651), .B(n4639), .Z(n4642) );
  NANDN U5879 ( .A(n4640), .B(n5347), .Z(n4641) );
  AND U5880 ( .A(n4642), .B(n4641), .Z(n4745) );
  AND U5881 ( .A(y[1840]), .B(x[225]), .Z(n4644) );
  NAND U5882 ( .A(y[1832]), .B(x[233]), .Z(n4643) );
  XNOR U5883 ( .A(n4644), .B(n4643), .Z(n4762) );
  ANDN U5884 ( .B(o[48]), .A(n4645), .Z(n4761) );
  XOR U5885 ( .A(n4762), .B(n4761), .Z(n4743) );
  AND U5886 ( .A(y[1826]), .B(x[239]), .Z(n4647) );
  NAND U5887 ( .A(y[1829]), .B(x[236]), .Z(n4646) );
  XNOR U5888 ( .A(n4647), .B(n4646), .Z(n4719) );
  AND U5889 ( .A(x[238]), .B(y[1827]), .Z(n4718) );
  XOR U5890 ( .A(n4719), .B(n4718), .Z(n4742) );
  XOR U5891 ( .A(n4743), .B(n4742), .Z(n4744) );
  XNOR U5892 ( .A(n4745), .B(n4744), .Z(n4790) );
  NAND U5893 ( .A(x[231]), .B(y[1834]), .Z(n4773) );
  NANDN U5894 ( .A(n4773), .B(n4648), .Z(n4652) );
  NAND U5895 ( .A(n4650), .B(n4649), .Z(n4651) );
  AND U5896 ( .A(n4652), .B(n4651), .Z(n4751) );
  NAND U5897 ( .A(x[232]), .B(y[1839]), .Z(n5441) );
  AND U5898 ( .A(x[225]), .B(y[1832]), .Z(n4842) );
  XNOR U5899 ( .A(n4751), .B(n4750), .Z(n4752) );
  NANDN U5900 ( .A(n4656), .B(n4655), .Z(n4660) );
  NANDN U5901 ( .A(n4658), .B(n4657), .Z(n4659) );
  AND U5902 ( .A(n4660), .B(n4659), .Z(n4749) );
  AND U5903 ( .A(x[224]), .B(y[1841]), .Z(n4733) );
  AND U5904 ( .A(x[241]), .B(y[1824]), .Z(n4732) );
  XOR U5905 ( .A(n4733), .B(n4732), .Z(n4735) );
  AND U5906 ( .A(x[240]), .B(y[1825]), .Z(n4729) );
  XOR U5907 ( .A(n4729), .B(o[49]), .Z(n4734) );
  XOR U5908 ( .A(n4735), .B(n4734), .Z(n4747) );
  AND U5909 ( .A(y[1839]), .B(x[226]), .Z(n4662) );
  NAND U5910 ( .A(y[1831]), .B(x[234]), .Z(n4661) );
  XNOR U5911 ( .A(n4662), .B(n4661), .Z(n4766) );
  AND U5912 ( .A(x[227]), .B(y[1838]), .Z(n4767) );
  XOR U5913 ( .A(n4766), .B(n4767), .Z(n4746) );
  XOR U5914 ( .A(n4747), .B(n4746), .Z(n4748) );
  XOR U5915 ( .A(n4749), .B(n4748), .Z(n4753) );
  XOR U5916 ( .A(n4752), .B(n4753), .Z(n4791) );
  XNOR U5917 ( .A(n4790), .B(n4791), .Z(n4792) );
  XOR U5918 ( .A(n4793), .B(n4792), .Z(n4712) );
  NAND U5919 ( .A(n4664), .B(n4663), .Z(n4668) );
  NAND U5920 ( .A(n4666), .B(n4665), .Z(n4667) );
  AND U5921 ( .A(n4668), .B(n4667), .Z(n4713) );
  XNOR U5922 ( .A(n4712), .B(n4713), .Z(n4715) );
  NAND U5923 ( .A(n4670), .B(n4669), .Z(n4674) );
  NAND U5924 ( .A(n4672), .B(n4671), .Z(n4673) );
  NAND U5925 ( .A(n4674), .B(n4673), .Z(n4708) );
  NANDN U5926 ( .A(n4676), .B(n4675), .Z(n4680) );
  NAND U5927 ( .A(n4678), .B(n4677), .Z(n4679) );
  AND U5928 ( .A(n4680), .B(n4679), .Z(n4787) );
  NANDN U5929 ( .A(n4682), .B(n4681), .Z(n4686) );
  NANDN U5930 ( .A(n4684), .B(n4683), .Z(n4685) );
  AND U5931 ( .A(n4686), .B(n4685), .Z(n4785) );
  NAND U5932 ( .A(x[238]), .B(y[1829]), .Z(n4982) );
  NANDN U5933 ( .A(n4982), .B(n5186), .Z(n4690) );
  NANDN U5934 ( .A(n4688), .B(n4687), .Z(n4689) );
  AND U5935 ( .A(n4690), .B(n4689), .Z(n4779) );
  AND U5936 ( .A(x[233]), .B(y[1838]), .Z(n5632) );
  NAND U5937 ( .A(n4765), .B(n5632), .Z(n4694) );
  NANDN U5938 ( .A(n4692), .B(n4691), .Z(n4693) );
  NAND U5939 ( .A(n4694), .B(n4693), .Z(n4778) );
  XNOR U5940 ( .A(n4779), .B(n4778), .Z(n4780) );
  AND U5941 ( .A(x[229]), .B(y[1836]), .Z(n4824) );
  NAND U5942 ( .A(y[1833]), .B(x[232]), .Z(n4695) );
  XNOR U5943 ( .A(n4824), .B(n4695), .Z(n4757) );
  XOR U5944 ( .A(n4757), .B(n4696), .Z(n4772) );
  XNOR U5945 ( .A(n4772), .B(n4773), .Z(n4774) );
  NAND U5946 ( .A(y[1837]), .B(x[228]), .Z(n4697) );
  XNOR U5947 ( .A(n4698), .B(n4697), .Z(n4723) );
  NAND U5948 ( .A(x[235]), .B(y[1830]), .Z(n4724) );
  XOR U5949 ( .A(n4723), .B(n4724), .Z(n4775) );
  XOR U5950 ( .A(n4774), .B(n4775), .Z(n4781) );
  XNOR U5951 ( .A(n4780), .B(n4781), .Z(n4784) );
  XNOR U5952 ( .A(n4785), .B(n4784), .Z(n4786) );
  XOR U5953 ( .A(n4787), .B(n4786), .Z(n4707) );
  NAND U5954 ( .A(n4700), .B(n4699), .Z(n4704) );
  NAND U5955 ( .A(n4702), .B(n4701), .Z(n4703) );
  NAND U5956 ( .A(n4704), .B(n4703), .Z(n4706) );
  XNOR U5957 ( .A(n4707), .B(n4706), .Z(n4709) );
  XOR U5958 ( .A(n4708), .B(n4709), .Z(n4796) );
  XOR U5959 ( .A(n4797), .B(n4796), .Z(n4798) );
  XOR U5960 ( .A(n4799), .B(n4798), .Z(n4804) );
  XNOR U5961 ( .A(n4803), .B(n4804), .Z(n4705) );
  XOR U5962 ( .A(n4802), .B(n4705), .Z(N114) );
  NAND U5963 ( .A(n4707), .B(n4706), .Z(n4711) );
  NANDN U5964 ( .A(n4709), .B(n4708), .Z(n4710) );
  AND U5965 ( .A(n4711), .B(n4710), .Z(n4911) );
  NAND U5966 ( .A(n4713), .B(n4712), .Z(n4717) );
  NANDN U5967 ( .A(n4715), .B(n4714), .Z(n4716) );
  AND U5968 ( .A(n4717), .B(n4716), .Z(n4909) );
  AND U5969 ( .A(x[236]), .B(y[1826]), .Z(n5045) );
  AND U5970 ( .A(x[239]), .B(y[1829]), .Z(n4956) );
  NAND U5971 ( .A(n5045), .B(n4956), .Z(n4721) );
  NAND U5972 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U5973 ( .A(n4721), .B(n4720), .Z(n4890) );
  NAND U5974 ( .A(n5987), .B(n4722), .Z(n4726) );
  NANDN U5975 ( .A(n4724), .B(n4723), .Z(n4725) );
  NAND U5976 ( .A(n4726), .B(n4725), .Z(n4881) );
  AND U5977 ( .A(y[1841]), .B(x[225]), .Z(n4728) );
  NAND U5978 ( .A(y[1832]), .B(x[234]), .Z(n4727) );
  XNOR U5979 ( .A(n4728), .B(n4727), .Z(n4843) );
  AND U5980 ( .A(n4729), .B(o[49]), .Z(n4844) );
  XOR U5981 ( .A(n4843), .B(n4844), .Z(n4879) );
  AND U5982 ( .A(y[1827]), .B(x[239]), .Z(n4731) );
  NAND U5983 ( .A(y[1833]), .B(x[233]), .Z(n4730) );
  XNOR U5984 ( .A(n4731), .B(n4730), .Z(n4834) );
  AND U5985 ( .A(x[238]), .B(y[1828]), .Z(n4835) );
  XOR U5986 ( .A(n4834), .B(n4835), .Z(n4878) );
  XOR U5987 ( .A(n4879), .B(n4878), .Z(n4880) );
  XOR U5988 ( .A(n4881), .B(n4880), .Z(n4891) );
  XOR U5989 ( .A(n4890), .B(n4891), .Z(n4893) );
  NAND U5990 ( .A(n4733), .B(n4732), .Z(n4737) );
  NAND U5991 ( .A(n4735), .B(n4734), .Z(n4736) );
  NAND U5992 ( .A(n4737), .B(n4736), .Z(n4902) );
  AND U5993 ( .A(y[1826]), .B(x[240]), .Z(n4739) );
  NAND U5994 ( .A(y[1831]), .B(x[235]), .Z(n4738) );
  XNOR U5995 ( .A(n4739), .B(n4738), .Z(n4830) );
  AND U5996 ( .A(x[226]), .B(y[1840]), .Z(n4831) );
  XOR U5997 ( .A(n4830), .B(n4831), .Z(n4903) );
  XOR U5998 ( .A(n4902), .B(n4903), .Z(n4905) );
  AND U5999 ( .A(y[1837]), .B(x[229]), .Z(n4964) );
  NAND U6000 ( .A(y[1836]), .B(x[230]), .Z(n4740) );
  XNOR U6001 ( .A(n4964), .B(n4740), .Z(n4827) );
  NAND U6002 ( .A(y[1838]), .B(x[228]), .Z(n4741) );
  XNOR U6003 ( .A(n5637), .B(n4741), .Z(n4865) );
  AND U6004 ( .A(x[231]), .B(y[1835]), .Z(n4866) );
  XOR U6005 ( .A(n4865), .B(n4866), .Z(n4826) );
  XOR U6006 ( .A(n4827), .B(n4826), .Z(n4904) );
  XOR U6007 ( .A(n4905), .B(n4904), .Z(n4892) );
  XOR U6008 ( .A(n4893), .B(n4892), .Z(n4813) );
  XOR U6009 ( .A(n4885), .B(n4884), .Z(n4887) );
  NANDN U6010 ( .A(n4751), .B(n4750), .Z(n4755) );
  NANDN U6011 ( .A(n4753), .B(n4752), .Z(n4754) );
  AND U6012 ( .A(n4755), .B(n4754), .Z(n4886) );
  XOR U6013 ( .A(n4887), .B(n4886), .Z(n4812) );
  XNOR U6014 ( .A(n4813), .B(n4812), .Z(n4815) );
  AND U6015 ( .A(x[232]), .B(y[1836]), .Z(n5085) );
  NAND U6016 ( .A(n5085), .B(n4756), .Z(n4760) );
  NANDN U6017 ( .A(n4758), .B(n4757), .Z(n4759) );
  NAND U6018 ( .A(n4760), .B(n4759), .Z(n4897) );
  AND U6019 ( .A(x[233]), .B(y[1840]), .Z(n5730) );
  NAND U6020 ( .A(n5730), .B(n4842), .Z(n4764) );
  NAND U6021 ( .A(n4762), .B(n4761), .Z(n4763) );
  NAND U6022 ( .A(n4764), .B(n4763), .Z(n4896) );
  XOR U6023 ( .A(n4897), .B(n4896), .Z(n4899) );
  AND U6024 ( .A(x[234]), .B(y[1839]), .Z(n5660) );
  IV U6025 ( .A(n5660), .Z(n5729) );
  NANDN U6026 ( .A(n5729), .B(n4765), .Z(n4769) );
  NAND U6027 ( .A(n4767), .B(n4766), .Z(n4768) );
  AND U6028 ( .A(n4769), .B(n4768), .Z(n4875) );
  AND U6029 ( .A(x[224]), .B(y[1842]), .Z(n4847) );
  AND U6030 ( .A(x[242]), .B(y[1824]), .Z(n4848) );
  XOR U6031 ( .A(n4847), .B(n4848), .Z(n4850) );
  AND U6032 ( .A(x[241]), .B(y[1825]), .Z(n4869) );
  XOR U6033 ( .A(o[50]), .B(n4869), .Z(n4849) );
  XOR U6034 ( .A(n4850), .B(n4849), .Z(n4873) );
  AND U6035 ( .A(y[1829]), .B(x[237]), .Z(n4771) );
  NAND U6036 ( .A(y[1839]), .B(x[227]), .Z(n4770) );
  XNOR U6037 ( .A(n4771), .B(n4770), .Z(n4855) );
  AND U6038 ( .A(x[236]), .B(y[1830]), .Z(n4856) );
  XOR U6039 ( .A(n4855), .B(n4856), .Z(n4872) );
  XOR U6040 ( .A(n4873), .B(n4872), .Z(n4874) );
  XNOR U6041 ( .A(n4899), .B(n4898), .Z(n4819) );
  NANDN U6042 ( .A(n4773), .B(n4772), .Z(n4777) );
  NANDN U6043 ( .A(n4775), .B(n4774), .Z(n4776) );
  AND U6044 ( .A(n4777), .B(n4776), .Z(n4818) );
  XOR U6045 ( .A(n4819), .B(n4818), .Z(n4820) );
  NANDN U6046 ( .A(n4779), .B(n4778), .Z(n4783) );
  NANDN U6047 ( .A(n4781), .B(n4780), .Z(n4782) );
  AND U6048 ( .A(n4783), .B(n4782), .Z(n4821) );
  XOR U6049 ( .A(n4820), .B(n4821), .Z(n4814) );
  XOR U6050 ( .A(n4815), .B(n4814), .Z(n4808) );
  NANDN U6051 ( .A(n4785), .B(n4784), .Z(n4789) );
  NANDN U6052 ( .A(n4787), .B(n4786), .Z(n4788) );
  AND U6053 ( .A(n4789), .B(n4788), .Z(n4807) );
  NANDN U6054 ( .A(n4791), .B(n4790), .Z(n4795) );
  NANDN U6055 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U6056 ( .A(n4795), .B(n4794), .Z(n4806) );
  XOR U6057 ( .A(n4807), .B(n4806), .Z(n4809) );
  XOR U6058 ( .A(n4808), .B(n4809), .Z(n4908) );
  XOR U6059 ( .A(n4909), .B(n4908), .Z(n4910) );
  XNOR U6060 ( .A(n4911), .B(n4910), .Z(n4916) );
  NAND U6061 ( .A(n4797), .B(n4796), .Z(n4801) );
  NAND U6062 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U6063 ( .A(n4801), .B(n4800), .Z(n4915) );
  XOR U6064 ( .A(n4915), .B(n4914), .Z(n4805) );
  XNOR U6065 ( .A(n4916), .B(n4805), .Z(N115) );
  NANDN U6066 ( .A(n4807), .B(n4806), .Z(n4811) );
  OR U6067 ( .A(n4809), .B(n4808), .Z(n4810) );
  AND U6068 ( .A(n4811), .B(n4810), .Z(n4924) );
  NANDN U6069 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U6070 ( .A(n4815), .B(n4814), .Z(n4816) );
  AND U6071 ( .A(n4817), .B(n4816), .Z(n4922) );
  NAND U6072 ( .A(n4819), .B(n4818), .Z(n4823) );
  NAND U6073 ( .A(n4821), .B(n4820), .Z(n4822) );
  AND U6074 ( .A(n4823), .B(n4822), .Z(n4928) );
  AND U6075 ( .A(x[230]), .B(y[1837]), .Z(n4825) );
  NAND U6076 ( .A(n4825), .B(n4824), .Z(n4829) );
  NAND U6077 ( .A(n4827), .B(n4826), .Z(n4828) );
  AND U6078 ( .A(n4829), .B(n4828), .Z(n5017) );
  AND U6079 ( .A(x[240]), .B(y[1831]), .Z(n5363) );
  NAND U6080 ( .A(n5363), .B(n5186), .Z(n4833) );
  NAND U6081 ( .A(n4831), .B(n4830), .Z(n4832) );
  AND U6082 ( .A(n4833), .B(n4832), .Z(n5015) );
  AND U6083 ( .A(x[239]), .B(y[1833]), .Z(n5665) );
  NAND U6084 ( .A(n5665), .B(n4943), .Z(n4837) );
  NAND U6085 ( .A(n4835), .B(n4834), .Z(n4836) );
  NAND U6086 ( .A(n4837), .B(n4836), .Z(n4934) );
  AND U6087 ( .A(y[1842]), .B(x[225]), .Z(n4839) );
  NAND U6088 ( .A(y[1835]), .B(x[232]), .Z(n4838) );
  XNOR U6089 ( .A(n4839), .B(n4838), .Z(n4981) );
  AND U6090 ( .A(y[1830]), .B(x[237]), .Z(n4841) );
  NAND U6091 ( .A(y[1841]), .B(x[226]), .Z(n4840) );
  XNOR U6092 ( .A(n4841), .B(n4840), .Z(n4949) );
  XOR U6093 ( .A(n4932), .B(n4931), .Z(n4933) );
  XOR U6094 ( .A(n4934), .B(n4933), .Z(n5014) );
  AND U6095 ( .A(x[234]), .B(y[1841]), .Z(n6075) );
  NAND U6096 ( .A(n6075), .B(n4842), .Z(n4846) );
  NAND U6097 ( .A(n4844), .B(n4843), .Z(n4845) );
  NAND U6098 ( .A(n4846), .B(n4845), .Z(n4993) );
  NAND U6099 ( .A(n4848), .B(n4847), .Z(n4852) );
  NAND U6100 ( .A(n4850), .B(n4849), .Z(n4851) );
  NAND U6101 ( .A(n4852), .B(n4851), .Z(n4991) );
  AND U6102 ( .A(y[1827]), .B(x[240]), .Z(n5603) );
  NAND U6103 ( .A(y[1834]), .B(x[233]), .Z(n4853) );
  XNOR U6104 ( .A(n5603), .B(n4853), .Z(n4944) );
  AND U6105 ( .A(x[239]), .B(y[1828]), .Z(n4945) );
  XOR U6106 ( .A(n4944), .B(n4945), .Z(n4990) );
  XOR U6107 ( .A(n4991), .B(n4990), .Z(n4992) );
  XNOR U6108 ( .A(n4993), .B(n4992), .Z(n5010) );
  AND U6109 ( .A(x[237]), .B(y[1839]), .Z(n6289) );
  NANDN U6110 ( .A(n4854), .B(n6289), .Z(n4858) );
  NAND U6111 ( .A(n4856), .B(n4855), .Z(n4857) );
  NAND U6112 ( .A(n4858), .B(n4857), .Z(n4999) );
  AND U6113 ( .A(y[1833]), .B(x[234]), .Z(n4860) );
  NAND U6114 ( .A(y[1826]), .B(x[241]), .Z(n4859) );
  XNOR U6115 ( .A(n4860), .B(n4859), .Z(n4987) );
  AND U6116 ( .A(x[242]), .B(y[1825]), .Z(n4963) );
  XOR U6117 ( .A(o[51]), .B(n4963), .Z(n4986) );
  XOR U6118 ( .A(n4987), .B(n4986), .Z(n4997) );
  NAND U6119 ( .A(y[1840]), .B(x[227]), .Z(n4861) );
  XNOR U6120 ( .A(n4862), .B(n4861), .Z(n4957) );
  XOR U6121 ( .A(n4997), .B(n4996), .Z(n4998) );
  XNOR U6122 ( .A(n4999), .B(n4998), .Z(n5009) );
  NAND U6123 ( .A(n4864), .B(n4863), .Z(n4868) );
  NAND U6124 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U6125 ( .A(n4868), .B(n4867), .Z(n4940) );
  AND U6126 ( .A(x[224]), .B(y[1843]), .Z(n4968) );
  AND U6127 ( .A(x[243]), .B(y[1824]), .Z(n4969) );
  XOR U6128 ( .A(n4968), .B(n4969), .Z(n4971) );
  AND U6129 ( .A(o[50]), .B(n4869), .Z(n4970) );
  XOR U6130 ( .A(n4971), .B(n4970), .Z(n4938) );
  AND U6131 ( .A(x[228]), .B(y[1839]), .Z(n5099) );
  AND U6132 ( .A(y[1838]), .B(x[229]), .Z(n4871) );
  NAND U6133 ( .A(y[1837]), .B(x[230]), .Z(n4870) );
  XNOR U6134 ( .A(n4871), .B(n4870), .Z(n4965) );
  XOR U6135 ( .A(n5099), .B(n4965), .Z(n4937) );
  XOR U6136 ( .A(n4938), .B(n4937), .Z(n4939) );
  XOR U6137 ( .A(n4940), .B(n4939), .Z(n5008) );
  XOR U6138 ( .A(n5009), .B(n5008), .Z(n5011) );
  XNOR U6139 ( .A(n5010), .B(n5011), .Z(n5004) );
  NAND U6140 ( .A(n4873), .B(n4872), .Z(n4877) );
  NANDN U6141 ( .A(n4875), .B(n4874), .Z(n4876) );
  AND U6142 ( .A(n4877), .B(n4876), .Z(n5003) );
  NAND U6143 ( .A(n4879), .B(n4878), .Z(n4883) );
  NAND U6144 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U6145 ( .A(n4883), .B(n4882), .Z(n5002) );
  XNOR U6146 ( .A(n5004), .B(n5005), .Z(n4925) );
  XOR U6147 ( .A(n4926), .B(n4925), .Z(n4927) );
  NAND U6148 ( .A(n4885), .B(n4884), .Z(n4889) );
  NAND U6149 ( .A(n4887), .B(n4886), .Z(n4888) );
  AND U6150 ( .A(n4889), .B(n4888), .Z(n5026) );
  NAND U6151 ( .A(n4891), .B(n4890), .Z(n4895) );
  NAND U6152 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U6153 ( .A(n4895), .B(n4894), .Z(n5022) );
  NAND U6154 ( .A(n4897), .B(n4896), .Z(n4901) );
  NAND U6155 ( .A(n4899), .B(n4898), .Z(n4900) );
  NAND U6156 ( .A(n4901), .B(n4900), .Z(n5021) );
  NAND U6157 ( .A(n4903), .B(n4902), .Z(n4907) );
  NAND U6158 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U6159 ( .A(n4907), .B(n4906), .Z(n5020) );
  XNOR U6160 ( .A(n5021), .B(n5020), .Z(n5023) );
  XNOR U6161 ( .A(n5026), .B(n5027), .Z(n5028) );
  XOR U6162 ( .A(n4922), .B(n4921), .Z(n4923) );
  XNOR U6163 ( .A(n4924), .B(n4923), .Z(n4920) );
  NAND U6164 ( .A(n4909), .B(n4908), .Z(n4913) );
  NAND U6165 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U6166 ( .A(n4913), .B(n4912), .Z(n4919) );
  XNOR U6167 ( .A(n4919), .B(n4918), .Z(n4917) );
  XNOR U6168 ( .A(n4920), .B(n4917), .Z(N116) );
  NAND U6169 ( .A(n4926), .B(n4925), .Z(n4930) );
  NANDN U6170 ( .A(n4928), .B(n4927), .Z(n4929) );
  AND U6171 ( .A(n4930), .B(n4929), .Z(n5137) );
  NAND U6172 ( .A(n4932), .B(n4931), .Z(n4936) );
  NAND U6173 ( .A(n4934), .B(n4933), .Z(n4935) );
  NAND U6174 ( .A(n4936), .B(n4935), .Z(n5034) );
  NAND U6175 ( .A(n4938), .B(n4937), .Z(n4942) );
  NANDN U6176 ( .A(n4940), .B(n4939), .Z(n4941) );
  NAND U6177 ( .A(n4942), .B(n4941), .Z(n5033) );
  XOR U6178 ( .A(n5034), .B(n5033), .Z(n5036) );
  AND U6179 ( .A(x[240]), .B(y[1834]), .Z(n5900) );
  NAND U6180 ( .A(n5900), .B(n4943), .Z(n4947) );
  NAND U6181 ( .A(n4945), .B(n4944), .Z(n4946) );
  NAND U6182 ( .A(n4947), .B(n4946), .Z(n5074) );
  AND U6183 ( .A(x[237]), .B(y[1841]), .Z(n6514) );
  NAND U6184 ( .A(n6514), .B(n4948), .Z(n4952) );
  NANDN U6185 ( .A(n4950), .B(n4949), .Z(n4951) );
  NAND U6186 ( .A(n4952), .B(n4951), .Z(n5119) );
  AND U6187 ( .A(y[1828]), .B(x[240]), .Z(n4954) );
  NAND U6188 ( .A(y[1834]), .B(x[234]), .Z(n4953) );
  XNOR U6189 ( .A(n4954), .B(n4953), .Z(n5080) );
  AND U6190 ( .A(x[226]), .B(y[1842]), .Z(n5081) );
  XOR U6191 ( .A(n5080), .B(n5081), .Z(n5117) );
  NAND U6192 ( .A(y[1835]), .B(x[233]), .Z(n4955) );
  XNOR U6193 ( .A(n4956), .B(n4955), .Z(n5040) );
  AND U6194 ( .A(x[238]), .B(y[1830]), .Z(n5041) );
  XOR U6195 ( .A(n5040), .B(n5041), .Z(n5116) );
  XOR U6196 ( .A(n5117), .B(n5116), .Z(n5118) );
  XOR U6197 ( .A(n5119), .B(n5118), .Z(n5073) );
  XOR U6198 ( .A(n5074), .B(n5073), .Z(n5076) );
  AND U6199 ( .A(x[235]), .B(y[1840]), .Z(n6077) );
  IV U6200 ( .A(n6077), .Z(n5948) );
  NANDN U6201 ( .A(n5948), .B(n5213), .Z(n4960) );
  NANDN U6202 ( .A(n4958), .B(n4957), .Z(n4959) );
  NAND U6203 ( .A(n4960), .B(n4959), .Z(n5125) );
  AND U6204 ( .A(y[1833]), .B(x[235]), .Z(n4962) );
  NAND U6205 ( .A(y[1843]), .B(x[225]), .Z(n4961) );
  XNOR U6206 ( .A(n4962), .B(n4961), .Z(n5052) );
  AND U6207 ( .A(x[243]), .B(y[1825]), .Z(n5044) );
  XOR U6208 ( .A(o[52]), .B(n5044), .Z(n5051) );
  XOR U6209 ( .A(n5052), .B(n5051), .Z(n5123) );
  AND U6210 ( .A(x[224]), .B(y[1844]), .Z(n5104) );
  AND U6211 ( .A(x[244]), .B(y[1824]), .Z(n5105) );
  XOR U6212 ( .A(n5104), .B(n5105), .Z(n5107) );
  AND U6213 ( .A(o[51]), .B(n4963), .Z(n5106) );
  XOR U6214 ( .A(n5107), .B(n5106), .Z(n5122) );
  XOR U6215 ( .A(n5123), .B(n5122), .Z(n5124) );
  XOR U6216 ( .A(n5125), .B(n5124), .Z(n5075) );
  XOR U6217 ( .A(n5076), .B(n5075), .Z(n5035) );
  XNOR U6218 ( .A(n5036), .B(n5035), .Z(n5131) );
  NAND U6219 ( .A(x[230]), .B(y[1838]), .Z(n5056) );
  NANDN U6220 ( .A(n5056), .B(n4964), .Z(n4967) );
  NAND U6221 ( .A(n4965), .B(n5099), .Z(n4966) );
  NAND U6222 ( .A(n4967), .B(n4966), .Z(n5064) );
  NAND U6223 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U6224 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U6225 ( .A(n4973), .B(n4972), .Z(n5062) );
  AND U6226 ( .A(y[1826]), .B(x[242]), .Z(n4975) );
  NAND U6227 ( .A(y[1832]), .B(x[236]), .Z(n4974) );
  XNOR U6228 ( .A(n4975), .B(n4974), .Z(n5046) );
  AND U6229 ( .A(x[241]), .B(y[1827]), .Z(n5047) );
  XOR U6230 ( .A(n5046), .B(n5047), .Z(n5061) );
  XOR U6231 ( .A(n5062), .B(n5061), .Z(n5063) );
  XNOR U6232 ( .A(n5064), .B(n5063), .Z(n5068) );
  AND U6233 ( .A(y[1831]), .B(x[237]), .Z(n4977) );
  NAND U6234 ( .A(y[1841]), .B(x[227]), .Z(n4976) );
  XNOR U6235 ( .A(n4977), .B(n4976), .Z(n5086) );
  XNOR U6236 ( .A(n5086), .B(n5085), .Z(n5058) );
  AND U6237 ( .A(y[1839]), .B(x[229]), .Z(n4979) );
  NAND U6238 ( .A(y[1840]), .B(x[228]), .Z(n4978) );
  XNOR U6239 ( .A(n4979), .B(n4978), .Z(n5101) );
  AND U6240 ( .A(x[231]), .B(y[1837]), .Z(n5100) );
  XNOR U6241 ( .A(n5101), .B(n5100), .Z(n5055) );
  XOR U6242 ( .A(n5056), .B(n5055), .Z(n5057) );
  XNOR U6243 ( .A(n5058), .B(n5057), .Z(n5112) );
  AND U6244 ( .A(x[232]), .B(y[1842]), .Z(n6241) );
  AND U6245 ( .A(x[225]), .B(y[1835]), .Z(n4980) );
  NAND U6246 ( .A(n6241), .B(n4980), .Z(n4984) );
  NANDN U6247 ( .A(n4982), .B(n4981), .Z(n4983) );
  NAND U6248 ( .A(n4984), .B(n4983), .Z(n5111) );
  NAND U6249 ( .A(x[241]), .B(y[1833]), .Z(n5908) );
  NANDN U6250 ( .A(n5908), .B(n4985), .Z(n4989) );
  NAND U6251 ( .A(n4987), .B(n4986), .Z(n4988) );
  NAND U6252 ( .A(n4989), .B(n4988), .Z(n5110) );
  XOR U6253 ( .A(n5111), .B(n5110), .Z(n5113) );
  XNOR U6254 ( .A(n5112), .B(n5113), .Z(n5067) );
  XOR U6255 ( .A(n5068), .B(n5067), .Z(n5069) );
  NAND U6256 ( .A(n4991), .B(n4990), .Z(n4995) );
  NAND U6257 ( .A(n4993), .B(n4992), .Z(n4994) );
  AND U6258 ( .A(n4995), .B(n4994), .Z(n5070) );
  XOR U6259 ( .A(n5069), .B(n5070), .Z(n5128) );
  NAND U6260 ( .A(n4997), .B(n4996), .Z(n5001) );
  NAND U6261 ( .A(n4999), .B(n4998), .Z(n5000) );
  AND U6262 ( .A(n5001), .B(n5000), .Z(n5129) );
  XOR U6263 ( .A(n5128), .B(n5129), .Z(n5130) );
  XNOR U6264 ( .A(n5131), .B(n5130), .Z(n5135) );
  NANDN U6265 ( .A(n5003), .B(n5002), .Z(n5007) );
  NAND U6266 ( .A(n5005), .B(n5004), .Z(n5006) );
  AND U6267 ( .A(n5007), .B(n5006), .Z(n5143) );
  NAND U6268 ( .A(n5009), .B(n5008), .Z(n5013) );
  NAND U6269 ( .A(n5011), .B(n5010), .Z(n5012) );
  AND U6270 ( .A(n5013), .B(n5012), .Z(n5141) );
  NANDN U6271 ( .A(n5015), .B(n5014), .Z(n5019) );
  NANDN U6272 ( .A(n5017), .B(n5016), .Z(n5018) );
  AND U6273 ( .A(n5019), .B(n5018), .Z(n5140) );
  XNOR U6274 ( .A(n5143), .B(n5142), .Z(n5134) );
  XOR U6275 ( .A(n5135), .B(n5134), .Z(n5136) );
  XOR U6276 ( .A(n5137), .B(n5136), .Z(n5152) );
  NAND U6277 ( .A(n5021), .B(n5020), .Z(n5025) );
  NANDN U6278 ( .A(n5023), .B(n5022), .Z(n5024) );
  AND U6279 ( .A(n5025), .B(n5024), .Z(n5150) );
  NANDN U6280 ( .A(n5027), .B(n5026), .Z(n5031) );
  NANDN U6281 ( .A(n5029), .B(n5028), .Z(n5030) );
  AND U6282 ( .A(n5031), .B(n5030), .Z(n5149) );
  XOR U6283 ( .A(n5150), .B(n5149), .Z(n5151) );
  XOR U6284 ( .A(n5146), .B(n5148), .Z(n5032) );
  XNOR U6285 ( .A(n5147), .B(n5032), .Z(N117) );
  NAND U6286 ( .A(n5034), .B(n5033), .Z(n5038) );
  NAND U6287 ( .A(n5036), .B(n5035), .Z(n5037) );
  NAND U6288 ( .A(n5038), .B(n5037), .Z(n5165) );
  AND U6289 ( .A(x[239]), .B(y[1835]), .Z(n5895) );
  NAND U6290 ( .A(n5895), .B(n5039), .Z(n5043) );
  NAND U6291 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U6292 ( .A(n5043), .B(n5042), .Z(n5199) );
  AND U6293 ( .A(x[224]), .B(y[1845]), .Z(n5219) );
  NAND U6294 ( .A(x[245]), .B(y[1824]), .Z(n5220) );
  AND U6295 ( .A(o[52]), .B(n5044), .Z(n5221) );
  XOR U6296 ( .A(n5222), .B(n5221), .Z(n5198) );
  AND U6297 ( .A(x[229]), .B(y[1840]), .Z(n5204) );
  AND U6298 ( .A(x[240]), .B(y[1829]), .Z(n5203) );
  XOR U6299 ( .A(n5204), .B(n5203), .Z(n5206) );
  AND U6300 ( .A(x[239]), .B(y[1830]), .Z(n5205) );
  XOR U6301 ( .A(n5206), .B(n5205), .Z(n5197) );
  XOR U6302 ( .A(n5198), .B(n5197), .Z(n5200) );
  XOR U6303 ( .A(n5199), .B(n5200), .Z(n5244) );
  AND U6304 ( .A(x[242]), .B(y[1832]), .Z(n5907) );
  NAND U6305 ( .A(n5907), .B(n5045), .Z(n5049) );
  NAND U6306 ( .A(n5047), .B(n5046), .Z(n5048) );
  AND U6307 ( .A(n5049), .B(n5048), .Z(n5242) );
  AND U6308 ( .A(x[235]), .B(y[1843]), .Z(n6561) );
  AND U6309 ( .A(x[225]), .B(y[1833]), .Z(n5050) );
  NAND U6310 ( .A(n6561), .B(n5050), .Z(n5054) );
  NAND U6311 ( .A(n5052), .B(n5051), .Z(n5053) );
  NAND U6312 ( .A(n5054), .B(n5053), .Z(n5241) );
  XNOR U6313 ( .A(n5244), .B(n5243), .Z(n5236) );
  NAND U6314 ( .A(n5056), .B(n5055), .Z(n5060) );
  NAND U6315 ( .A(n5058), .B(n5057), .Z(n5059) );
  NAND U6316 ( .A(n5060), .B(n5059), .Z(n5235) );
  XOR U6317 ( .A(n5236), .B(n5235), .Z(n5238) );
  NAND U6318 ( .A(n5062), .B(n5061), .Z(n5066) );
  NAND U6319 ( .A(n5064), .B(n5063), .Z(n5065) );
  AND U6320 ( .A(n5066), .B(n5065), .Z(n5237) );
  XNOR U6321 ( .A(n5238), .B(n5237), .Z(n5163) );
  NAND U6322 ( .A(n5068), .B(n5067), .Z(n5072) );
  NAND U6323 ( .A(n5070), .B(n5069), .Z(n5071) );
  AND U6324 ( .A(n5072), .B(n5071), .Z(n5162) );
  XOR U6325 ( .A(n5163), .B(n5162), .Z(n5164) );
  XNOR U6326 ( .A(n5165), .B(n5164), .Z(n5158) );
  NAND U6327 ( .A(n5074), .B(n5073), .Z(n5078) );
  NAND U6328 ( .A(n5076), .B(n5075), .Z(n5077) );
  NAND U6329 ( .A(n5078), .B(n5077), .Z(n5262) );
  NAND U6330 ( .A(n5900), .B(n5079), .Z(n5083) );
  NAND U6331 ( .A(n5081), .B(n5080), .Z(n5082) );
  NAND U6332 ( .A(n5083), .B(n5082), .Z(n5169) );
  NAND U6333 ( .A(n6514), .B(n5084), .Z(n5088) );
  NAND U6334 ( .A(n5086), .B(n5085), .Z(n5087) );
  NAND U6335 ( .A(n5088), .B(n5087), .Z(n5256) );
  AND U6336 ( .A(y[1826]), .B(x[243]), .Z(n5090) );
  NAND U6337 ( .A(y[1834]), .B(x[235]), .Z(n5089) );
  XNOR U6338 ( .A(n5090), .B(n5089), .Z(n5188) );
  AND U6339 ( .A(x[244]), .B(y[1825]), .Z(n5218) );
  XOR U6340 ( .A(n5218), .B(o[53]), .Z(n5187) );
  XOR U6341 ( .A(n5188), .B(n5187), .Z(n5254) );
  AND U6342 ( .A(y[1827]), .B(x[242]), .Z(n5092) );
  NAND U6343 ( .A(y[1835]), .B(x[234]), .Z(n5091) );
  XNOR U6344 ( .A(n5092), .B(n5091), .Z(n5226) );
  NAND U6345 ( .A(x[225]), .B(y[1844]), .Z(n5227) );
  XOR U6346 ( .A(n5254), .B(n5253), .Z(n5255) );
  XOR U6347 ( .A(n5256), .B(n5255), .Z(n5168) );
  XOR U6348 ( .A(n5169), .B(n5168), .Z(n5171) );
  AND U6349 ( .A(x[231]), .B(y[1838]), .Z(n5439) );
  AND U6350 ( .A(y[1839]), .B(x[230]), .Z(n5094) );
  NAND U6351 ( .A(y[1831]), .B(x[238]), .Z(n5093) );
  XOR U6352 ( .A(n5094), .B(n5093), .Z(n5230) );
  NAND U6353 ( .A(x[233]), .B(y[1836]), .Z(n5175) );
  NAND U6354 ( .A(x[232]), .B(y[1837]), .Z(n5174) );
  XOR U6355 ( .A(n5175), .B(n5174), .Z(n5176) );
  AND U6356 ( .A(y[1833]), .B(x[236]), .Z(n5096) );
  NAND U6357 ( .A(y[1828]), .B(x[241]), .Z(n5095) );
  XNOR U6358 ( .A(n5096), .B(n5095), .Z(n5180) );
  NAND U6359 ( .A(x[226]), .B(y[1843]), .Z(n5181) );
  AND U6360 ( .A(y[1832]), .B(x[237]), .Z(n5098) );
  NAND U6361 ( .A(y[1842]), .B(x[227]), .Z(n5097) );
  XNOR U6362 ( .A(n5098), .B(n5097), .Z(n5215) );
  AND U6363 ( .A(x[228]), .B(y[1841]), .Z(n5214) );
  XOR U6364 ( .A(n5215), .B(n5214), .Z(n5191) );
  XOR U6365 ( .A(n5192), .B(n5191), .Z(n5193) );
  NAND U6366 ( .A(n5204), .B(n5099), .Z(n5103) );
  NAND U6367 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U6368 ( .A(n5103), .B(n5102), .Z(n5248) );
  NAND U6369 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U6370 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U6371 ( .A(n5109), .B(n5108), .Z(n5247) );
  XOR U6372 ( .A(n5248), .B(n5247), .Z(n5249) );
  XOR U6373 ( .A(n5250), .B(n5249), .Z(n5170) );
  XOR U6374 ( .A(n5171), .B(n5170), .Z(n5260) );
  NAND U6375 ( .A(n5111), .B(n5110), .Z(n5115) );
  NAND U6376 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U6377 ( .A(n5115), .B(n5114), .Z(n5267) );
  NAND U6378 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U6379 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U6380 ( .A(n5121), .B(n5120), .Z(n5266) );
  NAND U6381 ( .A(n5123), .B(n5122), .Z(n5127) );
  NAND U6382 ( .A(n5125), .B(n5124), .Z(n5126) );
  NAND U6383 ( .A(n5127), .B(n5126), .Z(n5265) );
  XOR U6384 ( .A(n5266), .B(n5265), .Z(n5268) );
  XOR U6385 ( .A(n5267), .B(n5268), .Z(n5259) );
  XOR U6386 ( .A(n5260), .B(n5259), .Z(n5261) );
  XNOR U6387 ( .A(n5262), .B(n5261), .Z(n5157) );
  NAND U6388 ( .A(n5129), .B(n5128), .Z(n5133) );
  NAND U6389 ( .A(n5131), .B(n5130), .Z(n5132) );
  NAND U6390 ( .A(n5133), .B(n5132), .Z(n5156) );
  XOR U6391 ( .A(n5157), .B(n5156), .Z(n5159) );
  XNOR U6392 ( .A(n5158), .B(n5159), .Z(n5280) );
  NAND U6393 ( .A(n5135), .B(n5134), .Z(n5139) );
  NAND U6394 ( .A(n5137), .B(n5136), .Z(n5138) );
  AND U6395 ( .A(n5139), .B(n5138), .Z(n5279) );
  NANDN U6396 ( .A(n5141), .B(n5140), .Z(n5145) );
  NAND U6397 ( .A(n5143), .B(n5142), .Z(n5144) );
  AND U6398 ( .A(n5145), .B(n5144), .Z(n5278) );
  XNOR U6399 ( .A(n5280), .B(n5281), .Z(n5274) );
  NAND U6400 ( .A(n5150), .B(n5149), .Z(n5154) );
  NANDN U6401 ( .A(n5152), .B(n5151), .Z(n5153) );
  AND U6402 ( .A(n5154), .B(n5153), .Z(n5272) );
  IV U6403 ( .A(n5272), .Z(n5271) );
  XOR U6404 ( .A(n5273), .B(n5271), .Z(n5155) );
  XNOR U6405 ( .A(n5274), .B(n5155), .Z(N118) );
  NAND U6406 ( .A(n5157), .B(n5156), .Z(n5161) );
  NAND U6407 ( .A(n5159), .B(n5158), .Z(n5160) );
  AND U6408 ( .A(n5161), .B(n5160), .Z(n5415) );
  NAND U6409 ( .A(n5163), .B(n5162), .Z(n5167) );
  NAND U6410 ( .A(n5165), .B(n5164), .Z(n5166) );
  NAND U6411 ( .A(n5167), .B(n5166), .Z(n5413) );
  NAND U6412 ( .A(n5169), .B(n5168), .Z(n5173) );
  NAND U6413 ( .A(n5171), .B(n5170), .Z(n5172) );
  AND U6414 ( .A(n5173), .B(n5172), .Z(n5402) );
  NAND U6415 ( .A(n5175), .B(n5174), .Z(n5179) );
  NANDN U6416 ( .A(n5177), .B(n5176), .Z(n5178) );
  AND U6417 ( .A(n5179), .B(n5178), .Z(n5396) );
  NANDN U6418 ( .A(n5908), .B(n5347), .Z(n5183) );
  NANDN U6419 ( .A(n5181), .B(n5180), .Z(n5182) );
  AND U6420 ( .A(n5183), .B(n5182), .Z(n5324) );
  AND U6421 ( .A(x[229]), .B(y[1841]), .Z(n5369) );
  NAND U6422 ( .A(x[241]), .B(y[1829]), .Z(n5370) );
  NAND U6423 ( .A(x[240]), .B(y[1830]), .Z(n5372) );
  AND U6424 ( .A(y[1828]), .B(x[242]), .Z(n5185) );
  NAND U6425 ( .A(y[1834]), .B(x[236]), .Z(n5184) );
  XNOR U6426 ( .A(n5185), .B(n5184), .Z(n5348) );
  NAND U6427 ( .A(x[228]), .B(y[1842]), .Z(n5349) );
  XOR U6428 ( .A(n5322), .B(n5321), .Z(n5323) );
  AND U6429 ( .A(x[243]), .B(y[1834]), .Z(n6419) );
  NAND U6430 ( .A(n6419), .B(n5186), .Z(n5190) );
  NAND U6431 ( .A(n5188), .B(n5187), .Z(n5189) );
  AND U6432 ( .A(n5190), .B(n5189), .Z(n5394) );
  XOR U6433 ( .A(n5393), .B(n5394), .Z(n5395) );
  NAND U6434 ( .A(n5192), .B(n5191), .Z(n5196) );
  NANDN U6435 ( .A(n5194), .B(n5193), .Z(n5195) );
  AND U6436 ( .A(n5196), .B(n5195), .Z(n5382) );
  NAND U6437 ( .A(n5198), .B(n5197), .Z(n5202) );
  NAND U6438 ( .A(n5200), .B(n5199), .Z(n5201) );
  NAND U6439 ( .A(n5202), .B(n5201), .Z(n5381) );
  NAND U6440 ( .A(n5204), .B(n5203), .Z(n5208) );
  AND U6441 ( .A(n5206), .B(n5205), .Z(n5207) );
  ANDN U6442 ( .B(n5208), .A(n5207), .Z(n5344) );
  AND U6443 ( .A(y[1833]), .B(x[237]), .Z(n5210) );
  NAND U6444 ( .A(y[1826]), .B(x[244]), .Z(n5209) );
  XNOR U6445 ( .A(n5210), .B(n5209), .Z(n5365) );
  NAND U6446 ( .A(x[226]), .B(y[1844]), .Z(n5366) );
  AND U6447 ( .A(y[1840]), .B(x[230]), .Z(n5212) );
  NAND U6448 ( .A(y[1831]), .B(x[239]), .Z(n5211) );
  XNOR U6449 ( .A(n5212), .B(n5211), .Z(n5377) );
  XOR U6450 ( .A(n5342), .B(n5341), .Z(n5343) );
  AND U6451 ( .A(x[237]), .B(y[1842]), .Z(n6572) );
  NAND U6452 ( .A(n5213), .B(n6572), .Z(n5217) );
  NAND U6453 ( .A(n5215), .B(n5214), .Z(n5216) );
  AND U6454 ( .A(n5217), .B(n5216), .Z(n5312) );
  AND U6455 ( .A(x[225]), .B(y[1845]), .Z(n5335) );
  XOR U6456 ( .A(n5336), .B(n5335), .Z(n5334) );
  AND U6457 ( .A(n5218), .B(o[53]), .Z(n5333) );
  XOR U6458 ( .A(n5334), .B(n5333), .Z(n5310) );
  AND U6459 ( .A(x[238]), .B(y[1832]), .Z(n5327) );
  AND U6460 ( .A(x[227]), .B(y[1843]), .Z(n5328) );
  XOR U6461 ( .A(n5327), .B(n5328), .Z(n5329) );
  AND U6462 ( .A(x[243]), .B(y[1827]), .Z(n5330) );
  XOR U6463 ( .A(n5329), .B(n5330), .Z(n5309) );
  XOR U6464 ( .A(n5310), .B(n5309), .Z(n5311) );
  XOR U6465 ( .A(n5388), .B(n5387), .Z(n5390) );
  NANDN U6466 ( .A(n5220), .B(n5219), .Z(n5224) );
  NAND U6467 ( .A(n5222), .B(n5221), .Z(n5223) );
  AND U6468 ( .A(n5224), .B(n5223), .Z(n5304) );
  AND U6469 ( .A(x[242]), .B(y[1835]), .Z(n6422) );
  NAND U6470 ( .A(n6422), .B(n5225), .Z(n5229) );
  NANDN U6471 ( .A(n5227), .B(n5226), .Z(n5228) );
  NAND U6472 ( .A(n5229), .B(n5228), .Z(n5303) );
  AND U6473 ( .A(x[238]), .B(y[1839]), .Z(n6432) );
  NAND U6474 ( .A(n6432), .B(n5376), .Z(n5232) );
  NANDN U6475 ( .A(n5230), .B(n5439), .Z(n5231) );
  NAND U6476 ( .A(n5232), .B(n5231), .Z(n5317) );
  AND U6477 ( .A(x[224]), .B(y[1846]), .Z(n5352) );
  NAND U6478 ( .A(x[246]), .B(y[1824]), .Z(n5353) );
  AND U6479 ( .A(x[245]), .B(y[1825]), .Z(n5375) );
  XOR U6480 ( .A(o[54]), .B(n5375), .Z(n5354) );
  XOR U6481 ( .A(n5355), .B(n5354), .Z(n5316) );
  AND U6482 ( .A(y[1839]), .B(x[231]), .Z(n5234) );
  NAND U6483 ( .A(y[1838]), .B(x[232]), .Z(n5233) );
  XNOR U6484 ( .A(n5234), .B(n5233), .Z(n5359) );
  XOR U6485 ( .A(n5359), .B(n5358), .Z(n5315) );
  XOR U6486 ( .A(n5316), .B(n5315), .Z(n5318) );
  XOR U6487 ( .A(n5317), .B(n5318), .Z(n5305) );
  XOR U6488 ( .A(n5306), .B(n5305), .Z(n5389) );
  XOR U6489 ( .A(n5390), .B(n5389), .Z(n5383) );
  XOR U6490 ( .A(n5384), .B(n5383), .Z(n5400) );
  XOR U6491 ( .A(n5399), .B(n5400), .Z(n5401) );
  NAND U6492 ( .A(n5236), .B(n5235), .Z(n5240) );
  NAND U6493 ( .A(n5238), .B(n5237), .Z(n5239) );
  NAND U6494 ( .A(n5240), .B(n5239), .Z(n5292) );
  NANDN U6495 ( .A(n5242), .B(n5241), .Z(n5246) );
  NAND U6496 ( .A(n5244), .B(n5243), .Z(n5245) );
  AND U6497 ( .A(n5246), .B(n5245), .Z(n5300) );
  NAND U6498 ( .A(n5248), .B(n5247), .Z(n5252) );
  NAND U6499 ( .A(n5250), .B(n5249), .Z(n5251) );
  AND U6500 ( .A(n5252), .B(n5251), .Z(n5298) );
  NAND U6501 ( .A(n5254), .B(n5253), .Z(n5258) );
  NAND U6502 ( .A(n5256), .B(n5255), .Z(n5257) );
  NAND U6503 ( .A(n5258), .B(n5257), .Z(n5297) );
  XOR U6504 ( .A(n5300), .B(n5299), .Z(n5291) );
  XOR U6505 ( .A(n5292), .B(n5291), .Z(n5294) );
  XNOR U6506 ( .A(n5293), .B(n5294), .Z(n5287) );
  NAND U6507 ( .A(n5260), .B(n5259), .Z(n5264) );
  NAND U6508 ( .A(n5262), .B(n5261), .Z(n5263) );
  NAND U6509 ( .A(n5264), .B(n5263), .Z(n5286) );
  NAND U6510 ( .A(n5266), .B(n5265), .Z(n5270) );
  NAND U6511 ( .A(n5268), .B(n5267), .Z(n5269) );
  NAND U6512 ( .A(n5270), .B(n5269), .Z(n5285) );
  XOR U6513 ( .A(n5286), .B(n5285), .Z(n5288) );
  XOR U6514 ( .A(n5287), .B(n5288), .Z(n5412) );
  XOR U6515 ( .A(n5413), .B(n5412), .Z(n5414) );
  XNOR U6516 ( .A(n5415), .B(n5414), .Z(n5408) );
  OR U6517 ( .A(n5273), .B(n5271), .Z(n5277) );
  ANDN U6518 ( .B(n5273), .A(n5272), .Z(n5275) );
  OR U6519 ( .A(n5275), .B(n5274), .Z(n5276) );
  AND U6520 ( .A(n5277), .B(n5276), .Z(n5407) );
  NANDN U6521 ( .A(n5279), .B(n5278), .Z(n5283) );
  NAND U6522 ( .A(n5281), .B(n5280), .Z(n5282) );
  NAND U6523 ( .A(n5283), .B(n5282), .Z(n5406) );
  IV U6524 ( .A(n5406), .Z(n5405) );
  XOR U6525 ( .A(n5407), .B(n5405), .Z(n5284) );
  XNOR U6526 ( .A(n5408), .B(n5284), .Z(N119) );
  NAND U6527 ( .A(n5286), .B(n5285), .Z(n5290) );
  NAND U6528 ( .A(n5288), .B(n5287), .Z(n5289) );
  AND U6529 ( .A(n5290), .B(n5289), .Z(n5560) );
  NAND U6530 ( .A(n5292), .B(n5291), .Z(n5296) );
  NAND U6531 ( .A(n5294), .B(n5293), .Z(n5295) );
  NAND U6532 ( .A(n5296), .B(n5295), .Z(n5558) );
  NANDN U6533 ( .A(n5298), .B(n5297), .Z(n5302) );
  NANDN U6534 ( .A(n5300), .B(n5299), .Z(n5301) );
  AND U6535 ( .A(n5302), .B(n5301), .Z(n5535) );
  NANDN U6536 ( .A(n5304), .B(n5303), .Z(n5308) );
  NAND U6537 ( .A(n5306), .B(n5305), .Z(n5307) );
  NAND U6538 ( .A(n5308), .B(n5307), .Z(n5528) );
  NAND U6539 ( .A(n5310), .B(n5309), .Z(n5314) );
  NANDN U6540 ( .A(n5312), .B(n5311), .Z(n5313) );
  NAND U6541 ( .A(n5314), .B(n5313), .Z(n5527) );
  NAND U6542 ( .A(n5316), .B(n5315), .Z(n5320) );
  NAND U6543 ( .A(n5318), .B(n5317), .Z(n5319) );
  NAND U6544 ( .A(n5320), .B(n5319), .Z(n5526) );
  XOR U6545 ( .A(n5527), .B(n5526), .Z(n5529) );
  XOR U6546 ( .A(n5528), .B(n5529), .Z(n5546) );
  NAND U6547 ( .A(n5322), .B(n5321), .Z(n5326) );
  NANDN U6548 ( .A(n5324), .B(n5323), .Z(n5325) );
  NAND U6549 ( .A(n5326), .B(n5325), .Z(n5544) );
  NAND U6550 ( .A(n5328), .B(n5327), .Z(n5332) );
  NAND U6551 ( .A(n5330), .B(n5329), .Z(n5331) );
  NAND U6552 ( .A(n5332), .B(n5331), .Z(n5473) );
  AND U6553 ( .A(n5334), .B(n5333), .Z(n5338) );
  NAND U6554 ( .A(n5336), .B(n5335), .Z(n5337) );
  NANDN U6555 ( .A(n5338), .B(n5337), .Z(n5472) );
  XOR U6556 ( .A(n5473), .B(n5472), .Z(n5475) );
  AND U6557 ( .A(y[1840]), .B(x[231]), .Z(n5340) );
  NAND U6558 ( .A(y[1838]), .B(x[233]), .Z(n5339) );
  XNOR U6559 ( .A(n5340), .B(n5339), .Z(n5440) );
  AND U6560 ( .A(x[234]), .B(y[1837]), .Z(n5479) );
  XOR U6561 ( .A(n5478), .B(n5479), .Z(n5481) );
  AND U6562 ( .A(x[230]), .B(y[1841]), .Z(n5431) );
  AND U6563 ( .A(x[239]), .B(y[1832]), .Z(n5432) );
  XOR U6564 ( .A(n5431), .B(n5432), .Z(n5433) );
  AND U6565 ( .A(x[235]), .B(y[1836]), .Z(n5434) );
  XOR U6566 ( .A(n5433), .B(n5434), .Z(n5480) );
  XOR U6567 ( .A(n5481), .B(n5480), .Z(n5474) );
  XOR U6568 ( .A(n5475), .B(n5474), .Z(n5545) );
  XNOR U6569 ( .A(n5544), .B(n5545), .Z(n5547) );
  NAND U6570 ( .A(n5342), .B(n5341), .Z(n5346) );
  NANDN U6571 ( .A(n5344), .B(n5343), .Z(n5345) );
  AND U6572 ( .A(n5346), .B(n5345), .Z(n5467) );
  NAND U6573 ( .A(x[242]), .B(y[1834]), .Z(n6272) );
  NANDN U6574 ( .A(n6272), .B(n5347), .Z(n5351) );
  NANDN U6575 ( .A(n5349), .B(n5348), .Z(n5350) );
  AND U6576 ( .A(n5351), .B(n5350), .Z(n5503) );
  NANDN U6577 ( .A(n5353), .B(n5352), .Z(n5357) );
  NAND U6578 ( .A(n5355), .B(n5354), .Z(n5356) );
  NAND U6579 ( .A(n5357), .B(n5356), .Z(n5502) );
  NANDN U6580 ( .A(n5441), .B(n5439), .Z(n5361) );
  NAND U6581 ( .A(n5359), .B(n5358), .Z(n5360) );
  AND U6582 ( .A(n5361), .B(n5360), .Z(n5517) );
  AND U6583 ( .A(x[224]), .B(y[1847]), .Z(n5450) );
  AND U6584 ( .A(x[247]), .B(y[1824]), .Z(n5451) );
  XOR U6585 ( .A(n5450), .B(n5451), .Z(n5453) );
  AND U6586 ( .A(x[246]), .B(y[1825]), .Z(n5430) );
  XOR U6587 ( .A(o[55]), .B(n5430), .Z(n5452) );
  XOR U6588 ( .A(n5453), .B(n5452), .Z(n5515) );
  NAND U6589 ( .A(y[1827]), .B(x[244]), .Z(n5362) );
  XNOR U6590 ( .A(n5363), .B(n5362), .Z(n5426) );
  AND U6591 ( .A(x[243]), .B(y[1828]), .Z(n5427) );
  XOR U6592 ( .A(n5426), .B(n5427), .Z(n5514) );
  XOR U6593 ( .A(n5515), .B(n5514), .Z(n5516) );
  XOR U6594 ( .A(n5505), .B(n5504), .Z(n5466) );
  NAND U6595 ( .A(x[244]), .B(y[1833]), .Z(n6444) );
  AND U6596 ( .A(x[237]), .B(y[1826]), .Z(n5364) );
  NANDN U6597 ( .A(n6444), .B(n5364), .Z(n5368) );
  NANDN U6598 ( .A(n5366), .B(n5365), .Z(n5367) );
  AND U6599 ( .A(n5368), .B(n5367), .Z(n5461) );
  NANDN U6600 ( .A(n5370), .B(n5369), .Z(n5374) );
  NANDN U6601 ( .A(n5372), .B(n5371), .Z(n5373) );
  AND U6602 ( .A(n5374), .B(n5373), .Z(n5523) );
  AND U6603 ( .A(x[237]), .B(y[1834]), .Z(n5496) );
  AND U6604 ( .A(x[226]), .B(y[1845]), .Z(n5497) );
  XOR U6605 ( .A(n5496), .B(n5497), .Z(n5498) );
  AND U6606 ( .A(x[245]), .B(y[1826]), .Z(n5499) );
  XOR U6607 ( .A(n5498), .B(n5499), .Z(n5521) );
  AND U6608 ( .A(x[236]), .B(y[1835]), .Z(n5444) );
  AND U6609 ( .A(x[225]), .B(y[1846]), .Z(n5445) );
  XOR U6610 ( .A(n5444), .B(n5445), .Z(n5447) );
  AND U6611 ( .A(o[54]), .B(n5375), .Z(n5446) );
  XOR U6612 ( .A(n5447), .B(n5446), .Z(n5520) );
  XOR U6613 ( .A(n5521), .B(n5520), .Z(n5522) );
  AND U6614 ( .A(x[239]), .B(y[1840]), .Z(n6712) );
  NAND U6615 ( .A(n6712), .B(n5376), .Z(n5380) );
  NANDN U6616 ( .A(n5378), .B(n5377), .Z(n5379) );
  AND U6617 ( .A(n5380), .B(n5379), .Z(n5511) );
  AND U6618 ( .A(x[238]), .B(y[1833]), .Z(n5490) );
  AND U6619 ( .A(x[227]), .B(y[1844]), .Z(n5491) );
  XOR U6620 ( .A(n5490), .B(n5491), .Z(n5492) );
  AND U6621 ( .A(x[228]), .B(y[1843]), .Z(n5493) );
  XOR U6622 ( .A(n5492), .B(n5493), .Z(n5509) );
  AND U6623 ( .A(x[229]), .B(y[1842]), .Z(n5484) );
  AND U6624 ( .A(x[242]), .B(y[1829]), .Z(n5485) );
  XOR U6625 ( .A(n5484), .B(n5485), .Z(n5486) );
  AND U6626 ( .A(x[241]), .B(y[1830]), .Z(n5487) );
  XOR U6627 ( .A(n5486), .B(n5487), .Z(n5508) );
  XOR U6628 ( .A(n5509), .B(n5508), .Z(n5510) );
  XOR U6629 ( .A(n5463), .B(n5462), .Z(n5468) );
  XOR U6630 ( .A(n5469), .B(n5468), .Z(n5532) );
  XOR U6631 ( .A(n5533), .B(n5532), .Z(n5534) );
  NANDN U6632 ( .A(n5382), .B(n5381), .Z(n5386) );
  NAND U6633 ( .A(n5384), .B(n5383), .Z(n5385) );
  AND U6634 ( .A(n5386), .B(n5385), .Z(n5541) );
  NAND U6635 ( .A(n5388), .B(n5387), .Z(n5392) );
  NAND U6636 ( .A(n5390), .B(n5389), .Z(n5391) );
  AND U6637 ( .A(n5392), .B(n5391), .Z(n5539) );
  NAND U6638 ( .A(n5394), .B(n5393), .Z(n5398) );
  NANDN U6639 ( .A(n5396), .B(n5395), .Z(n5397) );
  AND U6640 ( .A(n5398), .B(n5397), .Z(n5538) );
  NAND U6641 ( .A(n5400), .B(n5399), .Z(n5404) );
  NANDN U6642 ( .A(n5402), .B(n5401), .Z(n5403) );
  AND U6643 ( .A(n5404), .B(n5403), .Z(n5420) );
  XOR U6644 ( .A(n5419), .B(n5420), .Z(n5422) );
  XOR U6645 ( .A(n5421), .B(n5422), .Z(n5557) );
  XOR U6646 ( .A(n5558), .B(n5557), .Z(n5559) );
  XNOR U6647 ( .A(n5560), .B(n5559), .Z(n5553) );
  OR U6648 ( .A(n5407), .B(n5405), .Z(n5411) );
  ANDN U6649 ( .B(n5407), .A(n5406), .Z(n5409) );
  OR U6650 ( .A(n5409), .B(n5408), .Z(n5410) );
  AND U6651 ( .A(n5411), .B(n5410), .Z(n5551) );
  NAND U6652 ( .A(n5413), .B(n5412), .Z(n5417) );
  NAND U6653 ( .A(n5415), .B(n5414), .Z(n5416) );
  AND U6654 ( .A(n5417), .B(n5416), .Z(n5552) );
  IV U6655 ( .A(n5552), .Z(n5550) );
  XOR U6656 ( .A(n5551), .B(n5550), .Z(n5418) );
  XNOR U6657 ( .A(n5553), .B(n5418), .Z(N120) );
  NAND U6658 ( .A(n5420), .B(n5419), .Z(n5424) );
  NAND U6659 ( .A(n5422), .B(n5421), .Z(n5423) );
  AND U6660 ( .A(n5424), .B(n5423), .Z(n5567) );
  AND U6661 ( .A(x[244]), .B(y[1831]), .Z(n5425) );
  NAND U6662 ( .A(n5425), .B(n5603), .Z(n5429) );
  NAND U6663 ( .A(n5427), .B(n5426), .Z(n5428) );
  NAND U6664 ( .A(n5429), .B(n5428), .Z(n5623) );
  AND U6665 ( .A(x[246]), .B(y[1826]), .Z(n5644) );
  XOR U6666 ( .A(n5645), .B(n5644), .Z(n5643) );
  AND U6667 ( .A(x[226]), .B(y[1846]), .Z(n5642) );
  XOR U6668 ( .A(n5643), .B(n5642), .Z(n5621) );
  AND U6669 ( .A(x[225]), .B(y[1847]), .Z(n5650) );
  XOR U6670 ( .A(n5651), .B(n5650), .Z(n5649) );
  AND U6671 ( .A(o[55]), .B(n5430), .Z(n5648) );
  XOR U6672 ( .A(n5649), .B(n5648), .Z(n5620) );
  XOR U6673 ( .A(n5621), .B(n5620), .Z(n5622) );
  XOR U6674 ( .A(n5623), .B(n5622), .Z(n5681) );
  NAND U6675 ( .A(n5432), .B(n5431), .Z(n5436) );
  NAND U6676 ( .A(n5434), .B(n5433), .Z(n5435) );
  NAND U6677 ( .A(n5436), .B(n5435), .Z(n5617) );
  AND U6678 ( .A(y[1832]), .B(x[240]), .Z(n5438) );
  NAND U6679 ( .A(y[1827]), .B(x[245]), .Z(n5437) );
  XNOR U6680 ( .A(n5438), .B(n5437), .Z(n5605) );
  AND U6681 ( .A(x[229]), .B(y[1843]), .Z(n5604) );
  XOR U6682 ( .A(n5605), .B(n5604), .Z(n5615) );
  AND U6683 ( .A(x[230]), .B(y[1842]), .Z(n5998) );
  AND U6684 ( .A(x[244]), .B(y[1828]), .Z(n5804) );
  XOR U6685 ( .A(n5998), .B(n5804), .Z(n5611) );
  AND U6686 ( .A(x[243]), .B(y[1829]), .Z(n5610) );
  XOR U6687 ( .A(n5611), .B(n5610), .Z(n5614) );
  XOR U6688 ( .A(n5615), .B(n5614), .Z(n5616) );
  XOR U6689 ( .A(n5617), .B(n5616), .Z(n5594) );
  NAND U6690 ( .A(n5730), .B(n5439), .Z(n5443) );
  NANDN U6691 ( .A(n5441), .B(n5440), .Z(n5442) );
  NAND U6692 ( .A(n5443), .B(n5442), .Z(n5592) );
  NAND U6693 ( .A(n5445), .B(n5444), .Z(n5449) );
  NAND U6694 ( .A(n5447), .B(n5446), .Z(n5448) );
  NAND U6695 ( .A(n5449), .B(n5448), .Z(n5591) );
  XOR U6696 ( .A(n5592), .B(n5591), .Z(n5593) );
  XOR U6697 ( .A(n5594), .B(n5593), .Z(n5680) );
  XOR U6698 ( .A(n5681), .B(n5680), .Z(n5683) );
  NAND U6699 ( .A(n5451), .B(n5450), .Z(n5455) );
  NAND U6700 ( .A(n5453), .B(n5452), .Z(n5454) );
  AND U6701 ( .A(n5455), .B(n5454), .Z(n5675) );
  AND U6702 ( .A(x[227]), .B(y[1845]), .Z(n5664) );
  XOR U6703 ( .A(n5665), .B(n5664), .Z(n5663) );
  AND U6704 ( .A(x[228]), .B(y[1844]), .Z(n5662) );
  XOR U6705 ( .A(n5663), .B(n5662), .Z(n5674) );
  AND U6706 ( .A(y[1839]), .B(x[233]), .Z(n5457) );
  NAND U6707 ( .A(y[1838]), .B(x[234]), .Z(n5456) );
  XNOR U6708 ( .A(n5457), .B(n5456), .Z(n5634) );
  AND U6709 ( .A(y[1834]), .B(x[238]), .Z(n5459) );
  NAND U6710 ( .A(y[1840]), .B(x[232]), .Z(n5458) );
  XNOR U6711 ( .A(n5459), .B(n5458), .Z(n5638) );
  NAND U6712 ( .A(x[235]), .B(y[1837]), .Z(n5639) );
  XOR U6713 ( .A(n5634), .B(n5633), .Z(n5676) );
  XOR U6714 ( .A(n5677), .B(n5676), .Z(n5682) );
  XOR U6715 ( .A(n5683), .B(n5682), .Z(n5693) );
  NANDN U6716 ( .A(n5461), .B(n5460), .Z(n5465) );
  NAND U6717 ( .A(n5463), .B(n5462), .Z(n5464) );
  AND U6718 ( .A(n5465), .B(n5464), .Z(n5692) );
  NANDN U6719 ( .A(n5467), .B(n5466), .Z(n5471) );
  NAND U6720 ( .A(n5469), .B(n5468), .Z(n5470) );
  NAND U6721 ( .A(n5471), .B(n5470), .Z(n5695) );
  NAND U6722 ( .A(n5473), .B(n5472), .Z(n5477) );
  NAND U6723 ( .A(n5475), .B(n5474), .Z(n5476) );
  NAND U6724 ( .A(n5477), .B(n5476), .Z(n5689) );
  NAND U6725 ( .A(n5479), .B(n5478), .Z(n5483) );
  NAND U6726 ( .A(n5481), .B(n5480), .Z(n5482) );
  NAND U6727 ( .A(n5483), .B(n5482), .Z(n5687) );
  NAND U6728 ( .A(n5485), .B(n5484), .Z(n5489) );
  NAND U6729 ( .A(n5487), .B(n5486), .Z(n5488) );
  NAND U6730 ( .A(n5489), .B(n5488), .Z(n5600) );
  AND U6731 ( .A(x[224]), .B(y[1848]), .Z(n5669) );
  AND U6732 ( .A(x[248]), .B(y[1824]), .Z(n5668) );
  XOR U6733 ( .A(n5669), .B(n5668), .Z(n5671) );
  AND U6734 ( .A(x[247]), .B(y[1825]), .Z(n5661) );
  XOR U6735 ( .A(n5661), .B(o[56]), .Z(n5670) );
  XOR U6736 ( .A(n5671), .B(n5670), .Z(n5598) );
  AND U6737 ( .A(x[231]), .B(y[1841]), .Z(n5655) );
  AND U6738 ( .A(x[242]), .B(y[1830]), .Z(n5654) );
  XOR U6739 ( .A(n5655), .B(n5654), .Z(n5657) );
  AND U6740 ( .A(x[241]), .B(y[1831]), .Z(n5656) );
  XOR U6741 ( .A(n5657), .B(n5656), .Z(n5597) );
  XOR U6742 ( .A(n5598), .B(n5597), .Z(n5599) );
  XOR U6743 ( .A(n5600), .B(n5599), .Z(n5588) );
  NAND U6744 ( .A(n5491), .B(n5490), .Z(n5495) );
  NAND U6745 ( .A(n5493), .B(n5492), .Z(n5494) );
  NAND U6746 ( .A(n5495), .B(n5494), .Z(n5586) );
  NAND U6747 ( .A(n5497), .B(n5496), .Z(n5501) );
  NAND U6748 ( .A(n5499), .B(n5498), .Z(n5500) );
  NAND U6749 ( .A(n5501), .B(n5500), .Z(n5585) );
  XOR U6750 ( .A(n5586), .B(n5585), .Z(n5587) );
  XOR U6751 ( .A(n5588), .B(n5587), .Z(n5686) );
  XOR U6752 ( .A(n5687), .B(n5686), .Z(n5688) );
  XNOR U6753 ( .A(n5689), .B(n5688), .Z(n5581) );
  NANDN U6754 ( .A(n5503), .B(n5502), .Z(n5507) );
  NAND U6755 ( .A(n5505), .B(n5504), .Z(n5506) );
  AND U6756 ( .A(n5507), .B(n5506), .Z(n5629) );
  NAND U6757 ( .A(n5509), .B(n5508), .Z(n5513) );
  NANDN U6758 ( .A(n5511), .B(n5510), .Z(n5512) );
  AND U6759 ( .A(n5513), .B(n5512), .Z(n5626) );
  NAND U6760 ( .A(n5515), .B(n5514), .Z(n5519) );
  NANDN U6761 ( .A(n5517), .B(n5516), .Z(n5518) );
  NAND U6762 ( .A(n5519), .B(n5518), .Z(n5627) );
  XOR U6763 ( .A(n5629), .B(n5628), .Z(n5579) );
  NAND U6764 ( .A(n5521), .B(n5520), .Z(n5525) );
  NANDN U6765 ( .A(n5523), .B(n5522), .Z(n5524) );
  NAND U6766 ( .A(n5525), .B(n5524), .Z(n5580) );
  XOR U6767 ( .A(n5581), .B(n5582), .Z(n5699) );
  NAND U6768 ( .A(n5527), .B(n5526), .Z(n5531) );
  NAND U6769 ( .A(n5529), .B(n5528), .Z(n5530) );
  AND U6770 ( .A(n5531), .B(n5530), .Z(n5698) );
  XOR U6771 ( .A(n5699), .B(n5698), .Z(n5700) );
  XOR U6772 ( .A(n5701), .B(n5700), .Z(n5565) );
  NAND U6773 ( .A(n5533), .B(n5532), .Z(n5537) );
  NANDN U6774 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U6775 ( .A(n5537), .B(n5536), .Z(n5575) );
  NANDN U6776 ( .A(n5539), .B(n5538), .Z(n5543) );
  NANDN U6777 ( .A(n5541), .B(n5540), .Z(n5542) );
  NAND U6778 ( .A(n5543), .B(n5542), .Z(n5574) );
  NAND U6779 ( .A(n5545), .B(n5544), .Z(n5549) );
  NANDN U6780 ( .A(n5547), .B(n5546), .Z(n5548) );
  NAND U6781 ( .A(n5549), .B(n5548), .Z(n5573) );
  XOR U6782 ( .A(n5574), .B(n5573), .Z(n5576) );
  XOR U6783 ( .A(n5575), .B(n5576), .Z(n5564) );
  XNOR U6784 ( .A(n5567), .B(n5566), .Z(n5572) );
  NANDN U6785 ( .A(n5550), .B(n5551), .Z(n5556) );
  NOR U6786 ( .A(n5552), .B(n5551), .Z(n5554) );
  OR U6787 ( .A(n5554), .B(n5553), .Z(n5555) );
  AND U6788 ( .A(n5556), .B(n5555), .Z(n5570) );
  NAND U6789 ( .A(n5558), .B(n5557), .Z(n5562) );
  NAND U6790 ( .A(n5560), .B(n5559), .Z(n5561) );
  AND U6791 ( .A(n5562), .B(n5561), .Z(n5571) );
  XOR U6792 ( .A(n5570), .B(n5571), .Z(n5563) );
  XNOR U6793 ( .A(n5572), .B(n5563), .Z(N121) );
  NANDN U6794 ( .A(n5565), .B(n5564), .Z(n5569) );
  NAND U6795 ( .A(n5567), .B(n5566), .Z(n5568) );
  NAND U6796 ( .A(n5569), .B(n5568), .Z(n5846) );
  IV U6797 ( .A(n5846), .Z(n5845) );
  NAND U6798 ( .A(n5574), .B(n5573), .Z(n5578) );
  NAND U6799 ( .A(n5576), .B(n5575), .Z(n5577) );
  AND U6800 ( .A(n5578), .B(n5577), .Z(n5854) );
  NANDN U6801 ( .A(n5580), .B(n5579), .Z(n5584) );
  NAND U6802 ( .A(n5582), .B(n5581), .Z(n5583) );
  AND U6803 ( .A(n5584), .B(n5583), .Z(n5714) );
  NAND U6804 ( .A(n5586), .B(n5585), .Z(n5590) );
  NAND U6805 ( .A(n5588), .B(n5587), .Z(n5589) );
  NAND U6806 ( .A(n5590), .B(n5589), .Z(n5718) );
  NAND U6807 ( .A(n5592), .B(n5591), .Z(n5596) );
  NAND U6808 ( .A(n5594), .B(n5593), .Z(n5595) );
  NAND U6809 ( .A(n5596), .B(n5595), .Z(n5717) );
  XOR U6810 ( .A(n5718), .B(n5717), .Z(n5720) );
  NAND U6811 ( .A(n5598), .B(n5597), .Z(n5602) );
  NAND U6812 ( .A(n5600), .B(n5599), .Z(n5601) );
  AND U6813 ( .A(n5602), .B(n5601), .Z(n5750) );
  NAND U6814 ( .A(x[245]), .B(y[1832]), .Z(n6684) );
  NANDN U6815 ( .A(n6684), .B(n5603), .Z(n5607) );
  NAND U6816 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U6817 ( .A(n5607), .B(n5606), .Z(n5823) );
  AND U6818 ( .A(x[246]), .B(y[1827]), .Z(n5794) );
  AND U6819 ( .A(x[229]), .B(y[1844]), .Z(n5792) );
  NAND U6820 ( .A(x[241]), .B(y[1832]), .Z(n5791) );
  XNOR U6821 ( .A(n5792), .B(n5791), .Z(n5793) );
  XOR U6822 ( .A(n5794), .B(n5793), .Z(n5821) );
  AND U6823 ( .A(y[1829]), .B(x[244]), .Z(n5609) );
  NAND U6824 ( .A(y[1828]), .B(x[245]), .Z(n5608) );
  XNOR U6825 ( .A(n5609), .B(n5608), .Z(n5806) );
  AND U6826 ( .A(x[243]), .B(y[1830]), .Z(n5805) );
  XOR U6827 ( .A(n5806), .B(n5805), .Z(n5822) );
  XOR U6828 ( .A(n5821), .B(n5822), .Z(n5824) );
  XNOR U6829 ( .A(n5823), .B(n5824), .Z(n5748) );
  NAND U6830 ( .A(n5998), .B(n5804), .Z(n5613) );
  NAND U6831 ( .A(n5611), .B(n5610), .Z(n5612) );
  NAND U6832 ( .A(n5613), .B(n5612), .Z(n5829) );
  AND U6833 ( .A(x[239]), .B(y[1834]), .Z(n5812) );
  AND U6834 ( .A(x[242]), .B(y[1831]), .Z(n5810) );
  NAND U6835 ( .A(x[230]), .B(y[1843]), .Z(n5809) );
  XNOR U6836 ( .A(n5810), .B(n5809), .Z(n5811) );
  XOR U6837 ( .A(n5812), .B(n5811), .Z(n5828) );
  AND U6838 ( .A(x[247]), .B(y[1826]), .Z(n5788) );
  AND U6839 ( .A(x[228]), .B(y[1845]), .Z(n5786) );
  NAND U6840 ( .A(x[240]), .B(y[1833]), .Z(n5785) );
  XNOR U6841 ( .A(n5786), .B(n5785), .Z(n5787) );
  XOR U6842 ( .A(n5788), .B(n5787), .Z(n5827) );
  XNOR U6843 ( .A(n5828), .B(n5827), .Z(n5830) );
  XOR U6844 ( .A(n5829), .B(n5830), .Z(n5747) );
  XOR U6845 ( .A(n5748), .B(n5747), .Z(n5749) );
  XNOR U6846 ( .A(n5750), .B(n5749), .Z(n5762) );
  NAND U6847 ( .A(n5615), .B(n5614), .Z(n5619) );
  NAND U6848 ( .A(n5617), .B(n5616), .Z(n5618) );
  NAND U6849 ( .A(n5619), .B(n5618), .Z(n5760) );
  NAND U6850 ( .A(n5621), .B(n5620), .Z(n5625) );
  NAND U6851 ( .A(n5623), .B(n5622), .Z(n5624) );
  NAND U6852 ( .A(n5625), .B(n5624), .Z(n5759) );
  XOR U6853 ( .A(n5760), .B(n5759), .Z(n5761) );
  XOR U6854 ( .A(n5762), .B(n5761), .Z(n5719) );
  XOR U6855 ( .A(n5720), .B(n5719), .Z(n5712) );
  NANDN U6856 ( .A(n5627), .B(n5626), .Z(n5631) );
  NAND U6857 ( .A(n5629), .B(n5628), .Z(n5630) );
  NAND U6858 ( .A(n5631), .B(n5630), .Z(n5711) );
  NANDN U6859 ( .A(n5729), .B(n5632), .Z(n5636) );
  NAND U6860 ( .A(n5634), .B(n5633), .Z(n5635) );
  NAND U6861 ( .A(n5636), .B(n5635), .Z(n5754) );
  AND U6862 ( .A(x[238]), .B(y[1840]), .Z(n6726) );
  NAND U6863 ( .A(n6726), .B(n5637), .Z(n5641) );
  NANDN U6864 ( .A(n5639), .B(n5638), .Z(n5640) );
  AND U6865 ( .A(n5641), .B(n5640), .Z(n5782) );
  AND U6866 ( .A(x[235]), .B(y[1838]), .Z(n5800) );
  AND U6867 ( .A(x[236]), .B(y[1837]), .Z(n5799) );
  NAND U6868 ( .A(x[231]), .B(y[1842]), .Z(n5798) );
  XOR U6869 ( .A(n5799), .B(n5798), .Z(n5801) );
  XOR U6870 ( .A(n5800), .B(n5801), .Z(n5780) );
  NAND U6871 ( .A(x[248]), .B(y[1825]), .Z(n5797) );
  XNOR U6872 ( .A(o[57]), .B(n5797), .Z(n5767) );
  NAND U6873 ( .A(x[225]), .B(y[1848]), .Z(n5768) );
  NAND U6874 ( .A(x[237]), .B(y[1836]), .Z(n5770) );
  XOR U6875 ( .A(n5754), .B(n5753), .Z(n5756) );
  AND U6876 ( .A(n5643), .B(n5642), .Z(n5647) );
  NAND U6877 ( .A(n5645), .B(n5644), .Z(n5646) );
  NANDN U6878 ( .A(n5647), .B(n5646), .Z(n5742) );
  AND U6879 ( .A(n5649), .B(n5648), .Z(n5653) );
  NAND U6880 ( .A(n5651), .B(n5650), .Z(n5652) );
  NANDN U6881 ( .A(n5653), .B(n5652), .Z(n5741) );
  XOR U6882 ( .A(n5742), .B(n5741), .Z(n5744) );
  NAND U6883 ( .A(n5655), .B(n5654), .Z(n5659) );
  NAND U6884 ( .A(n5657), .B(n5656), .Z(n5658) );
  NAND U6885 ( .A(n5659), .B(n5658), .Z(n5738) );
  AND U6886 ( .A(x[232]), .B(y[1841]), .Z(n5732) );
  XOR U6887 ( .A(n5730), .B(n5660), .Z(n5731) );
  XOR U6888 ( .A(n5732), .B(n5731), .Z(n5736) );
  AND U6889 ( .A(n5661), .B(o[56]), .Z(n5725) );
  AND U6890 ( .A(x[249]), .B(y[1824]), .Z(n5724) );
  NAND U6891 ( .A(x[224]), .B(y[1849]), .Z(n5723) );
  XOR U6892 ( .A(n5724), .B(n5723), .Z(n5726) );
  XNOR U6893 ( .A(n5725), .B(n5726), .Z(n5735) );
  XOR U6894 ( .A(n5736), .B(n5735), .Z(n5737) );
  XOR U6895 ( .A(n5738), .B(n5737), .Z(n5743) );
  XOR U6896 ( .A(n5744), .B(n5743), .Z(n5755) );
  XOR U6897 ( .A(n5756), .B(n5755), .Z(n5836) );
  AND U6898 ( .A(n5663), .B(n5662), .Z(n5667) );
  NAND U6899 ( .A(n5665), .B(n5664), .Z(n5666) );
  NANDN U6900 ( .A(n5667), .B(n5666), .Z(n5818) );
  NAND U6901 ( .A(n5669), .B(n5668), .Z(n5673) );
  NAND U6902 ( .A(n5671), .B(n5670), .Z(n5672) );
  NAND U6903 ( .A(n5673), .B(n5672), .Z(n5816) );
  AND U6904 ( .A(x[238]), .B(y[1835]), .Z(n5773) );
  AND U6905 ( .A(x[226]), .B(y[1847]), .Z(n5774) );
  XOR U6906 ( .A(n5773), .B(n5774), .Z(n5775) );
  AND U6907 ( .A(x[227]), .B(y[1846]), .Z(n5776) );
  XOR U6908 ( .A(n5775), .B(n5776), .Z(n5815) );
  XOR U6909 ( .A(n5816), .B(n5815), .Z(n5817) );
  XNOR U6910 ( .A(n5818), .B(n5817), .Z(n5833) );
  NANDN U6911 ( .A(n5675), .B(n5674), .Z(n5679) );
  NAND U6912 ( .A(n5677), .B(n5676), .Z(n5678) );
  AND U6913 ( .A(n5679), .B(n5678), .Z(n5834) );
  XOR U6914 ( .A(n5833), .B(n5834), .Z(n5835) );
  NAND U6915 ( .A(n5681), .B(n5680), .Z(n5685) );
  NAND U6916 ( .A(n5683), .B(n5682), .Z(n5684) );
  AND U6917 ( .A(n5685), .B(n5684), .Z(n5840) );
  XOR U6918 ( .A(n5839), .B(n5840), .Z(n5842) );
  NAND U6919 ( .A(n5687), .B(n5686), .Z(n5691) );
  NAND U6920 ( .A(n5689), .B(n5688), .Z(n5690) );
  AND U6921 ( .A(n5691), .B(n5690), .Z(n5841) );
  XOR U6922 ( .A(n5842), .B(n5841), .Z(n5706) );
  NANDN U6923 ( .A(n5693), .B(n5692), .Z(n5697) );
  NANDN U6924 ( .A(n5695), .B(n5694), .Z(n5696) );
  AND U6925 ( .A(n5697), .B(n5696), .Z(n5705) );
  XOR U6926 ( .A(n5707), .B(n5708), .Z(n5853) );
  NAND U6927 ( .A(n5699), .B(n5698), .Z(n5703) );
  NAND U6928 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U6929 ( .A(n5703), .B(n5702), .Z(n5852) );
  XNOR U6930 ( .A(n5854), .B(n5855), .Z(n5848) );
  XNOR U6931 ( .A(n5847), .B(n5848), .Z(n5704) );
  XOR U6932 ( .A(n5845), .B(n5704), .Z(N122) );
  NANDN U6933 ( .A(n5706), .B(n5705), .Z(n5710) );
  NAND U6934 ( .A(n5708), .B(n5707), .Z(n5709) );
  AND U6935 ( .A(n5710), .B(n5709), .Z(n5860) );
  NANDN U6936 ( .A(n5712), .B(n5711), .Z(n5716) );
  NANDN U6937 ( .A(n5714), .B(n5713), .Z(n5715) );
  AND U6938 ( .A(n5716), .B(n5715), .Z(n5859) );
  NAND U6939 ( .A(n5718), .B(n5717), .Z(n5722) );
  NAND U6940 ( .A(n5720), .B(n5719), .Z(n5721) );
  NAND U6941 ( .A(n5722), .B(n5721), .Z(n5881) );
  AND U6942 ( .A(x[226]), .B(y[1848]), .Z(n5894) );
  XOR U6943 ( .A(n5895), .B(n5894), .Z(n5897) );
  NAND U6944 ( .A(x[248]), .B(y[1826]), .Z(n5896) );
  XNOR U6945 ( .A(n5897), .B(n5896), .Z(n5936) );
  NANDN U6946 ( .A(n5724), .B(n5723), .Z(n5728) );
  OR U6947 ( .A(n5726), .B(n5725), .Z(n5727) );
  NAND U6948 ( .A(n5728), .B(n5727), .Z(n5937) );
  XNOR U6949 ( .A(n5936), .B(n5937), .Z(n5938) );
  NANDN U6950 ( .A(n5730), .B(n5729), .Z(n5734) );
  NANDN U6951 ( .A(n5732), .B(n5731), .Z(n5733) );
  NAND U6952 ( .A(n5734), .B(n5733), .Z(n5939) );
  XOR U6953 ( .A(n5938), .B(n5939), .Z(n5974) );
  NAND U6954 ( .A(n5736), .B(n5735), .Z(n5740) );
  NAND U6955 ( .A(n5738), .B(n5737), .Z(n5739) );
  AND U6956 ( .A(n5740), .B(n5739), .Z(n5975) );
  XOR U6957 ( .A(n5974), .B(n5975), .Z(n5977) );
  NAND U6958 ( .A(n5742), .B(n5741), .Z(n5746) );
  NAND U6959 ( .A(n5744), .B(n5743), .Z(n5745) );
  AND U6960 ( .A(n5746), .B(n5745), .Z(n5976) );
  XOR U6961 ( .A(n5977), .B(n5976), .Z(n5971) );
  NAND U6962 ( .A(n5748), .B(n5747), .Z(n5752) );
  NAND U6963 ( .A(n5750), .B(n5749), .Z(n5751) );
  NAND U6964 ( .A(n5752), .B(n5751), .Z(n5968) );
  NAND U6965 ( .A(n5754), .B(n5753), .Z(n5758) );
  NAND U6966 ( .A(n5756), .B(n5755), .Z(n5757) );
  AND U6967 ( .A(n5758), .B(n5757), .Z(n5969) );
  XOR U6968 ( .A(n5968), .B(n5969), .Z(n5970) );
  XNOR U6969 ( .A(n5971), .B(n5970), .Z(n5879) );
  NAND U6970 ( .A(n5760), .B(n5759), .Z(n5764) );
  NAND U6971 ( .A(n5762), .B(n5761), .Z(n5763) );
  NAND U6972 ( .A(n5764), .B(n5763), .Z(n5964) );
  AND U6973 ( .A(x[236]), .B(y[1838]), .Z(n6086) );
  AND U6974 ( .A(x[229]), .B(y[1845]), .Z(n5951) );
  XOR U6975 ( .A(n6086), .B(n5951), .Z(n5953) );
  NAND U6976 ( .A(x[234]), .B(y[1840]), .Z(n5952) );
  XNOR U6977 ( .A(n5953), .B(n5952), .Z(n5983) );
  AND U6978 ( .A(x[231]), .B(y[1843]), .Z(n5981) );
  AND U6979 ( .A(y[1844]), .B(x[230]), .Z(n5766) );
  NAND U6980 ( .A(y[1842]), .B(x[232]), .Z(n5765) );
  XNOR U6981 ( .A(n5766), .B(n5765), .Z(n5999) );
  NAND U6982 ( .A(x[233]), .B(y[1841]), .Z(n6000) );
  XNOR U6983 ( .A(n5999), .B(n6000), .Z(n5980) );
  XOR U6984 ( .A(n5981), .B(n5980), .Z(n5982) );
  XOR U6985 ( .A(n5983), .B(n5982), .Z(n5920) );
  NANDN U6986 ( .A(n5768), .B(n5767), .Z(n5772) );
  NANDN U6987 ( .A(n5770), .B(n5769), .Z(n5771) );
  NAND U6988 ( .A(n5772), .B(n5771), .Z(n5919) );
  NAND U6989 ( .A(n5774), .B(n5773), .Z(n5778) );
  NAND U6990 ( .A(n5776), .B(n5775), .Z(n5777) );
  NAND U6991 ( .A(n5778), .B(n5777), .Z(n5918) );
  XNOR U6992 ( .A(n5919), .B(n5918), .Z(n5921) );
  NANDN U6993 ( .A(n5780), .B(n5779), .Z(n5784) );
  NANDN U6994 ( .A(n5782), .B(n5781), .Z(n5783) );
  AND U6995 ( .A(n5784), .B(n5783), .Z(n5924) );
  NANDN U6996 ( .A(n5786), .B(n5785), .Z(n5790) );
  NANDN U6997 ( .A(n5788), .B(n5787), .Z(n5789) );
  AND U6998 ( .A(n5790), .B(n5789), .Z(n5884) );
  NANDN U6999 ( .A(n5792), .B(n5791), .Z(n5796) );
  NANDN U7000 ( .A(n5794), .B(n5793), .Z(n5795) );
  NAND U7001 ( .A(n5796), .B(n5795), .Z(n5885) );
  XNOR U7002 ( .A(n5884), .B(n5885), .Z(n5886) );
  ANDN U7003 ( .B(o[57]), .A(n5797), .Z(n5992) );
  NAND U7004 ( .A(x[238]), .B(y[1836]), .Z(n5993) );
  XNOR U7005 ( .A(n5992), .B(n5993), .Z(n5994) );
  NAND U7006 ( .A(x[225]), .B(y[1849]), .Z(n5995) );
  XNOR U7007 ( .A(n5994), .B(n5995), .Z(n5942) );
  NAND U7008 ( .A(x[249]), .B(y[1825]), .Z(n6003) );
  XNOR U7009 ( .A(o[58]), .B(n6003), .Z(n5956) );
  NAND U7010 ( .A(x[250]), .B(y[1824]), .Z(n5957) );
  XNOR U7011 ( .A(n5956), .B(n5957), .Z(n5958) );
  NAND U7012 ( .A(x[224]), .B(y[1850]), .Z(n5959) );
  XOR U7013 ( .A(n5958), .B(n5959), .Z(n5943) );
  XNOR U7014 ( .A(n5942), .B(n5943), .Z(n5944) );
  NANDN U7015 ( .A(n5799), .B(n5798), .Z(n5803) );
  OR U7016 ( .A(n5801), .B(n5800), .Z(n5802) );
  NAND U7017 ( .A(n5803), .B(n5802), .Z(n5945) );
  XOR U7018 ( .A(n5944), .B(n5945), .Z(n5887) );
  XOR U7019 ( .A(n5886), .B(n5887), .Z(n5932) );
  AND U7020 ( .A(x[245]), .B(y[1829]), .Z(n5986) );
  NAND U7021 ( .A(n5986), .B(n5804), .Z(n5808) );
  NAND U7022 ( .A(n5806), .B(n5805), .Z(n5807) );
  NAND U7023 ( .A(n5808), .B(n5807), .Z(n5914) );
  XOR U7024 ( .A(n5987), .B(n5986), .Z(n5989) );
  NAND U7025 ( .A(x[244]), .B(y[1830]), .Z(n5988) );
  XNOR U7026 ( .A(n5989), .B(n5988), .Z(n5913) );
  NAND U7027 ( .A(x[247]), .B(y[1827]), .Z(n5901) );
  XNOR U7028 ( .A(n5900), .B(n5901), .Z(n5903) );
  AND U7029 ( .A(x[246]), .B(y[1828]), .Z(n5902) );
  XOR U7030 ( .A(n5903), .B(n5902), .Z(n5912) );
  XOR U7031 ( .A(n5913), .B(n5912), .Z(n5915) );
  XOR U7032 ( .A(n5914), .B(n5915), .Z(n5931) );
  AND U7033 ( .A(x[243]), .B(y[1831]), .Z(n6004) );
  NAND U7034 ( .A(x[227]), .B(y[1847]), .Z(n6005) );
  XNOR U7035 ( .A(n6004), .B(n6005), .Z(n6006) );
  NAND U7036 ( .A(x[235]), .B(y[1839]), .Z(n6007) );
  XNOR U7037 ( .A(n6006), .B(n6007), .Z(n5891) );
  AND U7038 ( .A(x[228]), .B(y[1846]), .Z(n5906) );
  XOR U7039 ( .A(n5907), .B(n5906), .Z(n5909) );
  XOR U7040 ( .A(n5891), .B(n5890), .Z(n5892) );
  NANDN U7041 ( .A(n5810), .B(n5809), .Z(n5814) );
  NANDN U7042 ( .A(n5812), .B(n5811), .Z(n5813) );
  NAND U7043 ( .A(n5814), .B(n5813), .Z(n5893) );
  XOR U7044 ( .A(n5892), .B(n5893), .Z(n5930) );
  XOR U7045 ( .A(n5932), .B(n5933), .Z(n5927) );
  XNOR U7046 ( .A(n5926), .B(n5927), .Z(n5963) );
  NAND U7047 ( .A(n5816), .B(n5815), .Z(n5820) );
  NAND U7048 ( .A(n5818), .B(n5817), .Z(n5819) );
  NAND U7049 ( .A(n5820), .B(n5819), .Z(n6014) );
  NAND U7050 ( .A(n5822), .B(n5821), .Z(n5826) );
  NAND U7051 ( .A(n5824), .B(n5823), .Z(n5825) );
  NAND U7052 ( .A(n5826), .B(n5825), .Z(n6013) );
  NAND U7053 ( .A(n5828), .B(n5827), .Z(n5832) );
  NANDN U7054 ( .A(n5830), .B(n5829), .Z(n5831) );
  NAND U7055 ( .A(n5832), .B(n5831), .Z(n6012) );
  XOR U7056 ( .A(n6013), .B(n6012), .Z(n6015) );
  XOR U7057 ( .A(n6014), .B(n6015), .Z(n5962) );
  XOR U7058 ( .A(n5964), .B(n5965), .Z(n5878) );
  XOR U7059 ( .A(n5879), .B(n5878), .Z(n5880) );
  XOR U7060 ( .A(n5881), .B(n5880), .Z(n5875) );
  NAND U7061 ( .A(n5834), .B(n5833), .Z(n5838) );
  NANDN U7062 ( .A(n5836), .B(n5835), .Z(n5837) );
  AND U7063 ( .A(n5838), .B(n5837), .Z(n5872) );
  NAND U7064 ( .A(n5840), .B(n5839), .Z(n5844) );
  NAND U7065 ( .A(n5842), .B(n5841), .Z(n5843) );
  AND U7066 ( .A(n5844), .B(n5843), .Z(n5873) );
  XOR U7067 ( .A(n5872), .B(n5873), .Z(n5874) );
  XOR U7068 ( .A(n5875), .B(n5874), .Z(n5861) );
  XNOR U7069 ( .A(n5862), .B(n5861), .Z(n5868) );
  OR U7070 ( .A(n5847), .B(n5845), .Z(n5851) );
  ANDN U7071 ( .B(n5847), .A(n5846), .Z(n5849) );
  OR U7072 ( .A(n5849), .B(n5848), .Z(n5850) );
  AND U7073 ( .A(n5851), .B(n5850), .Z(n5867) );
  NANDN U7074 ( .A(n5853), .B(n5852), .Z(n5857) );
  NANDN U7075 ( .A(n5855), .B(n5854), .Z(n5856) );
  AND U7076 ( .A(n5857), .B(n5856), .Z(n5866) );
  IV U7077 ( .A(n5866), .Z(n5865) );
  XOR U7078 ( .A(n5867), .B(n5865), .Z(n5858) );
  XNOR U7079 ( .A(n5868), .B(n5858), .Z(N123) );
  NANDN U7080 ( .A(n5860), .B(n5859), .Z(n5864) );
  NAND U7081 ( .A(n5862), .B(n5861), .Z(n5863) );
  NAND U7082 ( .A(n5864), .B(n5863), .Z(n6026) );
  IV U7083 ( .A(n6026), .Z(n6025) );
  OR U7084 ( .A(n5867), .B(n5865), .Z(n5871) );
  ANDN U7085 ( .B(n5867), .A(n5866), .Z(n5869) );
  OR U7086 ( .A(n5869), .B(n5868), .Z(n5870) );
  AND U7087 ( .A(n5871), .B(n5870), .Z(n6027) );
  NAND U7088 ( .A(n5873), .B(n5872), .Z(n5877) );
  NAND U7089 ( .A(n5875), .B(n5874), .Z(n5876) );
  AND U7090 ( .A(n5877), .B(n5876), .Z(n6022) );
  NAND U7091 ( .A(n5879), .B(n5878), .Z(n5883) );
  NAND U7092 ( .A(n5881), .B(n5880), .Z(n5882) );
  AND U7093 ( .A(n5883), .B(n5882), .Z(n6020) );
  NANDN U7094 ( .A(n5885), .B(n5884), .Z(n5889) );
  NANDN U7095 ( .A(n5887), .B(n5886), .Z(n5888) );
  AND U7096 ( .A(n5889), .B(n5888), .Z(n6158) );
  NAND U7097 ( .A(n5895), .B(n5894), .Z(n5899) );
  ANDN U7098 ( .B(n5897), .A(n5896), .Z(n5898) );
  ANDN U7099 ( .B(n5899), .A(n5898), .Z(n6057) );
  NANDN U7100 ( .A(n5901), .B(n5900), .Z(n5905) );
  NAND U7101 ( .A(n5903), .B(n5902), .Z(n5904) );
  NAND U7102 ( .A(n5905), .B(n5904), .Z(n6056) );
  XNOR U7103 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U7104 ( .A(n5907), .B(n5906), .Z(n5911) );
  ANDN U7105 ( .B(n5909), .A(n5908), .Z(n5910) );
  ANDN U7106 ( .B(n5911), .A(n5910), .Z(n6071) );
  AND U7107 ( .A(x[224]), .B(y[1851]), .Z(n6143) );
  NAND U7108 ( .A(x[251]), .B(y[1824]), .Z(n6144) );
  XNOR U7109 ( .A(n6143), .B(n6144), .Z(n6145) );
  NAND U7110 ( .A(x[250]), .B(y[1825]), .Z(n6134) );
  XOR U7111 ( .A(o[59]), .B(n6134), .Z(n6146) );
  XNOR U7112 ( .A(n6145), .B(n6146), .Z(n6068) );
  AND U7113 ( .A(x[233]), .B(y[1842]), .Z(n6128) );
  NAND U7114 ( .A(x[245]), .B(y[1830]), .Z(n6129) );
  XNOR U7115 ( .A(n6128), .B(n6129), .Z(n6130) );
  NAND U7116 ( .A(x[242]), .B(y[1833]), .Z(n6131) );
  XOR U7117 ( .A(n6130), .B(n6131), .Z(n6069) );
  XNOR U7118 ( .A(n6068), .B(n6069), .Z(n6070) );
  XOR U7119 ( .A(n6071), .B(n6070), .Z(n6059) );
  XNOR U7120 ( .A(n6058), .B(n6059), .Z(n6155) );
  XNOR U7121 ( .A(n6156), .B(n6155), .Z(n6157) );
  XOR U7122 ( .A(n6158), .B(n6157), .Z(n6175) );
  NAND U7123 ( .A(n5913), .B(n5912), .Z(n5917) );
  NAND U7124 ( .A(n5915), .B(n5914), .Z(n5916) );
  AND U7125 ( .A(n5917), .B(n5916), .Z(n6174) );
  NAND U7126 ( .A(n5919), .B(n5918), .Z(n5923) );
  NANDN U7127 ( .A(n5921), .B(n5920), .Z(n5922) );
  AND U7128 ( .A(n5923), .B(n5922), .Z(n6173) );
  XOR U7129 ( .A(n6174), .B(n6173), .Z(n6176) );
  XOR U7130 ( .A(n6175), .B(n6176), .Z(n6033) );
  NANDN U7131 ( .A(n5925), .B(n5924), .Z(n5929) );
  NANDN U7132 ( .A(n5927), .B(n5926), .Z(n5928) );
  AND U7133 ( .A(n5929), .B(n5928), .Z(n6164) );
  NANDN U7134 ( .A(n5931), .B(n5930), .Z(n5935) );
  NANDN U7135 ( .A(n5933), .B(n5932), .Z(n5934) );
  AND U7136 ( .A(n5935), .B(n5934), .Z(n6162) );
  NANDN U7137 ( .A(n5937), .B(n5936), .Z(n5941) );
  NANDN U7138 ( .A(n5939), .B(n5938), .Z(n5940) );
  AND U7139 ( .A(n5941), .B(n5940), .Z(n6152) );
  NANDN U7140 ( .A(n5943), .B(n5942), .Z(n5947) );
  NANDN U7141 ( .A(n5945), .B(n5944), .Z(n5946) );
  AND U7142 ( .A(n5947), .B(n5946), .Z(n6150) );
  AND U7143 ( .A(x[243]), .B(y[1832]), .Z(n6122) );
  NAND U7144 ( .A(x[249]), .B(y[1826]), .Z(n6123) );
  XNOR U7145 ( .A(n6122), .B(n6123), .Z(n6124) );
  NAND U7146 ( .A(x[230]), .B(y[1845]), .Z(n6125) );
  XNOR U7147 ( .A(n6124), .B(n6125), .Z(n6111) );
  AND U7148 ( .A(x[239]), .B(y[1836]), .Z(n6091) );
  NAND U7149 ( .A(x[226]), .B(y[1849]), .Z(n6092) );
  NAND U7150 ( .A(x[227]), .B(y[1848]), .Z(n6094) );
  XNOR U7151 ( .A(n6111), .B(n6112), .Z(n6113) );
  NAND U7152 ( .A(x[240]), .B(y[1835]), .Z(n6074) );
  XNOR U7153 ( .A(n6074), .B(n6075), .Z(n6076) );
  XNOR U7154 ( .A(n5948), .B(n6076), .Z(n6087) );
  AND U7155 ( .A(y[1838]), .B(x[237]), .Z(n5950) );
  NAND U7156 ( .A(y[1839]), .B(x[236]), .Z(n5949) );
  XNOR U7157 ( .A(n5950), .B(n5949), .Z(n6088) );
  XNOR U7158 ( .A(n6087), .B(n6088), .Z(n6114) );
  XNOR U7159 ( .A(n6113), .B(n6114), .Z(n6052) );
  NAND U7160 ( .A(n6086), .B(n5951), .Z(n5955) );
  ANDN U7161 ( .B(n5953), .A(n5952), .Z(n5954) );
  ANDN U7162 ( .B(n5955), .A(n5954), .Z(n6051) );
  NANDN U7163 ( .A(n5957), .B(n5956), .Z(n5961) );
  NANDN U7164 ( .A(n5959), .B(n5958), .Z(n5960) );
  NAND U7165 ( .A(n5961), .B(n5960), .Z(n6050) );
  XOR U7166 ( .A(n6051), .B(n6050), .Z(n6053) );
  XNOR U7167 ( .A(n6052), .B(n6053), .Z(n6149) );
  XNOR U7168 ( .A(n6150), .B(n6149), .Z(n6151) );
  XNOR U7169 ( .A(n6152), .B(n6151), .Z(n6161) );
  XOR U7170 ( .A(n6162), .B(n6161), .Z(n6163) );
  XOR U7171 ( .A(n6164), .B(n6163), .Z(n6032) );
  NANDN U7172 ( .A(n5963), .B(n5962), .Z(n5967) );
  NAND U7173 ( .A(n5965), .B(n5964), .Z(n5966) );
  NAND U7174 ( .A(n5967), .B(n5966), .Z(n6034) );
  XOR U7175 ( .A(n6035), .B(n6034), .Z(n6041) );
  NAND U7176 ( .A(n5969), .B(n5968), .Z(n5973) );
  NAND U7177 ( .A(n5971), .B(n5970), .Z(n5972) );
  NAND U7178 ( .A(n5973), .B(n5972), .Z(n6038) );
  NAND U7179 ( .A(n5975), .B(n5974), .Z(n5979) );
  NAND U7180 ( .A(n5977), .B(n5976), .Z(n5978) );
  NAND U7181 ( .A(n5979), .B(n5978), .Z(n6045) );
  NAND U7182 ( .A(n5981), .B(n5980), .Z(n5985) );
  NAND U7183 ( .A(n5983), .B(n5982), .Z(n5984) );
  NAND U7184 ( .A(n5985), .B(n5984), .Z(n6169) );
  NAND U7185 ( .A(n5987), .B(n5986), .Z(n5991) );
  ANDN U7186 ( .B(n5989), .A(n5988), .Z(n5990) );
  ANDN U7187 ( .B(n5991), .A(n5990), .Z(n6104) );
  NANDN U7188 ( .A(n5993), .B(n5992), .Z(n5997) );
  NANDN U7189 ( .A(n5995), .B(n5994), .Z(n5996) );
  NAND U7190 ( .A(n5997), .B(n5996), .Z(n6103) );
  XNOR U7191 ( .A(n6104), .B(n6103), .Z(n6106) );
  AND U7192 ( .A(y[1844]), .B(x[232]), .Z(n6136) );
  NAND U7193 ( .A(n5998), .B(n6136), .Z(n6002) );
  NANDN U7194 ( .A(n6000), .B(n5999), .Z(n6001) );
  NAND U7195 ( .A(n6002), .B(n6001), .Z(n6064) );
  AND U7196 ( .A(x[238]), .B(y[1837]), .Z(n6097) );
  NAND U7197 ( .A(x[225]), .B(y[1850]), .Z(n6098) );
  ANDN U7198 ( .B(o[58]), .A(n6003), .Z(n6099) );
  XOR U7199 ( .A(n6100), .B(n6099), .Z(n6063) );
  AND U7200 ( .A(x[241]), .B(y[1834]), .Z(n6137) );
  NAND U7201 ( .A(x[228]), .B(y[1847]), .Z(n6138) );
  XNOR U7202 ( .A(n6137), .B(n6138), .Z(n6140) );
  AND U7203 ( .A(x[229]), .B(y[1846]), .Z(n6139) );
  XOR U7204 ( .A(n6140), .B(n6139), .Z(n6062) );
  XOR U7205 ( .A(n6063), .B(n6062), .Z(n6065) );
  XOR U7206 ( .A(n6064), .B(n6065), .Z(n6105) );
  XOR U7207 ( .A(n6106), .B(n6105), .Z(n6168) );
  NANDN U7208 ( .A(n6005), .B(n6004), .Z(n6009) );
  NANDN U7209 ( .A(n6007), .B(n6006), .Z(n6008) );
  AND U7210 ( .A(n6009), .B(n6008), .Z(n6110) );
  AND U7211 ( .A(y[1827]), .B(x[248]), .Z(n6011) );
  NAND U7212 ( .A(y[1831]), .B(x[244]), .Z(n6010) );
  XNOR U7213 ( .A(n6011), .B(n6010), .Z(n6118) );
  NAND U7214 ( .A(x[231]), .B(y[1844]), .Z(n6119) );
  XNOR U7215 ( .A(n6118), .B(n6119), .Z(n6108) );
  AND U7216 ( .A(x[232]), .B(y[1843]), .Z(n6080) );
  AND U7217 ( .A(x[247]), .B(y[1828]), .Z(n6081) );
  XOR U7218 ( .A(n6080), .B(n6081), .Z(n6082) );
  AND U7219 ( .A(x[246]), .B(y[1829]), .Z(n6083) );
  XOR U7220 ( .A(n6082), .B(n6083), .Z(n6107) );
  XOR U7221 ( .A(n6108), .B(n6107), .Z(n6109) );
  XNOR U7222 ( .A(n6110), .B(n6109), .Z(n6167) );
  XOR U7223 ( .A(n6168), .B(n6167), .Z(n6170) );
  XNOR U7224 ( .A(n6169), .B(n6170), .Z(n6044) );
  XOR U7225 ( .A(n6045), .B(n6044), .Z(n6047) );
  NAND U7226 ( .A(n6013), .B(n6012), .Z(n6017) );
  NAND U7227 ( .A(n6015), .B(n6014), .Z(n6016) );
  AND U7228 ( .A(n6017), .B(n6016), .Z(n6046) );
  XOR U7229 ( .A(n6047), .B(n6046), .Z(n6039) );
  XOR U7230 ( .A(n6038), .B(n6039), .Z(n6040) );
  XOR U7231 ( .A(n6020), .B(n6019), .Z(n6021) );
  XOR U7232 ( .A(n6022), .B(n6021), .Z(n6028) );
  XNOR U7233 ( .A(n6027), .B(n6028), .Z(n6018) );
  XOR U7234 ( .A(n6025), .B(n6018), .Z(N124) );
  NAND U7235 ( .A(n6020), .B(n6019), .Z(n6024) );
  NAND U7236 ( .A(n6022), .B(n6021), .Z(n6023) );
  NAND U7237 ( .A(n6024), .B(n6023), .Z(n6188) );
  IV U7238 ( .A(n6188), .Z(n6186) );
  OR U7239 ( .A(n6027), .B(n6025), .Z(n6031) );
  ANDN U7240 ( .B(n6027), .A(n6026), .Z(n6029) );
  OR U7241 ( .A(n6029), .B(n6028), .Z(n6030) );
  AND U7242 ( .A(n6031), .B(n6030), .Z(n6187) );
  NANDN U7243 ( .A(n6033), .B(n6032), .Z(n6037) );
  NAND U7244 ( .A(n6035), .B(n6034), .Z(n6036) );
  NAND U7245 ( .A(n6037), .B(n6036), .Z(n6180) );
  NAND U7246 ( .A(n6039), .B(n6038), .Z(n6043) );
  NANDN U7247 ( .A(n6041), .B(n6040), .Z(n6042) );
  AND U7248 ( .A(n6043), .B(n6042), .Z(n6181) );
  XOR U7249 ( .A(n6180), .B(n6181), .Z(n6183) );
  NAND U7250 ( .A(n6045), .B(n6044), .Z(n6049) );
  NAND U7251 ( .A(n6047), .B(n6046), .Z(n6048) );
  AND U7252 ( .A(n6049), .B(n6048), .Z(n6194) );
  NANDN U7253 ( .A(n6051), .B(n6050), .Z(n6055) );
  NANDN U7254 ( .A(n6053), .B(n6052), .Z(n6054) );
  AND U7255 ( .A(n6055), .B(n6054), .Z(n6218) );
  NANDN U7256 ( .A(n6057), .B(n6056), .Z(n6061) );
  NANDN U7257 ( .A(n6059), .B(n6058), .Z(n6060) );
  AND U7258 ( .A(n6061), .B(n6060), .Z(n6324) );
  NAND U7259 ( .A(n6063), .B(n6062), .Z(n6067) );
  NAND U7260 ( .A(n6065), .B(n6064), .Z(n6066) );
  AND U7261 ( .A(n6067), .B(n6066), .Z(n6322) );
  NANDN U7262 ( .A(n6069), .B(n6068), .Z(n6073) );
  NANDN U7263 ( .A(n6071), .B(n6070), .Z(n6072) );
  NAND U7264 ( .A(n6073), .B(n6072), .Z(n6321) );
  XNOR U7265 ( .A(n6322), .B(n6321), .Z(n6323) );
  XNOR U7266 ( .A(n6324), .B(n6323), .Z(n6217) );
  XNOR U7267 ( .A(n6218), .B(n6217), .Z(n6220) );
  NANDN U7268 ( .A(n6075), .B(n6074), .Z(n6079) );
  NANDN U7269 ( .A(n6077), .B(n6076), .Z(n6078) );
  AND U7270 ( .A(n6079), .B(n6078), .Z(n6285) );
  AND U7271 ( .A(x[239]), .B(y[1837]), .Z(n6297) );
  NAND U7272 ( .A(x[251]), .B(y[1825]), .Z(n6281) );
  AND U7273 ( .A(x[250]), .B(y[1826]), .Z(n6294) );
  XOR U7274 ( .A(n6295), .B(n6294), .Z(n6296) );
  XOR U7275 ( .A(n6297), .B(n6296), .Z(n6283) );
  AND U7276 ( .A(x[231]), .B(y[1845]), .Z(n6264) );
  NAND U7277 ( .A(x[236]), .B(y[1840]), .Z(n6265) );
  AND U7278 ( .A(x[235]), .B(y[1841]), .Z(n6266) );
  XNOR U7279 ( .A(n6267), .B(n6266), .Z(n6282) );
  AND U7280 ( .A(x[241]), .B(y[1835]), .Z(n6230) );
  AND U7281 ( .A(x[246]), .B(y[1830]), .Z(n6229) );
  XOR U7282 ( .A(n6230), .B(n6229), .Z(n6232) );
  AND U7283 ( .A(x[228]), .B(y[1848]), .Z(n6231) );
  XOR U7284 ( .A(n6232), .B(n6231), .Z(n6304) );
  AND U7285 ( .A(x[230]), .B(y[1846]), .Z(n6461) );
  NAND U7286 ( .A(x[243]), .B(y[1833]), .Z(n6270) );
  XOR U7287 ( .A(n6304), .B(n6303), .Z(n6305) );
  NAND U7288 ( .A(n6081), .B(n6080), .Z(n6085) );
  NAND U7289 ( .A(n6083), .B(n6082), .Z(n6084) );
  AND U7290 ( .A(n6085), .B(n6084), .Z(n6306) );
  XOR U7291 ( .A(n6328), .B(n6327), .Z(n6329) );
  NAND U7292 ( .A(n6289), .B(n6086), .Z(n6090) );
  NAND U7293 ( .A(n6088), .B(n6087), .Z(n6089) );
  AND U7294 ( .A(n6090), .B(n6089), .Z(n6249) );
  NANDN U7295 ( .A(n6092), .B(n6091), .Z(n6096) );
  NANDN U7296 ( .A(n6094), .B(n6093), .Z(n6095) );
  AND U7297 ( .A(n6096), .B(n6095), .Z(n6247) );
  NANDN U7298 ( .A(n6098), .B(n6097), .Z(n6102) );
  NAND U7299 ( .A(n6100), .B(n6099), .Z(n6101) );
  NAND U7300 ( .A(n6102), .B(n6101), .Z(n6246) );
  XNOR U7301 ( .A(n6329), .B(n6330), .Z(n6219) );
  XOR U7302 ( .A(n6220), .B(n6219), .Z(n6213) );
  NANDN U7303 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U7304 ( .A(n6114), .B(n6113), .Z(n6115) );
  NAND U7305 ( .A(n6116), .B(n6115), .Z(n6309) );
  XOR U7306 ( .A(n6310), .B(n6309), .Z(n6312) );
  XOR U7307 ( .A(n6311), .B(n6312), .Z(n6212) );
  AND U7308 ( .A(x[248]), .B(y[1831]), .Z(n6592) );
  AND U7309 ( .A(x[244]), .B(y[1827]), .Z(n6117) );
  NAND U7310 ( .A(n6592), .B(n6117), .Z(n6121) );
  NANDN U7311 ( .A(n6119), .B(n6118), .Z(n6120) );
  AND U7312 ( .A(n6121), .B(n6120), .Z(n6348) );
  AND U7313 ( .A(x[249]), .B(y[1827]), .Z(n6260) );
  XOR U7314 ( .A(n6261), .B(n6260), .Z(n6259) );
  AND U7315 ( .A(x[225]), .B(y[1851]), .Z(n6258) );
  XOR U7316 ( .A(n6259), .B(n6258), .Z(n6346) );
  AND U7317 ( .A(x[240]), .B(y[1836]), .Z(n6253) );
  AND U7318 ( .A(x[248]), .B(y[1828]), .Z(n6252) );
  XOR U7319 ( .A(n6253), .B(n6252), .Z(n6255) );
  AND U7320 ( .A(x[226]), .B(y[1850]), .Z(n6254) );
  XOR U7321 ( .A(n6255), .B(n6254), .Z(n6345) );
  XOR U7322 ( .A(n6346), .B(n6345), .Z(n6347) );
  NANDN U7323 ( .A(n6123), .B(n6122), .Z(n6127) );
  NANDN U7324 ( .A(n6125), .B(n6124), .Z(n6126) );
  AND U7325 ( .A(n6127), .B(n6126), .Z(n6342) );
  AND U7326 ( .A(x[227]), .B(y[1849]), .Z(n6288) );
  XOR U7327 ( .A(n6289), .B(n6288), .Z(n6291) );
  AND U7328 ( .A(x[247]), .B(y[1829]), .Z(n6290) );
  XOR U7329 ( .A(n6291), .B(n6290), .Z(n6340) );
  AND U7330 ( .A(x[229]), .B(y[1847]), .Z(n6276) );
  AND U7331 ( .A(x[245]), .B(y[1831]), .Z(n6275) );
  XOR U7332 ( .A(n6276), .B(n6275), .Z(n6278) );
  AND U7333 ( .A(x[244]), .B(y[1832]), .Z(n6277) );
  XOR U7334 ( .A(n6278), .B(n6277), .Z(n6339) );
  XOR U7335 ( .A(n6340), .B(n6339), .Z(n6341) );
  NANDN U7336 ( .A(n6129), .B(n6128), .Z(n6133) );
  NANDN U7337 ( .A(n6131), .B(n6130), .Z(n6132) );
  NAND U7338 ( .A(n6133), .B(n6132), .Z(n6225) );
  AND U7339 ( .A(x[224]), .B(y[1852]), .Z(n6236) );
  AND U7340 ( .A(x[252]), .B(y[1824]), .Z(n6235) );
  XOR U7341 ( .A(n6236), .B(n6235), .Z(n6238) );
  ANDN U7342 ( .B(o[59]), .A(n6134), .Z(n6237) );
  XOR U7343 ( .A(n6238), .B(n6237), .Z(n6224) );
  NAND U7344 ( .A(y[1842]), .B(x[234]), .Z(n6135) );
  XNOR U7345 ( .A(n6136), .B(n6135), .Z(n6243) );
  AND U7346 ( .A(x[233]), .B(y[1843]), .Z(n6242) );
  XOR U7347 ( .A(n6243), .B(n6242), .Z(n6223) );
  XOR U7348 ( .A(n6224), .B(n6223), .Z(n6226) );
  XOR U7349 ( .A(n6225), .B(n6226), .Z(n6336) );
  NANDN U7350 ( .A(n6138), .B(n6137), .Z(n6142) );
  NAND U7351 ( .A(n6140), .B(n6139), .Z(n6141) );
  AND U7352 ( .A(n6142), .B(n6141), .Z(n6334) );
  NANDN U7353 ( .A(n6144), .B(n6143), .Z(n6148) );
  NANDN U7354 ( .A(n6146), .B(n6145), .Z(n6147) );
  NAND U7355 ( .A(n6148), .B(n6147), .Z(n6333) );
  XNOR U7356 ( .A(n6336), .B(n6335), .Z(n6315) );
  XOR U7357 ( .A(n6316), .B(n6315), .Z(n6317) );
  XOR U7358 ( .A(n6318), .B(n6317), .Z(n6211) );
  XOR U7359 ( .A(n6212), .B(n6211), .Z(n6214) );
  XOR U7360 ( .A(n6213), .B(n6214), .Z(n6207) );
  NANDN U7361 ( .A(n6150), .B(n6149), .Z(n6154) );
  NANDN U7362 ( .A(n6152), .B(n6151), .Z(n6153) );
  AND U7363 ( .A(n6154), .B(n6153), .Z(n6206) );
  NANDN U7364 ( .A(n6156), .B(n6155), .Z(n6160) );
  NANDN U7365 ( .A(n6158), .B(n6157), .Z(n6159) );
  NAND U7366 ( .A(n6160), .B(n6159), .Z(n6205) );
  XOR U7367 ( .A(n6206), .B(n6205), .Z(n6208) );
  XOR U7368 ( .A(n6207), .B(n6208), .Z(n6193) );
  XOR U7369 ( .A(n6194), .B(n6193), .Z(n6196) );
  NAND U7370 ( .A(n6162), .B(n6161), .Z(n6166) );
  NAND U7371 ( .A(n6164), .B(n6163), .Z(n6165) );
  NAND U7372 ( .A(n6166), .B(n6165), .Z(n6201) );
  NAND U7373 ( .A(n6168), .B(n6167), .Z(n6172) );
  NAND U7374 ( .A(n6170), .B(n6169), .Z(n6171) );
  NAND U7375 ( .A(n6172), .B(n6171), .Z(n6199) );
  NAND U7376 ( .A(n6174), .B(n6173), .Z(n6178) );
  NAND U7377 ( .A(n6176), .B(n6175), .Z(n6177) );
  AND U7378 ( .A(n6178), .B(n6177), .Z(n6200) );
  XOR U7379 ( .A(n6199), .B(n6200), .Z(n6202) );
  XOR U7380 ( .A(n6201), .B(n6202), .Z(n6195) );
  XOR U7381 ( .A(n6196), .B(n6195), .Z(n6182) );
  XOR U7382 ( .A(n6183), .B(n6182), .Z(n6189) );
  XNOR U7383 ( .A(n6187), .B(n6189), .Z(n6179) );
  XOR U7384 ( .A(n6186), .B(n6179), .Z(N125) );
  NAND U7385 ( .A(n6181), .B(n6180), .Z(n6185) );
  NAND U7386 ( .A(n6183), .B(n6182), .Z(n6184) );
  AND U7387 ( .A(n6185), .B(n6184), .Z(n6352) );
  NANDN U7388 ( .A(n6186), .B(n6187), .Z(n6192) );
  NOR U7389 ( .A(n6188), .B(n6187), .Z(n6190) );
  OR U7390 ( .A(n6190), .B(n6189), .Z(n6191) );
  AND U7391 ( .A(n6192), .B(n6191), .Z(n6353) );
  NAND U7392 ( .A(n6194), .B(n6193), .Z(n6198) );
  NAND U7393 ( .A(n6196), .B(n6195), .Z(n6197) );
  NAND U7394 ( .A(n6198), .B(n6197), .Z(n6357) );
  NAND U7395 ( .A(n6200), .B(n6199), .Z(n6204) );
  NAND U7396 ( .A(n6202), .B(n6201), .Z(n6203) );
  NAND U7397 ( .A(n6204), .B(n6203), .Z(n6355) );
  NANDN U7398 ( .A(n6206), .B(n6205), .Z(n6210) );
  OR U7399 ( .A(n6208), .B(n6207), .Z(n6209) );
  AND U7400 ( .A(n6210), .B(n6209), .Z(n6362) );
  NANDN U7401 ( .A(n6212), .B(n6211), .Z(n6216) );
  OR U7402 ( .A(n6214), .B(n6213), .Z(n6215) );
  AND U7403 ( .A(n6216), .B(n6215), .Z(n6361) );
  XNOR U7404 ( .A(n6362), .B(n6361), .Z(n6364) );
  NANDN U7405 ( .A(n6218), .B(n6217), .Z(n6222) );
  NAND U7406 ( .A(n6220), .B(n6219), .Z(n6221) );
  AND U7407 ( .A(n6222), .B(n6221), .Z(n6372) );
  NAND U7408 ( .A(n6224), .B(n6223), .Z(n6228) );
  NAND U7409 ( .A(n6226), .B(n6225), .Z(n6227) );
  AND U7410 ( .A(n6228), .B(n6227), .Z(n6481) );
  NAND U7411 ( .A(n6230), .B(n6229), .Z(n6234) );
  NAND U7412 ( .A(n6232), .B(n6231), .Z(n6233) );
  NAND U7413 ( .A(n6234), .B(n6233), .Z(n6518) );
  NAND U7414 ( .A(n6236), .B(n6235), .Z(n6240) );
  NAND U7415 ( .A(n6238), .B(n6237), .Z(n6239) );
  NAND U7416 ( .A(n6240), .B(n6239), .Z(n6517) );
  XOR U7417 ( .A(n6518), .B(n6517), .Z(n6519) );
  AND U7418 ( .A(y[1844]), .B(x[234]), .Z(n6515) );
  NAND U7419 ( .A(n6241), .B(n6515), .Z(n6245) );
  NAND U7420 ( .A(n6243), .B(n6242), .Z(n6244) );
  NAND U7421 ( .A(n6245), .B(n6244), .Z(n6489) );
  AND U7422 ( .A(x[246]), .B(y[1831]), .Z(n6439) );
  AND U7423 ( .A(x[236]), .B(y[1841]), .Z(n6559) );
  AND U7424 ( .A(x[225]), .B(y[1852]), .Z(n6437) );
  XOR U7425 ( .A(n6559), .B(n6437), .Z(n6438) );
  XOR U7426 ( .A(n6439), .B(n6438), .Z(n6488) );
  AND U7427 ( .A(x[239]), .B(y[1838]), .Z(n6442) );
  XOR U7428 ( .A(n6488), .B(n6487), .Z(n6490) );
  XNOR U7429 ( .A(n6489), .B(n6490), .Z(n6520) );
  NANDN U7430 ( .A(n6247), .B(n6246), .Z(n6251) );
  NANDN U7431 ( .A(n6249), .B(n6248), .Z(n6250) );
  AND U7432 ( .A(n6251), .B(n6250), .Z(n6483) );
  XOR U7433 ( .A(n6484), .B(n6483), .Z(n6478) );
  NAND U7434 ( .A(n6253), .B(n6252), .Z(n6257) );
  NAND U7435 ( .A(n6255), .B(n6254), .Z(n6256) );
  NAND U7436 ( .A(n6257), .B(n6256), .Z(n6494) );
  AND U7437 ( .A(n6259), .B(n6258), .Z(n6263) );
  NAND U7438 ( .A(n6261), .B(n6260), .Z(n6262) );
  NANDN U7439 ( .A(n6263), .B(n6262), .Z(n6493) );
  XOR U7440 ( .A(n6494), .B(n6493), .Z(n6496) );
  NANDN U7441 ( .A(n6265), .B(n6264), .Z(n6269) );
  NAND U7442 ( .A(n6267), .B(n6266), .Z(n6268) );
  NAND U7443 ( .A(n6269), .B(n6268), .Z(n6403) );
  AND U7444 ( .A(x[235]), .B(y[1842]), .Z(n6458) );
  AND U7445 ( .A(x[227]), .B(y[1850]), .Z(n6456) );
  AND U7446 ( .A(x[241]), .B(y[1836]), .Z(n6455) );
  XOR U7447 ( .A(n6456), .B(n6455), .Z(n6457) );
  XOR U7448 ( .A(n6458), .B(n6457), .Z(n6402) );
  AND U7449 ( .A(x[247]), .B(y[1830]), .Z(n6452) );
  AND U7450 ( .A(x[237]), .B(y[1840]), .Z(n6450) );
  AND U7451 ( .A(x[248]), .B(y[1829]), .Z(n6690) );
  XOR U7452 ( .A(n6450), .B(n6690), .Z(n6451) );
  XOR U7453 ( .A(n6452), .B(n6451), .Z(n6401) );
  XOR U7454 ( .A(n6402), .B(n6401), .Z(n6404) );
  XOR U7455 ( .A(n6403), .B(n6404), .Z(n6495) );
  XOR U7456 ( .A(n6496), .B(n6495), .Z(n6392) );
  NANDN U7457 ( .A(n6270), .B(n6461), .Z(n6274) );
  NANDN U7458 ( .A(n6272), .B(n6271), .Z(n6273) );
  NAND U7459 ( .A(n6274), .B(n6273), .Z(n6502) );
  AND U7460 ( .A(x[249]), .B(y[1828]), .Z(n6434) );
  AND U7461 ( .A(x[250]), .B(y[1827]), .Z(n6431) );
  XOR U7462 ( .A(n6432), .B(n6431), .Z(n6433) );
  XOR U7463 ( .A(n6434), .B(n6433), .Z(n6500) );
  AND U7464 ( .A(x[252]), .B(y[1825]), .Z(n6449) );
  XOR U7465 ( .A(o[61]), .B(n6449), .Z(n6510) );
  AND U7466 ( .A(x[224]), .B(y[1853]), .Z(n6508) );
  AND U7467 ( .A(x[253]), .B(y[1824]), .Z(n6507) );
  XOR U7468 ( .A(n6508), .B(n6507), .Z(n6509) );
  XNOR U7469 ( .A(n6510), .B(n6509), .Z(n6499) );
  XOR U7470 ( .A(n6502), .B(n6501), .Z(n6390) );
  NAND U7471 ( .A(n6276), .B(n6275), .Z(n6280) );
  NAND U7472 ( .A(n6278), .B(n6277), .Z(n6279) );
  NAND U7473 ( .A(n6280), .B(n6279), .Z(n6470) );
  ANDN U7474 ( .B(o[60]), .A(n6281), .Z(n6410) );
  AND U7475 ( .A(x[240]), .B(y[1837]), .Z(n6408) );
  AND U7476 ( .A(x[251]), .B(y[1826]), .Z(n6407) );
  XOR U7477 ( .A(n6408), .B(n6407), .Z(n6409) );
  XOR U7478 ( .A(n6410), .B(n6409), .Z(n6469) );
  AND U7479 ( .A(x[226]), .B(y[1851]), .Z(n6420) );
  XOR U7480 ( .A(n6420), .B(n6419), .Z(n6421) );
  XOR U7481 ( .A(n6422), .B(n6421), .Z(n6468) );
  XOR U7482 ( .A(n6469), .B(n6468), .Z(n6471) );
  XNOR U7483 ( .A(n6470), .B(n6471), .Z(n6389) );
  XOR U7484 ( .A(n6390), .B(n6389), .Z(n6391) );
  NANDN U7485 ( .A(n6283), .B(n6282), .Z(n6287) );
  NANDN U7486 ( .A(n6285), .B(n6284), .Z(n6286) );
  AND U7487 ( .A(n6287), .B(n6286), .Z(n6396) );
  NAND U7488 ( .A(n6289), .B(n6288), .Z(n6293) );
  NAND U7489 ( .A(n6291), .B(n6290), .Z(n6292) );
  NAND U7490 ( .A(n6293), .B(n6292), .Z(n6426) );
  NAND U7491 ( .A(n6295), .B(n6294), .Z(n6299) );
  NAND U7492 ( .A(n6297), .B(n6296), .Z(n6298) );
  NAND U7493 ( .A(n6299), .B(n6298), .Z(n6425) );
  XOR U7494 ( .A(n6426), .B(n6425), .Z(n6428) );
  AND U7495 ( .A(x[232]), .B(y[1845]), .Z(n6463) );
  AND U7496 ( .A(y[1847]), .B(x[230]), .Z(n6301) );
  NAND U7497 ( .A(y[1846]), .B(x[231]), .Z(n6300) );
  XNOR U7498 ( .A(n6301), .B(n6300), .Z(n6462) );
  XNOR U7499 ( .A(n6463), .B(n6462), .Z(n6505) );
  NAND U7500 ( .A(x[233]), .B(y[1844]), .Z(n6608) );
  AND U7501 ( .A(x[229]), .B(y[1848]), .Z(n6416) );
  AND U7502 ( .A(x[228]), .B(y[1849]), .Z(n6414) );
  AND U7503 ( .A(x[234]), .B(y[1843]), .Z(n6413) );
  XOR U7504 ( .A(n6414), .B(n6413), .Z(n6415) );
  XNOR U7505 ( .A(n6416), .B(n6415), .Z(n6506) );
  XOR U7506 ( .A(n6608), .B(n6506), .Z(n6302) );
  XNOR U7507 ( .A(n6505), .B(n6302), .Z(n6427) );
  XNOR U7508 ( .A(n6428), .B(n6427), .Z(n6395) );
  XOR U7509 ( .A(n6398), .B(n6397), .Z(n6476) );
  NAND U7510 ( .A(n6304), .B(n6303), .Z(n6308) );
  NANDN U7511 ( .A(n6306), .B(n6305), .Z(n6307) );
  NAND U7512 ( .A(n6308), .B(n6307), .Z(n6475) );
  XNOR U7513 ( .A(n6372), .B(n6371), .Z(n6373) );
  NANDN U7514 ( .A(n6310), .B(n6309), .Z(n6314) );
  OR U7515 ( .A(n6312), .B(n6311), .Z(n6313) );
  AND U7516 ( .A(n6314), .B(n6313), .Z(n6366) );
  NAND U7517 ( .A(n6316), .B(n6315), .Z(n6320) );
  NAND U7518 ( .A(n6318), .B(n6317), .Z(n6319) );
  AND U7519 ( .A(n6320), .B(n6319), .Z(n6365) );
  XNOR U7520 ( .A(n6366), .B(n6365), .Z(n6367) );
  NANDN U7521 ( .A(n6322), .B(n6321), .Z(n6326) );
  NANDN U7522 ( .A(n6324), .B(n6323), .Z(n6325) );
  NAND U7523 ( .A(n6326), .B(n6325), .Z(n6379) );
  NAND U7524 ( .A(n6328), .B(n6327), .Z(n6332) );
  NANDN U7525 ( .A(n6330), .B(n6329), .Z(n6331) );
  NAND U7526 ( .A(n6332), .B(n6331), .Z(n6377) );
  NANDN U7527 ( .A(n6334), .B(n6333), .Z(n6338) );
  NAND U7528 ( .A(n6336), .B(n6335), .Z(n6337) );
  AND U7529 ( .A(n6338), .B(n6337), .Z(n6386) );
  NAND U7530 ( .A(n6340), .B(n6339), .Z(n6344) );
  NANDN U7531 ( .A(n6342), .B(n6341), .Z(n6343) );
  AND U7532 ( .A(n6344), .B(n6343), .Z(n6384) );
  NAND U7533 ( .A(n6346), .B(n6345), .Z(n6350) );
  NANDN U7534 ( .A(n6348), .B(n6347), .Z(n6349) );
  NAND U7535 ( .A(n6350), .B(n6349), .Z(n6383) );
  XOR U7536 ( .A(n6377), .B(n6378), .Z(n6380) );
  XNOR U7537 ( .A(n6379), .B(n6380), .Z(n6368) );
  XOR U7538 ( .A(n6367), .B(n6368), .Z(n6374) );
  XNOR U7539 ( .A(n6373), .B(n6374), .Z(n6363) );
  XOR U7540 ( .A(n6364), .B(n6363), .Z(n6356) );
  XOR U7541 ( .A(n6355), .B(n6356), .Z(n6358) );
  XOR U7542 ( .A(n6357), .B(n6358), .Z(n6354) );
  XNOR U7543 ( .A(n6353), .B(n6354), .Z(n6351) );
  XOR U7544 ( .A(n6352), .B(n6351), .Z(N126) );
  NAND U7545 ( .A(n6356), .B(n6355), .Z(n6360) );
  NAND U7546 ( .A(n6358), .B(n6357), .Z(n6359) );
  AND U7547 ( .A(n6360), .B(n6359), .Z(n6809) );
  XNOR U7548 ( .A(n6810), .B(n6809), .Z(n6808) );
  NANDN U7549 ( .A(n6366), .B(n6365), .Z(n6370) );
  NANDN U7550 ( .A(n6368), .B(n6367), .Z(n6369) );
  AND U7551 ( .A(n6370), .B(n6369), .Z(n6798) );
  NANDN U7552 ( .A(n6372), .B(n6371), .Z(n6376) );
  NANDN U7553 ( .A(n6374), .B(n6373), .Z(n6375) );
  AND U7554 ( .A(n6376), .B(n6375), .Z(n6797) );
  XOR U7555 ( .A(n6798), .B(n6797), .Z(n6796) );
  NAND U7556 ( .A(n6378), .B(n6377), .Z(n6382) );
  NAND U7557 ( .A(n6380), .B(n6379), .Z(n6381) );
  AND U7558 ( .A(n6382), .B(n6381), .Z(n6795) );
  XOR U7559 ( .A(n6796), .B(n6795), .Z(n6526) );
  NANDN U7560 ( .A(n6384), .B(n6383), .Z(n6388) );
  NANDN U7561 ( .A(n6386), .B(n6385), .Z(n6387) );
  AND U7562 ( .A(n6388), .B(n6387), .Z(n6792) );
  NAND U7563 ( .A(n6390), .B(n6389), .Z(n6394) );
  NANDN U7564 ( .A(n6392), .B(n6391), .Z(n6393) );
  NAND U7565 ( .A(n6394), .B(n6393), .Z(n6791) );
  XOR U7566 ( .A(n6792), .B(n6791), .Z(n6789) );
  NANDN U7567 ( .A(n6396), .B(n6395), .Z(n6400) );
  NAND U7568 ( .A(n6398), .B(n6397), .Z(n6399) );
  AND U7569 ( .A(n6400), .B(n6399), .Z(n6529) );
  NAND U7570 ( .A(n6402), .B(n6401), .Z(n6406) );
  NAND U7571 ( .A(n6404), .B(n6403), .Z(n6405) );
  AND U7572 ( .A(n6406), .B(n6405), .Z(n6779) );
  NAND U7573 ( .A(n6408), .B(n6407), .Z(n6412) );
  NAND U7574 ( .A(n6410), .B(n6409), .Z(n6411) );
  NAND U7575 ( .A(n6412), .B(n6411), .Z(n6667) );
  NAND U7576 ( .A(n6414), .B(n6413), .Z(n6418) );
  NAND U7577 ( .A(n6416), .B(n6415), .Z(n6417) );
  NAND U7578 ( .A(n6418), .B(n6417), .Z(n6670) );
  AND U7579 ( .A(x[230]), .B(y[1848]), .Z(n6554) );
  AND U7580 ( .A(x[229]), .B(y[1849]), .Z(n6556) );
  AND U7581 ( .A(x[243]), .B(y[1835]), .Z(n6555) );
  XOR U7582 ( .A(n6556), .B(n6555), .Z(n6553) );
  XNOR U7583 ( .A(n6554), .B(n6553), .Z(n6633) );
  AND U7584 ( .A(x[228]), .B(y[1850]), .Z(n6738) );
  AND U7585 ( .A(x[227]), .B(y[1851]), .Z(n6740) );
  AND U7586 ( .A(x[242]), .B(y[1836]), .Z(n6739) );
  XOR U7587 ( .A(n6740), .B(n6739), .Z(n6737) );
  XOR U7588 ( .A(n6738), .B(n6737), .Z(n6636) );
  NAND U7589 ( .A(n6420), .B(n6419), .Z(n6424) );
  NAND U7590 ( .A(n6422), .B(n6421), .Z(n6423) );
  AND U7591 ( .A(n6424), .B(n6423), .Z(n6635) );
  XOR U7592 ( .A(n6633), .B(n6634), .Z(n6669) );
  XOR U7593 ( .A(n6670), .B(n6669), .Z(n6668) );
  XOR U7594 ( .A(n6667), .B(n6668), .Z(n6780) );
  NAND U7595 ( .A(n6426), .B(n6425), .Z(n6430) );
  NAND U7596 ( .A(n6428), .B(n6427), .Z(n6429) );
  AND U7597 ( .A(n6430), .B(n6429), .Z(n6777) );
  XOR U7598 ( .A(n6778), .B(n6777), .Z(n6532) );
  IV U7599 ( .A(n6532), .Z(n6474) );
  AND U7600 ( .A(n6432), .B(n6431), .Z(n6436) );
  NAND U7601 ( .A(n6434), .B(n6433), .Z(n6435) );
  NANDN U7602 ( .A(n6436), .B(n6435), .Z(n6661) );
  AND U7603 ( .A(n6559), .B(n6437), .Z(n6441) );
  NAND U7604 ( .A(n6439), .B(n6438), .Z(n6440) );
  NANDN U7605 ( .A(n6441), .B(n6440), .Z(n6664) );
  NANDN U7606 ( .A(n6684), .B(n6442), .Z(n6446) );
  NANDN U7607 ( .A(n6444), .B(n6443), .Z(n6445) );
  AND U7608 ( .A(n6446), .B(n6445), .Z(n6642) );
  AND U7609 ( .A(x[247]), .B(y[1831]), .Z(n6688) );
  AND U7610 ( .A(y[1830]), .B(x[248]), .Z(n6448) );
  AND U7611 ( .A(y[1829]), .B(x[249]), .Z(n6447) );
  XOR U7612 ( .A(n6448), .B(n6447), .Z(n6687) );
  XOR U7613 ( .A(n6688), .B(n6687), .Z(n6644) );
  AND U7614 ( .A(n6449), .B(o[61]), .Z(n6732) );
  AND U7615 ( .A(x[252]), .B(y[1826]), .Z(n6734) );
  AND U7616 ( .A(x[240]), .B(y[1838]), .Z(n6733) );
  XOR U7617 ( .A(n6734), .B(n6733), .Z(n6731) );
  XNOR U7618 ( .A(n6732), .B(n6731), .Z(n6643) );
  XNOR U7619 ( .A(n6642), .B(n6641), .Z(n6663) );
  XOR U7620 ( .A(n6664), .B(n6663), .Z(n6662) );
  XOR U7621 ( .A(n6661), .B(n6662), .Z(n6772) );
  NAND U7622 ( .A(n6450), .B(n6690), .Z(n6454) );
  NAND U7623 ( .A(n6452), .B(n6451), .Z(n6453) );
  NAND U7624 ( .A(n6454), .B(n6453), .Z(n6762) );
  NAND U7625 ( .A(n6456), .B(n6455), .Z(n6460) );
  NAND U7626 ( .A(n6458), .B(n6457), .Z(n6459) );
  AND U7627 ( .A(n6460), .B(n6459), .Z(n6550) );
  AND U7628 ( .A(x[224]), .B(y[1854]), .Z(n6612) );
  AND U7629 ( .A(x[253]), .B(y[1825]), .Z(n6591) );
  XOR U7630 ( .A(o[62]), .B(n6591), .Z(n6614) );
  AND U7631 ( .A(x[254]), .B(y[1824]), .Z(n6613) );
  XOR U7632 ( .A(n6614), .B(n6613), .Z(n6611) );
  XOR U7633 ( .A(n6612), .B(n6611), .Z(n6547) );
  AND U7634 ( .A(x[244]), .B(y[1834]), .Z(n6725) );
  XOR U7635 ( .A(n6726), .B(n6725), .Z(n6724) );
  AND U7636 ( .A(x[232]), .B(y[1846]), .Z(n6723) );
  XNOR U7637 ( .A(n6724), .B(n6723), .Z(n6548) );
  XNOR U7638 ( .A(n6550), .B(n6549), .Z(n6761) );
  XOR U7639 ( .A(n6762), .B(n6761), .Z(n6759) );
  AND U7640 ( .A(x[231]), .B(y[1847]), .Z(n6682) );
  NAND U7641 ( .A(n6461), .B(n6682), .Z(n6465) );
  NAND U7642 ( .A(n6463), .B(n6462), .Z(n6464) );
  AND U7643 ( .A(n6465), .B(n6464), .Z(n6653) );
  AND U7644 ( .A(y[1833]), .B(x[245]), .Z(n6467) );
  AND U7645 ( .A(y[1832]), .B(x[246]), .Z(n6466) );
  XOR U7646 ( .A(n6467), .B(n6466), .Z(n6681) );
  XOR U7647 ( .A(n6682), .B(n6681), .Z(n6656) );
  AND U7648 ( .A(x[241]), .B(y[1837]), .Z(n6718) );
  AND U7649 ( .A(x[226]), .B(y[1852]), .Z(n6720) );
  AND U7650 ( .A(x[250]), .B(y[1828]), .Z(n6719) );
  XOR U7651 ( .A(n6720), .B(n6719), .Z(n6717) );
  XNOR U7652 ( .A(n6718), .B(n6717), .Z(n6655) );
  XNOR U7653 ( .A(n6653), .B(n6654), .Z(n6760) );
  NAND U7654 ( .A(n6469), .B(n6468), .Z(n6473) );
  NAND U7655 ( .A(n6471), .B(n6470), .Z(n6472) );
  NAND U7656 ( .A(n6473), .B(n6472), .Z(n6773) );
  XOR U7657 ( .A(n6774), .B(n6773), .Z(n6771) );
  XOR U7658 ( .A(n6772), .B(n6771), .Z(n6531) );
  XNOR U7659 ( .A(n6474), .B(n6531), .Z(n6530) );
  XNOR U7660 ( .A(n6529), .B(n6530), .Z(n6790) );
  NANDN U7661 ( .A(n6476), .B(n6475), .Z(n6480) );
  NANDN U7662 ( .A(n6478), .B(n6477), .Z(n6479) );
  NAND U7663 ( .A(n6480), .B(n6479), .Z(n6815) );
  NANDN U7664 ( .A(n6482), .B(n6481), .Z(n6486) );
  NAND U7665 ( .A(n6484), .B(n6483), .Z(n6485) );
  AND U7666 ( .A(n6486), .B(n6485), .Z(n6535) );
  NAND U7667 ( .A(n6488), .B(n6487), .Z(n6492) );
  NAND U7668 ( .A(n6490), .B(n6489), .Z(n6491) );
  AND U7669 ( .A(n6492), .B(n6491), .Z(n6544) );
  NAND U7670 ( .A(n6494), .B(n6493), .Z(n6498) );
  NAND U7671 ( .A(n6496), .B(n6495), .Z(n6497) );
  AND U7672 ( .A(n6498), .B(n6497), .Z(n6543) );
  XOR U7673 ( .A(n6544), .B(n6543), .Z(n6542) );
  NANDN U7674 ( .A(n6500), .B(n6499), .Z(n6504) );
  OR U7675 ( .A(n6502), .B(n6501), .Z(n6503) );
  NAND U7676 ( .A(n6504), .B(n6503), .Z(n6541) );
  XOR U7677 ( .A(n6542), .B(n6541), .Z(n6538) );
  NAND U7678 ( .A(n6508), .B(n6507), .Z(n6512) );
  NAND U7679 ( .A(n6510), .B(n6509), .Z(n6511) );
  NAND U7680 ( .A(n6512), .B(n6511), .Z(n6647) );
  AND U7681 ( .A(y[1842]), .B(x[236]), .Z(n6513) );
  XOR U7682 ( .A(n6514), .B(n6513), .Z(n6560) );
  XOR U7683 ( .A(n6561), .B(n6560), .Z(n6606) );
  AND U7684 ( .A(y[1845]), .B(x[233]), .Z(n6516) );
  XOR U7685 ( .A(n6516), .B(n6515), .Z(n6605) );
  XOR U7686 ( .A(n6606), .B(n6605), .Z(n6650) );
  AND U7687 ( .A(x[251]), .B(y[1827]), .Z(n6700) );
  AND U7688 ( .A(x[225]), .B(y[1853]), .Z(n6699) );
  XOR U7689 ( .A(n6700), .B(n6699), .Z(n6697) );
  XOR U7690 ( .A(n6698), .B(n6697), .Z(n6649) );
  XOR U7691 ( .A(n6650), .B(n6649), .Z(n6648) );
  XOR U7692 ( .A(n6647), .B(n6648), .Z(n6756) );
  NAND U7693 ( .A(n6518), .B(n6517), .Z(n6522) );
  NANDN U7694 ( .A(n6520), .B(n6519), .Z(n6521) );
  AND U7695 ( .A(n6522), .B(n6521), .Z(n6753) );
  XNOR U7696 ( .A(n6754), .B(n6753), .Z(n6537) );
  XNOR U7697 ( .A(n6535), .B(n6536), .Z(n6816) );
  XOR U7698 ( .A(n6815), .B(n6816), .Z(n6813) );
  XOR U7699 ( .A(n6524), .B(n6523), .Z(n6807) );
  XNOR U7700 ( .A(n6808), .B(n6807), .Z(N127) );
  NANDN U7701 ( .A(n6524), .B(n6523), .Z(n6528) );
  NANDN U7702 ( .A(n6526), .B(n6525), .Z(n6527) );
  AND U7703 ( .A(n6528), .B(n6527), .Z(n6824) );
  NANDN U7704 ( .A(n6530), .B(n6529), .Z(n6534) );
  NANDN U7705 ( .A(n6532), .B(n6531), .Z(n6533) );
  AND U7706 ( .A(n6534), .B(n6533), .Z(n6806) );
  NANDN U7707 ( .A(n6536), .B(n6535), .Z(n6540) );
  NANDN U7708 ( .A(n6538), .B(n6537), .Z(n6539) );
  AND U7709 ( .A(n6540), .B(n6539), .Z(n6788) );
  NAND U7710 ( .A(n6542), .B(n6541), .Z(n6546) );
  NAND U7711 ( .A(n6544), .B(n6543), .Z(n6545) );
  AND U7712 ( .A(n6546), .B(n6545), .Z(n6770) );
  ANDN U7713 ( .B(n6548), .A(n6547), .Z(n6552) );
  AND U7714 ( .A(n6550), .B(n6549), .Z(n6551) );
  NOR U7715 ( .A(n6552), .B(n6551), .Z(n6632) );
  NAND U7716 ( .A(n6554), .B(n6553), .Z(n6558) );
  NAND U7717 ( .A(n6556), .B(n6555), .Z(n6557) );
  AND U7718 ( .A(n6558), .B(n6557), .Z(n6565) );
  NAND U7719 ( .A(n6559), .B(n6572), .Z(n6563) );
  NAND U7720 ( .A(n6561), .B(n6560), .Z(n6562) );
  AND U7721 ( .A(n6563), .B(n6562), .Z(n6564) );
  XNOR U7722 ( .A(n6565), .B(n6564), .Z(n6630) );
  AND U7723 ( .A(y[1828]), .B(x[251]), .Z(n6567) );
  NAND U7724 ( .A(y[1838]), .B(x[241]), .Z(n6566) );
  XNOR U7725 ( .A(n6567), .B(n6566), .Z(n6571) );
  AND U7726 ( .A(y[1824]), .B(x[255]), .Z(n6569) );
  NAND U7727 ( .A(y[1852]), .B(x[227]), .Z(n6568) );
  XNOR U7728 ( .A(n6569), .B(n6568), .Z(n6570) );
  XOR U7729 ( .A(n6571), .B(n6570), .Z(n6574) );
  AND U7730 ( .A(x[234]), .B(y[1845]), .Z(n6607) );
  XNOR U7731 ( .A(n6572), .B(n6607), .Z(n6573) );
  XNOR U7732 ( .A(n6574), .B(n6573), .Z(n6590) );
  AND U7733 ( .A(y[1836]), .B(x[243]), .Z(n6576) );
  NAND U7734 ( .A(y[1851]), .B(x[228]), .Z(n6575) );
  XNOR U7735 ( .A(n6576), .B(n6575), .Z(n6580) );
  AND U7736 ( .A(y[1834]), .B(x[245]), .Z(n6578) );
  NAND U7737 ( .A(y[1847]), .B(x[232]), .Z(n6577) );
  XNOR U7738 ( .A(n6578), .B(n6577), .Z(n6579) );
  XOR U7739 ( .A(n6580), .B(n6579), .Z(n6588) );
  AND U7740 ( .A(y[1850]), .B(x[229]), .Z(n6582) );
  NAND U7741 ( .A(y[1837]), .B(x[242]), .Z(n6581) );
  XNOR U7742 ( .A(n6582), .B(n6581), .Z(n6586) );
  AND U7743 ( .A(y[1849]), .B(x[230]), .Z(n6584) );
  NAND U7744 ( .A(y[1848]), .B(x[231]), .Z(n6583) );
  XNOR U7745 ( .A(n6584), .B(n6583), .Z(n6585) );
  XNOR U7746 ( .A(n6586), .B(n6585), .Z(n6587) );
  XNOR U7747 ( .A(n6588), .B(n6587), .Z(n6589) );
  XOR U7748 ( .A(n6590), .B(n6589), .Z(n6604) );
  AND U7749 ( .A(y[1841]), .B(x[238]), .Z(n6598) );
  AND U7750 ( .A(n6591), .B(o[62]), .Z(n6596) );
  AND U7751 ( .A(x[246]), .B(y[1833]), .Z(n6683) );
  XOR U7752 ( .A(n6683), .B(o[63]), .Z(n6594) );
  AND U7753 ( .A(x[249]), .B(y[1830]), .Z(n6689) );
  XNOR U7754 ( .A(n6592), .B(n6689), .Z(n6593) );
  XNOR U7755 ( .A(n6594), .B(n6593), .Z(n6595) );
  XNOR U7756 ( .A(n6596), .B(n6595), .Z(n6597) );
  XNOR U7757 ( .A(n6598), .B(n6597), .Z(n6602) );
  AND U7758 ( .A(y[1832]), .B(x[247]), .Z(n6600) );
  NAND U7759 ( .A(y[1853]), .B(x[226]), .Z(n6599) );
  XNOR U7760 ( .A(n6600), .B(n6599), .Z(n6601) );
  XNOR U7761 ( .A(n6602), .B(n6601), .Z(n6603) );
  XNOR U7762 ( .A(n6604), .B(n6603), .Z(n6620) );
  NAND U7763 ( .A(n6606), .B(n6605), .Z(n6610) );
  NANDN U7764 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U7765 ( .A(n6610), .B(n6609), .Z(n6618) );
  NAND U7766 ( .A(n6612), .B(n6611), .Z(n6616) );
  NAND U7767 ( .A(n6614), .B(n6613), .Z(n6615) );
  NAND U7768 ( .A(n6616), .B(n6615), .Z(n6617) );
  XNOR U7769 ( .A(n6618), .B(n6617), .Z(n6619) );
  XOR U7770 ( .A(n6620), .B(n6619), .Z(n6628) );
  AND U7771 ( .A(y[1854]), .B(x[225]), .Z(n6622) );
  NAND U7772 ( .A(y[1846]), .B(x[233]), .Z(n6621) );
  XNOR U7773 ( .A(n6622), .B(n6621), .Z(n6626) );
  AND U7774 ( .A(y[1827]), .B(x[252]), .Z(n6624) );
  NAND U7775 ( .A(y[1855]), .B(x[224]), .Z(n6623) );
  XNOR U7776 ( .A(n6624), .B(n6623), .Z(n6625) );
  XNOR U7777 ( .A(n6626), .B(n6625), .Z(n6627) );
  XNOR U7778 ( .A(n6628), .B(n6627), .Z(n6629) );
  XOR U7779 ( .A(n6630), .B(n6629), .Z(n6631) );
  XNOR U7780 ( .A(n6632), .B(n6631), .Z(n6640) );
  NANDN U7781 ( .A(n6634), .B(n6633), .Z(n6638) );
  NANDN U7782 ( .A(n6636), .B(n6635), .Z(n6637) );
  NAND U7783 ( .A(n6638), .B(n6637), .Z(n6639) );
  XNOR U7784 ( .A(n6640), .B(n6639), .Z(n6680) );
  NAND U7785 ( .A(n6642), .B(n6641), .Z(n6646) );
  NANDN U7786 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U7787 ( .A(n6646), .B(n6645), .Z(n6678) );
  NAND U7788 ( .A(n6648), .B(n6647), .Z(n6652) );
  NAND U7789 ( .A(n6650), .B(n6649), .Z(n6651) );
  AND U7790 ( .A(n6652), .B(n6651), .Z(n6660) );
  NANDN U7791 ( .A(n6654), .B(n6653), .Z(n6658) );
  NANDN U7792 ( .A(n6656), .B(n6655), .Z(n6657) );
  NAND U7793 ( .A(n6658), .B(n6657), .Z(n6659) );
  XNOR U7794 ( .A(n6660), .B(n6659), .Z(n6676) );
  NAND U7795 ( .A(n6662), .B(n6661), .Z(n6666) );
  NAND U7796 ( .A(n6664), .B(n6663), .Z(n6665) );
  AND U7797 ( .A(n6666), .B(n6665), .Z(n6674) );
  NAND U7798 ( .A(n6668), .B(n6667), .Z(n6672) );
  NAND U7799 ( .A(n6670), .B(n6669), .Z(n6671) );
  NAND U7800 ( .A(n6672), .B(n6671), .Z(n6673) );
  XNOR U7801 ( .A(n6674), .B(n6673), .Z(n6675) );
  XNOR U7802 ( .A(n6676), .B(n6675), .Z(n6677) );
  XNOR U7803 ( .A(n6678), .B(n6677), .Z(n6679) );
  XOR U7804 ( .A(n6680), .B(n6679), .Z(n6752) );
  NAND U7805 ( .A(n6682), .B(n6681), .Z(n6686) );
  NANDN U7806 ( .A(n6684), .B(n6683), .Z(n6685) );
  AND U7807 ( .A(n6686), .B(n6685), .Z(n6694) );
  NAND U7808 ( .A(n6688), .B(n6687), .Z(n6692) );
  NAND U7809 ( .A(n6690), .B(n6689), .Z(n6691) );
  NAND U7810 ( .A(n6692), .B(n6691), .Z(n6693) );
  XNOR U7811 ( .A(n6694), .B(n6693), .Z(n6750) );
  AND U7812 ( .A(y[1825]), .B(x[254]), .Z(n6696) );
  NAND U7813 ( .A(y[1839]), .B(x[240]), .Z(n6695) );
  XNOR U7814 ( .A(n6696), .B(n6695), .Z(n6716) );
  AND U7815 ( .A(y[1835]), .B(x[244]), .Z(n6714) );
  NAND U7816 ( .A(n6698), .B(n6697), .Z(n6702) );
  NAND U7817 ( .A(n6700), .B(n6699), .Z(n6701) );
  AND U7818 ( .A(n6702), .B(n6701), .Z(n6710) );
  AND U7819 ( .A(y[1826]), .B(x[253]), .Z(n6704) );
  NAND U7820 ( .A(y[1829]), .B(x[250]), .Z(n6703) );
  XNOR U7821 ( .A(n6704), .B(n6703), .Z(n6708) );
  AND U7822 ( .A(y[1844]), .B(x[235]), .Z(n6706) );
  NAND U7823 ( .A(y[1843]), .B(x[236]), .Z(n6705) );
  XNOR U7824 ( .A(n6706), .B(n6705), .Z(n6707) );
  XNOR U7825 ( .A(n6708), .B(n6707), .Z(n6709) );
  XNOR U7826 ( .A(n6710), .B(n6709), .Z(n6711) );
  XNOR U7827 ( .A(n6712), .B(n6711), .Z(n6713) );
  XNOR U7828 ( .A(n6714), .B(n6713), .Z(n6715) );
  XOR U7829 ( .A(n6716), .B(n6715), .Z(n6748) );
  NAND U7830 ( .A(n6718), .B(n6717), .Z(n6722) );
  NAND U7831 ( .A(n6720), .B(n6719), .Z(n6721) );
  AND U7832 ( .A(n6722), .B(n6721), .Z(n6730) );
  NAND U7833 ( .A(n6724), .B(n6723), .Z(n6728) );
  NAND U7834 ( .A(n6726), .B(n6725), .Z(n6727) );
  NAND U7835 ( .A(n6728), .B(n6727), .Z(n6729) );
  XNOR U7836 ( .A(n6730), .B(n6729), .Z(n6746) );
  NAND U7837 ( .A(n6732), .B(n6731), .Z(n6736) );
  NAND U7838 ( .A(n6734), .B(n6733), .Z(n6735) );
  AND U7839 ( .A(n6736), .B(n6735), .Z(n6744) );
  NAND U7840 ( .A(n6738), .B(n6737), .Z(n6742) );
  NAND U7841 ( .A(n6740), .B(n6739), .Z(n6741) );
  NAND U7842 ( .A(n6742), .B(n6741), .Z(n6743) );
  XNOR U7843 ( .A(n6744), .B(n6743), .Z(n6745) );
  XNOR U7844 ( .A(n6746), .B(n6745), .Z(n6747) );
  XNOR U7845 ( .A(n6748), .B(n6747), .Z(n6749) );
  XNOR U7846 ( .A(n6750), .B(n6749), .Z(n6751) );
  XNOR U7847 ( .A(n6752), .B(n6751), .Z(n6768) );
  NAND U7848 ( .A(n6754), .B(n6753), .Z(n6758) );
  NANDN U7849 ( .A(n6756), .B(n6755), .Z(n6757) );
  AND U7850 ( .A(n6758), .B(n6757), .Z(n6766) );
  NANDN U7851 ( .A(n6760), .B(n6759), .Z(n6764) );
  NAND U7852 ( .A(n6762), .B(n6761), .Z(n6763) );
  NAND U7853 ( .A(n6764), .B(n6763), .Z(n6765) );
  XNOR U7854 ( .A(n6766), .B(n6765), .Z(n6767) );
  XNOR U7855 ( .A(n6768), .B(n6767), .Z(n6769) );
  XNOR U7856 ( .A(n6770), .B(n6769), .Z(n6786) );
  NAND U7857 ( .A(n6772), .B(n6771), .Z(n6776) );
  NAND U7858 ( .A(n6774), .B(n6773), .Z(n6775) );
  AND U7859 ( .A(n6776), .B(n6775), .Z(n6784) );
  NAND U7860 ( .A(n6778), .B(n6777), .Z(n6782) );
  NANDN U7861 ( .A(n6780), .B(n6779), .Z(n6781) );
  NAND U7862 ( .A(n6782), .B(n6781), .Z(n6783) );
  XNOR U7863 ( .A(n6784), .B(n6783), .Z(n6785) );
  XNOR U7864 ( .A(n6786), .B(n6785), .Z(n6787) );
  XNOR U7865 ( .A(n6788), .B(n6787), .Z(n6804) );
  NANDN U7866 ( .A(n6790), .B(n6789), .Z(n6794) );
  NAND U7867 ( .A(n6792), .B(n6791), .Z(n6793) );
  AND U7868 ( .A(n6794), .B(n6793), .Z(n6802) );
  NAND U7869 ( .A(n6796), .B(n6795), .Z(n6800) );
  NAND U7870 ( .A(n6798), .B(n6797), .Z(n6799) );
  NAND U7871 ( .A(n6800), .B(n6799), .Z(n6801) );
  XNOR U7872 ( .A(n6802), .B(n6801), .Z(n6803) );
  XNOR U7873 ( .A(n6804), .B(n6803), .Z(n6805) );
  XNOR U7874 ( .A(n6806), .B(n6805), .Z(n6822) );
  NAND U7875 ( .A(n6808), .B(n6807), .Z(n6812) );
  NANDN U7876 ( .A(n6810), .B(n6809), .Z(n6811) );
  AND U7877 ( .A(n6812), .B(n6811), .Z(n6820) );
  NANDN U7878 ( .A(n6814), .B(n6813), .Z(n6818) );
  NAND U7879 ( .A(n6816), .B(n6815), .Z(n6817) );
  NAND U7880 ( .A(n6818), .B(n6817), .Z(n6819) );
  XNOR U7881 ( .A(n6820), .B(n6819), .Z(n6821) );
  XNOR U7882 ( .A(n6822), .B(n6821), .Z(n6823) );
  XNOR U7883 ( .A(n6824), .B(n6823), .Z(N128) );
  AND U7884 ( .A(x[224]), .B(y[1856]), .Z(n7479) );
  XOR U7885 ( .A(n7479), .B(o[64]), .Z(N161) );
  AND U7886 ( .A(x[225]), .B(y[1856]), .Z(n6833) );
  AND U7887 ( .A(x[224]), .B(y[1857]), .Z(n6832) );
  XNOR U7888 ( .A(n6832), .B(o[65]), .Z(n6825) );
  XNOR U7889 ( .A(n6833), .B(n6825), .Z(n6827) );
  NAND U7890 ( .A(n7479), .B(o[64]), .Z(n6826) );
  XNOR U7891 ( .A(n6827), .B(n6826), .Z(N162) );
  NANDN U7892 ( .A(n6833), .B(n6825), .Z(n6829) );
  NAND U7893 ( .A(n6827), .B(n6826), .Z(n6828) );
  AND U7894 ( .A(n6829), .B(n6828), .Z(n6839) );
  AND U7895 ( .A(x[224]), .B(y[1858]), .Z(n6846) );
  XNOR U7896 ( .A(n6846), .B(o[66]), .Z(n6838) );
  XNOR U7897 ( .A(n6839), .B(n6838), .Z(n6841) );
  AND U7898 ( .A(y[1856]), .B(x[226]), .Z(n6831) );
  NAND U7899 ( .A(y[1857]), .B(x[225]), .Z(n6830) );
  XNOR U7900 ( .A(n6831), .B(n6830), .Z(n6835) );
  AND U7901 ( .A(n6832), .B(o[65]), .Z(n6834) );
  XNOR U7902 ( .A(n6835), .B(n6834), .Z(n6840) );
  XNOR U7903 ( .A(n6841), .B(n6840), .Z(N163) );
  NAND U7904 ( .A(x[226]), .B(y[1857]), .Z(n6853) );
  NANDN U7905 ( .A(n6853), .B(n6833), .Z(n6837) );
  NAND U7906 ( .A(n6835), .B(n6834), .Z(n6836) );
  AND U7907 ( .A(n6837), .B(n6836), .Z(n6859) );
  NANDN U7908 ( .A(n6839), .B(n6838), .Z(n6843) );
  NAND U7909 ( .A(n6841), .B(n6840), .Z(n6842) );
  AND U7910 ( .A(n6843), .B(n6842), .Z(n6858) );
  XNOR U7911 ( .A(n6859), .B(n6858), .Z(n6861) );
  AND U7912 ( .A(x[225]), .B(y[1858]), .Z(n6966) );
  XOR U7913 ( .A(n6966), .B(n6855), .Z(n6857) );
  AND U7914 ( .A(y[1856]), .B(x[227]), .Z(n6845) );
  NAND U7915 ( .A(y[1859]), .B(x[224]), .Z(n6844) );
  XNOR U7916 ( .A(n6845), .B(n6844), .Z(n6848) );
  AND U7917 ( .A(n6846), .B(o[66]), .Z(n6847) );
  XOR U7918 ( .A(n6848), .B(n6847), .Z(n6856) );
  XOR U7919 ( .A(n6857), .B(n6856), .Z(n6860) );
  XOR U7920 ( .A(n6861), .B(n6860), .Z(N164) );
  AND U7921 ( .A(x[227]), .B(y[1859]), .Z(n6901) );
  NAND U7922 ( .A(n7479), .B(n6901), .Z(n6850) );
  NAND U7923 ( .A(n6848), .B(n6847), .Z(n6849) );
  NAND U7924 ( .A(n6850), .B(n6849), .Z(n6879) );
  AND U7925 ( .A(y[1860]), .B(x[224]), .Z(n6852) );
  NAND U7926 ( .A(y[1856]), .B(x[228]), .Z(n6851) );
  XNOR U7927 ( .A(n6852), .B(n6851), .Z(n6873) );
  ANDN U7928 ( .B(o[67]), .A(n6853), .Z(n6874) );
  XOR U7929 ( .A(n6873), .B(n6874), .Z(n6878) );
  AND U7930 ( .A(y[1858]), .B(x[226]), .Z(n7013) );
  NAND U7931 ( .A(y[1859]), .B(x[225]), .Z(n6854) );
  XNOR U7932 ( .A(n7013), .B(n6854), .Z(n6872) );
  AND U7933 ( .A(x[227]), .B(y[1857]), .Z(n6867) );
  XOR U7934 ( .A(o[68]), .B(n6867), .Z(n6871) );
  XOR U7935 ( .A(n6872), .B(n6871), .Z(n6877) );
  XOR U7936 ( .A(n6878), .B(n6877), .Z(n6880) );
  XNOR U7937 ( .A(n6879), .B(n6880), .Z(n6885) );
  NANDN U7938 ( .A(n6859), .B(n6858), .Z(n6863) );
  NAND U7939 ( .A(n6861), .B(n6860), .Z(n6862) );
  NAND U7940 ( .A(n6863), .B(n6862), .Z(n6884) );
  XOR U7941 ( .A(n6883), .B(n6884), .Z(n6864) );
  XNOR U7942 ( .A(n6885), .B(n6864), .Z(N165) );
  AND U7943 ( .A(y[1858]), .B(x[227]), .Z(n6866) );
  NAND U7944 ( .A(y[1860]), .B(x[225]), .Z(n6865) );
  XNOR U7945 ( .A(n6866), .B(n6865), .Z(n6888) );
  AND U7946 ( .A(x[228]), .B(y[1857]), .Z(n6897) );
  XOR U7947 ( .A(n6897), .B(o[69]), .Z(n6887) );
  XNOR U7948 ( .A(n6888), .B(n6887), .Z(n6891) );
  NAND U7949 ( .A(x[226]), .B(y[1859]), .Z(n6975) );
  AND U7950 ( .A(o[68]), .B(n6867), .Z(n6893) );
  AND U7951 ( .A(y[1856]), .B(x[229]), .Z(n6869) );
  NAND U7952 ( .A(y[1861]), .B(x[224]), .Z(n6868) );
  XNOR U7953 ( .A(n6869), .B(n6868), .Z(n6894) );
  XOR U7954 ( .A(n6893), .B(n6894), .Z(n6892) );
  XOR U7955 ( .A(n6975), .B(n6892), .Z(n6870) );
  XOR U7956 ( .A(n6891), .B(n6870), .Z(n6905) );
  AND U7957 ( .A(x[228]), .B(y[1860]), .Z(n7690) );
  NAND U7958 ( .A(n7690), .B(n7479), .Z(n6876) );
  NAND U7959 ( .A(n6874), .B(n6873), .Z(n6875) );
  NAND U7960 ( .A(n6876), .B(n6875), .Z(n6903) );
  XOR U7961 ( .A(n6904), .B(n6903), .Z(n6906) );
  XNOR U7962 ( .A(n6905), .B(n6906), .Z(n6911) );
  NAND U7963 ( .A(n6878), .B(n6877), .Z(n6882) );
  NAND U7964 ( .A(n6880), .B(n6879), .Z(n6881) );
  AND U7965 ( .A(n6882), .B(n6881), .Z(n6910) );
  XNOR U7966 ( .A(n6910), .B(n6909), .Z(n6886) );
  XNOR U7967 ( .A(n6911), .B(n6886), .Z(N166) );
  AND U7968 ( .A(x[227]), .B(y[1860]), .Z(n6976) );
  NAND U7969 ( .A(n6976), .B(n6966), .Z(n6890) );
  NAND U7970 ( .A(n6888), .B(n6887), .Z(n6889) );
  NAND U7971 ( .A(n6890), .B(n6889), .Z(n6941) );
  XOR U7972 ( .A(n6941), .B(n6940), .Z(n6943) );
  AND U7973 ( .A(x[229]), .B(y[1861]), .Z(n7150) );
  NAND U7974 ( .A(n7479), .B(n7150), .Z(n6896) );
  NAND U7975 ( .A(n6894), .B(n6893), .Z(n6895) );
  NAND U7976 ( .A(n6896), .B(n6895), .Z(n6914) );
  AND U7977 ( .A(n6897), .B(o[69]), .Z(n6920) );
  AND U7978 ( .A(y[1856]), .B(x[230]), .Z(n6899) );
  NAND U7979 ( .A(y[1862]), .B(x[224]), .Z(n6898) );
  XNOR U7980 ( .A(n6899), .B(n6898), .Z(n6921) );
  XOR U7981 ( .A(n6920), .B(n6921), .Z(n6913) );
  XOR U7982 ( .A(n6914), .B(n6913), .Z(n6916) );
  NAND U7983 ( .A(y[1860]), .B(x[226]), .Z(n6900) );
  XNOR U7984 ( .A(n6901), .B(n6900), .Z(n6925) );
  AND U7985 ( .A(y[1861]), .B(x[225]), .Z(n7171) );
  NAND U7986 ( .A(y[1858]), .B(x[228]), .Z(n6902) );
  XNOR U7987 ( .A(n7171), .B(n6902), .Z(n6929) );
  NAND U7988 ( .A(x[229]), .B(y[1857]), .Z(n6936) );
  XOR U7989 ( .A(n6929), .B(n6928), .Z(n6924) );
  XOR U7990 ( .A(n6925), .B(n6924), .Z(n6915) );
  XOR U7991 ( .A(n6916), .B(n6915), .Z(n6942) );
  XNOR U7992 ( .A(n6943), .B(n6942), .Z(n6939) );
  NANDN U7993 ( .A(n6904), .B(n6903), .Z(n6908) );
  NANDN U7994 ( .A(n6906), .B(n6905), .Z(n6907) );
  NAND U7995 ( .A(n6908), .B(n6907), .Z(n6937) );
  XOR U7996 ( .A(n6937), .B(n6938), .Z(n6912) );
  XNOR U7997 ( .A(n6939), .B(n6912), .Z(N167) );
  NAND U7998 ( .A(n6914), .B(n6913), .Z(n6918) );
  NAND U7999 ( .A(n6916), .B(n6915), .Z(n6917) );
  AND U8000 ( .A(n6918), .B(n6917), .Z(n6950) );
  AND U8001 ( .A(y[1858]), .B(x[229]), .Z(n7058) );
  NAND U8002 ( .A(y[1862]), .B(x[225]), .Z(n6919) );
  XNOR U8003 ( .A(n7058), .B(n6919), .Z(n6968) );
  AND U8004 ( .A(x[230]), .B(y[1857]), .Z(n6972) );
  XOR U8005 ( .A(o[71]), .B(n6972), .Z(n6967) );
  XOR U8006 ( .A(n6968), .B(n6967), .Z(n6987) );
  AND U8007 ( .A(x[230]), .B(y[1862]), .Z(n7192) );
  NAND U8008 ( .A(n7479), .B(n7192), .Z(n6923) );
  NAND U8009 ( .A(n6921), .B(n6920), .Z(n6922) );
  AND U8010 ( .A(n6923), .B(n6922), .Z(n6986) );
  NANDN U8011 ( .A(n6975), .B(n6976), .Z(n6927) );
  NAND U8012 ( .A(n6925), .B(n6924), .Z(n6926) );
  AND U8013 ( .A(n6927), .B(n6926), .Z(n6988) );
  XOR U8014 ( .A(n6989), .B(n6988), .Z(n6948) );
  AND U8015 ( .A(x[228]), .B(y[1861]), .Z(n7484) );
  NAND U8016 ( .A(n7484), .B(n6966), .Z(n6931) );
  NAND U8017 ( .A(n6929), .B(n6928), .Z(n6930) );
  AND U8018 ( .A(n6931), .B(n6930), .Z(n6963) );
  AND U8019 ( .A(y[1861]), .B(x[226]), .Z(n6933) );
  NAND U8020 ( .A(y[1859]), .B(x[228]), .Z(n6932) );
  XNOR U8021 ( .A(n6933), .B(n6932), .Z(n6977) );
  XOR U8022 ( .A(n6977), .B(n6976), .Z(n6961) );
  AND U8023 ( .A(y[1856]), .B(x[231]), .Z(n6935) );
  NAND U8024 ( .A(y[1863]), .B(x[224]), .Z(n6934) );
  XNOR U8025 ( .A(n6935), .B(n6934), .Z(n6981) );
  ANDN U8026 ( .B(o[70]), .A(n6936), .Z(n6980) );
  XNOR U8027 ( .A(n6981), .B(n6980), .Z(n6960) );
  XOR U8028 ( .A(n6963), .B(n6962), .Z(n6947) );
  XOR U8029 ( .A(n6948), .B(n6947), .Z(n6949) );
  XNOR U8030 ( .A(n6950), .B(n6949), .Z(n6956) );
  NAND U8031 ( .A(n6941), .B(n6940), .Z(n6945) );
  NAND U8032 ( .A(n6943), .B(n6942), .Z(n6944) );
  AND U8033 ( .A(n6945), .B(n6944), .Z(n6955) );
  IV U8034 ( .A(n6955), .Z(n6953) );
  XOR U8035 ( .A(n6954), .B(n6953), .Z(n6946) );
  XNOR U8036 ( .A(n6956), .B(n6946), .Z(N168) );
  NAND U8037 ( .A(n6948), .B(n6947), .Z(n6952) );
  NAND U8038 ( .A(n6950), .B(n6949), .Z(n6951) );
  AND U8039 ( .A(n6952), .B(n6951), .Z(n7030) );
  NANDN U8040 ( .A(n6953), .B(n6954), .Z(n6959) );
  NOR U8041 ( .A(n6955), .B(n6954), .Z(n6957) );
  OR U8042 ( .A(n6957), .B(n6956), .Z(n6958) );
  AND U8043 ( .A(n6959), .B(n6958), .Z(n7029) );
  NANDN U8044 ( .A(n6961), .B(n6960), .Z(n6965) );
  NAND U8045 ( .A(n6963), .B(n6962), .Z(n6964) );
  AND U8046 ( .A(n6965), .B(n6964), .Z(n7026) );
  AND U8047 ( .A(x[229]), .B(y[1862]), .Z(n7142) );
  NAND U8048 ( .A(n7142), .B(n6966), .Z(n6970) );
  NAND U8049 ( .A(n6968), .B(n6967), .Z(n6969) );
  AND U8050 ( .A(n6970), .B(n6969), .Z(n7024) );
  AND U8051 ( .A(y[1859]), .B(x[229]), .Z(n7597) );
  NAND U8052 ( .A(y[1863]), .B(x[225]), .Z(n6971) );
  XNOR U8053 ( .A(n7597), .B(n6971), .Z(n7005) );
  AND U8054 ( .A(o[71]), .B(n6972), .Z(n7004) );
  XOR U8055 ( .A(n7005), .B(n7004), .Z(n7010) );
  NAND U8056 ( .A(x[227]), .B(y[1861]), .Z(n7815) );
  AND U8057 ( .A(y[1858]), .B(x[230]), .Z(n6974) );
  NAND U8058 ( .A(y[1862]), .B(x[226]), .Z(n6973) );
  XNOR U8059 ( .A(n6974), .B(n6973), .Z(n7014) );
  XNOR U8060 ( .A(n7690), .B(n7014), .Z(n7008) );
  XOR U8061 ( .A(n7815), .B(n7008), .Z(n7009) );
  XOR U8062 ( .A(n7010), .B(n7009), .Z(n7023) );
  XOR U8063 ( .A(n7026), .B(n7025), .Z(n7035) );
  NANDN U8064 ( .A(n6975), .B(n7484), .Z(n6979) );
  NAND U8065 ( .A(n6977), .B(n6976), .Z(n6978) );
  AND U8066 ( .A(n6979), .B(n6978), .Z(n7020) );
  AND U8067 ( .A(x[231]), .B(y[1863]), .Z(n7367) );
  NAND U8068 ( .A(n7479), .B(n7367), .Z(n6983) );
  NAND U8069 ( .A(n6981), .B(n6980), .Z(n6982) );
  AND U8070 ( .A(n6983), .B(n6982), .Z(n7018) );
  AND U8071 ( .A(y[1856]), .B(x[232]), .Z(n6985) );
  NAND U8072 ( .A(y[1864]), .B(x[224]), .Z(n6984) );
  XNOR U8073 ( .A(n6985), .B(n6984), .Z(n6995) );
  AND U8074 ( .A(x[231]), .B(y[1857]), .Z(n7000) );
  XOR U8075 ( .A(o[72]), .B(n7000), .Z(n6994) );
  XOR U8076 ( .A(n6995), .B(n6994), .Z(n7017) );
  NANDN U8077 ( .A(n6987), .B(n6986), .Z(n6991) );
  NAND U8078 ( .A(n6989), .B(n6988), .Z(n6990) );
  NAND U8079 ( .A(n6991), .B(n6990), .Z(n7032) );
  XNOR U8080 ( .A(n7029), .B(n7031), .Z(n6992) );
  XOR U8081 ( .A(n7030), .B(n6992), .Z(N169) );
  AND U8082 ( .A(x[232]), .B(y[1864]), .Z(n6993) );
  NAND U8083 ( .A(n6993), .B(n7479), .Z(n6997) );
  NAND U8084 ( .A(n6995), .B(n6994), .Z(n6996) );
  AND U8085 ( .A(n6997), .B(n6996), .Z(n7087) );
  AND U8086 ( .A(y[1860]), .B(x[229]), .Z(n6999) );
  NAND U8087 ( .A(y[1858]), .B(x[231]), .Z(n6998) );
  XNOR U8088 ( .A(n6999), .B(n6998), .Z(n7060) );
  AND U8089 ( .A(o[72]), .B(n7000), .Z(n7059) );
  XNOR U8090 ( .A(n7060), .B(n7059), .Z(n7085) );
  AND U8091 ( .A(y[1856]), .B(x[233]), .Z(n7002) );
  NAND U8092 ( .A(y[1865]), .B(x[224]), .Z(n7001) );
  XNOR U8093 ( .A(n7002), .B(n7001), .Z(n7067) );
  AND U8094 ( .A(x[232]), .B(y[1857]), .Z(n7076) );
  XOR U8095 ( .A(o[73]), .B(n7076), .Z(n7066) );
  XNOR U8096 ( .A(n7067), .B(n7066), .Z(n7084) );
  XOR U8097 ( .A(n7085), .B(n7084), .Z(n7086) );
  XNOR U8098 ( .A(n7087), .B(n7086), .Z(n7081) );
  AND U8099 ( .A(y[1859]), .B(x[230]), .Z(n7423) );
  NAND U8100 ( .A(y[1864]), .B(x[225]), .Z(n7003) );
  XNOR U8101 ( .A(n7423), .B(n7003), .Z(n7071) );
  XNOR U8102 ( .A(n7484), .B(n7071), .Z(n7091) );
  NAND U8103 ( .A(x[226]), .B(y[1863]), .Z(n7737) );
  AND U8104 ( .A(x[227]), .B(y[1862]), .Z(n7433) );
  XNOR U8105 ( .A(n7737), .B(n7433), .Z(n7090) );
  XNOR U8106 ( .A(n7091), .B(n7090), .Z(n7079) );
  NAND U8107 ( .A(x[229]), .B(y[1863]), .Z(n7258) );
  AND U8108 ( .A(x[225]), .B(y[1859]), .Z(n7070) );
  NANDN U8109 ( .A(n7258), .B(n7070), .Z(n7007) );
  NAND U8110 ( .A(n7005), .B(n7004), .Z(n7006) );
  NAND U8111 ( .A(n7007), .B(n7006), .Z(n7078) );
  XOR U8112 ( .A(n7079), .B(n7078), .Z(n7080) );
  XNOR U8113 ( .A(n7081), .B(n7080), .Z(n7054) );
  NAND U8114 ( .A(n7815), .B(n7008), .Z(n7012) );
  NANDN U8115 ( .A(n7010), .B(n7009), .Z(n7011) );
  NAND U8116 ( .A(n7012), .B(n7011), .Z(n7053) );
  NAND U8117 ( .A(n7192), .B(n7013), .Z(n7016) );
  NAND U8118 ( .A(n7690), .B(n7014), .Z(n7015) );
  AND U8119 ( .A(n7016), .B(n7015), .Z(n7052) );
  XOR U8120 ( .A(n7053), .B(n7052), .Z(n7055) );
  XNOR U8121 ( .A(n7054), .B(n7055), .Z(n7041) );
  NANDN U8122 ( .A(n7018), .B(n7017), .Z(n7022) );
  NANDN U8123 ( .A(n7020), .B(n7019), .Z(n7021) );
  AND U8124 ( .A(n7022), .B(n7021), .Z(n7040) );
  NANDN U8125 ( .A(n7024), .B(n7023), .Z(n7028) );
  NAND U8126 ( .A(n7026), .B(n7025), .Z(n7027) );
  NAND U8127 ( .A(n7028), .B(n7027), .Z(n7039) );
  XNOR U8128 ( .A(n7041), .B(n7042), .Z(n7048) );
  NANDN U8129 ( .A(n7033), .B(n7032), .Z(n7037) );
  NANDN U8130 ( .A(n7035), .B(n7034), .Z(n7036) );
  AND U8131 ( .A(n7037), .B(n7036), .Z(n7046) );
  IV U8132 ( .A(n7046), .Z(n7045) );
  XOR U8133 ( .A(n7047), .B(n7045), .Z(n7038) );
  XNOR U8134 ( .A(n7048), .B(n7038), .Z(N170) );
  NANDN U8135 ( .A(n7040), .B(n7039), .Z(n7044) );
  NAND U8136 ( .A(n7042), .B(n7041), .Z(n7043) );
  NAND U8137 ( .A(n7044), .B(n7043), .Z(n7102) );
  IV U8138 ( .A(n7102), .Z(n7101) );
  OR U8139 ( .A(n7047), .B(n7045), .Z(n7051) );
  ANDN U8140 ( .B(n7047), .A(n7046), .Z(n7049) );
  OR U8141 ( .A(n7049), .B(n7048), .Z(n7050) );
  AND U8142 ( .A(n7051), .B(n7050), .Z(n7103) );
  NAND U8143 ( .A(n7053), .B(n7052), .Z(n7057) );
  NAND U8144 ( .A(n7055), .B(n7054), .Z(n7056) );
  NAND U8145 ( .A(n7057), .B(n7056), .Z(n7098) );
  AND U8146 ( .A(x[231]), .B(y[1860]), .Z(n7144) );
  NAND U8147 ( .A(n7144), .B(n7058), .Z(n7062) );
  NAND U8148 ( .A(n7060), .B(n7059), .Z(n7061) );
  AND U8149 ( .A(n7062), .B(n7061), .Z(n7157) );
  AND U8150 ( .A(y[1859]), .B(x[231]), .Z(n7064) );
  NAND U8151 ( .A(y[1862]), .B(x[228]), .Z(n7063) );
  XNOR U8152 ( .A(n7064), .B(n7063), .Z(n7127) );
  AND U8153 ( .A(x[230]), .B(y[1860]), .Z(n7128) );
  XOR U8154 ( .A(n7127), .B(n7128), .Z(n7155) );
  AND U8155 ( .A(x[232]), .B(y[1858]), .Z(n7340) );
  AND U8156 ( .A(x[233]), .B(y[1857]), .Z(n7138) );
  XOR U8157 ( .A(o[74]), .B(n7138), .Z(n7149) );
  XOR U8158 ( .A(n7340), .B(n7149), .Z(n7151) );
  XNOR U8159 ( .A(n7151), .B(n7150), .Z(n7154) );
  XNOR U8160 ( .A(n7157), .B(n7156), .Z(n7117) );
  AND U8161 ( .A(x[233]), .B(y[1865]), .Z(n7065) );
  NAND U8162 ( .A(n7065), .B(n7479), .Z(n7069) );
  NAND U8163 ( .A(n7067), .B(n7066), .Z(n7068) );
  NAND U8164 ( .A(n7069), .B(n7068), .Z(n7115) );
  AND U8165 ( .A(x[230]), .B(y[1864]), .Z(n7377) );
  NAND U8166 ( .A(n7377), .B(n7070), .Z(n7073) );
  NAND U8167 ( .A(n7484), .B(n7071), .Z(n7072) );
  NAND U8168 ( .A(n7073), .B(n7072), .Z(n7123) );
  AND U8169 ( .A(y[1856]), .B(x[234]), .Z(n7075) );
  NAND U8170 ( .A(y[1866]), .B(x[224]), .Z(n7074) );
  XNOR U8171 ( .A(n7075), .B(n7074), .Z(n7133) );
  AND U8172 ( .A(o[73]), .B(n7076), .Z(n7132) );
  XOR U8173 ( .A(n7133), .B(n7132), .Z(n7121) );
  AND U8174 ( .A(y[1863]), .B(x[227]), .Z(n8048) );
  NAND U8175 ( .A(y[1865]), .B(x[225]), .Z(n7077) );
  XNOR U8176 ( .A(n8048), .B(n7077), .Z(n7145) );
  AND U8177 ( .A(x[226]), .B(y[1864]), .Z(n7146) );
  XOR U8178 ( .A(n7145), .B(n7146), .Z(n7120) );
  XOR U8179 ( .A(n7121), .B(n7120), .Z(n7122) );
  XOR U8180 ( .A(n7123), .B(n7122), .Z(n7114) );
  XOR U8181 ( .A(n7115), .B(n7114), .Z(n7116) );
  XNOR U8182 ( .A(n7117), .B(n7116), .Z(n7096) );
  NAND U8183 ( .A(n7079), .B(n7078), .Z(n7083) );
  NAND U8184 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U8185 ( .A(n7083), .B(n7082), .Z(n7111) );
  NAND U8186 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U8187 ( .A(n7087), .B(n7086), .Z(n7088) );
  AND U8188 ( .A(n7089), .B(n7088), .Z(n7108) );
  NAND U8189 ( .A(n7091), .B(n7090), .Z(n7093) );
  ANDN U8190 ( .B(n7737), .A(n7433), .Z(n7092) );
  ANDN U8191 ( .B(n7093), .A(n7092), .Z(n7109) );
  XOR U8192 ( .A(n7108), .B(n7109), .Z(n7110) );
  XOR U8193 ( .A(n7111), .B(n7110), .Z(n7095) );
  XOR U8194 ( .A(n7096), .B(n7095), .Z(n7097) );
  XOR U8195 ( .A(n7098), .B(n7097), .Z(n7104) );
  XNOR U8196 ( .A(n7103), .B(n7104), .Z(n7094) );
  XOR U8197 ( .A(n7101), .B(n7094), .Z(N171) );
  NAND U8198 ( .A(n7096), .B(n7095), .Z(n7100) );
  NAND U8199 ( .A(n7098), .B(n7097), .Z(n7099) );
  NAND U8200 ( .A(n7100), .B(n7099), .Z(n7224) );
  IV U8201 ( .A(n7224), .Z(n7222) );
  OR U8202 ( .A(n7103), .B(n7101), .Z(n7107) );
  ANDN U8203 ( .B(n7103), .A(n7102), .Z(n7105) );
  OR U8204 ( .A(n7105), .B(n7104), .Z(n7106) );
  AND U8205 ( .A(n7107), .B(n7106), .Z(n7223) );
  NAND U8206 ( .A(n7109), .B(n7108), .Z(n7113) );
  NANDN U8207 ( .A(n7111), .B(n7110), .Z(n7112) );
  NAND U8208 ( .A(n7113), .B(n7112), .Z(n7219) );
  NAND U8209 ( .A(n7115), .B(n7114), .Z(n7119) );
  NAND U8210 ( .A(n7117), .B(n7116), .Z(n7118) );
  NAND U8211 ( .A(n7119), .B(n7118), .Z(n7217) );
  NAND U8212 ( .A(n7121), .B(n7120), .Z(n7125) );
  NAND U8213 ( .A(n7123), .B(n7122), .Z(n7124) );
  NAND U8214 ( .A(n7125), .B(n7124), .Z(n7213) );
  AND U8215 ( .A(x[231]), .B(y[1862]), .Z(n7254) );
  AND U8216 ( .A(x[228]), .B(y[1859]), .Z(n7126) );
  NAND U8217 ( .A(n7254), .B(n7126), .Z(n7130) );
  NAND U8218 ( .A(n7128), .B(n7127), .Z(n7129) );
  NAND U8219 ( .A(n7130), .B(n7129), .Z(n7211) );
  AND U8220 ( .A(x[234]), .B(y[1866]), .Z(n7131) );
  NAND U8221 ( .A(n7131), .B(n7479), .Z(n7135) );
  NAND U8222 ( .A(n7133), .B(n7132), .Z(n7134) );
  NAND U8223 ( .A(n7135), .B(n7134), .Z(n7207) );
  AND U8224 ( .A(y[1856]), .B(x[235]), .Z(n7137) );
  NAND U8225 ( .A(y[1867]), .B(x[224]), .Z(n7136) );
  XNOR U8226 ( .A(n7137), .B(n7136), .Z(n7182) );
  AND U8227 ( .A(o[74]), .B(n7138), .Z(n7181) );
  XOR U8228 ( .A(n7182), .B(n7181), .Z(n7205) );
  AND U8229 ( .A(y[1861]), .B(x[230]), .Z(n7140) );
  NAND U8230 ( .A(y[1866]), .B(x[225]), .Z(n7139) );
  XNOR U8231 ( .A(n7140), .B(n7139), .Z(n7173) );
  AND U8232 ( .A(x[234]), .B(y[1857]), .Z(n7190) );
  XOR U8233 ( .A(o[75]), .B(n7190), .Z(n7172) );
  XOR U8234 ( .A(n7173), .B(n7172), .Z(n7204) );
  XOR U8235 ( .A(n7205), .B(n7204), .Z(n7206) );
  XOR U8236 ( .A(n7207), .B(n7206), .Z(n7210) );
  XOR U8237 ( .A(n7211), .B(n7210), .Z(n7212) );
  XNOR U8238 ( .A(n7213), .B(n7212), .Z(n7195) );
  AND U8239 ( .A(x[227]), .B(y[1864]), .Z(n8181) );
  NAND U8240 ( .A(y[1865]), .B(x[226]), .Z(n7141) );
  XNOR U8241 ( .A(n7142), .B(n7141), .Z(n7168) );
  AND U8242 ( .A(x[228]), .B(y[1863]), .Z(n7167) );
  XNOR U8243 ( .A(n7168), .B(n7167), .Z(n7199) );
  XNOR U8244 ( .A(n8181), .B(n7199), .Z(n7201) );
  NAND U8245 ( .A(y[1858]), .B(x[233]), .Z(n7143) );
  XNOR U8246 ( .A(n7144), .B(n7143), .Z(n7187) );
  AND U8247 ( .A(x[232]), .B(y[1859]), .Z(n7186) );
  XNOR U8248 ( .A(n7187), .B(n7186), .Z(n7200) );
  XNOR U8249 ( .A(n7201), .B(n7200), .Z(n7164) );
  NAND U8250 ( .A(x[227]), .B(y[1865]), .Z(n7249) );
  AND U8251 ( .A(x[225]), .B(y[1863]), .Z(n7474) );
  NANDN U8252 ( .A(n7249), .B(n7474), .Z(n7148) );
  NAND U8253 ( .A(n7146), .B(n7145), .Z(n7147) );
  NAND U8254 ( .A(n7148), .B(n7147), .Z(n7162) );
  NAND U8255 ( .A(n7340), .B(n7149), .Z(n7153) );
  NAND U8256 ( .A(n7151), .B(n7150), .Z(n7152) );
  NAND U8257 ( .A(n7153), .B(n7152), .Z(n7161) );
  XOR U8258 ( .A(n7162), .B(n7161), .Z(n7163) );
  XOR U8259 ( .A(n7164), .B(n7163), .Z(n7194) );
  NANDN U8260 ( .A(n7155), .B(n7154), .Z(n7159) );
  NAND U8261 ( .A(n7157), .B(n7156), .Z(n7158) );
  NAND U8262 ( .A(n7159), .B(n7158), .Z(n7193) );
  XOR U8263 ( .A(n7195), .B(n7196), .Z(n7216) );
  XOR U8264 ( .A(n7217), .B(n7216), .Z(n7218) );
  XOR U8265 ( .A(n7219), .B(n7218), .Z(n7225) );
  XNOR U8266 ( .A(n7223), .B(n7225), .Z(n7160) );
  XOR U8267 ( .A(n7222), .B(n7160), .Z(N172) );
  NAND U8268 ( .A(n7162), .B(n7161), .Z(n7166) );
  NAND U8269 ( .A(n7164), .B(n7163), .Z(n7165) );
  NAND U8270 ( .A(n7166), .B(n7165), .Z(n7290) );
  AND U8271 ( .A(x[226]), .B(y[1862]), .Z(n7929) );
  AND U8272 ( .A(x[229]), .B(y[1865]), .Z(n7728) );
  NAND U8273 ( .A(n7929), .B(n7728), .Z(n7170) );
  NAND U8274 ( .A(n7168), .B(n7167), .Z(n7169) );
  NAND U8275 ( .A(n7170), .B(n7169), .Z(n7237) );
  AND U8276 ( .A(x[230]), .B(y[1866]), .Z(n7491) );
  NAND U8277 ( .A(n7491), .B(n7171), .Z(n7175) );
  NAND U8278 ( .A(n7173), .B(n7172), .Z(n7174) );
  NAND U8279 ( .A(n7175), .B(n7174), .Z(n7236) );
  XOR U8280 ( .A(n7237), .B(n7236), .Z(n7239) );
  AND U8281 ( .A(x[233]), .B(y[1859]), .Z(n7924) );
  AND U8282 ( .A(y[1858]), .B(x[234]), .Z(n7907) );
  NAND U8283 ( .A(y[1864]), .B(x[228]), .Z(n7176) );
  XNOR U8284 ( .A(n7907), .B(n7176), .Z(n7280) );
  XOR U8285 ( .A(n7924), .B(n7280), .Z(n7259) );
  NAND U8286 ( .A(x[231]), .B(y[1861]), .Z(n7257) );
  XOR U8287 ( .A(n7258), .B(n7257), .Z(n7260) );
  AND U8288 ( .A(y[1856]), .B(x[236]), .Z(n7178) );
  NAND U8289 ( .A(y[1868]), .B(x[224]), .Z(n7177) );
  XNOR U8290 ( .A(n7178), .B(n7177), .Z(n7274) );
  AND U8291 ( .A(x[235]), .B(y[1857]), .Z(n7252) );
  XOR U8292 ( .A(o[76]), .B(n7252), .Z(n7273) );
  XOR U8293 ( .A(n7274), .B(n7273), .Z(n7243) );
  AND U8294 ( .A(y[1866]), .B(x[226]), .Z(n7180) );
  NAND U8295 ( .A(y[1860]), .B(x[232]), .Z(n7179) );
  XNOR U8296 ( .A(n7180), .B(n7179), .Z(n7248) );
  XOR U8297 ( .A(n7243), .B(n7242), .Z(n7245) );
  XOR U8298 ( .A(n7244), .B(n7245), .Z(n7238) );
  XOR U8299 ( .A(n7239), .B(n7238), .Z(n7288) );
  AND U8300 ( .A(x[235]), .B(y[1867]), .Z(n8309) );
  NAND U8301 ( .A(n8309), .B(n7479), .Z(n7184) );
  NAND U8302 ( .A(n7182), .B(n7181), .Z(n7183) );
  NAND U8303 ( .A(n7184), .B(n7183), .Z(n7266) );
  AND U8304 ( .A(x[231]), .B(y[1858]), .Z(n7409) );
  AND U8305 ( .A(x[233]), .B(y[1860]), .Z(n7185) );
  NAND U8306 ( .A(n7409), .B(n7185), .Z(n7189) );
  NAND U8307 ( .A(n7187), .B(n7186), .Z(n7188) );
  NAND U8308 ( .A(n7189), .B(n7188), .Z(n7264) );
  AND U8309 ( .A(o[75]), .B(n7190), .Z(n7269) );
  NAND U8310 ( .A(y[1867]), .B(x[225]), .Z(n7191) );
  XNOR U8311 ( .A(n7192), .B(n7191), .Z(n7270) );
  XOR U8312 ( .A(n7269), .B(n7270), .Z(n7263) );
  XOR U8313 ( .A(n7264), .B(n7263), .Z(n7265) );
  XOR U8314 ( .A(n7266), .B(n7265), .Z(n7287) );
  XOR U8315 ( .A(n7288), .B(n7287), .Z(n7289) );
  XOR U8316 ( .A(n7290), .B(n7289), .Z(n7297) );
  NANDN U8317 ( .A(n7194), .B(n7193), .Z(n7198) );
  NANDN U8318 ( .A(n7196), .B(n7195), .Z(n7197) );
  NAND U8319 ( .A(n7198), .B(n7197), .Z(n7296) );
  NANDN U8320 ( .A(n8181), .B(n7199), .Z(n7203) );
  NAND U8321 ( .A(n7201), .B(n7200), .Z(n7202) );
  NAND U8322 ( .A(n7203), .B(n7202), .Z(n7231) );
  NAND U8323 ( .A(n7205), .B(n7204), .Z(n7209) );
  NAND U8324 ( .A(n7207), .B(n7206), .Z(n7208) );
  AND U8325 ( .A(n7209), .B(n7208), .Z(n7230) );
  XOR U8326 ( .A(n7231), .B(n7230), .Z(n7233) );
  NAND U8327 ( .A(n7211), .B(n7210), .Z(n7215) );
  NAND U8328 ( .A(n7213), .B(n7212), .Z(n7214) );
  AND U8329 ( .A(n7215), .B(n7214), .Z(n7232) );
  XOR U8330 ( .A(n7233), .B(n7232), .Z(n7298) );
  XOR U8331 ( .A(n7299), .B(n7298), .Z(n7295) );
  NAND U8332 ( .A(n7217), .B(n7216), .Z(n7221) );
  NAND U8333 ( .A(n7219), .B(n7218), .Z(n7220) );
  NAND U8334 ( .A(n7221), .B(n7220), .Z(n7294) );
  NANDN U8335 ( .A(n7222), .B(n7223), .Z(n7228) );
  NOR U8336 ( .A(n7224), .B(n7223), .Z(n7226) );
  OR U8337 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U8338 ( .A(n7228), .B(n7227), .Z(n7293) );
  XOR U8339 ( .A(n7294), .B(n7293), .Z(n7229) );
  XNOR U8340 ( .A(n7295), .B(n7229), .Z(N173) );
  NAND U8341 ( .A(n7231), .B(n7230), .Z(n7235) );
  NAND U8342 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U8343 ( .A(n7235), .B(n7234), .Z(n7306) );
  NAND U8344 ( .A(n7237), .B(n7236), .Z(n7241) );
  NAND U8345 ( .A(n7239), .B(n7238), .Z(n7240) );
  NAND U8346 ( .A(n7241), .B(n7240), .Z(n7317) );
  NAND U8347 ( .A(n7243), .B(n7242), .Z(n7247) );
  NAND U8348 ( .A(n7245), .B(n7244), .Z(n7246) );
  NAND U8349 ( .A(n7247), .B(n7246), .Z(n7324) );
  AND U8350 ( .A(y[1866]), .B(x[232]), .Z(n8549) );
  AND U8351 ( .A(x[226]), .B(y[1860]), .Z(n7419) );
  NAND U8352 ( .A(n8549), .B(n7419), .Z(n7251) );
  NANDN U8353 ( .A(n7249), .B(n7248), .Z(n7250) );
  NAND U8354 ( .A(n7251), .B(n7250), .Z(n7356) );
  AND U8355 ( .A(o[76]), .B(n7252), .Z(n7346) );
  AND U8356 ( .A(y[1868]), .B(x[225]), .Z(n7253) );
  XOR U8357 ( .A(n7254), .B(n7253), .Z(n7345) );
  XOR U8358 ( .A(n7346), .B(n7345), .Z(n7354) );
  AND U8359 ( .A(x[230]), .B(y[1863]), .Z(n8349) );
  AND U8360 ( .A(y[1867]), .B(x[226]), .Z(n7256) );
  NAND U8361 ( .A(y[1860]), .B(x[233]), .Z(n7255) );
  XNOR U8362 ( .A(n7256), .B(n7255), .Z(n7360) );
  XOR U8363 ( .A(n8349), .B(n7360), .Z(n7353) );
  XOR U8364 ( .A(n7354), .B(n7353), .Z(n7355) );
  XOR U8365 ( .A(n7356), .B(n7355), .Z(n7323) );
  NAND U8366 ( .A(n7258), .B(n7257), .Z(n7262) );
  ANDN U8367 ( .B(n7260), .A(n7259), .Z(n7261) );
  ANDN U8368 ( .B(n7262), .A(n7261), .Z(n7322) );
  XOR U8369 ( .A(n7323), .B(n7322), .Z(n7325) );
  XOR U8370 ( .A(n7324), .B(n7325), .Z(n7316) );
  XOR U8371 ( .A(n7317), .B(n7316), .Z(n7319) );
  NAND U8372 ( .A(n7264), .B(n7263), .Z(n7268) );
  NAND U8373 ( .A(n7266), .B(n7265), .Z(n7267) );
  NAND U8374 ( .A(n7268), .B(n7267), .Z(n7331) );
  AND U8375 ( .A(x[230]), .B(y[1867]), .Z(n7729) );
  AND U8376 ( .A(x[225]), .B(y[1862]), .Z(n7344) );
  NAND U8377 ( .A(n7729), .B(n7344), .Z(n7272) );
  NAND U8378 ( .A(n7270), .B(n7269), .Z(n7271) );
  NAND U8379 ( .A(n7272), .B(n7271), .Z(n7337) );
  AND U8380 ( .A(x[236]), .B(y[1868]), .Z(n8555) );
  NAND U8381 ( .A(n8555), .B(n7479), .Z(n7276) );
  NAND U8382 ( .A(n7274), .B(n7273), .Z(n7275) );
  NAND U8383 ( .A(n7276), .B(n7275), .Z(n7335) );
  AND U8384 ( .A(x[234]), .B(y[1859]), .Z(n8193) );
  AND U8385 ( .A(y[1858]), .B(x[235]), .Z(n8154) );
  NAND U8386 ( .A(y[1861]), .B(x[232]), .Z(n7277) );
  XNOR U8387 ( .A(n8154), .B(n7277), .Z(n7341) );
  XOR U8388 ( .A(n8193), .B(n7341), .Z(n7334) );
  XOR U8389 ( .A(n7335), .B(n7334), .Z(n7336) );
  XOR U8390 ( .A(n7337), .B(n7336), .Z(n7329) );
  AND U8391 ( .A(x[234]), .B(y[1864]), .Z(n7279) );
  AND U8392 ( .A(x[228]), .B(y[1858]), .Z(n7278) );
  NAND U8393 ( .A(n7279), .B(n7278), .Z(n7282) );
  NAND U8394 ( .A(n7280), .B(n7924), .Z(n7281) );
  NAND U8395 ( .A(n7282), .B(n7281), .Z(n7381) );
  AND U8396 ( .A(y[1856]), .B(x[237]), .Z(n7284) );
  NAND U8397 ( .A(y[1869]), .B(x[224]), .Z(n7283) );
  XNOR U8398 ( .A(n7284), .B(n7283), .Z(n7373) );
  AND U8399 ( .A(x[236]), .B(y[1857]), .Z(n7365) );
  XOR U8400 ( .A(o[77]), .B(n7365), .Z(n7372) );
  XOR U8401 ( .A(n7373), .B(n7372), .Z(n7379) );
  AND U8402 ( .A(y[1864]), .B(x[229]), .Z(n7286) );
  NAND U8403 ( .A(y[1866]), .B(x[227]), .Z(n7285) );
  XNOR U8404 ( .A(n7286), .B(n7285), .Z(n7368) );
  AND U8405 ( .A(x[228]), .B(y[1865]), .Z(n7369) );
  XOR U8406 ( .A(n7368), .B(n7369), .Z(n7378) );
  XOR U8407 ( .A(n7379), .B(n7378), .Z(n7380) );
  XOR U8408 ( .A(n7381), .B(n7380), .Z(n7328) );
  XOR U8409 ( .A(n7329), .B(n7328), .Z(n7330) );
  XOR U8410 ( .A(n7331), .B(n7330), .Z(n7318) );
  XNOR U8411 ( .A(n7319), .B(n7318), .Z(n7304) );
  NAND U8412 ( .A(n7288), .B(n7287), .Z(n7292) );
  NAND U8413 ( .A(n7290), .B(n7289), .Z(n7291) );
  AND U8414 ( .A(n7292), .B(n7291), .Z(n7303) );
  XOR U8415 ( .A(n7304), .B(n7303), .Z(n7305) );
  XOR U8416 ( .A(n7306), .B(n7305), .Z(n7312) );
  NANDN U8417 ( .A(n7297), .B(n7296), .Z(n7301) );
  NAND U8418 ( .A(n7299), .B(n7298), .Z(n7300) );
  AND U8419 ( .A(n7301), .B(n7300), .Z(n7310) );
  IV U8420 ( .A(n7310), .Z(n7309) );
  XOR U8421 ( .A(n7311), .B(n7309), .Z(n7302) );
  XNOR U8422 ( .A(n7312), .B(n7302), .Z(N174) );
  NAND U8423 ( .A(n7304), .B(n7303), .Z(n7308) );
  NAND U8424 ( .A(n7306), .B(n7305), .Z(n7307) );
  NAND U8425 ( .A(n7308), .B(n7307), .Z(n7468) );
  IV U8426 ( .A(n7468), .Z(n7466) );
  OR U8427 ( .A(n7311), .B(n7309), .Z(n7315) );
  ANDN U8428 ( .B(n7311), .A(n7310), .Z(n7313) );
  OR U8429 ( .A(n7313), .B(n7312), .Z(n7314) );
  AND U8430 ( .A(n7315), .B(n7314), .Z(n7467) );
  NAND U8431 ( .A(n7317), .B(n7316), .Z(n7321) );
  NAND U8432 ( .A(n7319), .B(n7318), .Z(n7320) );
  NAND U8433 ( .A(n7321), .B(n7320), .Z(n7461) );
  NAND U8434 ( .A(n7323), .B(n7322), .Z(n7327) );
  NAND U8435 ( .A(n7325), .B(n7324), .Z(n7326) );
  NAND U8436 ( .A(n7327), .B(n7326), .Z(n7460) );
  XOR U8437 ( .A(n7461), .B(n7460), .Z(n7463) );
  NAND U8438 ( .A(n7329), .B(n7328), .Z(n7333) );
  NAND U8439 ( .A(n7331), .B(n7330), .Z(n7332) );
  NAND U8440 ( .A(n7333), .B(n7332), .Z(n7388) );
  NAND U8441 ( .A(n7335), .B(n7334), .Z(n7339) );
  NAND U8442 ( .A(n7337), .B(n7336), .Z(n7338) );
  AND U8443 ( .A(n7339), .B(n7338), .Z(n7394) );
  AND U8444 ( .A(x[235]), .B(y[1861]), .Z(n7505) );
  NAND U8445 ( .A(n7505), .B(n7340), .Z(n7343) );
  NAND U8446 ( .A(n7341), .B(n8193), .Z(n7342) );
  NAND U8447 ( .A(n7343), .B(n7342), .Z(n7449) );
  NAND U8448 ( .A(x[231]), .B(y[1868]), .Z(n7939) );
  NANDN U8449 ( .A(n7939), .B(n7344), .Z(n7348) );
  NAND U8450 ( .A(n7346), .B(n7345), .Z(n7347) );
  NAND U8451 ( .A(n7348), .B(n7347), .Z(n7448) );
  XOR U8452 ( .A(n7449), .B(n7448), .Z(n7451) );
  AND U8453 ( .A(x[228]), .B(y[1866]), .Z(n7824) );
  AND U8454 ( .A(y[1867]), .B(x[227]), .Z(n7350) );
  NAND U8455 ( .A(y[1862]), .B(x[232]), .Z(n7349) );
  XNOR U8456 ( .A(n7350), .B(n7349), .Z(n7434) );
  XOR U8457 ( .A(n7728), .B(n7434), .Z(n7443) );
  XOR U8458 ( .A(n7824), .B(n7443), .Z(n7445) );
  AND U8459 ( .A(x[233]), .B(y[1861]), .Z(n8013) );
  AND U8460 ( .A(y[1868]), .B(x[226]), .Z(n7352) );
  NAND U8461 ( .A(y[1860]), .B(x[234]), .Z(n7351) );
  XNOR U8462 ( .A(n7352), .B(n7351), .Z(n7420) );
  XOR U8463 ( .A(n8013), .B(n7420), .Z(n7444) );
  XOR U8464 ( .A(n7445), .B(n7444), .Z(n7450) );
  XNOR U8465 ( .A(n7451), .B(n7450), .Z(n7392) );
  NAND U8466 ( .A(n7354), .B(n7353), .Z(n7358) );
  NAND U8467 ( .A(n7356), .B(n7355), .Z(n7357) );
  AND U8468 ( .A(n7358), .B(n7357), .Z(n7391) );
  XOR U8469 ( .A(n7392), .B(n7391), .Z(n7393) );
  XNOR U8470 ( .A(n7394), .B(n7393), .Z(n7386) );
  AND U8471 ( .A(x[233]), .B(y[1867]), .Z(n7359) );
  NAND U8472 ( .A(n7359), .B(n7419), .Z(n7362) );
  NAND U8473 ( .A(n7360), .B(n8349), .Z(n7361) );
  NAND U8474 ( .A(n7362), .B(n7361), .Z(n7405) );
  AND U8475 ( .A(y[1856]), .B(x[238]), .Z(n7364) );
  NAND U8476 ( .A(y[1870]), .B(x[224]), .Z(n7363) );
  XNOR U8477 ( .A(n7364), .B(n7363), .Z(n7429) );
  AND U8478 ( .A(o[77]), .B(n7365), .Z(n7428) );
  XOR U8479 ( .A(n7429), .B(n7428), .Z(n7404) );
  NAND U8480 ( .A(y[1858]), .B(x[236]), .Z(n7366) );
  XNOR U8481 ( .A(n7367), .B(n7366), .Z(n7411) );
  AND U8482 ( .A(x[237]), .B(y[1857]), .Z(n7418) );
  XOR U8483 ( .A(o[78]), .B(n7418), .Z(n7410) );
  XOR U8484 ( .A(n7411), .B(n7410), .Z(n7403) );
  XOR U8485 ( .A(n7404), .B(n7403), .Z(n7406) );
  XNOR U8486 ( .A(n7405), .B(n7406), .Z(n7455) );
  AND U8487 ( .A(x[229]), .B(y[1866]), .Z(n7492) );
  NAND U8488 ( .A(n8181), .B(n7492), .Z(n7371) );
  NAND U8489 ( .A(n7369), .B(n7368), .Z(n7370) );
  NAND U8490 ( .A(n7371), .B(n7370), .Z(n7399) );
  AND U8491 ( .A(x[237]), .B(y[1869]), .Z(n8944) );
  NAND U8492 ( .A(n8944), .B(n7479), .Z(n7375) );
  NAND U8493 ( .A(n7373), .B(n7372), .Z(n7374) );
  NAND U8494 ( .A(n7375), .B(n7374), .Z(n7397) );
  NAND U8495 ( .A(y[1859]), .B(x[235]), .Z(n7376) );
  XNOR U8496 ( .A(n7377), .B(n7376), .Z(n7425) );
  AND U8497 ( .A(x[225]), .B(y[1869]), .Z(n7424) );
  XOR U8498 ( .A(n7425), .B(n7424), .Z(n7398) );
  XNOR U8499 ( .A(n7397), .B(n7398), .Z(n7400) );
  XOR U8500 ( .A(n7399), .B(n7400), .Z(n7454) );
  XOR U8501 ( .A(n7455), .B(n7454), .Z(n7457) );
  NAND U8502 ( .A(n7379), .B(n7378), .Z(n7383) );
  NAND U8503 ( .A(n7381), .B(n7380), .Z(n7382) );
  AND U8504 ( .A(n7383), .B(n7382), .Z(n7456) );
  XNOR U8505 ( .A(n7457), .B(n7456), .Z(n7385) );
  XOR U8506 ( .A(n7386), .B(n7385), .Z(n7387) );
  XOR U8507 ( .A(n7388), .B(n7387), .Z(n7462) );
  XOR U8508 ( .A(n7463), .B(n7462), .Z(n7469) );
  XNOR U8509 ( .A(n7467), .B(n7469), .Z(n7384) );
  XOR U8510 ( .A(n7466), .B(n7384), .Z(N175) );
  NAND U8511 ( .A(n7386), .B(n7385), .Z(n7390) );
  NAND U8512 ( .A(n7388), .B(n7387), .Z(n7389) );
  AND U8513 ( .A(n7390), .B(n7389), .Z(n7562) );
  NAND U8514 ( .A(n7392), .B(n7391), .Z(n7396) );
  NAND U8515 ( .A(n7394), .B(n7393), .Z(n7395) );
  NAND U8516 ( .A(n7396), .B(n7395), .Z(n7534) );
  NAND U8517 ( .A(n7398), .B(n7397), .Z(n7402) );
  NANDN U8518 ( .A(n7400), .B(n7399), .Z(n7401) );
  NAND U8519 ( .A(n7402), .B(n7401), .Z(n7540) );
  NAND U8520 ( .A(n7404), .B(n7403), .Z(n7408) );
  NAND U8521 ( .A(n7406), .B(n7405), .Z(n7407) );
  NAND U8522 ( .A(n7408), .B(n7407), .Z(n7538) );
  NAND U8523 ( .A(x[236]), .B(y[1863]), .Z(n7931) );
  NANDN U8524 ( .A(n7931), .B(n7409), .Z(n7413) );
  NAND U8525 ( .A(n7411), .B(n7410), .Z(n7412) );
  AND U8526 ( .A(n7413), .B(n7412), .Z(n7515) );
  AND U8527 ( .A(y[1860]), .B(x[235]), .Z(n7415) );
  NAND U8528 ( .A(y[1858]), .B(x[237]), .Z(n7414) );
  XNOR U8529 ( .A(n7415), .B(n7414), .Z(n7519) );
  AND U8530 ( .A(x[236]), .B(y[1859]), .Z(n7518) );
  XNOR U8531 ( .A(n7519), .B(n7518), .Z(n7513) );
  AND U8532 ( .A(y[1856]), .B(x[239]), .Z(n7417) );
  NAND U8533 ( .A(y[1871]), .B(x[224]), .Z(n7416) );
  XNOR U8534 ( .A(n7417), .B(n7416), .Z(n7481) );
  AND U8535 ( .A(o[78]), .B(n7418), .Z(n7480) );
  XNOR U8536 ( .A(n7481), .B(n7480), .Z(n7512) );
  XOR U8537 ( .A(n7513), .B(n7512), .Z(n7514) );
  XOR U8538 ( .A(n7515), .B(n7514), .Z(n7547) );
  NAND U8539 ( .A(x[234]), .B(y[1868]), .Z(n8351) );
  NANDN U8540 ( .A(n8351), .B(n7419), .Z(n7422) );
  NAND U8541 ( .A(n8013), .B(n7420), .Z(n7421) );
  NAND U8542 ( .A(n7422), .B(n7421), .Z(n7545) );
  AND U8543 ( .A(x[235]), .B(y[1864]), .Z(n7823) );
  NAND U8544 ( .A(n7823), .B(n7423), .Z(n7427) );
  NAND U8545 ( .A(n7425), .B(n7424), .Z(n7426) );
  NAND U8546 ( .A(n7427), .B(n7426), .Z(n7544) );
  XOR U8547 ( .A(n7545), .B(n7544), .Z(n7546) );
  XOR U8548 ( .A(n7538), .B(n7539), .Z(n7541) );
  XOR U8549 ( .A(n7540), .B(n7541), .Z(n7533) );
  AND U8550 ( .A(x[238]), .B(y[1870]), .Z(n9209) );
  NAND U8551 ( .A(n9209), .B(n7479), .Z(n7431) );
  NAND U8552 ( .A(n7429), .B(n7428), .Z(n7430) );
  NAND U8553 ( .A(n7431), .B(n7430), .Z(n7507) );
  AND U8554 ( .A(x[232]), .B(y[1867]), .Z(n7432) );
  NAND U8555 ( .A(n7433), .B(n7432), .Z(n7436) );
  NAND U8556 ( .A(n7728), .B(n7434), .Z(n7435) );
  NAND U8557 ( .A(n7436), .B(n7435), .Z(n7506) );
  XOR U8558 ( .A(n7507), .B(n7506), .Z(n7509) );
  AND U8559 ( .A(y[1861]), .B(x[234]), .Z(n7438) );
  NAND U8560 ( .A(y[1867]), .B(x[228]), .Z(n7437) );
  XNOR U8561 ( .A(n7438), .B(n7437), .Z(n7487) );
  AND U8562 ( .A(x[231]), .B(y[1864]), .Z(n7486) );
  XNOR U8563 ( .A(n7487), .B(n7486), .Z(n7494) );
  NAND U8564 ( .A(x[230]), .B(y[1865]), .Z(n7606) );
  XNOR U8565 ( .A(n7606), .B(n7492), .Z(n7493) );
  XNOR U8566 ( .A(n7494), .B(n7493), .Z(n7528) );
  AND U8567 ( .A(y[1869]), .B(x[226]), .Z(n7440) );
  NAND U8568 ( .A(y[1862]), .B(x[233]), .Z(n7439) );
  XNOR U8569 ( .A(n7440), .B(n7439), .Z(n7497) );
  AND U8570 ( .A(x[227]), .B(y[1868]), .Z(n7498) );
  XOR U8571 ( .A(n7497), .B(n7498), .Z(n7527) );
  AND U8572 ( .A(y[1870]), .B(x[225]), .Z(n7442) );
  NAND U8573 ( .A(y[1863]), .B(x[232]), .Z(n7441) );
  XNOR U8574 ( .A(n7442), .B(n7441), .Z(n7476) );
  AND U8575 ( .A(x[238]), .B(y[1857]), .Z(n7503) );
  XOR U8576 ( .A(o[79]), .B(n7503), .Z(n7475) );
  XOR U8577 ( .A(n7476), .B(n7475), .Z(n7526) );
  XOR U8578 ( .A(n7527), .B(n7526), .Z(n7529) );
  XOR U8579 ( .A(n7528), .B(n7529), .Z(n7508) );
  XOR U8580 ( .A(n7509), .B(n7508), .Z(n7551) );
  NAND U8581 ( .A(n7824), .B(n7443), .Z(n7447) );
  NAND U8582 ( .A(n7445), .B(n7444), .Z(n7446) );
  AND U8583 ( .A(n7447), .B(n7446), .Z(n7550) );
  NAND U8584 ( .A(n7449), .B(n7448), .Z(n7453) );
  NAND U8585 ( .A(n7451), .B(n7450), .Z(n7452) );
  AND U8586 ( .A(n7453), .B(n7452), .Z(n7552) );
  XOR U8587 ( .A(n7553), .B(n7552), .Z(n7532) );
  XOR U8588 ( .A(n7534), .B(n7535), .Z(n7559) );
  NAND U8589 ( .A(n7455), .B(n7454), .Z(n7459) );
  NAND U8590 ( .A(n7457), .B(n7456), .Z(n7458) );
  AND U8591 ( .A(n7459), .B(n7458), .Z(n7560) );
  XOR U8592 ( .A(n7559), .B(n7560), .Z(n7561) );
  XOR U8593 ( .A(n7562), .B(n7561), .Z(n7558) );
  NAND U8594 ( .A(n7461), .B(n7460), .Z(n7465) );
  NAND U8595 ( .A(n7463), .B(n7462), .Z(n7464) );
  NAND U8596 ( .A(n7465), .B(n7464), .Z(n7557) );
  NANDN U8597 ( .A(n7466), .B(n7467), .Z(n7472) );
  NOR U8598 ( .A(n7468), .B(n7467), .Z(n7470) );
  OR U8599 ( .A(n7470), .B(n7469), .Z(n7471) );
  AND U8600 ( .A(n7472), .B(n7471), .Z(n7556) );
  XOR U8601 ( .A(n7557), .B(n7556), .Z(n7473) );
  XNOR U8602 ( .A(n7558), .B(n7473), .Z(N176) );
  AND U8603 ( .A(x[232]), .B(y[1870]), .Z(n7825) );
  NAND U8604 ( .A(n7825), .B(n7474), .Z(n7478) );
  NAND U8605 ( .A(n7476), .B(n7475), .Z(n7477) );
  NAND U8606 ( .A(n7478), .B(n7477), .Z(n7636) );
  AND U8607 ( .A(x[239]), .B(y[1871]), .Z(n9638) );
  NAND U8608 ( .A(n9638), .B(n7479), .Z(n7483) );
  NAND U8609 ( .A(n7481), .B(n7480), .Z(n7482) );
  NAND U8610 ( .A(n7483), .B(n7482), .Z(n7635) );
  XOR U8611 ( .A(n7636), .B(n7635), .Z(n7638) );
  AND U8612 ( .A(x[234]), .B(y[1867]), .Z(n7485) );
  NAND U8613 ( .A(n7485), .B(n7484), .Z(n7489) );
  NAND U8614 ( .A(n7487), .B(n7486), .Z(n7488) );
  NAND U8615 ( .A(n7489), .B(n7488), .Z(n7593) );
  AND U8616 ( .A(x[224]), .B(y[1872]), .Z(n7615) );
  AND U8617 ( .A(x[240]), .B(y[1856]), .Z(n7616) );
  XOR U8618 ( .A(n7615), .B(n7616), .Z(n7617) );
  NAND U8619 ( .A(x[239]), .B(y[1857]), .Z(n7603) );
  XNOR U8620 ( .A(o[80]), .B(n7603), .Z(n7618) );
  XOR U8621 ( .A(n7617), .B(n7618), .Z(n7592) );
  NAND U8622 ( .A(y[1865]), .B(x[231]), .Z(n7490) );
  XNOR U8623 ( .A(n7491), .B(n7490), .Z(n7608) );
  AND U8624 ( .A(x[234]), .B(y[1862]), .Z(n7607) );
  XOR U8625 ( .A(n7608), .B(n7607), .Z(n7591) );
  XOR U8626 ( .A(n7592), .B(n7591), .Z(n7594) );
  XOR U8627 ( .A(n7593), .B(n7594), .Z(n7637) );
  XNOR U8628 ( .A(n7638), .B(n7637), .Z(n7588) );
  NANDN U8629 ( .A(n7492), .B(n7606), .Z(n7496) );
  NAND U8630 ( .A(n7494), .B(n7493), .Z(n7495) );
  NAND U8631 ( .A(n7496), .B(n7495), .Z(n7586) );
  NAND U8632 ( .A(x[233]), .B(y[1869]), .Z(n8332) );
  NANDN U8633 ( .A(n8332), .B(n7929), .Z(n7500) );
  NAND U8634 ( .A(n7498), .B(n7497), .Z(n7499) );
  AND U8635 ( .A(n7500), .B(n7499), .Z(n7626) );
  AND U8636 ( .A(y[1871]), .B(x[225]), .Z(n7502) );
  NAND U8637 ( .A(y[1864]), .B(x[232]), .Z(n7501) );
  XNOR U8638 ( .A(n7502), .B(n7501), .Z(n7612) );
  AND U8639 ( .A(o[79]), .B(n7503), .Z(n7611) );
  XOR U8640 ( .A(n7612), .B(n7611), .Z(n7623) );
  NAND U8641 ( .A(y[1858]), .B(x[238]), .Z(n7504) );
  XNOR U8642 ( .A(n7505), .B(n7504), .Z(n7647) );
  NAND U8643 ( .A(x[228]), .B(y[1868]), .Z(n7648) );
  XNOR U8644 ( .A(n7647), .B(n7648), .Z(n7624) );
  XOR U8645 ( .A(n7623), .B(n7624), .Z(n7625) );
  XOR U8646 ( .A(n7626), .B(n7625), .Z(n7585) );
  XOR U8647 ( .A(n7586), .B(n7585), .Z(n7587) );
  XOR U8648 ( .A(n7588), .B(n7587), .Z(n7629) );
  NAND U8649 ( .A(n7507), .B(n7506), .Z(n7511) );
  NAND U8650 ( .A(n7509), .B(n7508), .Z(n7510) );
  AND U8651 ( .A(n7511), .B(n7510), .Z(n7630) );
  XOR U8652 ( .A(n7629), .B(n7630), .Z(n7632) );
  NAND U8653 ( .A(n7513), .B(n7512), .Z(n7517) );
  NAND U8654 ( .A(n7515), .B(n7514), .Z(n7516) );
  NAND U8655 ( .A(n7517), .B(n7516), .Z(n7661) );
  AND U8656 ( .A(x[237]), .B(y[1860]), .Z(n7657) );
  NAND U8657 ( .A(n8154), .B(n7657), .Z(n7521) );
  NAND U8658 ( .A(n7519), .B(n7518), .Z(n7520) );
  NAND U8659 ( .A(n7521), .B(n7520), .Z(n7644) );
  AND U8660 ( .A(y[1870]), .B(x[226]), .Z(n7523) );
  NAND U8661 ( .A(y[1863]), .B(x[233]), .Z(n7522) );
  XNOR U8662 ( .A(n7523), .B(n7522), .Z(n7651) );
  NAND U8663 ( .A(x[227]), .B(y[1869]), .Z(n7652) );
  XNOR U8664 ( .A(n7651), .B(n7652), .Z(n7642) );
  AND U8665 ( .A(x[236]), .B(y[1860]), .Z(n8320) );
  AND U8666 ( .A(y[1867]), .B(x[229]), .Z(n7525) );
  NAND U8667 ( .A(y[1859]), .B(x[237]), .Z(n7524) );
  XNOR U8668 ( .A(n7525), .B(n7524), .Z(n7598) );
  XOR U8669 ( .A(n8320), .B(n7598), .Z(n7641) );
  XOR U8670 ( .A(n7642), .B(n7641), .Z(n7643) );
  XNOR U8671 ( .A(n7644), .B(n7643), .Z(n7658) );
  NAND U8672 ( .A(n7527), .B(n7526), .Z(n7531) );
  NAND U8673 ( .A(n7529), .B(n7528), .Z(n7530) );
  AND U8674 ( .A(n7531), .B(n7530), .Z(n7659) );
  XOR U8675 ( .A(n7658), .B(n7659), .Z(n7660) );
  XOR U8676 ( .A(n7661), .B(n7660), .Z(n7631) );
  XOR U8677 ( .A(n7632), .B(n7631), .Z(n7567) );
  NANDN U8678 ( .A(n7533), .B(n7532), .Z(n7537) );
  NANDN U8679 ( .A(n7535), .B(n7534), .Z(n7536) );
  AND U8680 ( .A(n7537), .B(n7536), .Z(n7566) );
  NAND U8681 ( .A(n7539), .B(n7538), .Z(n7543) );
  NAND U8682 ( .A(n7541), .B(n7540), .Z(n7542) );
  NAND U8683 ( .A(n7543), .B(n7542), .Z(n7581) );
  NAND U8684 ( .A(n7545), .B(n7544), .Z(n7549) );
  NANDN U8685 ( .A(n7547), .B(n7546), .Z(n7548) );
  NAND U8686 ( .A(n7549), .B(n7548), .Z(n7579) );
  NANDN U8687 ( .A(n7551), .B(n7550), .Z(n7555) );
  NAND U8688 ( .A(n7553), .B(n7552), .Z(n7554) );
  AND U8689 ( .A(n7555), .B(n7554), .Z(n7580) );
  XNOR U8690 ( .A(n7579), .B(n7580), .Z(n7582) );
  XNOR U8691 ( .A(n7568), .B(n7569), .Z(n7575) );
  NAND U8692 ( .A(n7560), .B(n7559), .Z(n7564) );
  NANDN U8693 ( .A(n7562), .B(n7561), .Z(n7563) );
  AND U8694 ( .A(n7564), .B(n7563), .Z(n7574) );
  IV U8695 ( .A(n7574), .Z(n7572) );
  XOR U8696 ( .A(n7573), .B(n7572), .Z(n7565) );
  XNOR U8697 ( .A(n7575), .B(n7565), .Z(N177) );
  NANDN U8698 ( .A(n7567), .B(n7566), .Z(n7571) );
  NANDN U8699 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U8700 ( .A(n7571), .B(n7570), .Z(n7671) );
  NANDN U8701 ( .A(n7572), .B(n7573), .Z(n7578) );
  NOR U8702 ( .A(n7574), .B(n7573), .Z(n7576) );
  OR U8703 ( .A(n7576), .B(n7575), .Z(n7577) );
  AND U8704 ( .A(n7578), .B(n7577), .Z(n7672) );
  NAND U8705 ( .A(n7580), .B(n7579), .Z(n7584) );
  NANDN U8706 ( .A(n7582), .B(n7581), .Z(n7583) );
  NAND U8707 ( .A(n7584), .B(n7583), .Z(n7667) );
  NAND U8708 ( .A(n7586), .B(n7585), .Z(n7590) );
  NAND U8709 ( .A(n7588), .B(n7587), .Z(n7589) );
  NAND U8710 ( .A(n7590), .B(n7589), .Z(n7683) );
  NAND U8711 ( .A(n7592), .B(n7591), .Z(n7596) );
  NAND U8712 ( .A(n7594), .B(n7593), .Z(n7595) );
  NAND U8713 ( .A(n7596), .B(n7595), .Z(n7763) );
  AND U8714 ( .A(x[237]), .B(y[1867]), .Z(n8563) );
  NAND U8715 ( .A(n8563), .B(n7597), .Z(n7600) );
  NAND U8716 ( .A(n7598), .B(n8320), .Z(n7599) );
  NAND U8717 ( .A(n7600), .B(n7599), .Z(n7713) );
  AND U8718 ( .A(y[1872]), .B(x[225]), .Z(n7602) );
  NAND U8719 ( .A(y[1864]), .B(x[233]), .Z(n7601) );
  XNOR U8720 ( .A(n7602), .B(n7601), .Z(n7733) );
  NANDN U8721 ( .A(n7603), .B(o[80]), .Z(n7734) );
  XNOR U8722 ( .A(n7733), .B(n7734), .Z(n7711) );
  AND U8723 ( .A(y[1858]), .B(x[239]), .Z(n7605) );
  NAND U8724 ( .A(y[1861]), .B(x[236]), .Z(n7604) );
  XNOR U8725 ( .A(n7605), .B(n7604), .Z(n7686) );
  NAND U8726 ( .A(x[238]), .B(y[1859]), .Z(n7687) );
  XOR U8727 ( .A(n7711), .B(n7710), .Z(n7712) );
  XOR U8728 ( .A(n7713), .B(n7712), .Z(n7761) );
  AND U8729 ( .A(x[231]), .B(y[1866]), .Z(n7743) );
  NANDN U8730 ( .A(n7606), .B(n7743), .Z(n7610) );
  NAND U8731 ( .A(n7608), .B(n7607), .Z(n7609) );
  NAND U8732 ( .A(n7610), .B(n7609), .Z(n7723) );
  NAND U8733 ( .A(x[232]), .B(y[1871]), .Z(n8401) );
  AND U8734 ( .A(x[225]), .B(y[1864]), .Z(n7803) );
  NANDN U8735 ( .A(n8401), .B(n7803), .Z(n7614) );
  NAND U8736 ( .A(n7612), .B(n7611), .Z(n7613) );
  NAND U8737 ( .A(n7614), .B(n7613), .Z(n7722) );
  XOR U8738 ( .A(n7723), .B(n7722), .Z(n7725) );
  NAND U8739 ( .A(n7616), .B(n7615), .Z(n7620) );
  NAND U8740 ( .A(n7618), .B(n7617), .Z(n7619) );
  NAND U8741 ( .A(n7620), .B(n7619), .Z(n7719) );
  AND U8742 ( .A(x[224]), .B(y[1873]), .Z(n7700) );
  NAND U8743 ( .A(x[241]), .B(y[1856]), .Z(n7701) );
  NAND U8744 ( .A(x[240]), .B(y[1857]), .Z(n7697) );
  XOR U8745 ( .A(o[81]), .B(n7697), .Z(n7703) );
  AND U8746 ( .A(y[1871]), .B(x[226]), .Z(n7622) );
  NAND U8747 ( .A(y[1863]), .B(x[234]), .Z(n7621) );
  XNOR U8748 ( .A(n7622), .B(n7621), .Z(n7738) );
  NAND U8749 ( .A(x[227]), .B(y[1870]), .Z(n7739) );
  XNOR U8750 ( .A(n7738), .B(n7739), .Z(n7717) );
  XOR U8751 ( .A(n7716), .B(n7717), .Z(n7718) );
  XOR U8752 ( .A(n7719), .B(n7718), .Z(n7724) );
  XOR U8753 ( .A(n7725), .B(n7724), .Z(n7760) );
  XOR U8754 ( .A(n7761), .B(n7760), .Z(n7762) );
  XNOR U8755 ( .A(n7763), .B(n7762), .Z(n7680) );
  NAND U8756 ( .A(n7624), .B(n7623), .Z(n7628) );
  NANDN U8757 ( .A(n7626), .B(n7625), .Z(n7627) );
  AND U8758 ( .A(n7628), .B(n7627), .Z(n7681) );
  XOR U8759 ( .A(n7680), .B(n7681), .Z(n7682) );
  XOR U8760 ( .A(n7683), .B(n7682), .Z(n7666) );
  NAND U8761 ( .A(n7630), .B(n7629), .Z(n7634) );
  NAND U8762 ( .A(n7632), .B(n7631), .Z(n7633) );
  AND U8763 ( .A(n7634), .B(n7633), .Z(n7677) );
  NAND U8764 ( .A(n7636), .B(n7635), .Z(n7640) );
  NAND U8765 ( .A(n7638), .B(n7637), .Z(n7639) );
  NAND U8766 ( .A(n7640), .B(n7639), .Z(n7757) );
  NAND U8767 ( .A(n7642), .B(n7641), .Z(n7646) );
  NAND U8768 ( .A(n7644), .B(n7643), .Z(n7645) );
  NAND U8769 ( .A(n7646), .B(n7645), .Z(n7755) );
  NAND U8770 ( .A(x[238]), .B(y[1861]), .Z(n7904) );
  NANDN U8771 ( .A(n7904), .B(n8154), .Z(n7650) );
  NANDN U8772 ( .A(n7648), .B(n7647), .Z(n7649) );
  AND U8773 ( .A(n7650), .B(n7649), .Z(n7749) );
  AND U8774 ( .A(x[233]), .B(y[1870]), .Z(n8544) );
  NANDN U8775 ( .A(n7737), .B(n8544), .Z(n7654) );
  NANDN U8776 ( .A(n7652), .B(n7651), .Z(n7653) );
  NAND U8777 ( .A(n7654), .B(n7653), .Z(n7748) );
  XNOR U8778 ( .A(n7749), .B(n7748), .Z(n7750) );
  AND U8779 ( .A(x[229]), .B(y[1868]), .Z(n7785) );
  NAND U8780 ( .A(y[1865]), .B(x[232]), .Z(n7655) );
  XNOR U8781 ( .A(n7785), .B(n7655), .Z(n7730) );
  XOR U8782 ( .A(n7730), .B(n7729), .Z(n7742) );
  XOR U8783 ( .A(n7742), .B(n7743), .Z(n7744) );
  NAND U8784 ( .A(y[1869]), .B(x[228]), .Z(n7656) );
  XNOR U8785 ( .A(n7657), .B(n7656), .Z(n7691) );
  NAND U8786 ( .A(x[235]), .B(y[1862]), .Z(n7692) );
  XOR U8787 ( .A(n7691), .B(n7692), .Z(n7745) );
  XOR U8788 ( .A(n7744), .B(n7745), .Z(n7751) );
  XNOR U8789 ( .A(n7750), .B(n7751), .Z(n7754) );
  XOR U8790 ( .A(n7755), .B(n7754), .Z(n7756) );
  XNOR U8791 ( .A(n7757), .B(n7756), .Z(n7675) );
  NAND U8792 ( .A(n7659), .B(n7658), .Z(n7663) );
  NAND U8793 ( .A(n7661), .B(n7660), .Z(n7662) );
  NAND U8794 ( .A(n7663), .B(n7662), .Z(n7674) );
  XOR U8795 ( .A(n7675), .B(n7674), .Z(n7676) );
  XOR U8796 ( .A(n7677), .B(n7676), .Z(n7665) );
  XOR U8797 ( .A(n7667), .B(n7668), .Z(n7673) );
  XNOR U8798 ( .A(n7672), .B(n7673), .Z(n7664) );
  XOR U8799 ( .A(n7671), .B(n7664), .Z(N178) );
  NANDN U8800 ( .A(n7666), .B(n7665), .Z(n7670) );
  NAND U8801 ( .A(n7668), .B(n7667), .Z(n7669) );
  AND U8802 ( .A(n7670), .B(n7669), .Z(n7875) );
  NAND U8803 ( .A(n7675), .B(n7674), .Z(n7679) );
  NANDN U8804 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U8805 ( .A(n7679), .B(n7678), .Z(n7872) );
  NAND U8806 ( .A(n7681), .B(n7680), .Z(n7685) );
  NAND U8807 ( .A(n7683), .B(n7682), .Z(n7684) );
  AND U8808 ( .A(n7685), .B(n7684), .Z(n7870) );
  AND U8809 ( .A(x[236]), .B(y[1858]), .Z(n8003) );
  AND U8810 ( .A(x[239]), .B(y[1861]), .Z(n7937) );
  NAND U8811 ( .A(n8003), .B(n7937), .Z(n7689) );
  NANDN U8812 ( .A(n7687), .B(n7686), .Z(n7688) );
  NAND U8813 ( .A(n7689), .B(n7688), .Z(n7852) );
  NAND U8814 ( .A(n8944), .B(n7690), .Z(n7694) );
  NANDN U8815 ( .A(n7692), .B(n7691), .Z(n7693) );
  AND U8816 ( .A(n7694), .B(n7693), .Z(n7842) );
  AND U8817 ( .A(y[1873]), .B(x[225]), .Z(n7696) );
  NAND U8818 ( .A(y[1864]), .B(x[234]), .Z(n7695) );
  XNOR U8819 ( .A(n7696), .B(n7695), .Z(n7804) );
  NANDN U8820 ( .A(n7697), .B(o[81]), .Z(n7805) );
  XNOR U8821 ( .A(n7804), .B(n7805), .Z(n7839) );
  AND U8822 ( .A(y[1859]), .B(x[239]), .Z(n7699) );
  NAND U8823 ( .A(y[1865]), .B(x[233]), .Z(n7698) );
  XNOR U8824 ( .A(n7699), .B(n7698), .Z(n7795) );
  NAND U8825 ( .A(x[238]), .B(y[1860]), .Z(n7796) );
  XOR U8826 ( .A(n7795), .B(n7796), .Z(n7840) );
  XNOR U8827 ( .A(n7839), .B(n7840), .Z(n7841) );
  XNOR U8828 ( .A(n7842), .B(n7841), .Z(n7851) );
  XOR U8829 ( .A(n7852), .B(n7851), .Z(n7854) );
  NANDN U8830 ( .A(n7701), .B(n7700), .Z(n7705) );
  NANDN U8831 ( .A(n7703), .B(n7702), .Z(n7704) );
  AND U8832 ( .A(n7705), .B(n7704), .Z(n7864) );
  AND U8833 ( .A(y[1858]), .B(x[240]), .Z(n7707) );
  NAND U8834 ( .A(y[1863]), .B(x[235]), .Z(n7706) );
  XNOR U8835 ( .A(n7707), .B(n7706), .Z(n7791) );
  NAND U8836 ( .A(x[226]), .B(y[1872]), .Z(n7792) );
  XNOR U8837 ( .A(n7791), .B(n7792), .Z(n7863) );
  AND U8838 ( .A(x[229]), .B(y[1869]), .Z(n7885) );
  NAND U8839 ( .A(y[1868]), .B(x[230]), .Z(n7708) );
  XNOR U8840 ( .A(n7885), .B(n7708), .Z(n7787) );
  NAND U8841 ( .A(y[1870]), .B(x[228]), .Z(n7709) );
  XNOR U8842 ( .A(n8549), .B(n7709), .Z(n7826) );
  NAND U8843 ( .A(x[231]), .B(y[1867]), .Z(n7827) );
  XNOR U8844 ( .A(n7787), .B(n7788), .Z(n7865) );
  XOR U8845 ( .A(n7866), .B(n7865), .Z(n7853) );
  XNOR U8846 ( .A(n7854), .B(n7853), .Z(n7774) );
  NAND U8847 ( .A(n7711), .B(n7710), .Z(n7715) );
  NAND U8848 ( .A(n7713), .B(n7712), .Z(n7714) );
  AND U8849 ( .A(n7715), .B(n7714), .Z(n7845) );
  NAND U8850 ( .A(n7717), .B(n7716), .Z(n7721) );
  NAND U8851 ( .A(n7719), .B(n7718), .Z(n7720) );
  AND U8852 ( .A(n7721), .B(n7720), .Z(n7846) );
  XOR U8853 ( .A(n7845), .B(n7846), .Z(n7847) );
  NAND U8854 ( .A(n7723), .B(n7722), .Z(n7727) );
  NAND U8855 ( .A(n7725), .B(n7724), .Z(n7726) );
  AND U8856 ( .A(n7727), .B(n7726), .Z(n7848) );
  XOR U8857 ( .A(n7847), .B(n7848), .Z(n7773) );
  XOR U8858 ( .A(n7774), .B(n7773), .Z(n7776) );
  AND U8859 ( .A(x[232]), .B(y[1868]), .Z(n8049) );
  NAND U8860 ( .A(n8049), .B(n7728), .Z(n7732) );
  NAND U8861 ( .A(n7730), .B(n7729), .Z(n7731) );
  NAND U8862 ( .A(n7732), .B(n7731), .Z(n7858) );
  NAND U8863 ( .A(x[233]), .B(y[1872]), .Z(n8696) );
  NANDN U8864 ( .A(n8696), .B(n7803), .Z(n7736) );
  NANDN U8865 ( .A(n7734), .B(n7733), .Z(n7735) );
  NAND U8866 ( .A(n7736), .B(n7735), .Z(n7857) );
  XOR U8867 ( .A(n7858), .B(n7857), .Z(n7860) );
  NAND U8868 ( .A(x[234]), .B(y[1871]), .Z(n8695) );
  AND U8869 ( .A(x[224]), .B(y[1874]), .Z(n7808) );
  NAND U8870 ( .A(x[242]), .B(y[1856]), .Z(n7809) );
  XNOR U8871 ( .A(n7808), .B(n7809), .Z(n7810) );
  NAND U8872 ( .A(x[241]), .B(y[1857]), .Z(n7830) );
  XOR U8873 ( .A(o[82]), .B(n7830), .Z(n7811) );
  XNOR U8874 ( .A(n7810), .B(n7811), .Z(n7833) );
  AND U8875 ( .A(y[1861]), .B(x[237]), .Z(n7741) );
  NAND U8876 ( .A(y[1871]), .B(x[227]), .Z(n7740) );
  XNOR U8877 ( .A(n7741), .B(n7740), .Z(n7816) );
  NAND U8878 ( .A(x[236]), .B(y[1862]), .Z(n7817) );
  XOR U8879 ( .A(n7816), .B(n7817), .Z(n7834) );
  XNOR U8880 ( .A(n7833), .B(n7834), .Z(n7835) );
  XNOR U8881 ( .A(n7836), .B(n7835), .Z(n7859) );
  XOR U8882 ( .A(n7860), .B(n7859), .Z(n7780) );
  NAND U8883 ( .A(n7743), .B(n7742), .Z(n7747) );
  NANDN U8884 ( .A(n7745), .B(n7744), .Z(n7746) );
  AND U8885 ( .A(n7747), .B(n7746), .Z(n7779) );
  XNOR U8886 ( .A(n7780), .B(n7779), .Z(n7781) );
  NANDN U8887 ( .A(n7749), .B(n7748), .Z(n7753) );
  NANDN U8888 ( .A(n7751), .B(n7750), .Z(n7752) );
  NAND U8889 ( .A(n7753), .B(n7752), .Z(n7782) );
  XNOR U8890 ( .A(n7781), .B(n7782), .Z(n7775) );
  XNOR U8891 ( .A(n7776), .B(n7775), .Z(n7770) );
  NAND U8892 ( .A(n7755), .B(n7754), .Z(n7759) );
  NAND U8893 ( .A(n7757), .B(n7756), .Z(n7758) );
  NAND U8894 ( .A(n7759), .B(n7758), .Z(n7768) );
  NAND U8895 ( .A(n7761), .B(n7760), .Z(n7765) );
  NAND U8896 ( .A(n7763), .B(n7762), .Z(n7764) );
  NAND U8897 ( .A(n7765), .B(n7764), .Z(n7767) );
  XOR U8898 ( .A(n7768), .B(n7767), .Z(n7769) );
  XOR U8899 ( .A(n7770), .B(n7769), .Z(n7869) );
  XOR U8900 ( .A(n7870), .B(n7869), .Z(n7871) );
  XOR U8901 ( .A(n7872), .B(n7871), .Z(n7877) );
  XNOR U8902 ( .A(n7876), .B(n7877), .Z(n7766) );
  XOR U8903 ( .A(n7875), .B(n7766), .Z(N179) );
  NAND U8904 ( .A(n7768), .B(n7767), .Z(n7772) );
  NAND U8905 ( .A(n7770), .B(n7769), .Z(n7771) );
  AND U8906 ( .A(n7772), .B(n7771), .Z(n7993) );
  NAND U8907 ( .A(n7774), .B(n7773), .Z(n7778) );
  NAND U8908 ( .A(n7776), .B(n7775), .Z(n7777) );
  AND U8909 ( .A(n7778), .B(n7777), .Z(n7991) );
  NANDN U8910 ( .A(n7780), .B(n7779), .Z(n7784) );
  NANDN U8911 ( .A(n7782), .B(n7781), .Z(n7783) );
  AND U8912 ( .A(n7784), .B(n7783), .Z(n7881) );
  AND U8913 ( .A(x[230]), .B(y[1869]), .Z(n7786) );
  NAND U8914 ( .A(n7786), .B(n7785), .Z(n7790) );
  NANDN U8915 ( .A(n7788), .B(n7787), .Z(n7789) );
  AND U8916 ( .A(n7790), .B(n7789), .Z(n7971) );
  AND U8917 ( .A(x[240]), .B(y[1863]), .Z(n8336) );
  NAND U8918 ( .A(n8336), .B(n8154), .Z(n7794) );
  NANDN U8919 ( .A(n7792), .B(n7791), .Z(n7793) );
  AND U8920 ( .A(n7794), .B(n7793), .Z(n7970) );
  AND U8921 ( .A(x[239]), .B(y[1865]), .Z(n8580) );
  NAND U8922 ( .A(n8580), .B(n7924), .Z(n7798) );
  NANDN U8923 ( .A(n7796), .B(n7795), .Z(n7797) );
  AND U8924 ( .A(n7798), .B(n7797), .Z(n7954) );
  AND U8925 ( .A(y[1874]), .B(x[225]), .Z(n7800) );
  NAND U8926 ( .A(y[1867]), .B(x[232]), .Z(n7799) );
  XNOR U8927 ( .A(n7800), .B(n7799), .Z(n7903) );
  AND U8928 ( .A(y[1862]), .B(x[237]), .Z(n7802) );
  NAND U8929 ( .A(y[1873]), .B(x[226]), .Z(n7801) );
  XNOR U8930 ( .A(n7802), .B(n7801), .Z(n7930) );
  XOR U8931 ( .A(n7952), .B(n7951), .Z(n7953) );
  XOR U8932 ( .A(n7970), .B(n7969), .Z(n7972) );
  XOR U8933 ( .A(n7971), .B(n7972), .Z(n7880) );
  NAND U8934 ( .A(x[234]), .B(y[1873]), .Z(n9026) );
  NANDN U8935 ( .A(n9026), .B(n7803), .Z(n7807) );
  NANDN U8936 ( .A(n7805), .B(n7804), .Z(n7806) );
  AND U8937 ( .A(n7807), .B(n7806), .Z(n7915) );
  NANDN U8938 ( .A(n7809), .B(n7808), .Z(n7813) );
  NANDN U8939 ( .A(n7811), .B(n7810), .Z(n7812) );
  AND U8940 ( .A(n7813), .B(n7812), .Z(n7913) );
  AND U8941 ( .A(y[1859]), .B(x[240]), .Z(n8627) );
  NAND U8942 ( .A(y[1866]), .B(x[233]), .Z(n7814) );
  XNOR U8943 ( .A(n8627), .B(n7814), .Z(n7925) );
  NAND U8944 ( .A(x[239]), .B(y[1860]), .Z(n7926) );
  AND U8945 ( .A(x[237]), .B(y[1871]), .Z(n9234) );
  NANDN U8946 ( .A(n7815), .B(n9234), .Z(n7819) );
  NANDN U8947 ( .A(n7817), .B(n7816), .Z(n7818) );
  AND U8948 ( .A(n7819), .B(n7818), .Z(n7921) );
  AND U8949 ( .A(y[1865]), .B(x[234]), .Z(n7821) );
  NAND U8950 ( .A(y[1858]), .B(x[241]), .Z(n7820) );
  XNOR U8951 ( .A(n7821), .B(n7820), .Z(n7909) );
  AND U8952 ( .A(x[242]), .B(y[1857]), .Z(n7944) );
  XOR U8953 ( .A(o[83]), .B(n7944), .Z(n7908) );
  XOR U8954 ( .A(n7909), .B(n7908), .Z(n7919) );
  NAND U8955 ( .A(y[1872]), .B(x[227]), .Z(n7822) );
  XNOR U8956 ( .A(n7823), .B(n7822), .Z(n7938) );
  XOR U8957 ( .A(n7919), .B(n7918), .Z(n7920) );
  NAND U8958 ( .A(n7825), .B(n7824), .Z(n7829) );
  NANDN U8959 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U8960 ( .A(n7829), .B(n7828), .Z(n7948) );
  AND U8961 ( .A(x[224]), .B(y[1875]), .Z(n7889) );
  NAND U8962 ( .A(x[243]), .B(y[1856]), .Z(n7890) );
  ANDN U8963 ( .B(o[82]), .A(n7830), .Z(n7891) );
  XOR U8964 ( .A(n7892), .B(n7891), .Z(n7946) );
  AND U8965 ( .A(x[228]), .B(y[1871]), .Z(n8063) );
  AND U8966 ( .A(y[1870]), .B(x[229]), .Z(n7832) );
  NAND U8967 ( .A(y[1869]), .B(x[230]), .Z(n7831) );
  XOR U8968 ( .A(n7832), .B(n7831), .Z(n7886) );
  XOR U8969 ( .A(n7946), .B(n7945), .Z(n7947) );
  XOR U8970 ( .A(n7948), .B(n7947), .Z(n7963) );
  XNOR U8971 ( .A(n7964), .B(n7963), .Z(n7966) );
  XOR U8972 ( .A(n7965), .B(n7966), .Z(n7959) );
  NANDN U8973 ( .A(n7834), .B(n7833), .Z(n7838) );
  NANDN U8974 ( .A(n7836), .B(n7835), .Z(n7837) );
  AND U8975 ( .A(n7838), .B(n7837), .Z(n7958) );
  NANDN U8976 ( .A(n7840), .B(n7839), .Z(n7844) );
  NANDN U8977 ( .A(n7842), .B(n7841), .Z(n7843) );
  NAND U8978 ( .A(n7844), .B(n7843), .Z(n7957) );
  XOR U8979 ( .A(n7958), .B(n7957), .Z(n7960) );
  XOR U8980 ( .A(n7959), .B(n7960), .Z(n7879) );
  XOR U8981 ( .A(n7880), .B(n7879), .Z(n7882) );
  XNOR U8982 ( .A(n7881), .B(n7882), .Z(n7984) );
  NAND U8983 ( .A(n7846), .B(n7845), .Z(n7850) );
  NAND U8984 ( .A(n7848), .B(n7847), .Z(n7849) );
  AND U8985 ( .A(n7850), .B(n7849), .Z(n7982) );
  NAND U8986 ( .A(n7852), .B(n7851), .Z(n7856) );
  NAND U8987 ( .A(n7854), .B(n7853), .Z(n7855) );
  AND U8988 ( .A(n7856), .B(n7855), .Z(n7978) );
  NAND U8989 ( .A(n7858), .B(n7857), .Z(n7862) );
  NAND U8990 ( .A(n7860), .B(n7859), .Z(n7861) );
  AND U8991 ( .A(n7862), .B(n7861), .Z(n7976) );
  NANDN U8992 ( .A(n7864), .B(n7863), .Z(n7868) );
  NAND U8993 ( .A(n7866), .B(n7865), .Z(n7867) );
  NAND U8994 ( .A(n7868), .B(n7867), .Z(n7975) );
  XOR U8995 ( .A(n7982), .B(n7981), .Z(n7983) );
  XOR U8996 ( .A(n7984), .B(n7983), .Z(n7990) );
  XOR U8997 ( .A(n7991), .B(n7990), .Z(n7992) );
  XOR U8998 ( .A(n7993), .B(n7992), .Z(n7989) );
  NAND U8999 ( .A(n7870), .B(n7869), .Z(n7874) );
  NAND U9000 ( .A(n7872), .B(n7871), .Z(n7873) );
  NAND U9001 ( .A(n7874), .B(n7873), .Z(n7988) );
  XOR U9002 ( .A(n7988), .B(n7987), .Z(n7878) );
  XNOR U9003 ( .A(n7989), .B(n7878), .Z(N180) );
  NANDN U9004 ( .A(n7880), .B(n7879), .Z(n7884) );
  OR U9005 ( .A(n7882), .B(n7881), .Z(n7883) );
  AND U9006 ( .A(n7884), .B(n7883), .Z(n8101) );
  AND U9007 ( .A(x[230]), .B(y[1870]), .Z(n8020) );
  IV U9008 ( .A(n8020), .Z(n7901) );
  NANDN U9009 ( .A(n7901), .B(n7885), .Z(n7888) );
  NANDN U9010 ( .A(n7886), .B(n8063), .Z(n7887) );
  AND U9011 ( .A(n7888), .B(n7887), .Z(n8028) );
  NANDN U9012 ( .A(n7890), .B(n7889), .Z(n7894) );
  NAND U9013 ( .A(n7892), .B(n7891), .Z(n7893) );
  AND U9014 ( .A(n7894), .B(n7893), .Z(n8026) );
  AND U9015 ( .A(y[1858]), .B(x[242]), .Z(n7896) );
  NAND U9016 ( .A(y[1864]), .B(x[236]), .Z(n7895) );
  XNOR U9017 ( .A(n7896), .B(n7895), .Z(n8004) );
  AND U9018 ( .A(x[241]), .B(y[1859]), .Z(n8005) );
  XOR U9019 ( .A(n8004), .B(n8005), .Z(n8025) );
  AND U9020 ( .A(y[1863]), .B(x[237]), .Z(n7898) );
  NAND U9021 ( .A(y[1873]), .B(x[227]), .Z(n7897) );
  XNOR U9022 ( .A(n7898), .B(n7897), .Z(n8050) );
  XOR U9023 ( .A(n8050), .B(n8049), .Z(n8022) );
  AND U9024 ( .A(y[1871]), .B(x[229]), .Z(n7900) );
  NAND U9025 ( .A(y[1872]), .B(x[228]), .Z(n7899) );
  XNOR U9026 ( .A(n7900), .B(n7899), .Z(n8065) );
  AND U9027 ( .A(x[231]), .B(y[1869]), .Z(n8064) );
  XNOR U9028 ( .A(n8065), .B(n8064), .Z(n8019) );
  XOR U9029 ( .A(n7901), .B(n8019), .Z(n8021) );
  AND U9030 ( .A(x[232]), .B(y[1874]), .Z(n9190) );
  AND U9031 ( .A(x[225]), .B(y[1867]), .Z(n7902) );
  NAND U9032 ( .A(n9190), .B(n7902), .Z(n7906) );
  NANDN U9033 ( .A(n7904), .B(n7903), .Z(n7905) );
  AND U9034 ( .A(n7906), .B(n7905), .Z(n8075) );
  NAND U9035 ( .A(x[241]), .B(y[1865]), .Z(n8879) );
  NANDN U9036 ( .A(n8879), .B(n7907), .Z(n7911) );
  NAND U9037 ( .A(n7909), .B(n7908), .Z(n7910) );
  NAND U9038 ( .A(n7911), .B(n7910), .Z(n8074) );
  XNOR U9039 ( .A(n8076), .B(n8077), .Z(n8031) );
  XOR U9040 ( .A(n8032), .B(n8031), .Z(n8033) );
  NANDN U9041 ( .A(n7913), .B(n7912), .Z(n7917) );
  NANDN U9042 ( .A(n7915), .B(n7914), .Z(n7916) );
  NAND U9043 ( .A(n7917), .B(n7916), .Z(n8034) );
  NAND U9044 ( .A(n7919), .B(n7918), .Z(n7923) );
  NANDN U9045 ( .A(n7921), .B(n7920), .Z(n7922) );
  NAND U9046 ( .A(n7923), .B(n7922), .Z(n8093) );
  AND U9047 ( .A(x[240]), .B(y[1866]), .Z(n8871) );
  NAND U9048 ( .A(n8871), .B(n7924), .Z(n7928) );
  NANDN U9049 ( .A(n7926), .B(n7925), .Z(n7927) );
  AND U9050 ( .A(n7928), .B(n7927), .Z(n8038) );
  AND U9051 ( .A(x[237]), .B(y[1873]), .Z(n9458) );
  NAND U9052 ( .A(n9458), .B(n7929), .Z(n7933) );
  NANDN U9053 ( .A(n7931), .B(n7930), .Z(n7932) );
  AND U9054 ( .A(n7933), .B(n7932), .Z(n8083) );
  AND U9055 ( .A(y[1860]), .B(x[240]), .Z(n7935) );
  NAND U9056 ( .A(y[1866]), .B(x[234]), .Z(n7934) );
  XNOR U9057 ( .A(n7935), .B(n7934), .Z(n8044) );
  AND U9058 ( .A(x[226]), .B(y[1874]), .Z(n8045) );
  XOR U9059 ( .A(n8044), .B(n8045), .Z(n8081) );
  NAND U9060 ( .A(y[1867]), .B(x[233]), .Z(n7936) );
  XNOR U9061 ( .A(n7937), .B(n7936), .Z(n8014) );
  AND U9062 ( .A(x[238]), .B(y[1862]), .Z(n8015) );
  XOR U9063 ( .A(n8014), .B(n8015), .Z(n8080) );
  XOR U9064 ( .A(n8081), .B(n8080), .Z(n8082) );
  NAND U9065 ( .A(x[235]), .B(y[1872]), .Z(n9027) );
  NANDN U9066 ( .A(n9027), .B(n8181), .Z(n7941) );
  NANDN U9067 ( .A(n7939), .B(n7938), .Z(n7940) );
  AND U9068 ( .A(n7941), .B(n7940), .Z(n8089) );
  AND U9069 ( .A(y[1865]), .B(x[235]), .Z(n7943) );
  NAND U9070 ( .A(y[1875]), .B(x[225]), .Z(n7942) );
  XNOR U9071 ( .A(n7943), .B(n7942), .Z(n8010) );
  AND U9072 ( .A(x[243]), .B(y[1857]), .Z(n8018) );
  XOR U9073 ( .A(o[84]), .B(n8018), .Z(n8009) );
  XOR U9074 ( .A(n8010), .B(n8009), .Z(n8087) );
  AND U9075 ( .A(o[83]), .B(n7944), .Z(n8071) );
  AND U9076 ( .A(x[224]), .B(y[1876]), .Z(n8068) );
  AND U9077 ( .A(x[244]), .B(y[1856]), .Z(n8069) );
  XOR U9078 ( .A(n8068), .B(n8069), .Z(n8070) );
  XOR U9079 ( .A(n8071), .B(n8070), .Z(n8086) );
  XOR U9080 ( .A(n8087), .B(n8086), .Z(n8088) );
  XOR U9081 ( .A(n8040), .B(n8039), .Z(n8000) );
  NAND U9082 ( .A(n7946), .B(n7945), .Z(n7950) );
  NANDN U9083 ( .A(n7948), .B(n7947), .Z(n7949) );
  AND U9084 ( .A(n7950), .B(n7949), .Z(n7997) );
  NAND U9085 ( .A(n7952), .B(n7951), .Z(n7956) );
  NANDN U9086 ( .A(n7954), .B(n7953), .Z(n7955) );
  NAND U9087 ( .A(n7956), .B(n7955), .Z(n7998) );
  XOR U9088 ( .A(n8095), .B(n8094), .Z(n8099) );
  NANDN U9089 ( .A(n7958), .B(n7957), .Z(n7962) );
  NANDN U9090 ( .A(n7960), .B(n7959), .Z(n7961) );
  AND U9091 ( .A(n7962), .B(n7961), .Z(n8107) );
  NAND U9092 ( .A(n7964), .B(n7963), .Z(n7968) );
  NANDN U9093 ( .A(n7966), .B(n7965), .Z(n7967) );
  AND U9094 ( .A(n7968), .B(n7967), .Z(n8105) );
  NANDN U9095 ( .A(n7970), .B(n7969), .Z(n7974) );
  OR U9096 ( .A(n7972), .B(n7971), .Z(n7973) );
  AND U9097 ( .A(n7974), .B(n7973), .Z(n8104) );
  XNOR U9098 ( .A(n8105), .B(n8104), .Z(n8106) );
  XNOR U9099 ( .A(n8107), .B(n8106), .Z(n8098) );
  XNOR U9100 ( .A(n8099), .B(n8098), .Z(n8100) );
  XOR U9101 ( .A(n8101), .B(n8100), .Z(n8120) );
  NANDN U9102 ( .A(n7976), .B(n7975), .Z(n7980) );
  NANDN U9103 ( .A(n7978), .B(n7977), .Z(n7979) );
  AND U9104 ( .A(n7980), .B(n7979), .Z(n8117) );
  NAND U9105 ( .A(n7982), .B(n7981), .Z(n7986) );
  NAND U9106 ( .A(n7984), .B(n7983), .Z(n7985) );
  AND U9107 ( .A(n7986), .B(n7985), .Z(n8118) );
  XOR U9108 ( .A(n8117), .B(n8118), .Z(n8119) );
  XOR U9109 ( .A(n8120), .B(n8119), .Z(n8113) );
  NAND U9110 ( .A(n7991), .B(n7990), .Z(n7995) );
  NANDN U9111 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U9112 ( .A(n7995), .B(n7994), .Z(n8112) );
  IV U9113 ( .A(n8112), .Z(n8110) );
  XOR U9114 ( .A(n8111), .B(n8110), .Z(n7996) );
  XNOR U9115 ( .A(n8113), .B(n7996), .Z(N181) );
  NANDN U9116 ( .A(n7998), .B(n7997), .Z(n8002) );
  NANDN U9117 ( .A(n8000), .B(n7999), .Z(n8001) );
  AND U9118 ( .A(n8002), .B(n8001), .Z(n8133) );
  AND U9119 ( .A(x[242]), .B(y[1864]), .Z(n8878) );
  NAND U9120 ( .A(n8878), .B(n8003), .Z(n8007) );
  NAND U9121 ( .A(n8005), .B(n8004), .Z(n8006) );
  NAND U9122 ( .A(n8007), .B(n8006), .Z(n8204) );
  AND U9123 ( .A(x[235]), .B(y[1875]), .Z(n9644) );
  AND U9124 ( .A(x[225]), .B(y[1865]), .Z(n8008) );
  NAND U9125 ( .A(n9644), .B(n8008), .Z(n8012) );
  NAND U9126 ( .A(n8010), .B(n8009), .Z(n8011) );
  NAND U9127 ( .A(n8012), .B(n8011), .Z(n8203) );
  XOR U9128 ( .A(n8204), .B(n8203), .Z(n8206) );
  AND U9129 ( .A(x[239]), .B(y[1867]), .Z(n8866) );
  NAND U9130 ( .A(n8866), .B(n8013), .Z(n8017) );
  NAND U9131 ( .A(n8015), .B(n8014), .Z(n8016) );
  NAND U9132 ( .A(n8017), .B(n8016), .Z(n8168) );
  AND U9133 ( .A(o[84]), .B(n8018), .Z(n8190) );
  AND U9134 ( .A(x[224]), .B(y[1877]), .Z(n8187) );
  AND U9135 ( .A(x[245]), .B(y[1856]), .Z(n8188) );
  XOR U9136 ( .A(n8187), .B(n8188), .Z(n8189) );
  XOR U9137 ( .A(n8190), .B(n8189), .Z(n8166) );
  AND U9138 ( .A(x[229]), .B(y[1872]), .Z(n8174) );
  AND U9139 ( .A(x[240]), .B(y[1861]), .Z(n8173) );
  XOR U9140 ( .A(n8174), .B(n8173), .Z(n8172) );
  AND U9141 ( .A(x[239]), .B(y[1862]), .Z(n8171) );
  XOR U9142 ( .A(n8172), .B(n8171), .Z(n8165) );
  XOR U9143 ( .A(n8166), .B(n8165), .Z(n8167) );
  XOR U9144 ( .A(n8168), .B(n8167), .Z(n8205) );
  XOR U9145 ( .A(n8206), .B(n8205), .Z(n8222) );
  NANDN U9146 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U9147 ( .A(n8022), .B(n8021), .Z(n8023) );
  NAND U9148 ( .A(n8024), .B(n8023), .Z(n8221) );
  NANDN U9149 ( .A(n8026), .B(n8025), .Z(n8030) );
  NANDN U9150 ( .A(n8028), .B(n8027), .Z(n8029) );
  AND U9151 ( .A(n8030), .B(n8029), .Z(n8223) );
  XOR U9152 ( .A(n8224), .B(n8223), .Z(n8131) );
  NAND U9153 ( .A(n8032), .B(n8031), .Z(n8036) );
  NANDN U9154 ( .A(n8034), .B(n8033), .Z(n8035) );
  AND U9155 ( .A(n8036), .B(n8035), .Z(n8130) );
  XOR U9156 ( .A(n8133), .B(n8132), .Z(n8127) );
  NANDN U9157 ( .A(n8038), .B(n8037), .Z(n8042) );
  NAND U9158 ( .A(n8040), .B(n8039), .Z(n8041) );
  AND U9159 ( .A(n8042), .B(n8041), .Z(n8230) );
  AND U9160 ( .A(x[234]), .B(y[1860]), .Z(n8043) );
  NAND U9161 ( .A(n8871), .B(n8043), .Z(n8047) );
  NAND U9162 ( .A(n8045), .B(n8044), .Z(n8046) );
  NAND U9163 ( .A(n8047), .B(n8046), .Z(n8137) );
  NAND U9164 ( .A(n9458), .B(n8048), .Z(n8052) );
  NAND U9165 ( .A(n8050), .B(n8049), .Z(n8051) );
  NAND U9166 ( .A(n8052), .B(n8051), .Z(n8218) );
  AND U9167 ( .A(y[1858]), .B(x[243]), .Z(n8054) );
  NAND U9168 ( .A(y[1866]), .B(x[235]), .Z(n8053) );
  XNOR U9169 ( .A(n8054), .B(n8053), .Z(n8156) );
  AND U9170 ( .A(x[244]), .B(y[1857]), .Z(n8186) );
  XOR U9171 ( .A(o[85]), .B(n8186), .Z(n8155) );
  XOR U9172 ( .A(n8156), .B(n8155), .Z(n8216) );
  AND U9173 ( .A(y[1859]), .B(x[242]), .Z(n8056) );
  NAND U9174 ( .A(y[1867]), .B(x[234]), .Z(n8055) );
  XNOR U9175 ( .A(n8056), .B(n8055), .Z(n8194) );
  AND U9176 ( .A(x[225]), .B(y[1876]), .Z(n8195) );
  XOR U9177 ( .A(n8194), .B(n8195), .Z(n8215) );
  XOR U9178 ( .A(n8216), .B(n8215), .Z(n8217) );
  XOR U9179 ( .A(n8218), .B(n8217), .Z(n8136) );
  XOR U9180 ( .A(n8137), .B(n8136), .Z(n8139) );
  AND U9181 ( .A(x[231]), .B(y[1870]), .Z(n8399) );
  AND U9182 ( .A(y[1871]), .B(x[230]), .Z(n8058) );
  NAND U9183 ( .A(y[1863]), .B(x[238]), .Z(n8057) );
  XNOR U9184 ( .A(n8058), .B(n8057), .Z(n8198) );
  XNOR U9185 ( .A(n8399), .B(n8198), .Z(n8145) );
  NAND U9186 ( .A(x[233]), .B(y[1868]), .Z(n8143) );
  NAND U9187 ( .A(x[232]), .B(y[1869]), .Z(n8142) );
  XOR U9188 ( .A(n8143), .B(n8142), .Z(n8144) );
  XNOR U9189 ( .A(n8145), .B(n8144), .Z(n8161) );
  AND U9190 ( .A(y[1865]), .B(x[236]), .Z(n8060) );
  NAND U9191 ( .A(y[1860]), .B(x[241]), .Z(n8059) );
  XNOR U9192 ( .A(n8060), .B(n8059), .Z(n8148) );
  AND U9193 ( .A(x[226]), .B(y[1875]), .Z(n8149) );
  XOR U9194 ( .A(n8148), .B(n8149), .Z(n8160) );
  AND U9195 ( .A(y[1864]), .B(x[237]), .Z(n8062) );
  NAND U9196 ( .A(y[1874]), .B(x[227]), .Z(n8061) );
  XNOR U9197 ( .A(n8062), .B(n8061), .Z(n8182) );
  AND U9198 ( .A(x[228]), .B(y[1873]), .Z(n8183) );
  XOR U9199 ( .A(n8182), .B(n8183), .Z(n8159) );
  XOR U9200 ( .A(n8160), .B(n8159), .Z(n8162) );
  XOR U9201 ( .A(n8161), .B(n8162), .Z(n8212) );
  NAND U9202 ( .A(n8174), .B(n8063), .Z(n8067) );
  NAND U9203 ( .A(n8065), .B(n8064), .Z(n8066) );
  NAND U9204 ( .A(n8067), .B(n8066), .Z(n8210) );
  NAND U9205 ( .A(n8069), .B(n8068), .Z(n8073) );
  NAND U9206 ( .A(n8071), .B(n8070), .Z(n8072) );
  NAND U9207 ( .A(n8073), .B(n8072), .Z(n8209) );
  XOR U9208 ( .A(n8210), .B(n8209), .Z(n8211) );
  XOR U9209 ( .A(n8212), .B(n8211), .Z(n8138) );
  XOR U9210 ( .A(n8139), .B(n8138), .Z(n8228) );
  NANDN U9211 ( .A(n8075), .B(n8074), .Z(n8079) );
  NAND U9212 ( .A(n8077), .B(n8076), .Z(n8078) );
  NAND U9213 ( .A(n8079), .B(n8078), .Z(n8235) );
  NAND U9214 ( .A(n8081), .B(n8080), .Z(n8085) );
  NANDN U9215 ( .A(n8083), .B(n8082), .Z(n8084) );
  NAND U9216 ( .A(n8085), .B(n8084), .Z(n8234) );
  NAND U9217 ( .A(n8087), .B(n8086), .Z(n8091) );
  NANDN U9218 ( .A(n8089), .B(n8088), .Z(n8090) );
  NAND U9219 ( .A(n8091), .B(n8090), .Z(n8233) );
  XOR U9220 ( .A(n8234), .B(n8233), .Z(n8236) );
  XOR U9221 ( .A(n8235), .B(n8236), .Z(n8227) );
  XOR U9222 ( .A(n8228), .B(n8227), .Z(n8229) );
  NANDN U9223 ( .A(n8093), .B(n8092), .Z(n8097) );
  NAND U9224 ( .A(n8095), .B(n8094), .Z(n8096) );
  NAND U9225 ( .A(n8097), .B(n8096), .Z(n8124) );
  XOR U9226 ( .A(n8125), .B(n8124), .Z(n8126) );
  NANDN U9227 ( .A(n8099), .B(n8098), .Z(n8103) );
  NAND U9228 ( .A(n8101), .B(n8100), .Z(n8102) );
  AND U9229 ( .A(n8103), .B(n8102), .Z(n8243) );
  NANDN U9230 ( .A(n8105), .B(n8104), .Z(n8109) );
  NAND U9231 ( .A(n8107), .B(n8106), .Z(n8108) );
  AND U9232 ( .A(n8109), .B(n8108), .Z(n8242) );
  XOR U9233 ( .A(n8243), .B(n8242), .Z(n8245) );
  XOR U9234 ( .A(n8244), .B(n8245), .Z(n8241) );
  NANDN U9235 ( .A(n8110), .B(n8111), .Z(n8116) );
  NOR U9236 ( .A(n8112), .B(n8111), .Z(n8114) );
  OR U9237 ( .A(n8114), .B(n8113), .Z(n8115) );
  AND U9238 ( .A(n8116), .B(n8115), .Z(n8239) );
  NAND U9239 ( .A(n8118), .B(n8117), .Z(n8122) );
  NANDN U9240 ( .A(n8120), .B(n8119), .Z(n8121) );
  AND U9241 ( .A(n8122), .B(n8121), .Z(n8240) );
  XOR U9242 ( .A(n8239), .B(n8240), .Z(n8123) );
  XNOR U9243 ( .A(n8241), .B(n8123), .Z(N182) );
  NAND U9244 ( .A(n8125), .B(n8124), .Z(n8129) );
  NANDN U9245 ( .A(n8127), .B(n8126), .Z(n8128) );
  AND U9246 ( .A(n8129), .B(n8128), .Z(n8252) );
  NANDN U9247 ( .A(n8131), .B(n8130), .Z(n8135) );
  NAND U9248 ( .A(n8133), .B(n8132), .Z(n8134) );
  AND U9249 ( .A(n8135), .B(n8134), .Z(n8250) );
  NAND U9250 ( .A(n8137), .B(n8136), .Z(n8141) );
  NAND U9251 ( .A(n8139), .B(n8138), .Z(n8140) );
  NAND U9252 ( .A(n8141), .B(n8140), .Z(n8375) );
  NAND U9253 ( .A(n8143), .B(n8142), .Z(n8147) );
  NAND U9254 ( .A(n8145), .B(n8144), .Z(n8146) );
  NAND U9255 ( .A(n8147), .B(n8146), .Z(n8369) );
  NANDN U9256 ( .A(n8879), .B(n8320), .Z(n8151) );
  NAND U9257 ( .A(n8149), .B(n8148), .Z(n8150) );
  NAND U9258 ( .A(n8151), .B(n8150), .Z(n8296) );
  AND U9259 ( .A(x[229]), .B(y[1873]), .Z(n8342) );
  AND U9260 ( .A(x[241]), .B(y[1861]), .Z(n8343) );
  XOR U9261 ( .A(n8342), .B(n8343), .Z(n8344) );
  AND U9262 ( .A(x[240]), .B(y[1862]), .Z(n8345) );
  XOR U9263 ( .A(n8344), .B(n8345), .Z(n8295) );
  AND U9264 ( .A(y[1860]), .B(x[242]), .Z(n8153) );
  NAND U9265 ( .A(y[1866]), .B(x[236]), .Z(n8152) );
  XNOR U9266 ( .A(n8153), .B(n8152), .Z(n8321) );
  AND U9267 ( .A(x[228]), .B(y[1874]), .Z(n8322) );
  XOR U9268 ( .A(n8321), .B(n8322), .Z(n8294) );
  XOR U9269 ( .A(n8295), .B(n8294), .Z(n8297) );
  XNOR U9270 ( .A(n8296), .B(n8297), .Z(n8366) );
  AND U9271 ( .A(x[243]), .B(y[1866]), .Z(n9360) );
  NAND U9272 ( .A(n9360), .B(n8154), .Z(n8158) );
  NAND U9273 ( .A(n8156), .B(n8155), .Z(n8157) );
  AND U9274 ( .A(n8158), .B(n8157), .Z(n8367) );
  XOR U9275 ( .A(n8366), .B(n8367), .Z(n8368) );
  XNOR U9276 ( .A(n8369), .B(n8368), .Z(n8372) );
  NAND U9277 ( .A(n8160), .B(n8159), .Z(n8164) );
  NAND U9278 ( .A(n8162), .B(n8161), .Z(n8163) );
  NAND U9279 ( .A(n8164), .B(n8163), .Z(n8355) );
  NAND U9280 ( .A(n8166), .B(n8165), .Z(n8170) );
  NAND U9281 ( .A(n8168), .B(n8167), .Z(n8169) );
  NAND U9282 ( .A(n8170), .B(n8169), .Z(n8354) );
  XOR U9283 ( .A(n8355), .B(n8354), .Z(n8357) );
  AND U9284 ( .A(n8172), .B(n8171), .Z(n8176) );
  NAND U9285 ( .A(n8174), .B(n8173), .Z(n8175) );
  NANDN U9286 ( .A(n8176), .B(n8175), .Z(n8317) );
  AND U9287 ( .A(y[1865]), .B(x[237]), .Z(n8178) );
  NAND U9288 ( .A(y[1858]), .B(x[244]), .Z(n8177) );
  XNOR U9289 ( .A(n8178), .B(n8177), .Z(n8338) );
  AND U9290 ( .A(x[226]), .B(y[1876]), .Z(n8339) );
  XOR U9291 ( .A(n8338), .B(n8339), .Z(n8315) );
  AND U9292 ( .A(y[1872]), .B(x[230]), .Z(n8180) );
  NAND U9293 ( .A(y[1863]), .B(x[239]), .Z(n8179) );
  XNOR U9294 ( .A(n8180), .B(n8179), .Z(n8350) );
  XOR U9295 ( .A(n8315), .B(n8314), .Z(n8316) );
  XOR U9296 ( .A(n8317), .B(n8316), .Z(n8361) );
  AND U9297 ( .A(x[237]), .B(y[1874]), .Z(n9645) );
  NAND U9298 ( .A(n8181), .B(n9645), .Z(n8185) );
  NAND U9299 ( .A(n8183), .B(n8182), .Z(n8184) );
  NAND U9300 ( .A(n8185), .B(n8184), .Z(n8285) );
  AND U9301 ( .A(x[225]), .B(y[1877]), .Z(n8308) );
  XOR U9302 ( .A(n8309), .B(n8308), .Z(n8307) );
  AND U9303 ( .A(o[85]), .B(n8186), .Z(n8306) );
  XOR U9304 ( .A(n8307), .B(n8306), .Z(n8283) );
  AND U9305 ( .A(x[238]), .B(y[1864]), .Z(n8300) );
  AND U9306 ( .A(x[227]), .B(y[1875]), .Z(n8301) );
  XOR U9307 ( .A(n8300), .B(n8301), .Z(n8302) );
  AND U9308 ( .A(x[243]), .B(y[1859]), .Z(n8303) );
  XOR U9309 ( .A(n8302), .B(n8303), .Z(n8282) );
  XOR U9310 ( .A(n8283), .B(n8282), .Z(n8284) );
  XOR U9311 ( .A(n8285), .B(n8284), .Z(n8360) );
  XOR U9312 ( .A(n8361), .B(n8360), .Z(n8363) );
  NAND U9313 ( .A(n8188), .B(n8187), .Z(n8192) );
  NAND U9314 ( .A(n8190), .B(n8189), .Z(n8191) );
  NAND U9315 ( .A(n8192), .B(n8191), .Z(n8277) );
  AND U9316 ( .A(x[242]), .B(y[1867]), .Z(n9363) );
  NAND U9317 ( .A(n9363), .B(n8193), .Z(n8197) );
  NAND U9318 ( .A(n8195), .B(n8194), .Z(n8196) );
  NAND U9319 ( .A(n8197), .B(n8196), .Z(n8276) );
  XOR U9320 ( .A(n8277), .B(n8276), .Z(n8279) );
  AND U9321 ( .A(x[238]), .B(y[1871]), .Z(n9373) );
  NAND U9322 ( .A(n9373), .B(n8349), .Z(n8200) );
  NAND U9323 ( .A(n8399), .B(n8198), .Z(n8199) );
  NAND U9324 ( .A(n8200), .B(n8199), .Z(n8291) );
  AND U9325 ( .A(x[224]), .B(y[1878]), .Z(n8325) );
  AND U9326 ( .A(x[246]), .B(y[1856]), .Z(n8326) );
  XOR U9327 ( .A(n8325), .B(n8326), .Z(n8328) );
  NAND U9328 ( .A(x[245]), .B(y[1857]), .Z(n8348) );
  XOR U9329 ( .A(n8328), .B(n8327), .Z(n8289) );
  AND U9330 ( .A(y[1871]), .B(x[231]), .Z(n8202) );
  NAND U9331 ( .A(y[1870]), .B(x[232]), .Z(n8201) );
  XNOR U9332 ( .A(n8202), .B(n8201), .Z(n8331) );
  XOR U9333 ( .A(n8289), .B(n8288), .Z(n8290) );
  XOR U9334 ( .A(n8291), .B(n8290), .Z(n8278) );
  XOR U9335 ( .A(n8279), .B(n8278), .Z(n8362) );
  XOR U9336 ( .A(n8363), .B(n8362), .Z(n8356) );
  XOR U9337 ( .A(n8357), .B(n8356), .Z(n8373) );
  XOR U9338 ( .A(n8372), .B(n8373), .Z(n8374) );
  XOR U9339 ( .A(n8375), .B(n8374), .Z(n8267) );
  NAND U9340 ( .A(n8204), .B(n8203), .Z(n8208) );
  NAND U9341 ( .A(n8206), .B(n8205), .Z(n8207) );
  NAND U9342 ( .A(n8208), .B(n8207), .Z(n8273) );
  NAND U9343 ( .A(n8210), .B(n8209), .Z(n8214) );
  NAND U9344 ( .A(n8212), .B(n8211), .Z(n8213) );
  NAND U9345 ( .A(n8214), .B(n8213), .Z(n8271) );
  NAND U9346 ( .A(n8216), .B(n8215), .Z(n8220) );
  NAND U9347 ( .A(n8218), .B(n8217), .Z(n8219) );
  NAND U9348 ( .A(n8220), .B(n8219), .Z(n8270) );
  XOR U9349 ( .A(n8271), .B(n8270), .Z(n8272) );
  XOR U9350 ( .A(n8273), .B(n8272), .Z(n8265) );
  NANDN U9351 ( .A(n8222), .B(n8221), .Z(n8226) );
  NAND U9352 ( .A(n8224), .B(n8223), .Z(n8225) );
  NAND U9353 ( .A(n8226), .B(n8225), .Z(n8264) );
  NAND U9354 ( .A(n8228), .B(n8227), .Z(n8232) );
  NANDN U9355 ( .A(n8230), .B(n8229), .Z(n8231) );
  NAND U9356 ( .A(n8232), .B(n8231), .Z(n8259) );
  NAND U9357 ( .A(n8234), .B(n8233), .Z(n8238) );
  NAND U9358 ( .A(n8236), .B(n8235), .Z(n8237) );
  NAND U9359 ( .A(n8238), .B(n8237), .Z(n8258) );
  XOR U9360 ( .A(n8259), .B(n8258), .Z(n8260) );
  XNOR U9361 ( .A(n8252), .B(n8251), .Z(n8255) );
  NANDN U9362 ( .A(n8243), .B(n8242), .Z(n8247) );
  NANDN U9363 ( .A(n8245), .B(n8244), .Z(n8246) );
  AND U9364 ( .A(n8247), .B(n8246), .Z(n8257) );
  XOR U9365 ( .A(n8256), .B(n8257), .Z(n8248) );
  XNOR U9366 ( .A(n8255), .B(n8248), .Z(N183) );
  NANDN U9367 ( .A(n8250), .B(n8249), .Z(n8254) );
  NAND U9368 ( .A(n8252), .B(n8251), .Z(n8253) );
  NAND U9369 ( .A(n8254), .B(n8253), .Z(n8512) );
  IV U9370 ( .A(n8512), .Z(n8511) );
  NAND U9371 ( .A(n8259), .B(n8258), .Z(n8263) );
  NANDN U9372 ( .A(n8261), .B(n8260), .Z(n8262) );
  AND U9373 ( .A(n8263), .B(n8262), .Z(n8520) );
  NANDN U9374 ( .A(n8265), .B(n8264), .Z(n8269) );
  NANDN U9375 ( .A(n8267), .B(n8266), .Z(n8268) );
  NAND U9376 ( .A(n8269), .B(n8268), .Z(n8518) );
  NAND U9377 ( .A(n8271), .B(n8270), .Z(n8275) );
  NAND U9378 ( .A(n8273), .B(n8272), .Z(n8274) );
  NAND U9379 ( .A(n8275), .B(n8274), .Z(n8496) );
  NAND U9380 ( .A(n8277), .B(n8276), .Z(n8281) );
  NAND U9381 ( .A(n8279), .B(n8278), .Z(n8280) );
  NAND U9382 ( .A(n8281), .B(n8280), .Z(n8489) );
  NAND U9383 ( .A(n8283), .B(n8282), .Z(n8287) );
  NAND U9384 ( .A(n8285), .B(n8284), .Z(n8286) );
  NAND U9385 ( .A(n8287), .B(n8286), .Z(n8487) );
  NAND U9386 ( .A(n8289), .B(n8288), .Z(n8293) );
  NAND U9387 ( .A(n8291), .B(n8290), .Z(n8292) );
  NAND U9388 ( .A(n8293), .B(n8292), .Z(n8486) );
  XOR U9389 ( .A(n8487), .B(n8486), .Z(n8488) );
  XOR U9390 ( .A(n8489), .B(n8488), .Z(n8508) );
  NAND U9391 ( .A(n8295), .B(n8294), .Z(n8299) );
  NAND U9392 ( .A(n8297), .B(n8296), .Z(n8298) );
  NAND U9393 ( .A(n8299), .B(n8298), .Z(n8506) );
  NAND U9394 ( .A(n8301), .B(n8300), .Z(n8305) );
  NAND U9395 ( .A(n8303), .B(n8302), .Z(n8304) );
  NAND U9396 ( .A(n8305), .B(n8304), .Z(n8433) );
  AND U9397 ( .A(n8307), .B(n8306), .Z(n8311) );
  NAND U9398 ( .A(n8309), .B(n8308), .Z(n8310) );
  NANDN U9399 ( .A(n8311), .B(n8310), .Z(n8432) );
  XOR U9400 ( .A(n8433), .B(n8432), .Z(n8435) );
  AND U9401 ( .A(y[1872]), .B(x[231]), .Z(n8313) );
  NAND U9402 ( .A(y[1870]), .B(x[233]), .Z(n8312) );
  XNOR U9403 ( .A(n8313), .B(n8312), .Z(n8400) );
  NAND U9404 ( .A(x[234]), .B(y[1869]), .Z(n8439) );
  AND U9405 ( .A(x[230]), .B(y[1873]), .Z(n8391) );
  NAND U9406 ( .A(x[239]), .B(y[1864]), .Z(n8392) );
  NAND U9407 ( .A(x[235]), .B(y[1868]), .Z(n8394) );
  XOR U9408 ( .A(n8441), .B(n8440), .Z(n8434) );
  XOR U9409 ( .A(n8435), .B(n8434), .Z(n8505) );
  XOR U9410 ( .A(n8506), .B(n8505), .Z(n8507) );
  XOR U9411 ( .A(n8508), .B(n8507), .Z(n8494) );
  NAND U9412 ( .A(n8315), .B(n8314), .Z(n8319) );
  NAND U9413 ( .A(n8317), .B(n8316), .Z(n8318) );
  NAND U9414 ( .A(n8319), .B(n8318), .Z(n8427) );
  AND U9415 ( .A(x[242]), .B(y[1866]), .Z(n9220) );
  NAND U9416 ( .A(n9220), .B(n8320), .Z(n8324) );
  NAND U9417 ( .A(n8322), .B(n8321), .Z(n8323) );
  NAND U9418 ( .A(n8324), .B(n8323), .Z(n8463) );
  NAND U9419 ( .A(n8326), .B(n8325), .Z(n8330) );
  NAND U9420 ( .A(n8328), .B(n8327), .Z(n8329) );
  NAND U9421 ( .A(n8330), .B(n8329), .Z(n8462) );
  XOR U9422 ( .A(n8463), .B(n8462), .Z(n8464) );
  NANDN U9423 ( .A(n8401), .B(n8399), .Z(n8334) );
  NANDN U9424 ( .A(n8332), .B(n8331), .Z(n8333) );
  NAND U9425 ( .A(n8334), .B(n8333), .Z(n8476) );
  AND U9426 ( .A(x[224]), .B(y[1879]), .Z(n8410) );
  NAND U9427 ( .A(x[247]), .B(y[1856]), .Z(n8411) );
  NAND U9428 ( .A(x[246]), .B(y[1857]), .Z(n8390) );
  XOR U9429 ( .A(n8413), .B(n8412), .Z(n8475) );
  NAND U9430 ( .A(y[1859]), .B(x[244]), .Z(n8335) );
  XNOR U9431 ( .A(n8336), .B(n8335), .Z(n8386) );
  NAND U9432 ( .A(x[243]), .B(y[1860]), .Z(n8387) );
  XOR U9433 ( .A(n8475), .B(n8474), .Z(n8477) );
  XOR U9434 ( .A(n8476), .B(n8477), .Z(n8465) );
  XOR U9435 ( .A(n8464), .B(n8465), .Z(n8426) );
  XOR U9436 ( .A(n8427), .B(n8426), .Z(n8429) );
  AND U9437 ( .A(x[244]), .B(y[1865]), .Z(n9196) );
  IV U9438 ( .A(n9196), .Z(n9383) );
  AND U9439 ( .A(x[237]), .B(y[1858]), .Z(n8337) );
  NANDN U9440 ( .A(n9383), .B(n8337), .Z(n8341) );
  NAND U9441 ( .A(n8339), .B(n8338), .Z(n8340) );
  NAND U9442 ( .A(n8341), .B(n8340), .Z(n8421) );
  NAND U9443 ( .A(n8343), .B(n8342), .Z(n8347) );
  NAND U9444 ( .A(n8345), .B(n8344), .Z(n8346) );
  NAND U9445 ( .A(n8347), .B(n8346), .Z(n8482) );
  AND U9446 ( .A(x[237]), .B(y[1866]), .Z(n8456) );
  AND U9447 ( .A(x[226]), .B(y[1877]), .Z(n8457) );
  XOR U9448 ( .A(n8456), .B(n8457), .Z(n8458) );
  AND U9449 ( .A(x[245]), .B(y[1858]), .Z(n8459) );
  XOR U9450 ( .A(n8458), .B(n8459), .Z(n8481) );
  AND U9451 ( .A(x[236]), .B(y[1867]), .Z(n8404) );
  NAND U9452 ( .A(x[225]), .B(y[1878]), .Z(n8405) );
  ANDN U9453 ( .B(o[86]), .A(n8348), .Z(n8406) );
  XOR U9454 ( .A(n8407), .B(n8406), .Z(n8480) );
  XOR U9455 ( .A(n8481), .B(n8480), .Z(n8483) );
  XOR U9456 ( .A(n8482), .B(n8483), .Z(n8420) );
  XOR U9457 ( .A(n8421), .B(n8420), .Z(n8423) );
  AND U9458 ( .A(x[239]), .B(y[1872]), .Z(n9618) );
  NAND U9459 ( .A(n9618), .B(n8349), .Z(n8353) );
  NANDN U9460 ( .A(n8351), .B(n8350), .Z(n8352) );
  NAND U9461 ( .A(n8353), .B(n8352), .Z(n8470) );
  AND U9462 ( .A(x[238]), .B(y[1865]), .Z(n8450) );
  AND U9463 ( .A(x[227]), .B(y[1876]), .Z(n8451) );
  XOR U9464 ( .A(n8450), .B(n8451), .Z(n8452) );
  AND U9465 ( .A(x[228]), .B(y[1875]), .Z(n8453) );
  XOR U9466 ( .A(n8452), .B(n8453), .Z(n8469) );
  AND U9467 ( .A(x[229]), .B(y[1874]), .Z(n8444) );
  AND U9468 ( .A(x[242]), .B(y[1861]), .Z(n8445) );
  XOR U9469 ( .A(n8444), .B(n8445), .Z(n8447) );
  AND U9470 ( .A(x[241]), .B(y[1862]), .Z(n8446) );
  XOR U9471 ( .A(n8447), .B(n8446), .Z(n8468) );
  XOR U9472 ( .A(n8469), .B(n8468), .Z(n8471) );
  XOR U9473 ( .A(n8470), .B(n8471), .Z(n8422) );
  XOR U9474 ( .A(n8423), .B(n8422), .Z(n8428) );
  XOR U9475 ( .A(n8429), .B(n8428), .Z(n8493) );
  XOR U9476 ( .A(n8494), .B(n8493), .Z(n8495) );
  XNOR U9477 ( .A(n8496), .B(n8495), .Z(n8381) );
  NAND U9478 ( .A(n8355), .B(n8354), .Z(n8359) );
  NAND U9479 ( .A(n8357), .B(n8356), .Z(n8358) );
  NAND U9480 ( .A(n8359), .B(n8358), .Z(n8502) );
  NAND U9481 ( .A(n8361), .B(n8360), .Z(n8365) );
  NAND U9482 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U9483 ( .A(n8365), .B(n8364), .Z(n8500) );
  NAND U9484 ( .A(n8367), .B(n8366), .Z(n8371) );
  NAND U9485 ( .A(n8369), .B(n8368), .Z(n8370) );
  AND U9486 ( .A(n8371), .B(n8370), .Z(n8499) );
  XOR U9487 ( .A(n8500), .B(n8499), .Z(n8501) );
  XNOR U9488 ( .A(n8502), .B(n8501), .Z(n8379) );
  NAND U9489 ( .A(n8373), .B(n8372), .Z(n8377) );
  NAND U9490 ( .A(n8375), .B(n8374), .Z(n8376) );
  AND U9491 ( .A(n8377), .B(n8376), .Z(n8380) );
  XOR U9492 ( .A(n8379), .B(n8380), .Z(n8382) );
  XNOR U9493 ( .A(n8381), .B(n8382), .Z(n8519) );
  XNOR U9494 ( .A(n8520), .B(n8521), .Z(n8514) );
  XNOR U9495 ( .A(n8513), .B(n8514), .Z(n8378) );
  XOR U9496 ( .A(n8511), .B(n8378), .Z(N184) );
  NAND U9497 ( .A(n8380), .B(n8379), .Z(n8384) );
  NAND U9498 ( .A(n8382), .B(n8381), .Z(n8383) );
  AND U9499 ( .A(n8384), .B(n8383), .Z(n8667) );
  AND U9500 ( .A(x[244]), .B(y[1863]), .Z(n8385) );
  NAND U9501 ( .A(n8385), .B(n8627), .Z(n8389) );
  NANDN U9502 ( .A(n8387), .B(n8386), .Z(n8388) );
  AND U9503 ( .A(n8389), .B(n8388), .Z(n8648) );
  AND U9504 ( .A(x[246]), .B(y[1858]), .Z(n8554) );
  XOR U9505 ( .A(n8555), .B(n8554), .Z(n8557) );
  NAND U9506 ( .A(x[226]), .B(y[1878]), .Z(n8556) );
  AND U9507 ( .A(x[225]), .B(y[1879]), .Z(n8562) );
  XOR U9508 ( .A(n8563), .B(n8562), .Z(n8561) );
  ANDN U9509 ( .B(o[87]), .A(n8390), .Z(n8560) );
  XOR U9510 ( .A(n8561), .B(n8560), .Z(n8645) );
  XOR U9511 ( .A(n8646), .B(n8645), .Z(n8647) );
  NANDN U9512 ( .A(n8392), .B(n8391), .Z(n8396) );
  NANDN U9513 ( .A(n8394), .B(n8393), .Z(n8395) );
  AND U9514 ( .A(n8396), .B(n8395), .Z(n8642) );
  AND U9515 ( .A(y[1864]), .B(x[240]), .Z(n8398) );
  NAND U9516 ( .A(y[1859]), .B(x[245]), .Z(n8397) );
  XNOR U9517 ( .A(n8398), .B(n8397), .Z(n8628) );
  NAND U9518 ( .A(x[229]), .B(y[1875]), .Z(n8629) );
  AND U9519 ( .A(x[230]), .B(y[1874]), .Z(n8956) );
  NAND U9520 ( .A(x[244]), .B(y[1860]), .Z(n8634) );
  IV U9521 ( .A(n8634), .Z(n8770) );
  XOR U9522 ( .A(n8956), .B(n8770), .Z(n8635) );
  NAND U9523 ( .A(x[243]), .B(y[1861]), .Z(n8636) );
  XOR U9524 ( .A(n8640), .B(n8639), .Z(n8641) );
  NANDN U9525 ( .A(n8696), .B(n8399), .Z(n8403) );
  NANDN U9526 ( .A(n8401), .B(n8400), .Z(n8402) );
  NAND U9527 ( .A(n8403), .B(n8402), .Z(n8616) );
  NANDN U9528 ( .A(n8405), .B(n8404), .Z(n8409) );
  NAND U9529 ( .A(n8407), .B(n8406), .Z(n8408) );
  NAND U9530 ( .A(n8409), .B(n8408), .Z(n8615) );
  XNOR U9531 ( .A(n8616), .B(n8615), .Z(n8618) );
  XOR U9532 ( .A(n8592), .B(n8591), .Z(n8594) );
  NANDN U9533 ( .A(n8411), .B(n8410), .Z(n8415) );
  NAND U9534 ( .A(n8413), .B(n8412), .Z(n8414) );
  AND U9535 ( .A(n8415), .B(n8414), .Z(n8574) );
  AND U9536 ( .A(x[227]), .B(y[1877]), .Z(n8579) );
  XOR U9537 ( .A(n8580), .B(n8579), .Z(n8582) );
  NAND U9538 ( .A(x[228]), .B(y[1876]), .Z(n8581) );
  AND U9539 ( .A(y[1871]), .B(x[233]), .Z(n8417) );
  NAND U9540 ( .A(y[1870]), .B(x[234]), .Z(n8416) );
  XNOR U9541 ( .A(n8417), .B(n8416), .Z(n8546) );
  AND U9542 ( .A(y[1866]), .B(x[238]), .Z(n8419) );
  NAND U9543 ( .A(y[1872]), .B(x[232]), .Z(n8418) );
  XNOR U9544 ( .A(n8419), .B(n8418), .Z(n8550) );
  NAND U9545 ( .A(x[235]), .B(y[1869]), .Z(n8551) );
  XOR U9546 ( .A(n8546), .B(n8545), .Z(n8575) );
  XOR U9547 ( .A(n8576), .B(n8575), .Z(n8593) );
  XOR U9548 ( .A(n8594), .B(n8593), .Z(n8539) );
  NAND U9549 ( .A(n8421), .B(n8420), .Z(n8425) );
  NAND U9550 ( .A(n8423), .B(n8422), .Z(n8424) );
  AND U9551 ( .A(n8425), .B(n8424), .Z(n8538) );
  NAND U9552 ( .A(n8427), .B(n8426), .Z(n8431) );
  NAND U9553 ( .A(n8429), .B(n8428), .Z(n8430) );
  NAND U9554 ( .A(n8431), .B(n8430), .Z(n8541) );
  NAND U9555 ( .A(n8433), .B(n8432), .Z(n8437) );
  NAND U9556 ( .A(n8435), .B(n8434), .Z(n8436) );
  AND U9557 ( .A(n8437), .B(n8436), .Z(n8600) );
  NANDN U9558 ( .A(n8439), .B(n8438), .Z(n8443) );
  NAND U9559 ( .A(n8441), .B(n8440), .Z(n8442) );
  AND U9560 ( .A(n8443), .B(n8442), .Z(n8598) );
  NAND U9561 ( .A(n8445), .B(n8444), .Z(n8449) );
  NAND U9562 ( .A(n8447), .B(n8446), .Z(n8448) );
  AND U9563 ( .A(n8449), .B(n8448), .Z(n8624) );
  AND U9564 ( .A(x[224]), .B(y[1880]), .Z(n8585) );
  NAND U9565 ( .A(x[248]), .B(y[1856]), .Z(n8586) );
  NAND U9566 ( .A(x[247]), .B(y[1857]), .Z(n8572) );
  XOR U9567 ( .A(n8588), .B(n8587), .Z(n8622) );
  AND U9568 ( .A(x[231]), .B(y[1873]), .Z(n8566) );
  NAND U9569 ( .A(x[242]), .B(y[1862]), .Z(n8567) );
  NAND U9570 ( .A(x[241]), .B(y[1863]), .Z(n8569) );
  XOR U9571 ( .A(n8622), .B(n8621), .Z(n8623) );
  NAND U9572 ( .A(n8451), .B(n8450), .Z(n8455) );
  NAND U9573 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U9574 ( .A(n8455), .B(n8454), .Z(n8610) );
  NAND U9575 ( .A(n8457), .B(n8456), .Z(n8461) );
  NAND U9576 ( .A(n8459), .B(n8458), .Z(n8460) );
  NAND U9577 ( .A(n8461), .B(n8460), .Z(n8609) );
  XNOR U9578 ( .A(n8610), .B(n8609), .Z(n8612) );
  NAND U9579 ( .A(n8463), .B(n8462), .Z(n8467) );
  NAND U9580 ( .A(n8465), .B(n8464), .Z(n8466) );
  AND U9581 ( .A(n8467), .B(n8466), .Z(n8654) );
  NAND U9582 ( .A(n8469), .B(n8468), .Z(n8473) );
  NAND U9583 ( .A(n8471), .B(n8470), .Z(n8472) );
  AND U9584 ( .A(n8473), .B(n8472), .Z(n8652) );
  NAND U9585 ( .A(n8475), .B(n8474), .Z(n8479) );
  NAND U9586 ( .A(n8477), .B(n8476), .Z(n8478) );
  AND U9587 ( .A(n8479), .B(n8478), .Z(n8651) );
  XOR U9588 ( .A(n8652), .B(n8651), .Z(n8653) );
  XOR U9589 ( .A(n8654), .B(n8653), .Z(n8603) );
  NAND U9590 ( .A(n8481), .B(n8480), .Z(n8485) );
  NAND U9591 ( .A(n8483), .B(n8482), .Z(n8484) );
  NAND U9592 ( .A(n8485), .B(n8484), .Z(n8604) );
  XOR U9593 ( .A(n8605), .B(n8606), .Z(n8532) );
  IV U9594 ( .A(n8532), .Z(n8531) );
  NAND U9595 ( .A(n8487), .B(n8486), .Z(n8491) );
  NAND U9596 ( .A(n8489), .B(n8488), .Z(n8490) );
  AND U9597 ( .A(n8491), .B(n8490), .Z(n8533) );
  XOR U9598 ( .A(n8531), .B(n8533), .Z(n8492) );
  XOR U9599 ( .A(n8535), .B(n8492), .Z(n8664) );
  NAND U9600 ( .A(n8494), .B(n8493), .Z(n8498) );
  NAND U9601 ( .A(n8496), .B(n8495), .Z(n8497) );
  NAND U9602 ( .A(n8498), .B(n8497), .Z(n8528) );
  NAND U9603 ( .A(n8500), .B(n8499), .Z(n8504) );
  NAND U9604 ( .A(n8502), .B(n8501), .Z(n8503) );
  NAND U9605 ( .A(n8504), .B(n8503), .Z(n8526) );
  NAND U9606 ( .A(n8506), .B(n8505), .Z(n8510) );
  NAND U9607 ( .A(n8508), .B(n8507), .Z(n8509) );
  NAND U9608 ( .A(n8510), .B(n8509), .Z(n8525) );
  XOR U9609 ( .A(n8526), .B(n8525), .Z(n8527) );
  XOR U9610 ( .A(n8528), .B(n8527), .Z(n8665) );
  XOR U9611 ( .A(n8664), .B(n8665), .Z(n8666) );
  XNOR U9612 ( .A(n8667), .B(n8666), .Z(n8660) );
  OR U9613 ( .A(n8513), .B(n8511), .Z(n8517) );
  ANDN U9614 ( .B(n8513), .A(n8512), .Z(n8515) );
  OR U9615 ( .A(n8515), .B(n8514), .Z(n8516) );
  AND U9616 ( .A(n8517), .B(n8516), .Z(n8659) );
  NANDN U9617 ( .A(n8519), .B(n8518), .Z(n8523) );
  NANDN U9618 ( .A(n8521), .B(n8520), .Z(n8522) );
  AND U9619 ( .A(n8523), .B(n8522), .Z(n8658) );
  IV U9620 ( .A(n8658), .Z(n8657) );
  XOR U9621 ( .A(n8659), .B(n8657), .Z(n8524) );
  XNOR U9622 ( .A(n8660), .B(n8524), .Z(N185) );
  NAND U9623 ( .A(n8526), .B(n8525), .Z(n8530) );
  NAND U9624 ( .A(n8528), .B(n8527), .Z(n8529) );
  AND U9625 ( .A(n8530), .B(n8529), .Z(n8822) );
  NANDN U9626 ( .A(n8531), .B(n8533), .Z(n8537) );
  OR U9627 ( .A(n8533), .B(n8532), .Z(n8534) );
  NAND U9628 ( .A(n8535), .B(n8534), .Z(n8536) );
  NAND U9629 ( .A(n8537), .B(n8536), .Z(n8820) );
  NANDN U9630 ( .A(n8539), .B(n8538), .Z(n8543) );
  NANDN U9631 ( .A(n8541), .B(n8540), .Z(n8542) );
  AND U9632 ( .A(n8543), .B(n8542), .Z(n8672) );
  NANDN U9633 ( .A(n8695), .B(n8544), .Z(n8548) );
  NAND U9634 ( .A(n8546), .B(n8545), .Z(n8547) );
  AND U9635 ( .A(n8548), .B(n8547), .Z(n8720) );
  AND U9636 ( .A(x[238]), .B(y[1872]), .Z(n9606) );
  NAND U9637 ( .A(n9606), .B(n8549), .Z(n8553) );
  NANDN U9638 ( .A(n8551), .B(n8550), .Z(n8552) );
  NAND U9639 ( .A(n8553), .B(n8552), .Z(n8747) );
  NAND U9640 ( .A(x[235]), .B(y[1870]), .Z(n8766) );
  NAND U9641 ( .A(x[236]), .B(y[1869]), .Z(n8765) );
  NAND U9642 ( .A(x[231]), .B(y[1874]), .Z(n8764) );
  XOR U9643 ( .A(n8765), .B(n8764), .Z(n8767) );
  XOR U9644 ( .A(n8766), .B(n8767), .Z(n8746) );
  NAND U9645 ( .A(x[248]), .B(y[1857]), .Z(n8763) );
  AND U9646 ( .A(x[225]), .B(y[1880]), .Z(n8733) );
  XOR U9647 ( .A(n8734), .B(n8733), .Z(n8736) );
  AND U9648 ( .A(x[237]), .B(y[1868]), .Z(n8735) );
  XOR U9649 ( .A(n8736), .B(n8735), .Z(n8745) );
  XOR U9650 ( .A(n8747), .B(n8748), .Z(n8719) );
  NAND U9651 ( .A(n8555), .B(n8554), .Z(n8559) );
  ANDN U9652 ( .B(n8557), .A(n8556), .Z(n8558) );
  ANDN U9653 ( .B(n8559), .A(n8558), .Z(n8708) );
  AND U9654 ( .A(n8561), .B(n8560), .Z(n8565) );
  NAND U9655 ( .A(n8563), .B(n8562), .Z(n8564) );
  NANDN U9656 ( .A(n8565), .B(n8564), .Z(n8707) );
  NANDN U9657 ( .A(n8567), .B(n8566), .Z(n8571) );
  NANDN U9658 ( .A(n8569), .B(n8568), .Z(n8570) );
  AND U9659 ( .A(n8571), .B(n8570), .Z(n8704) );
  NAND U9660 ( .A(x[232]), .B(y[1873]), .Z(n8697) );
  XNOR U9661 ( .A(n8696), .B(n8695), .Z(n8698) );
  NANDN U9662 ( .A(n8572), .B(o[88]), .Z(n8691) );
  NAND U9663 ( .A(x[249]), .B(y[1856]), .Z(n8690) );
  NAND U9664 ( .A(x[224]), .B(y[1881]), .Z(n8689) );
  XNOR U9665 ( .A(n8690), .B(n8689), .Z(n8692) );
  XOR U9666 ( .A(n8691), .B(n8692), .Z(n8701) );
  XOR U9667 ( .A(n8702), .B(n8701), .Z(n8703) );
  XOR U9668 ( .A(n8710), .B(n8709), .Z(n8721) );
  XOR U9669 ( .A(n8722), .B(n8721), .Z(n8803) );
  NANDN U9670 ( .A(n8574), .B(n8573), .Z(n8578) );
  NAND U9671 ( .A(n8576), .B(n8575), .Z(n8577) );
  AND U9672 ( .A(n8578), .B(n8577), .Z(n8800) );
  NAND U9673 ( .A(n8580), .B(n8579), .Z(n8584) );
  ANDN U9674 ( .B(n8582), .A(n8581), .Z(n8583) );
  ANDN U9675 ( .B(n8584), .A(n8583), .Z(n8785) );
  NANDN U9676 ( .A(n8586), .B(n8585), .Z(n8590) );
  NAND U9677 ( .A(n8588), .B(n8587), .Z(n8589) );
  AND U9678 ( .A(n8590), .B(n8589), .Z(n8783) );
  AND U9679 ( .A(x[238]), .B(y[1867]), .Z(n8740) );
  AND U9680 ( .A(x[226]), .B(y[1879]), .Z(n8739) );
  XOR U9681 ( .A(n8740), .B(n8739), .Z(n8742) );
  AND U9682 ( .A(x[227]), .B(y[1878]), .Z(n8741) );
  XOR U9683 ( .A(n8742), .B(n8741), .Z(n8782) );
  NAND U9684 ( .A(n8592), .B(n8591), .Z(n8596) );
  NAND U9685 ( .A(n8594), .B(n8593), .Z(n8595) );
  AND U9686 ( .A(n8596), .B(n8595), .Z(n8806) );
  XOR U9687 ( .A(n8807), .B(n8806), .Z(n8809) );
  NANDN U9688 ( .A(n8598), .B(n8597), .Z(n8602) );
  NANDN U9689 ( .A(n8600), .B(n8599), .Z(n8601) );
  AND U9690 ( .A(n8602), .B(n8601), .Z(n8808) );
  XOR U9691 ( .A(n8809), .B(n8808), .Z(n8671) );
  NANDN U9692 ( .A(n8604), .B(n8603), .Z(n8608) );
  NAND U9693 ( .A(n8606), .B(n8605), .Z(n8607) );
  NAND U9694 ( .A(n8608), .B(n8607), .Z(n8679) );
  NAND U9695 ( .A(n8610), .B(n8609), .Z(n8614) );
  NANDN U9696 ( .A(n8612), .B(n8611), .Z(n8613) );
  NAND U9697 ( .A(n8614), .B(n8613), .Z(n8684) );
  NAND U9698 ( .A(n8616), .B(n8615), .Z(n8620) );
  NANDN U9699 ( .A(n8618), .B(n8617), .Z(n8619) );
  NAND U9700 ( .A(n8620), .B(n8619), .Z(n8683) );
  XOR U9701 ( .A(n8684), .B(n8683), .Z(n8685) );
  NAND U9702 ( .A(n8622), .B(n8621), .Z(n8626) );
  NANDN U9703 ( .A(n8624), .B(n8623), .Z(n8625) );
  AND U9704 ( .A(n8626), .B(n8625), .Z(n8716) );
  AND U9705 ( .A(x[245]), .B(y[1864]), .Z(n9195) );
  IV U9706 ( .A(n9195), .Z(n9626) );
  NANDN U9707 ( .A(n9626), .B(n8627), .Z(n8631) );
  NANDN U9708 ( .A(n8629), .B(n8628), .Z(n8630) );
  AND U9709 ( .A(n8631), .B(n8630), .Z(n8791) );
  NAND U9710 ( .A(x[246]), .B(y[1859]), .Z(n8759) );
  NAND U9711 ( .A(x[229]), .B(y[1876]), .Z(n8758) );
  NAND U9712 ( .A(x[241]), .B(y[1864]), .Z(n8757) );
  XNOR U9713 ( .A(n8758), .B(n8757), .Z(n8760) );
  AND U9714 ( .A(y[1861]), .B(x[244]), .Z(n8633) );
  NAND U9715 ( .A(y[1860]), .B(x[245]), .Z(n8632) );
  XNOR U9716 ( .A(n8633), .B(n8632), .Z(n8772) );
  AND U9717 ( .A(x[243]), .B(y[1862]), .Z(n8771) );
  XOR U9718 ( .A(n8772), .B(n8771), .Z(n8789) );
  XOR U9719 ( .A(n8788), .B(n8789), .Z(n8790) );
  NANDN U9720 ( .A(n8634), .B(n8956), .Z(n8638) );
  NANDN U9721 ( .A(n8636), .B(n8635), .Z(n8637) );
  AND U9722 ( .A(n8638), .B(n8637), .Z(n8797) );
  NAND U9723 ( .A(x[239]), .B(y[1866]), .Z(n8778) );
  NAND U9724 ( .A(x[242]), .B(y[1863]), .Z(n8777) );
  NAND U9725 ( .A(x[230]), .B(y[1875]), .Z(n8776) );
  XNOR U9726 ( .A(n8777), .B(n8776), .Z(n8779) );
  NAND U9727 ( .A(x[247]), .B(y[1858]), .Z(n8753) );
  NAND U9728 ( .A(x[228]), .B(y[1877]), .Z(n8752) );
  NAND U9729 ( .A(x[240]), .B(y[1865]), .Z(n8751) );
  XNOR U9730 ( .A(n8752), .B(n8751), .Z(n8754) );
  XOR U9731 ( .A(n8753), .B(n8754), .Z(n8794) );
  XOR U9732 ( .A(n8795), .B(n8794), .Z(n8796) );
  XOR U9733 ( .A(n8797), .B(n8796), .Z(n8713) );
  XOR U9734 ( .A(n8714), .B(n8713), .Z(n8715) );
  XOR U9735 ( .A(n8716), .B(n8715), .Z(n8728) );
  NAND U9736 ( .A(n8640), .B(n8639), .Z(n8644) );
  NANDN U9737 ( .A(n8642), .B(n8641), .Z(n8643) );
  AND U9738 ( .A(n8644), .B(n8643), .Z(n8726) );
  NAND U9739 ( .A(n8646), .B(n8645), .Z(n8650) );
  NANDN U9740 ( .A(n8648), .B(n8647), .Z(n8649) );
  NAND U9741 ( .A(n8650), .B(n8649), .Z(n8725) );
  XNOR U9742 ( .A(n8685), .B(n8686), .Z(n8678) );
  NAND U9743 ( .A(n8652), .B(n8651), .Z(n8656) );
  NAND U9744 ( .A(n8654), .B(n8653), .Z(n8655) );
  NAND U9745 ( .A(n8656), .B(n8655), .Z(n8677) );
  XOR U9746 ( .A(n8679), .B(n8680), .Z(n8673) );
  XOR U9747 ( .A(n8674), .B(n8673), .Z(n8819) );
  XOR U9748 ( .A(n8820), .B(n8819), .Z(n8821) );
  XNOR U9749 ( .A(n8822), .B(n8821), .Z(n8815) );
  OR U9750 ( .A(n8659), .B(n8657), .Z(n8663) );
  ANDN U9751 ( .B(n8659), .A(n8658), .Z(n8661) );
  OR U9752 ( .A(n8661), .B(n8660), .Z(n8662) );
  AND U9753 ( .A(n8663), .B(n8662), .Z(n8813) );
  NAND U9754 ( .A(n8665), .B(n8664), .Z(n8669) );
  NAND U9755 ( .A(n8667), .B(n8666), .Z(n8668) );
  AND U9756 ( .A(n8669), .B(n8668), .Z(n8814) );
  IV U9757 ( .A(n8814), .Z(n8812) );
  XOR U9758 ( .A(n8813), .B(n8812), .Z(n8670) );
  XNOR U9759 ( .A(n8815), .B(n8670), .Z(N186) );
  NANDN U9760 ( .A(n8672), .B(n8671), .Z(n8676) );
  NAND U9761 ( .A(n8674), .B(n8673), .Z(n8675) );
  AND U9762 ( .A(n8676), .B(n8675), .Z(n8826) );
  NANDN U9763 ( .A(n8678), .B(n8677), .Z(n8682) );
  NAND U9764 ( .A(n8680), .B(n8679), .Z(n8681) );
  NAND U9765 ( .A(n8682), .B(n8681), .Z(n8827) );
  NAND U9766 ( .A(n8684), .B(n8683), .Z(n8688) );
  NANDN U9767 ( .A(n8686), .B(n8685), .Z(n8687) );
  NAND U9768 ( .A(n8688), .B(n8687), .Z(n8843) );
  AND U9769 ( .A(x[226]), .B(y[1880]), .Z(n8865) );
  XOR U9770 ( .A(n8866), .B(n8865), .Z(n8868) );
  NAND U9771 ( .A(x[248]), .B(y[1858]), .Z(n8867) );
  NAND U9772 ( .A(n8690), .B(n8689), .Z(n8694) );
  NANDN U9773 ( .A(n8692), .B(n8691), .Z(n8693) );
  AND U9774 ( .A(n8694), .B(n8693), .Z(n8907) );
  XOR U9775 ( .A(n8908), .B(n8907), .Z(n8910) );
  NAND U9776 ( .A(n8696), .B(n8695), .Z(n8700) );
  NANDN U9777 ( .A(n8698), .B(n8697), .Z(n8699) );
  AND U9778 ( .A(n8700), .B(n8699), .Z(n8909) );
  XOR U9779 ( .A(n8910), .B(n8909), .Z(n8971) );
  NAND U9780 ( .A(n8702), .B(n8701), .Z(n8706) );
  NANDN U9781 ( .A(n8704), .B(n8703), .Z(n8705) );
  AND U9782 ( .A(n8706), .B(n8705), .Z(n8970) );
  NANDN U9783 ( .A(n8708), .B(n8707), .Z(n8712) );
  NAND U9784 ( .A(n8710), .B(n8709), .Z(n8711) );
  NAND U9785 ( .A(n8712), .B(n8711), .Z(n8973) );
  NAND U9786 ( .A(n8714), .B(n8713), .Z(n8718) );
  NAND U9787 ( .A(n8716), .B(n8715), .Z(n8717) );
  AND U9788 ( .A(n8718), .B(n8717), .Z(n8933) );
  NANDN U9789 ( .A(n8720), .B(n8719), .Z(n8724) );
  NAND U9790 ( .A(n8722), .B(n8721), .Z(n8723) );
  AND U9791 ( .A(n8724), .B(n8723), .Z(n8932) );
  XOR U9792 ( .A(n8935), .B(n8934), .Z(n8842) );
  NANDN U9793 ( .A(n8726), .B(n8725), .Z(n8730) );
  NANDN U9794 ( .A(n8728), .B(n8727), .Z(n8729) );
  AND U9795 ( .A(n8730), .B(n8729), .Z(n8850) );
  AND U9796 ( .A(x[236]), .B(y[1870]), .Z(n9033) );
  AND U9797 ( .A(x[229]), .B(y[1877]), .Z(n8921) );
  XOR U9798 ( .A(n9033), .B(n8921), .Z(n8923) );
  NAND U9799 ( .A(x[234]), .B(y[1872]), .Z(n8922) );
  AND U9800 ( .A(x[231]), .B(y[1875]), .Z(n8939) );
  AND U9801 ( .A(y[1876]), .B(x[230]), .Z(n8732) );
  NAND U9802 ( .A(y[1874]), .B(x[232]), .Z(n8731) );
  XNOR U9803 ( .A(n8732), .B(n8731), .Z(n8957) );
  NAND U9804 ( .A(x[233]), .B(y[1873]), .Z(n8958) );
  XOR U9805 ( .A(n8939), .B(n8938), .Z(n8940) );
  XOR U9806 ( .A(n8941), .B(n8940), .Z(n8891) );
  NAND U9807 ( .A(n8734), .B(n8733), .Z(n8738) );
  NAND U9808 ( .A(n8736), .B(n8735), .Z(n8737) );
  NAND U9809 ( .A(n8738), .B(n8737), .Z(n8890) );
  NAND U9810 ( .A(n8740), .B(n8739), .Z(n8744) );
  NAND U9811 ( .A(n8742), .B(n8741), .Z(n8743) );
  NAND U9812 ( .A(n8744), .B(n8743), .Z(n8889) );
  XNOR U9813 ( .A(n8890), .B(n8889), .Z(n8892) );
  NANDN U9814 ( .A(n8746), .B(n8745), .Z(n8750) );
  NAND U9815 ( .A(n8748), .B(n8747), .Z(n8749) );
  AND U9816 ( .A(n8750), .B(n8749), .Z(n8895) );
  NAND U9817 ( .A(n8752), .B(n8751), .Z(n8756) );
  NANDN U9818 ( .A(n8754), .B(n8753), .Z(n8755) );
  AND U9819 ( .A(n8756), .B(n8755), .Z(n8854) );
  NAND U9820 ( .A(n8758), .B(n8757), .Z(n8762) );
  NANDN U9821 ( .A(n8760), .B(n8759), .Z(n8761) );
  AND U9822 ( .A(n8762), .B(n8761), .Z(n8853) );
  XOR U9823 ( .A(n8854), .B(n8853), .Z(n8856) );
  ANDN U9824 ( .B(o[89]), .A(n8763), .Z(n8950) );
  NAND U9825 ( .A(x[238]), .B(y[1868]), .Z(n8951) );
  NAND U9826 ( .A(x[225]), .B(y[1881]), .Z(n8953) );
  NAND U9827 ( .A(x[249]), .B(y[1857]), .Z(n8961) );
  XNOR U9828 ( .A(o[90]), .B(n8961), .Z(n8926) );
  NAND U9829 ( .A(x[250]), .B(y[1856]), .Z(n8927) );
  AND U9830 ( .A(x[224]), .B(y[1882]), .Z(n8928) );
  XOR U9831 ( .A(n8929), .B(n8928), .Z(n8913) );
  XOR U9832 ( .A(n8914), .B(n8913), .Z(n8916) );
  NAND U9833 ( .A(n8765), .B(n8764), .Z(n8769) );
  NAND U9834 ( .A(n8767), .B(n8766), .Z(n8768) );
  AND U9835 ( .A(n8769), .B(n8768), .Z(n8915) );
  XOR U9836 ( .A(n8916), .B(n8915), .Z(n8855) );
  XOR U9837 ( .A(n8856), .B(n8855), .Z(n8904) );
  AND U9838 ( .A(x[245]), .B(y[1861]), .Z(n8775) );
  IV U9839 ( .A(n8775), .Z(n8945) );
  NANDN U9840 ( .A(n8945), .B(n8770), .Z(n8774) );
  NAND U9841 ( .A(n8772), .B(n8771), .Z(n8773) );
  NAND U9842 ( .A(n8774), .B(n8773), .Z(n8885) );
  XOR U9843 ( .A(n8944), .B(n8775), .Z(n8947) );
  NAND U9844 ( .A(x[244]), .B(y[1862]), .Z(n8946) );
  NAND U9845 ( .A(x[247]), .B(y[1859]), .Z(n8872) );
  AND U9846 ( .A(x[246]), .B(y[1860]), .Z(n8873) );
  XOR U9847 ( .A(n8874), .B(n8873), .Z(n8883) );
  XOR U9848 ( .A(n8884), .B(n8883), .Z(n8886) );
  XOR U9849 ( .A(n8885), .B(n8886), .Z(n8902) );
  AND U9850 ( .A(x[228]), .B(y[1878]), .Z(n8877) );
  XOR U9851 ( .A(n8878), .B(n8877), .Z(n8880) );
  AND U9852 ( .A(x[227]), .B(y[1879]), .Z(n8962) );
  NAND U9853 ( .A(x[243]), .B(y[1863]), .Z(n8963) );
  AND U9854 ( .A(x[235]), .B(y[1871]), .Z(n8964) );
  XOR U9855 ( .A(n8965), .B(n8964), .Z(n8859) );
  XOR U9856 ( .A(n8860), .B(n8859), .Z(n8862) );
  NAND U9857 ( .A(n8777), .B(n8776), .Z(n8781) );
  NANDN U9858 ( .A(n8779), .B(n8778), .Z(n8780) );
  AND U9859 ( .A(n8781), .B(n8780), .Z(n8861) );
  XNOR U9860 ( .A(n8862), .B(n8861), .Z(n8901) );
  XOR U9861 ( .A(n8898), .B(n8897), .Z(n8848) );
  NANDN U9862 ( .A(n8783), .B(n8782), .Z(n8787) );
  NANDN U9863 ( .A(n8785), .B(n8784), .Z(n8786) );
  AND U9864 ( .A(n8787), .B(n8786), .Z(n8979) );
  NAND U9865 ( .A(n8789), .B(n8788), .Z(n8793) );
  NANDN U9866 ( .A(n8791), .B(n8790), .Z(n8792) );
  AND U9867 ( .A(n8793), .B(n8792), .Z(n8977) );
  NAND U9868 ( .A(n8795), .B(n8794), .Z(n8799) );
  NANDN U9869 ( .A(n8797), .B(n8796), .Z(n8798) );
  NAND U9870 ( .A(n8799), .B(n8798), .Z(n8976) );
  XOR U9871 ( .A(n8843), .B(n8844), .Z(n8838) );
  NANDN U9872 ( .A(n8801), .B(n8800), .Z(n8805) );
  NANDN U9873 ( .A(n8803), .B(n8802), .Z(n8804) );
  AND U9874 ( .A(n8805), .B(n8804), .Z(n8836) );
  NAND U9875 ( .A(n8807), .B(n8806), .Z(n8811) );
  NAND U9876 ( .A(n8809), .B(n8808), .Z(n8810) );
  AND U9877 ( .A(n8811), .B(n8810), .Z(n8835) );
  XOR U9878 ( .A(n8836), .B(n8835), .Z(n8837) );
  XOR U9879 ( .A(n8838), .B(n8837), .Z(n8828) );
  XNOR U9880 ( .A(n8829), .B(n8828), .Z(n8834) );
  NANDN U9881 ( .A(n8812), .B(n8813), .Z(n8818) );
  NOR U9882 ( .A(n8814), .B(n8813), .Z(n8816) );
  OR U9883 ( .A(n8816), .B(n8815), .Z(n8817) );
  AND U9884 ( .A(n8818), .B(n8817), .Z(n8832) );
  NAND U9885 ( .A(n8820), .B(n8819), .Z(n8824) );
  NAND U9886 ( .A(n8822), .B(n8821), .Z(n8823) );
  AND U9887 ( .A(n8824), .B(n8823), .Z(n8833) );
  XOR U9888 ( .A(n8832), .B(n8833), .Z(n8825) );
  XNOR U9889 ( .A(n8834), .B(n8825), .Z(N187) );
  NANDN U9890 ( .A(n8827), .B(n8826), .Z(n8831) );
  NAND U9891 ( .A(n8829), .B(n8828), .Z(n8830) );
  NAND U9892 ( .A(n8831), .B(n8830), .Z(n9127) );
  IV U9893 ( .A(n9127), .Z(n9126) );
  NAND U9894 ( .A(n8836), .B(n8835), .Z(n8840) );
  NAND U9895 ( .A(n8838), .B(n8837), .Z(n8839) );
  AND U9896 ( .A(n8840), .B(n8839), .Z(n9136) );
  NANDN U9897 ( .A(n8842), .B(n8841), .Z(n8846) );
  NAND U9898 ( .A(n8844), .B(n8843), .Z(n8845) );
  AND U9899 ( .A(n8846), .B(n8845), .Z(n9134) );
  NANDN U9900 ( .A(n8848), .B(n8847), .Z(n8852) );
  NANDN U9901 ( .A(n8850), .B(n8849), .Z(n8851) );
  NAND U9902 ( .A(n8852), .B(n8851), .Z(n8985) );
  NAND U9903 ( .A(n8854), .B(n8853), .Z(n8858) );
  NAND U9904 ( .A(n8856), .B(n8855), .Z(n8857) );
  NAND U9905 ( .A(n8858), .B(n8857), .Z(n9104) );
  NAND U9906 ( .A(n8860), .B(n8859), .Z(n8864) );
  NAND U9907 ( .A(n8862), .B(n8861), .Z(n8863) );
  NAND U9908 ( .A(n8864), .B(n8863), .Z(n9102) );
  NAND U9909 ( .A(n8866), .B(n8865), .Z(n8870) );
  ANDN U9910 ( .B(n8868), .A(n8867), .Z(n8869) );
  ANDN U9911 ( .B(n8870), .A(n8869), .Z(n9008) );
  NANDN U9912 ( .A(n8872), .B(n8871), .Z(n8876) );
  NAND U9913 ( .A(n8874), .B(n8873), .Z(n8875) );
  NAND U9914 ( .A(n8876), .B(n8875), .Z(n9007) );
  NAND U9915 ( .A(n8878), .B(n8877), .Z(n8882) );
  ANDN U9916 ( .B(n8880), .A(n8879), .Z(n8881) );
  ANDN U9917 ( .B(n8882), .A(n8881), .Z(n9022) );
  AND U9918 ( .A(x[224]), .B(y[1883]), .Z(n9090) );
  NAND U9919 ( .A(x[251]), .B(y[1856]), .Z(n9091) );
  XNOR U9920 ( .A(n9090), .B(n9091), .Z(n9092) );
  NAND U9921 ( .A(x[250]), .B(y[1857]), .Z(n9081) );
  XOR U9922 ( .A(o[91]), .B(n9081), .Z(n9093) );
  XNOR U9923 ( .A(n9092), .B(n9093), .Z(n9019) );
  AND U9924 ( .A(x[233]), .B(y[1874]), .Z(n9075) );
  NAND U9925 ( .A(x[245]), .B(y[1862]), .Z(n9076) );
  XNOR U9926 ( .A(n9075), .B(n9076), .Z(n9077) );
  NAND U9927 ( .A(x[242]), .B(y[1865]), .Z(n9078) );
  XOR U9928 ( .A(n9077), .B(n9078), .Z(n9020) );
  XOR U9929 ( .A(n9010), .B(n9009), .Z(n9103) );
  XOR U9930 ( .A(n9102), .B(n9103), .Z(n9105) );
  XOR U9931 ( .A(n9104), .B(n9105), .Z(n9123) );
  NAND U9932 ( .A(n8884), .B(n8883), .Z(n8888) );
  NAND U9933 ( .A(n8886), .B(n8885), .Z(n8887) );
  AND U9934 ( .A(n8888), .B(n8887), .Z(n9121) );
  NAND U9935 ( .A(n8890), .B(n8889), .Z(n8894) );
  NANDN U9936 ( .A(n8892), .B(n8891), .Z(n8893) );
  AND U9937 ( .A(n8894), .B(n8893), .Z(n9120) );
  XOR U9938 ( .A(n9121), .B(n9120), .Z(n9122) );
  NANDN U9939 ( .A(n8896), .B(n8895), .Z(n8900) );
  NAND U9940 ( .A(n8898), .B(n8897), .Z(n8899) );
  AND U9941 ( .A(n8900), .B(n8899), .Z(n9111) );
  NANDN U9942 ( .A(n8902), .B(n8901), .Z(n8906) );
  NANDN U9943 ( .A(n8904), .B(n8903), .Z(n8905) );
  AND U9944 ( .A(n8906), .B(n8905), .Z(n9108) );
  NAND U9945 ( .A(n8908), .B(n8907), .Z(n8912) );
  NAND U9946 ( .A(n8910), .B(n8909), .Z(n8911) );
  NAND U9947 ( .A(n8912), .B(n8911), .Z(n9098) );
  NAND U9948 ( .A(n8914), .B(n8913), .Z(n8918) );
  NAND U9949 ( .A(n8916), .B(n8915), .Z(n8917) );
  NAND U9950 ( .A(n8918), .B(n8917), .Z(n9096) );
  AND U9951 ( .A(x[243]), .B(y[1864]), .Z(n9069) );
  NAND U9952 ( .A(x[249]), .B(y[1858]), .Z(n9070) );
  XNOR U9953 ( .A(n9069), .B(n9070), .Z(n9071) );
  NAND U9954 ( .A(x[230]), .B(y[1877]), .Z(n9072) );
  XNOR U9955 ( .A(n9071), .B(n9072), .Z(n9059) );
  AND U9956 ( .A(x[239]), .B(y[1868]), .Z(n9039) );
  AND U9957 ( .A(x[226]), .B(y[1881]), .Z(n9038) );
  XOR U9958 ( .A(n9039), .B(n9038), .Z(n9041) );
  AND U9959 ( .A(x[227]), .B(y[1880]), .Z(n9040) );
  XOR U9960 ( .A(n9041), .B(n9040), .Z(n9058) );
  XOR U9961 ( .A(n9059), .B(n9058), .Z(n9060) );
  NAND U9962 ( .A(x[240]), .B(y[1867]), .Z(n9025) );
  XOR U9963 ( .A(n9025), .B(n9026), .Z(n9028) );
  XOR U9964 ( .A(n9027), .B(n9028), .Z(n9035) );
  AND U9965 ( .A(y[1870]), .B(x[237]), .Z(n8920) );
  NAND U9966 ( .A(y[1871]), .B(x[236]), .Z(n8919) );
  XNOR U9967 ( .A(n8920), .B(n8919), .Z(n9034) );
  XOR U9968 ( .A(n9035), .B(n9034), .Z(n9061) );
  NAND U9969 ( .A(n9033), .B(n8921), .Z(n8925) );
  ANDN U9970 ( .B(n8923), .A(n8922), .Z(n8924) );
  ANDN U9971 ( .B(n8925), .A(n8924), .Z(n9002) );
  NANDN U9972 ( .A(n8927), .B(n8926), .Z(n8931) );
  NAND U9973 ( .A(n8929), .B(n8928), .Z(n8930) );
  NAND U9974 ( .A(n8931), .B(n8930), .Z(n9001) );
  XOR U9975 ( .A(n9004), .B(n9003), .Z(n9097) );
  XNOR U9976 ( .A(n9096), .B(n9097), .Z(n9099) );
  XNOR U9977 ( .A(n9108), .B(n9109), .Z(n9110) );
  XOR U9978 ( .A(n9111), .B(n9110), .Z(n8983) );
  XOR U9979 ( .A(n8985), .B(n8986), .Z(n8991) );
  NANDN U9980 ( .A(n8933), .B(n8932), .Z(n8937) );
  NAND U9981 ( .A(n8935), .B(n8934), .Z(n8936) );
  AND U9982 ( .A(n8937), .B(n8936), .Z(n8990) );
  NAND U9983 ( .A(n8939), .B(n8938), .Z(n8943) );
  NAND U9984 ( .A(n8941), .B(n8940), .Z(n8942) );
  NAND U9985 ( .A(n8943), .B(n8942), .Z(n9116) );
  NANDN U9986 ( .A(n8945), .B(n8944), .Z(n8949) );
  ANDN U9987 ( .B(n8947), .A(n8946), .Z(n8948) );
  ANDN U9988 ( .B(n8949), .A(n8948), .Z(n9047) );
  NANDN U9989 ( .A(n8951), .B(n8950), .Z(n8955) );
  NANDN U9990 ( .A(n8953), .B(n8952), .Z(n8954) );
  NAND U9991 ( .A(n8955), .B(n8954), .Z(n9046) );
  AND U9992 ( .A(x[232]), .B(y[1876]), .Z(n9083) );
  NAND U9993 ( .A(n9083), .B(n8956), .Z(n8960) );
  NANDN U9994 ( .A(n8958), .B(n8957), .Z(n8959) );
  NAND U9995 ( .A(n8960), .B(n8959), .Z(n9015) );
  AND U9996 ( .A(x[238]), .B(y[1869]), .Z(n9043) );
  AND U9997 ( .A(x[225]), .B(y[1882]), .Z(n9042) );
  XOR U9998 ( .A(n9043), .B(n9042), .Z(n9045) );
  ANDN U9999 ( .B(o[90]), .A(n8961), .Z(n9044) );
  XOR U10000 ( .A(n9045), .B(n9044), .Z(n9014) );
  AND U10001 ( .A(x[241]), .B(y[1866]), .Z(n9084) );
  NAND U10002 ( .A(x[228]), .B(y[1879]), .Z(n9085) );
  XNOR U10003 ( .A(n9084), .B(n9085), .Z(n9087) );
  AND U10004 ( .A(x[229]), .B(y[1878]), .Z(n9086) );
  XOR U10005 ( .A(n9087), .B(n9086), .Z(n9013) );
  XOR U10006 ( .A(n9014), .B(n9013), .Z(n9016) );
  XOR U10007 ( .A(n9015), .B(n9016), .Z(n9048) );
  XOR U10008 ( .A(n9049), .B(n9048), .Z(n9114) );
  NANDN U10009 ( .A(n8963), .B(n8962), .Z(n8967) );
  NAND U10010 ( .A(n8965), .B(n8964), .Z(n8966) );
  AND U10011 ( .A(n8967), .B(n8966), .Z(n9055) );
  AND U10012 ( .A(y[1859]), .B(x[248]), .Z(n8969) );
  NAND U10013 ( .A(y[1863]), .B(x[244]), .Z(n8968) );
  XNOR U10014 ( .A(n8969), .B(n8968), .Z(n9065) );
  NAND U10015 ( .A(x[231]), .B(y[1876]), .Z(n9066) );
  XNOR U10016 ( .A(n9065), .B(n9066), .Z(n9053) );
  AND U10017 ( .A(x[232]), .B(y[1875]), .Z(n9030) );
  AND U10018 ( .A(x[247]), .B(y[1860]), .Z(n9029) );
  XOR U10019 ( .A(n9030), .B(n9029), .Z(n9032) );
  AND U10020 ( .A(x[246]), .B(y[1861]), .Z(n9031) );
  XOR U10021 ( .A(n9032), .B(n9031), .Z(n9052) );
  XOR U10022 ( .A(n9053), .B(n9052), .Z(n9054) );
  XNOR U10023 ( .A(n9114), .B(n9115), .Z(n9117) );
  XOR U10024 ( .A(n9116), .B(n9117), .Z(n8996) );
  NANDN U10025 ( .A(n8971), .B(n8970), .Z(n8975) );
  NANDN U10026 ( .A(n8973), .B(n8972), .Z(n8974) );
  NAND U10027 ( .A(n8975), .B(n8974), .Z(n8995) );
  NANDN U10028 ( .A(n8977), .B(n8976), .Z(n8981) );
  NANDN U10029 ( .A(n8979), .B(n8978), .Z(n8980) );
  AND U10030 ( .A(n8981), .B(n8980), .Z(n8997) );
  XOR U10031 ( .A(n8998), .B(n8997), .Z(n8989) );
  XOR U10032 ( .A(n8991), .B(n8992), .Z(n9133) );
  XOR U10033 ( .A(n9134), .B(n9133), .Z(n9135) );
  XOR U10034 ( .A(n9136), .B(n9135), .Z(n9129) );
  XNOR U10035 ( .A(n9128), .B(n9129), .Z(n8982) );
  XOR U10036 ( .A(n9126), .B(n8982), .Z(N188) );
  NANDN U10037 ( .A(n8984), .B(n8983), .Z(n8988) );
  NANDN U10038 ( .A(n8986), .B(n8985), .Z(n8987) );
  AND U10039 ( .A(n8988), .B(n8987), .Z(n9293) );
  NANDN U10040 ( .A(n8990), .B(n8989), .Z(n8994) );
  NAND U10041 ( .A(n8992), .B(n8991), .Z(n8993) );
  AND U10042 ( .A(n8994), .B(n8993), .Z(n9292) );
  NANDN U10043 ( .A(n8996), .B(n8995), .Z(n9000) );
  NAND U10044 ( .A(n8998), .B(n8997), .Z(n8999) );
  AND U10045 ( .A(n9000), .B(n8999), .Z(n9140) );
  NANDN U10046 ( .A(n9002), .B(n9001), .Z(n9006) );
  NAND U10047 ( .A(n9004), .B(n9003), .Z(n9005) );
  AND U10048 ( .A(n9006), .B(n9005), .Z(n9165) );
  NANDN U10049 ( .A(n9008), .B(n9007), .Z(n9012) );
  NAND U10050 ( .A(n9010), .B(n9009), .Z(n9011) );
  AND U10051 ( .A(n9012), .B(n9011), .Z(n9264) );
  NAND U10052 ( .A(n9014), .B(n9013), .Z(n9018) );
  NAND U10053 ( .A(n9016), .B(n9015), .Z(n9017) );
  AND U10054 ( .A(n9018), .B(n9017), .Z(n9262) );
  NANDN U10055 ( .A(n9020), .B(n9019), .Z(n9024) );
  NANDN U10056 ( .A(n9022), .B(n9021), .Z(n9023) );
  NAND U10057 ( .A(n9024), .B(n9023), .Z(n9261) );
  AND U10058 ( .A(x[231]), .B(y[1877]), .Z(n9213) );
  AND U10059 ( .A(x[236]), .B(y[1872]), .Z(n9212) );
  XOR U10060 ( .A(n9213), .B(n9212), .Z(n9215) );
  AND U10061 ( .A(x[235]), .B(y[1873]), .Z(n9214) );
  XOR U10062 ( .A(n9215), .B(n9214), .Z(n9230) );
  AND U10063 ( .A(x[239]), .B(y[1869]), .Z(n9240) );
  AND U10064 ( .A(x[251]), .B(y[1857]), .Z(n9228) );
  XOR U10065 ( .A(o[92]), .B(n9228), .Z(n9238) );
  AND U10066 ( .A(x[250]), .B(y[1858]), .Z(n9237) );
  XOR U10067 ( .A(n9238), .B(n9237), .Z(n9239) );
  XOR U10068 ( .A(n9240), .B(n9239), .Z(n9229) );
  XOR U10069 ( .A(n9230), .B(n9229), .Z(n9231) );
  XNOR U10070 ( .A(n9232), .B(n9231), .Z(n9267) );
  AND U10071 ( .A(x[241]), .B(y[1867]), .Z(n9179) );
  AND U10072 ( .A(x[246]), .B(y[1862]), .Z(n9178) );
  XOR U10073 ( .A(n9179), .B(n9178), .Z(n9181) );
  AND U10074 ( .A(x[228]), .B(y[1880]), .Z(n9180) );
  XOR U10075 ( .A(n9181), .B(n9180), .Z(n9246) );
  AND U10076 ( .A(x[230]), .B(y[1878]), .Z(n9400) );
  AND U10077 ( .A(x[243]), .B(y[1865]), .Z(n9218) );
  XOR U10078 ( .A(n9400), .B(n9218), .Z(n9221) );
  XOR U10079 ( .A(n9221), .B(n9220), .Z(n9245) );
  XOR U10080 ( .A(n9246), .B(n9245), .Z(n9248) );
  XOR U10081 ( .A(n9247), .B(n9248), .Z(n9268) );
  XOR U10082 ( .A(n9267), .B(n9268), .Z(n9270) );
  NAND U10083 ( .A(n9234), .B(n9033), .Z(n9037) );
  NANDN U10084 ( .A(n9035), .B(n9034), .Z(n9036) );
  NAND U10085 ( .A(n9037), .B(n9036), .Z(n9199) );
  XOR U10086 ( .A(n9197), .B(n9198), .Z(n9200) );
  XOR U10087 ( .A(n9199), .B(n9200), .Z(n9269) );
  XOR U10088 ( .A(n9270), .B(n9269), .Z(n9166) );
  XNOR U10089 ( .A(n9167), .B(n9166), .Z(n9161) );
  NANDN U10090 ( .A(n9047), .B(n9046), .Z(n9051) );
  NAND U10091 ( .A(n9049), .B(n9048), .Z(n9050) );
  AND U10092 ( .A(n9051), .B(n9050), .Z(n9252) );
  NAND U10093 ( .A(n9053), .B(n9052), .Z(n9057) );
  NANDN U10094 ( .A(n9055), .B(n9054), .Z(n9056) );
  AND U10095 ( .A(n9057), .B(n9056), .Z(n9250) );
  NAND U10096 ( .A(n9059), .B(n9058), .Z(n9063) );
  NANDN U10097 ( .A(n9061), .B(n9060), .Z(n9062) );
  NAND U10098 ( .A(n9063), .B(n9062), .Z(n9249) );
  AND U10099 ( .A(x[248]), .B(y[1863]), .Z(n9528) );
  AND U10100 ( .A(x[244]), .B(y[1859]), .Z(n9064) );
  NAND U10101 ( .A(n9528), .B(n9064), .Z(n9068) );
  NANDN U10102 ( .A(n9066), .B(n9065), .Z(n9067) );
  NAND U10103 ( .A(n9068), .B(n9067), .Z(n9284) );
  AND U10104 ( .A(x[249]), .B(y[1859]), .Z(n9208) );
  XOR U10105 ( .A(n9209), .B(n9208), .Z(n9207) );
  AND U10106 ( .A(x[225]), .B(y[1883]), .Z(n9205) );
  XOR U10107 ( .A(n9207), .B(n9205), .Z(n9282) );
  AND U10108 ( .A(x[240]), .B(y[1868]), .Z(n9202) );
  AND U10109 ( .A(x[248]), .B(y[1860]), .Z(n9201) );
  XOR U10110 ( .A(n9202), .B(n9201), .Z(n9204) );
  AND U10111 ( .A(x[226]), .B(y[1882]), .Z(n9203) );
  XOR U10112 ( .A(n9204), .B(n9203), .Z(n9281) );
  XOR U10113 ( .A(n9282), .B(n9281), .Z(n9283) );
  XNOR U10114 ( .A(n9284), .B(n9283), .Z(n9257) );
  NANDN U10115 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U10116 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U10117 ( .A(n9074), .B(n9073), .Z(n9280) );
  AND U10118 ( .A(x[227]), .B(y[1881]), .Z(n9233) );
  XOR U10119 ( .A(n9234), .B(n9233), .Z(n9236) );
  AND U10120 ( .A(x[247]), .B(y[1861]), .Z(n9235) );
  XOR U10121 ( .A(n9236), .B(n9235), .Z(n9278) );
  AND U10122 ( .A(x[229]), .B(y[1879]), .Z(n9225) );
  AND U10123 ( .A(x[245]), .B(y[1863]), .Z(n9224) );
  XOR U10124 ( .A(n9225), .B(n9224), .Z(n9227) );
  AND U10125 ( .A(x[244]), .B(y[1864]), .Z(n9226) );
  XOR U10126 ( .A(n9227), .B(n9226), .Z(n9277) );
  XOR U10127 ( .A(n9278), .B(n9277), .Z(n9279) );
  XNOR U10128 ( .A(n9280), .B(n9279), .Z(n9256) );
  NANDN U10129 ( .A(n9076), .B(n9075), .Z(n9080) );
  NANDN U10130 ( .A(n9078), .B(n9077), .Z(n9079) );
  NAND U10131 ( .A(n9080), .B(n9079), .Z(n9173) );
  AND U10132 ( .A(x[224]), .B(y[1884]), .Z(n9183) );
  AND U10133 ( .A(x[252]), .B(y[1856]), .Z(n9182) );
  XOR U10134 ( .A(n9183), .B(n9182), .Z(n9186) );
  ANDN U10135 ( .B(o[91]), .A(n9081), .Z(n9185) );
  XOR U10136 ( .A(n9186), .B(n9185), .Z(n9171) );
  NAND U10137 ( .A(y[1874]), .B(x[234]), .Z(n9082) );
  XNOR U10138 ( .A(n9083), .B(n9082), .Z(n9192) );
  AND U10139 ( .A(x[233]), .B(y[1875]), .Z(n9191) );
  XOR U10140 ( .A(n9192), .B(n9191), .Z(n9170) );
  XOR U10141 ( .A(n9171), .B(n9170), .Z(n9174) );
  XOR U10142 ( .A(n9173), .B(n9174), .Z(n9276) );
  NANDN U10143 ( .A(n9085), .B(n9084), .Z(n9089) );
  NAND U10144 ( .A(n9087), .B(n9086), .Z(n9088) );
  NAND U10145 ( .A(n9089), .B(n9088), .Z(n9273) );
  NANDN U10146 ( .A(n9091), .B(n9090), .Z(n9095) );
  NANDN U10147 ( .A(n9093), .B(n9092), .Z(n9094) );
  NAND U10148 ( .A(n9095), .B(n9094), .Z(n9274) );
  XOR U10149 ( .A(n9273), .B(n9274), .Z(n9275) );
  XNOR U10150 ( .A(n9276), .B(n9275), .Z(n9255) );
  XOR U10151 ( .A(n9256), .B(n9255), .Z(n9258) );
  XOR U10152 ( .A(n9257), .B(n9258), .Z(n9158) );
  XNOR U10153 ( .A(n9161), .B(n9160), .Z(n9154) );
  NAND U10154 ( .A(n9097), .B(n9096), .Z(n9101) );
  NANDN U10155 ( .A(n9099), .B(n9098), .Z(n9100) );
  NAND U10156 ( .A(n9101), .B(n9100), .Z(n9153) );
  NAND U10157 ( .A(n9103), .B(n9102), .Z(n9107) );
  NAND U10158 ( .A(n9105), .B(n9104), .Z(n9106) );
  NAND U10159 ( .A(n9107), .B(n9106), .Z(n9152) );
  XNOR U10160 ( .A(n9153), .B(n9152), .Z(n9155) );
  XNOR U10161 ( .A(n9140), .B(n9141), .Z(n9142) );
  NANDN U10162 ( .A(n9109), .B(n9108), .Z(n9113) );
  NAND U10163 ( .A(n9111), .B(n9110), .Z(n9112) );
  NAND U10164 ( .A(n9113), .B(n9112), .Z(n9148) );
  NANDN U10165 ( .A(n9115), .B(n9114), .Z(n9119) );
  NAND U10166 ( .A(n9117), .B(n9116), .Z(n9118) );
  NAND U10167 ( .A(n9119), .B(n9118), .Z(n9146) );
  NAND U10168 ( .A(n9121), .B(n9120), .Z(n9125) );
  NANDN U10169 ( .A(n9123), .B(n9122), .Z(n9124) );
  AND U10170 ( .A(n9125), .B(n9124), .Z(n9147) );
  XNOR U10171 ( .A(n9146), .B(n9147), .Z(n9149) );
  XNOR U10172 ( .A(n9142), .B(n9143), .Z(n9294) );
  XNOR U10173 ( .A(n9295), .B(n9294), .Z(n9288) );
  OR U10174 ( .A(n9128), .B(n9126), .Z(n9132) );
  ANDN U10175 ( .B(n9128), .A(n9127), .Z(n9130) );
  OR U10176 ( .A(n9130), .B(n9129), .Z(n9131) );
  AND U10177 ( .A(n9132), .B(n9131), .Z(n9287) );
  NAND U10178 ( .A(n9134), .B(n9133), .Z(n9138) );
  NAND U10179 ( .A(n9136), .B(n9135), .Z(n9137) );
  AND U10180 ( .A(n9138), .B(n9137), .Z(n9286) );
  IV U10181 ( .A(n9286), .Z(n9285) );
  XOR U10182 ( .A(n9287), .B(n9285), .Z(n9139) );
  XNOR U10183 ( .A(n9288), .B(n9139), .Z(N189) );
  NANDN U10184 ( .A(n9141), .B(n9140), .Z(n9145) );
  NANDN U10185 ( .A(n9143), .B(n9142), .Z(n9144) );
  NAND U10186 ( .A(n9145), .B(n9144), .Z(n9308) );
  NAND U10187 ( .A(n9147), .B(n9146), .Z(n9151) );
  NANDN U10188 ( .A(n9149), .B(n9148), .Z(n9150) );
  NAND U10189 ( .A(n9151), .B(n9150), .Z(n9306) );
  NAND U10190 ( .A(n9153), .B(n9152), .Z(n9157) );
  NANDN U10191 ( .A(n9155), .B(n9154), .Z(n9156) );
  NAND U10192 ( .A(n9157), .B(n9156), .Z(n9312) );
  NANDN U10193 ( .A(n9159), .B(n9158), .Z(n9163) );
  NAND U10194 ( .A(n9161), .B(n9160), .Z(n9162) );
  AND U10195 ( .A(n9163), .B(n9162), .Z(n9313) );
  XOR U10196 ( .A(n9312), .B(n9313), .Z(n9315) );
  NANDN U10197 ( .A(n9165), .B(n9164), .Z(n9169) );
  NAND U10198 ( .A(n9167), .B(n9166), .Z(n9168) );
  AND U10199 ( .A(n9169), .B(n9168), .Z(n9331) );
  IV U10200 ( .A(n9170), .Z(n9172) );
  NANDN U10201 ( .A(n9172), .B(n9171), .Z(n9177) );
  IV U10202 ( .A(n9173), .Z(n9175) );
  NANDN U10203 ( .A(n9175), .B(n9174), .Z(n9176) );
  AND U10204 ( .A(n9177), .B(n9176), .Z(n9428) );
  IV U10205 ( .A(n9182), .Z(n9184) );
  NANDN U10206 ( .A(n9184), .B(n9183), .Z(n9189) );
  IV U10207 ( .A(n9185), .Z(n9187) );
  NANDN U10208 ( .A(n9187), .B(n9186), .Z(n9188) );
  NAND U10209 ( .A(n9189), .B(n9188), .Z(n9462) );
  XOR U10210 ( .A(n9461), .B(n9462), .Z(n9463) );
  AND U10211 ( .A(x[234]), .B(y[1876]), .Z(n9459) );
  NAND U10212 ( .A(n9190), .B(n9459), .Z(n9194) );
  NAND U10213 ( .A(n9192), .B(n9191), .Z(n9193) );
  NAND U10214 ( .A(n9194), .B(n9193), .Z(n9433) );
  AND U10215 ( .A(x[246]), .B(y[1863]), .Z(n9380) );
  AND U10216 ( .A(x[236]), .B(y[1873]), .Z(n9646) );
  AND U10217 ( .A(x[225]), .B(y[1884]), .Z(n9378) );
  XOR U10218 ( .A(n9646), .B(n9378), .Z(n9379) );
  XOR U10219 ( .A(n9380), .B(n9379), .Z(n9432) );
  AND U10220 ( .A(x[239]), .B(y[1870]), .Z(n9381) );
  XOR U10221 ( .A(n9381), .B(n9195), .Z(n9382) );
  XOR U10222 ( .A(n9382), .B(n9196), .Z(n9431) );
  XOR U10223 ( .A(n9432), .B(n9431), .Z(n9434) );
  XNOR U10224 ( .A(n9433), .B(n9434), .Z(n9464) );
  XOR U10225 ( .A(n9463), .B(n9464), .Z(n9427) );
  XOR U10226 ( .A(n9428), .B(n9427), .Z(n9430) );
  XOR U10227 ( .A(n9430), .B(n9429), .Z(n9426) );
  IV U10228 ( .A(n9205), .Z(n9206) );
  ANDN U10229 ( .B(n9207), .A(n9206), .Z(n9211) );
  NAND U10230 ( .A(n9209), .B(n9208), .Z(n9210) );
  NANDN U10231 ( .A(n9211), .B(n9210), .Z(n9437) );
  XOR U10232 ( .A(n9438), .B(n9437), .Z(n9439) );
  NAND U10233 ( .A(n9213), .B(n9212), .Z(n9217) );
  NAND U10234 ( .A(n9215), .B(n9214), .Z(n9216) );
  NAND U10235 ( .A(n9217), .B(n9216), .Z(n9344) );
  AND U10236 ( .A(x[235]), .B(y[1874]), .Z(n9397) );
  AND U10237 ( .A(x[227]), .B(y[1882]), .Z(n9395) );
  AND U10238 ( .A(x[241]), .B(y[1868]), .Z(n9394) );
  XOR U10239 ( .A(n9395), .B(n9394), .Z(n9396) );
  XOR U10240 ( .A(n9397), .B(n9396), .Z(n9343) );
  AND U10241 ( .A(x[247]), .B(y[1862]), .Z(n9391) );
  AND U10242 ( .A(x[237]), .B(y[1872]), .Z(n9389) );
  AND U10243 ( .A(x[248]), .B(y[1861]), .Z(n9511) );
  XOR U10244 ( .A(n9389), .B(n9511), .Z(n9390) );
  XOR U10245 ( .A(n9391), .B(n9390), .Z(n9342) );
  XOR U10246 ( .A(n9343), .B(n9342), .Z(n9345) );
  XNOR U10247 ( .A(n9344), .B(n9345), .Z(n9440) );
  IV U10248 ( .A(n9218), .Z(n9219) );
  NANDN U10249 ( .A(n9219), .B(n9400), .Z(n9223) );
  NAND U10250 ( .A(n9221), .B(n9220), .Z(n9222) );
  NAND U10251 ( .A(n9223), .B(n9222), .Z(n9446) );
  AND U10252 ( .A(x[249]), .B(y[1860]), .Z(n9375) );
  AND U10253 ( .A(x[250]), .B(y[1859]), .Z(n9372) );
  XOR U10254 ( .A(n9373), .B(n9372), .Z(n9374) );
  XOR U10255 ( .A(n9375), .B(n9374), .Z(n9444) );
  AND U10256 ( .A(x[252]), .B(y[1857]), .Z(n9388) );
  XOR U10257 ( .A(o[93]), .B(n9388), .Z(n9454) );
  AND U10258 ( .A(x[224]), .B(y[1885]), .Z(n9452) );
  AND U10259 ( .A(x[253]), .B(y[1856]), .Z(n9451) );
  XOR U10260 ( .A(n9452), .B(n9451), .Z(n9453) );
  XNOR U10261 ( .A(n9454), .B(n9453), .Z(n9443) );
  XOR U10262 ( .A(n9446), .B(n9445), .Z(n9417) );
  AND U10263 ( .A(n9228), .B(o[92]), .Z(n9351) );
  AND U10264 ( .A(x[240]), .B(y[1869]), .Z(n9349) );
  AND U10265 ( .A(x[251]), .B(y[1858]), .Z(n9348) );
  XOR U10266 ( .A(n9349), .B(n9348), .Z(n9350) );
  XOR U10267 ( .A(n9351), .B(n9350), .Z(n9408) );
  AND U10268 ( .A(x[226]), .B(y[1883]), .Z(n9361) );
  XOR U10269 ( .A(n9361), .B(n9360), .Z(n9362) );
  XOR U10270 ( .A(n9363), .B(n9362), .Z(n9407) );
  XOR U10271 ( .A(n9408), .B(n9407), .Z(n9410) );
  XOR U10272 ( .A(n9409), .B(n9410), .Z(n9418) );
  NAND U10273 ( .A(n9238), .B(n9237), .Z(n9242) );
  NAND U10274 ( .A(n9240), .B(n9239), .Z(n9241) );
  NAND U10275 ( .A(n9242), .B(n9241), .Z(n9366) );
  XOR U10276 ( .A(n9367), .B(n9366), .Z(n9368) );
  AND U10277 ( .A(x[232]), .B(y[1877]), .Z(n9402) );
  AND U10278 ( .A(y[1879]), .B(x[230]), .Z(n9244) );
  NAND U10279 ( .A(y[1878]), .B(x[231]), .Z(n9243) );
  XNOR U10280 ( .A(n9244), .B(n9243), .Z(n9401) );
  XNOR U10281 ( .A(n9402), .B(n9401), .Z(n9449) );
  AND U10282 ( .A(x[229]), .B(y[1880]), .Z(n9357) );
  AND U10283 ( .A(x[228]), .B(y[1881]), .Z(n9355) );
  AND U10284 ( .A(x[234]), .B(y[1875]), .Z(n9354) );
  XOR U10285 ( .A(n9355), .B(n9354), .Z(n9356) );
  XOR U10286 ( .A(n9357), .B(n9356), .Z(n9450) );
  AND U10287 ( .A(x[233]), .B(y[1876]), .Z(n9564) );
  XOR U10288 ( .A(n9368), .B(n9369), .Z(n9337) );
  XOR U10289 ( .A(n9336), .B(n9337), .Z(n9339) );
  XOR U10290 ( .A(n9338), .B(n9339), .Z(n9423) );
  XOR U10291 ( .A(n9423), .B(n9424), .Z(n9425) );
  XNOR U10292 ( .A(n9426), .B(n9425), .Z(n9330) );
  NANDN U10293 ( .A(n9250), .B(n9249), .Z(n9254) );
  NANDN U10294 ( .A(n9252), .B(n9251), .Z(n9253) );
  AND U10295 ( .A(n9254), .B(n9253), .Z(n9325) );
  NAND U10296 ( .A(n9256), .B(n9255), .Z(n9260) );
  NAND U10297 ( .A(n9258), .B(n9257), .Z(n9259) );
  AND U10298 ( .A(n9260), .B(n9259), .Z(n9324) );
  NANDN U10299 ( .A(n9262), .B(n9261), .Z(n9266) );
  NANDN U10300 ( .A(n9264), .B(n9263), .Z(n9265) );
  NAND U10301 ( .A(n9266), .B(n9265), .Z(n9320) );
  NAND U10302 ( .A(n9268), .B(n9267), .Z(n9272) );
  NAND U10303 ( .A(n9270), .B(n9269), .Z(n9271) );
  NAND U10304 ( .A(n9272), .B(n9271), .Z(n9318) );
  XOR U10305 ( .A(n9413), .B(n9414), .Z(n9416) );
  XOR U10306 ( .A(n9415), .B(n9416), .Z(n9319) );
  XOR U10307 ( .A(n9318), .B(n9319), .Z(n9321) );
  XOR U10308 ( .A(n9320), .B(n9321), .Z(n9326) );
  XOR U10309 ( .A(n9327), .B(n9326), .Z(n9332) );
  XOR U10310 ( .A(n9333), .B(n9332), .Z(n9314) );
  XOR U10311 ( .A(n9315), .B(n9314), .Z(n9307) );
  XNOR U10312 ( .A(n9306), .B(n9307), .Z(n9309) );
  XOR U10313 ( .A(n9308), .B(n9309), .Z(n9302) );
  OR U10314 ( .A(n9287), .B(n9285), .Z(n9291) );
  ANDN U10315 ( .B(n9287), .A(n9286), .Z(n9289) );
  OR U10316 ( .A(n9289), .B(n9288), .Z(n9290) );
  AND U10317 ( .A(n9291), .B(n9290), .Z(n9301) );
  NANDN U10318 ( .A(n9293), .B(n9292), .Z(n9297) );
  NAND U10319 ( .A(n9295), .B(n9294), .Z(n9296) );
  NAND U10320 ( .A(n9297), .B(n9296), .Z(n9300) );
  IV U10321 ( .A(n9300), .Z(n9299) );
  XOR U10322 ( .A(n9301), .B(n9299), .Z(n9298) );
  XNOR U10323 ( .A(n9302), .B(n9298), .Z(N190) );
  OR U10324 ( .A(n9301), .B(n9299), .Z(n9305) );
  ANDN U10325 ( .B(n9301), .A(n9300), .Z(n9303) );
  OR U10326 ( .A(n9303), .B(n9302), .Z(n9304) );
  AND U10327 ( .A(n9305), .B(n9304), .Z(n9717) );
  NAND U10328 ( .A(n9307), .B(n9306), .Z(n9311) );
  NANDN U10329 ( .A(n9309), .B(n9308), .Z(n9310) );
  NAND U10330 ( .A(n9311), .B(n9310), .Z(n9718) );
  NAND U10331 ( .A(n9313), .B(n9312), .Z(n9317) );
  NAND U10332 ( .A(n9315), .B(n9314), .Z(n9316) );
  NAND U10333 ( .A(n9317), .B(n9316), .Z(n9721) );
  NAND U10334 ( .A(n9319), .B(n9318), .Z(n9323) );
  NAND U10335 ( .A(n9321), .B(n9320), .Z(n9322) );
  AND U10336 ( .A(n9323), .B(n9322), .Z(n9728) );
  NANDN U10337 ( .A(n9325), .B(n9324), .Z(n9329) );
  NAND U10338 ( .A(n9327), .B(n9326), .Z(n9328) );
  AND U10339 ( .A(n9329), .B(n9328), .Z(n9729) );
  NANDN U10340 ( .A(n9331), .B(n9330), .Z(n9335) );
  NAND U10341 ( .A(n9333), .B(n9332), .Z(n9334) );
  NAND U10342 ( .A(n9335), .B(n9334), .Z(n9730) );
  XOR U10343 ( .A(n9728), .B(n9727), .Z(n9724) );
  NANDN U10344 ( .A(n9337), .B(n9336), .Z(n9341) );
  NANDN U10345 ( .A(n9339), .B(n9338), .Z(n9340) );
  AND U10346 ( .A(n9341), .B(n9340), .Z(n9466) );
  NAND U10347 ( .A(n9343), .B(n9342), .Z(n9347) );
  NAND U10348 ( .A(n9345), .B(n9344), .Z(n9346) );
  AND U10349 ( .A(n9347), .B(n9346), .Z(n9472) );
  NAND U10350 ( .A(n9349), .B(n9348), .Z(n9353) );
  NAND U10351 ( .A(n9351), .B(n9350), .Z(n9352) );
  NAND U10352 ( .A(n9353), .B(n9352), .Z(n9479) );
  NAND U10353 ( .A(n9355), .B(n9354), .Z(n9359) );
  NAND U10354 ( .A(n9357), .B(n9356), .Z(n9358) );
  NAND U10355 ( .A(n9359), .B(n9358), .Z(n9482) );
  AND U10356 ( .A(x[230]), .B(y[1880]), .Z(n9515) );
  AND U10357 ( .A(x[229]), .B(y[1881]), .Z(n9517) );
  AND U10358 ( .A(x[243]), .B(y[1867]), .Z(n9516) );
  XOR U10359 ( .A(n9517), .B(n9516), .Z(n9514) );
  XNOR U10360 ( .A(n9515), .B(n9514), .Z(n9483) );
  AND U10361 ( .A(x[228]), .B(y[1882]), .Z(n9630) );
  AND U10362 ( .A(x[227]), .B(y[1883]), .Z(n9632) );
  AND U10363 ( .A(x[242]), .B(y[1868]), .Z(n9631) );
  XOR U10364 ( .A(n9632), .B(n9631), .Z(n9629) );
  XOR U10365 ( .A(n9630), .B(n9629), .Z(n9486) );
  NAND U10366 ( .A(n9361), .B(n9360), .Z(n9365) );
  NAND U10367 ( .A(n9363), .B(n9362), .Z(n9364) );
  AND U10368 ( .A(n9365), .B(n9364), .Z(n9485) );
  XOR U10369 ( .A(n9483), .B(n9484), .Z(n9481) );
  XOR U10370 ( .A(n9482), .B(n9481), .Z(n9480) );
  XOR U10371 ( .A(n9479), .B(n9480), .Z(n9471) );
  NAND U10372 ( .A(n9367), .B(n9366), .Z(n9371) );
  NAND U10373 ( .A(n9369), .B(n9368), .Z(n9370) );
  AND U10374 ( .A(n9371), .B(n9370), .Z(n9469) );
  XOR U10375 ( .A(n9470), .B(n9469), .Z(n9468) );
  AND U10376 ( .A(n9373), .B(n9372), .Z(n9377) );
  NAND U10377 ( .A(n9375), .B(n9374), .Z(n9376) );
  NANDN U10378 ( .A(n9377), .B(n9376), .Z(n9503) );
  NANDN U10379 ( .A(n9626), .B(n9381), .Z(n9385) );
  NANDN U10380 ( .A(n9383), .B(n9382), .Z(n9384) );
  AND U10381 ( .A(n9385), .B(n9384), .Z(n9666) );
  AND U10382 ( .A(x[247]), .B(y[1863]), .Z(n9510) );
  AND U10383 ( .A(y[1862]), .B(x[248]), .Z(n9387) );
  AND U10384 ( .A(y[1861]), .B(x[249]), .Z(n9386) );
  XOR U10385 ( .A(n9387), .B(n9386), .Z(n9509) );
  XOR U10386 ( .A(n9510), .B(n9509), .Z(n9668) );
  AND U10387 ( .A(n9388), .B(o[93]), .Z(n9594) );
  AND U10388 ( .A(x[252]), .B(y[1858]), .Z(n9596) );
  AND U10389 ( .A(x[240]), .B(y[1870]), .Z(n9595) );
  XOR U10390 ( .A(n9596), .B(n9595), .Z(n9593) );
  XNOR U10391 ( .A(n9594), .B(n9593), .Z(n9667) );
  XNOR U10392 ( .A(n9666), .B(n9665), .Z(n9505) );
  XOR U10393 ( .A(n9506), .B(n9505), .Z(n9504) );
  XOR U10394 ( .A(n9503), .B(n9504), .Z(n9696) );
  NAND U10395 ( .A(n9389), .B(n9511), .Z(n9393) );
  NAND U10396 ( .A(n9391), .B(n9390), .Z(n9392) );
  NAND U10397 ( .A(n9393), .B(n9392), .Z(n9476) );
  NAND U10398 ( .A(n9395), .B(n9394), .Z(n9399) );
  NAND U10399 ( .A(n9397), .B(n9396), .Z(n9398) );
  AND U10400 ( .A(n9399), .B(n9398), .Z(n9660) );
  AND U10401 ( .A(x[224]), .B(y[1886]), .Z(n9568) );
  AND U10402 ( .A(x[253]), .B(y[1857]), .Z(n9547) );
  XOR U10403 ( .A(o[94]), .B(n9547), .Z(n9570) );
  AND U10404 ( .A(x[254]), .B(y[1856]), .Z(n9569) );
  XOR U10405 ( .A(n9570), .B(n9569), .Z(n9567) );
  XOR U10406 ( .A(n9568), .B(n9567), .Z(n9662) );
  AND U10407 ( .A(x[244]), .B(y[1866]), .Z(n9605) );
  XOR U10408 ( .A(n9606), .B(n9605), .Z(n9604) );
  AND U10409 ( .A(x[232]), .B(y[1878]), .Z(n9603) );
  XNOR U10410 ( .A(n9604), .B(n9603), .Z(n9661) );
  XNOR U10411 ( .A(n9660), .B(n9659), .Z(n9475) );
  XOR U10412 ( .A(n9476), .B(n9475), .Z(n9473) );
  AND U10413 ( .A(x[231]), .B(y[1879]), .Z(n9624) );
  NAND U10414 ( .A(n9400), .B(n9624), .Z(n9404) );
  NAND U10415 ( .A(n9402), .B(n9401), .Z(n9403) );
  AND U10416 ( .A(n9404), .B(n9403), .Z(n9495) );
  AND U10417 ( .A(y[1865]), .B(x[245]), .Z(n9406) );
  AND U10418 ( .A(y[1864]), .B(x[246]), .Z(n9405) );
  XOR U10419 ( .A(n9406), .B(n9405), .Z(n9623) );
  XOR U10420 ( .A(n9624), .B(n9623), .Z(n9498) );
  AND U10421 ( .A(x[241]), .B(y[1869]), .Z(n9588) );
  AND U10422 ( .A(x[226]), .B(y[1884]), .Z(n9590) );
  AND U10423 ( .A(x[250]), .B(y[1860]), .Z(n9589) );
  XOR U10424 ( .A(n9590), .B(n9589), .Z(n9587) );
  XNOR U10425 ( .A(n9588), .B(n9587), .Z(n9497) );
  XNOR U10426 ( .A(n9495), .B(n9496), .Z(n9474) );
  NAND U10427 ( .A(n9408), .B(n9407), .Z(n9412) );
  NAND U10428 ( .A(n9410), .B(n9409), .Z(n9411) );
  NAND U10429 ( .A(n9412), .B(n9411), .Z(n9697) );
  XOR U10430 ( .A(n9698), .B(n9697), .Z(n9695) );
  XOR U10431 ( .A(n9696), .B(n9695), .Z(n9467) );
  XOR U10432 ( .A(n9466), .B(n9465), .Z(n9708) );
  NANDN U10433 ( .A(n9418), .B(n9417), .Z(n9422) );
  NANDN U10434 ( .A(n9420), .B(n9419), .Z(n9421) );
  NAND U10435 ( .A(n9422), .B(n9421), .Z(n9709) );
  XOR U10436 ( .A(n9710), .B(n9709), .Z(n9707) );
  NAND U10437 ( .A(n9432), .B(n9431), .Z(n9436) );
  NAND U10438 ( .A(n9434), .B(n9433), .Z(n9435) );
  AND U10439 ( .A(n9436), .B(n9435), .Z(n9687) );
  NAND U10440 ( .A(n9438), .B(n9437), .Z(n9442) );
  NANDN U10441 ( .A(n9440), .B(n9439), .Z(n9441) );
  NAND U10442 ( .A(n9442), .B(n9441), .Z(n9688) );
  NANDN U10443 ( .A(n9444), .B(n9443), .Z(n9448) );
  OR U10444 ( .A(n9446), .B(n9445), .Z(n9447) );
  NAND U10445 ( .A(n9448), .B(n9447), .Z(n9685) );
  XOR U10446 ( .A(n9686), .B(n9685), .Z(n9694) );
  NAND U10447 ( .A(n9452), .B(n9451), .Z(n9456) );
  NAND U10448 ( .A(n9454), .B(n9453), .Z(n9455) );
  AND U10449 ( .A(n9456), .B(n9455), .Z(n9490) );
  AND U10450 ( .A(y[1874]), .B(x[236]), .Z(n9457) );
  XOR U10451 ( .A(n9458), .B(n9457), .Z(n9643) );
  XOR U10452 ( .A(n9644), .B(n9643), .Z(n9562) );
  AND U10453 ( .A(y[1877]), .B(x[233]), .Z(n9460) );
  XOR U10454 ( .A(n9460), .B(n9459), .Z(n9561) );
  XOR U10455 ( .A(n9562), .B(n9561), .Z(n9492) );
  AND U10456 ( .A(x[251]), .B(y[1859]), .Z(n9640) );
  AND U10457 ( .A(x[225]), .B(y[1885]), .Z(n9639) );
  XOR U10458 ( .A(n9640), .B(n9639), .Z(n9637) );
  XOR U10459 ( .A(n9638), .B(n9637), .Z(n9491) );
  XOR U10460 ( .A(n9492), .B(n9491), .Z(n9489) );
  XOR U10461 ( .A(n9490), .B(n9489), .Z(n9681) );
  XOR U10462 ( .A(n9682), .B(n9681), .Z(n9680) );
  XNOR U10463 ( .A(n9680), .B(n9679), .Z(n9693) );
  XOR U10464 ( .A(n9692), .B(n9691), .Z(n9703) );
  XOR U10465 ( .A(n9702), .B(n9701), .Z(n9723) );
  XOR U10466 ( .A(n9721), .B(n9722), .Z(n9715) );
  XNOR U10467 ( .A(n9716), .B(n9715), .Z(N191) );
  NANDN U10468 ( .A(n9474), .B(n9473), .Z(n9478) );
  NAND U10469 ( .A(n9476), .B(n9475), .Z(n9477) );
  AND U10470 ( .A(n9478), .B(n9477), .Z(n9700) );
  NANDN U10471 ( .A(n9484), .B(n9483), .Z(n9488) );
  NANDN U10472 ( .A(n9486), .B(n9485), .Z(n9487) );
  NANDN U10473 ( .A(n9490), .B(n9489), .Z(n9494) );
  NAND U10474 ( .A(n9492), .B(n9491), .Z(n9493) );
  AND U10475 ( .A(n9494), .B(n9493), .Z(n9502) );
  NANDN U10476 ( .A(n9496), .B(n9495), .Z(n9500) );
  NANDN U10477 ( .A(n9498), .B(n9497), .Z(n9499) );
  NAND U10478 ( .A(n9500), .B(n9499), .Z(n9501) );
  XNOR U10479 ( .A(n9502), .B(n9501), .Z(n9678) );
  NAND U10480 ( .A(n9504), .B(n9503), .Z(n9508) );
  NAND U10481 ( .A(n9506), .B(n9505), .Z(n9507) );
  AND U10482 ( .A(n9508), .B(n9507), .Z(n9676) );
  NAND U10483 ( .A(n9510), .B(n9509), .Z(n9513) );
  AND U10484 ( .A(x[249]), .B(y[1862]), .Z(n9548) );
  NAND U10485 ( .A(n9511), .B(n9548), .Z(n9512) );
  AND U10486 ( .A(n9513), .B(n9512), .Z(n9521) );
  NAND U10487 ( .A(n9515), .B(n9514), .Z(n9519) );
  NAND U10488 ( .A(n9517), .B(n9516), .Z(n9518) );
  NAND U10489 ( .A(n9519), .B(n9518), .Z(n9520) );
  XNOR U10490 ( .A(n9521), .B(n9520), .Z(n9586) );
  AND U10491 ( .A(y[1871]), .B(x[240]), .Z(n9523) );
  NAND U10492 ( .A(y[1867]), .B(x[244]), .Z(n9522) );
  XNOR U10493 ( .A(n9523), .B(n9522), .Z(n9527) );
  AND U10494 ( .A(y[1876]), .B(x[235]), .Z(n9525) );
  NAND U10495 ( .A(y[1861]), .B(x[250]), .Z(n9524) );
  XNOR U10496 ( .A(n9525), .B(n9524), .Z(n9526) );
  XOR U10497 ( .A(n9527), .B(n9526), .Z(n9530) );
  AND U10498 ( .A(x[246]), .B(y[1865]), .Z(n9625) );
  XNOR U10499 ( .A(n9528), .B(n9625), .Z(n9529) );
  XNOR U10500 ( .A(n9530), .B(n9529), .Z(n9546) );
  AND U10501 ( .A(y[1880]), .B(x[231]), .Z(n9532) );
  NAND U10502 ( .A(y[1884]), .B(x[227]), .Z(n9531) );
  XNOR U10503 ( .A(n9532), .B(n9531), .Z(n9536) );
  AND U10504 ( .A(y[1882]), .B(x[229]), .Z(n9534) );
  NAND U10505 ( .A(y[1881]), .B(x[230]), .Z(n9533) );
  XNOR U10506 ( .A(n9534), .B(n9533), .Z(n9535) );
  XOR U10507 ( .A(n9536), .B(n9535), .Z(n9544) );
  AND U10508 ( .A(y[1864]), .B(x[247]), .Z(n9538) );
  NAND U10509 ( .A(y[1875]), .B(x[236]), .Z(n9537) );
  XNOR U10510 ( .A(n9538), .B(n9537), .Z(n9542) );
  AND U10511 ( .A(y[1860]), .B(x[251]), .Z(n9540) );
  NAND U10512 ( .A(y[1869]), .B(x[242]), .Z(n9539) );
  XNOR U10513 ( .A(n9540), .B(n9539), .Z(n9541) );
  XNOR U10514 ( .A(n9542), .B(n9541), .Z(n9543) );
  XNOR U10515 ( .A(n9544), .B(n9543), .Z(n9545) );
  XOR U10516 ( .A(n9546), .B(n9545), .Z(n9560) );
  AND U10517 ( .A(y[1878]), .B(x[233]), .Z(n9554) );
  AND U10518 ( .A(n9547), .B(o[94]), .Z(n9552) );
  AND U10519 ( .A(x[234]), .B(y[1877]), .Z(n9563) );
  XOR U10520 ( .A(n9563), .B(o[95]), .Z(n9550) );
  XNOR U10521 ( .A(n9548), .B(n9645), .Z(n9549) );
  XNOR U10522 ( .A(n9550), .B(n9549), .Z(n9551) );
  XNOR U10523 ( .A(n9552), .B(n9551), .Z(n9553) );
  XNOR U10524 ( .A(n9554), .B(n9553), .Z(n9558) );
  AND U10525 ( .A(y[1857]), .B(x[254]), .Z(n9556) );
  NAND U10526 ( .A(y[1858]), .B(x[253]), .Z(n9555) );
  XNOR U10527 ( .A(n9556), .B(n9555), .Z(n9557) );
  XNOR U10528 ( .A(n9558), .B(n9557), .Z(n9559) );
  XNOR U10529 ( .A(n9560), .B(n9559), .Z(n9576) );
  NAND U10530 ( .A(n9562), .B(n9561), .Z(n9566) );
  NAND U10531 ( .A(n9564), .B(n9563), .Z(n9565) );
  AND U10532 ( .A(n9566), .B(n9565), .Z(n9574) );
  NAND U10533 ( .A(n9568), .B(n9567), .Z(n9572) );
  NAND U10534 ( .A(n9570), .B(n9569), .Z(n9571) );
  NAND U10535 ( .A(n9572), .B(n9571), .Z(n9573) );
  XNOR U10536 ( .A(n9574), .B(n9573), .Z(n9575) );
  XOR U10537 ( .A(n9576), .B(n9575), .Z(n9584) );
  AND U10538 ( .A(y[1873]), .B(x[238]), .Z(n9578) );
  NAND U10539 ( .A(y[1887]), .B(x[224]), .Z(n9577) );
  XNOR U10540 ( .A(n9578), .B(n9577), .Z(n9582) );
  AND U10541 ( .A(y[1886]), .B(x[225]), .Z(n9580) );
  NAND U10542 ( .A(y[1859]), .B(x[252]), .Z(n9579) );
  XNOR U10543 ( .A(n9580), .B(n9579), .Z(n9581) );
  XNOR U10544 ( .A(n9582), .B(n9581), .Z(n9583) );
  XNOR U10545 ( .A(n9584), .B(n9583), .Z(n9585) );
  XOR U10546 ( .A(n9586), .B(n9585), .Z(n9658) );
  NAND U10547 ( .A(n9588), .B(n9587), .Z(n9592) );
  NAND U10548 ( .A(n9590), .B(n9589), .Z(n9591) );
  AND U10549 ( .A(n9592), .B(n9591), .Z(n9600) );
  NAND U10550 ( .A(n9594), .B(n9593), .Z(n9598) );
  NAND U10551 ( .A(n9596), .B(n9595), .Z(n9597) );
  NAND U10552 ( .A(n9598), .B(n9597), .Z(n9599) );
  XNOR U10553 ( .A(n9600), .B(n9599), .Z(n9656) );
  AND U10554 ( .A(y[1866]), .B(x[245]), .Z(n9602) );
  NAND U10555 ( .A(y[1879]), .B(x[232]), .Z(n9601) );
  XNOR U10556 ( .A(n9602), .B(n9601), .Z(n9622) );
  AND U10557 ( .A(y[1868]), .B(x[243]), .Z(n9620) );
  NAND U10558 ( .A(n9604), .B(n9603), .Z(n9608) );
  NAND U10559 ( .A(n9606), .B(n9605), .Z(n9607) );
  AND U10560 ( .A(n9608), .B(n9607), .Z(n9616) );
  AND U10561 ( .A(y[1885]), .B(x[226]), .Z(n9610) );
  NAND U10562 ( .A(y[1870]), .B(x[241]), .Z(n9609) );
  XNOR U10563 ( .A(n9610), .B(n9609), .Z(n9614) );
  AND U10564 ( .A(y[1856]), .B(x[255]), .Z(n9612) );
  NAND U10565 ( .A(y[1883]), .B(x[228]), .Z(n9611) );
  XNOR U10566 ( .A(n9612), .B(n9611), .Z(n9613) );
  XNOR U10567 ( .A(n9614), .B(n9613), .Z(n9615) );
  XNOR U10568 ( .A(n9616), .B(n9615), .Z(n9617) );
  XNOR U10569 ( .A(n9618), .B(n9617), .Z(n9619) );
  XNOR U10570 ( .A(n9620), .B(n9619), .Z(n9621) );
  XOR U10571 ( .A(n9622), .B(n9621), .Z(n9654) );
  NAND U10572 ( .A(n9624), .B(n9623), .Z(n9628) );
  NANDN U10573 ( .A(n9626), .B(n9625), .Z(n9627) );
  AND U10574 ( .A(n9628), .B(n9627), .Z(n9636) );
  NAND U10575 ( .A(n9630), .B(n9629), .Z(n9634) );
  NAND U10576 ( .A(n9632), .B(n9631), .Z(n9633) );
  NAND U10577 ( .A(n9634), .B(n9633), .Z(n9635) );
  XNOR U10578 ( .A(n9636), .B(n9635), .Z(n9652) );
  NAND U10579 ( .A(n9638), .B(n9637), .Z(n9642) );
  NAND U10580 ( .A(n9640), .B(n9639), .Z(n9641) );
  AND U10581 ( .A(n9642), .B(n9641), .Z(n9650) );
  NAND U10582 ( .A(n9644), .B(n9643), .Z(n9648) );
  NAND U10583 ( .A(n9646), .B(n9645), .Z(n9647) );
  NAND U10584 ( .A(n9648), .B(n9647), .Z(n9649) );
  XNOR U10585 ( .A(n9650), .B(n9649), .Z(n9651) );
  XNOR U10586 ( .A(n9652), .B(n9651), .Z(n9653) );
  XNOR U10587 ( .A(n9654), .B(n9653), .Z(n9655) );
  XNOR U10588 ( .A(n9656), .B(n9655), .Z(n9657) );
  XNOR U10589 ( .A(n9658), .B(n9657), .Z(n9674) );
  NAND U10590 ( .A(n9660), .B(n9659), .Z(n9664) );
  NANDN U10591 ( .A(n9662), .B(n9661), .Z(n9663) );
  AND U10592 ( .A(n9664), .B(n9663), .Z(n9672) );
  NAND U10593 ( .A(n9666), .B(n9665), .Z(n9670) );
  NANDN U10594 ( .A(n9668), .B(n9667), .Z(n9669) );
  NAND U10595 ( .A(n9670), .B(n9669), .Z(n9671) );
  XNOR U10596 ( .A(n9672), .B(n9671), .Z(n9673) );
  XNOR U10597 ( .A(n9674), .B(n9673), .Z(n9675) );
  XNOR U10598 ( .A(n9676), .B(n9675), .Z(n9677) );
  NAND U10599 ( .A(n9680), .B(n9679), .Z(n9684) );
  NAND U10600 ( .A(n9682), .B(n9681), .Z(n9683) );
  NAND U10601 ( .A(n9686), .B(n9685), .Z(n9690) );
  NANDN U10602 ( .A(n9688), .B(n9687), .Z(n9689) );
  NAND U10603 ( .A(n9702), .B(n9701), .Z(n9706) );
  NANDN U10604 ( .A(n9704), .B(n9703), .Z(n9705) );
  AND U10605 ( .A(n9706), .B(n9705), .Z(n9714) );
  NANDN U10606 ( .A(n9708), .B(n9707), .Z(n9712) );
  NAND U10607 ( .A(n9710), .B(n9709), .Z(n9711) );
  NAND U10608 ( .A(n9712), .B(n9711), .Z(n9713) );
  NAND U10609 ( .A(n9716), .B(n9715), .Z(n9720) );
  NANDN U10610 ( .A(n9718), .B(n9717), .Z(n9719) );
  NANDN U10611 ( .A(n9722), .B(n9721), .Z(n9726) );
  NANDN U10612 ( .A(n9724), .B(n9723), .Z(n9725) );
  AND U10613 ( .A(x[224]), .B(y[1888]), .Z(n10376) );
  XOR U10614 ( .A(n10376), .B(o[96]), .Z(N225) );
  NAND U10615 ( .A(x[225]), .B(y[1888]), .Z(n9731) );
  AND U10616 ( .A(x[224]), .B(y[1889]), .Z(n9737) );
  XNOR U10617 ( .A(n9737), .B(o[97]), .Z(n9732) );
  XOR U10618 ( .A(n9731), .B(n9732), .Z(n9734) );
  NAND U10619 ( .A(n10376), .B(o[96]), .Z(n9733) );
  XNOR U10620 ( .A(n9734), .B(n9733), .Z(N226) );
  IV U10621 ( .A(n9731), .Z(n9749) );
  NANDN U10622 ( .A(n9749), .B(n9732), .Z(n9736) );
  NAND U10623 ( .A(n9734), .B(n9733), .Z(n9735) );
  AND U10624 ( .A(n9736), .B(n9735), .Z(n9744) );
  AND U10625 ( .A(x[224]), .B(y[1890]), .Z(n9742) );
  XNOR U10626 ( .A(n9742), .B(o[98]), .Z(n9743) );
  XNOR U10627 ( .A(n9744), .B(n9743), .Z(n9746) );
  AND U10628 ( .A(n9737), .B(o[97]), .Z(n9751) );
  AND U10629 ( .A(y[1888]), .B(x[226]), .Z(n9739) );
  NAND U10630 ( .A(y[1889]), .B(x[225]), .Z(n9738) );
  XNOR U10631 ( .A(n9739), .B(n9738), .Z(n9750) );
  XNOR U10632 ( .A(n9751), .B(n9750), .Z(n9745) );
  XNOR U10633 ( .A(n9746), .B(n9745), .Z(N227) );
  AND U10634 ( .A(x[225]), .B(y[1890]), .Z(n9883) );
  NAND U10635 ( .A(x[226]), .B(y[1889]), .Z(n9761) );
  XOR U10636 ( .A(n9883), .B(n9763), .Z(n9765) );
  AND U10637 ( .A(y[1888]), .B(x[227]), .Z(n9741) );
  NAND U10638 ( .A(y[1891]), .B(x[224]), .Z(n9740) );
  XNOR U10639 ( .A(n9741), .B(n9740), .Z(n9755) );
  NAND U10640 ( .A(n9742), .B(o[98]), .Z(n9756) );
  XNOR U10641 ( .A(n9765), .B(n9764), .Z(n9770) );
  NANDN U10642 ( .A(n9744), .B(n9743), .Z(n9748) );
  NAND U10643 ( .A(n9746), .B(n9745), .Z(n9747) );
  AND U10644 ( .A(n9748), .B(n9747), .Z(n9769) );
  NANDN U10645 ( .A(n9761), .B(n9749), .Z(n9753) );
  NAND U10646 ( .A(n9751), .B(n9750), .Z(n9752) );
  NAND U10647 ( .A(n9753), .B(n9752), .Z(n9768) );
  XOR U10648 ( .A(n9769), .B(n9768), .Z(n9754) );
  XNOR U10649 ( .A(n9770), .B(n9754), .Z(N228) );
  AND U10650 ( .A(x[227]), .B(y[1891]), .Z(n9810) );
  NAND U10651 ( .A(n10376), .B(n9810), .Z(n9758) );
  NANDN U10652 ( .A(n9756), .B(n9755), .Z(n9757) );
  AND U10653 ( .A(n9758), .B(n9757), .Z(n9792) );
  AND U10654 ( .A(y[1892]), .B(x[224]), .Z(n9760) );
  NAND U10655 ( .A(y[1888]), .B(x[228]), .Z(n9759) );
  XNOR U10656 ( .A(n9760), .B(n9759), .Z(n9783) );
  ANDN U10657 ( .B(o[99]), .A(n9761), .Z(n9782) );
  XOR U10658 ( .A(n9783), .B(n9782), .Z(n9790) );
  AND U10659 ( .A(y[1890]), .B(x[226]), .Z(n9938) );
  NAND U10660 ( .A(y[1891]), .B(x[225]), .Z(n9762) );
  XNOR U10661 ( .A(n9938), .B(n9762), .Z(n9779) );
  AND U10662 ( .A(x[227]), .B(y[1889]), .Z(n9774) );
  XOR U10663 ( .A(o[100]), .B(n9774), .Z(n9778) );
  XOR U10664 ( .A(n9779), .B(n9778), .Z(n9789) );
  XOR U10665 ( .A(n9790), .B(n9789), .Z(n9791) );
  XOR U10666 ( .A(n9792), .B(n9791), .Z(n9788) );
  NAND U10667 ( .A(n9883), .B(n9763), .Z(n9767) );
  NAND U10668 ( .A(n9765), .B(n9764), .Z(n9766) );
  NAND U10669 ( .A(n9767), .B(n9766), .Z(n9786) );
  XOR U10670 ( .A(n9786), .B(n9787), .Z(n9771) );
  XNOR U10671 ( .A(n9788), .B(n9771), .Z(N229) );
  AND U10672 ( .A(y[1890]), .B(x[227]), .Z(n9773) );
  NAND U10673 ( .A(y[1892]), .B(x[225]), .Z(n9772) );
  XNOR U10674 ( .A(n9773), .B(n9772), .Z(n9797) );
  AND U10675 ( .A(x[228]), .B(y[1889]), .Z(n9808) );
  XOR U10676 ( .A(n9808), .B(o[101]), .Z(n9796) );
  XNOR U10677 ( .A(n9797), .B(n9796), .Z(n9800) );
  NAND U10678 ( .A(x[226]), .B(y[1891]), .Z(n9891) );
  AND U10679 ( .A(o[100]), .B(n9774), .Z(n9802) );
  AND U10680 ( .A(y[1888]), .B(x[229]), .Z(n9776) );
  NAND U10681 ( .A(y[1893]), .B(x[224]), .Z(n9775) );
  XNOR U10682 ( .A(n9776), .B(n9775), .Z(n9803) );
  XOR U10683 ( .A(n9802), .B(n9803), .Z(n9801) );
  XOR U10684 ( .A(n9891), .B(n9801), .Z(n9777) );
  XOR U10685 ( .A(n9800), .B(n9777), .Z(n9822) );
  NANDN U10686 ( .A(n9891), .B(n9883), .Z(n9781) );
  NAND U10687 ( .A(n9779), .B(n9778), .Z(n9780) );
  AND U10688 ( .A(n9781), .B(n9780), .Z(n9820) );
  AND U10689 ( .A(x[228]), .B(y[1892]), .Z(n10581) );
  NAND U10690 ( .A(n10581), .B(n10376), .Z(n9785) );
  NAND U10691 ( .A(n9783), .B(n9782), .Z(n9784) );
  NAND U10692 ( .A(n9785), .B(n9784), .Z(n9819) );
  XNOR U10693 ( .A(n9822), .B(n9821), .Z(n9815) );
  NAND U10694 ( .A(n9790), .B(n9789), .Z(n9794) );
  NANDN U10695 ( .A(n9792), .B(n9791), .Z(n9793) );
  NAND U10696 ( .A(n9794), .B(n9793), .Z(n9813) );
  IV U10697 ( .A(n9813), .Z(n9812) );
  XOR U10698 ( .A(n9814), .B(n9812), .Z(n9795) );
  XNOR U10699 ( .A(n9815), .B(n9795), .Z(N230) );
  AND U10700 ( .A(x[227]), .B(y[1892]), .Z(n9892) );
  NAND U10701 ( .A(n9892), .B(n9883), .Z(n9799) );
  NAND U10702 ( .A(n9797), .B(n9796), .Z(n9798) );
  NAND U10703 ( .A(n9799), .B(n9798), .Z(n9858) );
  XOR U10704 ( .A(n9858), .B(n9857), .Z(n9860) );
  AND U10705 ( .A(x[229]), .B(y[1893]), .Z(n10060) );
  NAND U10706 ( .A(n10376), .B(n10060), .Z(n9805) );
  NAND U10707 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U10708 ( .A(n9805), .B(n9804), .Z(n9827) );
  AND U10709 ( .A(y[1888]), .B(x[230]), .Z(n9807) );
  NAND U10710 ( .A(y[1894]), .B(x[224]), .Z(n9806) );
  XNOR U10711 ( .A(n9807), .B(n9806), .Z(n9833) );
  AND U10712 ( .A(n9808), .B(o[101]), .Z(n9834) );
  XOR U10713 ( .A(n9833), .B(n9834), .Z(n9826) );
  XOR U10714 ( .A(n9827), .B(n9826), .Z(n9829) );
  NAND U10715 ( .A(y[1892]), .B(x[226]), .Z(n9809) );
  XNOR U10716 ( .A(n9810), .B(n9809), .Z(n9838) );
  AND U10717 ( .A(y[1893]), .B(x[225]), .Z(n10092) );
  NAND U10718 ( .A(y[1890]), .B(x[228]), .Z(n9811) );
  XNOR U10719 ( .A(n10092), .B(n9811), .Z(n9842) );
  AND U10720 ( .A(x[229]), .B(y[1889]), .Z(n9849) );
  XOR U10721 ( .A(o[102]), .B(n9849), .Z(n9841) );
  XOR U10722 ( .A(n9842), .B(n9841), .Z(n9837) );
  XOR U10723 ( .A(n9838), .B(n9837), .Z(n9828) );
  XOR U10724 ( .A(n9829), .B(n9828), .Z(n9859) );
  XNOR U10725 ( .A(n9860), .B(n9859), .Z(n9853) );
  OR U10726 ( .A(n9814), .B(n9812), .Z(n9818) );
  ANDN U10727 ( .B(n9814), .A(n9813), .Z(n9816) );
  OR U10728 ( .A(n9816), .B(n9815), .Z(n9817) );
  AND U10729 ( .A(n9818), .B(n9817), .Z(n9852) );
  NANDN U10730 ( .A(n9820), .B(n9819), .Z(n9824) );
  NAND U10731 ( .A(n9822), .B(n9821), .Z(n9823) );
  NAND U10732 ( .A(n9824), .B(n9823), .Z(n9851) );
  IV U10733 ( .A(n9851), .Z(n9850) );
  XOR U10734 ( .A(n9852), .B(n9850), .Z(n9825) );
  XNOR U10735 ( .A(n9853), .B(n9825), .Z(N231) );
  NAND U10736 ( .A(n9827), .B(n9826), .Z(n9831) );
  NAND U10737 ( .A(n9829), .B(n9828), .Z(n9830) );
  AND U10738 ( .A(n9831), .B(n9830), .Z(n9867) );
  AND U10739 ( .A(y[1890]), .B(x[229]), .Z(n9961) );
  NAND U10740 ( .A(y[1894]), .B(x[225]), .Z(n9832) );
  XNOR U10741 ( .A(n9961), .B(n9832), .Z(n9885) );
  NAND U10742 ( .A(x[230]), .B(y[1889]), .Z(n9889) );
  XNOR U10743 ( .A(o[103]), .B(n9889), .Z(n9884) );
  XNOR U10744 ( .A(n9885), .B(n9884), .Z(n9903) );
  AND U10745 ( .A(x[230]), .B(y[1894]), .Z(n10112) );
  NAND U10746 ( .A(n10376), .B(n10112), .Z(n9836) );
  NAND U10747 ( .A(n9834), .B(n9833), .Z(n9835) );
  AND U10748 ( .A(n9836), .B(n9835), .Z(n9902) );
  XOR U10749 ( .A(n9903), .B(n9902), .Z(n9904) );
  NANDN U10750 ( .A(n9891), .B(n9892), .Z(n9840) );
  NAND U10751 ( .A(n9838), .B(n9837), .Z(n9839) );
  AND U10752 ( .A(n9840), .B(n9839), .Z(n9905) );
  XOR U10753 ( .A(n9904), .B(n9905), .Z(n9865) );
  AND U10754 ( .A(x[228]), .B(y[1893]), .Z(n10381) );
  NAND U10755 ( .A(n10381), .B(n9883), .Z(n9844) );
  NAND U10756 ( .A(n9842), .B(n9841), .Z(n9843) );
  AND U10757 ( .A(n9844), .B(n9843), .Z(n9880) );
  AND U10758 ( .A(y[1893]), .B(x[226]), .Z(n9846) );
  NAND U10759 ( .A(y[1891]), .B(x[228]), .Z(n9845) );
  XNOR U10760 ( .A(n9846), .B(n9845), .Z(n9893) );
  XNOR U10761 ( .A(n9893), .B(n9892), .Z(n9878) );
  AND U10762 ( .A(y[1888]), .B(x[231]), .Z(n9848) );
  NAND U10763 ( .A(y[1895]), .B(x[224]), .Z(n9847) );
  XNOR U10764 ( .A(n9848), .B(n9847), .Z(n9897) );
  AND U10765 ( .A(o[102]), .B(n9849), .Z(n9896) );
  XNOR U10766 ( .A(n9897), .B(n9896), .Z(n9877) );
  XOR U10767 ( .A(n9878), .B(n9877), .Z(n9879) );
  XOR U10768 ( .A(n9880), .B(n9879), .Z(n9864) );
  XOR U10769 ( .A(n9865), .B(n9864), .Z(n9866) );
  XNOR U10770 ( .A(n9867), .B(n9866), .Z(n9873) );
  OR U10771 ( .A(n9852), .B(n9850), .Z(n9856) );
  ANDN U10772 ( .B(n9852), .A(n9851), .Z(n9854) );
  OR U10773 ( .A(n9854), .B(n9853), .Z(n9855) );
  AND U10774 ( .A(n9856), .B(n9855), .Z(n9871) );
  NAND U10775 ( .A(n9858), .B(n9857), .Z(n9862) );
  NAND U10776 ( .A(n9860), .B(n9859), .Z(n9861) );
  AND U10777 ( .A(n9862), .B(n9861), .Z(n9872) );
  IV U10778 ( .A(n9872), .Z(n9870) );
  XOR U10779 ( .A(n9871), .B(n9870), .Z(n9863) );
  XNOR U10780 ( .A(n9873), .B(n9863), .Z(N232) );
  NAND U10781 ( .A(n9865), .B(n9864), .Z(n9869) );
  NAND U10782 ( .A(n9867), .B(n9866), .Z(n9868) );
  AND U10783 ( .A(n9869), .B(n9868), .Z(n9916) );
  NANDN U10784 ( .A(n9870), .B(n9871), .Z(n9876) );
  NOR U10785 ( .A(n9872), .B(n9871), .Z(n9874) );
  OR U10786 ( .A(n9874), .B(n9873), .Z(n9875) );
  AND U10787 ( .A(n9876), .B(n9875), .Z(n9915) );
  NAND U10788 ( .A(n9878), .B(n9877), .Z(n9882) );
  NAND U10789 ( .A(n9880), .B(n9879), .Z(n9881) );
  AND U10790 ( .A(n9882), .B(n9881), .Z(n9951) );
  AND U10791 ( .A(x[229]), .B(y[1894]), .Z(n10052) );
  NAND U10792 ( .A(n10052), .B(n9883), .Z(n9887) );
  NAND U10793 ( .A(n9885), .B(n9884), .Z(n9886) );
  NAND U10794 ( .A(n9887), .B(n9886), .Z(n9949) );
  AND U10795 ( .A(y[1891]), .B(x[229]), .Z(n10485) );
  NAND U10796 ( .A(y[1895]), .B(x[225]), .Z(n9888) );
  XNOR U10797 ( .A(n10485), .B(n9888), .Z(n9929) );
  ANDN U10798 ( .B(o[103]), .A(n9889), .Z(n9930) );
  XNOR U10799 ( .A(n9929), .B(n9930), .Z(n9934) );
  NAND U10800 ( .A(x[227]), .B(y[1893]), .Z(n10717) );
  AND U10801 ( .A(x[230]), .B(y[1890]), .Z(n9890) );
  AND U10802 ( .A(y[1894]), .B(x[226]), .Z(n10798) );
  XOR U10803 ( .A(n9890), .B(n10798), .Z(n9939) );
  XOR U10804 ( .A(n10581), .B(n9939), .Z(n9933) );
  XOR U10805 ( .A(n9934), .B(n9935), .Z(n9948) );
  XOR U10806 ( .A(n9949), .B(n9948), .Z(n9950) );
  XNOR U10807 ( .A(n9951), .B(n9950), .Z(n9912) );
  NANDN U10808 ( .A(n9891), .B(n10381), .Z(n9895) );
  NAND U10809 ( .A(n9893), .B(n9892), .Z(n9894) );
  NAND U10810 ( .A(n9895), .B(n9894), .Z(n9945) );
  AND U10811 ( .A(x[231]), .B(y[1895]), .Z(n10259) );
  NAND U10812 ( .A(n10376), .B(n10259), .Z(n9899) );
  NAND U10813 ( .A(n9897), .B(n9896), .Z(n9898) );
  NAND U10814 ( .A(n9899), .B(n9898), .Z(n9943) );
  AND U10815 ( .A(y[1888]), .B(x[232]), .Z(n9901) );
  NAND U10816 ( .A(y[1896]), .B(x[224]), .Z(n9900) );
  XNOR U10817 ( .A(n9901), .B(n9900), .Z(n9919) );
  NAND U10818 ( .A(x[231]), .B(y[1889]), .Z(n9925) );
  XOR U10819 ( .A(o[104]), .B(n9925), .Z(n9920) );
  XNOR U10820 ( .A(n9919), .B(n9920), .Z(n9942) );
  XOR U10821 ( .A(n9943), .B(n9942), .Z(n9944) );
  XNOR U10822 ( .A(n9945), .B(n9944), .Z(n9910) );
  NAND U10823 ( .A(n9903), .B(n9902), .Z(n9907) );
  NAND U10824 ( .A(n9905), .B(n9904), .Z(n9906) );
  NAND U10825 ( .A(n9907), .B(n9906), .Z(n9909) );
  XOR U10826 ( .A(n9910), .B(n9909), .Z(n9911) );
  XOR U10827 ( .A(n9912), .B(n9911), .Z(n9917) );
  XNOR U10828 ( .A(n9915), .B(n9917), .Z(n9908) );
  XOR U10829 ( .A(n9916), .B(n9908), .Z(N233) );
  NAND U10830 ( .A(n9910), .B(n9909), .Z(n9914) );
  NAND U10831 ( .A(n9912), .B(n9911), .Z(n9913) );
  NAND U10832 ( .A(n9914), .B(n9913), .Z(n10003) );
  IV U10833 ( .A(n10003), .Z(n10001) );
  AND U10834 ( .A(x[232]), .B(y[1896]), .Z(n9918) );
  NAND U10835 ( .A(n9918), .B(n10376), .Z(n9922) );
  NANDN U10836 ( .A(n9920), .B(n9919), .Z(n9921) );
  AND U10837 ( .A(n9922), .B(n9921), .Z(n9988) );
  AND U10838 ( .A(y[1892]), .B(x[229]), .Z(n9924) );
  NAND U10839 ( .A(y[1890]), .B(x[231]), .Z(n9923) );
  XNOR U10840 ( .A(n9924), .B(n9923), .Z(n9963) );
  ANDN U10841 ( .B(o[104]), .A(n9925), .Z(n9962) );
  XOR U10842 ( .A(n9963), .B(n9962), .Z(n9986) );
  AND U10843 ( .A(y[1888]), .B(x[233]), .Z(n9927) );
  NAND U10844 ( .A(y[1897]), .B(x[224]), .Z(n9926) );
  XNOR U10845 ( .A(n9927), .B(n9926), .Z(n9970) );
  NAND U10846 ( .A(x[232]), .B(y[1889]), .Z(n9979) );
  XNOR U10847 ( .A(o[105]), .B(n9979), .Z(n9969) );
  XNOR U10848 ( .A(n9970), .B(n9969), .Z(n9985) );
  XNOR U10849 ( .A(n9986), .B(n9985), .Z(n9987) );
  XOR U10850 ( .A(n9988), .B(n9987), .Z(n9984) );
  AND U10851 ( .A(y[1891]), .B(x[230]), .Z(n10328) );
  NAND U10852 ( .A(y[1896]), .B(x[225]), .Z(n9928) );
  XNOR U10853 ( .A(n10328), .B(n9928), .Z(n9974) );
  XOR U10854 ( .A(n10381), .B(n9974), .Z(n9992) );
  NAND U10855 ( .A(x[226]), .B(y[1895]), .Z(n10537) );
  NAND U10856 ( .A(x[227]), .B(y[1894]), .Z(n10336) );
  XOR U10857 ( .A(n10537), .B(n10336), .Z(n9991) );
  XOR U10858 ( .A(n9992), .B(n9991), .Z(n9981) );
  NAND U10859 ( .A(x[229]), .B(y[1895]), .Z(n10166) );
  AND U10860 ( .A(x[225]), .B(y[1891]), .Z(n9973) );
  NANDN U10861 ( .A(n10166), .B(n9973), .Z(n9932) );
  NAND U10862 ( .A(n9930), .B(n9929), .Z(n9931) );
  NAND U10863 ( .A(n9932), .B(n9931), .Z(n9982) );
  XOR U10864 ( .A(n9981), .B(n9982), .Z(n9983) );
  XOR U10865 ( .A(n9984), .B(n9983), .Z(n9957) );
  NANDN U10866 ( .A(n9933), .B(n10717), .Z(n9937) );
  NANDN U10867 ( .A(n9935), .B(n9934), .Z(n9936) );
  NAND U10868 ( .A(n9937), .B(n9936), .Z(n9955) );
  NAND U10869 ( .A(n10112), .B(n9938), .Z(n9941) );
  NAND U10870 ( .A(n10581), .B(n9939), .Z(n9940) );
  AND U10871 ( .A(n9941), .B(n9940), .Z(n9956) );
  XNOR U10872 ( .A(n9955), .B(n9956), .Z(n9958) );
  NAND U10873 ( .A(n9943), .B(n9942), .Z(n9947) );
  NAND U10874 ( .A(n9945), .B(n9944), .Z(n9946) );
  NAND U10875 ( .A(n9947), .B(n9946), .Z(n9996) );
  NAND U10876 ( .A(n9949), .B(n9948), .Z(n9953) );
  NAND U10877 ( .A(n9951), .B(n9950), .Z(n9952) );
  NAND U10878 ( .A(n9953), .B(n9952), .Z(n9995) );
  XOR U10879 ( .A(n9996), .B(n9995), .Z(n9998) );
  XOR U10880 ( .A(n9997), .B(n9998), .Z(n10004) );
  XNOR U10881 ( .A(n10002), .B(n10004), .Z(n9954) );
  XOR U10882 ( .A(n10001), .B(n9954), .Z(N234) );
  NAND U10883 ( .A(n9956), .B(n9955), .Z(n9960) );
  NANDN U10884 ( .A(n9958), .B(n9957), .Z(n9959) );
  NAND U10885 ( .A(n9960), .B(n9959), .Z(n10014) );
  AND U10886 ( .A(x[231]), .B(y[1892]), .Z(n10054) );
  NAND U10887 ( .A(n10054), .B(n9961), .Z(n9965) );
  NAND U10888 ( .A(n9963), .B(n9962), .Z(n9964) );
  AND U10889 ( .A(n9965), .B(n9964), .Z(n10067) );
  AND U10890 ( .A(y[1891]), .B(x[231]), .Z(n9967) );
  NAND U10891 ( .A(y[1894]), .B(x[228]), .Z(n9966) );
  XNOR U10892 ( .A(n9967), .B(n9966), .Z(n10038) );
  AND U10893 ( .A(x[230]), .B(y[1892]), .Z(n10037) );
  XNOR U10894 ( .A(n10038), .B(n10037), .Z(n10065) );
  AND U10895 ( .A(x[232]), .B(y[1890]), .Z(n10235) );
  AND U10896 ( .A(x[233]), .B(y[1889]), .Z(n10048) );
  XOR U10897 ( .A(o[106]), .B(n10048), .Z(n10059) );
  XOR U10898 ( .A(n10235), .B(n10059), .Z(n10061) );
  XNOR U10899 ( .A(n10061), .B(n10060), .Z(n10064) );
  XOR U10900 ( .A(n10065), .B(n10064), .Z(n10066) );
  XOR U10901 ( .A(n10067), .B(n10066), .Z(n10027) );
  AND U10902 ( .A(x[233]), .B(y[1897]), .Z(n9968) );
  NAND U10903 ( .A(n9968), .B(n10376), .Z(n9972) );
  NAND U10904 ( .A(n9970), .B(n9969), .Z(n9971) );
  AND U10905 ( .A(n9972), .B(n9971), .Z(n10025) );
  AND U10906 ( .A(x[230]), .B(y[1896]), .Z(n10269) );
  NAND U10907 ( .A(n10269), .B(n9973), .Z(n9976) );
  NAND U10908 ( .A(n10381), .B(n9974), .Z(n9975) );
  NAND U10909 ( .A(n9976), .B(n9975), .Z(n10033) );
  AND U10910 ( .A(y[1888]), .B(x[234]), .Z(n9978) );
  NAND U10911 ( .A(y[1898]), .B(x[224]), .Z(n9977) );
  XNOR U10912 ( .A(n9978), .B(n9977), .Z(n10043) );
  ANDN U10913 ( .B(o[105]), .A(n9979), .Z(n10042) );
  XOR U10914 ( .A(n10043), .B(n10042), .Z(n10031) );
  AND U10915 ( .A(y[1895]), .B(x[227]), .Z(n10954) );
  NAND U10916 ( .A(y[1897]), .B(x[225]), .Z(n9980) );
  XNOR U10917 ( .A(n10954), .B(n9980), .Z(n10055) );
  AND U10918 ( .A(x[226]), .B(y[1896]), .Z(n10056) );
  XOR U10919 ( .A(n10055), .B(n10056), .Z(n10030) );
  XOR U10920 ( .A(n10031), .B(n10030), .Z(n10032) );
  XOR U10921 ( .A(n10033), .B(n10032), .Z(n10024) );
  XNOR U10922 ( .A(n10025), .B(n10024), .Z(n10026) );
  XOR U10923 ( .A(n10027), .B(n10026), .Z(n10013) );
  NANDN U10924 ( .A(n9986), .B(n9985), .Z(n9990) );
  NAND U10925 ( .A(n9988), .B(n9987), .Z(n9989) );
  AND U10926 ( .A(n9990), .B(n9989), .Z(n10018) );
  IV U10927 ( .A(n10537), .Z(n10628) );
  ANDN U10928 ( .B(n10336), .A(n10628), .Z(n9994) );
  NANDN U10929 ( .A(n9992), .B(n9991), .Z(n9993) );
  NANDN U10930 ( .A(n9994), .B(n9993), .Z(n10019) );
  XOR U10931 ( .A(n10018), .B(n10019), .Z(n10021) );
  XNOR U10932 ( .A(n10020), .B(n10021), .Z(n10012) );
  XOR U10933 ( .A(n10013), .B(n10012), .Z(n10015) );
  XOR U10934 ( .A(n10014), .B(n10015), .Z(n10011) );
  NAND U10935 ( .A(n9996), .B(n9995), .Z(n10000) );
  NAND U10936 ( .A(n9998), .B(n9997), .Z(n9999) );
  NAND U10937 ( .A(n10000), .B(n9999), .Z(n10010) );
  NANDN U10938 ( .A(n10001), .B(n10002), .Z(n10007) );
  NOR U10939 ( .A(n10003), .B(n10002), .Z(n10005) );
  OR U10940 ( .A(n10005), .B(n10004), .Z(n10006) );
  AND U10941 ( .A(n10007), .B(n10006), .Z(n10009) );
  XOR U10942 ( .A(n10010), .B(n10009), .Z(n10008) );
  XNOR U10943 ( .A(n10011), .B(n10008), .Z(N235) );
  NAND U10944 ( .A(n10013), .B(n10012), .Z(n10017) );
  NAND U10945 ( .A(n10015), .B(n10014), .Z(n10016) );
  AND U10946 ( .A(n10017), .B(n10016), .Z(n10070) );
  XNOR U10947 ( .A(n10071), .B(n10070), .Z(n10073) );
  NANDN U10948 ( .A(n10019), .B(n10018), .Z(n10023) );
  OR U10949 ( .A(n10021), .B(n10020), .Z(n10022) );
  AND U10950 ( .A(n10023), .B(n10022), .Z(n10079) );
  NANDN U10951 ( .A(n10025), .B(n10024), .Z(n10029) );
  NANDN U10952 ( .A(n10027), .B(n10026), .Z(n10028) );
  AND U10953 ( .A(n10029), .B(n10028), .Z(n10077) );
  NAND U10954 ( .A(n10031), .B(n10030), .Z(n10035) );
  NAND U10955 ( .A(n10033), .B(n10032), .Z(n10034) );
  NAND U10956 ( .A(n10035), .B(n10034), .Z(n10134) );
  AND U10957 ( .A(x[231]), .B(y[1894]), .Z(n10161) );
  AND U10958 ( .A(x[228]), .B(y[1891]), .Z(n10036) );
  NAND U10959 ( .A(n10161), .B(n10036), .Z(n10040) );
  NAND U10960 ( .A(n10038), .B(n10037), .Z(n10039) );
  NAND U10961 ( .A(n10040), .B(n10039), .Z(n10132) );
  AND U10962 ( .A(x[234]), .B(y[1898]), .Z(n10041) );
  NAND U10963 ( .A(n10041), .B(n10376), .Z(n10045) );
  NAND U10964 ( .A(n10043), .B(n10042), .Z(n10044) );
  NAND U10965 ( .A(n10045), .B(n10044), .Z(n10128) );
  AND U10966 ( .A(y[1888]), .B(x[235]), .Z(n10047) );
  NAND U10967 ( .A(y[1899]), .B(x[224]), .Z(n10046) );
  XNOR U10968 ( .A(n10047), .B(n10046), .Z(n10103) );
  AND U10969 ( .A(o[106]), .B(n10048), .Z(n10102) );
  XOR U10970 ( .A(n10103), .B(n10102), .Z(n10126) );
  AND U10971 ( .A(y[1893]), .B(x[230]), .Z(n10050) );
  NAND U10972 ( .A(y[1898]), .B(x[225]), .Z(n10049) );
  XNOR U10973 ( .A(n10050), .B(n10049), .Z(n10094) );
  NAND U10974 ( .A(x[234]), .B(y[1889]), .Z(n10113) );
  XOR U10975 ( .A(n10094), .B(n10093), .Z(n10125) );
  XOR U10976 ( .A(n10126), .B(n10125), .Z(n10127) );
  XOR U10977 ( .A(n10128), .B(n10127), .Z(n10131) );
  XOR U10978 ( .A(n10132), .B(n10131), .Z(n10133) );
  XNOR U10979 ( .A(n10134), .B(n10133), .Z(n10116) );
  AND U10980 ( .A(x[227]), .B(y[1896]), .Z(n11083) );
  NAND U10981 ( .A(y[1897]), .B(x[226]), .Z(n10051) );
  XNOR U10982 ( .A(n10052), .B(n10051), .Z(n10089) );
  AND U10983 ( .A(x[228]), .B(y[1895]), .Z(n10088) );
  XNOR U10984 ( .A(n10089), .B(n10088), .Z(n10120) );
  XNOR U10985 ( .A(n11083), .B(n10120), .Z(n10122) );
  NAND U10986 ( .A(y[1890]), .B(x[233]), .Z(n10053) );
  XNOR U10987 ( .A(n10054), .B(n10053), .Z(n10108) );
  AND U10988 ( .A(x[232]), .B(y[1891]), .Z(n10107) );
  XNOR U10989 ( .A(n10108), .B(n10107), .Z(n10121) );
  XNOR U10990 ( .A(n10122), .B(n10121), .Z(n10085) );
  NAND U10991 ( .A(x[227]), .B(y[1897]), .Z(n10157) );
  AND U10992 ( .A(x[225]), .B(y[1895]), .Z(n10371) );
  NANDN U10993 ( .A(n10157), .B(n10371), .Z(n10058) );
  NAND U10994 ( .A(n10056), .B(n10055), .Z(n10057) );
  NAND U10995 ( .A(n10058), .B(n10057), .Z(n10083) );
  NAND U10996 ( .A(n10235), .B(n10059), .Z(n10063) );
  NAND U10997 ( .A(n10061), .B(n10060), .Z(n10062) );
  NAND U10998 ( .A(n10063), .B(n10062), .Z(n10082) );
  XOR U10999 ( .A(n10083), .B(n10082), .Z(n10084) );
  XNOR U11000 ( .A(n10085), .B(n10084), .Z(n10115) );
  NAND U11001 ( .A(n10065), .B(n10064), .Z(n10069) );
  NAND U11002 ( .A(n10067), .B(n10066), .Z(n10068) );
  NAND U11003 ( .A(n10069), .B(n10068), .Z(n10114) );
  XOR U11004 ( .A(n10115), .B(n10114), .Z(n10117) );
  XNOR U11005 ( .A(n10116), .B(n10117), .Z(n10076) );
  XNOR U11006 ( .A(n10077), .B(n10076), .Z(n10078) );
  XNOR U11007 ( .A(n10079), .B(n10078), .Z(n10072) );
  XOR U11008 ( .A(n10073), .B(n10072), .Z(N236) );
  NANDN U11009 ( .A(n10071), .B(n10070), .Z(n10075) );
  NAND U11010 ( .A(n10073), .B(n10072), .Z(n10074) );
  NAND U11011 ( .A(n10075), .B(n10074), .Z(n10202) );
  NANDN U11012 ( .A(n10077), .B(n10076), .Z(n10081) );
  NANDN U11013 ( .A(n10079), .B(n10078), .Z(n10080) );
  NAND U11014 ( .A(n10081), .B(n10080), .Z(n10201) );
  NAND U11015 ( .A(n10083), .B(n10082), .Z(n10087) );
  NAND U11016 ( .A(n10085), .B(n10084), .Z(n10086) );
  NAND U11017 ( .A(n10087), .B(n10086), .Z(n10198) );
  AND U11018 ( .A(x[229]), .B(y[1897]), .Z(n10619) );
  NAND U11019 ( .A(n10798), .B(n10619), .Z(n10091) );
  NAND U11020 ( .A(n10089), .B(n10088), .Z(n10090) );
  NAND U11021 ( .A(n10091), .B(n10090), .Z(n10145) );
  AND U11022 ( .A(x[230]), .B(y[1898]), .Z(n10388) );
  NAND U11023 ( .A(n10388), .B(n10092), .Z(n10096) );
  NAND U11024 ( .A(n10094), .B(n10093), .Z(n10095) );
  NAND U11025 ( .A(n10096), .B(n10095), .Z(n10144) );
  XOR U11026 ( .A(n10145), .B(n10144), .Z(n10147) );
  AND U11027 ( .A(x[233]), .B(y[1891]), .Z(n10793) );
  AND U11028 ( .A(x[234]), .B(y[1890]), .Z(n10848) );
  NAND U11029 ( .A(y[1896]), .B(x[228]), .Z(n10097) );
  XOR U11030 ( .A(n10848), .B(n10097), .Z(n10188) );
  NAND U11031 ( .A(x[231]), .B(y[1893]), .Z(n10165) );
  XOR U11032 ( .A(n10166), .B(n10165), .Z(n10168) );
  AND U11033 ( .A(y[1888]), .B(x[236]), .Z(n10099) );
  NAND U11034 ( .A(y[1900]), .B(x[224]), .Z(n10098) );
  XNOR U11035 ( .A(n10099), .B(n10098), .Z(n10181) );
  NAND U11036 ( .A(x[235]), .B(y[1889]), .Z(n10162) );
  XOR U11037 ( .A(o[108]), .B(n10162), .Z(n10182) );
  AND U11038 ( .A(y[1898]), .B(x[226]), .Z(n10101) );
  NAND U11039 ( .A(y[1892]), .B(x[232]), .Z(n10100) );
  XNOR U11040 ( .A(n10101), .B(n10100), .Z(n10156) );
  XOR U11041 ( .A(n10151), .B(n10150), .Z(n10153) );
  XOR U11042 ( .A(n10152), .B(n10153), .Z(n10146) );
  XOR U11043 ( .A(n10147), .B(n10146), .Z(n10196) );
  AND U11044 ( .A(x[235]), .B(y[1899]), .Z(n11215) );
  NAND U11045 ( .A(n11215), .B(n10376), .Z(n10105) );
  NAND U11046 ( .A(n10103), .B(n10102), .Z(n10104) );
  NAND U11047 ( .A(n10105), .B(n10104), .Z(n10174) );
  AND U11048 ( .A(x[231]), .B(y[1890]), .Z(n10314) );
  AND U11049 ( .A(x[233]), .B(y[1892]), .Z(n10106) );
  NAND U11050 ( .A(n10314), .B(n10106), .Z(n10110) );
  NAND U11051 ( .A(n10108), .B(n10107), .Z(n10109) );
  NAND U11052 ( .A(n10110), .B(n10109), .Z(n10172) );
  NAND U11053 ( .A(y[1899]), .B(x[225]), .Z(n10111) );
  XNOR U11054 ( .A(n10112), .B(n10111), .Z(n10178) );
  ANDN U11055 ( .B(o[107]), .A(n10113), .Z(n10177) );
  XOR U11056 ( .A(n10178), .B(n10177), .Z(n10171) );
  XOR U11057 ( .A(n10172), .B(n10171), .Z(n10173) );
  XOR U11058 ( .A(n10174), .B(n10173), .Z(n10195) );
  XOR U11059 ( .A(n10196), .B(n10195), .Z(n10197) );
  XNOR U11060 ( .A(n10198), .B(n10197), .Z(n10205) );
  NAND U11061 ( .A(n10115), .B(n10114), .Z(n10119) );
  NAND U11062 ( .A(n10117), .B(n10116), .Z(n10118) );
  NAND U11063 ( .A(n10119), .B(n10118), .Z(n10204) );
  XOR U11064 ( .A(n10205), .B(n10204), .Z(n10207) );
  NANDN U11065 ( .A(n11083), .B(n10120), .Z(n10124) );
  NAND U11066 ( .A(n10122), .B(n10121), .Z(n10123) );
  NAND U11067 ( .A(n10124), .B(n10123), .Z(n10139) );
  NAND U11068 ( .A(n10126), .B(n10125), .Z(n10130) );
  NAND U11069 ( .A(n10128), .B(n10127), .Z(n10129) );
  AND U11070 ( .A(n10130), .B(n10129), .Z(n10138) );
  XOR U11071 ( .A(n10139), .B(n10138), .Z(n10140) );
  NAND U11072 ( .A(n10132), .B(n10131), .Z(n10136) );
  NAND U11073 ( .A(n10134), .B(n10133), .Z(n10135) );
  AND U11074 ( .A(n10136), .B(n10135), .Z(n10141) );
  XOR U11075 ( .A(n10140), .B(n10141), .Z(n10206) );
  XOR U11076 ( .A(n10207), .B(n10206), .Z(n10203) );
  XOR U11077 ( .A(n10201), .B(n10203), .Z(n10137) );
  XNOR U11078 ( .A(n10202), .B(n10137), .Z(N237) );
  NAND U11079 ( .A(n10139), .B(n10138), .Z(n10143) );
  NAND U11080 ( .A(n10141), .B(n10140), .Z(n10142) );
  AND U11081 ( .A(n10143), .B(n10142), .Z(n10286) );
  NAND U11082 ( .A(n10145), .B(n10144), .Z(n10149) );
  NAND U11083 ( .A(n10147), .B(n10146), .Z(n10148) );
  AND U11084 ( .A(n10149), .B(n10148), .Z(n10212) );
  NAND U11085 ( .A(n10151), .B(n10150), .Z(n10155) );
  NAND U11086 ( .A(n10153), .B(n10152), .Z(n10154) );
  NAND U11087 ( .A(n10155), .B(n10154), .Z(n10219) );
  AND U11088 ( .A(y[1898]), .B(x[232]), .Z(n11487) );
  AND U11089 ( .A(x[226]), .B(y[1892]), .Z(n10324) );
  NAND U11090 ( .A(n11487), .B(n10324), .Z(n10159) );
  NANDN U11091 ( .A(n10157), .B(n10156), .Z(n10158) );
  AND U11092 ( .A(n10159), .B(n10158), .Z(n10248) );
  NAND U11093 ( .A(y[1900]), .B(x[225]), .Z(n10160) );
  XNOR U11094 ( .A(n10161), .B(n10160), .Z(n10241) );
  ANDN U11095 ( .B(o[108]), .A(n10162), .Z(n10240) );
  XOR U11096 ( .A(n10241), .B(n10240), .Z(n10245) );
  AND U11097 ( .A(x[230]), .B(y[1895]), .Z(n11253) );
  AND U11098 ( .A(y[1899]), .B(x[226]), .Z(n10164) );
  NAND U11099 ( .A(y[1892]), .B(x[233]), .Z(n10163) );
  XOR U11100 ( .A(n10164), .B(n10163), .Z(n10252) );
  XOR U11101 ( .A(n11253), .B(n10252), .Z(n10246) );
  NAND U11102 ( .A(n10166), .B(n10165), .Z(n10170) );
  ANDN U11103 ( .B(n10168), .A(n10167), .Z(n10169) );
  ANDN U11104 ( .B(n10170), .A(n10169), .Z(n10217) );
  XOR U11105 ( .A(n10218), .B(n10217), .Z(n10220) );
  XOR U11106 ( .A(n10219), .B(n10220), .Z(n10211) );
  NAND U11107 ( .A(n10172), .B(n10171), .Z(n10176) );
  NAND U11108 ( .A(n10174), .B(n10173), .Z(n10175) );
  AND U11109 ( .A(n10176), .B(n10175), .Z(n10226) );
  AND U11110 ( .A(x[230]), .B(y[1899]), .Z(n10620) );
  AND U11111 ( .A(x[225]), .B(y[1894]), .Z(n10239) );
  NAND U11112 ( .A(n10620), .B(n10239), .Z(n10180) );
  NAND U11113 ( .A(n10178), .B(n10177), .Z(n10179) );
  AND U11114 ( .A(n10180), .B(n10179), .Z(n10232) );
  AND U11115 ( .A(x[236]), .B(y[1900]), .Z(n11495) );
  NAND U11116 ( .A(n10376), .B(n11495), .Z(n10184) );
  NANDN U11117 ( .A(n10182), .B(n10181), .Z(n10183) );
  AND U11118 ( .A(n10184), .B(n10183), .Z(n10230) );
  AND U11119 ( .A(x[234]), .B(y[1891]), .Z(n11095) );
  AND U11120 ( .A(y[1890]), .B(x[235]), .Z(n11056) );
  NAND U11121 ( .A(y[1893]), .B(x[232]), .Z(n10185) );
  XOR U11122 ( .A(n11056), .B(n10185), .Z(n10236) );
  XNOR U11123 ( .A(n11095), .B(n10236), .Z(n10229) );
  AND U11124 ( .A(x[234]), .B(y[1896]), .Z(n10187) );
  AND U11125 ( .A(x[228]), .B(y[1890]), .Z(n10186) );
  NAND U11126 ( .A(n10187), .B(n10186), .Z(n10190) );
  NANDN U11127 ( .A(n10188), .B(n10793), .Z(n10189) );
  AND U11128 ( .A(n10190), .B(n10189), .Z(n10273) );
  AND U11129 ( .A(y[1888]), .B(x[237]), .Z(n10192) );
  NAND U11130 ( .A(y[1901]), .B(x[224]), .Z(n10191) );
  XNOR U11131 ( .A(n10192), .B(n10191), .Z(n10264) );
  NAND U11132 ( .A(x[236]), .B(y[1889]), .Z(n10257) );
  XOR U11133 ( .A(o[109]), .B(n10257), .Z(n10265) );
  XNOR U11134 ( .A(n10264), .B(n10265), .Z(n10270) );
  AND U11135 ( .A(y[1896]), .B(x[229]), .Z(n10194) );
  NAND U11136 ( .A(y[1898]), .B(x[227]), .Z(n10193) );
  XNOR U11137 ( .A(n10194), .B(n10193), .Z(n10260) );
  NAND U11138 ( .A(x[228]), .B(y[1897]), .Z(n10261) );
  XOR U11139 ( .A(n10260), .B(n10261), .Z(n10271) );
  XOR U11140 ( .A(n10224), .B(n10223), .Z(n10225) );
  XNOR U11141 ( .A(n10214), .B(n10213), .Z(n10284) );
  NAND U11142 ( .A(n10196), .B(n10195), .Z(n10200) );
  NAND U11143 ( .A(n10198), .B(n10197), .Z(n10199) );
  AND U11144 ( .A(n10200), .B(n10199), .Z(n10283) );
  XOR U11145 ( .A(n10284), .B(n10283), .Z(n10285) );
  XOR U11146 ( .A(n10286), .B(n10285), .Z(n10279) );
  NAND U11147 ( .A(n10205), .B(n10204), .Z(n10209) );
  NAND U11148 ( .A(n10207), .B(n10206), .Z(n10208) );
  NAND U11149 ( .A(n10209), .B(n10208), .Z(n10278) );
  IV U11150 ( .A(n10278), .Z(n10276) );
  XOR U11151 ( .A(n10277), .B(n10276), .Z(n10210) );
  XNOR U11152 ( .A(n10279), .B(n10210), .Z(N238) );
  NANDN U11153 ( .A(n10212), .B(n10211), .Z(n10216) );
  NAND U11154 ( .A(n10214), .B(n10213), .Z(n10215) );
  AND U11155 ( .A(n10216), .B(n10215), .Z(n10365) );
  NAND U11156 ( .A(n10218), .B(n10217), .Z(n10222) );
  NAND U11157 ( .A(n10220), .B(n10219), .Z(n10221) );
  NAND U11158 ( .A(n10222), .B(n10221), .Z(n10364) );
  NAND U11159 ( .A(n10224), .B(n10223), .Z(n10228) );
  NANDN U11160 ( .A(n10226), .B(n10225), .Z(n10227) );
  AND U11161 ( .A(n10228), .B(n10227), .Z(n10293) );
  NANDN U11162 ( .A(n10230), .B(n10229), .Z(n10234) );
  NANDN U11163 ( .A(n10232), .B(n10231), .Z(n10233) );
  AND U11164 ( .A(n10234), .B(n10233), .Z(n10299) );
  AND U11165 ( .A(x[235]), .B(y[1893]), .Z(n10402) );
  NAND U11166 ( .A(n10402), .B(n10235), .Z(n10238) );
  NANDN U11167 ( .A(n10236), .B(n11095), .Z(n10237) );
  AND U11168 ( .A(n10238), .B(n10237), .Z(n10350) );
  NAND U11169 ( .A(x[231]), .B(y[1900]), .Z(n10808) );
  XNOR U11170 ( .A(n10350), .B(n10349), .Z(n10352) );
  AND U11171 ( .A(x[228]), .B(y[1898]), .Z(n10727) );
  AND U11172 ( .A(y[1899]), .B(x[227]), .Z(n10243) );
  NAND U11173 ( .A(y[1894]), .B(x[232]), .Z(n10242) );
  XOR U11174 ( .A(n10243), .B(n10242), .Z(n10337) );
  XOR U11175 ( .A(n10619), .B(n10337), .Z(n10346) );
  XNOR U11176 ( .A(n10727), .B(n10346), .Z(n10348) );
  AND U11177 ( .A(x[233]), .B(y[1893]), .Z(n10919) );
  AND U11178 ( .A(y[1900]), .B(x[226]), .Z(n10244) );
  AND U11179 ( .A(y[1892]), .B(x[234]), .Z(n10949) );
  XOR U11180 ( .A(n10244), .B(n10949), .Z(n10325) );
  XOR U11181 ( .A(n10919), .B(n10325), .Z(n10347) );
  XOR U11182 ( .A(n10348), .B(n10347), .Z(n10351) );
  XOR U11183 ( .A(n10352), .B(n10351), .Z(n10297) );
  NANDN U11184 ( .A(n10246), .B(n10245), .Z(n10250) );
  NANDN U11185 ( .A(n10248), .B(n10247), .Z(n10249) );
  AND U11186 ( .A(n10250), .B(n10249), .Z(n10296) );
  XOR U11187 ( .A(n10299), .B(n10298), .Z(n10291) );
  AND U11188 ( .A(x[233]), .B(y[1899]), .Z(n10251) );
  NAND U11189 ( .A(n10251), .B(n10324), .Z(n10254) );
  NANDN U11190 ( .A(n10252), .B(n11253), .Z(n10253) );
  AND U11191 ( .A(n10254), .B(n10253), .Z(n10310) );
  AND U11192 ( .A(y[1888]), .B(x[238]), .Z(n10256) );
  NAND U11193 ( .A(y[1902]), .B(x[224]), .Z(n10255) );
  XNOR U11194 ( .A(n10256), .B(n10255), .Z(n10334) );
  ANDN U11195 ( .B(o[109]), .A(n10257), .Z(n10333) );
  XOR U11196 ( .A(n10334), .B(n10333), .Z(n10308) );
  NAND U11197 ( .A(y[1890]), .B(x[236]), .Z(n10258) );
  XNOR U11198 ( .A(n10259), .B(n10258), .Z(n10315) );
  NAND U11199 ( .A(x[237]), .B(y[1889]), .Z(n10323) );
  XOR U11200 ( .A(o[110]), .B(n10323), .Z(n10316) );
  XOR U11201 ( .A(n10315), .B(n10316), .Z(n10309) );
  XOR U11202 ( .A(n10308), .B(n10309), .Z(n10311) );
  XOR U11203 ( .A(n10310), .B(n10311), .Z(n10356) );
  AND U11204 ( .A(x[229]), .B(y[1898]), .Z(n10389) );
  NAND U11205 ( .A(n11083), .B(n10389), .Z(n10263) );
  NANDN U11206 ( .A(n10261), .B(n10260), .Z(n10262) );
  AND U11207 ( .A(n10263), .B(n10262), .Z(n10304) );
  AND U11208 ( .A(x[237]), .B(y[1901]), .Z(n11744) );
  NAND U11209 ( .A(n11744), .B(n10376), .Z(n10267) );
  NANDN U11210 ( .A(n10265), .B(n10264), .Z(n10266) );
  AND U11211 ( .A(n10267), .B(n10266), .Z(n10303) );
  NAND U11212 ( .A(y[1891]), .B(x[235]), .Z(n10268) );
  XNOR U11213 ( .A(n10269), .B(n10268), .Z(n10329) );
  NAND U11214 ( .A(x[225]), .B(y[1901]), .Z(n10330) );
  XNOR U11215 ( .A(n10329), .B(n10330), .Z(n10302) );
  XOR U11216 ( .A(n10303), .B(n10302), .Z(n10305) );
  XNOR U11217 ( .A(n10304), .B(n10305), .Z(n10355) );
  NANDN U11218 ( .A(n10271), .B(n10270), .Z(n10275) );
  NANDN U11219 ( .A(n10273), .B(n10272), .Z(n10274) );
  AND U11220 ( .A(n10275), .B(n10274), .Z(n10357) );
  XNOR U11221 ( .A(n10358), .B(n10357), .Z(n10290) );
  XNOR U11222 ( .A(n10367), .B(n10366), .Z(n10363) );
  NANDN U11223 ( .A(n10276), .B(n10277), .Z(n10282) );
  NOR U11224 ( .A(n10278), .B(n10277), .Z(n10280) );
  OR U11225 ( .A(n10280), .B(n10279), .Z(n10281) );
  AND U11226 ( .A(n10282), .B(n10281), .Z(n10361) );
  NAND U11227 ( .A(n10284), .B(n10283), .Z(n10288) );
  NANDN U11228 ( .A(n10286), .B(n10285), .Z(n10287) );
  AND U11229 ( .A(n10288), .B(n10287), .Z(n10362) );
  XOR U11230 ( .A(n10361), .B(n10362), .Z(n10289) );
  XNOR U11231 ( .A(n10363), .B(n10289), .Z(N239) );
  NANDN U11232 ( .A(n10291), .B(n10290), .Z(n10295) );
  NANDN U11233 ( .A(n10293), .B(n10292), .Z(n10294) );
  AND U11234 ( .A(n10295), .B(n10294), .Z(n10463) );
  NANDN U11235 ( .A(n10297), .B(n10296), .Z(n10301) );
  NAND U11236 ( .A(n10299), .B(n10298), .Z(n10300) );
  NAND U11237 ( .A(n10301), .B(n10300), .Z(n10431) );
  NANDN U11238 ( .A(n10303), .B(n10302), .Z(n10307) );
  OR U11239 ( .A(n10305), .B(n10304), .Z(n10306) );
  AND U11240 ( .A(n10307), .B(n10306), .Z(n10438) );
  NANDN U11241 ( .A(n10309), .B(n10308), .Z(n10313) );
  OR U11242 ( .A(n10311), .B(n10310), .Z(n10312) );
  AND U11243 ( .A(n10313), .B(n10312), .Z(n10436) );
  NAND U11244 ( .A(x[236]), .B(y[1895]), .Z(n10800) );
  NANDN U11245 ( .A(n10800), .B(n10314), .Z(n10318) );
  NANDN U11246 ( .A(n10316), .B(n10315), .Z(n10317) );
  AND U11247 ( .A(n10318), .B(n10317), .Z(n10412) );
  AND U11248 ( .A(y[1892]), .B(x[235]), .Z(n10320) );
  NAND U11249 ( .A(y[1890]), .B(x[237]), .Z(n10319) );
  XNOR U11250 ( .A(n10320), .B(n10319), .Z(n10416) );
  AND U11251 ( .A(x[236]), .B(y[1891]), .Z(n10415) );
  XOR U11252 ( .A(n10416), .B(n10415), .Z(n10410) );
  AND U11253 ( .A(y[1888]), .B(x[239]), .Z(n10322) );
  NAND U11254 ( .A(y[1903]), .B(x[224]), .Z(n10321) );
  XNOR U11255 ( .A(n10322), .B(n10321), .Z(n10378) );
  ANDN U11256 ( .B(o[110]), .A(n10323), .Z(n10377) );
  XNOR U11257 ( .A(n10378), .B(n10377), .Z(n10409) );
  XNOR U11258 ( .A(n10410), .B(n10409), .Z(n10411) );
  XOR U11259 ( .A(n10412), .B(n10411), .Z(n10444) );
  NAND U11260 ( .A(x[234]), .B(y[1900]), .Z(n11255) );
  NANDN U11261 ( .A(n11255), .B(n10324), .Z(n10327) );
  NAND U11262 ( .A(n10919), .B(n10325), .Z(n10326) );
  AND U11263 ( .A(n10327), .B(n10326), .Z(n10442) );
  AND U11264 ( .A(x[235]), .B(y[1896]), .Z(n10725) );
  NAND U11265 ( .A(n10725), .B(n10328), .Z(n10332) );
  NANDN U11266 ( .A(n10330), .B(n10329), .Z(n10331) );
  NAND U11267 ( .A(n10332), .B(n10331), .Z(n10441) );
  XNOR U11268 ( .A(n10442), .B(n10441), .Z(n10443) );
  XNOR U11269 ( .A(n10444), .B(n10443), .Z(n10435) );
  XNOR U11270 ( .A(n10436), .B(n10435), .Z(n10437) );
  XOR U11271 ( .A(n10438), .B(n10437), .Z(n10429) );
  AND U11272 ( .A(x[238]), .B(y[1902]), .Z(n12097) );
  AND U11273 ( .A(x[232]), .B(y[1899]), .Z(n10335) );
  NANDN U11274 ( .A(n10336), .B(n10335), .Z(n10339) );
  NANDN U11275 ( .A(n10337), .B(n10619), .Z(n10338) );
  NAND U11276 ( .A(n10339), .B(n10338), .Z(n10403) );
  XNOR U11277 ( .A(n10404), .B(n10403), .Z(n10406) );
  AND U11278 ( .A(y[1893]), .B(x[234]), .Z(n10341) );
  NAND U11279 ( .A(y[1899]), .B(x[228]), .Z(n10340) );
  XNOR U11280 ( .A(n10341), .B(n10340), .Z(n10384) );
  AND U11281 ( .A(x[231]), .B(y[1896]), .Z(n10383) );
  XOR U11282 ( .A(n10384), .B(n10383), .Z(n10391) );
  NAND U11283 ( .A(x[230]), .B(y[1897]), .Z(n10494) );
  XNOR U11284 ( .A(n10494), .B(n10389), .Z(n10390) );
  XOR U11285 ( .A(n10391), .B(n10390), .Z(n10425) );
  AND U11286 ( .A(y[1901]), .B(x[226]), .Z(n10343) );
  NAND U11287 ( .A(y[1894]), .B(x[233]), .Z(n10342) );
  XNOR U11288 ( .A(n10343), .B(n10342), .Z(n10394) );
  NAND U11289 ( .A(x[227]), .B(y[1900]), .Z(n10395) );
  XNOR U11290 ( .A(n10394), .B(n10395), .Z(n10423) );
  AND U11291 ( .A(y[1902]), .B(x[225]), .Z(n10345) );
  NAND U11292 ( .A(y[1895]), .B(x[232]), .Z(n10344) );
  XNOR U11293 ( .A(n10345), .B(n10344), .Z(n10372) );
  NAND U11294 ( .A(x[238]), .B(y[1889]), .Z(n10400) );
  XOR U11295 ( .A(o[111]), .B(n10400), .Z(n10373) );
  XNOR U11296 ( .A(n10372), .B(n10373), .Z(n10424) );
  XOR U11297 ( .A(n10423), .B(n10424), .Z(n10426) );
  XOR U11298 ( .A(n10425), .B(n10426), .Z(n10405) );
  XOR U11299 ( .A(n10406), .B(n10405), .Z(n10448) );
  XNOR U11300 ( .A(n10448), .B(n10447), .Z(n10450) );
  NANDN U11301 ( .A(n10350), .B(n10349), .Z(n10354) );
  NAND U11302 ( .A(n10352), .B(n10351), .Z(n10353) );
  AND U11303 ( .A(n10354), .B(n10353), .Z(n10449) );
  XOR U11304 ( .A(n10450), .B(n10449), .Z(n10430) );
  XNOR U11305 ( .A(n10429), .B(n10430), .Z(n10432) );
  NANDN U11306 ( .A(n10356), .B(n10355), .Z(n10360) );
  NAND U11307 ( .A(n10358), .B(n10357), .Z(n10359) );
  AND U11308 ( .A(n10360), .B(n10359), .Z(n10461) );
  XOR U11309 ( .A(n10460), .B(n10461), .Z(n10462) );
  XOR U11310 ( .A(n10463), .B(n10462), .Z(n10456) );
  NANDN U11311 ( .A(n10365), .B(n10364), .Z(n10369) );
  NAND U11312 ( .A(n10367), .B(n10366), .Z(n10368) );
  NAND U11313 ( .A(n10369), .B(n10368), .Z(n10454) );
  IV U11314 ( .A(n10454), .Z(n10453) );
  XOR U11315 ( .A(n10455), .B(n10453), .Z(n10370) );
  XNOR U11316 ( .A(n10456), .B(n10370), .Z(N240) );
  AND U11317 ( .A(x[232]), .B(y[1902]), .Z(n10726) );
  NAND U11318 ( .A(n10726), .B(n10371), .Z(n10375) );
  NANDN U11319 ( .A(n10373), .B(n10372), .Z(n10374) );
  NAND U11320 ( .A(n10375), .B(n10374), .Z(n10522) );
  AND U11321 ( .A(x[239]), .B(y[1903]), .Z(n12407) );
  NAND U11322 ( .A(n12407), .B(n10376), .Z(n10380) );
  NAND U11323 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND U11324 ( .A(n10380), .B(n10379), .Z(n10521) );
  XOR U11325 ( .A(n10522), .B(n10521), .Z(n10524) );
  AND U11326 ( .A(x[234]), .B(y[1899]), .Z(n10382) );
  NAND U11327 ( .A(n10382), .B(n10381), .Z(n10386) );
  NAND U11328 ( .A(n10384), .B(n10383), .Z(n10385) );
  NAND U11329 ( .A(n10386), .B(n10385), .Z(n10481) );
  AND U11330 ( .A(x[224]), .B(y[1904]), .Z(n10503) );
  AND U11331 ( .A(x[240]), .B(y[1888]), .Z(n10504) );
  XOR U11332 ( .A(n10503), .B(n10504), .Z(n10505) );
  NAND U11333 ( .A(x[239]), .B(y[1889]), .Z(n10491) );
  XNOR U11334 ( .A(o[112]), .B(n10491), .Z(n10506) );
  XOR U11335 ( .A(n10505), .B(n10506), .Z(n10480) );
  NAND U11336 ( .A(y[1897]), .B(x[231]), .Z(n10387) );
  XNOR U11337 ( .A(n10388), .B(n10387), .Z(n10496) );
  AND U11338 ( .A(x[234]), .B(y[1894]), .Z(n10495) );
  XOR U11339 ( .A(n10496), .B(n10495), .Z(n10479) );
  XOR U11340 ( .A(n10480), .B(n10479), .Z(n10482) );
  XOR U11341 ( .A(n10481), .B(n10482), .Z(n10523) );
  XOR U11342 ( .A(n10524), .B(n10523), .Z(n10476) );
  NANDN U11343 ( .A(n10389), .B(n10494), .Z(n10393) );
  NANDN U11344 ( .A(n10391), .B(n10390), .Z(n10392) );
  AND U11345 ( .A(n10393), .B(n10392), .Z(n10474) );
  NAND U11346 ( .A(x[233]), .B(y[1901]), .Z(n11236) );
  NANDN U11347 ( .A(n11236), .B(n10798), .Z(n10397) );
  NANDN U11348 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U11349 ( .A(n10397), .B(n10396), .Z(n10514) );
  AND U11350 ( .A(y[1903]), .B(x[225]), .Z(n10399) );
  NAND U11351 ( .A(y[1896]), .B(x[232]), .Z(n10398) );
  XNOR U11352 ( .A(n10399), .B(n10398), .Z(n10500) );
  ANDN U11353 ( .B(o[111]), .A(n10400), .Z(n10499) );
  XOR U11354 ( .A(n10500), .B(n10499), .Z(n10511) );
  NAND U11355 ( .A(y[1890]), .B(x[238]), .Z(n10401) );
  XNOR U11356 ( .A(n10402), .B(n10401), .Z(n10533) );
  NAND U11357 ( .A(x[228]), .B(y[1900]), .Z(n10534) );
  XNOR U11358 ( .A(n10533), .B(n10534), .Z(n10512) );
  XOR U11359 ( .A(n10511), .B(n10512), .Z(n10513) );
  XOR U11360 ( .A(n10514), .B(n10513), .Z(n10473) );
  XNOR U11361 ( .A(n10474), .B(n10473), .Z(n10475) );
  XNOR U11362 ( .A(n10476), .B(n10475), .Z(n10517) );
  NANDN U11363 ( .A(n10404), .B(n10403), .Z(n10408) );
  NAND U11364 ( .A(n10406), .B(n10405), .Z(n10407) );
  NAND U11365 ( .A(n10408), .B(n10407), .Z(n10518) );
  XNOR U11366 ( .A(n10517), .B(n10518), .Z(n10520) );
  NANDN U11367 ( .A(n10410), .B(n10409), .Z(n10414) );
  NAND U11368 ( .A(n10412), .B(n10411), .Z(n10413) );
  NAND U11369 ( .A(n10414), .B(n10413), .Z(n10548) );
  AND U11370 ( .A(x[237]), .B(y[1892]), .Z(n10544) );
  NAND U11371 ( .A(n11056), .B(n10544), .Z(n10418) );
  NAND U11372 ( .A(n10416), .B(n10415), .Z(n10417) );
  NAND U11373 ( .A(n10418), .B(n10417), .Z(n10530) );
  AND U11374 ( .A(y[1902]), .B(x[226]), .Z(n10420) );
  NAND U11375 ( .A(y[1895]), .B(x[233]), .Z(n10419) );
  XNOR U11376 ( .A(n10420), .B(n10419), .Z(n10538) );
  NAND U11377 ( .A(x[227]), .B(y[1901]), .Z(n10539) );
  XNOR U11378 ( .A(n10538), .B(n10539), .Z(n10527) );
  AND U11379 ( .A(x[236]), .B(y[1892]), .Z(n11224) );
  AND U11380 ( .A(y[1899]), .B(x[229]), .Z(n10422) );
  NAND U11381 ( .A(y[1891]), .B(x[237]), .Z(n10421) );
  XOR U11382 ( .A(n10422), .B(n10421), .Z(n10486) );
  XNOR U11383 ( .A(n11224), .B(n10486), .Z(n10528) );
  XOR U11384 ( .A(n10527), .B(n10528), .Z(n10529) );
  XNOR U11385 ( .A(n10530), .B(n10529), .Z(n10545) );
  NAND U11386 ( .A(n10424), .B(n10423), .Z(n10428) );
  NAND U11387 ( .A(n10426), .B(n10425), .Z(n10427) );
  AND U11388 ( .A(n10428), .B(n10427), .Z(n10546) );
  XOR U11389 ( .A(n10545), .B(n10546), .Z(n10547) );
  XOR U11390 ( .A(n10548), .B(n10547), .Z(n10519) );
  XOR U11391 ( .A(n10520), .B(n10519), .Z(n10552) );
  NAND U11392 ( .A(n10430), .B(n10429), .Z(n10434) );
  NANDN U11393 ( .A(n10432), .B(n10431), .Z(n10433) );
  AND U11394 ( .A(n10434), .B(n10433), .Z(n10551) );
  NANDN U11395 ( .A(n10436), .B(n10435), .Z(n10440) );
  NANDN U11396 ( .A(n10438), .B(n10437), .Z(n10439) );
  AND U11397 ( .A(n10440), .B(n10439), .Z(n10470) );
  NANDN U11398 ( .A(n10442), .B(n10441), .Z(n10446) );
  NANDN U11399 ( .A(n10444), .B(n10443), .Z(n10445) );
  AND U11400 ( .A(n10446), .B(n10445), .Z(n10468) );
  NANDN U11401 ( .A(n10448), .B(n10447), .Z(n10452) );
  NAND U11402 ( .A(n10450), .B(n10449), .Z(n10451) );
  AND U11403 ( .A(n10452), .B(n10451), .Z(n10467) );
  XNOR U11404 ( .A(n10468), .B(n10467), .Z(n10469) );
  XNOR U11405 ( .A(n10470), .B(n10469), .Z(n10553) );
  XNOR U11406 ( .A(n10554), .B(n10553), .Z(n10560) );
  OR U11407 ( .A(n10455), .B(n10453), .Z(n10459) );
  ANDN U11408 ( .B(n10455), .A(n10454), .Z(n10457) );
  OR U11409 ( .A(n10457), .B(n10456), .Z(n10458) );
  AND U11410 ( .A(n10459), .B(n10458), .Z(n10559) );
  NAND U11411 ( .A(n10461), .B(n10460), .Z(n10465) );
  NANDN U11412 ( .A(n10463), .B(n10462), .Z(n10464) );
  NAND U11413 ( .A(n10465), .B(n10464), .Z(n10558) );
  IV U11414 ( .A(n10558), .Z(n10557) );
  XOR U11415 ( .A(n10559), .B(n10557), .Z(n10466) );
  XNOR U11416 ( .A(n10560), .B(n10466), .Z(N241) );
  NANDN U11417 ( .A(n10468), .B(n10467), .Z(n10472) );
  NANDN U11418 ( .A(n10470), .B(n10469), .Z(n10471) );
  AND U11419 ( .A(n10472), .B(n10471), .Z(n10662) );
  NANDN U11420 ( .A(n10474), .B(n10473), .Z(n10478) );
  NANDN U11421 ( .A(n10476), .B(n10475), .Z(n10477) );
  NAND U11422 ( .A(n10478), .B(n10477), .Z(n10574) );
  NAND U11423 ( .A(n10480), .B(n10479), .Z(n10484) );
  NAND U11424 ( .A(n10482), .B(n10481), .Z(n10483) );
  NAND U11425 ( .A(n10484), .B(n10483), .Z(n10656) );
  AND U11426 ( .A(x[237]), .B(y[1899]), .Z(n11501) );
  NAND U11427 ( .A(n11501), .B(n10485), .Z(n10488) );
  NANDN U11428 ( .A(n10486), .B(n11224), .Z(n10487) );
  NAND U11429 ( .A(n10488), .B(n10487), .Z(n10604) );
  AND U11430 ( .A(y[1904]), .B(x[225]), .Z(n10490) );
  NAND U11431 ( .A(y[1896]), .B(x[233]), .Z(n10489) );
  XNOR U11432 ( .A(n10490), .B(n10489), .Z(n10624) );
  NANDN U11433 ( .A(n10491), .B(o[112]), .Z(n10625) );
  XNOR U11434 ( .A(n10624), .B(n10625), .Z(n10602) );
  AND U11435 ( .A(y[1890]), .B(x[239]), .Z(n10493) );
  NAND U11436 ( .A(y[1893]), .B(x[236]), .Z(n10492) );
  XNOR U11437 ( .A(n10493), .B(n10492), .Z(n10578) );
  AND U11438 ( .A(x[238]), .B(y[1891]), .Z(n10577) );
  XOR U11439 ( .A(n10578), .B(n10577), .Z(n10601) );
  XOR U11440 ( .A(n10602), .B(n10601), .Z(n10603) );
  XOR U11441 ( .A(n10604), .B(n10603), .Z(n10654) );
  AND U11442 ( .A(x[231]), .B(y[1898]), .Z(n10636) );
  NANDN U11443 ( .A(n10494), .B(n10636), .Z(n10498) );
  NAND U11444 ( .A(n10496), .B(n10495), .Z(n10497) );
  NAND U11445 ( .A(n10498), .B(n10497), .Z(n10614) );
  AND U11446 ( .A(x[225]), .B(y[1896]), .Z(n10705) );
  AND U11447 ( .A(x[232]), .B(y[1903]), .Z(n11303) );
  NAND U11448 ( .A(n10705), .B(n11303), .Z(n10502) );
  NAND U11449 ( .A(n10500), .B(n10499), .Z(n10501) );
  NAND U11450 ( .A(n10502), .B(n10501), .Z(n10613) );
  XOR U11451 ( .A(n10614), .B(n10613), .Z(n10616) );
  NAND U11452 ( .A(n10504), .B(n10503), .Z(n10508) );
  NAND U11453 ( .A(n10506), .B(n10505), .Z(n10507) );
  NAND U11454 ( .A(n10508), .B(n10507), .Z(n10610) );
  AND U11455 ( .A(x[224]), .B(y[1905]), .Z(n10592) );
  AND U11456 ( .A(x[241]), .B(y[1888]), .Z(n10591) );
  XOR U11457 ( .A(n10592), .B(n10591), .Z(n10594) );
  AND U11458 ( .A(x[240]), .B(y[1889]), .Z(n10588) );
  XOR U11459 ( .A(n10588), .B(o[113]), .Z(n10593) );
  XOR U11460 ( .A(n10594), .B(n10593), .Z(n10607) );
  AND U11461 ( .A(y[1903]), .B(x[226]), .Z(n10510) );
  NAND U11462 ( .A(y[1895]), .B(x[234]), .Z(n10509) );
  XNOR U11463 ( .A(n10510), .B(n10509), .Z(n10629) );
  NAND U11464 ( .A(x[227]), .B(y[1902]), .Z(n10630) );
  XNOR U11465 ( .A(n10629), .B(n10630), .Z(n10608) );
  XOR U11466 ( .A(n10607), .B(n10608), .Z(n10609) );
  XOR U11467 ( .A(n10610), .B(n10609), .Z(n10615) );
  XOR U11468 ( .A(n10616), .B(n10615), .Z(n10653) );
  XOR U11469 ( .A(n10654), .B(n10653), .Z(n10655) );
  XNOR U11470 ( .A(n10656), .B(n10655), .Z(n10571) );
  NAND U11471 ( .A(n10512), .B(n10511), .Z(n10516) );
  NANDN U11472 ( .A(n10514), .B(n10513), .Z(n10515) );
  AND U11473 ( .A(n10516), .B(n10515), .Z(n10572) );
  XOR U11474 ( .A(n10571), .B(n10572), .Z(n10573) );
  XNOR U11475 ( .A(n10574), .B(n10573), .Z(n10660) );
  NAND U11476 ( .A(n10522), .B(n10521), .Z(n10526) );
  NAND U11477 ( .A(n10524), .B(n10523), .Z(n10525) );
  NAND U11478 ( .A(n10526), .B(n10525), .Z(n10650) );
  NAND U11479 ( .A(n10528), .B(n10527), .Z(n10532) );
  NAND U11480 ( .A(n10530), .B(n10529), .Z(n10531) );
  NAND U11481 ( .A(n10532), .B(n10531), .Z(n10648) );
  NAND U11482 ( .A(x[238]), .B(y[1893]), .Z(n10845) );
  NANDN U11483 ( .A(n10845), .B(n11056), .Z(n10536) );
  NANDN U11484 ( .A(n10534), .B(n10533), .Z(n10535) );
  AND U11485 ( .A(n10536), .B(n10535), .Z(n10642) );
  AND U11486 ( .A(x[233]), .B(y[1902]), .Z(n11482) );
  NANDN U11487 ( .A(n10537), .B(n11482), .Z(n10541) );
  NANDN U11488 ( .A(n10539), .B(n10538), .Z(n10540) );
  NAND U11489 ( .A(n10541), .B(n10540), .Z(n10641) );
  XNOR U11490 ( .A(n10642), .B(n10641), .Z(n10643) );
  AND U11491 ( .A(x[229]), .B(y[1900]), .Z(n10687) );
  NAND U11492 ( .A(y[1897]), .B(x[232]), .Z(n10542) );
  XNOR U11493 ( .A(n10687), .B(n10542), .Z(n10621) );
  XOR U11494 ( .A(n10621), .B(n10620), .Z(n10635) );
  XOR U11495 ( .A(n10635), .B(n10636), .Z(n10637) );
  NAND U11496 ( .A(y[1901]), .B(x[228]), .Z(n10543) );
  XNOR U11497 ( .A(n10544), .B(n10543), .Z(n10582) );
  NAND U11498 ( .A(x[235]), .B(y[1894]), .Z(n10583) );
  XOR U11499 ( .A(n10582), .B(n10583), .Z(n10638) );
  XOR U11500 ( .A(n10637), .B(n10638), .Z(n10644) );
  XNOR U11501 ( .A(n10643), .B(n10644), .Z(n10647) );
  XOR U11502 ( .A(n10648), .B(n10647), .Z(n10649) );
  XNOR U11503 ( .A(n10650), .B(n10649), .Z(n10566) );
  NAND U11504 ( .A(n10546), .B(n10545), .Z(n10550) );
  NAND U11505 ( .A(n10548), .B(n10547), .Z(n10549) );
  NAND U11506 ( .A(n10550), .B(n10549), .Z(n10565) );
  XOR U11507 ( .A(n10566), .B(n10565), .Z(n10567) );
  XOR U11508 ( .A(n10568), .B(n10567), .Z(n10659) );
  XOR U11509 ( .A(n10660), .B(n10659), .Z(n10661) );
  XNOR U11510 ( .A(n10662), .B(n10661), .Z(n10667) );
  NANDN U11511 ( .A(n10552), .B(n10551), .Z(n10556) );
  NAND U11512 ( .A(n10554), .B(n10553), .Z(n10555) );
  AND U11513 ( .A(n10556), .B(n10555), .Z(n10666) );
  OR U11514 ( .A(n10559), .B(n10557), .Z(n10563) );
  ANDN U11515 ( .B(n10559), .A(n10558), .Z(n10561) );
  OR U11516 ( .A(n10561), .B(n10560), .Z(n10562) );
  AND U11517 ( .A(n10563), .B(n10562), .Z(n10665) );
  XNOR U11518 ( .A(n10666), .B(n10665), .Z(n10564) );
  XNOR U11519 ( .A(n10667), .B(n10564), .Z(N242) );
  NAND U11520 ( .A(n10566), .B(n10565), .Z(n10570) );
  NANDN U11521 ( .A(n10568), .B(n10567), .Z(n10569) );
  AND U11522 ( .A(n10570), .B(n10569), .Z(n10777) );
  NAND U11523 ( .A(n10572), .B(n10571), .Z(n10576) );
  NAND U11524 ( .A(n10574), .B(n10573), .Z(n10575) );
  AND U11525 ( .A(n10576), .B(n10575), .Z(n10775) );
  AND U11526 ( .A(x[236]), .B(y[1890]), .Z(n10909) );
  AND U11527 ( .A(x[239]), .B(y[1893]), .Z(n10806) );
  NAND U11528 ( .A(n10909), .B(n10806), .Z(n10580) );
  NAND U11529 ( .A(n10578), .B(n10577), .Z(n10579) );
  NAND U11530 ( .A(n10580), .B(n10579), .Z(n10753) );
  NAND U11531 ( .A(n11744), .B(n10581), .Z(n10585) );
  NANDN U11532 ( .A(n10583), .B(n10582), .Z(n10584) );
  AND U11533 ( .A(n10585), .B(n10584), .Z(n10744) );
  AND U11534 ( .A(y[1905]), .B(x[225]), .Z(n10587) );
  NAND U11535 ( .A(y[1896]), .B(x[234]), .Z(n10586) );
  XNOR U11536 ( .A(n10587), .B(n10586), .Z(n10706) );
  NAND U11537 ( .A(n10588), .B(o[113]), .Z(n10707) );
  XNOR U11538 ( .A(n10706), .B(n10707), .Z(n10741) );
  AND U11539 ( .A(y[1891]), .B(x[239]), .Z(n10590) );
  NAND U11540 ( .A(y[1897]), .B(x[233]), .Z(n10589) );
  XNOR U11541 ( .A(n10590), .B(n10589), .Z(n10697) );
  NAND U11542 ( .A(x[238]), .B(y[1892]), .Z(n10698) );
  XOR U11543 ( .A(n10697), .B(n10698), .Z(n10742) );
  XNOR U11544 ( .A(n10741), .B(n10742), .Z(n10743) );
  XNOR U11545 ( .A(n10744), .B(n10743), .Z(n10754) );
  XOR U11546 ( .A(n10753), .B(n10754), .Z(n10756) );
  NAND U11547 ( .A(n10592), .B(n10591), .Z(n10596) );
  NAND U11548 ( .A(n10594), .B(n10593), .Z(n10595) );
  NAND U11549 ( .A(n10596), .B(n10595), .Z(n10765) );
  AND U11550 ( .A(y[1890]), .B(x[240]), .Z(n10598) );
  NAND U11551 ( .A(y[1895]), .B(x[235]), .Z(n10597) );
  XNOR U11552 ( .A(n10598), .B(n10597), .Z(n10693) );
  NAND U11553 ( .A(x[226]), .B(y[1904]), .Z(n10694) );
  XNOR U11554 ( .A(n10693), .B(n10694), .Z(n10766) );
  XOR U11555 ( .A(n10765), .B(n10766), .Z(n10768) );
  AND U11556 ( .A(x[229]), .B(y[1901]), .Z(n10826) );
  NAND U11557 ( .A(y[1900]), .B(x[230]), .Z(n10599) );
  XNOR U11558 ( .A(n10826), .B(n10599), .Z(n10690) );
  NAND U11559 ( .A(y[1902]), .B(x[228]), .Z(n10600) );
  XNOR U11560 ( .A(n11487), .B(n10600), .Z(n10728) );
  NAND U11561 ( .A(x[231]), .B(y[1899]), .Z(n10729) );
  XOR U11562 ( .A(n10690), .B(n10689), .Z(n10767) );
  XOR U11563 ( .A(n10768), .B(n10767), .Z(n10755) );
  XNOR U11564 ( .A(n10756), .B(n10755), .Z(n10676) );
  NAND U11565 ( .A(n10602), .B(n10601), .Z(n10606) );
  NAND U11566 ( .A(n10604), .B(n10603), .Z(n10605) );
  AND U11567 ( .A(n10606), .B(n10605), .Z(n10748) );
  NAND U11568 ( .A(n10608), .B(n10607), .Z(n10612) );
  NAND U11569 ( .A(n10610), .B(n10609), .Z(n10611) );
  AND U11570 ( .A(n10612), .B(n10611), .Z(n10747) );
  XOR U11571 ( .A(n10748), .B(n10747), .Z(n10750) );
  NAND U11572 ( .A(n10614), .B(n10613), .Z(n10618) );
  NAND U11573 ( .A(n10616), .B(n10615), .Z(n10617) );
  AND U11574 ( .A(n10618), .B(n10617), .Z(n10749) );
  XOR U11575 ( .A(n10750), .B(n10749), .Z(n10675) );
  XOR U11576 ( .A(n10676), .B(n10675), .Z(n10678) );
  AND U11577 ( .A(x[232]), .B(y[1900]), .Z(n10955) );
  NAND U11578 ( .A(n10955), .B(n10619), .Z(n10623) );
  NAND U11579 ( .A(n10621), .B(n10620), .Z(n10622) );
  NAND U11580 ( .A(n10623), .B(n10622), .Z(n10760) );
  NAND U11581 ( .A(x[233]), .B(y[1904]), .Z(n11603) );
  NANDN U11582 ( .A(n11603), .B(n10705), .Z(n10627) );
  NANDN U11583 ( .A(n10625), .B(n10624), .Z(n10626) );
  NAND U11584 ( .A(n10627), .B(n10626), .Z(n10759) );
  XOR U11585 ( .A(n10760), .B(n10759), .Z(n10762) );
  NAND U11586 ( .A(x[234]), .B(y[1903]), .Z(n11604) );
  NANDN U11587 ( .A(n11604), .B(n10628), .Z(n10632) );
  NANDN U11588 ( .A(n10630), .B(n10629), .Z(n10631) );
  AND U11589 ( .A(n10632), .B(n10631), .Z(n10738) );
  AND U11590 ( .A(x[224]), .B(y[1906]), .Z(n10710) );
  NAND U11591 ( .A(x[242]), .B(y[1888]), .Z(n10711) );
  XNOR U11592 ( .A(n10710), .B(n10711), .Z(n10712) );
  NAND U11593 ( .A(x[241]), .B(y[1889]), .Z(n10732) );
  XOR U11594 ( .A(o[114]), .B(n10732), .Z(n10713) );
  XNOR U11595 ( .A(n10712), .B(n10713), .Z(n10735) );
  AND U11596 ( .A(y[1893]), .B(x[237]), .Z(n10634) );
  NAND U11597 ( .A(y[1903]), .B(x[227]), .Z(n10633) );
  XNOR U11598 ( .A(n10634), .B(n10633), .Z(n10718) );
  NAND U11599 ( .A(x[236]), .B(y[1894]), .Z(n10719) );
  XOR U11600 ( .A(n10718), .B(n10719), .Z(n10736) );
  XNOR U11601 ( .A(n10735), .B(n10736), .Z(n10737) );
  XNOR U11602 ( .A(n10738), .B(n10737), .Z(n10761) );
  XOR U11603 ( .A(n10762), .B(n10761), .Z(n10682) );
  NAND U11604 ( .A(n10636), .B(n10635), .Z(n10640) );
  NANDN U11605 ( .A(n10638), .B(n10637), .Z(n10639) );
  AND U11606 ( .A(n10640), .B(n10639), .Z(n10681) );
  XNOR U11607 ( .A(n10682), .B(n10681), .Z(n10683) );
  NANDN U11608 ( .A(n10642), .B(n10641), .Z(n10646) );
  NANDN U11609 ( .A(n10644), .B(n10643), .Z(n10645) );
  NAND U11610 ( .A(n10646), .B(n10645), .Z(n10684) );
  XNOR U11611 ( .A(n10683), .B(n10684), .Z(n10677) );
  XNOR U11612 ( .A(n10678), .B(n10677), .Z(n10672) );
  NAND U11613 ( .A(n10648), .B(n10647), .Z(n10652) );
  NAND U11614 ( .A(n10650), .B(n10649), .Z(n10651) );
  NAND U11615 ( .A(n10652), .B(n10651), .Z(n10670) );
  NAND U11616 ( .A(n10654), .B(n10653), .Z(n10658) );
  NAND U11617 ( .A(n10656), .B(n10655), .Z(n10657) );
  NAND U11618 ( .A(n10658), .B(n10657), .Z(n10669) );
  XOR U11619 ( .A(n10670), .B(n10669), .Z(n10671) );
  XOR U11620 ( .A(n10672), .B(n10671), .Z(n10774) );
  XOR U11621 ( .A(n10775), .B(n10774), .Z(n10776) );
  XNOR U11622 ( .A(n10777), .B(n10776), .Z(n10773) );
  NAND U11623 ( .A(n10660), .B(n10659), .Z(n10664) );
  NANDN U11624 ( .A(n10662), .B(n10661), .Z(n10663) );
  NAND U11625 ( .A(n10664), .B(n10663), .Z(n10771) );
  XOR U11626 ( .A(n10771), .B(n10772), .Z(n10668) );
  XNOR U11627 ( .A(n10773), .B(n10668), .Z(N243) );
  NAND U11628 ( .A(n10670), .B(n10669), .Z(n10674) );
  NAND U11629 ( .A(n10672), .B(n10671), .Z(n10673) );
  NAND U11630 ( .A(n10674), .B(n10673), .Z(n10892) );
  NAND U11631 ( .A(n10676), .B(n10675), .Z(n10680) );
  NAND U11632 ( .A(n10678), .B(n10677), .Z(n10679) );
  AND U11633 ( .A(n10680), .B(n10679), .Z(n10890) );
  NANDN U11634 ( .A(n10682), .B(n10681), .Z(n10686) );
  NANDN U11635 ( .A(n10684), .B(n10683), .Z(n10685) );
  AND U11636 ( .A(n10686), .B(n10685), .Z(n10874) );
  AND U11637 ( .A(x[230]), .B(y[1901]), .Z(n10688) );
  NAND U11638 ( .A(n10688), .B(n10687), .Z(n10692) );
  NAND U11639 ( .A(n10690), .B(n10689), .Z(n10691) );
  AND U11640 ( .A(n10692), .B(n10691), .Z(n10867) );
  AND U11641 ( .A(x[240]), .B(y[1895]), .Z(n11240) );
  NAND U11642 ( .A(n11056), .B(n11240), .Z(n10696) );
  NANDN U11643 ( .A(n10694), .B(n10693), .Z(n10695) );
  AND U11644 ( .A(n10696), .B(n10695), .Z(n10866) );
  AND U11645 ( .A(x[239]), .B(y[1897]), .Z(n11518) );
  NAND U11646 ( .A(n10793), .B(n11518), .Z(n10700) );
  NANDN U11647 ( .A(n10698), .B(n10697), .Z(n10699) );
  AND U11648 ( .A(n10700), .B(n10699), .Z(n10784) );
  AND U11649 ( .A(y[1906]), .B(x[225]), .Z(n10702) );
  NAND U11650 ( .A(y[1899]), .B(x[232]), .Z(n10701) );
  XNOR U11651 ( .A(n10702), .B(n10701), .Z(n10844) );
  AND U11652 ( .A(y[1894]), .B(x[237]), .Z(n10704) );
  NAND U11653 ( .A(y[1905]), .B(x[226]), .Z(n10703) );
  XNOR U11654 ( .A(n10704), .B(n10703), .Z(n10799) );
  XOR U11655 ( .A(n10782), .B(n10781), .Z(n10783) );
  XOR U11656 ( .A(n10866), .B(n10865), .Z(n10868) );
  XOR U11657 ( .A(n10867), .B(n10868), .Z(n10872) );
  AND U11658 ( .A(x[234]), .B(y[1905]), .Z(n11918) );
  IV U11659 ( .A(n11918), .Z(n11841) );
  NANDN U11660 ( .A(n11841), .B(n10705), .Z(n10709) );
  NANDN U11661 ( .A(n10707), .B(n10706), .Z(n10708) );
  AND U11662 ( .A(n10709), .B(n10708), .Z(n10823) );
  NANDN U11663 ( .A(n10711), .B(n10710), .Z(n10715) );
  NANDN U11664 ( .A(n10713), .B(n10712), .Z(n10714) );
  AND U11665 ( .A(n10715), .B(n10714), .Z(n10821) );
  AND U11666 ( .A(y[1891]), .B(x[240]), .Z(n11455) );
  NAND U11667 ( .A(y[1898]), .B(x[233]), .Z(n10716) );
  XNOR U11668 ( .A(n11455), .B(n10716), .Z(n10794) );
  NAND U11669 ( .A(x[239]), .B(y[1892]), .Z(n10795) );
  AND U11670 ( .A(x[237]), .B(y[1903]), .Z(n12125) );
  NANDN U11671 ( .A(n10717), .B(n12125), .Z(n10721) );
  NANDN U11672 ( .A(n10719), .B(n10718), .Z(n10720) );
  AND U11673 ( .A(n10721), .B(n10720), .Z(n10817) );
  AND U11674 ( .A(y[1897]), .B(x[234]), .Z(n10723) );
  NAND U11675 ( .A(y[1890]), .B(x[241]), .Z(n10722) );
  XNOR U11676 ( .A(n10723), .B(n10722), .Z(n10850) );
  AND U11677 ( .A(x[242]), .B(y[1889]), .Z(n10813) );
  XOR U11678 ( .A(o[115]), .B(n10813), .Z(n10849) );
  XOR U11679 ( .A(n10850), .B(n10849), .Z(n10815) );
  NAND U11680 ( .A(y[1904]), .B(x[227]), .Z(n10724) );
  XNOR U11681 ( .A(n10725), .B(n10724), .Z(n10807) );
  XOR U11682 ( .A(n10815), .B(n10814), .Z(n10816) );
  NAND U11683 ( .A(n10727), .B(n10726), .Z(n10731) );
  NANDN U11684 ( .A(n10729), .B(n10728), .Z(n10730) );
  AND U11685 ( .A(n10731), .B(n10730), .Z(n10790) );
  AND U11686 ( .A(x[224]), .B(y[1907]), .Z(n10830) );
  NAND U11687 ( .A(x[243]), .B(y[1888]), .Z(n10831) );
  ANDN U11688 ( .B(o[114]), .A(n10732), .Z(n10832) );
  XOR U11689 ( .A(n10833), .B(n10832), .Z(n10788) );
  AND U11690 ( .A(x[228]), .B(y[1903]), .Z(n10975) );
  AND U11691 ( .A(y[1902]), .B(x[229]), .Z(n10734) );
  NAND U11692 ( .A(y[1901]), .B(x[230]), .Z(n10733) );
  XOR U11693 ( .A(n10734), .B(n10733), .Z(n10827) );
  XOR U11694 ( .A(n10788), .B(n10787), .Z(n10789) );
  XOR U11695 ( .A(n10790), .B(n10789), .Z(n10859) );
  XNOR U11696 ( .A(n10860), .B(n10859), .Z(n10862) );
  XOR U11697 ( .A(n10861), .B(n10862), .Z(n10855) );
  NANDN U11698 ( .A(n10736), .B(n10735), .Z(n10740) );
  NANDN U11699 ( .A(n10738), .B(n10737), .Z(n10739) );
  AND U11700 ( .A(n10740), .B(n10739), .Z(n10854) );
  NANDN U11701 ( .A(n10742), .B(n10741), .Z(n10746) );
  NANDN U11702 ( .A(n10744), .B(n10743), .Z(n10745) );
  NAND U11703 ( .A(n10746), .B(n10745), .Z(n10853) );
  XOR U11704 ( .A(n10854), .B(n10853), .Z(n10856) );
  XOR U11705 ( .A(n10855), .B(n10856), .Z(n10871) );
  XNOR U11706 ( .A(n10872), .B(n10871), .Z(n10873) );
  XOR U11707 ( .A(n10874), .B(n10873), .Z(n10885) );
  NAND U11708 ( .A(n10748), .B(n10747), .Z(n10752) );
  NAND U11709 ( .A(n10750), .B(n10749), .Z(n10751) );
  AND U11710 ( .A(n10752), .B(n10751), .Z(n10883) );
  NAND U11711 ( .A(n10754), .B(n10753), .Z(n10758) );
  NAND U11712 ( .A(n10756), .B(n10755), .Z(n10757) );
  NAND U11713 ( .A(n10758), .B(n10757), .Z(n10879) );
  NAND U11714 ( .A(n10760), .B(n10759), .Z(n10764) );
  NAND U11715 ( .A(n10762), .B(n10761), .Z(n10763) );
  NAND U11716 ( .A(n10764), .B(n10763), .Z(n10878) );
  NAND U11717 ( .A(n10766), .B(n10765), .Z(n10770) );
  NAND U11718 ( .A(n10768), .B(n10767), .Z(n10769) );
  NAND U11719 ( .A(n10770), .B(n10769), .Z(n10877) );
  XNOR U11720 ( .A(n10878), .B(n10877), .Z(n10880) );
  XNOR U11721 ( .A(n10883), .B(n10884), .Z(n10886) );
  XOR U11722 ( .A(n10885), .B(n10886), .Z(n10889) );
  XOR U11723 ( .A(n10890), .B(n10889), .Z(n10891) );
  XOR U11724 ( .A(n10892), .B(n10891), .Z(n10898) );
  NAND U11725 ( .A(n10775), .B(n10774), .Z(n10779) );
  NAND U11726 ( .A(n10777), .B(n10776), .Z(n10778) );
  AND U11727 ( .A(n10779), .B(n10778), .Z(n10897) );
  IV U11728 ( .A(n10897), .Z(n10895) );
  XOR U11729 ( .A(n10896), .B(n10895), .Z(n10780) );
  XNOR U11730 ( .A(n10898), .B(n10780), .Z(N244) );
  NAND U11731 ( .A(n10782), .B(n10781), .Z(n10786) );
  NANDN U11732 ( .A(n10784), .B(n10783), .Z(n10785) );
  AND U11733 ( .A(n10786), .B(n10785), .Z(n10904) );
  NAND U11734 ( .A(n10788), .B(n10787), .Z(n10792) );
  NANDN U11735 ( .A(n10790), .B(n10789), .Z(n10791) );
  NAND U11736 ( .A(n10792), .B(n10791), .Z(n10903) );
  AND U11737 ( .A(x[240]), .B(y[1898]), .Z(n11799) );
  NAND U11738 ( .A(n11799), .B(n10793), .Z(n10797) );
  NANDN U11739 ( .A(n10795), .B(n10794), .Z(n10796) );
  AND U11740 ( .A(n10797), .B(n10796), .Z(n10944) );
  AND U11741 ( .A(x[237]), .B(y[1905]), .Z(n12365) );
  NAND U11742 ( .A(n12365), .B(n10798), .Z(n10802) );
  NANDN U11743 ( .A(n10800), .B(n10799), .Z(n10801) );
  AND U11744 ( .A(n10802), .B(n10801), .Z(n10989) );
  AND U11745 ( .A(y[1892]), .B(x[240]), .Z(n10804) );
  NAND U11746 ( .A(y[1898]), .B(x[234]), .Z(n10803) );
  XNOR U11747 ( .A(n10804), .B(n10803), .Z(n10950) );
  AND U11748 ( .A(x[226]), .B(y[1906]), .Z(n10951) );
  XOR U11749 ( .A(n10950), .B(n10951), .Z(n10987) );
  NAND U11750 ( .A(y[1899]), .B(x[233]), .Z(n10805) );
  XNOR U11751 ( .A(n10806), .B(n10805), .Z(n10920) );
  AND U11752 ( .A(x[238]), .B(y[1894]), .Z(n10921) );
  XOR U11753 ( .A(n10920), .B(n10921), .Z(n10986) );
  XOR U11754 ( .A(n10987), .B(n10986), .Z(n10988) );
  NAND U11755 ( .A(x[235]), .B(y[1904]), .Z(n11919) );
  NANDN U11756 ( .A(n11919), .B(n11083), .Z(n10810) );
  NANDN U11757 ( .A(n10808), .B(n10807), .Z(n10809) );
  AND U11758 ( .A(n10810), .B(n10809), .Z(n10995) );
  AND U11759 ( .A(y[1897]), .B(x[235]), .Z(n10812) );
  NAND U11760 ( .A(y[1907]), .B(x[225]), .Z(n10811) );
  XNOR U11761 ( .A(n10812), .B(n10811), .Z(n10916) );
  AND U11762 ( .A(x[243]), .B(y[1889]), .Z(n10924) );
  XOR U11763 ( .A(o[116]), .B(n10924), .Z(n10915) );
  XOR U11764 ( .A(n10916), .B(n10915), .Z(n10993) );
  AND U11765 ( .A(o[115]), .B(n10813), .Z(n10972) );
  AND U11766 ( .A(x[224]), .B(y[1908]), .Z(n10969) );
  AND U11767 ( .A(x[244]), .B(y[1888]), .Z(n10970) );
  XOR U11768 ( .A(n10969), .B(n10970), .Z(n10971) );
  XOR U11769 ( .A(n10972), .B(n10971), .Z(n10992) );
  XOR U11770 ( .A(n10993), .B(n10992), .Z(n10994) );
  XOR U11771 ( .A(n10946), .B(n10945), .Z(n10905) );
  XOR U11772 ( .A(n10906), .B(n10905), .Z(n11001) );
  NAND U11773 ( .A(n10815), .B(n10814), .Z(n10819) );
  NANDN U11774 ( .A(n10817), .B(n10816), .Z(n10818) );
  AND U11775 ( .A(n10819), .B(n10818), .Z(n10999) );
  NANDN U11776 ( .A(n10821), .B(n10820), .Z(n10825) );
  NANDN U11777 ( .A(n10823), .B(n10822), .Z(n10824) );
  AND U11778 ( .A(n10825), .B(n10824), .Z(n10940) );
  AND U11779 ( .A(x[230]), .B(y[1902]), .Z(n10926) );
  IV U11780 ( .A(n10926), .Z(n10842) );
  NANDN U11781 ( .A(n10842), .B(n10826), .Z(n10829) );
  NANDN U11782 ( .A(n10827), .B(n10975), .Z(n10828) );
  AND U11783 ( .A(n10829), .B(n10828), .Z(n10934) );
  NANDN U11784 ( .A(n10831), .B(n10830), .Z(n10835) );
  NAND U11785 ( .A(n10833), .B(n10832), .Z(n10834) );
  AND U11786 ( .A(n10835), .B(n10834), .Z(n10932) );
  AND U11787 ( .A(y[1890]), .B(x[242]), .Z(n10837) );
  NAND U11788 ( .A(y[1896]), .B(x[236]), .Z(n10836) );
  XNOR U11789 ( .A(n10837), .B(n10836), .Z(n10910) );
  AND U11790 ( .A(x[241]), .B(y[1891]), .Z(n10911) );
  XOR U11791 ( .A(n10910), .B(n10911), .Z(n10931) );
  AND U11792 ( .A(y[1895]), .B(x[237]), .Z(n10839) );
  NAND U11793 ( .A(y[1905]), .B(x[227]), .Z(n10838) );
  XNOR U11794 ( .A(n10839), .B(n10838), .Z(n10956) );
  XOR U11795 ( .A(n10956), .B(n10955), .Z(n10928) );
  AND U11796 ( .A(y[1903]), .B(x[229]), .Z(n10841) );
  NAND U11797 ( .A(y[1904]), .B(x[228]), .Z(n10840) );
  XNOR U11798 ( .A(n10841), .B(n10840), .Z(n10977) );
  AND U11799 ( .A(x[231]), .B(y[1901]), .Z(n10976) );
  XNOR U11800 ( .A(n10977), .B(n10976), .Z(n10925) );
  XOR U11801 ( .A(n10842), .B(n10925), .Z(n10927) );
  AND U11802 ( .A(x[232]), .B(y[1906]), .Z(n12077) );
  AND U11803 ( .A(x[225]), .B(y[1899]), .Z(n10843) );
  NAND U11804 ( .A(n12077), .B(n10843), .Z(n10847) );
  NANDN U11805 ( .A(n10845), .B(n10844), .Z(n10846) );
  AND U11806 ( .A(n10847), .B(n10846), .Z(n10981) );
  AND U11807 ( .A(x[241]), .B(y[1897]), .Z(n11807) );
  NAND U11808 ( .A(n11807), .B(n10848), .Z(n10852) );
  NAND U11809 ( .A(n10850), .B(n10849), .Z(n10851) );
  NAND U11810 ( .A(n10852), .B(n10851), .Z(n10980) );
  XNOR U11811 ( .A(n10982), .B(n10983), .Z(n10937) );
  XOR U11812 ( .A(n10938), .B(n10937), .Z(n10939) );
  XOR U11813 ( .A(n10940), .B(n10939), .Z(n10998) );
  XOR U11814 ( .A(n10999), .B(n10998), .Z(n11000) );
  NANDN U11815 ( .A(n10854), .B(n10853), .Z(n10858) );
  NANDN U11816 ( .A(n10856), .B(n10855), .Z(n10857) );
  AND U11817 ( .A(n10858), .B(n10857), .Z(n11013) );
  NAND U11818 ( .A(n10860), .B(n10859), .Z(n10864) );
  NANDN U11819 ( .A(n10862), .B(n10861), .Z(n10863) );
  AND U11820 ( .A(n10864), .B(n10863), .Z(n11011) );
  NANDN U11821 ( .A(n10866), .B(n10865), .Z(n10870) );
  OR U11822 ( .A(n10868), .B(n10867), .Z(n10869) );
  AND U11823 ( .A(n10870), .B(n10869), .Z(n11010) );
  XNOR U11824 ( .A(n11011), .B(n11010), .Z(n11012) );
  XNOR U11825 ( .A(n11013), .B(n11012), .Z(n11004) );
  XOR U11826 ( .A(n11005), .B(n11004), .Z(n11006) );
  NANDN U11827 ( .A(n10872), .B(n10871), .Z(n10876) );
  NANDN U11828 ( .A(n10874), .B(n10873), .Z(n10875) );
  NAND U11829 ( .A(n10876), .B(n10875), .Z(n11007) );
  XOR U11830 ( .A(n11006), .B(n11007), .Z(n11021) );
  NAND U11831 ( .A(n10878), .B(n10877), .Z(n10882) );
  NANDN U11832 ( .A(n10880), .B(n10879), .Z(n10881) );
  AND U11833 ( .A(n10882), .B(n10881), .Z(n11020) );
  NANDN U11834 ( .A(n10884), .B(n10883), .Z(n10888) );
  NAND U11835 ( .A(n10886), .B(n10885), .Z(n10887) );
  AND U11836 ( .A(n10888), .B(n10887), .Z(n11019) );
  XOR U11837 ( .A(n11020), .B(n11019), .Z(n11022) );
  XOR U11838 ( .A(n11021), .B(n11022), .Z(n11018) );
  NAND U11839 ( .A(n10890), .B(n10889), .Z(n10894) );
  NAND U11840 ( .A(n10892), .B(n10891), .Z(n10893) );
  NAND U11841 ( .A(n10894), .B(n10893), .Z(n11017) );
  NANDN U11842 ( .A(n10895), .B(n10896), .Z(n10901) );
  NOR U11843 ( .A(n10897), .B(n10896), .Z(n10899) );
  OR U11844 ( .A(n10899), .B(n10898), .Z(n10900) );
  AND U11845 ( .A(n10901), .B(n10900), .Z(n11016) );
  XOR U11846 ( .A(n11017), .B(n11016), .Z(n10902) );
  XNOR U11847 ( .A(n11018), .B(n10902), .Z(N245) );
  NANDN U11848 ( .A(n10904), .B(n10903), .Z(n10908) );
  NAND U11849 ( .A(n10906), .B(n10905), .Z(n10907) );
  AND U11850 ( .A(n10908), .B(n10907), .Z(n11035) );
  AND U11851 ( .A(x[242]), .B(y[1896]), .Z(n11806) );
  NAND U11852 ( .A(n11806), .B(n10909), .Z(n10913) );
  NAND U11853 ( .A(n10911), .B(n10910), .Z(n10912) );
  NAND U11854 ( .A(n10913), .B(n10912), .Z(n11106) );
  AND U11855 ( .A(x[235]), .B(y[1907]), .Z(n12525) );
  AND U11856 ( .A(x[225]), .B(y[1897]), .Z(n10914) );
  NAND U11857 ( .A(n12525), .B(n10914), .Z(n10918) );
  NAND U11858 ( .A(n10916), .B(n10915), .Z(n10917) );
  NAND U11859 ( .A(n10918), .B(n10917), .Z(n11105) );
  XOR U11860 ( .A(n11106), .B(n11105), .Z(n11108) );
  AND U11861 ( .A(x[239]), .B(y[1899]), .Z(n11794) );
  NAND U11862 ( .A(n11794), .B(n10919), .Z(n10923) );
  NAND U11863 ( .A(n10921), .B(n10920), .Z(n10922) );
  NAND U11864 ( .A(n10923), .B(n10922), .Z(n11070) );
  AND U11865 ( .A(o[116]), .B(n10924), .Z(n11092) );
  AND U11866 ( .A(x[224]), .B(y[1909]), .Z(n11089) );
  AND U11867 ( .A(x[245]), .B(y[1888]), .Z(n11090) );
  XOR U11868 ( .A(n11089), .B(n11090), .Z(n11091) );
  XOR U11869 ( .A(n11092), .B(n11091), .Z(n11068) );
  AND U11870 ( .A(x[229]), .B(y[1904]), .Z(n11076) );
  AND U11871 ( .A(x[240]), .B(y[1893]), .Z(n11075) );
  XOR U11872 ( .A(n11076), .B(n11075), .Z(n11074) );
  AND U11873 ( .A(x[239]), .B(y[1894]), .Z(n11073) );
  XOR U11874 ( .A(n11074), .B(n11073), .Z(n11067) );
  XOR U11875 ( .A(n11068), .B(n11067), .Z(n11069) );
  XOR U11876 ( .A(n11070), .B(n11069), .Z(n11107) );
  XOR U11877 ( .A(n11108), .B(n11107), .Z(n11124) );
  NANDN U11878 ( .A(n10926), .B(n10925), .Z(n10930) );
  NANDN U11879 ( .A(n10928), .B(n10927), .Z(n10929) );
  NAND U11880 ( .A(n10930), .B(n10929), .Z(n11123) );
  NANDN U11881 ( .A(n10932), .B(n10931), .Z(n10936) );
  NANDN U11882 ( .A(n10934), .B(n10933), .Z(n10935) );
  AND U11883 ( .A(n10936), .B(n10935), .Z(n11125) );
  XOR U11884 ( .A(n11126), .B(n11125), .Z(n11033) );
  NAND U11885 ( .A(n10938), .B(n10937), .Z(n10942) );
  NAND U11886 ( .A(n10940), .B(n10939), .Z(n10941) );
  AND U11887 ( .A(n10942), .B(n10941), .Z(n11032) );
  NANDN U11888 ( .A(n10944), .B(n10943), .Z(n10948) );
  NAND U11889 ( .A(n10946), .B(n10945), .Z(n10947) );
  AND U11890 ( .A(n10948), .B(n10947), .Z(n11132) );
  NAND U11891 ( .A(n11799), .B(n10949), .Z(n10953) );
  NAND U11892 ( .A(n10951), .B(n10950), .Z(n10952) );
  NAND U11893 ( .A(n10953), .B(n10952), .Z(n11039) );
  NAND U11894 ( .A(n12365), .B(n10954), .Z(n10958) );
  NAND U11895 ( .A(n10956), .B(n10955), .Z(n10957) );
  NAND U11896 ( .A(n10958), .B(n10957), .Z(n11120) );
  AND U11897 ( .A(y[1890]), .B(x[243]), .Z(n10960) );
  NAND U11898 ( .A(y[1898]), .B(x[235]), .Z(n10959) );
  XNOR U11899 ( .A(n10960), .B(n10959), .Z(n11057) );
  NAND U11900 ( .A(x[244]), .B(y[1889]), .Z(n11088) );
  XNOR U11901 ( .A(o[117]), .B(n11088), .Z(n11058) );
  XOR U11902 ( .A(n11057), .B(n11058), .Z(n11118) );
  AND U11903 ( .A(y[1891]), .B(x[242]), .Z(n10962) );
  NAND U11904 ( .A(y[1899]), .B(x[234]), .Z(n10961) );
  XNOR U11905 ( .A(n10962), .B(n10961), .Z(n11096) );
  AND U11906 ( .A(x[225]), .B(y[1908]), .Z(n11097) );
  XOR U11907 ( .A(n11096), .B(n11097), .Z(n11117) );
  XOR U11908 ( .A(n11118), .B(n11117), .Z(n11119) );
  XOR U11909 ( .A(n11120), .B(n11119), .Z(n11038) );
  XOR U11910 ( .A(n11039), .B(n11038), .Z(n11041) );
  AND U11911 ( .A(x[231]), .B(y[1902]), .Z(n11302) );
  AND U11912 ( .A(y[1903]), .B(x[230]), .Z(n10964) );
  NAND U11913 ( .A(y[1895]), .B(x[238]), .Z(n10963) );
  XNOR U11914 ( .A(n10964), .B(n10963), .Z(n11100) );
  XNOR U11915 ( .A(n11302), .B(n11100), .Z(n11047) );
  NAND U11916 ( .A(x[233]), .B(y[1900]), .Z(n11045) );
  NAND U11917 ( .A(x[232]), .B(y[1901]), .Z(n11044) );
  XOR U11918 ( .A(n11045), .B(n11044), .Z(n11046) );
  XNOR U11919 ( .A(n11047), .B(n11046), .Z(n11063) );
  AND U11920 ( .A(y[1897]), .B(x[236]), .Z(n10966) );
  NAND U11921 ( .A(y[1892]), .B(x[241]), .Z(n10965) );
  XNOR U11922 ( .A(n10966), .B(n10965), .Z(n11050) );
  AND U11923 ( .A(x[226]), .B(y[1907]), .Z(n11051) );
  XOR U11924 ( .A(n11050), .B(n11051), .Z(n11062) );
  AND U11925 ( .A(y[1896]), .B(x[237]), .Z(n10968) );
  NAND U11926 ( .A(y[1906]), .B(x[227]), .Z(n10967) );
  XNOR U11927 ( .A(n10968), .B(n10967), .Z(n11084) );
  AND U11928 ( .A(x[228]), .B(y[1905]), .Z(n11085) );
  XOR U11929 ( .A(n11084), .B(n11085), .Z(n11061) );
  XOR U11930 ( .A(n11062), .B(n11061), .Z(n11064) );
  XOR U11931 ( .A(n11063), .B(n11064), .Z(n11114) );
  NAND U11932 ( .A(n10970), .B(n10969), .Z(n10974) );
  NAND U11933 ( .A(n10972), .B(n10971), .Z(n10973) );
  NAND U11934 ( .A(n10974), .B(n10973), .Z(n11112) );
  NAND U11935 ( .A(n11076), .B(n10975), .Z(n10979) );
  NAND U11936 ( .A(n10977), .B(n10976), .Z(n10978) );
  NAND U11937 ( .A(n10979), .B(n10978), .Z(n11111) );
  XOR U11938 ( .A(n11112), .B(n11111), .Z(n11113) );
  XOR U11939 ( .A(n11114), .B(n11113), .Z(n11040) );
  XOR U11940 ( .A(n11041), .B(n11040), .Z(n11130) );
  NANDN U11941 ( .A(n10981), .B(n10980), .Z(n10985) );
  NAND U11942 ( .A(n10983), .B(n10982), .Z(n10984) );
  NAND U11943 ( .A(n10985), .B(n10984), .Z(n11137) );
  NAND U11944 ( .A(n10987), .B(n10986), .Z(n10991) );
  NANDN U11945 ( .A(n10989), .B(n10988), .Z(n10990) );
  NAND U11946 ( .A(n10991), .B(n10990), .Z(n11136) );
  NAND U11947 ( .A(n10993), .B(n10992), .Z(n10997) );
  NANDN U11948 ( .A(n10995), .B(n10994), .Z(n10996) );
  NAND U11949 ( .A(n10997), .B(n10996), .Z(n11135) );
  XOR U11950 ( .A(n11136), .B(n11135), .Z(n11138) );
  XOR U11951 ( .A(n11137), .B(n11138), .Z(n11129) );
  XOR U11952 ( .A(n11130), .B(n11129), .Z(n11131) );
  NAND U11953 ( .A(n10999), .B(n10998), .Z(n11003) );
  NANDN U11954 ( .A(n11001), .B(n11000), .Z(n11002) );
  NAND U11955 ( .A(n11003), .B(n11002), .Z(n11026) );
  XOR U11956 ( .A(n11027), .B(n11026), .Z(n11029) );
  XNOR U11957 ( .A(n11028), .B(n11029), .Z(n11150) );
  NAND U11958 ( .A(n11005), .B(n11004), .Z(n11009) );
  NANDN U11959 ( .A(n11007), .B(n11006), .Z(n11008) );
  AND U11960 ( .A(n11009), .B(n11008), .Z(n11149) );
  NANDN U11961 ( .A(n11011), .B(n11010), .Z(n11015) );
  NAND U11962 ( .A(n11013), .B(n11012), .Z(n11014) );
  AND U11963 ( .A(n11015), .B(n11014), .Z(n11148) );
  XOR U11964 ( .A(n11149), .B(n11148), .Z(n11151) );
  XOR U11965 ( .A(n11150), .B(n11151), .Z(n11144) );
  NAND U11966 ( .A(n11020), .B(n11019), .Z(n11024) );
  NAND U11967 ( .A(n11022), .B(n11021), .Z(n11023) );
  AND U11968 ( .A(n11024), .B(n11023), .Z(n11142) );
  IV U11969 ( .A(n11142), .Z(n11141) );
  XOR U11970 ( .A(n11143), .B(n11141), .Z(n11025) );
  XNOR U11971 ( .A(n11144), .B(n11025), .Z(N246) );
  NAND U11972 ( .A(n11027), .B(n11026), .Z(n11031) );
  NAND U11973 ( .A(n11029), .B(n11028), .Z(n11030) );
  AND U11974 ( .A(n11031), .B(n11030), .Z(n11158) );
  NANDN U11975 ( .A(n11033), .B(n11032), .Z(n11037) );
  NANDN U11976 ( .A(n11035), .B(n11034), .Z(n11036) );
  AND U11977 ( .A(n11037), .B(n11036), .Z(n11156) );
  NAND U11978 ( .A(n11039), .B(n11038), .Z(n11043) );
  NAND U11979 ( .A(n11041), .B(n11040), .Z(n11042) );
  NAND U11980 ( .A(n11043), .B(n11042), .Z(n11279) );
  NAND U11981 ( .A(n11045), .B(n11044), .Z(n11049) );
  NAND U11982 ( .A(n11047), .B(n11046), .Z(n11048) );
  NAND U11983 ( .A(n11049), .B(n11048), .Z(n11273) );
  NAND U11984 ( .A(n11807), .B(n11224), .Z(n11053) );
  NAND U11985 ( .A(n11051), .B(n11050), .Z(n11052) );
  NAND U11986 ( .A(n11053), .B(n11052), .Z(n11202) );
  AND U11987 ( .A(x[229]), .B(y[1905]), .Z(n11246) );
  AND U11988 ( .A(x[241]), .B(y[1893]), .Z(n11247) );
  XOR U11989 ( .A(n11246), .B(n11247), .Z(n11248) );
  AND U11990 ( .A(x[240]), .B(y[1894]), .Z(n11249) );
  XOR U11991 ( .A(n11248), .B(n11249), .Z(n11201) );
  AND U11992 ( .A(y[1892]), .B(x[242]), .Z(n11055) );
  NAND U11993 ( .A(y[1898]), .B(x[236]), .Z(n11054) );
  XNOR U11994 ( .A(n11055), .B(n11054), .Z(n11225) );
  AND U11995 ( .A(x[228]), .B(y[1906]), .Z(n11226) );
  XOR U11996 ( .A(n11225), .B(n11226), .Z(n11200) );
  XOR U11997 ( .A(n11201), .B(n11200), .Z(n11203) );
  XNOR U11998 ( .A(n11202), .B(n11203), .Z(n11270) );
  NAND U11999 ( .A(x[243]), .B(y[1898]), .Z(n12263) );
  NANDN U12000 ( .A(n12263), .B(n11056), .Z(n11060) );
  NAND U12001 ( .A(n11058), .B(n11057), .Z(n11059) );
  AND U12002 ( .A(n11060), .B(n11059), .Z(n11271) );
  XOR U12003 ( .A(n11270), .B(n11271), .Z(n11272) );
  XNOR U12004 ( .A(n11273), .B(n11272), .Z(n11276) );
  NAND U12005 ( .A(n11062), .B(n11061), .Z(n11066) );
  NAND U12006 ( .A(n11064), .B(n11063), .Z(n11065) );
  NAND U12007 ( .A(n11066), .B(n11065), .Z(n11259) );
  NAND U12008 ( .A(n11068), .B(n11067), .Z(n11072) );
  NAND U12009 ( .A(n11070), .B(n11069), .Z(n11071) );
  NAND U12010 ( .A(n11072), .B(n11071), .Z(n11258) );
  XOR U12011 ( .A(n11259), .B(n11258), .Z(n11261) );
  AND U12012 ( .A(n11074), .B(n11073), .Z(n11078) );
  NAND U12013 ( .A(n11076), .B(n11075), .Z(n11077) );
  NANDN U12014 ( .A(n11078), .B(n11077), .Z(n11221) );
  AND U12015 ( .A(y[1897]), .B(x[237]), .Z(n11080) );
  NAND U12016 ( .A(y[1890]), .B(x[244]), .Z(n11079) );
  XNOR U12017 ( .A(n11080), .B(n11079), .Z(n11242) );
  AND U12018 ( .A(x[226]), .B(y[1908]), .Z(n11243) );
  XOR U12019 ( .A(n11242), .B(n11243), .Z(n11219) );
  AND U12020 ( .A(y[1904]), .B(x[230]), .Z(n11082) );
  NAND U12021 ( .A(y[1895]), .B(x[239]), .Z(n11081) );
  XNOR U12022 ( .A(n11082), .B(n11081), .Z(n11254) );
  XOR U12023 ( .A(n11219), .B(n11218), .Z(n11220) );
  XOR U12024 ( .A(n11221), .B(n11220), .Z(n11265) );
  AND U12025 ( .A(x[237]), .B(y[1906]), .Z(n12526) );
  NAND U12026 ( .A(n11083), .B(n12526), .Z(n11087) );
  NAND U12027 ( .A(n11085), .B(n11084), .Z(n11086) );
  NAND U12028 ( .A(n11087), .B(n11086), .Z(n11191) );
  ANDN U12029 ( .B(o[117]), .A(n11088), .Z(n11213) );
  AND U12030 ( .A(x[225]), .B(y[1909]), .Z(n11214) );
  XOR U12031 ( .A(n11215), .B(n11214), .Z(n11212) );
  XOR U12032 ( .A(n11213), .B(n11212), .Z(n11188) );
  AND U12033 ( .A(x[238]), .B(y[1896]), .Z(n11206) );
  NAND U12034 ( .A(x[227]), .B(y[1907]), .Z(n11207) );
  XNOR U12035 ( .A(n11206), .B(n11207), .Z(n11208) );
  NAND U12036 ( .A(x[243]), .B(y[1891]), .Z(n11209) );
  XNOR U12037 ( .A(n11208), .B(n11209), .Z(n11189) );
  XOR U12038 ( .A(n11188), .B(n11189), .Z(n11190) );
  XOR U12039 ( .A(n11191), .B(n11190), .Z(n11264) );
  XOR U12040 ( .A(n11265), .B(n11264), .Z(n11267) );
  NAND U12041 ( .A(n11090), .B(n11089), .Z(n11094) );
  NAND U12042 ( .A(n11092), .B(n11091), .Z(n11093) );
  NAND U12043 ( .A(n11094), .B(n11093), .Z(n11183) );
  AND U12044 ( .A(x[242]), .B(y[1899]), .Z(n12265) );
  NAND U12045 ( .A(n12265), .B(n11095), .Z(n11099) );
  NAND U12046 ( .A(n11097), .B(n11096), .Z(n11098) );
  NAND U12047 ( .A(n11099), .B(n11098), .Z(n11182) );
  XOR U12048 ( .A(n11183), .B(n11182), .Z(n11185) );
  AND U12049 ( .A(x[238]), .B(y[1903]), .Z(n12275) );
  NAND U12050 ( .A(n12275), .B(n11253), .Z(n11102) );
  NAND U12051 ( .A(n11302), .B(n11100), .Z(n11101) );
  NAND U12052 ( .A(n11102), .B(n11101), .Z(n11197) );
  AND U12053 ( .A(x[224]), .B(y[1910]), .Z(n11229) );
  AND U12054 ( .A(x[246]), .B(y[1888]), .Z(n11230) );
  XOR U12055 ( .A(n11229), .B(n11230), .Z(n11231) );
  NAND U12056 ( .A(x[245]), .B(y[1889]), .Z(n11252) );
  XNOR U12057 ( .A(o[118]), .B(n11252), .Z(n11232) );
  XOR U12058 ( .A(n11231), .B(n11232), .Z(n11195) );
  AND U12059 ( .A(y[1903]), .B(x[231]), .Z(n11104) );
  NAND U12060 ( .A(y[1902]), .B(x[232]), .Z(n11103) );
  XNOR U12061 ( .A(n11104), .B(n11103), .Z(n11235) );
  XOR U12062 ( .A(n11195), .B(n11194), .Z(n11196) );
  XOR U12063 ( .A(n11197), .B(n11196), .Z(n11184) );
  XOR U12064 ( .A(n11185), .B(n11184), .Z(n11266) );
  XOR U12065 ( .A(n11267), .B(n11266), .Z(n11260) );
  XOR U12066 ( .A(n11261), .B(n11260), .Z(n11277) );
  XOR U12067 ( .A(n11276), .B(n11277), .Z(n11278) );
  XOR U12068 ( .A(n11279), .B(n11278), .Z(n11173) );
  NAND U12069 ( .A(n11106), .B(n11105), .Z(n11110) );
  NAND U12070 ( .A(n11108), .B(n11107), .Z(n11109) );
  NAND U12071 ( .A(n11110), .B(n11109), .Z(n11179) );
  NAND U12072 ( .A(n11112), .B(n11111), .Z(n11116) );
  NAND U12073 ( .A(n11114), .B(n11113), .Z(n11115) );
  NAND U12074 ( .A(n11116), .B(n11115), .Z(n11177) );
  NAND U12075 ( .A(n11118), .B(n11117), .Z(n11122) );
  NAND U12076 ( .A(n11120), .B(n11119), .Z(n11121) );
  NAND U12077 ( .A(n11122), .B(n11121), .Z(n11176) );
  XOR U12078 ( .A(n11177), .B(n11176), .Z(n11178) );
  XOR U12079 ( .A(n11179), .B(n11178), .Z(n11171) );
  NANDN U12080 ( .A(n11124), .B(n11123), .Z(n11128) );
  NAND U12081 ( .A(n11126), .B(n11125), .Z(n11127) );
  NAND U12082 ( .A(n11128), .B(n11127), .Z(n11170) );
  NAND U12083 ( .A(n11130), .B(n11129), .Z(n11134) );
  NANDN U12084 ( .A(n11132), .B(n11131), .Z(n11133) );
  NAND U12085 ( .A(n11134), .B(n11133), .Z(n11165) );
  NAND U12086 ( .A(n11136), .B(n11135), .Z(n11140) );
  NAND U12087 ( .A(n11138), .B(n11137), .Z(n11139) );
  NAND U12088 ( .A(n11140), .B(n11139), .Z(n11164) );
  XOR U12089 ( .A(n11165), .B(n11164), .Z(n11166) );
  XNOR U12090 ( .A(n11158), .B(n11157), .Z(n11161) );
  OR U12091 ( .A(n11143), .B(n11141), .Z(n11147) );
  ANDN U12092 ( .B(n11143), .A(n11142), .Z(n11145) );
  OR U12093 ( .A(n11145), .B(n11144), .Z(n11146) );
  AND U12094 ( .A(n11147), .B(n11146), .Z(n11162) );
  NANDN U12095 ( .A(n11149), .B(n11148), .Z(n11153) );
  NANDN U12096 ( .A(n11151), .B(n11150), .Z(n11152) );
  AND U12097 ( .A(n11153), .B(n11152), .Z(n11163) );
  XOR U12098 ( .A(n11162), .B(n11163), .Z(n11154) );
  XNOR U12099 ( .A(n11161), .B(n11154), .Z(N247) );
  NANDN U12100 ( .A(n11156), .B(n11155), .Z(n11160) );
  NAND U12101 ( .A(n11158), .B(n11157), .Z(n11159) );
  NAND U12102 ( .A(n11160), .B(n11159), .Z(n11414) );
  IV U12103 ( .A(n11414), .Z(n11413) );
  NAND U12104 ( .A(n11165), .B(n11164), .Z(n11169) );
  NANDN U12105 ( .A(n11167), .B(n11166), .Z(n11168) );
  AND U12106 ( .A(n11169), .B(n11168), .Z(n11422) );
  NANDN U12107 ( .A(n11171), .B(n11170), .Z(n11175) );
  NANDN U12108 ( .A(n11173), .B(n11172), .Z(n11174) );
  NAND U12109 ( .A(n11175), .B(n11174), .Z(n11420) );
  NAND U12110 ( .A(n11177), .B(n11176), .Z(n11181) );
  NAND U12111 ( .A(n11179), .B(n11178), .Z(n11180) );
  NAND U12112 ( .A(n11181), .B(n11180), .Z(n11398) );
  NAND U12113 ( .A(n11183), .B(n11182), .Z(n11187) );
  NAND U12114 ( .A(n11185), .B(n11184), .Z(n11186) );
  NAND U12115 ( .A(n11187), .B(n11186), .Z(n11392) );
  NAND U12116 ( .A(n11189), .B(n11188), .Z(n11193) );
  NAND U12117 ( .A(n11191), .B(n11190), .Z(n11192) );
  NAND U12118 ( .A(n11193), .B(n11192), .Z(n11390) );
  NAND U12119 ( .A(n11195), .B(n11194), .Z(n11199) );
  NAND U12120 ( .A(n11197), .B(n11196), .Z(n11198) );
  NAND U12121 ( .A(n11199), .B(n11198), .Z(n11389) );
  XOR U12122 ( .A(n11390), .B(n11389), .Z(n11391) );
  XOR U12123 ( .A(n11392), .B(n11391), .Z(n11410) );
  NAND U12124 ( .A(n11201), .B(n11200), .Z(n11205) );
  NAND U12125 ( .A(n11203), .B(n11202), .Z(n11204) );
  NAND U12126 ( .A(n11205), .B(n11204), .Z(n11408) );
  NANDN U12127 ( .A(n11207), .B(n11206), .Z(n11211) );
  NANDN U12128 ( .A(n11209), .B(n11208), .Z(n11210) );
  AND U12129 ( .A(n11211), .B(n11210), .Z(n11336) );
  XNOR U12130 ( .A(n11336), .B(n11335), .Z(n11337) );
  AND U12131 ( .A(y[1904]), .B(x[231]), .Z(n11217) );
  NAND U12132 ( .A(y[1902]), .B(x[233]), .Z(n11216) );
  XOR U12133 ( .A(n11217), .B(n11216), .Z(n11304) );
  XNOR U12134 ( .A(n11303), .B(n11304), .Z(n11341) );
  NAND U12135 ( .A(x[234]), .B(y[1901]), .Z(n11342) );
  XNOR U12136 ( .A(n11341), .B(n11342), .Z(n11343) );
  AND U12137 ( .A(x[230]), .B(y[1905]), .Z(n11294) );
  NAND U12138 ( .A(x[239]), .B(y[1896]), .Z(n11295) );
  XNOR U12139 ( .A(n11294), .B(n11295), .Z(n11296) );
  NAND U12140 ( .A(x[235]), .B(y[1900]), .Z(n11297) );
  XOR U12141 ( .A(n11296), .B(n11297), .Z(n11344) );
  XOR U12142 ( .A(n11343), .B(n11344), .Z(n11338) );
  XNOR U12143 ( .A(n11337), .B(n11338), .Z(n11407) );
  XOR U12144 ( .A(n11408), .B(n11407), .Z(n11409) );
  XOR U12145 ( .A(n11410), .B(n11409), .Z(n11396) );
  NAND U12146 ( .A(n11219), .B(n11218), .Z(n11223) );
  NAND U12147 ( .A(n11221), .B(n11220), .Z(n11222) );
  NAND U12148 ( .A(n11223), .B(n11222), .Z(n11330) );
  AND U12149 ( .A(x[242]), .B(y[1898]), .Z(n12107) );
  NAND U12150 ( .A(n12107), .B(n11224), .Z(n11228) );
  NAND U12151 ( .A(n11226), .B(n11225), .Z(n11227) );
  NAND U12152 ( .A(n11228), .B(n11227), .Z(n11366) );
  NAND U12153 ( .A(n11230), .B(n11229), .Z(n11234) );
  NAND U12154 ( .A(n11232), .B(n11231), .Z(n11233) );
  NAND U12155 ( .A(n11234), .B(n11233), .Z(n11365) );
  XOR U12156 ( .A(n11366), .B(n11365), .Z(n11368) );
  NAND U12157 ( .A(n11302), .B(n11303), .Z(n11238) );
  NANDN U12158 ( .A(n11236), .B(n11235), .Z(n11237) );
  NAND U12159 ( .A(n11238), .B(n11237), .Z(n11379) );
  AND U12160 ( .A(x[224]), .B(y[1911]), .Z(n11313) );
  NAND U12161 ( .A(x[247]), .B(y[1888]), .Z(n11314) );
  XNOR U12162 ( .A(n11313), .B(n11314), .Z(n11315) );
  NAND U12163 ( .A(x[246]), .B(y[1889]), .Z(n11293) );
  XOR U12164 ( .A(o[119]), .B(n11293), .Z(n11316) );
  XNOR U12165 ( .A(n11315), .B(n11316), .Z(n11378) );
  NAND U12166 ( .A(y[1891]), .B(x[244]), .Z(n11239) );
  XNOR U12167 ( .A(n11240), .B(n11239), .Z(n11290) );
  AND U12168 ( .A(x[243]), .B(y[1892]), .Z(n11289) );
  XOR U12169 ( .A(n11290), .B(n11289), .Z(n11377) );
  XOR U12170 ( .A(n11378), .B(n11377), .Z(n11380) );
  XOR U12171 ( .A(n11379), .B(n11380), .Z(n11367) );
  XOR U12172 ( .A(n11368), .B(n11367), .Z(n11329) );
  XOR U12173 ( .A(n11330), .B(n11329), .Z(n11332) );
  NAND U12174 ( .A(x[244]), .B(y[1897]), .Z(n12287) );
  AND U12175 ( .A(x[237]), .B(y[1890]), .Z(n11241) );
  NANDN U12176 ( .A(n12287), .B(n11241), .Z(n11245) );
  NAND U12177 ( .A(n11243), .B(n11242), .Z(n11244) );
  NAND U12178 ( .A(n11245), .B(n11244), .Z(n11324) );
  NAND U12179 ( .A(n11247), .B(n11246), .Z(n11251) );
  NAND U12180 ( .A(n11249), .B(n11248), .Z(n11250) );
  NAND U12181 ( .A(n11251), .B(n11250), .Z(n11386) );
  AND U12182 ( .A(x[237]), .B(y[1898]), .Z(n11359) );
  NAND U12183 ( .A(x[226]), .B(y[1909]), .Z(n11360) );
  XNOR U12184 ( .A(n11359), .B(n11360), .Z(n11361) );
  NAND U12185 ( .A(x[245]), .B(y[1890]), .Z(n11362) );
  XNOR U12186 ( .A(n11361), .B(n11362), .Z(n11383) );
  ANDN U12187 ( .B(o[118]), .A(n11252), .Z(n11309) );
  AND U12188 ( .A(x[236]), .B(y[1899]), .Z(n11307) );
  NAND U12189 ( .A(x[225]), .B(y[1910]), .Z(n11308) );
  XOR U12190 ( .A(n11307), .B(n11308), .Z(n11310) );
  XNOR U12191 ( .A(n11309), .B(n11310), .Z(n11384) );
  XOR U12192 ( .A(n11383), .B(n11384), .Z(n11385) );
  XOR U12193 ( .A(n11386), .B(n11385), .Z(n11323) );
  XOR U12194 ( .A(n11324), .B(n11323), .Z(n11326) );
  AND U12195 ( .A(x[239]), .B(y[1904]), .Z(n12480) );
  NAND U12196 ( .A(n11253), .B(n12480), .Z(n11257) );
  NANDN U12197 ( .A(n11255), .B(n11254), .Z(n11256) );
  NAND U12198 ( .A(n11257), .B(n11256), .Z(n11374) );
  AND U12199 ( .A(x[238]), .B(y[1897]), .Z(n11353) );
  NAND U12200 ( .A(x[227]), .B(y[1908]), .Z(n11354) );
  XNOR U12201 ( .A(n11353), .B(n11354), .Z(n11355) );
  NAND U12202 ( .A(x[228]), .B(y[1907]), .Z(n11356) );
  XNOR U12203 ( .A(n11355), .B(n11356), .Z(n11371) );
  AND U12204 ( .A(x[229]), .B(y[1906]), .Z(n11347) );
  NAND U12205 ( .A(x[242]), .B(y[1893]), .Z(n11348) );
  XNOR U12206 ( .A(n11347), .B(n11348), .Z(n11349) );
  NAND U12207 ( .A(x[241]), .B(y[1894]), .Z(n11350) );
  XNOR U12208 ( .A(n11349), .B(n11350), .Z(n11372) );
  XOR U12209 ( .A(n11371), .B(n11372), .Z(n11373) );
  XOR U12210 ( .A(n11374), .B(n11373), .Z(n11325) );
  XOR U12211 ( .A(n11326), .B(n11325), .Z(n11331) );
  XOR U12212 ( .A(n11332), .B(n11331), .Z(n11395) );
  XOR U12213 ( .A(n11396), .B(n11395), .Z(n11397) );
  XNOR U12214 ( .A(n11398), .B(n11397), .Z(n11285) );
  NAND U12215 ( .A(n11259), .B(n11258), .Z(n11263) );
  NAND U12216 ( .A(n11261), .B(n11260), .Z(n11262) );
  NAND U12217 ( .A(n11263), .B(n11262), .Z(n11404) );
  NAND U12218 ( .A(n11265), .B(n11264), .Z(n11269) );
  NAND U12219 ( .A(n11267), .B(n11266), .Z(n11268) );
  NAND U12220 ( .A(n11269), .B(n11268), .Z(n11402) );
  NAND U12221 ( .A(n11271), .B(n11270), .Z(n11275) );
  NAND U12222 ( .A(n11273), .B(n11272), .Z(n11274) );
  AND U12223 ( .A(n11275), .B(n11274), .Z(n11401) );
  XOR U12224 ( .A(n11402), .B(n11401), .Z(n11403) );
  XNOR U12225 ( .A(n11404), .B(n11403), .Z(n11283) );
  NAND U12226 ( .A(n11277), .B(n11276), .Z(n11281) );
  NAND U12227 ( .A(n11279), .B(n11278), .Z(n11280) );
  AND U12228 ( .A(n11281), .B(n11280), .Z(n11284) );
  XOR U12229 ( .A(n11283), .B(n11284), .Z(n11286) );
  XNOR U12230 ( .A(n11285), .B(n11286), .Z(n11421) );
  XNOR U12231 ( .A(n11422), .B(n11423), .Z(n11416) );
  XNOR U12232 ( .A(n11415), .B(n11416), .Z(n11282) );
  XOR U12233 ( .A(n11413), .B(n11282), .Z(N248) );
  NAND U12234 ( .A(n11284), .B(n11283), .Z(n11288) );
  NAND U12235 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U12236 ( .A(n11288), .B(n11287), .Z(n11563) );
  AND U12237 ( .A(x[244]), .B(y[1895]), .Z(n11767) );
  NAND U12238 ( .A(n11767), .B(n11455), .Z(n11292) );
  NAND U12239 ( .A(n11290), .B(n11289), .Z(n11291) );
  AND U12240 ( .A(n11292), .B(n11291), .Z(n11475) );
  AND U12241 ( .A(x[246]), .B(y[1890]), .Z(n11494) );
  XOR U12242 ( .A(n11495), .B(n11494), .Z(n11492) );
  AND U12243 ( .A(x[226]), .B(y[1910]), .Z(n11493) );
  XOR U12244 ( .A(n11492), .B(n11493), .Z(n11473) );
  ANDN U12245 ( .B(o[119]), .A(n11293), .Z(n11499) );
  AND U12246 ( .A(x[225]), .B(y[1911]), .Z(n11500) );
  XOR U12247 ( .A(n11501), .B(n11500), .Z(n11498) );
  XOR U12248 ( .A(n11499), .B(n11498), .Z(n11472) );
  XOR U12249 ( .A(n11473), .B(n11472), .Z(n11474) );
  XNOR U12250 ( .A(n11475), .B(n11474), .Z(n11529) );
  NANDN U12251 ( .A(n11295), .B(n11294), .Z(n11299) );
  NANDN U12252 ( .A(n11297), .B(n11296), .Z(n11298) );
  AND U12253 ( .A(n11299), .B(n11298), .Z(n11469) );
  AND U12254 ( .A(y[1896]), .B(x[240]), .Z(n11301) );
  NAND U12255 ( .A(y[1891]), .B(x[245]), .Z(n11300) );
  XNOR U12256 ( .A(n11301), .B(n11300), .Z(n11456) );
  NAND U12257 ( .A(x[229]), .B(y[1907]), .Z(n11457) );
  XNOR U12258 ( .A(n11456), .B(n11457), .Z(n11466) );
  AND U12259 ( .A(x[230]), .B(y[1906]), .Z(n11755) );
  NAND U12260 ( .A(x[244]), .B(y[1892]), .Z(n11676) );
  XNOR U12261 ( .A(n11755), .B(n11676), .Z(n11462) );
  NAND U12262 ( .A(x[243]), .B(y[1893]), .Z(n11463) );
  XOR U12263 ( .A(n11462), .B(n11463), .Z(n11467) );
  XNOR U12264 ( .A(n11466), .B(n11467), .Z(n11468) );
  XNOR U12265 ( .A(n11469), .B(n11468), .Z(n11447) );
  NANDN U12266 ( .A(n11603), .B(n11302), .Z(n11306) );
  NANDN U12267 ( .A(n11304), .B(n11303), .Z(n11305) );
  AND U12268 ( .A(n11306), .B(n11305), .Z(n11446) );
  NANDN U12269 ( .A(n11308), .B(n11307), .Z(n11312) );
  NANDN U12270 ( .A(n11310), .B(n11309), .Z(n11311) );
  NAND U12271 ( .A(n11312), .B(n11311), .Z(n11445) );
  XOR U12272 ( .A(n11446), .B(n11445), .Z(n11448) );
  XOR U12273 ( .A(n11447), .B(n11448), .Z(n11530) );
  XNOR U12274 ( .A(n11529), .B(n11530), .Z(n11532) );
  NANDN U12275 ( .A(n11314), .B(n11313), .Z(n11318) );
  NANDN U12276 ( .A(n11316), .B(n11315), .Z(n11317) );
  AND U12277 ( .A(n11318), .B(n11317), .Z(n11512) );
  AND U12278 ( .A(x[227]), .B(y[1909]), .Z(n11517) );
  XOR U12279 ( .A(n11518), .B(n11517), .Z(n11520) );
  NAND U12280 ( .A(x[228]), .B(y[1908]), .Z(n11519) );
  XNOR U12281 ( .A(n11520), .B(n11519), .Z(n11511) );
  XNOR U12282 ( .A(n11512), .B(n11511), .Z(n11513) );
  AND U12283 ( .A(y[1903]), .B(x[233]), .Z(n11320) );
  NAND U12284 ( .A(y[1902]), .B(x[234]), .Z(n11319) );
  XNOR U12285 ( .A(n11320), .B(n11319), .Z(n11483) );
  AND U12286 ( .A(y[1898]), .B(x[238]), .Z(n11322) );
  NAND U12287 ( .A(y[1904]), .B(x[232]), .Z(n11321) );
  XNOR U12288 ( .A(n11322), .B(n11321), .Z(n11488) );
  NAND U12289 ( .A(x[235]), .B(y[1901]), .Z(n11489) );
  XOR U12290 ( .A(n11488), .B(n11489), .Z(n11484) );
  XOR U12291 ( .A(n11483), .B(n11484), .Z(n11514) );
  XNOR U12292 ( .A(n11513), .B(n11514), .Z(n11531) );
  XNOR U12293 ( .A(n11532), .B(n11531), .Z(n11542) );
  NAND U12294 ( .A(n11324), .B(n11323), .Z(n11328) );
  NAND U12295 ( .A(n11326), .B(n11325), .Z(n11327) );
  AND U12296 ( .A(n11328), .B(n11327), .Z(n11541) );
  XOR U12297 ( .A(n11542), .B(n11541), .Z(n11543) );
  NAND U12298 ( .A(n11330), .B(n11329), .Z(n11334) );
  NAND U12299 ( .A(n11332), .B(n11331), .Z(n11333) );
  AND U12300 ( .A(n11334), .B(n11333), .Z(n11544) );
  XOR U12301 ( .A(n11543), .B(n11544), .Z(n11550) );
  NANDN U12302 ( .A(n11336), .B(n11335), .Z(n11340) );
  NANDN U12303 ( .A(n11338), .B(n11337), .Z(n11339) );
  AND U12304 ( .A(n11340), .B(n11339), .Z(n11537) );
  NANDN U12305 ( .A(n11342), .B(n11341), .Z(n11346) );
  NANDN U12306 ( .A(n11344), .B(n11343), .Z(n11345) );
  AND U12307 ( .A(n11346), .B(n11345), .Z(n11536) );
  NANDN U12308 ( .A(n11348), .B(n11347), .Z(n11352) );
  NANDN U12309 ( .A(n11350), .B(n11349), .Z(n11351) );
  AND U12310 ( .A(n11352), .B(n11351), .Z(n11454) );
  AND U12311 ( .A(x[224]), .B(y[1912]), .Z(n11523) );
  NAND U12312 ( .A(x[248]), .B(y[1888]), .Z(n11524) );
  XNOR U12313 ( .A(n11523), .B(n11524), .Z(n11525) );
  AND U12314 ( .A(x[247]), .B(y[1889]), .Z(n11510) );
  XNOR U12315 ( .A(n11510), .B(o[120]), .Z(n11526) );
  XNOR U12316 ( .A(n11525), .B(n11526), .Z(n11452) );
  AND U12317 ( .A(x[231]), .B(y[1905]), .Z(n11504) );
  NAND U12318 ( .A(x[242]), .B(y[1894]), .Z(n11505) );
  NAND U12319 ( .A(x[241]), .B(y[1895]), .Z(n11507) );
  XOR U12320 ( .A(n11452), .B(n11451), .Z(n11453) );
  XNOR U12321 ( .A(n11454), .B(n11453), .Z(n11441) );
  NANDN U12322 ( .A(n11354), .B(n11353), .Z(n11358) );
  NANDN U12323 ( .A(n11356), .B(n11355), .Z(n11357) );
  AND U12324 ( .A(n11358), .B(n11357), .Z(n11440) );
  NANDN U12325 ( .A(n11360), .B(n11359), .Z(n11364) );
  NANDN U12326 ( .A(n11362), .B(n11361), .Z(n11363) );
  NAND U12327 ( .A(n11364), .B(n11363), .Z(n11439) );
  XOR U12328 ( .A(n11440), .B(n11439), .Z(n11442) );
  XNOR U12329 ( .A(n11441), .B(n11442), .Z(n11535) );
  XOR U12330 ( .A(n11536), .B(n11535), .Z(n11538) );
  XNOR U12331 ( .A(n11537), .B(n11538), .Z(n11436) );
  NAND U12332 ( .A(n11366), .B(n11365), .Z(n11370) );
  NAND U12333 ( .A(n11368), .B(n11367), .Z(n11369) );
  AND U12334 ( .A(n11370), .B(n11369), .Z(n11479) );
  NAND U12335 ( .A(n11372), .B(n11371), .Z(n11376) );
  NAND U12336 ( .A(n11374), .B(n11373), .Z(n11375) );
  AND U12337 ( .A(n11376), .B(n11375), .Z(n11477) );
  NAND U12338 ( .A(n11378), .B(n11377), .Z(n11382) );
  NAND U12339 ( .A(n11380), .B(n11379), .Z(n11381) );
  AND U12340 ( .A(n11382), .B(n11381), .Z(n11476) );
  XOR U12341 ( .A(n11477), .B(n11476), .Z(n11478) );
  XOR U12342 ( .A(n11479), .B(n11478), .Z(n11433) );
  NAND U12343 ( .A(n11384), .B(n11383), .Z(n11388) );
  NAND U12344 ( .A(n11386), .B(n11385), .Z(n11387) );
  AND U12345 ( .A(n11388), .B(n11387), .Z(n11434) );
  XOR U12346 ( .A(n11433), .B(n11434), .Z(n11435) );
  XOR U12347 ( .A(n11436), .B(n11435), .Z(n11547) );
  NAND U12348 ( .A(n11390), .B(n11389), .Z(n11394) );
  NAND U12349 ( .A(n11392), .B(n11391), .Z(n11393) );
  AND U12350 ( .A(n11394), .B(n11393), .Z(n11548) );
  XOR U12351 ( .A(n11547), .B(n11548), .Z(n11549) );
  XNOR U12352 ( .A(n11550), .B(n11549), .Z(n11561) );
  NAND U12353 ( .A(n11396), .B(n11395), .Z(n11400) );
  NAND U12354 ( .A(n11398), .B(n11397), .Z(n11399) );
  NAND U12355 ( .A(n11400), .B(n11399), .Z(n11430) );
  NAND U12356 ( .A(n11402), .B(n11401), .Z(n11406) );
  NAND U12357 ( .A(n11404), .B(n11403), .Z(n11405) );
  NAND U12358 ( .A(n11406), .B(n11405), .Z(n11428) );
  NAND U12359 ( .A(n11408), .B(n11407), .Z(n11412) );
  NAND U12360 ( .A(n11410), .B(n11409), .Z(n11411) );
  NAND U12361 ( .A(n11412), .B(n11411), .Z(n11427) );
  XOR U12362 ( .A(n11428), .B(n11427), .Z(n11429) );
  XOR U12363 ( .A(n11430), .B(n11429), .Z(n11560) );
  XOR U12364 ( .A(n11561), .B(n11560), .Z(n11562) );
  XNOR U12365 ( .A(n11563), .B(n11562), .Z(n11556) );
  OR U12366 ( .A(n11415), .B(n11413), .Z(n11419) );
  ANDN U12367 ( .B(n11415), .A(n11414), .Z(n11417) );
  OR U12368 ( .A(n11417), .B(n11416), .Z(n11418) );
  AND U12369 ( .A(n11419), .B(n11418), .Z(n11555) );
  NANDN U12370 ( .A(n11421), .B(n11420), .Z(n11425) );
  NANDN U12371 ( .A(n11423), .B(n11422), .Z(n11424) );
  AND U12372 ( .A(n11425), .B(n11424), .Z(n11554) );
  IV U12373 ( .A(n11554), .Z(n11553) );
  XOR U12374 ( .A(n11555), .B(n11553), .Z(n11426) );
  XNOR U12375 ( .A(n11556), .B(n11426), .Z(N249) );
  NAND U12376 ( .A(n11428), .B(n11427), .Z(n11432) );
  NAND U12377 ( .A(n11430), .B(n11429), .Z(n11431) );
  AND U12378 ( .A(n11432), .B(n11431), .Z(n11715) );
  NAND U12379 ( .A(n11434), .B(n11433), .Z(n11438) );
  NAND U12380 ( .A(n11436), .B(n11435), .Z(n11437) );
  NAND U12381 ( .A(n11438), .B(n11437), .Z(n11575) );
  NANDN U12382 ( .A(n11440), .B(n11439), .Z(n11444) );
  NANDN U12383 ( .A(n11442), .B(n11441), .Z(n11443) );
  AND U12384 ( .A(n11444), .B(n11443), .Z(n11592) );
  NANDN U12385 ( .A(n11446), .B(n11445), .Z(n11450) );
  NANDN U12386 ( .A(n11448), .B(n11447), .Z(n11449) );
  NAND U12387 ( .A(n11450), .B(n11449), .Z(n11591) );
  XNOR U12388 ( .A(n11592), .B(n11591), .Z(n11593) );
  NAND U12389 ( .A(x[245]), .B(y[1896]), .Z(n12452) );
  NANDN U12390 ( .A(n12452), .B(n11455), .Z(n11459) );
  NANDN U12391 ( .A(n11457), .B(n11456), .Z(n11458) );
  NAND U12392 ( .A(n11459), .B(n11458), .Z(n11695) );
  AND U12393 ( .A(x[246]), .B(y[1891]), .Z(n11666) );
  AND U12394 ( .A(x[229]), .B(y[1908]), .Z(n11664) );
  NAND U12395 ( .A(x[241]), .B(y[1896]), .Z(n11663) );
  XNOR U12396 ( .A(n11664), .B(n11663), .Z(n11665) );
  XNOR U12397 ( .A(n11666), .B(n11665), .Z(n11694) );
  AND U12398 ( .A(y[1893]), .B(x[244]), .Z(n11461) );
  NAND U12399 ( .A(y[1892]), .B(x[245]), .Z(n11460) );
  XNOR U12400 ( .A(n11461), .B(n11460), .Z(n11678) );
  AND U12401 ( .A(x[243]), .B(y[1894]), .Z(n11677) );
  XOR U12402 ( .A(n11678), .B(n11677), .Z(n11693) );
  XOR U12403 ( .A(n11694), .B(n11693), .Z(n11696) );
  XOR U12404 ( .A(n11695), .B(n11696), .Z(n11620) );
  NANDN U12405 ( .A(n11676), .B(n11755), .Z(n11465) );
  NANDN U12406 ( .A(n11463), .B(n11462), .Z(n11464) );
  NAND U12407 ( .A(n11465), .B(n11464), .Z(n11701) );
  AND U12408 ( .A(x[239]), .B(y[1898]), .Z(n11684) );
  AND U12409 ( .A(x[242]), .B(y[1895]), .Z(n11682) );
  NAND U12410 ( .A(x[230]), .B(y[1907]), .Z(n11681) );
  XNOR U12411 ( .A(n11682), .B(n11681), .Z(n11683) );
  XNOR U12412 ( .A(n11684), .B(n11683), .Z(n11700) );
  AND U12413 ( .A(x[247]), .B(y[1890]), .Z(n11660) );
  AND U12414 ( .A(x[228]), .B(y[1909]), .Z(n11658) );
  NAND U12415 ( .A(x[240]), .B(y[1897]), .Z(n11657) );
  XNOR U12416 ( .A(n11658), .B(n11657), .Z(n11659) );
  XNOR U12417 ( .A(n11660), .B(n11659), .Z(n11699) );
  XNOR U12418 ( .A(n11700), .B(n11699), .Z(n11702) );
  XOR U12419 ( .A(n11701), .B(n11702), .Z(n11619) );
  XOR U12420 ( .A(n11620), .B(n11619), .Z(n11621) );
  XOR U12421 ( .A(n11622), .B(n11621), .Z(n11634) );
  NANDN U12422 ( .A(n11467), .B(n11466), .Z(n11471) );
  NANDN U12423 ( .A(n11469), .B(n11468), .Z(n11470) );
  AND U12424 ( .A(n11471), .B(n11470), .Z(n11632) );
  XNOR U12425 ( .A(n11632), .B(n11631), .Z(n11633) );
  XOR U12426 ( .A(n11634), .B(n11633), .Z(n11594) );
  XOR U12427 ( .A(n11593), .B(n11594), .Z(n11574) );
  NAND U12428 ( .A(n11477), .B(n11476), .Z(n11481) );
  NAND U12429 ( .A(n11479), .B(n11478), .Z(n11480) );
  NAND U12430 ( .A(n11481), .B(n11480), .Z(n11573) );
  XOR U12431 ( .A(n11574), .B(n11573), .Z(n11576) );
  XNOR U12432 ( .A(n11575), .B(n11576), .Z(n11569) );
  NANDN U12433 ( .A(n11604), .B(n11482), .Z(n11486) );
  NANDN U12434 ( .A(n11484), .B(n11483), .Z(n11485) );
  AND U12435 ( .A(n11486), .B(n11485), .Z(n11626) );
  AND U12436 ( .A(x[238]), .B(y[1904]), .Z(n12415) );
  NAND U12437 ( .A(n12415), .B(n11487), .Z(n11491) );
  NANDN U12438 ( .A(n11489), .B(n11488), .Z(n11490) );
  AND U12439 ( .A(n11491), .B(n11490), .Z(n11654) );
  AND U12440 ( .A(x[235]), .B(y[1902]), .Z(n11673) );
  AND U12441 ( .A(x[236]), .B(y[1901]), .Z(n11671) );
  NAND U12442 ( .A(x[231]), .B(y[1906]), .Z(n11670) );
  XNOR U12443 ( .A(n11671), .B(n11670), .Z(n11672) );
  XNOR U12444 ( .A(n11673), .B(n11672), .Z(n11652) );
  NAND U12445 ( .A(x[248]), .B(y[1889]), .Z(n11669) );
  XNOR U12446 ( .A(o[121]), .B(n11669), .Z(n11639) );
  NAND U12447 ( .A(x[225]), .B(y[1912]), .Z(n11640) );
  XNOR U12448 ( .A(n11639), .B(n11640), .Z(n11641) );
  NAND U12449 ( .A(x[237]), .B(y[1900]), .Z(n11642) );
  XNOR U12450 ( .A(n11641), .B(n11642), .Z(n11651) );
  XNOR U12451 ( .A(n11652), .B(n11651), .Z(n11653) );
  XNOR U12452 ( .A(n11654), .B(n11653), .Z(n11625) );
  XNOR U12453 ( .A(n11626), .B(n11625), .Z(n11628) );
  NAND U12454 ( .A(n11493), .B(n11492), .Z(n11497) );
  AND U12455 ( .A(n11495), .B(n11494), .Z(n11496) );
  ANDN U12456 ( .B(n11497), .A(n11496), .Z(n11614) );
  AND U12457 ( .A(n11499), .B(n11498), .Z(n11503) );
  NAND U12458 ( .A(n11501), .B(n11500), .Z(n11502) );
  NANDN U12459 ( .A(n11503), .B(n11502), .Z(n11613) );
  XNOR U12460 ( .A(n11614), .B(n11613), .Z(n11615) );
  NANDN U12461 ( .A(n11505), .B(n11504), .Z(n11509) );
  NANDN U12462 ( .A(n11507), .B(n11506), .Z(n11508) );
  NAND U12463 ( .A(n11509), .B(n11508), .Z(n11609) );
  AND U12464 ( .A(x[232]), .B(y[1905]), .Z(n11606) );
  XOR U12465 ( .A(n11603), .B(n11604), .Z(n11605) );
  XNOR U12466 ( .A(n11606), .B(n11605), .Z(n11608) );
  AND U12467 ( .A(n11510), .B(o[120]), .Z(n11600) );
  AND U12468 ( .A(x[249]), .B(y[1888]), .Z(n11598) );
  NAND U12469 ( .A(x[224]), .B(y[1913]), .Z(n11597) );
  XNOR U12470 ( .A(n11598), .B(n11597), .Z(n11599) );
  XNOR U12471 ( .A(n11600), .B(n11599), .Z(n11607) );
  XNOR U12472 ( .A(n11608), .B(n11607), .Z(n11610) );
  XOR U12473 ( .A(n11609), .B(n11610), .Z(n11616) );
  XNOR U12474 ( .A(n11615), .B(n11616), .Z(n11627) );
  XOR U12475 ( .A(n11628), .B(n11627), .Z(n11582) );
  NANDN U12476 ( .A(n11512), .B(n11511), .Z(n11516) );
  NANDN U12477 ( .A(n11514), .B(n11513), .Z(n11515) );
  AND U12478 ( .A(n11516), .B(n11515), .Z(n11579) );
  NAND U12479 ( .A(n11518), .B(n11517), .Z(n11522) );
  ANDN U12480 ( .B(n11520), .A(n11519), .Z(n11521) );
  ANDN U12481 ( .B(n11522), .A(n11521), .Z(n11689) );
  NANDN U12482 ( .A(n11524), .B(n11523), .Z(n11528) );
  NANDN U12483 ( .A(n11526), .B(n11525), .Z(n11527) );
  AND U12484 ( .A(n11528), .B(n11527), .Z(n11688) );
  AND U12485 ( .A(x[238]), .B(y[1899]), .Z(n11645) );
  NAND U12486 ( .A(x[226]), .B(y[1911]), .Z(n11646) );
  XNOR U12487 ( .A(n11645), .B(n11646), .Z(n11647) );
  NAND U12488 ( .A(x[227]), .B(y[1910]), .Z(n11648) );
  XNOR U12489 ( .A(n11647), .B(n11648), .Z(n11687) );
  XOR U12490 ( .A(n11688), .B(n11687), .Z(n11690) );
  XOR U12491 ( .A(n11689), .B(n11690), .Z(n11580) );
  XNOR U12492 ( .A(n11579), .B(n11580), .Z(n11581) );
  XNOR U12493 ( .A(n11582), .B(n11581), .Z(n11585) );
  NANDN U12494 ( .A(n11530), .B(n11529), .Z(n11534) );
  NAND U12495 ( .A(n11532), .B(n11531), .Z(n11533) );
  NAND U12496 ( .A(n11534), .B(n11533), .Z(n11586) );
  XNOR U12497 ( .A(n11585), .B(n11586), .Z(n11587) );
  NANDN U12498 ( .A(n11536), .B(n11535), .Z(n11540) );
  OR U12499 ( .A(n11538), .B(n11537), .Z(n11539) );
  NAND U12500 ( .A(n11540), .B(n11539), .Z(n11588) );
  XOR U12501 ( .A(n11587), .B(n11588), .Z(n11567) );
  NAND U12502 ( .A(n11542), .B(n11541), .Z(n11546) );
  NAND U12503 ( .A(n11544), .B(n11543), .Z(n11545) );
  AND U12504 ( .A(n11546), .B(n11545), .Z(n11568) );
  XOR U12505 ( .A(n11567), .B(n11568), .Z(n11570) );
  XNOR U12506 ( .A(n11569), .B(n11570), .Z(n11713) );
  NAND U12507 ( .A(n11548), .B(n11547), .Z(n11552) );
  NAND U12508 ( .A(n11550), .B(n11549), .Z(n11551) );
  NAND U12509 ( .A(n11552), .B(n11551), .Z(n11712) );
  XOR U12510 ( .A(n11713), .B(n11712), .Z(n11714) );
  XNOR U12511 ( .A(n11715), .B(n11714), .Z(n11708) );
  OR U12512 ( .A(n11555), .B(n11553), .Z(n11559) );
  ANDN U12513 ( .B(n11555), .A(n11554), .Z(n11557) );
  OR U12514 ( .A(n11557), .B(n11556), .Z(n11558) );
  AND U12515 ( .A(n11559), .B(n11558), .Z(n11706) );
  NAND U12516 ( .A(n11561), .B(n11560), .Z(n11565) );
  NAND U12517 ( .A(n11563), .B(n11562), .Z(n11564) );
  AND U12518 ( .A(n11565), .B(n11564), .Z(n11707) );
  IV U12519 ( .A(n11707), .Z(n11705) );
  XOR U12520 ( .A(n11706), .B(n11705), .Z(n11566) );
  XNOR U12521 ( .A(n11708), .B(n11566), .Z(N250) );
  NAND U12522 ( .A(n11568), .B(n11567), .Z(n11572) );
  NAND U12523 ( .A(n11570), .B(n11569), .Z(n11571) );
  NAND U12524 ( .A(n11572), .B(n11571), .Z(n11870) );
  NAND U12525 ( .A(n11574), .B(n11573), .Z(n11578) );
  NAND U12526 ( .A(n11576), .B(n11575), .Z(n11577) );
  AND U12527 ( .A(n11578), .B(n11577), .Z(n11871) );
  XOR U12528 ( .A(n11870), .B(n11871), .Z(n11873) );
  NANDN U12529 ( .A(n11580), .B(n11579), .Z(n11584) );
  NANDN U12530 ( .A(n11582), .B(n11581), .Z(n11583) );
  AND U12531 ( .A(n11584), .B(n11583), .Z(n11719) );
  NANDN U12532 ( .A(n11586), .B(n11585), .Z(n11590) );
  NANDN U12533 ( .A(n11588), .B(n11587), .Z(n11589) );
  NAND U12534 ( .A(n11590), .B(n11589), .Z(n11720) );
  XNOR U12535 ( .A(n11719), .B(n11720), .Z(n11721) );
  NANDN U12536 ( .A(n11592), .B(n11591), .Z(n11596) );
  NANDN U12537 ( .A(n11594), .B(n11593), .Z(n11595) );
  AND U12538 ( .A(n11596), .B(n11595), .Z(n11864) );
  AND U12539 ( .A(x[226]), .B(y[1912]), .Z(n11793) );
  XOR U12540 ( .A(n11794), .B(n11793), .Z(n11795) );
  NAND U12541 ( .A(x[248]), .B(y[1890]), .Z(n11796) );
  XNOR U12542 ( .A(n11795), .B(n11796), .Z(n11829) );
  NANDN U12543 ( .A(n11598), .B(n11597), .Z(n11602) );
  NANDN U12544 ( .A(n11600), .B(n11599), .Z(n11601) );
  NAND U12545 ( .A(n11602), .B(n11601), .Z(n11830) );
  XNOR U12546 ( .A(n11829), .B(n11830), .Z(n11831) );
  XNOR U12547 ( .A(n11831), .B(n11832), .Z(n11732) );
  OR U12548 ( .A(n11608), .B(n11607), .Z(n11612) );
  NANDN U12549 ( .A(n11610), .B(n11609), .Z(n11611) );
  AND U12550 ( .A(n11612), .B(n11611), .Z(n11731) );
  XNOR U12551 ( .A(n11732), .B(n11731), .Z(n11733) );
  NANDN U12552 ( .A(n11614), .B(n11613), .Z(n11618) );
  NANDN U12553 ( .A(n11616), .B(n11615), .Z(n11617) );
  NAND U12554 ( .A(n11618), .B(n11617), .Z(n11734) );
  XNOR U12555 ( .A(n11733), .B(n11734), .Z(n11728) );
  NAND U12556 ( .A(n11620), .B(n11619), .Z(n11624) );
  NAND U12557 ( .A(n11622), .B(n11621), .Z(n11623) );
  AND U12558 ( .A(n11624), .B(n11623), .Z(n11726) );
  NANDN U12559 ( .A(n11626), .B(n11625), .Z(n11630) );
  NAND U12560 ( .A(n11628), .B(n11627), .Z(n11629) );
  AND U12561 ( .A(n11630), .B(n11629), .Z(n11725) );
  XNOR U12562 ( .A(n11726), .B(n11725), .Z(n11727) );
  XOR U12563 ( .A(n11728), .B(n11727), .Z(n11862) );
  NANDN U12564 ( .A(n11632), .B(n11631), .Z(n11636) );
  NANDN U12565 ( .A(n11634), .B(n11633), .Z(n11635) );
  AND U12566 ( .A(n11636), .B(n11635), .Z(n11778) );
  AND U12567 ( .A(y[1908]), .B(x[230]), .Z(n11638) );
  NAND U12568 ( .A(y[1906]), .B(x[232]), .Z(n11637) );
  XNOR U12569 ( .A(n11638), .B(n11637), .Z(n11757) );
  AND U12570 ( .A(x[233]), .B(y[1905]), .Z(n11756) );
  XOR U12571 ( .A(n11757), .B(n11756), .Z(n11737) );
  AND U12572 ( .A(x[231]), .B(y[1907]), .Z(n11738) );
  XOR U12573 ( .A(n11737), .B(n11738), .Z(n11740) );
  AND U12574 ( .A(x[236]), .B(y[1902]), .Z(n11927) );
  AND U12575 ( .A(x[229]), .B(y[1909]), .Z(n11844) );
  XOR U12576 ( .A(n11927), .B(n11844), .Z(n11846) );
  AND U12577 ( .A(x[234]), .B(y[1904]), .Z(n11845) );
  XOR U12578 ( .A(n11846), .B(n11845), .Z(n11739) );
  XOR U12579 ( .A(n11740), .B(n11739), .Z(n11819) );
  NANDN U12580 ( .A(n11640), .B(n11639), .Z(n11644) );
  NANDN U12581 ( .A(n11642), .B(n11641), .Z(n11643) );
  AND U12582 ( .A(n11644), .B(n11643), .Z(n11818) );
  NANDN U12583 ( .A(n11646), .B(n11645), .Z(n11650) );
  NANDN U12584 ( .A(n11648), .B(n11647), .Z(n11649) );
  NAND U12585 ( .A(n11650), .B(n11649), .Z(n11817) );
  XOR U12586 ( .A(n11818), .B(n11817), .Z(n11820) );
  XNOR U12587 ( .A(n11819), .B(n11820), .Z(n11856) );
  NANDN U12588 ( .A(n11652), .B(n11651), .Z(n11656) );
  NANDN U12589 ( .A(n11654), .B(n11653), .Z(n11655) );
  AND U12590 ( .A(n11656), .B(n11655), .Z(n11855) );
  XNOR U12591 ( .A(n11856), .B(n11855), .Z(n11858) );
  NANDN U12592 ( .A(n11658), .B(n11657), .Z(n11662) );
  NANDN U12593 ( .A(n11660), .B(n11659), .Z(n11661) );
  AND U12594 ( .A(n11662), .B(n11661), .Z(n11781) );
  NANDN U12595 ( .A(n11664), .B(n11663), .Z(n11668) );
  NANDN U12596 ( .A(n11666), .B(n11665), .Z(n11667) );
  NAND U12597 ( .A(n11668), .B(n11667), .Z(n11782) );
  XNOR U12598 ( .A(n11781), .B(n11782), .Z(n11783) );
  ANDN U12599 ( .B(o[121]), .A(n11669), .Z(n11749) );
  AND U12600 ( .A(x[238]), .B(y[1900]), .Z(n11750) );
  XOR U12601 ( .A(n11749), .B(n11750), .Z(n11751) );
  AND U12602 ( .A(x[225]), .B(y[1913]), .Z(n11752) );
  XOR U12603 ( .A(n11751), .B(n11752), .Z(n11836) );
  AND U12604 ( .A(x[249]), .B(y[1889]), .Z(n11760) );
  XOR U12605 ( .A(o[122]), .B(n11760), .Z(n11850) );
  AND U12606 ( .A(x[250]), .B(y[1888]), .Z(n11849) );
  XOR U12607 ( .A(n11850), .B(n11849), .Z(n11852) );
  AND U12608 ( .A(x[224]), .B(y[1914]), .Z(n11851) );
  XOR U12609 ( .A(n11852), .B(n11851), .Z(n11835) );
  XOR U12610 ( .A(n11836), .B(n11835), .Z(n11838) );
  NANDN U12611 ( .A(n11671), .B(n11670), .Z(n11675) );
  NANDN U12612 ( .A(n11673), .B(n11672), .Z(n11674) );
  AND U12613 ( .A(n11675), .B(n11674), .Z(n11837) );
  XNOR U12614 ( .A(n11838), .B(n11837), .Z(n11784) );
  XNOR U12615 ( .A(n11783), .B(n11784), .Z(n11826) );
  AND U12616 ( .A(x[245]), .B(y[1893]), .Z(n11743) );
  NANDN U12617 ( .A(n11676), .B(n11743), .Z(n11680) );
  NAND U12618 ( .A(n11678), .B(n11677), .Z(n11679) );
  AND U12619 ( .A(n11680), .B(n11679), .Z(n11814) );
  XOR U12620 ( .A(n11744), .B(n11743), .Z(n11745) );
  AND U12621 ( .A(x[244]), .B(y[1894]), .Z(n11746) );
  XOR U12622 ( .A(n11745), .B(n11746), .Z(n11811) );
  NAND U12623 ( .A(x[247]), .B(y[1891]), .Z(n11800) );
  XNOR U12624 ( .A(n11799), .B(n11800), .Z(n11802) );
  AND U12625 ( .A(x[246]), .B(y[1892]), .Z(n11801) );
  XNOR U12626 ( .A(n11802), .B(n11801), .Z(n11812) );
  XNOR U12627 ( .A(n11811), .B(n11812), .Z(n11813) );
  XNOR U12628 ( .A(n11814), .B(n11813), .Z(n11824) );
  AND U12629 ( .A(x[228]), .B(y[1910]), .Z(n11805) );
  XOR U12630 ( .A(n11806), .B(n11805), .Z(n11808) );
  XOR U12631 ( .A(n11808), .B(n11807), .Z(n11787) );
  AND U12632 ( .A(x[235]), .B(y[1903]), .Z(n11761) );
  AND U12633 ( .A(x[227]), .B(y[1911]), .Z(n11762) );
  XOR U12634 ( .A(n11761), .B(n11762), .Z(n11764) );
  AND U12635 ( .A(x[243]), .B(y[1895]), .Z(n11763) );
  XNOR U12636 ( .A(n11764), .B(n11763), .Z(n11788) );
  XNOR U12637 ( .A(n11787), .B(n11788), .Z(n11790) );
  NANDN U12638 ( .A(n11682), .B(n11681), .Z(n11686) );
  NANDN U12639 ( .A(n11684), .B(n11683), .Z(n11685) );
  AND U12640 ( .A(n11686), .B(n11685), .Z(n11789) );
  XNOR U12641 ( .A(n11790), .B(n11789), .Z(n11823) );
  XNOR U12642 ( .A(n11824), .B(n11823), .Z(n11825) );
  XNOR U12643 ( .A(n11826), .B(n11825), .Z(n11857) );
  XOR U12644 ( .A(n11858), .B(n11857), .Z(n11776) );
  NANDN U12645 ( .A(n11688), .B(n11687), .Z(n11692) );
  OR U12646 ( .A(n11690), .B(n11689), .Z(n11691) );
  NAND U12647 ( .A(n11692), .B(n11691), .Z(n11772) );
  NANDN U12648 ( .A(n11694), .B(n11693), .Z(n11698) );
  NANDN U12649 ( .A(n11696), .B(n11695), .Z(n11697) );
  NAND U12650 ( .A(n11698), .B(n11697), .Z(n11770) );
  OR U12651 ( .A(n11700), .B(n11699), .Z(n11704) );
  NANDN U12652 ( .A(n11702), .B(n11701), .Z(n11703) );
  NAND U12653 ( .A(n11704), .B(n11703), .Z(n11769) );
  XOR U12654 ( .A(n11770), .B(n11769), .Z(n11771) );
  XOR U12655 ( .A(n11772), .B(n11771), .Z(n11775) );
  XNOR U12656 ( .A(n11776), .B(n11775), .Z(n11777) );
  XNOR U12657 ( .A(n11778), .B(n11777), .Z(n11861) );
  XNOR U12658 ( .A(n11862), .B(n11861), .Z(n11863) );
  XOR U12659 ( .A(n11864), .B(n11863), .Z(n11722) );
  XNOR U12660 ( .A(n11721), .B(n11722), .Z(n11872) );
  XNOR U12661 ( .A(n11873), .B(n11872), .Z(n11869) );
  NANDN U12662 ( .A(n11705), .B(n11706), .Z(n11711) );
  NOR U12663 ( .A(n11707), .B(n11706), .Z(n11709) );
  OR U12664 ( .A(n11709), .B(n11708), .Z(n11710) );
  AND U12665 ( .A(n11711), .B(n11710), .Z(n11867) );
  NAND U12666 ( .A(n11713), .B(n11712), .Z(n11717) );
  NAND U12667 ( .A(n11715), .B(n11714), .Z(n11716) );
  AND U12668 ( .A(n11717), .B(n11716), .Z(n11868) );
  XOR U12669 ( .A(n11867), .B(n11868), .Z(n11718) );
  XNOR U12670 ( .A(n11869), .B(n11718), .Z(N251) );
  NANDN U12671 ( .A(n11720), .B(n11719), .Z(n11724) );
  NANDN U12672 ( .A(n11722), .B(n11721), .Z(n11723) );
  AND U12673 ( .A(n11724), .B(n11723), .Z(n12029) );
  NANDN U12674 ( .A(n11726), .B(n11725), .Z(n11730) );
  NAND U12675 ( .A(n11728), .B(n11727), .Z(n11729) );
  NAND U12676 ( .A(n11730), .B(n11729), .Z(n11883) );
  NANDN U12677 ( .A(n11732), .B(n11731), .Z(n11736) );
  NANDN U12678 ( .A(n11734), .B(n11733), .Z(n11735) );
  NAND U12679 ( .A(n11736), .B(n11735), .Z(n11888) );
  NAND U12680 ( .A(n11738), .B(n11737), .Z(n11742) );
  NAND U12681 ( .A(n11740), .B(n11739), .Z(n11741) );
  NAND U12682 ( .A(n11742), .B(n11741), .Z(n12014) );
  AND U12683 ( .A(n11744), .B(n11743), .Z(n11748) );
  NAND U12684 ( .A(n11746), .B(n11745), .Z(n11747) );
  NANDN U12685 ( .A(n11748), .B(n11747), .Z(n11945) );
  NAND U12686 ( .A(n11750), .B(n11749), .Z(n11754) );
  NAND U12687 ( .A(n11752), .B(n11751), .Z(n11753) );
  NAND U12688 ( .A(n11754), .B(n11753), .Z(n11944) );
  XOR U12689 ( .A(n11945), .B(n11944), .Z(n11946) );
  AND U12690 ( .A(y[1908]), .B(x[232]), .Z(n11987) );
  NAND U12691 ( .A(n11755), .B(n11987), .Z(n11759) );
  NAND U12692 ( .A(n11757), .B(n11756), .Z(n11758) );
  NAND U12693 ( .A(n11759), .B(n11758), .Z(n11907) );
  AND U12694 ( .A(o[122]), .B(n11760), .Z(n11941) );
  AND U12695 ( .A(x[225]), .B(y[1914]), .Z(n11939) );
  AND U12696 ( .A(x[238]), .B(y[1901]), .Z(n11938) );
  XOR U12697 ( .A(n11939), .B(n11938), .Z(n11940) );
  XOR U12698 ( .A(n11941), .B(n11940), .Z(n11906) );
  AND U12699 ( .A(x[241]), .B(y[1898]), .Z(n11974) );
  AND U12700 ( .A(x[228]), .B(y[1911]), .Z(n11973) );
  XOR U12701 ( .A(n11974), .B(n11973), .Z(n11976) );
  AND U12702 ( .A(x[229]), .B(y[1910]), .Z(n11975) );
  XOR U12703 ( .A(n11976), .B(n11975), .Z(n11905) );
  XOR U12704 ( .A(n11906), .B(n11905), .Z(n11908) );
  XNOR U12705 ( .A(n11907), .B(n11908), .Z(n11947) );
  NAND U12706 ( .A(n11762), .B(n11761), .Z(n11766) );
  NAND U12707 ( .A(n11764), .B(n11763), .Z(n11765) );
  NAND U12708 ( .A(n11766), .B(n11765), .Z(n11952) );
  AND U12709 ( .A(x[231]), .B(y[1908]), .Z(n11964) );
  AND U12710 ( .A(y[1891]), .B(x[248]), .Z(n11768) );
  XOR U12711 ( .A(n11768), .B(n11767), .Z(n11963) );
  XOR U12712 ( .A(n11964), .B(n11963), .Z(n11951) );
  AND U12713 ( .A(x[246]), .B(y[1893]), .Z(n11924) );
  AND U12714 ( .A(x[232]), .B(y[1907]), .Z(n11922) );
  AND U12715 ( .A(x[247]), .B(y[1892]), .Z(n11921) );
  XOR U12716 ( .A(n11922), .B(n11921), .Z(n11923) );
  XOR U12717 ( .A(n11924), .B(n11923), .Z(n11950) );
  XOR U12718 ( .A(n11951), .B(n11950), .Z(n11953) );
  XOR U12719 ( .A(n11952), .B(n11953), .Z(n12012) );
  XOR U12720 ( .A(n12013), .B(n12012), .Z(n12015) );
  XNOR U12721 ( .A(n12014), .B(n12015), .Z(n11887) );
  XOR U12722 ( .A(n11888), .B(n11887), .Z(n11890) );
  NAND U12723 ( .A(n11770), .B(n11769), .Z(n11774) );
  NAND U12724 ( .A(n11772), .B(n11771), .Z(n11773) );
  AND U12725 ( .A(n11774), .B(n11773), .Z(n11889) );
  XOR U12726 ( .A(n11890), .B(n11889), .Z(n11884) );
  XOR U12727 ( .A(n11883), .B(n11884), .Z(n11886) );
  NANDN U12728 ( .A(n11776), .B(n11775), .Z(n11780) );
  NANDN U12729 ( .A(n11778), .B(n11777), .Z(n11779) );
  AND U12730 ( .A(n11780), .B(n11779), .Z(n11879) );
  NANDN U12731 ( .A(n11782), .B(n11781), .Z(n11786) );
  NANDN U12732 ( .A(n11784), .B(n11783), .Z(n11785) );
  NAND U12733 ( .A(n11786), .B(n11785), .Z(n12002) );
  NANDN U12734 ( .A(n11788), .B(n11787), .Z(n11792) );
  NAND U12735 ( .A(n11790), .B(n11789), .Z(n11791) );
  NAND U12736 ( .A(n11792), .B(n11791), .Z(n12000) );
  AND U12737 ( .A(n11794), .B(n11793), .Z(n11798) );
  NANDN U12738 ( .A(n11796), .B(n11795), .Z(n11797) );
  NANDN U12739 ( .A(n11798), .B(n11797), .Z(n11900) );
  NANDN U12740 ( .A(n11800), .B(n11799), .Z(n11804) );
  NAND U12741 ( .A(n11802), .B(n11801), .Z(n11803) );
  NAND U12742 ( .A(n11804), .B(n11803), .Z(n11899) );
  XOR U12743 ( .A(n11900), .B(n11899), .Z(n11901) );
  AND U12744 ( .A(n11806), .B(n11805), .Z(n11810) );
  NAND U12745 ( .A(n11808), .B(n11807), .Z(n11809) );
  NANDN U12746 ( .A(n11810), .B(n11809), .Z(n11913) );
  AND U12747 ( .A(x[224]), .B(y[1915]), .Z(n11980) );
  AND U12748 ( .A(x[251]), .B(y[1888]), .Z(n11979) );
  XOR U12749 ( .A(n11980), .B(n11979), .Z(n11982) );
  AND U12750 ( .A(x[250]), .B(y[1889]), .Z(n11985) );
  XOR U12751 ( .A(n11985), .B(o[123]), .Z(n11981) );
  XOR U12752 ( .A(n11982), .B(n11981), .Z(n11912) );
  AND U12753 ( .A(x[233]), .B(y[1906]), .Z(n11989) );
  AND U12754 ( .A(x[245]), .B(y[1894]), .Z(n11988) );
  XOR U12755 ( .A(n11989), .B(n11988), .Z(n11991) );
  AND U12756 ( .A(x[242]), .B(y[1897]), .Z(n11990) );
  XOR U12757 ( .A(n11991), .B(n11990), .Z(n11911) );
  XOR U12758 ( .A(n11912), .B(n11911), .Z(n11914) );
  XNOR U12759 ( .A(n11913), .B(n11914), .Z(n11902) );
  XOR U12760 ( .A(n12000), .B(n12001), .Z(n12003) );
  XOR U12761 ( .A(n12002), .B(n12003), .Z(n12021) );
  NANDN U12762 ( .A(n11812), .B(n11811), .Z(n11816) );
  NANDN U12763 ( .A(n11814), .B(n11813), .Z(n11815) );
  AND U12764 ( .A(n11816), .B(n11815), .Z(n12019) );
  NANDN U12765 ( .A(n11818), .B(n11817), .Z(n11822) );
  NANDN U12766 ( .A(n11820), .B(n11819), .Z(n11821) );
  AND U12767 ( .A(n11822), .B(n11821), .Z(n12018) );
  XOR U12768 ( .A(n12019), .B(n12018), .Z(n12020) );
  NANDN U12769 ( .A(n11824), .B(n11823), .Z(n11828) );
  NANDN U12770 ( .A(n11826), .B(n11825), .Z(n11827) );
  AND U12771 ( .A(n11828), .B(n11827), .Z(n12006) );
  NANDN U12772 ( .A(n11830), .B(n11829), .Z(n11834) );
  NANDN U12773 ( .A(n11832), .B(n11831), .Z(n11833) );
  NAND U12774 ( .A(n11834), .B(n11833), .Z(n11996) );
  NAND U12775 ( .A(n11836), .B(n11835), .Z(n11840) );
  NAND U12776 ( .A(n11838), .B(n11837), .Z(n11839) );
  NAND U12777 ( .A(n11840), .B(n11839), .Z(n11994) );
  AND U12778 ( .A(x[230]), .B(y[1909]), .Z(n11970) );
  AND U12779 ( .A(x[249]), .B(y[1890]), .Z(n11968) );
  AND U12780 ( .A(x[243]), .B(y[1896]), .Z(n11967) );
  XOR U12781 ( .A(n11968), .B(n11967), .Z(n11969) );
  XOR U12782 ( .A(n11970), .B(n11969), .Z(n11957) );
  AND U12783 ( .A(x[239]), .B(y[1900]), .Z(n11933) );
  AND U12784 ( .A(x[226]), .B(y[1913]), .Z(n11932) );
  XOR U12785 ( .A(n11933), .B(n11932), .Z(n11935) );
  AND U12786 ( .A(x[227]), .B(y[1912]), .Z(n11934) );
  XOR U12787 ( .A(n11935), .B(n11934), .Z(n11956) );
  XOR U12788 ( .A(n11957), .B(n11956), .Z(n11958) );
  NAND U12789 ( .A(x[240]), .B(y[1899]), .Z(n11917) );
  XOR U12790 ( .A(n11917), .B(n11841), .Z(n11920) );
  XOR U12791 ( .A(n11919), .B(n11920), .Z(n11929) );
  AND U12792 ( .A(y[1902]), .B(x[237]), .Z(n11843) );
  AND U12793 ( .A(y[1903]), .B(x[236]), .Z(n11842) );
  XOR U12794 ( .A(n11843), .B(n11842), .Z(n11928) );
  XNOR U12795 ( .A(n11958), .B(n11959), .Z(n11896) );
  AND U12796 ( .A(n11927), .B(n11844), .Z(n11848) );
  NAND U12797 ( .A(n11846), .B(n11845), .Z(n11847) );
  NANDN U12798 ( .A(n11848), .B(n11847), .Z(n11894) );
  NAND U12799 ( .A(n11850), .B(n11849), .Z(n11854) );
  NAND U12800 ( .A(n11852), .B(n11851), .Z(n11853) );
  NAND U12801 ( .A(n11854), .B(n11853), .Z(n11893) );
  XOR U12802 ( .A(n11894), .B(n11893), .Z(n11895) );
  XOR U12803 ( .A(n11896), .B(n11895), .Z(n11995) );
  XNOR U12804 ( .A(n11994), .B(n11995), .Z(n11997) );
  XNOR U12805 ( .A(n12006), .B(n12007), .Z(n12009) );
  NANDN U12806 ( .A(n11856), .B(n11855), .Z(n11860) );
  NAND U12807 ( .A(n11858), .B(n11857), .Z(n11859) );
  AND U12808 ( .A(n11860), .B(n11859), .Z(n12008) );
  XNOR U12809 ( .A(n12009), .B(n12008), .Z(n11877) );
  XNOR U12810 ( .A(n11878), .B(n11877), .Z(n11880) );
  XNOR U12811 ( .A(n11879), .B(n11880), .Z(n11885) );
  XOR U12812 ( .A(n11886), .B(n11885), .Z(n12028) );
  NANDN U12813 ( .A(n11862), .B(n11861), .Z(n11866) );
  NANDN U12814 ( .A(n11864), .B(n11863), .Z(n11865) );
  NAND U12815 ( .A(n11866), .B(n11865), .Z(n12027) );
  XOR U12816 ( .A(n12028), .B(n12027), .Z(n12030) );
  XNOR U12817 ( .A(n12029), .B(n12030), .Z(n12026) );
  NAND U12818 ( .A(n11871), .B(n11870), .Z(n11875) );
  NAND U12819 ( .A(n11873), .B(n11872), .Z(n11874) );
  NAND U12820 ( .A(n11875), .B(n11874), .Z(n12024) );
  XNOR U12821 ( .A(n12025), .B(n12024), .Z(n11876) );
  XNOR U12822 ( .A(n12026), .B(n11876), .Z(N252) );
  NAND U12823 ( .A(n11878), .B(n11877), .Z(n11882) );
  NANDN U12824 ( .A(n11880), .B(n11879), .Z(n11881) );
  AND U12825 ( .A(n11882), .B(n11881), .Z(n12035) );
  XOR U12826 ( .A(n12035), .B(n12034), .Z(n12037) );
  NAND U12827 ( .A(n11888), .B(n11887), .Z(n11892) );
  NAND U12828 ( .A(n11890), .B(n11889), .Z(n11891) );
  AND U12829 ( .A(n11892), .B(n11891), .Z(n12041) );
  NAND U12830 ( .A(n11894), .B(n11893), .Z(n11898) );
  NAND U12831 ( .A(n11896), .B(n11895), .Z(n11897) );
  NAND U12832 ( .A(n11898), .B(n11897), .Z(n12053) );
  NAND U12833 ( .A(n11900), .B(n11899), .Z(n11904) );
  NANDN U12834 ( .A(n11902), .B(n11901), .Z(n11903) );
  NAND U12835 ( .A(n11904), .B(n11903), .Z(n12158) );
  NAND U12836 ( .A(n11906), .B(n11905), .Z(n11910) );
  NAND U12837 ( .A(n11908), .B(n11907), .Z(n11909) );
  NAND U12838 ( .A(n11910), .B(n11909), .Z(n12157) );
  NAND U12839 ( .A(n11912), .B(n11911), .Z(n11916) );
  NAND U12840 ( .A(n11914), .B(n11913), .Z(n11915) );
  NAND U12841 ( .A(n11916), .B(n11915), .Z(n12156) );
  XOR U12842 ( .A(n12157), .B(n12156), .Z(n12159) );
  XOR U12843 ( .A(n12158), .B(n12159), .Z(n12054) );
  XOR U12844 ( .A(n12053), .B(n12054), .Z(n12056) );
  AND U12845 ( .A(x[239]), .B(y[1901]), .Z(n12133) );
  AND U12846 ( .A(x[251]), .B(y[1889]), .Z(n12117) );
  XOR U12847 ( .A(o[124]), .B(n12117), .Z(n12131) );
  AND U12848 ( .A(x[250]), .B(y[1890]), .Z(n12130) );
  XOR U12849 ( .A(n12131), .B(n12130), .Z(n12132) );
  XOR U12850 ( .A(n12133), .B(n12132), .Z(n12119) );
  AND U12851 ( .A(x[231]), .B(y[1909]), .Z(n12101) );
  AND U12852 ( .A(x[236]), .B(y[1904]), .Z(n12100) );
  XOR U12853 ( .A(n12101), .B(n12100), .Z(n12103) );
  AND U12854 ( .A(x[235]), .B(y[1905]), .Z(n12102) );
  XNOR U12855 ( .A(n12103), .B(n12102), .Z(n12118) );
  XOR U12856 ( .A(n12120), .B(n12121), .Z(n12163) );
  AND U12857 ( .A(x[241]), .B(y[1899]), .Z(n12066) );
  AND U12858 ( .A(x[246]), .B(y[1894]), .Z(n12065) );
  XOR U12859 ( .A(n12066), .B(n12065), .Z(n12068) );
  AND U12860 ( .A(x[228]), .B(y[1912]), .Z(n12067) );
  XOR U12861 ( .A(n12068), .B(n12067), .Z(n12139) );
  AND U12862 ( .A(x[230]), .B(y[1910]), .Z(n12293) );
  AND U12863 ( .A(x[243]), .B(y[1897]), .Z(n12106) );
  XOR U12864 ( .A(n12293), .B(n12106), .Z(n12108) );
  XOR U12865 ( .A(n12108), .B(n12107), .Z(n12138) );
  XOR U12866 ( .A(n12139), .B(n12138), .Z(n12141) );
  NAND U12867 ( .A(n11922), .B(n11921), .Z(n11926) );
  NAND U12868 ( .A(n11924), .B(n11923), .Z(n11925) );
  NAND U12869 ( .A(n11926), .B(n11925), .Z(n12140) );
  XOR U12870 ( .A(n12141), .B(n12140), .Z(n12162) );
  NAND U12871 ( .A(n11927), .B(n12125), .Z(n11931) );
  NANDN U12872 ( .A(n11929), .B(n11928), .Z(n11930) );
  NAND U12873 ( .A(n11931), .B(n11930), .Z(n12084) );
  NAND U12874 ( .A(n11933), .B(n11932), .Z(n11937) );
  NAND U12875 ( .A(n11935), .B(n11934), .Z(n11936) );
  NAND U12876 ( .A(n11937), .B(n11936), .Z(n12083) );
  NAND U12877 ( .A(n11939), .B(n11938), .Z(n11943) );
  NAND U12878 ( .A(n11941), .B(n11940), .Z(n11942) );
  NAND U12879 ( .A(n11943), .B(n11942), .Z(n12082) );
  XOR U12880 ( .A(n12083), .B(n12082), .Z(n12085) );
  XOR U12881 ( .A(n12084), .B(n12085), .Z(n12164) );
  XOR U12882 ( .A(n12165), .B(n12164), .Z(n12055) );
  XNOR U12883 ( .A(n12056), .B(n12055), .Z(n12189) );
  NAND U12884 ( .A(n11945), .B(n11944), .Z(n11949) );
  NANDN U12885 ( .A(n11947), .B(n11946), .Z(n11948) );
  NAND U12886 ( .A(n11949), .B(n11948), .Z(n12146) );
  NAND U12887 ( .A(n11951), .B(n11950), .Z(n11955) );
  NAND U12888 ( .A(n11953), .B(n11952), .Z(n11954) );
  NAND U12889 ( .A(n11955), .B(n11954), .Z(n12145) );
  NAND U12890 ( .A(n11957), .B(n11956), .Z(n11961) );
  NANDN U12891 ( .A(n11959), .B(n11958), .Z(n11960) );
  NAND U12892 ( .A(n11961), .B(n11960), .Z(n12144) );
  XOR U12893 ( .A(n12145), .B(n12144), .Z(n12147) );
  XOR U12894 ( .A(n12146), .B(n12147), .Z(n12187) );
  AND U12895 ( .A(x[248]), .B(y[1895]), .Z(n12470) );
  AND U12896 ( .A(x[244]), .B(y[1891]), .Z(n11962) );
  NAND U12897 ( .A(n12470), .B(n11962), .Z(n11966) );
  NAND U12898 ( .A(n11964), .B(n11963), .Z(n11965) );
  NAND U12899 ( .A(n11966), .B(n11965), .Z(n12182) );
  AND U12900 ( .A(x[249]), .B(y[1891]), .Z(n12096) );
  XOR U12901 ( .A(n12097), .B(n12096), .Z(n12095) );
  AND U12902 ( .A(x[225]), .B(y[1915]), .Z(n12094) );
  XOR U12903 ( .A(n12095), .B(n12094), .Z(n12181) );
  AND U12904 ( .A(x[240]), .B(y[1900]), .Z(n12089) );
  AND U12905 ( .A(x[248]), .B(y[1892]), .Z(n12088) );
  XOR U12906 ( .A(n12089), .B(n12088), .Z(n12091) );
  AND U12907 ( .A(x[226]), .B(y[1914]), .Z(n12090) );
  XOR U12908 ( .A(n12091), .B(n12090), .Z(n12180) );
  XOR U12909 ( .A(n12181), .B(n12180), .Z(n12183) );
  XOR U12910 ( .A(n12182), .B(n12183), .Z(n12153) );
  NAND U12911 ( .A(n11968), .B(n11967), .Z(n11972) );
  NAND U12912 ( .A(n11970), .B(n11969), .Z(n11971) );
  NAND U12913 ( .A(n11972), .B(n11971), .Z(n12176) );
  AND U12914 ( .A(x[227]), .B(y[1913]), .Z(n12124) );
  XOR U12915 ( .A(n12125), .B(n12124), .Z(n12127) );
  AND U12916 ( .A(x[247]), .B(y[1893]), .Z(n12126) );
  XOR U12917 ( .A(n12127), .B(n12126), .Z(n12175) );
  AND U12918 ( .A(x[229]), .B(y[1911]), .Z(n12112) );
  AND U12919 ( .A(x[245]), .B(y[1895]), .Z(n12111) );
  XOR U12920 ( .A(n12112), .B(n12111), .Z(n12114) );
  AND U12921 ( .A(x[244]), .B(y[1896]), .Z(n12113) );
  XOR U12922 ( .A(n12114), .B(n12113), .Z(n12174) );
  XOR U12923 ( .A(n12175), .B(n12174), .Z(n12177) );
  XOR U12924 ( .A(n12176), .B(n12177), .Z(n12151) );
  NAND U12925 ( .A(n11974), .B(n11973), .Z(n11978) );
  NAND U12926 ( .A(n11976), .B(n11975), .Z(n11977) );
  NAND U12927 ( .A(n11978), .B(n11977), .Z(n12169) );
  NAND U12928 ( .A(n11980), .B(n11979), .Z(n11984) );
  NAND U12929 ( .A(n11982), .B(n11981), .Z(n11983) );
  NAND U12930 ( .A(n11984), .B(n11983), .Z(n12168) );
  XOR U12931 ( .A(n12169), .B(n12168), .Z(n12171) );
  AND U12932 ( .A(n11985), .B(o[123]), .Z(n12074) );
  AND U12933 ( .A(x[224]), .B(y[1916]), .Z(n12072) );
  AND U12934 ( .A(x[252]), .B(y[1888]), .Z(n12071) );
  XOR U12935 ( .A(n12072), .B(n12071), .Z(n12073) );
  XOR U12936 ( .A(n12074), .B(n12073), .Z(n12060) );
  NAND U12937 ( .A(y[1906]), .B(x[234]), .Z(n11986) );
  XNOR U12938 ( .A(n11987), .B(n11986), .Z(n12079) );
  AND U12939 ( .A(x[233]), .B(y[1907]), .Z(n12078) );
  XOR U12940 ( .A(n12079), .B(n12078), .Z(n12059) );
  XOR U12941 ( .A(n12060), .B(n12059), .Z(n12062) );
  NAND U12942 ( .A(n11989), .B(n11988), .Z(n11993) );
  NAND U12943 ( .A(n11991), .B(n11990), .Z(n11992) );
  NAND U12944 ( .A(n11993), .B(n11992), .Z(n12061) );
  XOR U12945 ( .A(n12062), .B(n12061), .Z(n12170) );
  XNOR U12946 ( .A(n12171), .B(n12170), .Z(n12150) );
  XNOR U12947 ( .A(n12189), .B(n12188), .Z(n12194) );
  NAND U12948 ( .A(n11995), .B(n11994), .Z(n11999) );
  NANDN U12949 ( .A(n11997), .B(n11996), .Z(n11998) );
  NAND U12950 ( .A(n11999), .B(n11998), .Z(n12193) );
  NAND U12951 ( .A(n12001), .B(n12000), .Z(n12005) );
  NAND U12952 ( .A(n12003), .B(n12002), .Z(n12004) );
  NAND U12953 ( .A(n12005), .B(n12004), .Z(n12192) );
  XNOR U12954 ( .A(n12193), .B(n12192), .Z(n12195) );
  XNOR U12955 ( .A(n12041), .B(n12042), .Z(n12043) );
  NANDN U12956 ( .A(n12007), .B(n12006), .Z(n12011) );
  NAND U12957 ( .A(n12009), .B(n12008), .Z(n12010) );
  NAND U12958 ( .A(n12011), .B(n12010), .Z(n12049) );
  NAND U12959 ( .A(n12013), .B(n12012), .Z(n12017) );
  NAND U12960 ( .A(n12015), .B(n12014), .Z(n12016) );
  NAND U12961 ( .A(n12017), .B(n12016), .Z(n12047) );
  NAND U12962 ( .A(n12019), .B(n12018), .Z(n12023) );
  NANDN U12963 ( .A(n12021), .B(n12020), .Z(n12022) );
  AND U12964 ( .A(n12023), .B(n12022), .Z(n12048) );
  XNOR U12965 ( .A(n12047), .B(n12048), .Z(n12050) );
  XNOR U12966 ( .A(n12043), .B(n12044), .Z(n12036) );
  XNOR U12967 ( .A(n12037), .B(n12036), .Z(n12040) );
  NANDN U12968 ( .A(n12028), .B(n12027), .Z(n12032) );
  OR U12969 ( .A(n12030), .B(n12029), .Z(n12031) );
  NAND U12970 ( .A(n12032), .B(n12031), .Z(n12038) );
  XOR U12971 ( .A(n12039), .B(n12038), .Z(n12033) );
  XNOR U12972 ( .A(n12040), .B(n12033), .Z(N253) );
  NANDN U12973 ( .A(n12042), .B(n12041), .Z(n12046) );
  NANDN U12974 ( .A(n12044), .B(n12043), .Z(n12045) );
  NAND U12975 ( .A(n12046), .B(n12045), .Z(n12204) );
  NAND U12976 ( .A(n12048), .B(n12047), .Z(n12052) );
  NANDN U12977 ( .A(n12050), .B(n12049), .Z(n12051) );
  NAND U12978 ( .A(n12052), .B(n12051), .Z(n12203) );
  NAND U12979 ( .A(n12054), .B(n12053), .Z(n12058) );
  NAND U12980 ( .A(n12056), .B(n12055), .Z(n12057) );
  NAND U12981 ( .A(n12058), .B(n12057), .Z(n12220) );
  NAND U12982 ( .A(n12060), .B(n12059), .Z(n12064) );
  NAND U12983 ( .A(n12062), .B(n12061), .Z(n12063) );
  AND U12984 ( .A(n12064), .B(n12063), .Z(n12329) );
  NAND U12985 ( .A(n12066), .B(n12065), .Z(n12070) );
  NAND U12986 ( .A(n12068), .B(n12067), .Z(n12069) );
  NAND U12987 ( .A(n12070), .B(n12069), .Z(n12369) );
  NAND U12988 ( .A(n12072), .B(n12071), .Z(n12076) );
  NAND U12989 ( .A(n12074), .B(n12073), .Z(n12075) );
  NAND U12990 ( .A(n12076), .B(n12075), .Z(n12368) );
  XOR U12991 ( .A(n12369), .B(n12368), .Z(n12370) );
  AND U12992 ( .A(y[1908]), .B(x[234]), .Z(n12366) );
  NAND U12993 ( .A(n12077), .B(n12366), .Z(n12081) );
  NAND U12994 ( .A(n12079), .B(n12078), .Z(n12080) );
  NAND U12995 ( .A(n12081), .B(n12080), .Z(n12337) );
  AND U12996 ( .A(x[246]), .B(y[1895]), .Z(n12282) );
  AND U12997 ( .A(x[236]), .B(y[1905]), .Z(n12527) );
  AND U12998 ( .A(x[225]), .B(y[1916]), .Z(n12280) );
  XOR U12999 ( .A(n12527), .B(n12280), .Z(n12281) );
  XOR U13000 ( .A(n12282), .B(n12281), .Z(n12336) );
  AND U13001 ( .A(x[239]), .B(y[1902]), .Z(n12285) );
  XOR U13002 ( .A(n12336), .B(n12335), .Z(n12338) );
  XNOR U13003 ( .A(n12337), .B(n12338), .Z(n12371) );
  NAND U13004 ( .A(n12083), .B(n12082), .Z(n12087) );
  NAND U13005 ( .A(n12085), .B(n12084), .Z(n12086) );
  AND U13006 ( .A(n12087), .B(n12086), .Z(n12331) );
  XOR U13007 ( .A(n12332), .B(n12331), .Z(n12326) );
  NAND U13008 ( .A(n12089), .B(n12088), .Z(n12093) );
  NAND U13009 ( .A(n12091), .B(n12090), .Z(n12092) );
  NAND U13010 ( .A(n12093), .B(n12092), .Z(n12342) );
  AND U13011 ( .A(n12095), .B(n12094), .Z(n12099) );
  NAND U13012 ( .A(n12097), .B(n12096), .Z(n12098) );
  NANDN U13013 ( .A(n12099), .B(n12098), .Z(n12341) );
  XOR U13014 ( .A(n12342), .B(n12341), .Z(n12343) );
  NAND U13015 ( .A(n12101), .B(n12100), .Z(n12105) );
  NAND U13016 ( .A(n12103), .B(n12102), .Z(n12104) );
  NAND U13017 ( .A(n12105), .B(n12104), .Z(n12246) );
  AND U13018 ( .A(x[247]), .B(y[1894]), .Z(n12302) );
  AND U13019 ( .A(x[237]), .B(y[1904]), .Z(n12300) );
  AND U13020 ( .A(x[248]), .B(y[1893]), .Z(n12533) );
  XOR U13021 ( .A(n12300), .B(n12533), .Z(n12301) );
  XOR U13022 ( .A(n12302), .B(n12301), .Z(n12245) );
  AND U13023 ( .A(x[235]), .B(y[1906]), .Z(n12308) );
  AND U13024 ( .A(x[227]), .B(y[1914]), .Z(n12306) );
  AND U13025 ( .A(x[241]), .B(y[1900]), .Z(n12305) );
  XOR U13026 ( .A(n12306), .B(n12305), .Z(n12307) );
  XOR U13027 ( .A(n12308), .B(n12307), .Z(n12244) );
  XOR U13028 ( .A(n12245), .B(n12244), .Z(n12247) );
  XNOR U13029 ( .A(n12246), .B(n12247), .Z(n12344) );
  NAND U13030 ( .A(n12293), .B(n12106), .Z(n12110) );
  NAND U13031 ( .A(n12108), .B(n12107), .Z(n12109) );
  NAND U13032 ( .A(n12110), .B(n12109), .Z(n12350) );
  AND U13033 ( .A(x[249]), .B(y[1892]), .Z(n12277) );
  AND U13034 ( .A(x[250]), .B(y[1891]), .Z(n12274) );
  XOR U13035 ( .A(n12275), .B(n12274), .Z(n12276) );
  XOR U13036 ( .A(n12277), .B(n12276), .Z(n12348) );
  AND U13037 ( .A(x[252]), .B(y[1889]), .Z(n12292) );
  XOR U13038 ( .A(o[125]), .B(n12292), .Z(n12361) );
  AND U13039 ( .A(x[224]), .B(y[1917]), .Z(n12359) );
  AND U13040 ( .A(x[253]), .B(y[1888]), .Z(n12358) );
  XOR U13041 ( .A(n12359), .B(n12358), .Z(n12360) );
  XNOR U13042 ( .A(n12361), .B(n12360), .Z(n12347) );
  XOR U13043 ( .A(n12350), .B(n12349), .Z(n12232) );
  NAND U13044 ( .A(n12112), .B(n12111), .Z(n12116) );
  NAND U13045 ( .A(n12114), .B(n12113), .Z(n12115) );
  NAND U13046 ( .A(n12116), .B(n12115), .Z(n12313) );
  AND U13047 ( .A(n12117), .B(o[124]), .Z(n12253) );
  AND U13048 ( .A(x[240]), .B(y[1901]), .Z(n12251) );
  AND U13049 ( .A(x[251]), .B(y[1890]), .Z(n12250) );
  XOR U13050 ( .A(n12251), .B(n12250), .Z(n12252) );
  XOR U13051 ( .A(n12253), .B(n12252), .Z(n12312) );
  AND U13052 ( .A(x[226]), .B(y[1915]), .Z(n12262) );
  XOR U13053 ( .A(n12265), .B(n12264), .Z(n12311) );
  XOR U13054 ( .A(n12312), .B(n12311), .Z(n12314) );
  XOR U13055 ( .A(n12313), .B(n12314), .Z(n12233) );
  NANDN U13056 ( .A(n12119), .B(n12118), .Z(n12123) );
  NAND U13057 ( .A(n12121), .B(n12120), .Z(n12122) );
  NAND U13058 ( .A(n12123), .B(n12122), .Z(n12238) );
  NAND U13059 ( .A(n12125), .B(n12124), .Z(n12129) );
  NAND U13060 ( .A(n12127), .B(n12126), .Z(n12128) );
  NAND U13061 ( .A(n12129), .B(n12128), .Z(n12269) );
  NAND U13062 ( .A(n12131), .B(n12130), .Z(n12135) );
  NAND U13063 ( .A(n12133), .B(n12132), .Z(n12134) );
  NAND U13064 ( .A(n12135), .B(n12134), .Z(n12268) );
  XOR U13065 ( .A(n12269), .B(n12268), .Z(n12271) );
  AND U13066 ( .A(x[232]), .B(y[1909]), .Z(n12295) );
  AND U13067 ( .A(x[230]), .B(y[1911]), .Z(n12137) );
  AND U13068 ( .A(y[1910]), .B(x[231]), .Z(n12136) );
  XOR U13069 ( .A(n12137), .B(n12136), .Z(n12294) );
  XOR U13070 ( .A(n12295), .B(n12294), .Z(n12353) );
  AND U13071 ( .A(x[233]), .B(y[1908]), .Z(n12465) );
  XOR U13072 ( .A(n12353), .B(n12465), .Z(n12355) );
  AND U13073 ( .A(x[229]), .B(y[1912]), .Z(n12259) );
  AND U13074 ( .A(x[228]), .B(y[1913]), .Z(n12257) );
  AND U13075 ( .A(x[234]), .B(y[1907]), .Z(n12256) );
  XOR U13076 ( .A(n12257), .B(n12256), .Z(n12258) );
  XOR U13077 ( .A(n12259), .B(n12258), .Z(n12354) );
  XOR U13078 ( .A(n12355), .B(n12354), .Z(n12270) );
  XOR U13079 ( .A(n12271), .B(n12270), .Z(n12239) );
  XNOR U13080 ( .A(n12240), .B(n12241), .Z(n12324) );
  NAND U13081 ( .A(n12139), .B(n12138), .Z(n12143) );
  NAND U13082 ( .A(n12141), .B(n12140), .Z(n12142) );
  NAND U13083 ( .A(n12143), .B(n12142), .Z(n12323) );
  XOR U13084 ( .A(n12220), .B(n12221), .Z(n12223) );
  NAND U13085 ( .A(n12145), .B(n12144), .Z(n12149) );
  NAND U13086 ( .A(n12147), .B(n12146), .Z(n12148) );
  NAND U13087 ( .A(n12149), .B(n12148), .Z(n12214) );
  NANDN U13088 ( .A(n12151), .B(n12150), .Z(n12155) );
  NANDN U13089 ( .A(n12153), .B(n12152), .Z(n12154) );
  AND U13090 ( .A(n12155), .B(n12154), .Z(n12215) );
  XOR U13091 ( .A(n12214), .B(n12215), .Z(n12217) );
  NAND U13092 ( .A(n12157), .B(n12156), .Z(n12161) );
  NAND U13093 ( .A(n12159), .B(n12158), .Z(n12160) );
  NAND U13094 ( .A(n12161), .B(n12160), .Z(n12228) );
  NANDN U13095 ( .A(n12163), .B(n12162), .Z(n12167) );
  NAND U13096 ( .A(n12165), .B(n12164), .Z(n12166) );
  NAND U13097 ( .A(n12167), .B(n12166), .Z(n12226) );
  NAND U13098 ( .A(n12169), .B(n12168), .Z(n12173) );
  NAND U13099 ( .A(n12171), .B(n12170), .Z(n12172) );
  NAND U13100 ( .A(n12173), .B(n12172), .Z(n12319) );
  NAND U13101 ( .A(n12175), .B(n12174), .Z(n12179) );
  NAND U13102 ( .A(n12177), .B(n12176), .Z(n12178) );
  NAND U13103 ( .A(n12179), .B(n12178), .Z(n12318) );
  NAND U13104 ( .A(n12181), .B(n12180), .Z(n12185) );
  NAND U13105 ( .A(n12183), .B(n12182), .Z(n12184) );
  NAND U13106 ( .A(n12185), .B(n12184), .Z(n12317) );
  XOR U13107 ( .A(n12318), .B(n12317), .Z(n12320) );
  XOR U13108 ( .A(n12319), .B(n12320), .Z(n12227) );
  XOR U13109 ( .A(n12226), .B(n12227), .Z(n12229) );
  XOR U13110 ( .A(n12228), .B(n12229), .Z(n12216) );
  XOR U13111 ( .A(n12217), .B(n12216), .Z(n12222) );
  XNOR U13112 ( .A(n12223), .B(n12222), .Z(n12210) );
  NANDN U13113 ( .A(n12187), .B(n12186), .Z(n12191) );
  NAND U13114 ( .A(n12189), .B(n12188), .Z(n12190) );
  NAND U13115 ( .A(n12191), .B(n12190), .Z(n12208) );
  NAND U13116 ( .A(n12193), .B(n12192), .Z(n12197) );
  NANDN U13117 ( .A(n12195), .B(n12194), .Z(n12196) );
  AND U13118 ( .A(n12197), .B(n12196), .Z(n12209) );
  XNOR U13119 ( .A(n12208), .B(n12209), .Z(n12211) );
  XOR U13120 ( .A(n12210), .B(n12211), .Z(n12202) );
  XOR U13121 ( .A(n12203), .B(n12202), .Z(n12205) );
  XOR U13122 ( .A(n12204), .B(n12205), .Z(n12201) );
  XOR U13123 ( .A(n12199), .B(n12201), .Z(n12198) );
  XOR U13124 ( .A(n12200), .B(n12198), .Z(N254) );
  NAND U13125 ( .A(n12203), .B(n12202), .Z(n12207) );
  NAND U13126 ( .A(n12205), .B(n12204), .Z(n12206) );
  AND U13127 ( .A(n12207), .B(n12206), .Z(n12376) );
  XNOR U13128 ( .A(n12377), .B(n12376), .Z(n12375) );
  NAND U13129 ( .A(n12209), .B(n12208), .Z(n12213) );
  NANDN U13130 ( .A(n12211), .B(n12210), .Z(n12212) );
  AND U13131 ( .A(n12213), .B(n12212), .Z(n12661) );
  NAND U13132 ( .A(n12215), .B(n12214), .Z(n12219) );
  NAND U13133 ( .A(n12217), .B(n12216), .Z(n12218) );
  AND U13134 ( .A(n12219), .B(n12218), .Z(n12667) );
  NAND U13135 ( .A(n12221), .B(n12220), .Z(n12225) );
  NAND U13136 ( .A(n12223), .B(n12222), .Z(n12224) );
  AND U13137 ( .A(n12225), .B(n12224), .Z(n12666) );
  XOR U13138 ( .A(n12667), .B(n12666), .Z(n12669) );
  NAND U13139 ( .A(n12227), .B(n12226), .Z(n12231) );
  NAND U13140 ( .A(n12229), .B(n12228), .Z(n12230) );
  AND U13141 ( .A(n12231), .B(n12230), .Z(n12668) );
  XOR U13142 ( .A(n12669), .B(n12668), .Z(n12662) );
  NANDN U13143 ( .A(n12233), .B(n12232), .Z(n12237) );
  NANDN U13144 ( .A(n12235), .B(n12234), .Z(n12236) );
  AND U13145 ( .A(n12237), .B(n12236), .Z(n12648) );
  NANDN U13146 ( .A(n12239), .B(n12238), .Z(n12243) );
  NANDN U13147 ( .A(n12241), .B(n12240), .Z(n12242) );
  AND U13148 ( .A(n12243), .B(n12242), .Z(n12640) );
  NAND U13149 ( .A(n12245), .B(n12244), .Z(n12249) );
  NAND U13150 ( .A(n12247), .B(n12246), .Z(n12248) );
  AND U13151 ( .A(n12249), .B(n12248), .Z(n12624) );
  NAND U13152 ( .A(n12251), .B(n12250), .Z(n12255) );
  NAND U13153 ( .A(n12253), .B(n12252), .Z(n12254) );
  NAND U13154 ( .A(n12255), .B(n12254), .Z(n12582) );
  NAND U13155 ( .A(n12257), .B(n12256), .Z(n12261) );
  NAND U13156 ( .A(n12259), .B(n12258), .Z(n12260) );
  NAND U13157 ( .A(n12261), .B(n12260), .Z(n12585) );
  AND U13158 ( .A(x[230]), .B(y[1912]), .Z(n12545) );
  AND U13159 ( .A(x[229]), .B(y[1913]), .Z(n12547) );
  AND U13160 ( .A(x[243]), .B(y[1899]), .Z(n12546) );
  XOR U13161 ( .A(n12547), .B(n12546), .Z(n12544) );
  XNOR U13162 ( .A(n12545), .B(n12544), .Z(n12559) );
  AND U13163 ( .A(x[228]), .B(y[1914]), .Z(n12456) );
  AND U13164 ( .A(x[227]), .B(y[1915]), .Z(n12458) );
  AND U13165 ( .A(x[242]), .B(y[1900]), .Z(n12457) );
  XOR U13166 ( .A(n12458), .B(n12457), .Z(n12455) );
  XOR U13167 ( .A(n12456), .B(n12455), .Z(n12556) );
  NANDN U13168 ( .A(n12263), .B(n12262), .Z(n12267) );
  NAND U13169 ( .A(n12265), .B(n12264), .Z(n12266) );
  AND U13170 ( .A(n12267), .B(n12266), .Z(n12557) );
  XOR U13171 ( .A(n12559), .B(n12558), .Z(n12584) );
  XOR U13172 ( .A(n12585), .B(n12584), .Z(n12583) );
  XOR U13173 ( .A(n12582), .B(n12583), .Z(n12625) );
  NAND U13174 ( .A(n12269), .B(n12268), .Z(n12273) );
  NAND U13175 ( .A(n12271), .B(n12270), .Z(n12272) );
  AND U13176 ( .A(n12273), .B(n12272), .Z(n12622) );
  XOR U13177 ( .A(n12623), .B(n12622), .Z(n12643) );
  AND U13178 ( .A(n12275), .B(n12274), .Z(n12279) );
  NAND U13179 ( .A(n12277), .B(n12276), .Z(n12278) );
  NANDN U13180 ( .A(n12279), .B(n12278), .Z(n12576) );
  AND U13181 ( .A(n12527), .B(n12280), .Z(n12284) );
  NAND U13182 ( .A(n12282), .B(n12281), .Z(n12283) );
  NANDN U13183 ( .A(n12284), .B(n12283), .Z(n12579) );
  NANDN U13184 ( .A(n12452), .B(n12285), .Z(n12289) );
  NANDN U13185 ( .A(n12287), .B(n12286), .Z(n12288) );
  AND U13186 ( .A(n12289), .B(n12288), .Z(n12571) );
  AND U13187 ( .A(x[247]), .B(y[1895]), .Z(n12531) );
  AND U13188 ( .A(y[1894]), .B(x[248]), .Z(n12291) );
  AND U13189 ( .A(y[1893]), .B(x[249]), .Z(n12290) );
  XOR U13190 ( .A(n12291), .B(n12290), .Z(n12530) );
  XOR U13191 ( .A(n12531), .B(n12530), .Z(n12569) );
  AND U13192 ( .A(n12292), .B(o[125]), .Z(n12539) );
  AND U13193 ( .A(x[252]), .B(y[1890]), .Z(n12541) );
  AND U13194 ( .A(x[240]), .B(y[1902]), .Z(n12540) );
  XOR U13195 ( .A(n12541), .B(n12540), .Z(n12538) );
  XNOR U13196 ( .A(n12539), .B(n12538), .Z(n12568) );
  XNOR U13197 ( .A(n12571), .B(n12570), .Z(n12578) );
  XOR U13198 ( .A(n12579), .B(n12578), .Z(n12577) );
  XOR U13199 ( .A(n12576), .B(n12577), .Z(n12617) );
  AND U13200 ( .A(x[231]), .B(y[1911]), .Z(n12451) );
  NAND U13201 ( .A(n12293), .B(n12451), .Z(n12297) );
  NAND U13202 ( .A(n12295), .B(n12294), .Z(n12296) );
  AND U13203 ( .A(n12297), .B(n12296), .Z(n12395) );
  AND U13204 ( .A(y[1897]), .B(x[245]), .Z(n12299) );
  AND U13205 ( .A(y[1896]), .B(x[246]), .Z(n12298) );
  XOR U13206 ( .A(n12299), .B(n12298), .Z(n12450) );
  XOR U13207 ( .A(n12451), .B(n12450), .Z(n12393) );
  AND U13208 ( .A(x[241]), .B(y[1901]), .Z(n12419) );
  AND U13209 ( .A(x[226]), .B(y[1916]), .Z(n12421) );
  AND U13210 ( .A(x[250]), .B(y[1892]), .Z(n12420) );
  XOR U13211 ( .A(n12421), .B(n12420), .Z(n12418) );
  XNOR U13212 ( .A(n12419), .B(n12418), .Z(n12392) );
  XNOR U13213 ( .A(n12395), .B(n12394), .Z(n12387) );
  NAND U13214 ( .A(n12300), .B(n12533), .Z(n12304) );
  NAND U13215 ( .A(n12302), .B(n12301), .Z(n12303) );
  NAND U13216 ( .A(n12304), .B(n12303), .Z(n12389) );
  NAND U13217 ( .A(n12306), .B(n12305), .Z(n12310) );
  NAND U13218 ( .A(n12308), .B(n12307), .Z(n12309) );
  AND U13219 ( .A(n12310), .B(n12309), .Z(n12401) );
  AND U13220 ( .A(x[224]), .B(y[1918]), .Z(n12445) );
  AND U13221 ( .A(x[253]), .B(y[1889]), .Z(n12468) );
  XOR U13222 ( .A(o[126]), .B(n12468), .Z(n12447) );
  AND U13223 ( .A(x[254]), .B(y[1888]), .Z(n12446) );
  XOR U13224 ( .A(n12447), .B(n12446), .Z(n12444) );
  XOR U13225 ( .A(n12445), .B(n12444), .Z(n12399) );
  AND U13226 ( .A(x[244]), .B(y[1898]), .Z(n12414) );
  XOR U13227 ( .A(n12415), .B(n12414), .Z(n12413) );
  AND U13228 ( .A(x[232]), .B(y[1910]), .Z(n12412) );
  XNOR U13229 ( .A(n12413), .B(n12412), .Z(n12398) );
  XNOR U13230 ( .A(n12401), .B(n12400), .Z(n12388) );
  XOR U13231 ( .A(n12389), .B(n12388), .Z(n12386) );
  NAND U13232 ( .A(n12312), .B(n12311), .Z(n12316) );
  NAND U13233 ( .A(n12314), .B(n12313), .Z(n12315) );
  NAND U13234 ( .A(n12316), .B(n12315), .Z(n12618) );
  XOR U13235 ( .A(n12619), .B(n12618), .Z(n12616) );
  XOR U13236 ( .A(n12617), .B(n12616), .Z(n12642) );
  XNOR U13237 ( .A(n12640), .B(n12641), .Z(n12650) );
  NAND U13238 ( .A(n12318), .B(n12317), .Z(n12322) );
  NAND U13239 ( .A(n12320), .B(n12319), .Z(n12321) );
  AND U13240 ( .A(n12322), .B(n12321), .Z(n12649) );
  NANDN U13241 ( .A(n12324), .B(n12323), .Z(n12328) );
  NANDN U13242 ( .A(n12326), .B(n12325), .Z(n12327) );
  NAND U13243 ( .A(n12328), .B(n12327), .Z(n12636) );
  NANDN U13244 ( .A(n12330), .B(n12329), .Z(n12334) );
  NAND U13245 ( .A(n12332), .B(n12331), .Z(n12333) );
  AND U13246 ( .A(n12334), .B(n12333), .Z(n12381) );
  NAND U13247 ( .A(n12336), .B(n12335), .Z(n12340) );
  NAND U13248 ( .A(n12338), .B(n12337), .Z(n12339) );
  AND U13249 ( .A(n12340), .B(n12339), .Z(n12607) );
  NAND U13250 ( .A(n12342), .B(n12341), .Z(n12346) );
  NANDN U13251 ( .A(n12344), .B(n12343), .Z(n12345) );
  AND U13252 ( .A(n12346), .B(n12345), .Z(n12606) );
  XOR U13253 ( .A(n12607), .B(n12606), .Z(n12605) );
  NANDN U13254 ( .A(n12348), .B(n12347), .Z(n12352) );
  OR U13255 ( .A(n12350), .B(n12349), .Z(n12351) );
  NAND U13256 ( .A(n12352), .B(n12351), .Z(n12604) );
  XOR U13257 ( .A(n12605), .B(n12604), .Z(n12383) );
  NAND U13258 ( .A(n12353), .B(n12465), .Z(n12357) );
  NAND U13259 ( .A(n12355), .B(n12354), .Z(n12356) );
  AND U13260 ( .A(n12357), .B(n12356), .Z(n12600) );
  NAND U13261 ( .A(n12359), .B(n12358), .Z(n12363) );
  NAND U13262 ( .A(n12361), .B(n12360), .Z(n12362) );
  NAND U13263 ( .A(n12363), .B(n12362), .Z(n12564) );
  AND U13264 ( .A(y[1906]), .B(x[236]), .Z(n12364) );
  XOR U13265 ( .A(n12365), .B(n12364), .Z(n12524) );
  XOR U13266 ( .A(n12525), .B(n12524), .Z(n12464) );
  AND U13267 ( .A(y[1909]), .B(x[233]), .Z(n12367) );
  XOR U13268 ( .A(n12367), .B(n12366), .Z(n12463) );
  XOR U13269 ( .A(n12464), .B(n12463), .Z(n12563) );
  AND U13270 ( .A(x[251]), .B(y[1891]), .Z(n12409) );
  AND U13271 ( .A(x[225]), .B(y[1917]), .Z(n12408) );
  XOR U13272 ( .A(n12409), .B(n12408), .Z(n12406) );
  XOR U13273 ( .A(n12407), .B(n12406), .Z(n12562) );
  XOR U13274 ( .A(n12563), .B(n12562), .Z(n12565) );
  XOR U13275 ( .A(n12564), .B(n12565), .Z(n12601) );
  NAND U13276 ( .A(n12369), .B(n12368), .Z(n12373) );
  NANDN U13277 ( .A(n12371), .B(n12370), .Z(n12372) );
  AND U13278 ( .A(n12373), .B(n12372), .Z(n12598) );
  XNOR U13279 ( .A(n12599), .B(n12598), .Z(n12382) );
  XOR U13280 ( .A(n12381), .B(n12380), .Z(n12637) );
  XNOR U13281 ( .A(n12636), .B(n12637), .Z(n12635) );
  XNOR U13282 ( .A(n12661), .B(n12660), .Z(n12374) );
  XNOR U13283 ( .A(n12375), .B(n12374), .Z(N255) );
  NAND U13284 ( .A(n12375), .B(n12374), .Z(n12379) );
  NANDN U13285 ( .A(n12377), .B(n12376), .Z(n12378) );
  AND U13286 ( .A(n12379), .B(n12378), .Z(n12659) );
  NAND U13287 ( .A(n12381), .B(n12380), .Z(n12385) );
  NANDN U13288 ( .A(n12383), .B(n12382), .Z(n12384) );
  AND U13289 ( .A(n12385), .B(n12384), .Z(n12633) );
  NANDN U13290 ( .A(n12387), .B(n12386), .Z(n12391) );
  NAND U13291 ( .A(n12389), .B(n12388), .Z(n12390) );
  AND U13292 ( .A(n12391), .B(n12390), .Z(n12615) );
  NANDN U13293 ( .A(n12393), .B(n12392), .Z(n12397) );
  ANDN U13294 ( .B(n12395), .A(n12394), .Z(n12396) );
  ANDN U13295 ( .B(n12397), .A(n12396), .Z(n12405) );
  NANDN U13296 ( .A(n12399), .B(n12398), .Z(n12403) );
  AND U13297 ( .A(n12401), .B(n12400), .Z(n12402) );
  ANDN U13298 ( .B(n12403), .A(n12402), .Z(n12404) );
  XNOR U13299 ( .A(n12405), .B(n12404), .Z(n12597) );
  NAND U13300 ( .A(n12407), .B(n12406), .Z(n12411) );
  NAND U13301 ( .A(n12409), .B(n12408), .Z(n12410) );
  AND U13302 ( .A(n12411), .B(n12410), .Z(n12443) );
  NAND U13303 ( .A(n12413), .B(n12412), .Z(n12417) );
  NAND U13304 ( .A(n12415), .B(n12414), .Z(n12416) );
  AND U13305 ( .A(n12417), .B(n12416), .Z(n12425) );
  NAND U13306 ( .A(n12419), .B(n12418), .Z(n12423) );
  NAND U13307 ( .A(n12421), .B(n12420), .Z(n12422) );
  NAND U13308 ( .A(n12423), .B(n12422), .Z(n12424) );
  XNOR U13309 ( .A(n12425), .B(n12424), .Z(n12441) );
  AND U13310 ( .A(y[1892]), .B(x[251]), .Z(n12427) );
  NAND U13311 ( .A(y[1901]), .B(x[242]), .Z(n12426) );
  XNOR U13312 ( .A(n12427), .B(n12426), .Z(n12431) );
  AND U13313 ( .A(y[1900]), .B(x[243]), .Z(n12429) );
  NAND U13314 ( .A(y[1898]), .B(x[245]), .Z(n12428) );
  XNOR U13315 ( .A(n12429), .B(n12428), .Z(n12430) );
  XOR U13316 ( .A(n12431), .B(n12430), .Z(n12439) );
  AND U13317 ( .A(y[1916]), .B(x[227]), .Z(n12433) );
  NAND U13318 ( .A(y[1915]), .B(x[228]), .Z(n12432) );
  XNOR U13319 ( .A(n12433), .B(n12432), .Z(n12437) );
  AND U13320 ( .A(y[1888]), .B(x[255]), .Z(n12435) );
  NAND U13321 ( .A(y[1912]), .B(x[231]), .Z(n12434) );
  XNOR U13322 ( .A(n12435), .B(n12434), .Z(n12436) );
  XNOR U13323 ( .A(n12437), .B(n12436), .Z(n12438) );
  XNOR U13324 ( .A(n12439), .B(n12438), .Z(n12440) );
  XNOR U13325 ( .A(n12441), .B(n12440), .Z(n12442) );
  XNOR U13326 ( .A(n12443), .B(n12442), .Z(n12523) );
  NAND U13327 ( .A(n12445), .B(n12444), .Z(n12449) );
  NAND U13328 ( .A(n12447), .B(n12446), .Z(n12448) );
  AND U13329 ( .A(n12449), .B(n12448), .Z(n12521) );
  NAND U13330 ( .A(n12451), .B(n12450), .Z(n12454) );
  AND U13331 ( .A(x[246]), .B(y[1897]), .Z(n12469) );
  NANDN U13332 ( .A(n12452), .B(n12469), .Z(n12453) );
  AND U13333 ( .A(n12454), .B(n12453), .Z(n12462) );
  NAND U13334 ( .A(n12456), .B(n12455), .Z(n12460) );
  NAND U13335 ( .A(n12458), .B(n12457), .Z(n12459) );
  NAND U13336 ( .A(n12460), .B(n12459), .Z(n12461) );
  XNOR U13337 ( .A(n12462), .B(n12461), .Z(n12519) );
  NAND U13338 ( .A(n12464), .B(n12463), .Z(n12467) );
  AND U13339 ( .A(x[234]), .B(y[1909]), .Z(n12491) );
  NAND U13340 ( .A(n12465), .B(n12491), .Z(n12466) );
  AND U13341 ( .A(n12467), .B(n12466), .Z(n12517) );
  AND U13342 ( .A(y[1917]), .B(x[226]), .Z(n12476) );
  AND U13343 ( .A(n12468), .B(o[126]), .Z(n12474) );
  XOR U13344 ( .A(n12469), .B(o[127]), .Z(n12472) );
  AND U13345 ( .A(x[249]), .B(y[1894]), .Z(n12532) );
  XNOR U13346 ( .A(n12470), .B(n12532), .Z(n12471) );
  XNOR U13347 ( .A(n12472), .B(n12471), .Z(n12473) );
  XNOR U13348 ( .A(n12474), .B(n12473), .Z(n12475) );
  XNOR U13349 ( .A(n12476), .B(n12475), .Z(n12515) );
  AND U13350 ( .A(y[1891]), .B(x[252]), .Z(n12482) );
  AND U13351 ( .A(y[1899]), .B(x[244]), .Z(n12478) );
  NAND U13352 ( .A(y[1911]), .B(x[232]), .Z(n12477) );
  XNOR U13353 ( .A(n12478), .B(n12477), .Z(n12479) );
  XNOR U13354 ( .A(n12480), .B(n12479), .Z(n12481) );
  XNOR U13355 ( .A(n12482), .B(n12481), .Z(n12505) );
  AND U13356 ( .A(y[1889]), .B(x[254]), .Z(n12484) );
  NAND U13357 ( .A(y[1890]), .B(x[253]), .Z(n12483) );
  XNOR U13358 ( .A(n12484), .B(n12483), .Z(n12495) );
  AND U13359 ( .A(y[1908]), .B(x[235]), .Z(n12486) );
  NAND U13360 ( .A(y[1910]), .B(x[233]), .Z(n12485) );
  XNOR U13361 ( .A(n12486), .B(n12485), .Z(n12490) );
  AND U13362 ( .A(y[1907]), .B(x[236]), .Z(n12488) );
  NAND U13363 ( .A(y[1893]), .B(x[250]), .Z(n12487) );
  XNOR U13364 ( .A(n12488), .B(n12487), .Z(n12489) );
  XOR U13365 ( .A(n12490), .B(n12489), .Z(n12493) );
  XNOR U13366 ( .A(n12526), .B(n12491), .Z(n12492) );
  XNOR U13367 ( .A(n12493), .B(n12492), .Z(n12494) );
  XOR U13368 ( .A(n12495), .B(n12494), .Z(n12503) );
  AND U13369 ( .A(y[1896]), .B(x[247]), .Z(n12497) );
  NAND U13370 ( .A(y[1902]), .B(x[241]), .Z(n12496) );
  XNOR U13371 ( .A(n12497), .B(n12496), .Z(n12501) );
  AND U13372 ( .A(y[1914]), .B(x[229]), .Z(n12499) );
  NAND U13373 ( .A(y[1913]), .B(x[230]), .Z(n12498) );
  XNOR U13374 ( .A(n12499), .B(n12498), .Z(n12500) );
  XNOR U13375 ( .A(n12501), .B(n12500), .Z(n12502) );
  XNOR U13376 ( .A(n12503), .B(n12502), .Z(n12504) );
  XOR U13377 ( .A(n12505), .B(n12504), .Z(n12513) );
  AND U13378 ( .A(y[1918]), .B(x[225]), .Z(n12507) );
  NAND U13379 ( .A(y[1919]), .B(x[224]), .Z(n12506) );
  XNOR U13380 ( .A(n12507), .B(n12506), .Z(n12511) );
  AND U13381 ( .A(y[1903]), .B(x[240]), .Z(n12509) );
  NAND U13382 ( .A(y[1905]), .B(x[238]), .Z(n12508) );
  XNOR U13383 ( .A(n12509), .B(n12508), .Z(n12510) );
  XNOR U13384 ( .A(n12511), .B(n12510), .Z(n12512) );
  XNOR U13385 ( .A(n12513), .B(n12512), .Z(n12514) );
  XNOR U13386 ( .A(n12515), .B(n12514), .Z(n12516) );
  XNOR U13387 ( .A(n12517), .B(n12516), .Z(n12518) );
  XNOR U13388 ( .A(n12519), .B(n12518), .Z(n12520) );
  XNOR U13389 ( .A(n12521), .B(n12520), .Z(n12522) );
  XOR U13390 ( .A(n12523), .B(n12522), .Z(n12555) );
  NAND U13391 ( .A(n12525), .B(n12524), .Z(n12529) );
  NAND U13392 ( .A(n12527), .B(n12526), .Z(n12528) );
  AND U13393 ( .A(n12529), .B(n12528), .Z(n12537) );
  NAND U13394 ( .A(n12531), .B(n12530), .Z(n12535) );
  NAND U13395 ( .A(n12533), .B(n12532), .Z(n12534) );
  NAND U13396 ( .A(n12535), .B(n12534), .Z(n12536) );
  XNOR U13397 ( .A(n12537), .B(n12536), .Z(n12553) );
  NAND U13398 ( .A(n12539), .B(n12538), .Z(n12543) );
  NAND U13399 ( .A(n12541), .B(n12540), .Z(n12542) );
  AND U13400 ( .A(n12543), .B(n12542), .Z(n12551) );
  NAND U13401 ( .A(n12545), .B(n12544), .Z(n12549) );
  NAND U13402 ( .A(n12547), .B(n12546), .Z(n12548) );
  NAND U13403 ( .A(n12549), .B(n12548), .Z(n12550) );
  XNOR U13404 ( .A(n12551), .B(n12550), .Z(n12552) );
  XNOR U13405 ( .A(n12553), .B(n12552), .Z(n12554) );
  XNOR U13406 ( .A(n12555), .B(n12554), .Z(n12595) );
  ANDN U13407 ( .B(n12557), .A(n12556), .Z(n12561) );
  ANDN U13408 ( .B(n12559), .A(n12558), .Z(n12560) );
  NOR U13409 ( .A(n12561), .B(n12560), .Z(n12593) );
  AND U13410 ( .A(n12563), .B(n12562), .Z(n12567) );
  AND U13411 ( .A(n12565), .B(n12564), .Z(n12566) );
  NOR U13412 ( .A(n12567), .B(n12566), .Z(n12575) );
  NANDN U13413 ( .A(n12569), .B(n12568), .Z(n12573) );
  NAND U13414 ( .A(n12571), .B(n12570), .Z(n12572) );
  AND U13415 ( .A(n12573), .B(n12572), .Z(n12574) );
  XNOR U13416 ( .A(n12575), .B(n12574), .Z(n12591) );
  NAND U13417 ( .A(n12577), .B(n12576), .Z(n12581) );
  NAND U13418 ( .A(n12579), .B(n12578), .Z(n12580) );
  AND U13419 ( .A(n12581), .B(n12580), .Z(n12589) );
  NAND U13420 ( .A(n12583), .B(n12582), .Z(n12587) );
  NAND U13421 ( .A(n12585), .B(n12584), .Z(n12586) );
  NAND U13422 ( .A(n12587), .B(n12586), .Z(n12588) );
  XNOR U13423 ( .A(n12589), .B(n12588), .Z(n12590) );
  XOR U13424 ( .A(n12591), .B(n12590), .Z(n12592) );
  XNOR U13425 ( .A(n12593), .B(n12592), .Z(n12594) );
  XOR U13426 ( .A(n12595), .B(n12594), .Z(n12596) );
  XNOR U13427 ( .A(n12597), .B(n12596), .Z(n12613) );
  NAND U13428 ( .A(n12599), .B(n12598), .Z(n12603) );
  NANDN U13429 ( .A(n12601), .B(n12600), .Z(n12602) );
  AND U13430 ( .A(n12603), .B(n12602), .Z(n12611) );
  NAND U13431 ( .A(n12605), .B(n12604), .Z(n12609) );
  NAND U13432 ( .A(n12607), .B(n12606), .Z(n12608) );
  NAND U13433 ( .A(n12609), .B(n12608), .Z(n12610) );
  XNOR U13434 ( .A(n12611), .B(n12610), .Z(n12612) );
  XNOR U13435 ( .A(n12613), .B(n12612), .Z(n12614) );
  XNOR U13436 ( .A(n12615), .B(n12614), .Z(n12631) );
  NAND U13437 ( .A(n12617), .B(n12616), .Z(n12621) );
  NAND U13438 ( .A(n12619), .B(n12618), .Z(n12620) );
  AND U13439 ( .A(n12621), .B(n12620), .Z(n12629) );
  NAND U13440 ( .A(n12623), .B(n12622), .Z(n12627) );
  NANDN U13441 ( .A(n12625), .B(n12624), .Z(n12626) );
  NAND U13442 ( .A(n12627), .B(n12626), .Z(n12628) );
  XNOR U13443 ( .A(n12629), .B(n12628), .Z(n12630) );
  XNOR U13444 ( .A(n12631), .B(n12630), .Z(n12632) );
  XNOR U13445 ( .A(n12633), .B(n12632), .Z(n12657) );
  NANDN U13446 ( .A(n12635), .B(n12634), .Z(n12639) );
  NAND U13447 ( .A(n12637), .B(n12636), .Z(n12638) );
  AND U13448 ( .A(n12639), .B(n12638), .Z(n12647) );
  NANDN U13449 ( .A(n12641), .B(n12640), .Z(n12645) );
  NANDN U13450 ( .A(n12643), .B(n12642), .Z(n12644) );
  NAND U13451 ( .A(n12645), .B(n12644), .Z(n12646) );
  XNOR U13452 ( .A(n12647), .B(n12646), .Z(n12655) );
  ANDN U13453 ( .B(n12649), .A(n12648), .Z(n12651) );
  NANDN U13454 ( .A(n12651), .B(n12650), .Z(n12652) );
  NAND U13455 ( .A(n12653), .B(n12652), .Z(n12654) );
  XNOR U13456 ( .A(n12655), .B(n12654), .Z(n12656) );
  XNOR U13457 ( .A(n12657), .B(n12656), .Z(n12658) );
  XNOR U13458 ( .A(n12659), .B(n12658), .Z(n12675) );
  NAND U13459 ( .A(n12661), .B(n12660), .Z(n12665) );
  ANDN U13460 ( .B(n12663), .A(n12662), .Z(n12664) );
  ANDN U13461 ( .B(n12665), .A(n12664), .Z(n12673) );
  AND U13462 ( .A(n12667), .B(n12666), .Z(n12671) );
  AND U13463 ( .A(n12669), .B(n12668), .Z(n12670) );
  OR U13464 ( .A(n12671), .B(n12670), .Z(n12672) );
  XNOR U13465 ( .A(n12673), .B(n12672), .Z(n12674) );
  XNOR U13466 ( .A(n12675), .B(n12674), .Z(N256) );
  AND U13467 ( .A(x[224]), .B(y[1920]), .Z(n13329) );
  XOR U13468 ( .A(n13329), .B(o[128]), .Z(N289) );
  AND U13469 ( .A(x[225]), .B(y[1920]), .Z(n12684) );
  AND U13470 ( .A(x[224]), .B(y[1921]), .Z(n12683) );
  XNOR U13471 ( .A(n12683), .B(o[129]), .Z(n12676) );
  XNOR U13472 ( .A(n12684), .B(n12676), .Z(n12678) );
  NAND U13473 ( .A(n13329), .B(o[128]), .Z(n12677) );
  XNOR U13474 ( .A(n12678), .B(n12677), .Z(N290) );
  NANDN U13475 ( .A(n12684), .B(n12676), .Z(n12680) );
  NAND U13476 ( .A(n12678), .B(n12677), .Z(n12679) );
  AND U13477 ( .A(n12680), .B(n12679), .Z(n12690) );
  AND U13478 ( .A(x[224]), .B(y[1922]), .Z(n12697) );
  XNOR U13479 ( .A(n12697), .B(o[130]), .Z(n12689) );
  XNOR U13480 ( .A(n12690), .B(n12689), .Z(n12692) );
  AND U13481 ( .A(y[1920]), .B(x[226]), .Z(n12682) );
  NAND U13482 ( .A(y[1921]), .B(x[225]), .Z(n12681) );
  XNOR U13483 ( .A(n12682), .B(n12681), .Z(n12686) );
  AND U13484 ( .A(n12683), .B(o[129]), .Z(n12685) );
  XNOR U13485 ( .A(n12686), .B(n12685), .Z(n12691) );
  XNOR U13486 ( .A(n12692), .B(n12691), .Z(N291) );
  AND U13487 ( .A(x[226]), .B(y[1921]), .Z(n12704) );
  NAND U13488 ( .A(n12704), .B(n12684), .Z(n12688) );
  NAND U13489 ( .A(n12686), .B(n12685), .Z(n12687) );
  AND U13490 ( .A(n12688), .B(n12687), .Z(n12707) );
  NANDN U13491 ( .A(n12690), .B(n12689), .Z(n12694) );
  NAND U13492 ( .A(n12692), .B(n12691), .Z(n12693) );
  AND U13493 ( .A(n12694), .B(n12693), .Z(n12706) );
  XNOR U13494 ( .A(n12707), .B(n12706), .Z(n12709) );
  AND U13495 ( .A(x[225]), .B(y[1922]), .Z(n12822) );
  XOR U13496 ( .A(n12704), .B(o[131]), .Z(n12712) );
  XOR U13497 ( .A(n12822), .B(n12712), .Z(n12714) );
  AND U13498 ( .A(y[1920]), .B(x[227]), .Z(n12696) );
  NAND U13499 ( .A(y[1923]), .B(x[224]), .Z(n12695) );
  XNOR U13500 ( .A(n12696), .B(n12695), .Z(n12699) );
  AND U13501 ( .A(n12697), .B(o[130]), .Z(n12698) );
  XOR U13502 ( .A(n12699), .B(n12698), .Z(n12713) );
  XOR U13503 ( .A(n12714), .B(n12713), .Z(n12708) );
  XOR U13504 ( .A(n12709), .B(n12708), .Z(N292) );
  AND U13505 ( .A(x[227]), .B(y[1923]), .Z(n12757) );
  NAND U13506 ( .A(n13329), .B(n12757), .Z(n12701) );
  NAND U13507 ( .A(n12699), .B(n12698), .Z(n12700) );
  NAND U13508 ( .A(n12701), .B(n12700), .Z(n12735) );
  AND U13509 ( .A(y[1924]), .B(x[224]), .Z(n12703) );
  NAND U13510 ( .A(y[1920]), .B(x[228]), .Z(n12702) );
  XNOR U13511 ( .A(n12703), .B(n12702), .Z(n12728) );
  AND U13512 ( .A(n12704), .B(o[131]), .Z(n12729) );
  XOR U13513 ( .A(n12728), .B(n12729), .Z(n12733) );
  AND U13514 ( .A(y[1922]), .B(x[226]), .Z(n12858) );
  NAND U13515 ( .A(y[1923]), .B(x[225]), .Z(n12705) );
  XNOR U13516 ( .A(n12858), .B(n12705), .Z(n12725) );
  AND U13517 ( .A(x[227]), .B(y[1921]), .Z(n12720) );
  XOR U13518 ( .A(o[132]), .B(n12720), .Z(n12724) );
  XOR U13519 ( .A(n12725), .B(n12724), .Z(n12732) );
  XOR U13520 ( .A(n12733), .B(n12732), .Z(n12734) );
  XOR U13521 ( .A(n12735), .B(n12734), .Z(n12739) );
  NANDN U13522 ( .A(n12707), .B(n12706), .Z(n12711) );
  NAND U13523 ( .A(n12709), .B(n12708), .Z(n12710) );
  NAND U13524 ( .A(n12711), .B(n12710), .Z(n12740) );
  NAND U13525 ( .A(n12822), .B(n12712), .Z(n12716) );
  NAND U13526 ( .A(n12714), .B(n12713), .Z(n12715) );
  NAND U13527 ( .A(n12716), .B(n12715), .Z(n12741) );
  IV U13528 ( .A(n12741), .Z(n12738) );
  XOR U13529 ( .A(n12740), .B(n12738), .Z(n12717) );
  XNOR U13530 ( .A(n12739), .B(n12717), .Z(N293) );
  AND U13531 ( .A(y[1922]), .B(x[227]), .Z(n12719) );
  NAND U13532 ( .A(y[1924]), .B(x[225]), .Z(n12718) );
  XNOR U13533 ( .A(n12719), .B(n12718), .Z(n12744) );
  AND U13534 ( .A(x[228]), .B(y[1921]), .Z(n12755) );
  XOR U13535 ( .A(n12755), .B(o[133]), .Z(n12743) );
  XNOR U13536 ( .A(n12744), .B(n12743), .Z(n12747) );
  AND U13537 ( .A(x[226]), .B(y[1923]), .Z(n12831) );
  AND U13538 ( .A(o[132]), .B(n12720), .Z(n12749) );
  AND U13539 ( .A(y[1920]), .B(x[229]), .Z(n12722) );
  NAND U13540 ( .A(y[1925]), .B(x[224]), .Z(n12721) );
  XNOR U13541 ( .A(n12722), .B(n12721), .Z(n12750) );
  XOR U13542 ( .A(n12749), .B(n12750), .Z(n12748) );
  XNOR U13543 ( .A(n12831), .B(n12748), .Z(n12723) );
  XOR U13544 ( .A(n12747), .B(n12723), .Z(n12765) );
  NAND U13545 ( .A(n12831), .B(n12822), .Z(n12727) );
  NAND U13546 ( .A(n12725), .B(n12724), .Z(n12726) );
  NAND U13547 ( .A(n12727), .B(n12726), .Z(n12763) );
  AND U13548 ( .A(x[228]), .B(y[1924]), .Z(n13545) );
  NAND U13549 ( .A(n13545), .B(n13329), .Z(n12731) );
  NAND U13550 ( .A(n12729), .B(n12728), .Z(n12730) );
  NAND U13551 ( .A(n12731), .B(n12730), .Z(n12762) );
  XOR U13552 ( .A(n12763), .B(n12762), .Z(n12764) );
  XNOR U13553 ( .A(n12765), .B(n12764), .Z(n12761) );
  NAND U13554 ( .A(n12733), .B(n12732), .Z(n12737) );
  NAND U13555 ( .A(n12735), .B(n12734), .Z(n12736) );
  NAND U13556 ( .A(n12737), .B(n12736), .Z(n12760) );
  XOR U13557 ( .A(n12760), .B(n12759), .Z(n12742) );
  XNOR U13558 ( .A(n12761), .B(n12742), .Z(N294) );
  AND U13559 ( .A(x[227]), .B(y[1924]), .Z(n12832) );
  NAND U13560 ( .A(n12832), .B(n12822), .Z(n12746) );
  NAND U13561 ( .A(n12744), .B(n12743), .Z(n12745) );
  NAND U13562 ( .A(n12746), .B(n12745), .Z(n12800) );
  XOR U13563 ( .A(n12800), .B(n12801), .Z(n12803) );
  AND U13564 ( .A(x[229]), .B(y[1925]), .Z(n13000) );
  NAND U13565 ( .A(n13329), .B(n13000), .Z(n12752) );
  NAND U13566 ( .A(n12750), .B(n12749), .Z(n12751) );
  NAND U13567 ( .A(n12752), .B(n12751), .Z(n12770) );
  AND U13568 ( .A(y[1920]), .B(x[230]), .Z(n12754) );
  NAND U13569 ( .A(y[1926]), .B(x[224]), .Z(n12753) );
  XNOR U13570 ( .A(n12754), .B(n12753), .Z(n12776) );
  AND U13571 ( .A(n12755), .B(o[133]), .Z(n12777) );
  XOR U13572 ( .A(n12776), .B(n12777), .Z(n12769) );
  XOR U13573 ( .A(n12770), .B(n12769), .Z(n12772) );
  NAND U13574 ( .A(y[1924]), .B(x[226]), .Z(n12756) );
  XNOR U13575 ( .A(n12757), .B(n12756), .Z(n12781) );
  AND U13576 ( .A(x[225]), .B(y[1925]), .Z(n13021) );
  NAND U13577 ( .A(y[1922]), .B(x[228]), .Z(n12758) );
  XNOR U13578 ( .A(n13021), .B(n12758), .Z(n12785) );
  AND U13579 ( .A(x[229]), .B(y[1921]), .Z(n12792) );
  XOR U13580 ( .A(o[134]), .B(n12792), .Z(n12784) );
  XOR U13581 ( .A(n12785), .B(n12784), .Z(n12780) );
  XOR U13582 ( .A(n12781), .B(n12780), .Z(n12771) );
  XOR U13583 ( .A(n12772), .B(n12771), .Z(n12802) );
  XOR U13584 ( .A(n12803), .B(n12802), .Z(n12796) );
  NAND U13585 ( .A(n12763), .B(n12762), .Z(n12767) );
  NAND U13586 ( .A(n12765), .B(n12764), .Z(n12766) );
  AND U13587 ( .A(n12767), .B(n12766), .Z(n12795) );
  IV U13588 ( .A(n12795), .Z(n12793) );
  XOR U13589 ( .A(n12794), .B(n12793), .Z(n12768) );
  XNOR U13590 ( .A(n12796), .B(n12768), .Z(N295) );
  NAND U13591 ( .A(n12770), .B(n12769), .Z(n12774) );
  NAND U13592 ( .A(n12772), .B(n12771), .Z(n12773) );
  AND U13593 ( .A(n12774), .B(n12773), .Z(n12810) );
  AND U13594 ( .A(y[1922]), .B(x[229]), .Z(n12899) );
  NAND U13595 ( .A(y[1926]), .B(x[225]), .Z(n12775) );
  XNOR U13596 ( .A(n12899), .B(n12775), .Z(n12824) );
  AND U13597 ( .A(x[230]), .B(y[1921]), .Z(n12828) );
  XOR U13598 ( .A(o[135]), .B(n12828), .Z(n12823) );
  XNOR U13599 ( .A(n12824), .B(n12823), .Z(n12843) );
  AND U13600 ( .A(x[230]), .B(y[1926]), .Z(n13042) );
  NAND U13601 ( .A(n13329), .B(n13042), .Z(n12779) );
  NAND U13602 ( .A(n12777), .B(n12776), .Z(n12778) );
  AND U13603 ( .A(n12779), .B(n12778), .Z(n12842) );
  XOR U13604 ( .A(n12843), .B(n12842), .Z(n12844) );
  NAND U13605 ( .A(n12831), .B(n12832), .Z(n12783) );
  NAND U13606 ( .A(n12781), .B(n12780), .Z(n12782) );
  AND U13607 ( .A(n12783), .B(n12782), .Z(n12845) );
  XOR U13608 ( .A(n12844), .B(n12845), .Z(n12808) );
  AND U13609 ( .A(x[228]), .B(y[1925]), .Z(n13334) );
  NAND U13610 ( .A(n13334), .B(n12822), .Z(n12787) );
  NAND U13611 ( .A(n12785), .B(n12784), .Z(n12786) );
  AND U13612 ( .A(n12787), .B(n12786), .Z(n12819) );
  AND U13613 ( .A(y[1925]), .B(x[226]), .Z(n12789) );
  NAND U13614 ( .A(y[1923]), .B(x[228]), .Z(n12788) );
  XNOR U13615 ( .A(n12789), .B(n12788), .Z(n12833) );
  XNOR U13616 ( .A(n12833), .B(n12832), .Z(n12817) );
  AND U13617 ( .A(y[1920]), .B(x[231]), .Z(n12791) );
  NAND U13618 ( .A(y[1927]), .B(x[224]), .Z(n12790) );
  XNOR U13619 ( .A(n12791), .B(n12790), .Z(n12837) );
  AND U13620 ( .A(o[134]), .B(n12792), .Z(n12836) );
  XNOR U13621 ( .A(n12837), .B(n12836), .Z(n12816) );
  XOR U13622 ( .A(n12817), .B(n12816), .Z(n12818) );
  XOR U13623 ( .A(n12819), .B(n12818), .Z(n12807) );
  XOR U13624 ( .A(n12808), .B(n12807), .Z(n12809) );
  XNOR U13625 ( .A(n12810), .B(n12809), .Z(n12815) );
  NANDN U13626 ( .A(n12793), .B(n12794), .Z(n12799) );
  NOR U13627 ( .A(n12795), .B(n12794), .Z(n12797) );
  OR U13628 ( .A(n12797), .B(n12796), .Z(n12798) );
  AND U13629 ( .A(n12799), .B(n12798), .Z(n12814) );
  NAND U13630 ( .A(n12801), .B(n12800), .Z(n12805) );
  NAND U13631 ( .A(n12803), .B(n12802), .Z(n12804) );
  AND U13632 ( .A(n12805), .B(n12804), .Z(n12813) );
  XOR U13633 ( .A(n12814), .B(n12813), .Z(n12806) );
  XNOR U13634 ( .A(n12815), .B(n12806), .Z(N296) );
  NAND U13635 ( .A(n12808), .B(n12807), .Z(n12812) );
  NAND U13636 ( .A(n12810), .B(n12809), .Z(n12811) );
  AND U13637 ( .A(n12812), .B(n12811), .Z(n12856) );
  NAND U13638 ( .A(n12817), .B(n12816), .Z(n12821) );
  NAND U13639 ( .A(n12819), .B(n12818), .Z(n12820) );
  AND U13640 ( .A(n12821), .B(n12820), .Z(n12889) );
  AND U13641 ( .A(x[229]), .B(y[1926]), .Z(n12992) );
  NAND U13642 ( .A(n12992), .B(n12822), .Z(n12826) );
  NAND U13643 ( .A(n12824), .B(n12823), .Z(n12825) );
  NAND U13644 ( .A(n12826), .B(n12825), .Z(n12887) );
  AND U13645 ( .A(y[1923]), .B(x[229]), .Z(n13487) );
  NAND U13646 ( .A(y[1927]), .B(x[225]), .Z(n12827) );
  XNOR U13647 ( .A(n13487), .B(n12827), .Z(n12877) );
  AND U13648 ( .A(o[135]), .B(n12828), .Z(n12876) );
  XOR U13649 ( .A(n12877), .B(n12876), .Z(n12864) );
  NAND U13650 ( .A(x[227]), .B(y[1925]), .Z(n13672) );
  AND U13651 ( .A(y[1922]), .B(x[230]), .Z(n12830) );
  NAND U13652 ( .A(y[1926]), .B(x[226]), .Z(n12829) );
  XNOR U13653 ( .A(n12830), .B(n12829), .Z(n12859) );
  XNOR U13654 ( .A(n13545), .B(n12859), .Z(n12862) );
  XOR U13655 ( .A(n13672), .B(n12862), .Z(n12863) );
  XOR U13656 ( .A(n12864), .B(n12863), .Z(n12886) );
  XOR U13657 ( .A(n12887), .B(n12886), .Z(n12888) );
  XNOR U13658 ( .A(n12889), .B(n12888), .Z(n12852) );
  NAND U13659 ( .A(n12831), .B(n13334), .Z(n12835) );
  NAND U13660 ( .A(n12833), .B(n12832), .Z(n12834) );
  NAND U13661 ( .A(n12835), .B(n12834), .Z(n12883) );
  AND U13662 ( .A(x[231]), .B(y[1927]), .Z(n13204) );
  NAND U13663 ( .A(n13329), .B(n13204), .Z(n12839) );
  NAND U13664 ( .A(n12837), .B(n12836), .Z(n12838) );
  NAND U13665 ( .A(n12839), .B(n12838), .Z(n12881) );
  AND U13666 ( .A(y[1920]), .B(x[232]), .Z(n12841) );
  NAND U13667 ( .A(y[1928]), .B(x[224]), .Z(n12840) );
  XNOR U13668 ( .A(n12841), .B(n12840), .Z(n12867) );
  AND U13669 ( .A(x[231]), .B(y[1921]), .Z(n12872) );
  XOR U13670 ( .A(o[136]), .B(n12872), .Z(n12866) );
  XOR U13671 ( .A(n12867), .B(n12866), .Z(n12880) );
  XOR U13672 ( .A(n12881), .B(n12880), .Z(n12882) );
  XNOR U13673 ( .A(n12883), .B(n12882), .Z(n12850) );
  NAND U13674 ( .A(n12843), .B(n12842), .Z(n12847) );
  NAND U13675 ( .A(n12845), .B(n12844), .Z(n12846) );
  NAND U13676 ( .A(n12847), .B(n12846), .Z(n12849) );
  XOR U13677 ( .A(n12850), .B(n12849), .Z(n12851) );
  XOR U13678 ( .A(n12852), .B(n12851), .Z(n12857) );
  XNOR U13679 ( .A(n12855), .B(n12857), .Z(n12848) );
  XOR U13680 ( .A(n12856), .B(n12848), .Z(N297) );
  NAND U13681 ( .A(n12850), .B(n12849), .Z(n12854) );
  NAND U13682 ( .A(n12852), .B(n12851), .Z(n12853) );
  NAND U13683 ( .A(n12854), .B(n12853), .Z(n12943) );
  IV U13684 ( .A(n12943), .Z(n12941) );
  NAND U13685 ( .A(n13042), .B(n12858), .Z(n12861) );
  NAND U13686 ( .A(n13545), .B(n12859), .Z(n12860) );
  NAND U13687 ( .A(n12861), .B(n12860), .Z(n12894) );
  XOR U13688 ( .A(n12894), .B(n12893), .Z(n12896) );
  AND U13689 ( .A(x[232]), .B(y[1928]), .Z(n12865) );
  NAND U13690 ( .A(n12865), .B(n13329), .Z(n12869) );
  NAND U13691 ( .A(n12867), .B(n12866), .Z(n12868) );
  AND U13692 ( .A(n12869), .B(n12868), .Z(n12928) );
  AND U13693 ( .A(y[1924]), .B(x[229]), .Z(n12871) );
  NAND U13694 ( .A(y[1922]), .B(x[231]), .Z(n12870) );
  XNOR U13695 ( .A(n12871), .B(n12870), .Z(n12901) );
  AND U13696 ( .A(o[136]), .B(n12872), .Z(n12900) );
  XNOR U13697 ( .A(n12901), .B(n12900), .Z(n12926) );
  AND U13698 ( .A(y[1920]), .B(x[233]), .Z(n12874) );
  NAND U13699 ( .A(y[1929]), .B(x[224]), .Z(n12873) );
  XNOR U13700 ( .A(n12874), .B(n12873), .Z(n12908) );
  NAND U13701 ( .A(x[232]), .B(y[1921]), .Z(n12915) );
  XNOR U13702 ( .A(n12908), .B(n12907), .Z(n12925) );
  XOR U13703 ( .A(n12926), .B(n12925), .Z(n12927) );
  XNOR U13704 ( .A(n12928), .B(n12927), .Z(n12922) );
  AND U13705 ( .A(y[1923]), .B(x[230]), .Z(n13273) );
  NAND U13706 ( .A(y[1928]), .B(x[225]), .Z(n12875) );
  XNOR U13707 ( .A(n13273), .B(n12875), .Z(n12912) );
  XNOR U13708 ( .A(n13334), .B(n12912), .Z(n12932) );
  NAND U13709 ( .A(x[226]), .B(y[1927]), .Z(n13592) );
  AND U13710 ( .A(x[227]), .B(y[1926]), .Z(n13283) );
  XNOR U13711 ( .A(n13592), .B(n13283), .Z(n12931) );
  XNOR U13712 ( .A(n12932), .B(n12931), .Z(n12920) );
  NAND U13713 ( .A(x[229]), .B(y[1927]), .Z(n13108) );
  AND U13714 ( .A(x[225]), .B(y[1923]), .Z(n12911) );
  NANDN U13715 ( .A(n13108), .B(n12911), .Z(n12879) );
  NAND U13716 ( .A(n12877), .B(n12876), .Z(n12878) );
  NAND U13717 ( .A(n12879), .B(n12878), .Z(n12919) );
  XOR U13718 ( .A(n12920), .B(n12919), .Z(n12921) );
  XOR U13719 ( .A(n12922), .B(n12921), .Z(n12895) );
  XOR U13720 ( .A(n12896), .B(n12895), .Z(n12938) );
  NAND U13721 ( .A(n12881), .B(n12880), .Z(n12885) );
  NAND U13722 ( .A(n12883), .B(n12882), .Z(n12884) );
  NAND U13723 ( .A(n12885), .B(n12884), .Z(n12936) );
  NAND U13724 ( .A(n12887), .B(n12886), .Z(n12891) );
  NAND U13725 ( .A(n12889), .B(n12888), .Z(n12890) );
  NAND U13726 ( .A(n12891), .B(n12890), .Z(n12935) );
  XOR U13727 ( .A(n12936), .B(n12935), .Z(n12937) );
  XOR U13728 ( .A(n12938), .B(n12937), .Z(n12944) );
  XNOR U13729 ( .A(n12942), .B(n12944), .Z(n12892) );
  XOR U13730 ( .A(n12941), .B(n12892), .Z(N298) );
  NAND U13731 ( .A(n12894), .B(n12893), .Z(n12898) );
  NAND U13732 ( .A(n12896), .B(n12895), .Z(n12897) );
  AND U13733 ( .A(n12898), .B(n12897), .Z(n12952) );
  AND U13734 ( .A(x[231]), .B(y[1924]), .Z(n12994) );
  NAND U13735 ( .A(n12994), .B(n12899), .Z(n12903) );
  NAND U13736 ( .A(n12901), .B(n12900), .Z(n12902) );
  AND U13737 ( .A(n12903), .B(n12902), .Z(n13007) );
  AND U13738 ( .A(y[1923]), .B(x[231]), .Z(n12905) );
  NAND U13739 ( .A(y[1926]), .B(x[228]), .Z(n12904) );
  XNOR U13740 ( .A(n12905), .B(n12904), .Z(n12978) );
  AND U13741 ( .A(x[230]), .B(y[1924]), .Z(n12977) );
  XOR U13742 ( .A(n12978), .B(n12977), .Z(n13005) );
  AND U13743 ( .A(x[232]), .B(y[1922]), .Z(n13177) );
  AND U13744 ( .A(x[233]), .B(y[1921]), .Z(n12988) );
  XOR U13745 ( .A(n12988), .B(o[138]), .Z(n12999) );
  XOR U13746 ( .A(n13177), .B(n12999), .Z(n13001) );
  XNOR U13747 ( .A(n13001), .B(n13000), .Z(n13004) );
  XNOR U13748 ( .A(n13007), .B(n13006), .Z(n12967) );
  AND U13749 ( .A(x[233]), .B(y[1929]), .Z(n12906) );
  NAND U13750 ( .A(n12906), .B(n13329), .Z(n12910) );
  NAND U13751 ( .A(n12908), .B(n12907), .Z(n12909) );
  NAND U13752 ( .A(n12910), .B(n12909), .Z(n12965) );
  AND U13753 ( .A(x[230]), .B(y[1928]), .Z(n13214) );
  NAND U13754 ( .A(n13214), .B(n12911), .Z(n12914) );
  NAND U13755 ( .A(n13334), .B(n12912), .Z(n12913) );
  NAND U13756 ( .A(n12914), .B(n12913), .Z(n12972) );
  ANDN U13757 ( .B(o[137]), .A(n12915), .Z(n12983) );
  AND U13758 ( .A(y[1920]), .B(x[234]), .Z(n12917) );
  AND U13759 ( .A(y[1930]), .B(x[224]), .Z(n12916) );
  XOR U13760 ( .A(n12917), .B(n12916), .Z(n12982) );
  XOR U13761 ( .A(n12983), .B(n12982), .Z(n12971) );
  AND U13762 ( .A(y[1927]), .B(x[227]), .Z(n13900) );
  NAND U13763 ( .A(y[1929]), .B(x[225]), .Z(n12918) );
  XNOR U13764 ( .A(n13900), .B(n12918), .Z(n12996) );
  AND U13765 ( .A(x[226]), .B(y[1928]), .Z(n12995) );
  XOR U13766 ( .A(n12996), .B(n12995), .Z(n12970) );
  XOR U13767 ( .A(n12971), .B(n12970), .Z(n12973) );
  XOR U13768 ( .A(n12972), .B(n12973), .Z(n12964) );
  XOR U13769 ( .A(n12965), .B(n12964), .Z(n12966) );
  XNOR U13770 ( .A(n12967), .B(n12966), .Z(n12950) );
  NAND U13771 ( .A(n12920), .B(n12919), .Z(n12924) );
  NAND U13772 ( .A(n12922), .B(n12921), .Z(n12923) );
  AND U13773 ( .A(n12924), .B(n12923), .Z(n12961) );
  NAND U13774 ( .A(n12926), .B(n12925), .Z(n12930) );
  NAND U13775 ( .A(n12928), .B(n12927), .Z(n12929) );
  AND U13776 ( .A(n12930), .B(n12929), .Z(n12958) );
  NAND U13777 ( .A(n12932), .B(n12931), .Z(n12934) );
  ANDN U13778 ( .B(n13592), .A(n13283), .Z(n12933) );
  ANDN U13779 ( .B(n12934), .A(n12933), .Z(n12959) );
  XOR U13780 ( .A(n12958), .B(n12959), .Z(n12960) );
  XOR U13781 ( .A(n12961), .B(n12960), .Z(n12949) );
  XOR U13782 ( .A(n12950), .B(n12949), .Z(n12951) );
  XOR U13783 ( .A(n12952), .B(n12951), .Z(n12957) );
  NAND U13784 ( .A(n12936), .B(n12935), .Z(n12940) );
  NAND U13785 ( .A(n12938), .B(n12937), .Z(n12939) );
  NAND U13786 ( .A(n12940), .B(n12939), .Z(n12956) );
  NANDN U13787 ( .A(n12941), .B(n12942), .Z(n12947) );
  NOR U13788 ( .A(n12943), .B(n12942), .Z(n12945) );
  OR U13789 ( .A(n12945), .B(n12944), .Z(n12946) );
  AND U13790 ( .A(n12947), .B(n12946), .Z(n12955) );
  XOR U13791 ( .A(n12956), .B(n12955), .Z(n12948) );
  XNOR U13792 ( .A(n12957), .B(n12948), .Z(N299) );
  NAND U13793 ( .A(n12950), .B(n12949), .Z(n12954) );
  NAND U13794 ( .A(n12952), .B(n12951), .Z(n12953) );
  NAND U13795 ( .A(n12954), .B(n12953), .Z(n13074) );
  IV U13796 ( .A(n13074), .Z(n13072) );
  NAND U13797 ( .A(n12959), .B(n12958), .Z(n12963) );
  NANDN U13798 ( .A(n12961), .B(n12960), .Z(n12962) );
  NAND U13799 ( .A(n12963), .B(n12962), .Z(n13069) );
  NAND U13800 ( .A(n12965), .B(n12964), .Z(n12969) );
  NAND U13801 ( .A(n12967), .B(n12966), .Z(n12968) );
  NAND U13802 ( .A(n12969), .B(n12968), .Z(n13067) );
  NAND U13803 ( .A(n12971), .B(n12970), .Z(n12975) );
  NAND U13804 ( .A(n12973), .B(n12972), .Z(n12974) );
  NAND U13805 ( .A(n12975), .B(n12974), .Z(n13062) );
  AND U13806 ( .A(x[231]), .B(y[1926]), .Z(n13104) );
  AND U13807 ( .A(x[228]), .B(y[1923]), .Z(n12976) );
  NAND U13808 ( .A(n13104), .B(n12976), .Z(n12980) );
  NAND U13809 ( .A(n12978), .B(n12977), .Z(n12979) );
  NAND U13810 ( .A(n12980), .B(n12979), .Z(n13060) );
  AND U13811 ( .A(x[234]), .B(y[1930]), .Z(n12981) );
  NAND U13812 ( .A(n12981), .B(n13329), .Z(n12985) );
  NAND U13813 ( .A(n12983), .B(n12982), .Z(n12984) );
  NAND U13814 ( .A(n12985), .B(n12984), .Z(n13056) );
  AND U13815 ( .A(y[1920]), .B(x[235]), .Z(n12987) );
  NAND U13816 ( .A(y[1931]), .B(x[224]), .Z(n12986) );
  XNOR U13817 ( .A(n12987), .B(n12986), .Z(n13031) );
  AND U13818 ( .A(n12988), .B(o[138]), .Z(n13032) );
  XOR U13819 ( .A(n13031), .B(n13032), .Z(n13055) );
  AND U13820 ( .A(y[1925]), .B(x[230]), .Z(n12990) );
  NAND U13821 ( .A(y[1930]), .B(x[225]), .Z(n12989) );
  XNOR U13822 ( .A(n12990), .B(n12989), .Z(n13023) );
  AND U13823 ( .A(x[234]), .B(y[1921]), .Z(n13040) );
  XOR U13824 ( .A(o[139]), .B(n13040), .Z(n13022) );
  XOR U13825 ( .A(n13023), .B(n13022), .Z(n13054) );
  XOR U13826 ( .A(n13055), .B(n13054), .Z(n13057) );
  XOR U13827 ( .A(n13056), .B(n13057), .Z(n13061) );
  XOR U13828 ( .A(n13060), .B(n13061), .Z(n13063) );
  XNOR U13829 ( .A(n13062), .B(n13063), .Z(n13045) );
  NAND U13830 ( .A(x[227]), .B(y[1928]), .Z(n14006) );
  NAND U13831 ( .A(y[1929]), .B(x[226]), .Z(n12991) );
  XNOR U13832 ( .A(n12992), .B(n12991), .Z(n13018) );
  AND U13833 ( .A(x[228]), .B(y[1927]), .Z(n13017) );
  XNOR U13834 ( .A(n13018), .B(n13017), .Z(n13049) );
  XOR U13835 ( .A(n14006), .B(n13049), .Z(n13050) );
  NAND U13836 ( .A(y[1922]), .B(x[233]), .Z(n12993) );
  XNOR U13837 ( .A(n12994), .B(n12993), .Z(n13036) );
  AND U13838 ( .A(x[232]), .B(y[1923]), .Z(n13037) );
  XOR U13839 ( .A(n13036), .B(n13037), .Z(n13051) );
  AND U13840 ( .A(x[227]), .B(y[1929]), .Z(n13099) );
  AND U13841 ( .A(x[225]), .B(y[1927]), .Z(n13324) );
  NAND U13842 ( .A(n13099), .B(n13324), .Z(n12998) );
  NAND U13843 ( .A(n12996), .B(n12995), .Z(n12997) );
  NAND U13844 ( .A(n12998), .B(n12997), .Z(n13012) );
  NAND U13845 ( .A(n13177), .B(n12999), .Z(n13003) );
  NAND U13846 ( .A(n13001), .B(n13000), .Z(n13002) );
  NAND U13847 ( .A(n13003), .B(n13002), .Z(n13011) );
  XOR U13848 ( .A(n13012), .B(n13011), .Z(n13013) );
  NANDN U13849 ( .A(n13005), .B(n13004), .Z(n13009) );
  NAND U13850 ( .A(n13007), .B(n13006), .Z(n13008) );
  NAND U13851 ( .A(n13009), .B(n13008), .Z(n13043) );
  XOR U13852 ( .A(n13045), .B(n13046), .Z(n13066) );
  XOR U13853 ( .A(n13067), .B(n13066), .Z(n13068) );
  XOR U13854 ( .A(n13069), .B(n13068), .Z(n13075) );
  XNOR U13855 ( .A(n13073), .B(n13075), .Z(n13010) );
  XOR U13856 ( .A(n13072), .B(n13010), .Z(N300) );
  NAND U13857 ( .A(n13012), .B(n13011), .Z(n13016) );
  NANDN U13858 ( .A(n13014), .B(n13013), .Z(n13015) );
  NAND U13859 ( .A(n13016), .B(n13015), .Z(n13139) );
  AND U13860 ( .A(x[226]), .B(y[1926]), .Z(n13759) );
  AND U13861 ( .A(x[229]), .B(y[1929]), .Z(n13583) );
  NAND U13862 ( .A(n13759), .B(n13583), .Z(n13020) );
  NAND U13863 ( .A(n13018), .B(n13017), .Z(n13019) );
  AND U13864 ( .A(n13020), .B(n13019), .Z(n13087) );
  AND U13865 ( .A(x[230]), .B(y[1930]), .Z(n13341) );
  NAND U13866 ( .A(n13341), .B(n13021), .Z(n13025) );
  NAND U13867 ( .A(n13023), .B(n13022), .Z(n13024) );
  NAND U13868 ( .A(n13025), .B(n13024), .Z(n13086) );
  AND U13869 ( .A(x[233]), .B(y[1923]), .Z(n13754) );
  AND U13870 ( .A(y[1922]), .B(x[234]), .Z(n13795) );
  NAND U13871 ( .A(y[1928]), .B(x[228]), .Z(n13026) );
  XNOR U13872 ( .A(n13795), .B(n13026), .Z(n13130) );
  XOR U13873 ( .A(n13754), .B(n13130), .Z(n13109) );
  NAND U13874 ( .A(x[231]), .B(y[1925]), .Z(n13107) );
  XOR U13875 ( .A(n13108), .B(n13107), .Z(n13110) );
  AND U13876 ( .A(y[1920]), .B(x[236]), .Z(n13028) );
  NAND U13877 ( .A(y[1932]), .B(x[224]), .Z(n13027) );
  XNOR U13878 ( .A(n13028), .B(n13027), .Z(n13124) );
  AND U13879 ( .A(x[235]), .B(y[1921]), .Z(n13102) );
  XOR U13880 ( .A(o[140]), .B(n13102), .Z(n13123) );
  XOR U13881 ( .A(n13124), .B(n13123), .Z(n13093) );
  AND U13882 ( .A(y[1930]), .B(x[226]), .Z(n13030) );
  NAND U13883 ( .A(y[1924]), .B(x[232]), .Z(n13029) );
  XNOR U13884 ( .A(n13030), .B(n13029), .Z(n13098) );
  XOR U13885 ( .A(n13098), .B(n13099), .Z(n13092) );
  XOR U13886 ( .A(n13093), .B(n13092), .Z(n13095) );
  XOR U13887 ( .A(n13094), .B(n13095), .Z(n13088) );
  XOR U13888 ( .A(n13089), .B(n13088), .Z(n13137) );
  AND U13889 ( .A(x[235]), .B(y[1931]), .Z(n14146) );
  NAND U13890 ( .A(n14146), .B(n13329), .Z(n13034) );
  NAND U13891 ( .A(n13032), .B(n13031), .Z(n13033) );
  NAND U13892 ( .A(n13034), .B(n13033), .Z(n13116) );
  AND U13893 ( .A(x[231]), .B(y[1922]), .Z(n13259) );
  AND U13894 ( .A(x[233]), .B(y[1924]), .Z(n13035) );
  NAND U13895 ( .A(n13259), .B(n13035), .Z(n13039) );
  NAND U13896 ( .A(n13037), .B(n13036), .Z(n13038) );
  NAND U13897 ( .A(n13039), .B(n13038), .Z(n13114) );
  AND U13898 ( .A(o[139]), .B(n13040), .Z(n13119) );
  NAND U13899 ( .A(y[1931]), .B(x[225]), .Z(n13041) );
  XNOR U13900 ( .A(n13042), .B(n13041), .Z(n13120) );
  XOR U13901 ( .A(n13119), .B(n13120), .Z(n13113) );
  XOR U13902 ( .A(n13114), .B(n13113), .Z(n13115) );
  XNOR U13903 ( .A(n13116), .B(n13115), .Z(n13138) );
  XNOR U13904 ( .A(n13137), .B(n13138), .Z(n13140) );
  XOR U13905 ( .A(n13139), .B(n13140), .Z(n13147) );
  NANDN U13906 ( .A(n13044), .B(n13043), .Z(n13048) );
  NANDN U13907 ( .A(n13046), .B(n13045), .Z(n13047) );
  NAND U13908 ( .A(n13048), .B(n13047), .Z(n13146) );
  IV U13909 ( .A(n14006), .Z(n13768) );
  NANDN U13910 ( .A(n13768), .B(n13049), .Z(n13053) );
  NANDN U13911 ( .A(n13051), .B(n13050), .Z(n13052) );
  NAND U13912 ( .A(n13053), .B(n13052), .Z(n13080) );
  NAND U13913 ( .A(n13055), .B(n13054), .Z(n13059) );
  NAND U13914 ( .A(n13057), .B(n13056), .Z(n13058) );
  AND U13915 ( .A(n13059), .B(n13058), .Z(n13081) );
  XOR U13916 ( .A(n13080), .B(n13081), .Z(n13083) );
  NAND U13917 ( .A(n13061), .B(n13060), .Z(n13065) );
  NAND U13918 ( .A(n13063), .B(n13062), .Z(n13064) );
  AND U13919 ( .A(n13065), .B(n13064), .Z(n13082) );
  XOR U13920 ( .A(n13083), .B(n13082), .Z(n13148) );
  XOR U13921 ( .A(n13149), .B(n13148), .Z(n13145) );
  NAND U13922 ( .A(n13067), .B(n13066), .Z(n13071) );
  NAND U13923 ( .A(n13069), .B(n13068), .Z(n13070) );
  NAND U13924 ( .A(n13071), .B(n13070), .Z(n13144) );
  NANDN U13925 ( .A(n13072), .B(n13073), .Z(n13078) );
  NOR U13926 ( .A(n13074), .B(n13073), .Z(n13076) );
  OR U13927 ( .A(n13076), .B(n13075), .Z(n13077) );
  AND U13928 ( .A(n13078), .B(n13077), .Z(n13143) );
  XOR U13929 ( .A(n13144), .B(n13143), .Z(n13079) );
  XNOR U13930 ( .A(n13145), .B(n13079), .Z(N301) );
  NAND U13931 ( .A(n13081), .B(n13080), .Z(n13085) );
  NAND U13932 ( .A(n13083), .B(n13082), .Z(n13084) );
  NAND U13933 ( .A(n13085), .B(n13084), .Z(n13230) );
  NANDN U13934 ( .A(n13087), .B(n13086), .Z(n13091) );
  NAND U13935 ( .A(n13089), .B(n13088), .Z(n13090) );
  AND U13936 ( .A(n13091), .B(n13090), .Z(n13154) );
  NAND U13937 ( .A(n13093), .B(n13092), .Z(n13097) );
  NAND U13938 ( .A(n13095), .B(n13094), .Z(n13096) );
  NAND U13939 ( .A(n13097), .B(n13096), .Z(n13161) );
  AND U13940 ( .A(y[1930]), .B(x[232]), .Z(n14417) );
  AND U13941 ( .A(x[226]), .B(y[1924]), .Z(n13269) );
  NAND U13942 ( .A(n14417), .B(n13269), .Z(n13101) );
  NAND U13943 ( .A(n13099), .B(n13098), .Z(n13100) );
  NAND U13944 ( .A(n13101), .B(n13100), .Z(n13193) );
  AND U13945 ( .A(o[140]), .B(n13102), .Z(n13183) );
  AND U13946 ( .A(y[1932]), .B(x[225]), .Z(n13103) );
  XOR U13947 ( .A(n13104), .B(n13103), .Z(n13182) );
  XOR U13948 ( .A(n13183), .B(n13182), .Z(n13191) );
  AND U13949 ( .A(x[230]), .B(y[1927]), .Z(n14185) );
  AND U13950 ( .A(y[1931]), .B(x[226]), .Z(n13106) );
  NAND U13951 ( .A(y[1924]), .B(x[233]), .Z(n13105) );
  XNOR U13952 ( .A(n13106), .B(n13105), .Z(n13197) );
  XOR U13953 ( .A(n14185), .B(n13197), .Z(n13190) );
  XOR U13954 ( .A(n13191), .B(n13190), .Z(n13192) );
  XOR U13955 ( .A(n13193), .B(n13192), .Z(n13160) );
  NAND U13956 ( .A(n13108), .B(n13107), .Z(n13112) );
  ANDN U13957 ( .B(n13110), .A(n13109), .Z(n13111) );
  ANDN U13958 ( .B(n13112), .A(n13111), .Z(n13159) );
  XOR U13959 ( .A(n13160), .B(n13159), .Z(n13162) );
  XOR U13960 ( .A(n13161), .B(n13162), .Z(n13153) );
  NAND U13961 ( .A(n13114), .B(n13113), .Z(n13118) );
  NAND U13962 ( .A(n13116), .B(n13115), .Z(n13117) );
  NAND U13963 ( .A(n13118), .B(n13117), .Z(n13168) );
  AND U13964 ( .A(x[230]), .B(y[1931]), .Z(n13466) );
  IV U13965 ( .A(n13466), .Z(n13585) );
  AND U13966 ( .A(x[225]), .B(y[1926]), .Z(n13181) );
  NANDN U13967 ( .A(n13585), .B(n13181), .Z(n13122) );
  NAND U13968 ( .A(n13120), .B(n13119), .Z(n13121) );
  NAND U13969 ( .A(n13122), .B(n13121), .Z(n13174) );
  AND U13970 ( .A(x[236]), .B(y[1932]), .Z(n14423) );
  NAND U13971 ( .A(n14423), .B(n13329), .Z(n13126) );
  NAND U13972 ( .A(n13124), .B(n13123), .Z(n13125) );
  NAND U13973 ( .A(n13126), .B(n13125), .Z(n13172) );
  AND U13974 ( .A(x[234]), .B(y[1923]), .Z(n14018) );
  AND U13975 ( .A(y[1922]), .B(x[235]), .Z(n14028) );
  NAND U13976 ( .A(y[1925]), .B(x[232]), .Z(n13127) );
  XNOR U13977 ( .A(n14028), .B(n13127), .Z(n13178) );
  XOR U13978 ( .A(n14018), .B(n13178), .Z(n13171) );
  XOR U13979 ( .A(n13172), .B(n13171), .Z(n13173) );
  XOR U13980 ( .A(n13174), .B(n13173), .Z(n13166) );
  AND U13981 ( .A(x[234]), .B(y[1928]), .Z(n13129) );
  AND U13982 ( .A(x[228]), .B(y[1922]), .Z(n13128) );
  NAND U13983 ( .A(n13129), .B(n13128), .Z(n13132) );
  NAND U13984 ( .A(n13130), .B(n13754), .Z(n13131) );
  NAND U13985 ( .A(n13132), .B(n13131), .Z(n13218) );
  AND U13986 ( .A(y[1920]), .B(x[237]), .Z(n13134) );
  NAND U13987 ( .A(y[1933]), .B(x[224]), .Z(n13133) );
  XNOR U13988 ( .A(n13134), .B(n13133), .Z(n13210) );
  AND U13989 ( .A(x[236]), .B(y[1921]), .Z(n13202) );
  XOR U13990 ( .A(o[141]), .B(n13202), .Z(n13209) );
  XOR U13991 ( .A(n13210), .B(n13209), .Z(n13216) );
  AND U13992 ( .A(y[1928]), .B(x[229]), .Z(n13136) );
  NAND U13993 ( .A(y[1930]), .B(x[227]), .Z(n13135) );
  XNOR U13994 ( .A(n13136), .B(n13135), .Z(n13205) );
  AND U13995 ( .A(x[228]), .B(y[1929]), .Z(n13206) );
  XOR U13996 ( .A(n13205), .B(n13206), .Z(n13215) );
  XOR U13997 ( .A(n13216), .B(n13215), .Z(n13217) );
  XOR U13998 ( .A(n13218), .B(n13217), .Z(n13165) );
  XOR U13999 ( .A(n13166), .B(n13165), .Z(n13167) );
  XOR U14000 ( .A(n13168), .B(n13167), .Z(n13155) );
  XOR U14001 ( .A(n13156), .B(n13155), .Z(n13229) );
  NANDN U14002 ( .A(n13138), .B(n13137), .Z(n13142) );
  NAND U14003 ( .A(n13140), .B(n13139), .Z(n13141) );
  AND U14004 ( .A(n13142), .B(n13141), .Z(n13228) );
  XOR U14005 ( .A(n13230), .B(n13231), .Z(n13224) );
  NANDN U14006 ( .A(n13147), .B(n13146), .Z(n13151) );
  NAND U14007 ( .A(n13149), .B(n13148), .Z(n13150) );
  AND U14008 ( .A(n13151), .B(n13150), .Z(n13222) );
  IV U14009 ( .A(n13222), .Z(n13221) );
  XOR U14010 ( .A(n13223), .B(n13221), .Z(n13152) );
  XNOR U14011 ( .A(n13224), .B(n13152), .Z(N302) );
  NANDN U14012 ( .A(n13154), .B(n13153), .Z(n13158) );
  NAND U14013 ( .A(n13156), .B(n13155), .Z(n13157) );
  AND U14014 ( .A(n13158), .B(n13157), .Z(n13318) );
  NAND U14015 ( .A(n13160), .B(n13159), .Z(n13164) );
  NAND U14016 ( .A(n13162), .B(n13161), .Z(n13163) );
  NAND U14017 ( .A(n13164), .B(n13163), .Z(n13317) );
  NAND U14018 ( .A(n13166), .B(n13165), .Z(n13170) );
  NAND U14019 ( .A(n13168), .B(n13167), .Z(n13169) );
  NAND U14020 ( .A(n13170), .B(n13169), .Z(n13238) );
  NAND U14021 ( .A(n13172), .B(n13171), .Z(n13176) );
  NAND U14022 ( .A(n13174), .B(n13173), .Z(n13175) );
  AND U14023 ( .A(n13176), .B(n13175), .Z(n13244) );
  AND U14024 ( .A(x[235]), .B(y[1925]), .Z(n13355) );
  NAND U14025 ( .A(n13355), .B(n13177), .Z(n13180) );
  NAND U14026 ( .A(n13178), .B(n14018), .Z(n13179) );
  NAND U14027 ( .A(n13180), .B(n13179), .Z(n13299) );
  NAND U14028 ( .A(x[231]), .B(y[1932]), .Z(n13770) );
  NANDN U14029 ( .A(n13770), .B(n13181), .Z(n13185) );
  NAND U14030 ( .A(n13183), .B(n13182), .Z(n13184) );
  NAND U14031 ( .A(n13185), .B(n13184), .Z(n13298) );
  XOR U14032 ( .A(n13299), .B(n13298), .Z(n13301) );
  AND U14033 ( .A(x[228]), .B(y[1930]), .Z(n13681) );
  AND U14034 ( .A(y[1931]), .B(x[227]), .Z(n13187) );
  NAND U14035 ( .A(y[1926]), .B(x[232]), .Z(n13186) );
  XNOR U14036 ( .A(n13187), .B(n13186), .Z(n13284) );
  XOR U14037 ( .A(n13583), .B(n13284), .Z(n13293) );
  XOR U14038 ( .A(n13681), .B(n13293), .Z(n13295) );
  AND U14039 ( .A(x[233]), .B(y[1925]), .Z(n13871) );
  AND U14040 ( .A(y[1932]), .B(x[226]), .Z(n13189) );
  NAND U14041 ( .A(y[1924]), .B(x[234]), .Z(n13188) );
  XNOR U14042 ( .A(n13189), .B(n13188), .Z(n13270) );
  XOR U14043 ( .A(n13871), .B(n13270), .Z(n13294) );
  XOR U14044 ( .A(n13295), .B(n13294), .Z(n13300) );
  XNOR U14045 ( .A(n13301), .B(n13300), .Z(n13242) );
  NAND U14046 ( .A(n13191), .B(n13190), .Z(n13195) );
  NAND U14047 ( .A(n13193), .B(n13192), .Z(n13194) );
  AND U14048 ( .A(n13195), .B(n13194), .Z(n13241) );
  XOR U14049 ( .A(n13242), .B(n13241), .Z(n13243) );
  XNOR U14050 ( .A(n13244), .B(n13243), .Z(n13236) );
  AND U14051 ( .A(x[233]), .B(y[1931]), .Z(n13196) );
  NAND U14052 ( .A(n13196), .B(n13269), .Z(n13199) );
  NAND U14053 ( .A(n13197), .B(n14185), .Z(n13198) );
  NAND U14054 ( .A(n13199), .B(n13198), .Z(n13255) );
  AND U14055 ( .A(y[1920]), .B(x[238]), .Z(n13201) );
  NAND U14056 ( .A(y[1934]), .B(x[224]), .Z(n13200) );
  XNOR U14057 ( .A(n13201), .B(n13200), .Z(n13279) );
  AND U14058 ( .A(o[141]), .B(n13202), .Z(n13278) );
  XOR U14059 ( .A(n13279), .B(n13278), .Z(n13254) );
  NAND U14060 ( .A(y[1922]), .B(x[236]), .Z(n13203) );
  XNOR U14061 ( .A(n13204), .B(n13203), .Z(n13261) );
  AND U14062 ( .A(x[237]), .B(y[1921]), .Z(n13268) );
  XOR U14063 ( .A(o[142]), .B(n13268), .Z(n13260) );
  XOR U14064 ( .A(n13261), .B(n13260), .Z(n13253) );
  XOR U14065 ( .A(n13254), .B(n13253), .Z(n13256) );
  XNOR U14066 ( .A(n13255), .B(n13256), .Z(n13305) );
  AND U14067 ( .A(x[229]), .B(y[1930]), .Z(n13342) );
  NANDN U14068 ( .A(n14006), .B(n13342), .Z(n13208) );
  NAND U14069 ( .A(n13206), .B(n13205), .Z(n13207) );
  NAND U14070 ( .A(n13208), .B(n13207), .Z(n13249) );
  AND U14071 ( .A(x[237]), .B(y[1933]), .Z(n14719) );
  NAND U14072 ( .A(n14719), .B(n13329), .Z(n13212) );
  NAND U14073 ( .A(n13210), .B(n13209), .Z(n13211) );
  NAND U14074 ( .A(n13212), .B(n13211), .Z(n13247) );
  NAND U14075 ( .A(y[1923]), .B(x[235]), .Z(n13213) );
  XNOR U14076 ( .A(n13214), .B(n13213), .Z(n13275) );
  AND U14077 ( .A(x[225]), .B(y[1933]), .Z(n13274) );
  XOR U14078 ( .A(n13275), .B(n13274), .Z(n13248) );
  XNOR U14079 ( .A(n13247), .B(n13248), .Z(n13250) );
  XOR U14080 ( .A(n13249), .B(n13250), .Z(n13304) );
  XOR U14081 ( .A(n13305), .B(n13304), .Z(n13307) );
  NAND U14082 ( .A(n13216), .B(n13215), .Z(n13220) );
  NAND U14083 ( .A(n13218), .B(n13217), .Z(n13219) );
  AND U14084 ( .A(n13220), .B(n13219), .Z(n13306) );
  XNOR U14085 ( .A(n13307), .B(n13306), .Z(n13235) );
  XOR U14086 ( .A(n13236), .B(n13235), .Z(n13237) );
  XOR U14087 ( .A(n13238), .B(n13237), .Z(n13319) );
  XNOR U14088 ( .A(n13320), .B(n13319), .Z(n13313) );
  OR U14089 ( .A(n13223), .B(n13221), .Z(n13227) );
  ANDN U14090 ( .B(n13223), .A(n13222), .Z(n13225) );
  OR U14091 ( .A(n13225), .B(n13224), .Z(n13226) );
  AND U14092 ( .A(n13227), .B(n13226), .Z(n13312) );
  NANDN U14093 ( .A(n13229), .B(n13228), .Z(n13233) );
  NAND U14094 ( .A(n13231), .B(n13230), .Z(n13232) );
  AND U14095 ( .A(n13233), .B(n13232), .Z(n13311) );
  IV U14096 ( .A(n13311), .Z(n13310) );
  XOR U14097 ( .A(n13312), .B(n13310), .Z(n13234) );
  XNOR U14098 ( .A(n13313), .B(n13234), .Z(N303) );
  NAND U14099 ( .A(n13236), .B(n13235), .Z(n13240) );
  NAND U14100 ( .A(n13238), .B(n13237), .Z(n13239) );
  AND U14101 ( .A(n13240), .B(n13239), .Z(n13416) );
  NAND U14102 ( .A(n13242), .B(n13241), .Z(n13246) );
  NAND U14103 ( .A(n13244), .B(n13243), .Z(n13245) );
  NAND U14104 ( .A(n13246), .B(n13245), .Z(n13384) );
  NAND U14105 ( .A(n13248), .B(n13247), .Z(n13252) );
  NANDN U14106 ( .A(n13250), .B(n13249), .Z(n13251) );
  NAND U14107 ( .A(n13252), .B(n13251), .Z(n13390) );
  NAND U14108 ( .A(n13254), .B(n13253), .Z(n13258) );
  NAND U14109 ( .A(n13256), .B(n13255), .Z(n13257) );
  NAND U14110 ( .A(n13258), .B(n13257), .Z(n13388) );
  AND U14111 ( .A(x[236]), .B(y[1927]), .Z(n13760) );
  NAND U14112 ( .A(n13760), .B(n13259), .Z(n13263) );
  NAND U14113 ( .A(n13261), .B(n13260), .Z(n13262) );
  AND U14114 ( .A(n13263), .B(n13262), .Z(n13365) );
  AND U14115 ( .A(y[1924]), .B(x[235]), .Z(n13265) );
  NAND U14116 ( .A(y[1922]), .B(x[237]), .Z(n13264) );
  XNOR U14117 ( .A(n13265), .B(n13264), .Z(n13369) );
  AND U14118 ( .A(x[236]), .B(y[1923]), .Z(n13368) );
  XNOR U14119 ( .A(n13369), .B(n13368), .Z(n13363) );
  AND U14120 ( .A(y[1920]), .B(x[239]), .Z(n13267) );
  NAND U14121 ( .A(y[1935]), .B(x[224]), .Z(n13266) );
  XNOR U14122 ( .A(n13267), .B(n13266), .Z(n13331) );
  AND U14123 ( .A(o[142]), .B(n13268), .Z(n13330) );
  XNOR U14124 ( .A(n13331), .B(n13330), .Z(n13362) );
  XOR U14125 ( .A(n13363), .B(n13362), .Z(n13364) );
  XOR U14126 ( .A(n13365), .B(n13364), .Z(n13397) );
  AND U14127 ( .A(x[234]), .B(y[1932]), .Z(n14186) );
  NAND U14128 ( .A(n14186), .B(n13269), .Z(n13272) );
  NAND U14129 ( .A(n13871), .B(n13270), .Z(n13271) );
  NAND U14130 ( .A(n13272), .B(n13271), .Z(n13395) );
  AND U14131 ( .A(x[235]), .B(y[1928]), .Z(n13680) );
  NAND U14132 ( .A(n13680), .B(n13273), .Z(n13277) );
  NAND U14133 ( .A(n13275), .B(n13274), .Z(n13276) );
  NAND U14134 ( .A(n13277), .B(n13276), .Z(n13394) );
  XOR U14135 ( .A(n13395), .B(n13394), .Z(n13396) );
  XOR U14136 ( .A(n13388), .B(n13389), .Z(n13391) );
  XOR U14137 ( .A(n13390), .B(n13391), .Z(n13383) );
  AND U14138 ( .A(x[238]), .B(y[1934]), .Z(n14995) );
  NAND U14139 ( .A(n14995), .B(n13329), .Z(n13281) );
  NAND U14140 ( .A(n13279), .B(n13278), .Z(n13280) );
  NAND U14141 ( .A(n13281), .B(n13280), .Z(n13357) );
  AND U14142 ( .A(x[232]), .B(y[1931]), .Z(n13282) );
  NAND U14143 ( .A(n13283), .B(n13282), .Z(n13286) );
  NAND U14144 ( .A(n13583), .B(n13284), .Z(n13285) );
  NAND U14145 ( .A(n13286), .B(n13285), .Z(n13356) );
  XOR U14146 ( .A(n13357), .B(n13356), .Z(n13359) );
  AND U14147 ( .A(y[1925]), .B(x[234]), .Z(n13288) );
  NAND U14148 ( .A(y[1931]), .B(x[228]), .Z(n13287) );
  XNOR U14149 ( .A(n13288), .B(n13287), .Z(n13337) );
  AND U14150 ( .A(x[231]), .B(y[1928]), .Z(n13336) );
  XNOR U14151 ( .A(n13337), .B(n13336), .Z(n13344) );
  NAND U14152 ( .A(x[230]), .B(y[1929]), .Z(n13496) );
  XNOR U14153 ( .A(n13496), .B(n13342), .Z(n13343) );
  XNOR U14154 ( .A(n13344), .B(n13343), .Z(n13378) );
  AND U14155 ( .A(y[1933]), .B(x[226]), .Z(n13290) );
  NAND U14156 ( .A(y[1926]), .B(x[233]), .Z(n13289) );
  XNOR U14157 ( .A(n13290), .B(n13289), .Z(n13347) );
  AND U14158 ( .A(x[227]), .B(y[1932]), .Z(n13348) );
  XOR U14159 ( .A(n13347), .B(n13348), .Z(n13377) );
  AND U14160 ( .A(y[1934]), .B(x[225]), .Z(n13292) );
  NAND U14161 ( .A(y[1927]), .B(x[232]), .Z(n13291) );
  XNOR U14162 ( .A(n13292), .B(n13291), .Z(n13326) );
  AND U14163 ( .A(x[238]), .B(y[1921]), .Z(n13353) );
  XOR U14164 ( .A(o[143]), .B(n13353), .Z(n13325) );
  XOR U14165 ( .A(n13326), .B(n13325), .Z(n13376) );
  XOR U14166 ( .A(n13377), .B(n13376), .Z(n13379) );
  XOR U14167 ( .A(n13378), .B(n13379), .Z(n13358) );
  XOR U14168 ( .A(n13359), .B(n13358), .Z(n13401) );
  NAND U14169 ( .A(n13681), .B(n13293), .Z(n13297) );
  NAND U14170 ( .A(n13295), .B(n13294), .Z(n13296) );
  AND U14171 ( .A(n13297), .B(n13296), .Z(n13400) );
  NAND U14172 ( .A(n13299), .B(n13298), .Z(n13303) );
  NAND U14173 ( .A(n13301), .B(n13300), .Z(n13302) );
  AND U14174 ( .A(n13303), .B(n13302), .Z(n13402) );
  XOR U14175 ( .A(n13403), .B(n13402), .Z(n13382) );
  XOR U14176 ( .A(n13384), .B(n13385), .Z(n13413) );
  NAND U14177 ( .A(n13305), .B(n13304), .Z(n13309) );
  NAND U14178 ( .A(n13307), .B(n13306), .Z(n13308) );
  AND U14179 ( .A(n13309), .B(n13308), .Z(n13414) );
  XOR U14180 ( .A(n13413), .B(n13414), .Z(n13415) );
  XOR U14181 ( .A(n13416), .B(n13415), .Z(n13409) );
  OR U14182 ( .A(n13312), .B(n13310), .Z(n13316) );
  ANDN U14183 ( .B(n13312), .A(n13311), .Z(n13314) );
  OR U14184 ( .A(n13314), .B(n13313), .Z(n13315) );
  AND U14185 ( .A(n13316), .B(n13315), .Z(n13408) );
  NANDN U14186 ( .A(n13318), .B(n13317), .Z(n13322) );
  NAND U14187 ( .A(n13320), .B(n13319), .Z(n13321) );
  NAND U14188 ( .A(n13322), .B(n13321), .Z(n13407) );
  IV U14189 ( .A(n13407), .Z(n13406) );
  XOR U14190 ( .A(n13408), .B(n13406), .Z(n13323) );
  XNOR U14191 ( .A(n13409), .B(n13323), .Z(N304) );
  AND U14192 ( .A(x[232]), .B(y[1934]), .Z(n13682) );
  NAND U14193 ( .A(n13682), .B(n13324), .Z(n13328) );
  NAND U14194 ( .A(n13326), .B(n13325), .Z(n13327) );
  NAND U14195 ( .A(n13328), .B(n13327), .Z(n13446) );
  AND U14196 ( .A(x[239]), .B(y[1935]), .Z(n15360) );
  NAND U14197 ( .A(n15360), .B(n13329), .Z(n13333) );
  NAND U14198 ( .A(n13331), .B(n13330), .Z(n13332) );
  NAND U14199 ( .A(n13333), .B(n13332), .Z(n13445) );
  XOR U14200 ( .A(n13446), .B(n13445), .Z(n13448) );
  AND U14201 ( .A(x[234]), .B(y[1931]), .Z(n13335) );
  NAND U14202 ( .A(n13335), .B(n13334), .Z(n13339) );
  NAND U14203 ( .A(n13337), .B(n13336), .Z(n13338) );
  NAND U14204 ( .A(n13339), .B(n13338), .Z(n13483) );
  AND U14205 ( .A(x[224]), .B(y[1936]), .Z(n13505) );
  AND U14206 ( .A(x[240]), .B(y[1920]), .Z(n13506) );
  XOR U14207 ( .A(n13505), .B(n13506), .Z(n13508) );
  AND U14208 ( .A(x[239]), .B(y[1921]), .Z(n13493) );
  XOR U14209 ( .A(o[144]), .B(n13493), .Z(n13507) );
  XOR U14210 ( .A(n13508), .B(n13507), .Z(n13482) );
  NAND U14211 ( .A(y[1929]), .B(x[231]), .Z(n13340) );
  XNOR U14212 ( .A(n13341), .B(n13340), .Z(n13498) );
  AND U14213 ( .A(x[234]), .B(y[1926]), .Z(n13497) );
  XOR U14214 ( .A(n13498), .B(n13497), .Z(n13481) );
  XOR U14215 ( .A(n13482), .B(n13481), .Z(n13484) );
  XOR U14216 ( .A(n13483), .B(n13484), .Z(n13447) );
  XNOR U14217 ( .A(n13448), .B(n13447), .Z(n13478) );
  NANDN U14218 ( .A(n13342), .B(n13496), .Z(n13346) );
  NAND U14219 ( .A(n13344), .B(n13343), .Z(n13345) );
  NAND U14220 ( .A(n13346), .B(n13345), .Z(n13476) );
  AND U14221 ( .A(x[233]), .B(y[1933]), .Z(n14167) );
  NAND U14222 ( .A(n14167), .B(n13759), .Z(n13350) );
  NAND U14223 ( .A(n13348), .B(n13347), .Z(n13349) );
  AND U14224 ( .A(n13350), .B(n13349), .Z(n13516) );
  AND U14225 ( .A(y[1935]), .B(x[225]), .Z(n13352) );
  NAND U14226 ( .A(y[1928]), .B(x[232]), .Z(n13351) );
  XNOR U14227 ( .A(n13352), .B(n13351), .Z(n13502) );
  AND U14228 ( .A(o[143]), .B(n13353), .Z(n13501) );
  XOR U14229 ( .A(n13502), .B(n13501), .Z(n13514) );
  NAND U14230 ( .A(y[1922]), .B(x[238]), .Z(n13354) );
  XNOR U14231 ( .A(n13355), .B(n13354), .Z(n13457) );
  AND U14232 ( .A(x[228]), .B(y[1932]), .Z(n13458) );
  XOR U14233 ( .A(n13457), .B(n13458), .Z(n13513) );
  XOR U14234 ( .A(n13514), .B(n13513), .Z(n13515) );
  XOR U14235 ( .A(n13516), .B(n13515), .Z(n13475) );
  XOR U14236 ( .A(n13476), .B(n13475), .Z(n13477) );
  XOR U14237 ( .A(n13478), .B(n13477), .Z(n13439) );
  NAND U14238 ( .A(n13357), .B(n13356), .Z(n13361) );
  NAND U14239 ( .A(n13359), .B(n13358), .Z(n13360) );
  AND U14240 ( .A(n13361), .B(n13360), .Z(n13440) );
  XOR U14241 ( .A(n13439), .B(n13440), .Z(n13442) );
  NAND U14242 ( .A(n13363), .B(n13362), .Z(n13367) );
  NAND U14243 ( .A(n13365), .B(n13364), .Z(n13366) );
  NAND U14244 ( .A(n13367), .B(n13366), .Z(n13472) );
  AND U14245 ( .A(x[237]), .B(y[1924]), .Z(n13468) );
  NAND U14246 ( .A(n14028), .B(n13468), .Z(n13371) );
  NAND U14247 ( .A(n13369), .B(n13368), .Z(n13370) );
  NAND U14248 ( .A(n13371), .B(n13370), .Z(n13454) );
  AND U14249 ( .A(y[1934]), .B(x[226]), .Z(n13373) );
  NAND U14250 ( .A(y[1927]), .B(x[233]), .Z(n13372) );
  XNOR U14251 ( .A(n13373), .B(n13372), .Z(n13461) );
  AND U14252 ( .A(x[227]), .B(y[1933]), .Z(n13462) );
  XOR U14253 ( .A(n13461), .B(n13462), .Z(n13452) );
  AND U14254 ( .A(x[236]), .B(y[1924]), .Z(n14156) );
  AND U14255 ( .A(y[1931]), .B(x[229]), .Z(n13375) );
  NAND U14256 ( .A(y[1923]), .B(x[237]), .Z(n13374) );
  XNOR U14257 ( .A(n13375), .B(n13374), .Z(n13488) );
  XOR U14258 ( .A(n14156), .B(n13488), .Z(n13451) );
  XOR U14259 ( .A(n13452), .B(n13451), .Z(n13453) );
  XNOR U14260 ( .A(n13454), .B(n13453), .Z(n13469) );
  NAND U14261 ( .A(n13377), .B(n13376), .Z(n13381) );
  NAND U14262 ( .A(n13379), .B(n13378), .Z(n13380) );
  AND U14263 ( .A(n13381), .B(n13380), .Z(n13470) );
  XOR U14264 ( .A(n13469), .B(n13470), .Z(n13471) );
  XOR U14265 ( .A(n13472), .B(n13471), .Z(n13441) );
  XOR U14266 ( .A(n13442), .B(n13441), .Z(n13421) );
  NANDN U14267 ( .A(n13383), .B(n13382), .Z(n13387) );
  NANDN U14268 ( .A(n13385), .B(n13384), .Z(n13386) );
  AND U14269 ( .A(n13387), .B(n13386), .Z(n13420) );
  NAND U14270 ( .A(n13389), .B(n13388), .Z(n13393) );
  NAND U14271 ( .A(n13391), .B(n13390), .Z(n13392) );
  NAND U14272 ( .A(n13393), .B(n13392), .Z(n13435) );
  NAND U14273 ( .A(n13395), .B(n13394), .Z(n13399) );
  NANDN U14274 ( .A(n13397), .B(n13396), .Z(n13398) );
  NAND U14275 ( .A(n13399), .B(n13398), .Z(n13433) );
  NANDN U14276 ( .A(n13401), .B(n13400), .Z(n13405) );
  NAND U14277 ( .A(n13403), .B(n13402), .Z(n13404) );
  AND U14278 ( .A(n13405), .B(n13404), .Z(n13434) );
  XNOR U14279 ( .A(n13433), .B(n13434), .Z(n13436) );
  XNOR U14280 ( .A(n13422), .B(n13423), .Z(n13429) );
  OR U14281 ( .A(n13408), .B(n13406), .Z(n13412) );
  ANDN U14282 ( .B(n13408), .A(n13407), .Z(n13410) );
  OR U14283 ( .A(n13410), .B(n13409), .Z(n13411) );
  AND U14284 ( .A(n13412), .B(n13411), .Z(n13427) );
  NAND U14285 ( .A(n13414), .B(n13413), .Z(n13418) );
  NANDN U14286 ( .A(n13416), .B(n13415), .Z(n13417) );
  AND U14287 ( .A(n13418), .B(n13417), .Z(n13428) );
  IV U14288 ( .A(n13428), .Z(n13426) );
  XOR U14289 ( .A(n13427), .B(n13426), .Z(n13419) );
  XNOR U14290 ( .A(n13429), .B(n13419), .Z(N305) );
  NANDN U14291 ( .A(n13421), .B(n13420), .Z(n13425) );
  NANDN U14292 ( .A(n13423), .B(n13422), .Z(n13424) );
  AND U14293 ( .A(n13425), .B(n13424), .Z(n13526) );
  NANDN U14294 ( .A(n13426), .B(n13427), .Z(n13432) );
  NOR U14295 ( .A(n13428), .B(n13427), .Z(n13430) );
  OR U14296 ( .A(n13430), .B(n13429), .Z(n13431) );
  AND U14297 ( .A(n13432), .B(n13431), .Z(n13527) );
  NAND U14298 ( .A(n13434), .B(n13433), .Z(n13438) );
  NANDN U14299 ( .A(n13436), .B(n13435), .Z(n13437) );
  NAND U14300 ( .A(n13438), .B(n13437), .Z(n13522) );
  NAND U14301 ( .A(n13440), .B(n13439), .Z(n13444) );
  NAND U14302 ( .A(n13442), .B(n13441), .Z(n13443) );
  NAND U14303 ( .A(n13444), .B(n13443), .Z(n13532) );
  NAND U14304 ( .A(n13446), .B(n13445), .Z(n13450) );
  NAND U14305 ( .A(n13448), .B(n13447), .Z(n13449) );
  NAND U14306 ( .A(n13450), .B(n13449), .Z(n13614) );
  NAND U14307 ( .A(n13452), .B(n13451), .Z(n13456) );
  NAND U14308 ( .A(n13454), .B(n13453), .Z(n13455) );
  NAND U14309 ( .A(n13456), .B(n13455), .Z(n13612) );
  NAND U14310 ( .A(x[238]), .B(y[1925]), .Z(n13792) );
  NANDN U14311 ( .A(n13792), .B(n14028), .Z(n13460) );
  NAND U14312 ( .A(n13458), .B(n13457), .Z(n13459) );
  NAND U14313 ( .A(n13460), .B(n13459), .Z(n13606) );
  AND U14314 ( .A(x[233]), .B(y[1934]), .Z(n14412) );
  NANDN U14315 ( .A(n13592), .B(n14412), .Z(n13464) );
  NAND U14316 ( .A(n13462), .B(n13461), .Z(n13463) );
  NAND U14317 ( .A(n13464), .B(n13463), .Z(n13605) );
  XOR U14318 ( .A(n13606), .B(n13605), .Z(n13608) );
  AND U14319 ( .A(x[231]), .B(y[1930]), .Z(n13600) );
  AND U14320 ( .A(y[1932]), .B(x[229]), .Z(n13642) );
  NAND U14321 ( .A(y[1929]), .B(x[232]), .Z(n13465) );
  XNOR U14322 ( .A(n13642), .B(n13465), .Z(n13584) );
  XOR U14323 ( .A(n13584), .B(n13466), .Z(n13599) );
  XOR U14324 ( .A(n13600), .B(n13599), .Z(n13602) );
  NAND U14325 ( .A(y[1933]), .B(x[228]), .Z(n13467) );
  XNOR U14326 ( .A(n13468), .B(n13467), .Z(n13546) );
  AND U14327 ( .A(x[235]), .B(y[1926]), .Z(n13547) );
  XOR U14328 ( .A(n13546), .B(n13547), .Z(n13601) );
  XOR U14329 ( .A(n13602), .B(n13601), .Z(n13607) );
  XOR U14330 ( .A(n13608), .B(n13607), .Z(n13611) );
  XOR U14331 ( .A(n13612), .B(n13611), .Z(n13613) );
  XNOR U14332 ( .A(n13614), .B(n13613), .Z(n13530) );
  NAND U14333 ( .A(n13470), .B(n13469), .Z(n13474) );
  NAND U14334 ( .A(n13472), .B(n13471), .Z(n13473) );
  NAND U14335 ( .A(n13474), .B(n13473), .Z(n13529) );
  XOR U14336 ( .A(n13530), .B(n13529), .Z(n13531) );
  XOR U14337 ( .A(n13532), .B(n13531), .Z(n13521) );
  NAND U14338 ( .A(n13476), .B(n13475), .Z(n13480) );
  NAND U14339 ( .A(n13478), .B(n13477), .Z(n13479) );
  AND U14340 ( .A(n13480), .B(n13479), .Z(n13538) );
  NAND U14341 ( .A(n13482), .B(n13481), .Z(n13486) );
  NAND U14342 ( .A(n13484), .B(n13483), .Z(n13485) );
  NAND U14343 ( .A(n13486), .B(n13485), .Z(n13620) );
  AND U14344 ( .A(x[237]), .B(y[1931]), .Z(n14431) );
  NAND U14345 ( .A(n14431), .B(n13487), .Z(n13490) );
  NAND U14346 ( .A(n13488), .B(n14156), .Z(n13489) );
  NAND U14347 ( .A(n13490), .B(n13489), .Z(n13568) );
  AND U14348 ( .A(y[1936]), .B(x[225]), .Z(n13492) );
  NAND U14349 ( .A(y[1928]), .B(x[233]), .Z(n13491) );
  XNOR U14350 ( .A(n13492), .B(n13491), .Z(n13589) );
  AND U14351 ( .A(o[144]), .B(n13493), .Z(n13588) );
  XOR U14352 ( .A(n13589), .B(n13588), .Z(n13566) );
  AND U14353 ( .A(y[1922]), .B(x[239]), .Z(n13495) );
  NAND U14354 ( .A(y[1925]), .B(x[236]), .Z(n13494) );
  XNOR U14355 ( .A(n13495), .B(n13494), .Z(n13541) );
  AND U14356 ( .A(x[238]), .B(y[1923]), .Z(n13542) );
  XOR U14357 ( .A(n13541), .B(n13542), .Z(n13565) );
  XOR U14358 ( .A(n13566), .B(n13565), .Z(n13567) );
  XOR U14359 ( .A(n13568), .B(n13567), .Z(n13618) );
  NANDN U14360 ( .A(n13496), .B(n13600), .Z(n13500) );
  NAND U14361 ( .A(n13498), .B(n13497), .Z(n13499) );
  NAND U14362 ( .A(n13500), .B(n13499), .Z(n13578) );
  AND U14363 ( .A(x[232]), .B(y[1935]), .Z(n14151) );
  IV U14364 ( .A(n14151), .Z(n14237) );
  AND U14365 ( .A(x[225]), .B(y[1928]), .Z(n13660) );
  NANDN U14366 ( .A(n14237), .B(n13660), .Z(n13504) );
  NAND U14367 ( .A(n13502), .B(n13501), .Z(n13503) );
  NAND U14368 ( .A(n13504), .B(n13503), .Z(n13577) );
  XOR U14369 ( .A(n13578), .B(n13577), .Z(n13580) );
  NAND U14370 ( .A(n13506), .B(n13505), .Z(n13510) );
  NAND U14371 ( .A(n13508), .B(n13507), .Z(n13509) );
  NAND U14372 ( .A(n13510), .B(n13509), .Z(n13574) );
  AND U14373 ( .A(x[224]), .B(y[1937]), .Z(n13555) );
  AND U14374 ( .A(x[241]), .B(y[1920]), .Z(n13556) );
  XOR U14375 ( .A(n13555), .B(n13556), .Z(n13558) );
  AND U14376 ( .A(x[240]), .B(y[1921]), .Z(n13552) );
  XOR U14377 ( .A(o[145]), .B(n13552), .Z(n13557) );
  XOR U14378 ( .A(n13558), .B(n13557), .Z(n13572) );
  AND U14379 ( .A(y[1935]), .B(x[226]), .Z(n13512) );
  NAND U14380 ( .A(y[1927]), .B(x[234]), .Z(n13511) );
  XNOR U14381 ( .A(n13512), .B(n13511), .Z(n13593) );
  AND U14382 ( .A(x[227]), .B(y[1934]), .Z(n13594) );
  XOR U14383 ( .A(n13593), .B(n13594), .Z(n13571) );
  XOR U14384 ( .A(n13572), .B(n13571), .Z(n13573) );
  XOR U14385 ( .A(n13574), .B(n13573), .Z(n13579) );
  XOR U14386 ( .A(n13580), .B(n13579), .Z(n13617) );
  XOR U14387 ( .A(n13618), .B(n13617), .Z(n13619) );
  XNOR U14388 ( .A(n13620), .B(n13619), .Z(n13535) );
  NAND U14389 ( .A(n13514), .B(n13513), .Z(n13518) );
  NANDN U14390 ( .A(n13516), .B(n13515), .Z(n13517) );
  AND U14391 ( .A(n13518), .B(n13517), .Z(n13536) );
  XOR U14392 ( .A(n13535), .B(n13536), .Z(n13537) );
  XOR U14393 ( .A(n13538), .B(n13537), .Z(n13520) );
  XOR U14394 ( .A(n13522), .B(n13523), .Z(n13528) );
  XNOR U14395 ( .A(n13527), .B(n13528), .Z(n13519) );
  XOR U14396 ( .A(n13526), .B(n13519), .Z(N306) );
  NANDN U14397 ( .A(n13521), .B(n13520), .Z(n13525) );
  NAND U14398 ( .A(n13523), .B(n13522), .Z(n13524) );
  AND U14399 ( .A(n13525), .B(n13524), .Z(n13732) );
  NAND U14400 ( .A(n13530), .B(n13529), .Z(n13534) );
  NAND U14401 ( .A(n13532), .B(n13531), .Z(n13533) );
  AND U14402 ( .A(n13534), .B(n13533), .Z(n13729) );
  NAND U14403 ( .A(n13536), .B(n13535), .Z(n13540) );
  NANDN U14404 ( .A(n13538), .B(n13537), .Z(n13539) );
  AND U14405 ( .A(n13540), .B(n13539), .Z(n13727) );
  AND U14406 ( .A(x[236]), .B(y[1922]), .Z(n13864) );
  AND U14407 ( .A(x[239]), .B(y[1925]), .Z(n13767) );
  NAND U14408 ( .A(n13864), .B(n13767), .Z(n13544) );
  NAND U14409 ( .A(n13542), .B(n13541), .Z(n13543) );
  AND U14410 ( .A(n13544), .B(n13543), .Z(n13709) );
  NAND U14411 ( .A(n14719), .B(n13545), .Z(n13549) );
  NAND U14412 ( .A(n13547), .B(n13546), .Z(n13548) );
  NAND U14413 ( .A(n13549), .B(n13548), .Z(n13699) );
  AND U14414 ( .A(y[1937]), .B(x[225]), .Z(n13551) );
  NAND U14415 ( .A(y[1928]), .B(x[234]), .Z(n13550) );
  XNOR U14416 ( .A(n13551), .B(n13550), .Z(n13662) );
  AND U14417 ( .A(o[145]), .B(n13552), .Z(n13661) );
  XOR U14418 ( .A(n13662), .B(n13661), .Z(n13697) );
  AND U14419 ( .A(y[1923]), .B(x[239]), .Z(n13554) );
  NAND U14420 ( .A(y[1929]), .B(x[233]), .Z(n13553) );
  XNOR U14421 ( .A(n13554), .B(n13553), .Z(n13652) );
  AND U14422 ( .A(x[238]), .B(y[1924]), .Z(n13653) );
  XOR U14423 ( .A(n13652), .B(n13653), .Z(n13696) );
  XOR U14424 ( .A(n13697), .B(n13696), .Z(n13698) );
  XOR U14425 ( .A(n13699), .B(n13698), .Z(n13708) );
  NAND U14426 ( .A(n13556), .B(n13555), .Z(n13560) );
  NAND U14427 ( .A(n13558), .B(n13557), .Z(n13559) );
  AND U14428 ( .A(n13560), .B(n13559), .Z(n13721) );
  AND U14429 ( .A(y[1922]), .B(x[240]), .Z(n13562) );
  NAND U14430 ( .A(y[1927]), .B(x[235]), .Z(n13561) );
  XNOR U14431 ( .A(n13562), .B(n13561), .Z(n13648) );
  AND U14432 ( .A(x[226]), .B(y[1936]), .Z(n13649) );
  XOR U14433 ( .A(n13648), .B(n13649), .Z(n13720) );
  AND U14434 ( .A(y[1933]), .B(x[229]), .Z(n13776) );
  NAND U14435 ( .A(y[1932]), .B(x[230]), .Z(n13563) );
  XNOR U14436 ( .A(n13776), .B(n13563), .Z(n13645) );
  NAND U14437 ( .A(y[1934]), .B(x[228]), .Z(n13564) );
  XNOR U14438 ( .A(n14417), .B(n13564), .Z(n13684) );
  AND U14439 ( .A(x[231]), .B(y[1931]), .Z(n13683) );
  XOR U14440 ( .A(n13684), .B(n13683), .Z(n13644) );
  XOR U14441 ( .A(n13645), .B(n13644), .Z(n13722) );
  XOR U14442 ( .A(n13723), .B(n13722), .Z(n13710) );
  XNOR U14443 ( .A(n13711), .B(n13710), .Z(n13631) );
  NAND U14444 ( .A(n13566), .B(n13565), .Z(n13570) );
  NAND U14445 ( .A(n13568), .B(n13567), .Z(n13569) );
  AND U14446 ( .A(n13570), .B(n13569), .Z(n13702) );
  NAND U14447 ( .A(n13572), .B(n13571), .Z(n13576) );
  NAND U14448 ( .A(n13574), .B(n13573), .Z(n13575) );
  NAND U14449 ( .A(n13576), .B(n13575), .Z(n13703) );
  NAND U14450 ( .A(n13578), .B(n13577), .Z(n13582) );
  NAND U14451 ( .A(n13580), .B(n13579), .Z(n13581) );
  NAND U14452 ( .A(n13582), .B(n13581), .Z(n13705) );
  XOR U14453 ( .A(n13631), .B(n13630), .Z(n13633) );
  AND U14454 ( .A(x[232]), .B(y[1932]), .Z(n13901) );
  NAND U14455 ( .A(n13901), .B(n13583), .Z(n13587) );
  NANDN U14456 ( .A(n13585), .B(n13584), .Z(n13586) );
  NAND U14457 ( .A(n13587), .B(n13586), .Z(n13715) );
  NAND U14458 ( .A(x[233]), .B(y[1936]), .Z(n14491) );
  NANDN U14459 ( .A(n14491), .B(n13660), .Z(n13591) );
  NAND U14460 ( .A(n13589), .B(n13588), .Z(n13590) );
  NAND U14461 ( .A(n13591), .B(n13590), .Z(n13714) );
  XOR U14462 ( .A(n13715), .B(n13714), .Z(n13717) );
  NAND U14463 ( .A(x[234]), .B(y[1935]), .Z(n14492) );
  OR U14464 ( .A(n14492), .B(n13592), .Z(n13596) );
  NAND U14465 ( .A(n13594), .B(n13593), .Z(n13595) );
  NAND U14466 ( .A(n13596), .B(n13595), .Z(n13693) );
  AND U14467 ( .A(x[224]), .B(y[1938]), .Z(n13665) );
  AND U14468 ( .A(x[242]), .B(y[1920]), .Z(n13666) );
  XOR U14469 ( .A(n13665), .B(n13666), .Z(n13667) );
  NAND U14470 ( .A(x[241]), .B(y[1921]), .Z(n13687) );
  XNOR U14471 ( .A(o[146]), .B(n13687), .Z(n13668) );
  XOR U14472 ( .A(n13667), .B(n13668), .Z(n13691) );
  AND U14473 ( .A(y[1925]), .B(x[237]), .Z(n13598) );
  NAND U14474 ( .A(y[1935]), .B(x[227]), .Z(n13597) );
  XNOR U14475 ( .A(n13598), .B(n13597), .Z(n13673) );
  AND U14476 ( .A(x[236]), .B(y[1926]), .Z(n13674) );
  XOR U14477 ( .A(n13673), .B(n13674), .Z(n13690) );
  XOR U14478 ( .A(n13691), .B(n13690), .Z(n13692) );
  XOR U14479 ( .A(n13693), .B(n13692), .Z(n13716) );
  XNOR U14480 ( .A(n13717), .B(n13716), .Z(n13637) );
  NAND U14481 ( .A(n13600), .B(n13599), .Z(n13604) );
  NAND U14482 ( .A(n13602), .B(n13601), .Z(n13603) );
  AND U14483 ( .A(n13604), .B(n13603), .Z(n13636) );
  XOR U14484 ( .A(n13637), .B(n13636), .Z(n13638) );
  NAND U14485 ( .A(n13606), .B(n13605), .Z(n13610) );
  NAND U14486 ( .A(n13608), .B(n13607), .Z(n13609) );
  AND U14487 ( .A(n13610), .B(n13609), .Z(n13639) );
  XOR U14488 ( .A(n13638), .B(n13639), .Z(n13632) );
  XNOR U14489 ( .A(n13633), .B(n13632), .Z(n13627) );
  NAND U14490 ( .A(n13612), .B(n13611), .Z(n13616) );
  NAND U14491 ( .A(n13614), .B(n13613), .Z(n13615) );
  NAND U14492 ( .A(n13616), .B(n13615), .Z(n13625) );
  NAND U14493 ( .A(n13618), .B(n13617), .Z(n13622) );
  NAND U14494 ( .A(n13620), .B(n13619), .Z(n13621) );
  NAND U14495 ( .A(n13622), .B(n13621), .Z(n13624) );
  XOR U14496 ( .A(n13625), .B(n13624), .Z(n13626) );
  XOR U14497 ( .A(n13627), .B(n13626), .Z(n13726) );
  XOR U14498 ( .A(n13727), .B(n13726), .Z(n13728) );
  XOR U14499 ( .A(n13729), .B(n13728), .Z(n13734) );
  XNOR U14500 ( .A(n13733), .B(n13734), .Z(n13623) );
  XOR U14501 ( .A(n13732), .B(n13623), .Z(N307) );
  NAND U14502 ( .A(n13625), .B(n13624), .Z(n13629) );
  NAND U14503 ( .A(n13627), .B(n13626), .Z(n13628) );
  AND U14504 ( .A(n13629), .B(n13628), .Z(n13848) );
  NAND U14505 ( .A(n13631), .B(n13630), .Z(n13635) );
  NAND U14506 ( .A(n13633), .B(n13632), .Z(n13634) );
  AND U14507 ( .A(n13635), .B(n13634), .Z(n13846) );
  NAND U14508 ( .A(n13637), .B(n13636), .Z(n13641) );
  NAND U14509 ( .A(n13639), .B(n13638), .Z(n13640) );
  NAND U14510 ( .A(n13641), .B(n13640), .Z(n13739) );
  AND U14511 ( .A(x[230]), .B(y[1933]), .Z(n13643) );
  NAND U14512 ( .A(n13643), .B(n13642), .Z(n13647) );
  NAND U14513 ( .A(n13645), .B(n13644), .Z(n13646) );
  NAND U14514 ( .A(n13647), .B(n13646), .Z(n13821) );
  AND U14515 ( .A(x[240]), .B(y[1927]), .Z(n14172) );
  NAND U14516 ( .A(n14172), .B(n14028), .Z(n13651) );
  NAND U14517 ( .A(n13649), .B(n13648), .Z(n13650) );
  NAND U14518 ( .A(n13651), .B(n13650), .Z(n13819) );
  AND U14519 ( .A(x[239]), .B(y[1929]), .Z(n14401) );
  NAND U14520 ( .A(n14401), .B(n13754), .Z(n13655) );
  NAND U14521 ( .A(n13653), .B(n13652), .Z(n13654) );
  NAND U14522 ( .A(n13655), .B(n13654), .Z(n13744) );
  AND U14523 ( .A(y[1938]), .B(x[225]), .Z(n13657) );
  NAND U14524 ( .A(y[1931]), .B(x[232]), .Z(n13656) );
  XNOR U14525 ( .A(n13657), .B(n13656), .Z(n13791) );
  XNOR U14526 ( .A(n13791), .B(n13792), .Z(n13743) );
  AND U14527 ( .A(y[1926]), .B(x[237]), .Z(n13659) );
  NAND U14528 ( .A(y[1937]), .B(x[226]), .Z(n13658) );
  XNOR U14529 ( .A(n13659), .B(n13658), .Z(n13761) );
  XOR U14530 ( .A(n13761), .B(n13760), .Z(n13742) );
  XOR U14531 ( .A(n13743), .B(n13742), .Z(n13745) );
  XOR U14532 ( .A(n13744), .B(n13745), .Z(n13818) );
  XOR U14533 ( .A(n13819), .B(n13818), .Z(n13820) );
  XNOR U14534 ( .A(n13821), .B(n13820), .Z(n13737) );
  AND U14535 ( .A(x[234]), .B(y[1937]), .Z(n14809) );
  IV U14536 ( .A(n14809), .Z(n14672) );
  NANDN U14537 ( .A(n14672), .B(n13660), .Z(n13664) );
  NAND U14538 ( .A(n13662), .B(n13661), .Z(n13663) );
  NAND U14539 ( .A(n13664), .B(n13663), .Z(n13802) );
  NAND U14540 ( .A(n13666), .B(n13665), .Z(n13670) );
  NAND U14541 ( .A(n13668), .B(n13667), .Z(n13669) );
  NAND U14542 ( .A(n13670), .B(n13669), .Z(n13800) );
  AND U14543 ( .A(y[1923]), .B(x[240]), .Z(n14371) );
  NAND U14544 ( .A(y[1930]), .B(x[233]), .Z(n13671) );
  XNOR U14545 ( .A(n14371), .B(n13671), .Z(n13756) );
  AND U14546 ( .A(x[239]), .B(y[1924]), .Z(n13755) );
  XOR U14547 ( .A(n13756), .B(n13755), .Z(n13801) );
  XOR U14548 ( .A(n13800), .B(n13801), .Z(n13803) );
  XNOR U14549 ( .A(n13802), .B(n13803), .Z(n13814) );
  AND U14550 ( .A(x[237]), .B(y[1935]), .Z(n15017) );
  NANDN U14551 ( .A(n13672), .B(n15017), .Z(n13676) );
  NAND U14552 ( .A(n13674), .B(n13673), .Z(n13675) );
  NAND U14553 ( .A(n13676), .B(n13675), .Z(n13808) );
  AND U14554 ( .A(y[1929]), .B(x[234]), .Z(n13678) );
  NAND U14555 ( .A(y[1922]), .B(x[241]), .Z(n13677) );
  XNOR U14556 ( .A(n13678), .B(n13677), .Z(n13796) );
  NAND U14557 ( .A(x[242]), .B(y[1921]), .Z(n13775) );
  XOR U14558 ( .A(o[147]), .B(n13775), .Z(n13797) );
  XNOR U14559 ( .A(n13796), .B(n13797), .Z(n13807) );
  NAND U14560 ( .A(y[1936]), .B(x[227]), .Z(n13679) );
  XNOR U14561 ( .A(n13680), .B(n13679), .Z(n13769) );
  XNOR U14562 ( .A(n13769), .B(n13770), .Z(n13806) );
  XOR U14563 ( .A(n13807), .B(n13806), .Z(n13809) );
  XNOR U14564 ( .A(n13808), .B(n13809), .Z(n13813) );
  NAND U14565 ( .A(n13682), .B(n13681), .Z(n13686) );
  NAND U14566 ( .A(n13684), .B(n13683), .Z(n13685) );
  NAND U14567 ( .A(n13686), .B(n13685), .Z(n13750) );
  AND U14568 ( .A(x[224]), .B(y[1939]), .Z(n13780) );
  NAND U14569 ( .A(x[243]), .B(y[1920]), .Z(n13781) );
  XNOR U14570 ( .A(n13780), .B(n13781), .Z(n13783) );
  ANDN U14571 ( .B(o[146]), .A(n13687), .Z(n13782) );
  XOR U14572 ( .A(n13783), .B(n13782), .Z(n13749) );
  AND U14573 ( .A(x[228]), .B(y[1935]), .Z(n13915) );
  AND U14574 ( .A(y[1934]), .B(x[229]), .Z(n13689) );
  NAND U14575 ( .A(y[1933]), .B(x[230]), .Z(n13688) );
  XOR U14576 ( .A(n13689), .B(n13688), .Z(n13777) );
  XNOR U14577 ( .A(n13915), .B(n13777), .Z(n13748) );
  XOR U14578 ( .A(n13749), .B(n13748), .Z(n13751) );
  XNOR U14579 ( .A(n13750), .B(n13751), .Z(n13812) );
  XOR U14580 ( .A(n13813), .B(n13812), .Z(n13815) );
  XNOR U14581 ( .A(n13814), .B(n13815), .Z(n13826) );
  NAND U14582 ( .A(n13691), .B(n13690), .Z(n13695) );
  NAND U14583 ( .A(n13693), .B(n13692), .Z(n13694) );
  NAND U14584 ( .A(n13695), .B(n13694), .Z(n13825) );
  NAND U14585 ( .A(n13697), .B(n13696), .Z(n13701) );
  NAND U14586 ( .A(n13699), .B(n13698), .Z(n13700) );
  NAND U14587 ( .A(n13701), .B(n13700), .Z(n13824) );
  XOR U14588 ( .A(n13825), .B(n13824), .Z(n13827) );
  XNOR U14589 ( .A(n13826), .B(n13827), .Z(n13736) );
  XOR U14590 ( .A(n13737), .B(n13736), .Z(n13738) );
  XNOR U14591 ( .A(n13739), .B(n13738), .Z(n13838) );
  NANDN U14592 ( .A(n13703), .B(n13702), .Z(n13707) );
  NANDN U14593 ( .A(n13705), .B(n13704), .Z(n13706) );
  AND U14594 ( .A(n13707), .B(n13706), .Z(n13837) );
  NANDN U14595 ( .A(n13709), .B(n13708), .Z(n13713) );
  NAND U14596 ( .A(n13711), .B(n13710), .Z(n13712) );
  AND U14597 ( .A(n13713), .B(n13712), .Z(n13833) );
  NAND U14598 ( .A(n13715), .B(n13714), .Z(n13719) );
  NAND U14599 ( .A(n13717), .B(n13716), .Z(n13718) );
  AND U14600 ( .A(n13719), .B(n13718), .Z(n13831) );
  NANDN U14601 ( .A(n13721), .B(n13720), .Z(n13725) );
  NAND U14602 ( .A(n13723), .B(n13722), .Z(n13724) );
  NAND U14603 ( .A(n13725), .B(n13724), .Z(n13830) );
  XOR U14604 ( .A(n13837), .B(n13836), .Z(n13839) );
  XOR U14605 ( .A(n13838), .B(n13839), .Z(n13845) );
  XOR U14606 ( .A(n13846), .B(n13845), .Z(n13847) );
  XOR U14607 ( .A(n13848), .B(n13847), .Z(n13844) );
  NAND U14608 ( .A(n13727), .B(n13726), .Z(n13731) );
  NAND U14609 ( .A(n13729), .B(n13728), .Z(n13730) );
  NAND U14610 ( .A(n13731), .B(n13730), .Z(n13843) );
  XOR U14611 ( .A(n13843), .B(n13842), .Z(n13735) );
  XNOR U14612 ( .A(n13844), .B(n13735), .Z(N308) );
  NAND U14613 ( .A(n13737), .B(n13736), .Z(n13741) );
  NAND U14614 ( .A(n13739), .B(n13738), .Z(n13740) );
  AND U14615 ( .A(n13741), .B(n13740), .Z(n13949) );
  NAND U14616 ( .A(n13743), .B(n13742), .Z(n13747) );
  NAND U14617 ( .A(n13745), .B(n13744), .Z(n13746) );
  NAND U14618 ( .A(n13747), .B(n13746), .Z(n13853) );
  NAND U14619 ( .A(n13749), .B(n13748), .Z(n13753) );
  NAND U14620 ( .A(n13751), .B(n13750), .Z(n13752) );
  NAND U14621 ( .A(n13753), .B(n13752), .Z(n13852) );
  XOR U14622 ( .A(n13853), .B(n13852), .Z(n13855) );
  AND U14623 ( .A(x[240]), .B(y[1930]), .Z(n14630) );
  NAND U14624 ( .A(n14630), .B(n13754), .Z(n13758) );
  NAND U14625 ( .A(n13756), .B(n13755), .Z(n13757) );
  AND U14626 ( .A(n13758), .B(n13757), .Z(n13890) );
  AND U14627 ( .A(x[237]), .B(y[1937]), .Z(n15264) );
  NAND U14628 ( .A(n15264), .B(n13759), .Z(n13763) );
  NAND U14629 ( .A(n13761), .B(n13760), .Z(n13762) );
  AND U14630 ( .A(n13763), .B(n13762), .Z(n13933) );
  AND U14631 ( .A(y[1924]), .B(x[240]), .Z(n13765) );
  NAND U14632 ( .A(y[1930]), .B(x[234]), .Z(n13764) );
  XNOR U14633 ( .A(n13765), .B(n13764), .Z(n13896) );
  NAND U14634 ( .A(x[226]), .B(y[1938]), .Z(n13897) );
  XNOR U14635 ( .A(n13896), .B(n13897), .Z(n13930) );
  NAND U14636 ( .A(y[1931]), .B(x[233]), .Z(n13766) );
  XNOR U14637 ( .A(n13767), .B(n13766), .Z(n13872) );
  NAND U14638 ( .A(x[238]), .B(y[1926]), .Z(n13873) );
  XOR U14639 ( .A(n13872), .B(n13873), .Z(n13931) );
  XNOR U14640 ( .A(n13930), .B(n13931), .Z(n13932) );
  XNOR U14641 ( .A(n13933), .B(n13932), .Z(n13889) );
  XNOR U14642 ( .A(n13890), .B(n13889), .Z(n13892) );
  NAND U14643 ( .A(x[235]), .B(y[1936]), .Z(n14810) );
  NANDN U14644 ( .A(n14810), .B(n13768), .Z(n13772) );
  NANDN U14645 ( .A(n13770), .B(n13769), .Z(n13771) );
  AND U14646 ( .A(n13772), .B(n13771), .Z(n13939) );
  AND U14647 ( .A(y[1929]), .B(x[235]), .Z(n13774) );
  NAND U14648 ( .A(y[1939]), .B(x[225]), .Z(n13773) );
  XNOR U14649 ( .A(n13774), .B(n13773), .Z(n13870) );
  AND U14650 ( .A(x[243]), .B(y[1921]), .Z(n13876) );
  XOR U14651 ( .A(o[148]), .B(n13876), .Z(n13869) );
  XOR U14652 ( .A(n13870), .B(n13869), .Z(n13937) );
  AND U14653 ( .A(x[224]), .B(y[1940]), .Z(n13920) );
  NAND U14654 ( .A(x[244]), .B(y[1920]), .Z(n13921) );
  XNOR U14655 ( .A(n13920), .B(n13921), .Z(n13923) );
  ANDN U14656 ( .B(o[147]), .A(n13775), .Z(n13922) );
  XOR U14657 ( .A(n13923), .B(n13922), .Z(n13936) );
  XOR U14658 ( .A(n13937), .B(n13936), .Z(n13938) );
  XNOR U14659 ( .A(n13939), .B(n13938), .Z(n13891) );
  XOR U14660 ( .A(n13892), .B(n13891), .Z(n13854) );
  XNOR U14661 ( .A(n13855), .B(n13854), .Z(n13943) );
  AND U14662 ( .A(x[230]), .B(y[1934]), .Z(n13859) );
  NAND U14663 ( .A(n13859), .B(n13776), .Z(n13779) );
  NANDN U14664 ( .A(n13777), .B(n13915), .Z(n13778) );
  AND U14665 ( .A(n13779), .B(n13778), .Z(n13880) );
  AND U14666 ( .A(y[1922]), .B(x[242]), .Z(n13785) );
  NAND U14667 ( .A(y[1928]), .B(x[236]), .Z(n13784) );
  XNOR U14668 ( .A(n13785), .B(n13784), .Z(n13865) );
  NAND U14669 ( .A(x[241]), .B(y[1923]), .Z(n13866) );
  XNOR U14670 ( .A(n13865), .B(n13866), .Z(n13877) );
  XNOR U14671 ( .A(n13878), .B(n13877), .Z(n13879) );
  XOR U14672 ( .A(n13880), .B(n13879), .Z(n13884) );
  AND U14673 ( .A(y[1927]), .B(x[237]), .Z(n13787) );
  NAND U14674 ( .A(y[1937]), .B(x[227]), .Z(n13786) );
  XNOR U14675 ( .A(n13787), .B(n13786), .Z(n13902) );
  XOR U14676 ( .A(n13902), .B(n13901), .Z(n13860) );
  AND U14677 ( .A(y[1935]), .B(x[229]), .Z(n13789) );
  NAND U14678 ( .A(y[1936]), .B(x[228]), .Z(n13788) );
  XNOR U14679 ( .A(n13789), .B(n13788), .Z(n13917) );
  AND U14680 ( .A(x[231]), .B(y[1933]), .Z(n13916) );
  XNOR U14681 ( .A(n13917), .B(n13916), .Z(n13858) );
  XOR U14682 ( .A(n13859), .B(n13858), .Z(n13861) );
  XOR U14683 ( .A(n13860), .B(n13861), .Z(n13926) );
  AND U14684 ( .A(x[232]), .B(y[1938]), .Z(n14975) );
  AND U14685 ( .A(x[225]), .B(y[1931]), .Z(n13790) );
  NAND U14686 ( .A(n14975), .B(n13790), .Z(n13794) );
  NANDN U14687 ( .A(n13792), .B(n13791), .Z(n13793) );
  AND U14688 ( .A(n13794), .B(n13793), .Z(n13925) );
  AND U14689 ( .A(x[241]), .B(y[1929]), .Z(n14638) );
  NAND U14690 ( .A(n14638), .B(n13795), .Z(n13799) );
  NANDN U14691 ( .A(n13797), .B(n13796), .Z(n13798) );
  NAND U14692 ( .A(n13799), .B(n13798), .Z(n13924) );
  XOR U14693 ( .A(n13925), .B(n13924), .Z(n13927) );
  XNOR U14694 ( .A(n13926), .B(n13927), .Z(n13883) );
  XOR U14695 ( .A(n13884), .B(n13883), .Z(n13886) );
  NAND U14696 ( .A(n13801), .B(n13800), .Z(n13805) );
  NAND U14697 ( .A(n13803), .B(n13802), .Z(n13804) );
  AND U14698 ( .A(n13805), .B(n13804), .Z(n13885) );
  XOR U14699 ( .A(n13886), .B(n13885), .Z(n13941) );
  NAND U14700 ( .A(n13807), .B(n13806), .Z(n13811) );
  NAND U14701 ( .A(n13809), .B(n13808), .Z(n13810) );
  AND U14702 ( .A(n13811), .B(n13810), .Z(n13940) );
  XOR U14703 ( .A(n13941), .B(n13940), .Z(n13942) );
  XNOR U14704 ( .A(n13943), .B(n13942), .Z(n13947) );
  NAND U14705 ( .A(n13813), .B(n13812), .Z(n13817) );
  NAND U14706 ( .A(n13815), .B(n13814), .Z(n13816) );
  AND U14707 ( .A(n13817), .B(n13816), .Z(n13953) );
  NAND U14708 ( .A(n13819), .B(n13818), .Z(n13823) );
  NAND U14709 ( .A(n13821), .B(n13820), .Z(n13822) );
  AND U14710 ( .A(n13823), .B(n13822), .Z(n13952) );
  NAND U14711 ( .A(n13825), .B(n13824), .Z(n13829) );
  NAND U14712 ( .A(n13827), .B(n13826), .Z(n13828) );
  AND U14713 ( .A(n13829), .B(n13828), .Z(n13954) );
  XNOR U14714 ( .A(n13955), .B(n13954), .Z(n13946) );
  XOR U14715 ( .A(n13947), .B(n13946), .Z(n13948) );
  XOR U14716 ( .A(n13949), .B(n13948), .Z(n13961) );
  NANDN U14717 ( .A(n13831), .B(n13830), .Z(n13835) );
  NANDN U14718 ( .A(n13833), .B(n13832), .Z(n13834) );
  AND U14719 ( .A(n13835), .B(n13834), .Z(n13958) );
  NAND U14720 ( .A(n13837), .B(n13836), .Z(n13841) );
  NAND U14721 ( .A(n13839), .B(n13838), .Z(n13840) );
  NAND U14722 ( .A(n13841), .B(n13840), .Z(n13959) );
  XOR U14723 ( .A(n13961), .B(n13960), .Z(n13967) );
  NAND U14724 ( .A(n13846), .B(n13845), .Z(n13850) );
  NANDN U14725 ( .A(n13848), .B(n13847), .Z(n13849) );
  AND U14726 ( .A(n13850), .B(n13849), .Z(n13966) );
  IV U14727 ( .A(n13966), .Z(n13964) );
  XOR U14728 ( .A(n13965), .B(n13964), .Z(n13851) );
  XNOR U14729 ( .A(n13967), .B(n13851), .Z(N309) );
  NAND U14730 ( .A(n13853), .B(n13852), .Z(n13857) );
  NAND U14731 ( .A(n13855), .B(n13854), .Z(n13856) );
  NAND U14732 ( .A(n13857), .B(n13856), .Z(n13980) );
  NANDN U14733 ( .A(n13859), .B(n13858), .Z(n13863) );
  OR U14734 ( .A(n13861), .B(n13860), .Z(n13862) );
  AND U14735 ( .A(n13863), .B(n13862), .Z(n14068) );
  AND U14736 ( .A(x[242]), .B(y[1928]), .Z(n14637) );
  NAND U14737 ( .A(n14637), .B(n13864), .Z(n13868) );
  NANDN U14738 ( .A(n13866), .B(n13865), .Z(n13867) );
  AND U14739 ( .A(n13868), .B(n13867), .Z(n14052) );
  AND U14740 ( .A(x[235]), .B(y[1939]), .Z(n15313) );
  XNOR U14741 ( .A(n14052), .B(n14051), .Z(n14054) );
  AND U14742 ( .A(x[239]), .B(y[1931]), .Z(n14625) );
  NAND U14743 ( .A(n14625), .B(n13871), .Z(n13875) );
  NANDN U14744 ( .A(n13873), .B(n13872), .Z(n13874) );
  NAND U14745 ( .A(n13875), .B(n13874), .Z(n13992) );
  AND U14746 ( .A(x[224]), .B(y[1941]), .Z(n14012) );
  AND U14747 ( .A(x[245]), .B(y[1920]), .Z(n14013) );
  XOR U14748 ( .A(n14012), .B(n14013), .Z(n14015) );
  AND U14749 ( .A(o[148]), .B(n13876), .Z(n14014) );
  XOR U14750 ( .A(n14015), .B(n14014), .Z(n13991) );
  AND U14751 ( .A(x[229]), .B(y[1936]), .Z(n13997) );
  AND U14752 ( .A(x[240]), .B(y[1925]), .Z(n13996) );
  XOR U14753 ( .A(n13997), .B(n13996), .Z(n13999) );
  AND U14754 ( .A(x[239]), .B(y[1926]), .Z(n13998) );
  XOR U14755 ( .A(n13999), .B(n13998), .Z(n13990) );
  XOR U14756 ( .A(n13991), .B(n13990), .Z(n13993) );
  XOR U14757 ( .A(n13992), .B(n13993), .Z(n14053) );
  XNOR U14758 ( .A(n14054), .B(n14053), .Z(n14067) );
  XNOR U14759 ( .A(n14068), .B(n14067), .Z(n14069) );
  NANDN U14760 ( .A(n13878), .B(n13877), .Z(n13882) );
  NANDN U14761 ( .A(n13880), .B(n13879), .Z(n13881) );
  NAND U14762 ( .A(n13882), .B(n13881), .Z(n14070) );
  XOR U14763 ( .A(n14069), .B(n14070), .Z(n13978) );
  NAND U14764 ( .A(n13884), .B(n13883), .Z(n13888) );
  NAND U14765 ( .A(n13886), .B(n13885), .Z(n13887) );
  AND U14766 ( .A(n13888), .B(n13887), .Z(n13979) );
  XOR U14767 ( .A(n13978), .B(n13979), .Z(n13981) );
  XNOR U14768 ( .A(n13980), .B(n13981), .Z(n13974) );
  NANDN U14769 ( .A(n13890), .B(n13889), .Z(n13894) );
  NAND U14770 ( .A(n13892), .B(n13891), .Z(n13893) );
  AND U14771 ( .A(n13894), .B(n13893), .Z(n14076) );
  AND U14772 ( .A(x[234]), .B(y[1924]), .Z(n13895) );
  NAND U14773 ( .A(n14630), .B(n13895), .Z(n13899) );
  NANDN U14774 ( .A(n13897), .B(n13896), .Z(n13898) );
  AND U14775 ( .A(n13899), .B(n13898), .Z(n14046) );
  NAND U14776 ( .A(n15264), .B(n13900), .Z(n13904) );
  NAND U14777 ( .A(n13902), .B(n13901), .Z(n13903) );
  AND U14778 ( .A(n13904), .B(n13903), .Z(n14066) );
  AND U14779 ( .A(y[1922]), .B(x[243]), .Z(n13906) );
  NAND U14780 ( .A(y[1930]), .B(x[235]), .Z(n13905) );
  XNOR U14781 ( .A(n13906), .B(n13905), .Z(n14030) );
  AND U14782 ( .A(x[244]), .B(y[1921]), .Z(n14011) );
  XOR U14783 ( .A(n14011), .B(o[149]), .Z(n14029) );
  XOR U14784 ( .A(n14030), .B(n14029), .Z(n14064) );
  AND U14785 ( .A(y[1923]), .B(x[242]), .Z(n13908) );
  NAND U14786 ( .A(y[1931]), .B(x[234]), .Z(n13907) );
  XNOR U14787 ( .A(n13908), .B(n13907), .Z(n14019) );
  AND U14788 ( .A(x[225]), .B(y[1940]), .Z(n14020) );
  XOR U14789 ( .A(n14019), .B(n14020), .Z(n14063) );
  XOR U14790 ( .A(n14064), .B(n14063), .Z(n14065) );
  XNOR U14791 ( .A(n14066), .B(n14065), .Z(n14045) );
  XNOR U14792 ( .A(n14046), .B(n14045), .Z(n14047) );
  AND U14793 ( .A(x[231]), .B(y[1934]), .Z(n14235) );
  AND U14794 ( .A(y[1935]), .B(x[230]), .Z(n13910) );
  NAND U14795 ( .A(y[1927]), .B(x[238]), .Z(n13909) );
  XNOR U14796 ( .A(n13910), .B(n13909), .Z(n14023) );
  XOR U14797 ( .A(n14235), .B(n14023), .Z(n14042) );
  NAND U14798 ( .A(x[233]), .B(y[1932]), .Z(n14040) );
  NAND U14799 ( .A(x[232]), .B(y[1933]), .Z(n14039) );
  XOR U14800 ( .A(n14040), .B(n14039), .Z(n14041) );
  AND U14801 ( .A(y[1929]), .B(x[236]), .Z(n13912) );
  NAND U14802 ( .A(y[1924]), .B(x[241]), .Z(n13911) );
  XNOR U14803 ( .A(n13912), .B(n13911), .Z(n14033) );
  AND U14804 ( .A(x[226]), .B(y[1939]), .Z(n14034) );
  XOR U14805 ( .A(n14033), .B(n14034), .Z(n13985) );
  AND U14806 ( .A(y[1928]), .B(x[237]), .Z(n13914) );
  NAND U14807 ( .A(y[1938]), .B(x[227]), .Z(n13913) );
  XNOR U14808 ( .A(n13914), .B(n13913), .Z(n14008) );
  AND U14809 ( .A(x[228]), .B(y[1937]), .Z(n14007) );
  XOR U14810 ( .A(n14008), .B(n14007), .Z(n13984) );
  XOR U14811 ( .A(n13985), .B(n13984), .Z(n13986) );
  NAND U14812 ( .A(n13997), .B(n13915), .Z(n13919) );
  NAND U14813 ( .A(n13917), .B(n13916), .Z(n13918) );
  AND U14814 ( .A(n13919), .B(n13918), .Z(n14058) );
  XOR U14815 ( .A(n14058), .B(n14057), .Z(n14060) );
  XOR U14816 ( .A(n14059), .B(n14060), .Z(n14048) );
  XNOR U14817 ( .A(n14047), .B(n14048), .Z(n14074) );
  NANDN U14818 ( .A(n13925), .B(n13924), .Z(n13929) );
  OR U14819 ( .A(n13927), .B(n13926), .Z(n13928) );
  NAND U14820 ( .A(n13929), .B(n13928), .Z(n14079) );
  NANDN U14821 ( .A(n13931), .B(n13930), .Z(n13935) );
  NANDN U14822 ( .A(n13933), .B(n13932), .Z(n13934) );
  NAND U14823 ( .A(n13935), .B(n13934), .Z(n14078) );
  XOR U14824 ( .A(n14078), .B(n14077), .Z(n14080) );
  XOR U14825 ( .A(n14079), .B(n14080), .Z(n14073) );
  XOR U14826 ( .A(n14074), .B(n14073), .Z(n14075) );
  XOR U14827 ( .A(n14076), .B(n14075), .Z(n13973) );
  NAND U14828 ( .A(n13941), .B(n13940), .Z(n13945) );
  NAND U14829 ( .A(n13943), .B(n13942), .Z(n13944) );
  NAND U14830 ( .A(n13945), .B(n13944), .Z(n13972) );
  XOR U14831 ( .A(n13973), .B(n13972), .Z(n13975) );
  XNOR U14832 ( .A(n13974), .B(n13975), .Z(n14085) );
  NAND U14833 ( .A(n13947), .B(n13946), .Z(n13951) );
  NAND U14834 ( .A(n13949), .B(n13948), .Z(n13950) );
  NAND U14835 ( .A(n13951), .B(n13950), .Z(n14084) );
  NANDN U14836 ( .A(n13953), .B(n13952), .Z(n13957) );
  NAND U14837 ( .A(n13955), .B(n13954), .Z(n13956) );
  AND U14838 ( .A(n13957), .B(n13956), .Z(n14083) );
  XOR U14839 ( .A(n14084), .B(n14083), .Z(n14086) );
  XOR U14840 ( .A(n14085), .B(n14086), .Z(n14091) );
  NANDN U14841 ( .A(n13959), .B(n13958), .Z(n13963) );
  NANDN U14842 ( .A(n13961), .B(n13960), .Z(n13962) );
  NAND U14843 ( .A(n13963), .B(n13962), .Z(n14089) );
  NANDN U14844 ( .A(n13964), .B(n13965), .Z(n13970) );
  NOR U14845 ( .A(n13966), .B(n13965), .Z(n13968) );
  OR U14846 ( .A(n13968), .B(n13967), .Z(n13969) );
  AND U14847 ( .A(n13970), .B(n13969), .Z(n14090) );
  XOR U14848 ( .A(n14089), .B(n14090), .Z(n13971) );
  XNOR U14849 ( .A(n14091), .B(n13971), .Z(N310) );
  NAND U14850 ( .A(n13973), .B(n13972), .Z(n13977) );
  NAND U14851 ( .A(n13975), .B(n13974), .Z(n13976) );
  AND U14852 ( .A(n13977), .B(n13976), .Z(n14096) );
  NAND U14853 ( .A(n13979), .B(n13978), .Z(n13983) );
  NAND U14854 ( .A(n13981), .B(n13980), .Z(n13982) );
  NAND U14855 ( .A(n13983), .B(n13982), .Z(n14093) );
  NAND U14856 ( .A(n13985), .B(n13984), .Z(n13989) );
  NANDN U14857 ( .A(n13987), .B(n13986), .Z(n13988) );
  AND U14858 ( .A(n13989), .B(n13988), .Z(n14191) );
  NAND U14859 ( .A(n13991), .B(n13990), .Z(n13995) );
  NAND U14860 ( .A(n13993), .B(n13992), .Z(n13994) );
  NAND U14861 ( .A(n13995), .B(n13994), .Z(n14190) );
  XNOR U14862 ( .A(n14191), .B(n14190), .Z(n14193) );
  NAND U14863 ( .A(n13997), .B(n13996), .Z(n14001) );
  AND U14864 ( .A(n13999), .B(n13998), .Z(n14000) );
  ANDN U14865 ( .B(n14001), .A(n14000), .Z(n14155) );
  AND U14866 ( .A(y[1929]), .B(x[237]), .Z(n14003) );
  NAND U14867 ( .A(y[1922]), .B(x[244]), .Z(n14002) );
  XNOR U14868 ( .A(n14003), .B(n14002), .Z(n14175) );
  AND U14869 ( .A(x[226]), .B(y[1940]), .Z(n14174) );
  XOR U14870 ( .A(n14175), .B(n14174), .Z(n14153) );
  AND U14871 ( .A(y[1936]), .B(x[230]), .Z(n14005) );
  NAND U14872 ( .A(y[1927]), .B(x[239]), .Z(n14004) );
  XNOR U14873 ( .A(n14005), .B(n14004), .Z(n14187) );
  XOR U14874 ( .A(n14187), .B(n14186), .Z(n14152) );
  XOR U14875 ( .A(n14153), .B(n14152), .Z(n14154) );
  XNOR U14876 ( .A(n14155), .B(n14154), .Z(n14196) );
  AND U14877 ( .A(x[237]), .B(y[1938]), .Z(n15430) );
  NANDN U14878 ( .A(n14006), .B(n15430), .Z(n14010) );
  NAND U14879 ( .A(n14008), .B(n14007), .Z(n14009) );
  AND U14880 ( .A(n14010), .B(n14009), .Z(n14127) );
  AND U14881 ( .A(x[225]), .B(y[1941]), .Z(n14145) );
  XOR U14882 ( .A(n14146), .B(n14145), .Z(n14144) );
  AND U14883 ( .A(n14011), .B(o[149]), .Z(n14142) );
  XOR U14884 ( .A(n14144), .B(n14142), .Z(n14125) );
  AND U14885 ( .A(x[238]), .B(y[1928]), .Z(n14139) );
  AND U14886 ( .A(x[227]), .B(y[1939]), .Z(n14138) );
  XOR U14887 ( .A(n14139), .B(n14138), .Z(n14141) );
  AND U14888 ( .A(x[243]), .B(y[1923]), .Z(n14140) );
  XOR U14889 ( .A(n14141), .B(n14140), .Z(n14124) );
  XOR U14890 ( .A(n14125), .B(n14124), .Z(n14126) );
  XNOR U14891 ( .A(n14127), .B(n14126), .Z(n14197) );
  XOR U14892 ( .A(n14196), .B(n14197), .Z(n14199) );
  NAND U14893 ( .A(n14013), .B(n14012), .Z(n14017) );
  NAND U14894 ( .A(n14015), .B(n14014), .Z(n14016) );
  AND U14895 ( .A(n14017), .B(n14016), .Z(n14121) );
  AND U14896 ( .A(x[242]), .B(y[1931]), .Z(n15207) );
  NAND U14897 ( .A(n15207), .B(n14018), .Z(n14022) );
  NAND U14898 ( .A(n14020), .B(n14019), .Z(n14021) );
  NAND U14899 ( .A(n14022), .B(n14021), .Z(n14120) );
  XNOR U14900 ( .A(n14121), .B(n14120), .Z(n14123) );
  AND U14901 ( .A(x[238]), .B(y[1935]), .Z(n15144) );
  NAND U14902 ( .A(n15144), .B(n14185), .Z(n14025) );
  NAND U14903 ( .A(n14023), .B(n14235), .Z(n14024) );
  NAND U14904 ( .A(n14025), .B(n14024), .Z(n14130) );
  AND U14905 ( .A(x[224]), .B(y[1942]), .Z(n14162) );
  AND U14906 ( .A(x[246]), .B(y[1920]), .Z(n14161) );
  XOR U14907 ( .A(n14162), .B(n14161), .Z(n14164) );
  AND U14908 ( .A(x[245]), .B(y[1921]), .Z(n14184) );
  XOR U14909 ( .A(n14184), .B(o[150]), .Z(n14163) );
  XOR U14910 ( .A(n14164), .B(n14163), .Z(n14129) );
  AND U14911 ( .A(y[1935]), .B(x[231]), .Z(n14027) );
  NAND U14912 ( .A(y[1934]), .B(x[232]), .Z(n14026) );
  XNOR U14913 ( .A(n14027), .B(n14026), .Z(n14168) );
  XOR U14914 ( .A(n14168), .B(n14167), .Z(n14128) );
  XOR U14915 ( .A(n14129), .B(n14128), .Z(n14131) );
  XOR U14916 ( .A(n14130), .B(n14131), .Z(n14122) );
  XOR U14917 ( .A(n14123), .B(n14122), .Z(n14198) );
  XOR U14918 ( .A(n14199), .B(n14198), .Z(n14192) );
  XOR U14919 ( .A(n14193), .B(n14192), .Z(n14209) );
  NAND U14920 ( .A(x[243]), .B(y[1930]), .Z(n15205) );
  NANDN U14921 ( .A(n15205), .B(n14028), .Z(n14032) );
  NAND U14922 ( .A(n14030), .B(n14029), .Z(n14031) );
  AND U14923 ( .A(n14032), .B(n14031), .Z(n14203) );
  NAND U14924 ( .A(n14638), .B(n14156), .Z(n14036) );
  NAND U14925 ( .A(n14034), .B(n14033), .Z(n14035) );
  AND U14926 ( .A(n14036), .B(n14035), .Z(n14137) );
  AND U14927 ( .A(x[229]), .B(y[1937]), .Z(n14179) );
  AND U14928 ( .A(x[241]), .B(y[1925]), .Z(n14178) );
  XOR U14929 ( .A(n14179), .B(n14178), .Z(n14181) );
  AND U14930 ( .A(x[240]), .B(y[1926]), .Z(n14180) );
  XOR U14931 ( .A(n14181), .B(n14180), .Z(n14135) );
  AND U14932 ( .A(y[1924]), .B(x[242]), .Z(n14038) );
  NAND U14933 ( .A(y[1930]), .B(x[236]), .Z(n14037) );
  XNOR U14934 ( .A(n14038), .B(n14037), .Z(n14158) );
  AND U14935 ( .A(x[228]), .B(y[1938]), .Z(n14157) );
  XOR U14936 ( .A(n14158), .B(n14157), .Z(n14134) );
  XOR U14937 ( .A(n14135), .B(n14134), .Z(n14136) );
  XNOR U14938 ( .A(n14137), .B(n14136), .Z(n14202) );
  XNOR U14939 ( .A(n14203), .B(n14202), .Z(n14205) );
  NAND U14940 ( .A(n14040), .B(n14039), .Z(n14044) );
  NANDN U14941 ( .A(n14042), .B(n14041), .Z(n14043) );
  AND U14942 ( .A(n14044), .B(n14043), .Z(n14204) );
  XNOR U14943 ( .A(n14205), .B(n14204), .Z(n14208) );
  XNOR U14944 ( .A(n14209), .B(n14208), .Z(n14210) );
  NANDN U14945 ( .A(n14046), .B(n14045), .Z(n14050) );
  NANDN U14946 ( .A(n14048), .B(n14047), .Z(n14049) );
  NAND U14947 ( .A(n14050), .B(n14049), .Z(n14211) );
  XNOR U14948 ( .A(n14210), .B(n14211), .Z(n14111) );
  NANDN U14949 ( .A(n14052), .B(n14051), .Z(n14056) );
  NAND U14950 ( .A(n14054), .B(n14053), .Z(n14055) );
  AND U14951 ( .A(n14056), .B(n14055), .Z(n14116) );
  NANDN U14952 ( .A(n14058), .B(n14057), .Z(n14062) );
  NANDN U14953 ( .A(n14060), .B(n14059), .Z(n14061) );
  AND U14954 ( .A(n14062), .B(n14061), .Z(n14115) );
  XOR U14955 ( .A(n14115), .B(n14114), .Z(n14117) );
  XOR U14956 ( .A(n14116), .B(n14117), .Z(n14109) );
  NANDN U14957 ( .A(n14068), .B(n14067), .Z(n14072) );
  NANDN U14958 ( .A(n14070), .B(n14069), .Z(n14071) );
  NAND U14959 ( .A(n14072), .B(n14071), .Z(n14108) );
  XNOR U14960 ( .A(n14109), .B(n14108), .Z(n14110) );
  XOR U14961 ( .A(n14111), .B(n14110), .Z(n14105) );
  NAND U14962 ( .A(n14078), .B(n14077), .Z(n14082) );
  NAND U14963 ( .A(n14080), .B(n14079), .Z(n14081) );
  NAND U14964 ( .A(n14082), .B(n14081), .Z(n14102) );
  XNOR U14965 ( .A(n14103), .B(n14102), .Z(n14104) );
  XNOR U14966 ( .A(n14105), .B(n14104), .Z(n14094) );
  XOR U14967 ( .A(n14093), .B(n14094), .Z(n14095) );
  XNOR U14968 ( .A(n14096), .B(n14095), .Z(n14101) );
  NAND U14969 ( .A(n14084), .B(n14083), .Z(n14088) );
  NAND U14970 ( .A(n14086), .B(n14085), .Z(n14087) );
  NAND U14971 ( .A(n14088), .B(n14087), .Z(n14100) );
  XOR U14972 ( .A(n14100), .B(n14099), .Z(n14092) );
  XNOR U14973 ( .A(n14101), .B(n14092), .Z(N311) );
  NAND U14974 ( .A(n14094), .B(n14093), .Z(n14098) );
  NAND U14975 ( .A(n14096), .B(n14095), .Z(n14097) );
  NAND U14976 ( .A(n14098), .B(n14097), .Z(n14340) );
  NANDN U14977 ( .A(n14103), .B(n14102), .Z(n14107) );
  NANDN U14978 ( .A(n14105), .B(n14104), .Z(n14106) );
  AND U14979 ( .A(n14107), .B(n14106), .Z(n14336) );
  NANDN U14980 ( .A(n14109), .B(n14108), .Z(n14113) );
  NAND U14981 ( .A(n14111), .B(n14110), .Z(n14112) );
  AND U14982 ( .A(n14113), .B(n14112), .Z(n14335) );
  NANDN U14983 ( .A(n14115), .B(n14114), .Z(n14119) );
  OR U14984 ( .A(n14117), .B(n14116), .Z(n14118) );
  NAND U14985 ( .A(n14119), .B(n14118), .Z(n14319) );
  NAND U14986 ( .A(n14129), .B(n14128), .Z(n14133) );
  NAND U14987 ( .A(n14131), .B(n14130), .Z(n14132) );
  NAND U14988 ( .A(n14133), .B(n14132), .Z(n14310) );
  XOR U14989 ( .A(n14311), .B(n14310), .Z(n14313) );
  XOR U14990 ( .A(n14312), .B(n14313), .Z(n14330) );
  IV U14991 ( .A(n14142), .Z(n14143) );
  ANDN U14992 ( .B(n14144), .A(n14143), .Z(n14148) );
  NAND U14993 ( .A(n14146), .B(n14145), .Z(n14147) );
  NANDN U14994 ( .A(n14148), .B(n14147), .Z(n14265) );
  XOR U14995 ( .A(n14264), .B(n14265), .Z(n14267) );
  AND U14996 ( .A(y[1936]), .B(x[231]), .Z(n14150) );
  NAND U14997 ( .A(y[1934]), .B(x[233]), .Z(n14149) );
  XNOR U14998 ( .A(n14150), .B(n14149), .Z(n14236) );
  XOR U14999 ( .A(n14236), .B(n14151), .Z(n14269) );
  AND U15000 ( .A(x[234]), .B(y[1933]), .Z(n14268) );
  XOR U15001 ( .A(n14269), .B(n14268), .Z(n14271) );
  AND U15002 ( .A(x[230]), .B(y[1937]), .Z(n14227) );
  NAND U15003 ( .A(x[239]), .B(y[1928]), .Z(n14228) );
  XNOR U15004 ( .A(n14227), .B(n14228), .Z(n14230) );
  AND U15005 ( .A(x[235]), .B(y[1932]), .Z(n14229) );
  XOR U15006 ( .A(n14230), .B(n14229), .Z(n14270) );
  XOR U15007 ( .A(n14271), .B(n14270), .Z(n14266) );
  XOR U15008 ( .A(n14267), .B(n14266), .Z(n14329) );
  XNOR U15009 ( .A(n14328), .B(n14329), .Z(n14331) );
  AND U15010 ( .A(x[242]), .B(y[1930]), .Z(n15012) );
  NAND U15011 ( .A(n15012), .B(n14156), .Z(n14160) );
  NAND U15012 ( .A(n14158), .B(n14157), .Z(n14159) );
  NAND U15013 ( .A(n14160), .B(n14159), .Z(n14287) );
  NAND U15014 ( .A(n14162), .B(n14161), .Z(n14166) );
  NAND U15015 ( .A(n14164), .B(n14163), .Z(n14165) );
  NAND U15016 ( .A(n14166), .B(n14165), .Z(n14286) );
  XOR U15017 ( .A(n14287), .B(n14286), .Z(n14288) );
  NANDN U15018 ( .A(n14237), .B(n14235), .Z(n14170) );
  NAND U15019 ( .A(n14168), .B(n14167), .Z(n14169) );
  NAND U15020 ( .A(n14170), .B(n14169), .Z(n14300) );
  AND U15021 ( .A(x[224]), .B(y[1943]), .Z(n14245) );
  AND U15022 ( .A(x[247]), .B(y[1920]), .Z(n14244) );
  XOR U15023 ( .A(n14245), .B(n14244), .Z(n14247) );
  AND U15024 ( .A(x[246]), .B(y[1921]), .Z(n14226) );
  XOR U15025 ( .A(n14226), .B(o[151]), .Z(n14246) );
  XOR U15026 ( .A(n14247), .B(n14246), .Z(n14299) );
  NAND U15027 ( .A(y[1923]), .B(x[244]), .Z(n14171) );
  XNOR U15028 ( .A(n14172), .B(n14171), .Z(n14222) );
  NAND U15029 ( .A(x[243]), .B(y[1924]), .Z(n14223) );
  XNOR U15030 ( .A(n14222), .B(n14223), .Z(n14298) );
  XOR U15031 ( .A(n14299), .B(n14298), .Z(n14301) );
  XNOR U15032 ( .A(n14300), .B(n14301), .Z(n14289) );
  XOR U15033 ( .A(n14258), .B(n14259), .Z(n14261) );
  NAND U15034 ( .A(x[244]), .B(y[1929]), .Z(n15156) );
  AND U15035 ( .A(x[237]), .B(y[1922]), .Z(n14173) );
  NANDN U15036 ( .A(n15156), .B(n14173), .Z(n14177) );
  NAND U15037 ( .A(n14175), .B(n14174), .Z(n14176) );
  NAND U15038 ( .A(n14177), .B(n14176), .Z(n14252) );
  NAND U15039 ( .A(n14179), .B(n14178), .Z(n14183) );
  NAND U15040 ( .A(n14181), .B(n14180), .Z(n14182) );
  NAND U15041 ( .A(n14183), .B(n14182), .Z(n14306) );
  AND U15042 ( .A(x[237]), .B(y[1930]), .Z(n14283) );
  AND U15043 ( .A(x[226]), .B(y[1941]), .Z(n14282) );
  XOR U15044 ( .A(n14283), .B(n14282), .Z(n14285) );
  AND U15045 ( .A(x[245]), .B(y[1922]), .Z(n14284) );
  XOR U15046 ( .A(n14285), .B(n14284), .Z(n14305) );
  AND U15047 ( .A(x[236]), .B(y[1931]), .Z(n14241) );
  AND U15048 ( .A(x[225]), .B(y[1942]), .Z(n14240) );
  XOR U15049 ( .A(n14241), .B(n14240), .Z(n14243) );
  AND U15050 ( .A(n14184), .B(o[150]), .Z(n14242) );
  XOR U15051 ( .A(n14243), .B(n14242), .Z(n14304) );
  XOR U15052 ( .A(n14305), .B(n14304), .Z(n14307) );
  XOR U15053 ( .A(n14306), .B(n14307), .Z(n14253) );
  XOR U15054 ( .A(n14252), .B(n14253), .Z(n14255) );
  AND U15055 ( .A(x[239]), .B(y[1936]), .Z(n15340) );
  NAND U15056 ( .A(n15340), .B(n14185), .Z(n14189) );
  NAND U15057 ( .A(n14187), .B(n14186), .Z(n14188) );
  NAND U15058 ( .A(n14189), .B(n14188), .Z(n14294) );
  AND U15059 ( .A(x[238]), .B(y[1929]), .Z(n14279) );
  AND U15060 ( .A(x[227]), .B(y[1940]), .Z(n14278) );
  XOR U15061 ( .A(n14279), .B(n14278), .Z(n14281) );
  AND U15062 ( .A(x[228]), .B(y[1939]), .Z(n14280) );
  XOR U15063 ( .A(n14281), .B(n14280), .Z(n14293) );
  AND U15064 ( .A(x[229]), .B(y[1938]), .Z(n14272) );
  NAND U15065 ( .A(x[242]), .B(y[1925]), .Z(n14273) );
  XNOR U15066 ( .A(n14272), .B(n14273), .Z(n14275) );
  AND U15067 ( .A(x[241]), .B(y[1926]), .Z(n14274) );
  XOR U15068 ( .A(n14275), .B(n14274), .Z(n14292) );
  XOR U15069 ( .A(n14293), .B(n14292), .Z(n14295) );
  XOR U15070 ( .A(n14294), .B(n14295), .Z(n14254) );
  XOR U15071 ( .A(n14255), .B(n14254), .Z(n14260) );
  XOR U15072 ( .A(n14261), .B(n14260), .Z(n14316) );
  XOR U15073 ( .A(n14317), .B(n14316), .Z(n14318) );
  XNOR U15074 ( .A(n14319), .B(n14318), .Z(n14217) );
  NANDN U15075 ( .A(n14191), .B(n14190), .Z(n14195) );
  NAND U15076 ( .A(n14193), .B(n14192), .Z(n14194) );
  NAND U15077 ( .A(n14195), .B(n14194), .Z(n14325) );
  NAND U15078 ( .A(n14197), .B(n14196), .Z(n14201) );
  NAND U15079 ( .A(n14199), .B(n14198), .Z(n14200) );
  NAND U15080 ( .A(n14201), .B(n14200), .Z(n14323) );
  NANDN U15081 ( .A(n14203), .B(n14202), .Z(n14207) );
  NAND U15082 ( .A(n14205), .B(n14204), .Z(n14206) );
  NAND U15083 ( .A(n14207), .B(n14206), .Z(n14322) );
  XOR U15084 ( .A(n14323), .B(n14322), .Z(n14324) );
  XNOR U15085 ( .A(n14325), .B(n14324), .Z(n14216) );
  NANDN U15086 ( .A(n14209), .B(n14208), .Z(n14213) );
  NANDN U15087 ( .A(n14211), .B(n14210), .Z(n14212) );
  NAND U15088 ( .A(n14213), .B(n14212), .Z(n14215) );
  XOR U15089 ( .A(n14216), .B(n14215), .Z(n14218) );
  XOR U15090 ( .A(n14217), .B(n14218), .Z(n14334) );
  XOR U15091 ( .A(n14335), .B(n14334), .Z(n14337) );
  XNOR U15092 ( .A(n14336), .B(n14337), .Z(n14342) );
  XNOR U15093 ( .A(n14341), .B(n14342), .Z(n14214) );
  XNOR U15094 ( .A(n14340), .B(n14214), .Z(N312) );
  NAND U15095 ( .A(n14216), .B(n14215), .Z(n14220) );
  NAND U15096 ( .A(n14218), .B(n14217), .Z(n14219) );
  AND U15097 ( .A(n14220), .B(n14219), .Z(n14464) );
  AND U15098 ( .A(x[244]), .B(y[1927]), .Z(n14221) );
  NAND U15099 ( .A(n14221), .B(n14371), .Z(n14225) );
  NANDN U15100 ( .A(n14223), .B(n14222), .Z(n14224) );
  AND U15101 ( .A(n14225), .B(n14224), .Z(n14389) );
  AND U15102 ( .A(x[246]), .B(y[1922]), .Z(n14422) );
  XOR U15103 ( .A(n14423), .B(n14422), .Z(n14424) );
  AND U15104 ( .A(x[226]), .B(y[1942]), .Z(n14425) );
  XOR U15105 ( .A(n14424), .B(n14425), .Z(n14387) );
  AND U15106 ( .A(n14226), .B(o[151]), .Z(n14429) );
  AND U15107 ( .A(x[225]), .B(y[1943]), .Z(n14430) );
  XOR U15108 ( .A(n14431), .B(n14430), .Z(n14428) );
  XOR U15109 ( .A(n14429), .B(n14428), .Z(n14386) );
  XOR U15110 ( .A(n14387), .B(n14386), .Z(n14388) );
  XNOR U15111 ( .A(n14389), .B(n14388), .Z(n14442) );
  NANDN U15112 ( .A(n14228), .B(n14227), .Z(n14232) );
  NAND U15113 ( .A(n14230), .B(n14229), .Z(n14231) );
  AND U15114 ( .A(n14232), .B(n14231), .Z(n14385) );
  AND U15115 ( .A(y[1928]), .B(x[240]), .Z(n14234) );
  NAND U15116 ( .A(y[1923]), .B(x[245]), .Z(n14233) );
  XNOR U15117 ( .A(n14234), .B(n14233), .Z(n14372) );
  AND U15118 ( .A(x[229]), .B(y[1939]), .Z(n14373) );
  XOR U15119 ( .A(n14372), .B(n14373), .Z(n14383) );
  AND U15120 ( .A(x[230]), .B(y[1938]), .Z(n14730) );
  AND U15121 ( .A(x[244]), .B(y[1924]), .Z(n14560) );
  XOR U15122 ( .A(n14730), .B(n14560), .Z(n14378) );
  AND U15123 ( .A(x[243]), .B(y[1925]), .Z(n14379) );
  XOR U15124 ( .A(n14378), .B(n14379), .Z(n14382) );
  XOR U15125 ( .A(n14383), .B(n14382), .Z(n14384) );
  XNOR U15126 ( .A(n14385), .B(n14384), .Z(n14364) );
  NANDN U15127 ( .A(n14491), .B(n14235), .Z(n14239) );
  NANDN U15128 ( .A(n14237), .B(n14236), .Z(n14238) );
  NAND U15129 ( .A(n14239), .B(n14238), .Z(n14360) );
  XOR U15130 ( .A(n14360), .B(n14361), .Z(n14363) );
  XOR U15131 ( .A(n14364), .B(n14363), .Z(n14441) );
  XOR U15132 ( .A(n14442), .B(n14441), .Z(n14444) );
  AND U15133 ( .A(x[227]), .B(y[1941]), .Z(n14400) );
  XOR U15134 ( .A(n14401), .B(n14400), .Z(n14403) );
  NAND U15135 ( .A(x[228]), .B(y[1940]), .Z(n14402) );
  XNOR U15136 ( .A(n14403), .B(n14402), .Z(n14397) );
  XOR U15137 ( .A(n14396), .B(n14397), .Z(n14399) );
  AND U15138 ( .A(y[1935]), .B(x[233]), .Z(n14249) );
  NAND U15139 ( .A(y[1934]), .B(x[234]), .Z(n14248) );
  XNOR U15140 ( .A(n14249), .B(n14248), .Z(n14413) );
  AND U15141 ( .A(y[1930]), .B(x[238]), .Z(n14251) );
  NAND U15142 ( .A(y[1936]), .B(x[232]), .Z(n14250) );
  XNOR U15143 ( .A(n14251), .B(n14250), .Z(n14418) );
  NAND U15144 ( .A(x[235]), .B(y[1933]), .Z(n14419) );
  XOR U15145 ( .A(n14418), .B(n14419), .Z(n14414) );
  XNOR U15146 ( .A(n14413), .B(n14414), .Z(n14398) );
  XOR U15147 ( .A(n14399), .B(n14398), .Z(n14443) );
  XOR U15148 ( .A(n14444), .B(n14443), .Z(n14450) );
  NAND U15149 ( .A(n14253), .B(n14252), .Z(n14257) );
  NAND U15150 ( .A(n14255), .B(n14254), .Z(n14256) );
  AND U15151 ( .A(n14257), .B(n14256), .Z(n14449) );
  NAND U15152 ( .A(n14259), .B(n14258), .Z(n14263) );
  NAND U15153 ( .A(n14261), .B(n14260), .Z(n14262) );
  AND U15154 ( .A(n14263), .B(n14262), .Z(n14451) );
  XOR U15155 ( .A(n14452), .B(n14451), .Z(n14458) );
  NANDN U15156 ( .A(n14273), .B(n14272), .Z(n14277) );
  NAND U15157 ( .A(n14275), .B(n14274), .Z(n14276) );
  AND U15158 ( .A(n14277), .B(n14276), .Z(n14370) );
  AND U15159 ( .A(x[224]), .B(y[1944]), .Z(n14407) );
  AND U15160 ( .A(x[248]), .B(y[1920]), .Z(n14406) );
  XOR U15161 ( .A(n14407), .B(n14406), .Z(n14409) );
  AND U15162 ( .A(x[247]), .B(y[1921]), .Z(n14440) );
  XOR U15163 ( .A(n14440), .B(o[152]), .Z(n14408) );
  XOR U15164 ( .A(n14409), .B(n14408), .Z(n14368) );
  AND U15165 ( .A(x[231]), .B(y[1937]), .Z(n14434) );
  AND U15166 ( .A(x[242]), .B(y[1926]), .Z(n14435) );
  XOR U15167 ( .A(n14434), .B(n14435), .Z(n14436) );
  AND U15168 ( .A(x[241]), .B(y[1927]), .Z(n14437) );
  XOR U15169 ( .A(n14436), .B(n14437), .Z(n14367) );
  XOR U15170 ( .A(n14368), .B(n14367), .Z(n14369) );
  XNOR U15171 ( .A(n14370), .B(n14369), .Z(n14358) );
  XNOR U15172 ( .A(n14356), .B(n14357), .Z(n14359) );
  XNOR U15173 ( .A(n14358), .B(n14359), .Z(n14446) );
  XOR U15174 ( .A(n14445), .B(n14446), .Z(n14448) );
  XOR U15175 ( .A(n14447), .B(n14448), .Z(n14353) );
  NAND U15176 ( .A(n14287), .B(n14286), .Z(n14291) );
  NANDN U15177 ( .A(n14289), .B(n14288), .Z(n14290) );
  AND U15178 ( .A(n14291), .B(n14290), .Z(n14393) );
  NAND U15179 ( .A(n14293), .B(n14292), .Z(n14297) );
  NAND U15180 ( .A(n14295), .B(n14294), .Z(n14296) );
  AND U15181 ( .A(n14297), .B(n14296), .Z(n14391) );
  NAND U15182 ( .A(n14299), .B(n14298), .Z(n14303) );
  NAND U15183 ( .A(n14301), .B(n14300), .Z(n14302) );
  AND U15184 ( .A(n14303), .B(n14302), .Z(n14390) );
  XOR U15185 ( .A(n14391), .B(n14390), .Z(n14392) );
  XOR U15186 ( .A(n14393), .B(n14392), .Z(n14351) );
  NAND U15187 ( .A(n14305), .B(n14304), .Z(n14309) );
  NAND U15188 ( .A(n14307), .B(n14306), .Z(n14308) );
  AND U15189 ( .A(n14309), .B(n14308), .Z(n14350) );
  XOR U15190 ( .A(n14351), .B(n14350), .Z(n14352) );
  NAND U15191 ( .A(n14311), .B(n14310), .Z(n14315) );
  NAND U15192 ( .A(n14313), .B(n14312), .Z(n14314) );
  AND U15193 ( .A(n14315), .B(n14314), .Z(n14455) );
  XOR U15194 ( .A(n14456), .B(n14455), .Z(n14457) );
  XNOR U15195 ( .A(n14458), .B(n14457), .Z(n14462) );
  NAND U15196 ( .A(n14317), .B(n14316), .Z(n14321) );
  NAND U15197 ( .A(n14319), .B(n14318), .Z(n14320) );
  NAND U15198 ( .A(n14321), .B(n14320), .Z(n14346) );
  NAND U15199 ( .A(n14323), .B(n14322), .Z(n14327) );
  NAND U15200 ( .A(n14325), .B(n14324), .Z(n14326) );
  NAND U15201 ( .A(n14327), .B(n14326), .Z(n14345) );
  NAND U15202 ( .A(n14329), .B(n14328), .Z(n14333) );
  NANDN U15203 ( .A(n14331), .B(n14330), .Z(n14332) );
  NAND U15204 ( .A(n14333), .B(n14332), .Z(n14344) );
  XOR U15205 ( .A(n14345), .B(n14344), .Z(n14347) );
  XOR U15206 ( .A(n14346), .B(n14347), .Z(n14461) );
  XOR U15207 ( .A(n14462), .B(n14461), .Z(n14463) );
  XOR U15208 ( .A(n14464), .B(n14463), .Z(n14469) );
  NANDN U15209 ( .A(n14335), .B(n14334), .Z(n14339) );
  NANDN U15210 ( .A(n14337), .B(n14336), .Z(n14338) );
  AND U15211 ( .A(n14339), .B(n14338), .Z(n14468) );
  XOR U15212 ( .A(n14468), .B(n14467), .Z(n14343) );
  XNOR U15213 ( .A(n14469), .B(n14343), .Z(N313) );
  NAND U15214 ( .A(n14345), .B(n14344), .Z(n14349) );
  NAND U15215 ( .A(n14347), .B(n14346), .Z(n14348) );
  AND U15216 ( .A(n14349), .B(n14348), .Z(n14603) );
  NAND U15217 ( .A(n14351), .B(n14350), .Z(n14355) );
  NANDN U15218 ( .A(n14353), .B(n14352), .Z(n14354) );
  NAND U15219 ( .A(n14355), .B(n14354), .Z(n14479) );
  IV U15220 ( .A(n14360), .Z(n14362) );
  NANDN U15221 ( .A(n14362), .B(n14361), .Z(n14366) );
  NAND U15222 ( .A(n14364), .B(n14363), .Z(n14365) );
  NAND U15223 ( .A(n14366), .B(n14365), .Z(n14484) );
  XOR U15224 ( .A(n14483), .B(n14484), .Z(n14486) );
  NAND U15225 ( .A(x[245]), .B(y[1928]), .Z(n15316) );
  NANDN U15226 ( .A(n15316), .B(n14371), .Z(n14375) );
  NAND U15227 ( .A(n14373), .B(n14372), .Z(n14374) );
  NAND U15228 ( .A(n14375), .B(n14374), .Z(n14580) );
  NAND U15229 ( .A(x[246]), .B(y[1923]), .Z(n14549) );
  NAND U15230 ( .A(x[229]), .B(y[1940]), .Z(n14548) );
  NAND U15231 ( .A(x[241]), .B(y[1928]), .Z(n14547) );
  XOR U15232 ( .A(n14548), .B(n14547), .Z(n14550) );
  XNOR U15233 ( .A(n14549), .B(n14550), .Z(n14579) );
  AND U15234 ( .A(y[1925]), .B(x[244]), .Z(n14377) );
  NAND U15235 ( .A(y[1924]), .B(x[245]), .Z(n14376) );
  XNOR U15236 ( .A(n14377), .B(n14376), .Z(n14562) );
  AND U15237 ( .A(x[243]), .B(y[1926]), .Z(n14561) );
  XOR U15238 ( .A(n14562), .B(n14561), .Z(n14578) );
  XNOR U15239 ( .A(n14579), .B(n14578), .Z(n14581) );
  XOR U15240 ( .A(n14580), .B(n14581), .Z(n14504) );
  NAND U15241 ( .A(n14560), .B(n14730), .Z(n14381) );
  NAND U15242 ( .A(n14379), .B(n14378), .Z(n14380) );
  NAND U15243 ( .A(n14381), .B(n14380), .Z(n14586) );
  NAND U15244 ( .A(x[239]), .B(y[1930]), .Z(n14568) );
  NAND U15245 ( .A(x[242]), .B(y[1927]), .Z(n14567) );
  NAND U15246 ( .A(x[230]), .B(y[1939]), .Z(n14566) );
  XOR U15247 ( .A(n14567), .B(n14566), .Z(n14569) );
  XNOR U15248 ( .A(n14568), .B(n14569), .Z(n14585) );
  NAND U15249 ( .A(x[247]), .B(y[1922]), .Z(n14543) );
  NAND U15250 ( .A(x[228]), .B(y[1941]), .Z(n14542) );
  NAND U15251 ( .A(x[240]), .B(y[1929]), .Z(n14541) );
  XOR U15252 ( .A(n14542), .B(n14541), .Z(n14544) );
  XNOR U15253 ( .A(n14543), .B(n14544), .Z(n14584) );
  XNOR U15254 ( .A(n14585), .B(n14584), .Z(n14587) );
  XOR U15255 ( .A(n14586), .B(n14587), .Z(n14503) );
  XOR U15256 ( .A(n14504), .B(n14503), .Z(n14505) );
  XOR U15257 ( .A(n14506), .B(n14505), .Z(n14517) );
  XOR U15258 ( .A(n14516), .B(n14515), .Z(n14518) );
  XOR U15259 ( .A(n14517), .B(n14518), .Z(n14485) );
  XOR U15260 ( .A(n14486), .B(n14485), .Z(n14478) );
  NAND U15261 ( .A(n14391), .B(n14390), .Z(n14395) );
  NAND U15262 ( .A(n14393), .B(n14392), .Z(n14394) );
  NAND U15263 ( .A(n14395), .B(n14394), .Z(n14477) );
  XOR U15264 ( .A(n14479), .B(n14480), .Z(n14474) );
  NAND U15265 ( .A(n14401), .B(n14400), .Z(n14405) );
  ANDN U15266 ( .B(n14403), .A(n14402), .Z(n14404) );
  ANDN U15267 ( .B(n14405), .A(n14404), .Z(n14575) );
  NAND U15268 ( .A(n14407), .B(n14406), .Z(n14411) );
  NAND U15269 ( .A(n14409), .B(n14408), .Z(n14410) );
  AND U15270 ( .A(n14411), .B(n14410), .Z(n14573) );
  AND U15271 ( .A(x[238]), .B(y[1931]), .Z(n14529) );
  NAND U15272 ( .A(x[226]), .B(y[1943]), .Z(n14530) );
  XNOR U15273 ( .A(n14529), .B(n14530), .Z(n14531) );
  NAND U15274 ( .A(x[227]), .B(y[1942]), .Z(n14532) );
  XNOR U15275 ( .A(n14531), .B(n14532), .Z(n14572) );
  XNOR U15276 ( .A(n14573), .B(n14572), .Z(n14574) );
  XOR U15277 ( .A(n14575), .B(n14574), .Z(n14590) );
  XOR U15278 ( .A(n14591), .B(n14590), .Z(n14593) );
  NANDN U15279 ( .A(n14492), .B(n14412), .Z(n14416) );
  NANDN U15280 ( .A(n14414), .B(n14413), .Z(n14415) );
  AND U15281 ( .A(n14416), .B(n14415), .Z(n14510) );
  AND U15282 ( .A(x[238]), .B(y[1936]), .Z(n15354) );
  NAND U15283 ( .A(n15354), .B(n14417), .Z(n14421) );
  NANDN U15284 ( .A(n14419), .B(n14418), .Z(n14420) );
  AND U15285 ( .A(n14421), .B(n14420), .Z(n14538) );
  NAND U15286 ( .A(x[235]), .B(y[1934]), .Z(n14556) );
  NAND U15287 ( .A(x[236]), .B(y[1933]), .Z(n14555) );
  NAND U15288 ( .A(x[231]), .B(y[1938]), .Z(n14554) );
  XOR U15289 ( .A(n14555), .B(n14554), .Z(n14557) );
  XOR U15290 ( .A(n14556), .B(n14557), .Z(n14536) );
  AND U15291 ( .A(x[248]), .B(y[1921]), .Z(n14553) );
  XOR U15292 ( .A(o[153]), .B(n14553), .Z(n14523) );
  NAND U15293 ( .A(x[225]), .B(y[1944]), .Z(n14524) );
  XNOR U15294 ( .A(n14523), .B(n14524), .Z(n14525) );
  NAND U15295 ( .A(x[237]), .B(y[1932]), .Z(n14526) );
  XNOR U15296 ( .A(n14525), .B(n14526), .Z(n14535) );
  XNOR U15297 ( .A(n14536), .B(n14535), .Z(n14537) );
  XNOR U15298 ( .A(n14538), .B(n14537), .Z(n14509) );
  XNOR U15299 ( .A(n14510), .B(n14509), .Z(n14511) );
  AND U15300 ( .A(n14423), .B(n14422), .Z(n14427) );
  NAND U15301 ( .A(n14425), .B(n14424), .Z(n14426) );
  NANDN U15302 ( .A(n14427), .B(n14426), .Z(n14499) );
  AND U15303 ( .A(n14429), .B(n14428), .Z(n14433) );
  NAND U15304 ( .A(n14431), .B(n14430), .Z(n14432) );
  NANDN U15305 ( .A(n14433), .B(n14432), .Z(n14500) );
  XOR U15306 ( .A(n14499), .B(n14500), .Z(n14501) );
  NAND U15307 ( .A(n14435), .B(n14434), .Z(n14439) );
  NAND U15308 ( .A(n14437), .B(n14436), .Z(n14438) );
  NAND U15309 ( .A(n14439), .B(n14438), .Z(n14498) );
  NAND U15310 ( .A(x[232]), .B(y[1937]), .Z(n14493) );
  XOR U15311 ( .A(n14491), .B(n14492), .Z(n14494) );
  XOR U15312 ( .A(n14493), .B(n14494), .Z(n14496) );
  NAND U15313 ( .A(n14440), .B(o[152]), .Z(n14489) );
  NAND U15314 ( .A(x[249]), .B(y[1920]), .Z(n14487) );
  NAND U15315 ( .A(x[224]), .B(y[1945]), .Z(n14488) );
  XOR U15316 ( .A(n14487), .B(n14488), .Z(n14490) );
  XOR U15317 ( .A(n14489), .B(n14490), .Z(n14495) );
  XOR U15318 ( .A(n14496), .B(n14495), .Z(n14497) );
  XNOR U15319 ( .A(n14498), .B(n14497), .Z(n14502) );
  XOR U15320 ( .A(n14501), .B(n14502), .Z(n14512) );
  XOR U15321 ( .A(n14511), .B(n14512), .Z(n14592) );
  XOR U15322 ( .A(n14593), .B(n14592), .Z(n14595) );
  XOR U15323 ( .A(n14595), .B(n14594), .Z(n14597) );
  XOR U15324 ( .A(n14597), .B(n14596), .Z(n14472) );
  NANDN U15325 ( .A(n14450), .B(n14449), .Z(n14454) );
  NAND U15326 ( .A(n14452), .B(n14451), .Z(n14453) );
  AND U15327 ( .A(n14454), .B(n14453), .Z(n14471) );
  NAND U15328 ( .A(n14456), .B(n14455), .Z(n14460) );
  NAND U15329 ( .A(n14458), .B(n14457), .Z(n14459) );
  NAND U15330 ( .A(n14460), .B(n14459), .Z(n14601) );
  XNOR U15331 ( .A(n14603), .B(n14604), .Z(n14600) );
  NAND U15332 ( .A(n14462), .B(n14461), .Z(n14466) );
  NAND U15333 ( .A(n14464), .B(n14463), .Z(n14465) );
  NAND U15334 ( .A(n14466), .B(n14465), .Z(n14599) );
  XOR U15335 ( .A(n14599), .B(n14598), .Z(n14470) );
  XNOR U15336 ( .A(n14600), .B(n14470), .Z(N314) );
  NANDN U15337 ( .A(n14472), .B(n14471), .Z(n14476) );
  NANDN U15338 ( .A(n14474), .B(n14473), .Z(n14475) );
  NAND U15339 ( .A(n14476), .B(n14475), .Z(n14752) );
  NANDN U15340 ( .A(n14478), .B(n14477), .Z(n14482) );
  NAND U15341 ( .A(n14480), .B(n14479), .Z(n14481) );
  AND U15342 ( .A(n14482), .B(n14481), .Z(n14753) );
  XOR U15343 ( .A(n14752), .B(n14753), .Z(n14755) );
  AND U15344 ( .A(x[226]), .B(y[1944]), .Z(n14624) );
  XOR U15345 ( .A(n14625), .B(n14624), .Z(n14627) );
  AND U15346 ( .A(x[248]), .B(y[1922]), .Z(n14626) );
  XOR U15347 ( .A(n14627), .B(n14626), .Z(n14661) );
  XOR U15348 ( .A(n14661), .B(n14660), .Z(n14663) );
  XNOR U15349 ( .A(n14663), .B(n14662), .Z(n14699) );
  XOR U15350 ( .A(n14699), .B(n14698), .Z(n14701) );
  XOR U15351 ( .A(n14701), .B(n14700), .Z(n14745) );
  NAND U15352 ( .A(n14504), .B(n14503), .Z(n14508) );
  NAND U15353 ( .A(n14506), .B(n14505), .Z(n14507) );
  NAND U15354 ( .A(n14508), .B(n14507), .Z(n14743) );
  NANDN U15355 ( .A(n14510), .B(n14509), .Z(n14514) );
  NANDN U15356 ( .A(n14512), .B(n14511), .Z(n14513) );
  AND U15357 ( .A(n14514), .B(n14513), .Z(n14742) );
  XOR U15358 ( .A(n14743), .B(n14742), .Z(n14744) );
  XOR U15359 ( .A(n14745), .B(n14744), .Z(n14749) );
  NANDN U15360 ( .A(n14516), .B(n14515), .Z(n14520) );
  OR U15361 ( .A(n14518), .B(n14517), .Z(n14519) );
  NAND U15362 ( .A(n14520), .B(n14519), .Z(n14695) );
  AND U15363 ( .A(x[236]), .B(y[1934]), .Z(n14820) );
  AND U15364 ( .A(x[229]), .B(y[1941]), .Z(n14675) );
  XOR U15365 ( .A(n14820), .B(n14675), .Z(n14677) );
  AND U15366 ( .A(x[234]), .B(y[1936]), .Z(n14676) );
  XOR U15367 ( .A(n14677), .B(n14676), .Z(n14707) );
  AND U15368 ( .A(y[1940]), .B(x[230]), .Z(n14522) );
  NAND U15369 ( .A(y[1938]), .B(x[232]), .Z(n14521) );
  XNOR U15370 ( .A(n14522), .B(n14521), .Z(n14732) );
  AND U15371 ( .A(x[233]), .B(y[1937]), .Z(n14731) );
  XOR U15372 ( .A(n14732), .B(n14731), .Z(n14704) );
  AND U15373 ( .A(x[231]), .B(y[1939]), .Z(n14705) );
  XOR U15374 ( .A(n14704), .B(n14705), .Z(n14706) );
  XOR U15375 ( .A(n14707), .B(n14706), .Z(n14651) );
  NANDN U15376 ( .A(n14524), .B(n14523), .Z(n14528) );
  NANDN U15377 ( .A(n14526), .B(n14525), .Z(n14527) );
  NAND U15378 ( .A(n14528), .B(n14527), .Z(n14649) );
  NANDN U15379 ( .A(n14530), .B(n14529), .Z(n14534) );
  NANDN U15380 ( .A(n14532), .B(n14531), .Z(n14533) );
  NAND U15381 ( .A(n14534), .B(n14533), .Z(n14648) );
  XOR U15382 ( .A(n14649), .B(n14648), .Z(n14650) );
  XNOR U15383 ( .A(n14651), .B(n14650), .Z(n14687) );
  NANDN U15384 ( .A(n14536), .B(n14535), .Z(n14540) );
  NANDN U15385 ( .A(n14538), .B(n14537), .Z(n14539) );
  AND U15386 ( .A(n14540), .B(n14539), .Z(n14686) );
  XOR U15387 ( .A(n14687), .B(n14686), .Z(n14689) );
  NAND U15388 ( .A(n14542), .B(n14541), .Z(n14546) );
  NAND U15389 ( .A(n14544), .B(n14543), .Z(n14545) );
  AND U15390 ( .A(n14546), .B(n14545), .Z(n14612) );
  NAND U15391 ( .A(n14548), .B(n14547), .Z(n14552) );
  NAND U15392 ( .A(n14550), .B(n14549), .Z(n14551) );
  AND U15393 ( .A(n14552), .B(n14551), .Z(n14613) );
  XOR U15394 ( .A(n14612), .B(n14613), .Z(n14615) );
  AND U15395 ( .A(n14553), .B(o[153]), .Z(n14724) );
  AND U15396 ( .A(x[238]), .B(y[1932]), .Z(n14725) );
  XOR U15397 ( .A(n14724), .B(n14725), .Z(n14726) );
  AND U15398 ( .A(x[225]), .B(y[1945]), .Z(n14727) );
  XOR U15399 ( .A(n14726), .B(n14727), .Z(n14667) );
  AND U15400 ( .A(x[249]), .B(y[1921]), .Z(n14735) );
  XOR U15401 ( .A(o[154]), .B(n14735), .Z(n14681) );
  AND U15402 ( .A(x[250]), .B(y[1920]), .Z(n14680) );
  XOR U15403 ( .A(n14681), .B(n14680), .Z(n14683) );
  AND U15404 ( .A(x[224]), .B(y[1946]), .Z(n14682) );
  XOR U15405 ( .A(n14683), .B(n14682), .Z(n14666) );
  XOR U15406 ( .A(n14667), .B(n14666), .Z(n14669) );
  NAND U15407 ( .A(n14555), .B(n14554), .Z(n14559) );
  NAND U15408 ( .A(n14557), .B(n14556), .Z(n14558) );
  AND U15409 ( .A(n14559), .B(n14558), .Z(n14668) );
  XOR U15410 ( .A(n14669), .B(n14668), .Z(n14614) );
  XNOR U15411 ( .A(n14615), .B(n14614), .Z(n14657) );
  AND U15412 ( .A(x[245]), .B(y[1925]), .Z(n14565) );
  IV U15413 ( .A(n14565), .Z(n14718) );
  NANDN U15414 ( .A(n14718), .B(n14560), .Z(n14564) );
  NAND U15415 ( .A(n14562), .B(n14561), .Z(n14563) );
  NAND U15416 ( .A(n14564), .B(n14563), .Z(n14645) );
  XOR U15417 ( .A(n14719), .B(n14565), .Z(n14720) );
  AND U15418 ( .A(x[244]), .B(y[1926]), .Z(n14721) );
  XOR U15419 ( .A(n14720), .B(n14721), .Z(n14643) );
  AND U15420 ( .A(x[247]), .B(y[1923]), .Z(n14631) );
  XOR U15421 ( .A(n14630), .B(n14631), .Z(n14632) );
  AND U15422 ( .A(x[246]), .B(y[1924]), .Z(n14633) );
  XOR U15423 ( .A(n14632), .B(n14633), .Z(n14642) );
  XOR U15424 ( .A(n14643), .B(n14642), .Z(n14644) );
  XNOR U15425 ( .A(n14645), .B(n14644), .Z(n14655) );
  AND U15426 ( .A(x[228]), .B(y[1942]), .Z(n14636) );
  XOR U15427 ( .A(n14637), .B(n14636), .Z(n14639) );
  XOR U15428 ( .A(n14639), .B(n14638), .Z(n14619) );
  AND U15429 ( .A(x[227]), .B(y[1943]), .Z(n14710) );
  AND U15430 ( .A(x[243]), .B(y[1927]), .Z(n14711) );
  XOR U15431 ( .A(n14710), .B(n14711), .Z(n14712) );
  AND U15432 ( .A(x[235]), .B(y[1935]), .Z(n14713) );
  XOR U15433 ( .A(n14712), .B(n14713), .Z(n14618) );
  XOR U15434 ( .A(n14619), .B(n14618), .Z(n14621) );
  NAND U15435 ( .A(n14567), .B(n14566), .Z(n14571) );
  NAND U15436 ( .A(n14569), .B(n14568), .Z(n14570) );
  AND U15437 ( .A(n14571), .B(n14570), .Z(n14620) );
  XNOR U15438 ( .A(n14621), .B(n14620), .Z(n14654) );
  XOR U15439 ( .A(n14655), .B(n14654), .Z(n14656) );
  XOR U15440 ( .A(n14657), .B(n14656), .Z(n14688) );
  XNOR U15441 ( .A(n14689), .B(n14688), .Z(n14693) );
  NANDN U15442 ( .A(n14573), .B(n14572), .Z(n14577) );
  NANDN U15443 ( .A(n14575), .B(n14574), .Z(n14576) );
  NAND U15444 ( .A(n14577), .B(n14576), .Z(n14739) );
  NAND U15445 ( .A(n14579), .B(n14578), .Z(n14583) );
  NANDN U15446 ( .A(n14581), .B(n14580), .Z(n14582) );
  NAND U15447 ( .A(n14583), .B(n14582), .Z(n14737) );
  NAND U15448 ( .A(n14585), .B(n14584), .Z(n14589) );
  NANDN U15449 ( .A(n14587), .B(n14586), .Z(n14588) );
  NAND U15450 ( .A(n14589), .B(n14588), .Z(n14736) );
  XOR U15451 ( .A(n14737), .B(n14736), .Z(n14738) );
  XOR U15452 ( .A(n14739), .B(n14738), .Z(n14692) );
  XOR U15453 ( .A(n14693), .B(n14692), .Z(n14694) );
  XOR U15454 ( .A(n14695), .B(n14694), .Z(n14748) );
  XNOR U15455 ( .A(n14749), .B(n14748), .Z(n14751) );
  XOR U15456 ( .A(n14750), .B(n14751), .Z(n14611) );
  XOR U15457 ( .A(n14609), .B(n14608), .Z(n14610) );
  XOR U15458 ( .A(n14611), .B(n14610), .Z(n14754) );
  XNOR U15459 ( .A(n14755), .B(n14754), .Z(n14761) );
  NANDN U15460 ( .A(n14602), .B(n14601), .Z(n14606) );
  NANDN U15461 ( .A(n14604), .B(n14603), .Z(n14605) );
  AND U15462 ( .A(n14606), .B(n14605), .Z(n14759) );
  IV U15463 ( .A(n14759), .Z(n14758) );
  XOR U15464 ( .A(n14760), .B(n14758), .Z(n14607) );
  XNOR U15465 ( .A(n14761), .B(n14607), .Z(N315) );
  NAND U15466 ( .A(n14613), .B(n14612), .Z(n14617) );
  NAND U15467 ( .A(n14615), .B(n14614), .Z(n14616) );
  NAND U15468 ( .A(n14617), .B(n14616), .Z(n14895) );
  NAND U15469 ( .A(n14619), .B(n14618), .Z(n14623) );
  NAND U15470 ( .A(n14621), .B(n14620), .Z(n14622) );
  NAND U15471 ( .A(n14623), .B(n14622), .Z(n14893) );
  AND U15472 ( .A(n14625), .B(n14624), .Z(n14629) );
  NAND U15473 ( .A(n14627), .B(n14626), .Z(n14628) );
  NANDN U15474 ( .A(n14629), .B(n14628), .Z(n14791) );
  NAND U15475 ( .A(n14631), .B(n14630), .Z(n14635) );
  NAND U15476 ( .A(n14633), .B(n14632), .Z(n14634) );
  NAND U15477 ( .A(n14635), .B(n14634), .Z(n14790) );
  XOR U15478 ( .A(n14791), .B(n14790), .Z(n14792) );
  AND U15479 ( .A(n14637), .B(n14636), .Z(n14641) );
  NAND U15480 ( .A(n14639), .B(n14638), .Z(n14640) );
  NANDN U15481 ( .A(n14641), .B(n14640), .Z(n14804) );
  AND U15482 ( .A(x[224]), .B(y[1947]), .Z(n14882) );
  AND U15483 ( .A(x[251]), .B(y[1920]), .Z(n14881) );
  XOR U15484 ( .A(n14882), .B(n14881), .Z(n14884) );
  AND U15485 ( .A(x[250]), .B(y[1921]), .Z(n14872) );
  XOR U15486 ( .A(n14872), .B(o[155]), .Z(n14883) );
  XOR U15487 ( .A(n14884), .B(n14883), .Z(n14803) );
  AND U15488 ( .A(x[233]), .B(y[1938]), .Z(n14867) );
  AND U15489 ( .A(x[245]), .B(y[1926]), .Z(n14866) );
  XOR U15490 ( .A(n14867), .B(n14866), .Z(n14869) );
  AND U15491 ( .A(x[242]), .B(y[1929]), .Z(n14868) );
  XOR U15492 ( .A(n14869), .B(n14868), .Z(n14802) );
  XOR U15493 ( .A(n14803), .B(n14802), .Z(n14805) );
  XNOR U15494 ( .A(n14804), .B(n14805), .Z(n14793) );
  XOR U15495 ( .A(n14893), .B(n14894), .Z(n14896) );
  XOR U15496 ( .A(n14895), .B(n14896), .Z(n14914) );
  NAND U15497 ( .A(n14643), .B(n14642), .Z(n14647) );
  NAND U15498 ( .A(n14645), .B(n14644), .Z(n14646) );
  AND U15499 ( .A(n14647), .B(n14646), .Z(n14912) );
  NAND U15500 ( .A(n14649), .B(n14648), .Z(n14653) );
  NAND U15501 ( .A(n14651), .B(n14650), .Z(n14652) );
  AND U15502 ( .A(n14653), .B(n14652), .Z(n14911) );
  XOR U15503 ( .A(n14912), .B(n14911), .Z(n14913) );
  NAND U15504 ( .A(n14655), .B(n14654), .Z(n14659) );
  NAND U15505 ( .A(n14657), .B(n14656), .Z(n14658) );
  AND U15506 ( .A(n14659), .B(n14658), .Z(n14899) );
  NAND U15507 ( .A(n14661), .B(n14660), .Z(n14665) );
  NAND U15508 ( .A(n14663), .B(n14662), .Z(n14664) );
  NAND U15509 ( .A(n14665), .B(n14664), .Z(n14889) );
  NAND U15510 ( .A(n14667), .B(n14666), .Z(n14671) );
  NAND U15511 ( .A(n14669), .B(n14668), .Z(n14670) );
  NAND U15512 ( .A(n14671), .B(n14670), .Z(n14887) );
  AND U15513 ( .A(x[243]), .B(y[1928]), .Z(n14861) );
  AND U15514 ( .A(x[249]), .B(y[1922]), .Z(n14860) );
  XOR U15515 ( .A(n14861), .B(n14860), .Z(n14863) );
  AND U15516 ( .A(x[230]), .B(y[1941]), .Z(n14862) );
  XOR U15517 ( .A(n14863), .B(n14862), .Z(n14850) );
  AND U15518 ( .A(x[239]), .B(y[1932]), .Z(n14826) );
  AND U15519 ( .A(x[226]), .B(y[1945]), .Z(n14825) );
  XOR U15520 ( .A(n14826), .B(n14825), .Z(n14828) );
  AND U15521 ( .A(x[227]), .B(y[1944]), .Z(n14827) );
  XOR U15522 ( .A(n14828), .B(n14827), .Z(n14849) );
  XOR U15523 ( .A(n14850), .B(n14849), .Z(n14851) );
  NAND U15524 ( .A(x[240]), .B(y[1931]), .Z(n14808) );
  XOR U15525 ( .A(n14808), .B(n14672), .Z(n14811) );
  XOR U15526 ( .A(n14810), .B(n14811), .Z(n14822) );
  AND U15527 ( .A(y[1934]), .B(x[237]), .Z(n14674) );
  AND U15528 ( .A(y[1935]), .B(x[236]), .Z(n14673) );
  XOR U15529 ( .A(n14674), .B(n14673), .Z(n14821) );
  XNOR U15530 ( .A(n14851), .B(n14852), .Z(n14787) );
  AND U15531 ( .A(n14820), .B(n14675), .Z(n14679) );
  NAND U15532 ( .A(n14677), .B(n14676), .Z(n14678) );
  NANDN U15533 ( .A(n14679), .B(n14678), .Z(n14785) );
  NAND U15534 ( .A(n14681), .B(n14680), .Z(n14685) );
  NAND U15535 ( .A(n14683), .B(n14682), .Z(n14684) );
  NAND U15536 ( .A(n14685), .B(n14684), .Z(n14784) );
  XOR U15537 ( .A(n14785), .B(n14784), .Z(n14786) );
  XOR U15538 ( .A(n14787), .B(n14786), .Z(n14888) );
  XNOR U15539 ( .A(n14887), .B(n14888), .Z(n14890) );
  XNOR U15540 ( .A(n14899), .B(n14900), .Z(n14902) );
  NAND U15541 ( .A(n14687), .B(n14686), .Z(n14691) );
  NAND U15542 ( .A(n14689), .B(n14688), .Z(n14690) );
  AND U15543 ( .A(n14691), .B(n14690), .Z(n14901) );
  XOR U15544 ( .A(n14902), .B(n14901), .Z(n14772) );
  NAND U15545 ( .A(n14693), .B(n14692), .Z(n14697) );
  NAND U15546 ( .A(n14695), .B(n14694), .Z(n14696) );
  NAND U15547 ( .A(n14697), .B(n14696), .Z(n14774) );
  XOR U15548 ( .A(n14775), .B(n14774), .Z(n14769) );
  NAND U15549 ( .A(n14699), .B(n14698), .Z(n14703) );
  NAND U15550 ( .A(n14701), .B(n14700), .Z(n14702) );
  NAND U15551 ( .A(n14703), .B(n14702), .Z(n14778) );
  NAND U15552 ( .A(n14705), .B(n14704), .Z(n14709) );
  NAND U15553 ( .A(n14707), .B(n14706), .Z(n14708) );
  AND U15554 ( .A(n14709), .B(n14708), .Z(n14907) );
  NAND U15555 ( .A(n14711), .B(n14710), .Z(n14715) );
  NAND U15556 ( .A(n14713), .B(n14712), .Z(n14714) );
  NAND U15557 ( .A(n14715), .B(n14714), .Z(n14845) );
  AND U15558 ( .A(y[1923]), .B(x[248]), .Z(n14717) );
  NAND U15559 ( .A(y[1927]), .B(x[244]), .Z(n14716) );
  XNOR U15560 ( .A(n14717), .B(n14716), .Z(n14857) );
  AND U15561 ( .A(x[231]), .B(y[1940]), .Z(n14856) );
  XOR U15562 ( .A(n14857), .B(n14856), .Z(n14844) );
  AND U15563 ( .A(x[232]), .B(y[1939]), .Z(n14815) );
  AND U15564 ( .A(x[247]), .B(y[1924]), .Z(n14814) );
  XOR U15565 ( .A(n14815), .B(n14814), .Z(n14817) );
  AND U15566 ( .A(x[246]), .B(y[1925]), .Z(n14816) );
  XOR U15567 ( .A(n14817), .B(n14816), .Z(n14843) );
  XOR U15568 ( .A(n14844), .B(n14843), .Z(n14846) );
  XOR U15569 ( .A(n14845), .B(n14846), .Z(n14906) );
  ANDN U15570 ( .B(n14719), .A(n14718), .Z(n14723) );
  NAND U15571 ( .A(n14721), .B(n14720), .Z(n14722) );
  NANDN U15572 ( .A(n14723), .B(n14722), .Z(n14838) );
  NAND U15573 ( .A(n14725), .B(n14724), .Z(n14729) );
  NAND U15574 ( .A(n14727), .B(n14726), .Z(n14728) );
  NAND U15575 ( .A(n14729), .B(n14728), .Z(n14837) );
  XOR U15576 ( .A(n14838), .B(n14837), .Z(n14839) );
  AND U15577 ( .A(y[1940]), .B(x[232]), .Z(n14874) );
  NAND U15578 ( .A(n14874), .B(n14730), .Z(n14734) );
  NAND U15579 ( .A(n14732), .B(n14731), .Z(n14733) );
  NAND U15580 ( .A(n14734), .B(n14733), .Z(n14798) );
  AND U15581 ( .A(x[238]), .B(y[1933]), .Z(n14832) );
  AND U15582 ( .A(x[225]), .B(y[1946]), .Z(n14831) );
  XOR U15583 ( .A(n14832), .B(n14831), .Z(n14834) );
  AND U15584 ( .A(o[154]), .B(n14735), .Z(n14833) );
  XOR U15585 ( .A(n14834), .B(n14833), .Z(n14797) );
  AND U15586 ( .A(x[241]), .B(y[1930]), .Z(n14876) );
  AND U15587 ( .A(x[228]), .B(y[1943]), .Z(n14875) );
  XOR U15588 ( .A(n14876), .B(n14875), .Z(n14878) );
  AND U15589 ( .A(x[229]), .B(y[1942]), .Z(n14877) );
  XOR U15590 ( .A(n14878), .B(n14877), .Z(n14796) );
  XOR U15591 ( .A(n14797), .B(n14796), .Z(n14799) );
  XOR U15592 ( .A(n14798), .B(n14799), .Z(n14840) );
  XNOR U15593 ( .A(n14839), .B(n14840), .Z(n14905) );
  XNOR U15594 ( .A(n14907), .B(n14908), .Z(n14779) );
  XOR U15595 ( .A(n14778), .B(n14779), .Z(n14781) );
  NAND U15596 ( .A(n14737), .B(n14736), .Z(n14741) );
  NAND U15597 ( .A(n14739), .B(n14738), .Z(n14740) );
  AND U15598 ( .A(n14741), .B(n14740), .Z(n14780) );
  XNOR U15599 ( .A(n14781), .B(n14780), .Z(n14767) );
  NAND U15600 ( .A(n14743), .B(n14742), .Z(n14747) );
  NAND U15601 ( .A(n14745), .B(n14744), .Z(n14746) );
  AND U15602 ( .A(n14747), .B(n14746), .Z(n14766) );
  XOR U15603 ( .A(n14767), .B(n14766), .Z(n14768) );
  XOR U15604 ( .A(n14769), .B(n14768), .Z(n14921) );
  XNOR U15605 ( .A(n14921), .B(n14920), .Z(n14922) );
  XNOR U15606 ( .A(n14923), .B(n14922), .Z(n14919) );
  NAND U15607 ( .A(n14753), .B(n14752), .Z(n14757) );
  NAND U15608 ( .A(n14755), .B(n14754), .Z(n14756) );
  AND U15609 ( .A(n14757), .B(n14756), .Z(n14918) );
  OR U15610 ( .A(n14760), .B(n14758), .Z(n14764) );
  ANDN U15611 ( .B(n14760), .A(n14759), .Z(n14762) );
  OR U15612 ( .A(n14762), .B(n14761), .Z(n14763) );
  AND U15613 ( .A(n14764), .B(n14763), .Z(n14917) );
  XNOR U15614 ( .A(n14918), .B(n14917), .Z(n14765) );
  XNOR U15615 ( .A(n14919), .B(n14765), .Z(N316) );
  NAND U15616 ( .A(n14767), .B(n14766), .Z(n14771) );
  NAND U15617 ( .A(n14769), .B(n14768), .Z(n14770) );
  NAND U15618 ( .A(n14771), .B(n14770), .Z(n15088) );
  NANDN U15619 ( .A(n14773), .B(n14772), .Z(n14777) );
  NAND U15620 ( .A(n14775), .B(n14774), .Z(n14776) );
  NAND U15621 ( .A(n14777), .B(n14776), .Z(n15087) );
  XOR U15622 ( .A(n15088), .B(n15087), .Z(n15090) );
  NAND U15623 ( .A(n14779), .B(n14778), .Z(n14783) );
  NAND U15624 ( .A(n14781), .B(n14780), .Z(n14782) );
  AND U15625 ( .A(n14783), .B(n14782), .Z(n14927) );
  NAND U15626 ( .A(n14785), .B(n14784), .Z(n14789) );
  NAND U15627 ( .A(n14787), .B(n14786), .Z(n14788) );
  NAND U15628 ( .A(n14789), .B(n14788), .Z(n14951) );
  NAND U15629 ( .A(n14791), .B(n14790), .Z(n14795) );
  NANDN U15630 ( .A(n14793), .B(n14792), .Z(n14794) );
  NAND U15631 ( .A(n14795), .B(n14794), .Z(n15056) );
  NAND U15632 ( .A(n14797), .B(n14796), .Z(n14801) );
  NAND U15633 ( .A(n14799), .B(n14798), .Z(n14800) );
  NAND U15634 ( .A(n14801), .B(n14800), .Z(n15055) );
  NAND U15635 ( .A(n14803), .B(n14802), .Z(n14807) );
  NAND U15636 ( .A(n14805), .B(n14804), .Z(n14806) );
  NAND U15637 ( .A(n14807), .B(n14806), .Z(n15054) );
  XOR U15638 ( .A(n15055), .B(n15054), .Z(n15057) );
  XOR U15639 ( .A(n15056), .B(n15057), .Z(n14952) );
  XOR U15640 ( .A(n14951), .B(n14952), .Z(n14954) );
  NANDN U15641 ( .A(n14809), .B(n14808), .Z(n14813) );
  NAND U15642 ( .A(n14811), .B(n14810), .Z(n14812) );
  NAND U15643 ( .A(n14813), .B(n14812), .Z(n15032) );
  AND U15644 ( .A(x[231]), .B(y[1941]), .Z(n14999) );
  AND U15645 ( .A(x[236]), .B(y[1936]), .Z(n14998) );
  XOR U15646 ( .A(n14999), .B(n14998), .Z(n15001) );
  AND U15647 ( .A(x[235]), .B(y[1937]), .Z(n15000) );
  XOR U15648 ( .A(n15001), .B(n15000), .Z(n15031) );
  AND U15649 ( .A(x[251]), .B(y[1921]), .Z(n15010) );
  XOR U15650 ( .A(o[156]), .B(n15010), .Z(n15023) );
  AND U15651 ( .A(x[250]), .B(y[1922]), .Z(n15022) );
  XOR U15652 ( .A(n15023), .B(n15022), .Z(n15025) );
  AND U15653 ( .A(x[239]), .B(y[1933]), .Z(n15024) );
  XNOR U15654 ( .A(n15025), .B(n15024), .Z(n15030) );
  XOR U15655 ( .A(n15032), .B(n15033), .Z(n15061) );
  NAND U15656 ( .A(n14815), .B(n14814), .Z(n14819) );
  NAND U15657 ( .A(n14817), .B(n14816), .Z(n14818) );
  NAND U15658 ( .A(n14819), .B(n14818), .Z(n15038) );
  AND U15659 ( .A(x[241]), .B(y[1931]), .Z(n14964) );
  AND U15660 ( .A(x[246]), .B(y[1926]), .Z(n14963) );
  XOR U15661 ( .A(n14964), .B(n14963), .Z(n14966) );
  AND U15662 ( .A(x[228]), .B(y[1944]), .Z(n14965) );
  XOR U15663 ( .A(n14966), .B(n14965), .Z(n15037) );
  AND U15664 ( .A(x[230]), .B(y[1942]), .Z(n15173) );
  AND U15665 ( .A(x[243]), .B(y[1929]), .Z(n15011) );
  XOR U15666 ( .A(n15173), .B(n15011), .Z(n15013) );
  XOR U15667 ( .A(n15013), .B(n15012), .Z(n15036) );
  XOR U15668 ( .A(n15037), .B(n15036), .Z(n15039) );
  XOR U15669 ( .A(n15038), .B(n15039), .Z(n15060) );
  NAND U15670 ( .A(n15017), .B(n14820), .Z(n14824) );
  NANDN U15671 ( .A(n14822), .B(n14821), .Z(n14823) );
  NAND U15672 ( .A(n14824), .B(n14823), .Z(n14959) );
  NAND U15673 ( .A(n14826), .B(n14825), .Z(n14830) );
  NAND U15674 ( .A(n14828), .B(n14827), .Z(n14829) );
  NAND U15675 ( .A(n14830), .B(n14829), .Z(n14958) );
  NAND U15676 ( .A(n14832), .B(n14831), .Z(n14836) );
  NAND U15677 ( .A(n14834), .B(n14833), .Z(n14835) );
  NAND U15678 ( .A(n14836), .B(n14835), .Z(n14957) );
  XOR U15679 ( .A(n14958), .B(n14957), .Z(n14960) );
  XOR U15680 ( .A(n14959), .B(n14960), .Z(n15062) );
  XOR U15681 ( .A(n15063), .B(n15062), .Z(n14953) );
  XNOR U15682 ( .A(n14954), .B(n14953), .Z(n14948) );
  NAND U15683 ( .A(n14838), .B(n14837), .Z(n14842) );
  NAND U15684 ( .A(n14840), .B(n14839), .Z(n14841) );
  NAND U15685 ( .A(n14842), .B(n14841), .Z(n15044) );
  NAND U15686 ( .A(n14844), .B(n14843), .Z(n14848) );
  NAND U15687 ( .A(n14846), .B(n14845), .Z(n14847) );
  NAND U15688 ( .A(n14848), .B(n14847), .Z(n15043) );
  NAND U15689 ( .A(n14850), .B(n14849), .Z(n14854) );
  NANDN U15690 ( .A(n14852), .B(n14851), .Z(n14853) );
  NAND U15691 ( .A(n14854), .B(n14853), .Z(n15042) );
  XOR U15692 ( .A(n15043), .B(n15042), .Z(n15045) );
  XOR U15693 ( .A(n15044), .B(n15045), .Z(n14946) );
  AND U15694 ( .A(x[248]), .B(y[1927]), .Z(n15452) );
  AND U15695 ( .A(x[244]), .B(y[1923]), .Z(n14855) );
  NAND U15696 ( .A(n15452), .B(n14855), .Z(n14859) );
  NAND U15697 ( .A(n14857), .B(n14856), .Z(n14858) );
  NAND U15698 ( .A(n14859), .B(n14858), .Z(n15080) );
  AND U15699 ( .A(x[249]), .B(y[1923]), .Z(n14994) );
  XOR U15700 ( .A(n14995), .B(n14994), .Z(n14993) );
  AND U15701 ( .A(x[225]), .B(y[1947]), .Z(n14992) );
  XOR U15702 ( .A(n14993), .B(n14992), .Z(n15079) );
  AND U15703 ( .A(x[240]), .B(y[1932]), .Z(n14987) );
  AND U15704 ( .A(x[248]), .B(y[1924]), .Z(n14986) );
  XOR U15705 ( .A(n14987), .B(n14986), .Z(n14989) );
  AND U15706 ( .A(x[226]), .B(y[1946]), .Z(n14988) );
  XOR U15707 ( .A(n14989), .B(n14988), .Z(n15078) );
  XOR U15708 ( .A(n15079), .B(n15078), .Z(n15081) );
  XOR U15709 ( .A(n15080), .B(n15081), .Z(n15051) );
  NAND U15710 ( .A(n14861), .B(n14860), .Z(n14865) );
  NAND U15711 ( .A(n14863), .B(n14862), .Z(n14864) );
  NAND U15712 ( .A(n14865), .B(n14864), .Z(n15074) );
  AND U15713 ( .A(x[227]), .B(y[1945]), .Z(n15016) );
  XOR U15714 ( .A(n15017), .B(n15016), .Z(n15019) );
  AND U15715 ( .A(x[247]), .B(y[1925]), .Z(n15018) );
  XOR U15716 ( .A(n15019), .B(n15018), .Z(n15073) );
  AND U15717 ( .A(x[229]), .B(y[1943]), .Z(n15005) );
  AND U15718 ( .A(x[245]), .B(y[1927]), .Z(n15004) );
  XOR U15719 ( .A(n15005), .B(n15004), .Z(n15007) );
  AND U15720 ( .A(x[244]), .B(y[1928]), .Z(n15006) );
  XOR U15721 ( .A(n15007), .B(n15006), .Z(n15072) );
  XOR U15722 ( .A(n15073), .B(n15072), .Z(n15075) );
  XOR U15723 ( .A(n15074), .B(n15075), .Z(n15049) );
  NAND U15724 ( .A(n14867), .B(n14866), .Z(n14871) );
  NAND U15725 ( .A(n14869), .B(n14868), .Z(n14870) );
  NAND U15726 ( .A(n14871), .B(n14870), .Z(n14982) );
  AND U15727 ( .A(n14872), .B(o[155]), .Z(n14972) );
  AND U15728 ( .A(x[224]), .B(y[1948]), .Z(n14970) );
  AND U15729 ( .A(x[252]), .B(y[1920]), .Z(n14969) );
  XOR U15730 ( .A(n14970), .B(n14969), .Z(n14971) );
  XOR U15731 ( .A(n14972), .B(n14971), .Z(n14981) );
  NAND U15732 ( .A(y[1938]), .B(x[234]), .Z(n14873) );
  XNOR U15733 ( .A(n14874), .B(n14873), .Z(n14977) );
  AND U15734 ( .A(x[233]), .B(y[1939]), .Z(n14976) );
  XOR U15735 ( .A(n14977), .B(n14976), .Z(n14980) );
  XOR U15736 ( .A(n14981), .B(n14980), .Z(n14983) );
  XOR U15737 ( .A(n14982), .B(n14983), .Z(n15069) );
  NAND U15738 ( .A(n14876), .B(n14875), .Z(n14880) );
  NAND U15739 ( .A(n14878), .B(n14877), .Z(n14879) );
  NAND U15740 ( .A(n14880), .B(n14879), .Z(n15067) );
  NAND U15741 ( .A(n14882), .B(n14881), .Z(n14886) );
  NAND U15742 ( .A(n14884), .B(n14883), .Z(n14885) );
  NAND U15743 ( .A(n14886), .B(n14885), .Z(n15066) );
  XOR U15744 ( .A(n15067), .B(n15066), .Z(n15068) );
  XNOR U15745 ( .A(n15069), .B(n15068), .Z(n15048) );
  XNOR U15746 ( .A(n14948), .B(n14947), .Z(n14941) );
  NAND U15747 ( .A(n14888), .B(n14887), .Z(n14892) );
  NANDN U15748 ( .A(n14890), .B(n14889), .Z(n14891) );
  NAND U15749 ( .A(n14892), .B(n14891), .Z(n14940) );
  NAND U15750 ( .A(n14894), .B(n14893), .Z(n14898) );
  NAND U15751 ( .A(n14896), .B(n14895), .Z(n14897) );
  NAND U15752 ( .A(n14898), .B(n14897), .Z(n14939) );
  XNOR U15753 ( .A(n14940), .B(n14939), .Z(n14942) );
  XNOR U15754 ( .A(n14927), .B(n14928), .Z(n14929) );
  NANDN U15755 ( .A(n14900), .B(n14899), .Z(n14904) );
  NAND U15756 ( .A(n14902), .B(n14901), .Z(n14903) );
  NAND U15757 ( .A(n14904), .B(n14903), .Z(n14935) );
  NANDN U15758 ( .A(n14906), .B(n14905), .Z(n14910) );
  NANDN U15759 ( .A(n14908), .B(n14907), .Z(n14909) );
  AND U15760 ( .A(n14910), .B(n14909), .Z(n14934) );
  NAND U15761 ( .A(n14912), .B(n14911), .Z(n14916) );
  NANDN U15762 ( .A(n14914), .B(n14913), .Z(n14915) );
  AND U15763 ( .A(n14916), .B(n14915), .Z(n14933) );
  XOR U15764 ( .A(n14934), .B(n14933), .Z(n14936) );
  XNOR U15765 ( .A(n14935), .B(n14936), .Z(n14930) );
  XNOR U15766 ( .A(n15090), .B(n15089), .Z(n15086) );
  NANDN U15767 ( .A(n14921), .B(n14920), .Z(n14925) );
  NAND U15768 ( .A(n14923), .B(n14922), .Z(n14924) );
  AND U15769 ( .A(n14925), .B(n14924), .Z(n15085) );
  XOR U15770 ( .A(n15084), .B(n15085), .Z(n14926) );
  XNOR U15771 ( .A(n15086), .B(n14926), .Z(N317) );
  NANDN U15772 ( .A(n14928), .B(n14927), .Z(n14932) );
  NANDN U15773 ( .A(n14930), .B(n14929), .Z(n14931) );
  NAND U15774 ( .A(n14932), .B(n14931), .Z(n15103) );
  NAND U15775 ( .A(n14934), .B(n14933), .Z(n14938) );
  NAND U15776 ( .A(n14936), .B(n14935), .Z(n14937) );
  NAND U15777 ( .A(n14938), .B(n14937), .Z(n15101) );
  NAND U15778 ( .A(n14940), .B(n14939), .Z(n14944) );
  NANDN U15779 ( .A(n14942), .B(n14941), .Z(n14943) );
  NAND U15780 ( .A(n14944), .B(n14943), .Z(n15107) );
  NANDN U15781 ( .A(n14946), .B(n14945), .Z(n14950) );
  NAND U15782 ( .A(n14948), .B(n14947), .Z(n14949) );
  AND U15783 ( .A(n14950), .B(n14949), .Z(n15108) );
  XOR U15784 ( .A(n15107), .B(n15108), .Z(n15110) );
  NAND U15785 ( .A(n14952), .B(n14951), .Z(n14956) );
  NAND U15786 ( .A(n14954), .B(n14953), .Z(n14955) );
  NAND U15787 ( .A(n14956), .B(n14955), .Z(n15125) );
  NAND U15788 ( .A(n14958), .B(n14957), .Z(n14962) );
  NAND U15789 ( .A(n14960), .B(n14959), .Z(n14961) );
  AND U15790 ( .A(n14962), .B(n14961), .Z(n15230) );
  NAND U15791 ( .A(n14964), .B(n14963), .Z(n14968) );
  NAND U15792 ( .A(n14966), .B(n14965), .Z(n14967) );
  NAND U15793 ( .A(n14968), .B(n14967), .Z(n15268) );
  NAND U15794 ( .A(n14970), .B(n14969), .Z(n14974) );
  NAND U15795 ( .A(n14972), .B(n14971), .Z(n14973) );
  NAND U15796 ( .A(n14974), .B(n14973), .Z(n15267) );
  XOR U15797 ( .A(n15268), .B(n15267), .Z(n15269) );
  AND U15798 ( .A(y[1940]), .B(x[234]), .Z(n15265) );
  NAND U15799 ( .A(n14975), .B(n15265), .Z(n14979) );
  NAND U15800 ( .A(n14977), .B(n14976), .Z(n14978) );
  NAND U15801 ( .A(n14979), .B(n14978), .Z(n15236) );
  AND U15802 ( .A(x[236]), .B(y[1937]), .Z(n15311) );
  AND U15803 ( .A(x[225]), .B(y[1948]), .Z(n15149) );
  XOR U15804 ( .A(n15311), .B(n15149), .Z(n15151) );
  AND U15805 ( .A(x[246]), .B(y[1927]), .Z(n15150) );
  XOR U15806 ( .A(n15151), .B(n15150), .Z(n15235) );
  AND U15807 ( .A(x[239]), .B(y[1934]), .Z(n15154) );
  XOR U15808 ( .A(n15235), .B(n15234), .Z(n15237) );
  XNOR U15809 ( .A(n15236), .B(n15237), .Z(n15270) );
  NAND U15810 ( .A(n14981), .B(n14980), .Z(n14985) );
  NAND U15811 ( .A(n14983), .B(n14982), .Z(n14984) );
  AND U15812 ( .A(n14985), .B(n14984), .Z(n15228) );
  XNOR U15813 ( .A(n15230), .B(n15231), .Z(n15225) );
  NAND U15814 ( .A(n14987), .B(n14986), .Z(n14991) );
  NAND U15815 ( .A(n14989), .B(n14988), .Z(n14990) );
  NAND U15816 ( .A(n14991), .B(n14990), .Z(n15241) );
  AND U15817 ( .A(n14993), .B(n14992), .Z(n14997) );
  NAND U15818 ( .A(n14995), .B(n14994), .Z(n14996) );
  NANDN U15819 ( .A(n14997), .B(n14996), .Z(n15240) );
  XOR U15820 ( .A(n15241), .B(n15240), .Z(n15242) );
  NAND U15821 ( .A(n14999), .B(n14998), .Z(n15003) );
  NAND U15822 ( .A(n15001), .B(n15000), .Z(n15002) );
  NAND U15823 ( .A(n15003), .B(n15002), .Z(n15188) );
  AND U15824 ( .A(x[235]), .B(y[1938]), .Z(n15170) );
  AND U15825 ( .A(x[227]), .B(y[1946]), .Z(n15168) );
  AND U15826 ( .A(x[241]), .B(y[1932]), .Z(n15167) );
  XOR U15827 ( .A(n15168), .B(n15167), .Z(n15169) );
  XOR U15828 ( .A(n15170), .B(n15169), .Z(n15187) );
  AND U15829 ( .A(x[247]), .B(y[1926]), .Z(n15164) );
  AND U15830 ( .A(x[237]), .B(y[1936]), .Z(n15162) );
  AND U15831 ( .A(x[248]), .B(y[1925]), .Z(n15367) );
  XOR U15832 ( .A(n15162), .B(n15367), .Z(n15163) );
  XOR U15833 ( .A(n15164), .B(n15163), .Z(n15186) );
  XOR U15834 ( .A(n15187), .B(n15186), .Z(n15189) );
  XNOR U15835 ( .A(n15188), .B(n15189), .Z(n15243) );
  NAND U15836 ( .A(n15005), .B(n15004), .Z(n15009) );
  NAND U15837 ( .A(n15007), .B(n15006), .Z(n15008) );
  NAND U15838 ( .A(n15009), .B(n15008), .Z(n15182) );
  AND U15839 ( .A(n15010), .B(o[156]), .Z(n15195) );
  AND U15840 ( .A(x[240]), .B(y[1933]), .Z(n15193) );
  AND U15841 ( .A(x[251]), .B(y[1922]), .Z(n15192) );
  XOR U15842 ( .A(n15193), .B(n15192), .Z(n15194) );
  XOR U15843 ( .A(n15195), .B(n15194), .Z(n15181) );
  AND U15844 ( .A(x[226]), .B(y[1947]), .Z(n15204) );
  XOR U15845 ( .A(n15207), .B(n15206), .Z(n15180) );
  XOR U15846 ( .A(n15181), .B(n15180), .Z(n15183) );
  XOR U15847 ( .A(n15182), .B(n15183), .Z(n15132) );
  NAND U15848 ( .A(n15173), .B(n15011), .Z(n15015) );
  NAND U15849 ( .A(n15013), .B(n15012), .Z(n15014) );
  NAND U15850 ( .A(n15015), .B(n15014), .Z(n15249) );
  AND U15851 ( .A(x[249]), .B(y[1924]), .Z(n15146) );
  AND U15852 ( .A(x[250]), .B(y[1923]), .Z(n15143) );
  XOR U15853 ( .A(n15144), .B(n15143), .Z(n15145) );
  XOR U15854 ( .A(n15146), .B(n15145), .Z(n15247) );
  AND U15855 ( .A(x[252]), .B(y[1921]), .Z(n15161) );
  XOR U15856 ( .A(o[157]), .B(n15161), .Z(n15260) );
  AND U15857 ( .A(x[224]), .B(y[1949]), .Z(n15258) );
  AND U15858 ( .A(x[253]), .B(y[1920]), .Z(n15257) );
  XOR U15859 ( .A(n15258), .B(n15257), .Z(n15259) );
  XNOR U15860 ( .A(n15260), .B(n15259), .Z(n15246) );
  XOR U15861 ( .A(n15249), .B(n15248), .Z(n15131) );
  NAND U15862 ( .A(n15017), .B(n15016), .Z(n15021) );
  NAND U15863 ( .A(n15019), .B(n15018), .Z(n15020) );
  NAND U15864 ( .A(n15021), .B(n15020), .Z(n15211) );
  NAND U15865 ( .A(n15023), .B(n15022), .Z(n15027) );
  NAND U15866 ( .A(n15025), .B(n15024), .Z(n15026) );
  NAND U15867 ( .A(n15027), .B(n15026), .Z(n15210) );
  XOR U15868 ( .A(n15211), .B(n15210), .Z(n15213) );
  AND U15869 ( .A(x[232]), .B(y[1941]), .Z(n15175) );
  AND U15870 ( .A(x[230]), .B(y[1943]), .Z(n15029) );
  AND U15871 ( .A(y[1942]), .B(x[231]), .Z(n15028) );
  XOR U15872 ( .A(n15029), .B(n15028), .Z(n15174) );
  XOR U15873 ( .A(n15175), .B(n15174), .Z(n15252) );
  AND U15874 ( .A(x[233]), .B(y[1940]), .Z(n15468) );
  XOR U15875 ( .A(n15252), .B(n15468), .Z(n15254) );
  AND U15876 ( .A(x[229]), .B(y[1944]), .Z(n15201) );
  AND U15877 ( .A(x[228]), .B(y[1945]), .Z(n15199) );
  AND U15878 ( .A(x[234]), .B(y[1939]), .Z(n15198) );
  XOR U15879 ( .A(n15199), .B(n15198), .Z(n15200) );
  XOR U15880 ( .A(n15201), .B(n15200), .Z(n15253) );
  XOR U15881 ( .A(n15254), .B(n15253), .Z(n15212) );
  XOR U15882 ( .A(n15213), .B(n15212), .Z(n15138) );
  NANDN U15883 ( .A(n15031), .B(n15030), .Z(n15035) );
  NAND U15884 ( .A(n15033), .B(n15032), .Z(n15034) );
  NAND U15885 ( .A(n15035), .B(n15034), .Z(n15137) );
  XNOR U15886 ( .A(n15139), .B(n15140), .Z(n15223) );
  NAND U15887 ( .A(n15037), .B(n15036), .Z(n15041) );
  NAND U15888 ( .A(n15039), .B(n15038), .Z(n15040) );
  NAND U15889 ( .A(n15041), .B(n15040), .Z(n15222) );
  XOR U15890 ( .A(n15125), .B(n15126), .Z(n15128) );
  NAND U15891 ( .A(n15043), .B(n15042), .Z(n15047) );
  NAND U15892 ( .A(n15045), .B(n15044), .Z(n15046) );
  NAND U15893 ( .A(n15047), .B(n15046), .Z(n15119) );
  NANDN U15894 ( .A(n15049), .B(n15048), .Z(n15053) );
  NANDN U15895 ( .A(n15051), .B(n15050), .Z(n15052) );
  AND U15896 ( .A(n15053), .B(n15052), .Z(n15120) );
  XOR U15897 ( .A(n15119), .B(n15120), .Z(n15121) );
  NAND U15898 ( .A(n15055), .B(n15054), .Z(n15059) );
  NAND U15899 ( .A(n15057), .B(n15056), .Z(n15058) );
  NAND U15900 ( .A(n15059), .B(n15058), .Z(n15115) );
  NANDN U15901 ( .A(n15061), .B(n15060), .Z(n15065) );
  NAND U15902 ( .A(n15063), .B(n15062), .Z(n15064) );
  NAND U15903 ( .A(n15065), .B(n15064), .Z(n15113) );
  NAND U15904 ( .A(n15067), .B(n15066), .Z(n15071) );
  NAND U15905 ( .A(n15069), .B(n15068), .Z(n15070) );
  NAND U15906 ( .A(n15071), .B(n15070), .Z(n15218) );
  NAND U15907 ( .A(n15073), .B(n15072), .Z(n15077) );
  NAND U15908 ( .A(n15075), .B(n15074), .Z(n15076) );
  NAND U15909 ( .A(n15077), .B(n15076), .Z(n15217) );
  NAND U15910 ( .A(n15079), .B(n15078), .Z(n15083) );
  NAND U15911 ( .A(n15081), .B(n15080), .Z(n15082) );
  NAND U15912 ( .A(n15083), .B(n15082), .Z(n15216) );
  XNOR U15913 ( .A(n15217), .B(n15216), .Z(n15219) );
  XOR U15914 ( .A(n15113), .B(n15114), .Z(n15116) );
  XOR U15915 ( .A(n15115), .B(n15116), .Z(n15122) );
  XNOR U15916 ( .A(n15121), .B(n15122), .Z(n15127) );
  XOR U15917 ( .A(n15128), .B(n15127), .Z(n15109) );
  XOR U15918 ( .A(n15110), .B(n15109), .Z(n15102) );
  XOR U15919 ( .A(n15101), .B(n15102), .Z(n15104) );
  XOR U15920 ( .A(n15103), .B(n15104), .Z(n15097) );
  NAND U15921 ( .A(n15088), .B(n15087), .Z(n15092) );
  NAND U15922 ( .A(n15090), .B(n15089), .Z(n15091) );
  AND U15923 ( .A(n15092), .B(n15091), .Z(n15096) );
  IV U15924 ( .A(n15096), .Z(n15094) );
  XOR U15925 ( .A(n15095), .B(n15094), .Z(n15093) );
  XNOR U15926 ( .A(n15097), .B(n15093), .Z(N318) );
  NANDN U15927 ( .A(n15094), .B(n15095), .Z(n15100) );
  NOR U15928 ( .A(n15096), .B(n15095), .Z(n15098) );
  OR U15929 ( .A(n15098), .B(n15097), .Z(n15099) );
  AND U15930 ( .A(n15100), .B(n15099), .Z(n15276) );
  NAND U15931 ( .A(n15102), .B(n15101), .Z(n15106) );
  NAND U15932 ( .A(n15104), .B(n15103), .Z(n15105) );
  AND U15933 ( .A(n15106), .B(n15105), .Z(n15275) );
  XNOR U15934 ( .A(n15276), .B(n15275), .Z(n15274) );
  NAND U15935 ( .A(n15108), .B(n15107), .Z(n15112) );
  NAND U15936 ( .A(n15110), .B(n15109), .Z(n15111) );
  NAND U15937 ( .A(n15112), .B(n15111), .Z(n15562) );
  NANDN U15938 ( .A(n15114), .B(n15113), .Z(n15118) );
  NANDN U15939 ( .A(n15116), .B(n15115), .Z(n15117) );
  AND U15940 ( .A(n15118), .B(n15117), .Z(n15568) );
  NAND U15941 ( .A(n15120), .B(n15119), .Z(n15124) );
  NANDN U15942 ( .A(n15122), .B(n15121), .Z(n15123) );
  AND U15943 ( .A(n15124), .B(n15123), .Z(n15566) );
  NAND U15944 ( .A(n15126), .B(n15125), .Z(n15130) );
  NAND U15945 ( .A(n15128), .B(n15127), .Z(n15129) );
  AND U15946 ( .A(n15130), .B(n15129), .Z(n15565) );
  XOR U15947 ( .A(n15566), .B(n15565), .Z(n15567) );
  XOR U15948 ( .A(n15568), .B(n15567), .Z(n15559) );
  NANDN U15949 ( .A(n15132), .B(n15131), .Z(n15136) );
  NANDN U15950 ( .A(n15134), .B(n15133), .Z(n15135) );
  AND U15951 ( .A(n15136), .B(n15135), .Z(n15547) );
  NANDN U15952 ( .A(n15138), .B(n15137), .Z(n15142) );
  NANDN U15953 ( .A(n15140), .B(n15139), .Z(n15141) );
  AND U15954 ( .A(n15142), .B(n15141), .Z(n15540) );
  AND U15955 ( .A(n15144), .B(n15143), .Z(n15148) );
  NAND U15956 ( .A(n15146), .B(n15145), .Z(n15147) );
  NANDN U15957 ( .A(n15148), .B(n15147), .Z(n15400) );
  AND U15958 ( .A(n15311), .B(n15149), .Z(n15153) );
  NAND U15959 ( .A(n15151), .B(n15150), .Z(n15152) );
  NANDN U15960 ( .A(n15153), .B(n15152), .Z(n15403) );
  NANDN U15961 ( .A(n15316), .B(n15154), .Z(n15158) );
  NANDN U15962 ( .A(n15156), .B(n15155), .Z(n15157) );
  AND U15963 ( .A(n15158), .B(n15157), .Z(n15292) );
  AND U15964 ( .A(x[247]), .B(y[1927]), .Z(n15366) );
  AND U15965 ( .A(y[1926]), .B(x[248]), .Z(n15160) );
  AND U15966 ( .A(y[1925]), .B(x[249]), .Z(n15159) );
  XOR U15967 ( .A(n15160), .B(n15159), .Z(n15365) );
  XOR U15968 ( .A(n15366), .B(n15365), .Z(n15294) );
  AND U15969 ( .A(n15161), .B(o[157]), .Z(n15326) );
  AND U15970 ( .A(x[252]), .B(y[1922]), .Z(n15328) );
  AND U15971 ( .A(x[240]), .B(y[1934]), .Z(n15327) );
  XOR U15972 ( .A(n15328), .B(n15327), .Z(n15325) );
  XNOR U15973 ( .A(n15326), .B(n15325), .Z(n15293) );
  XNOR U15974 ( .A(n15292), .B(n15291), .Z(n15402) );
  XOR U15975 ( .A(n15403), .B(n15402), .Z(n15401) );
  XOR U15976 ( .A(n15400), .B(n15401), .Z(n15522) );
  NAND U15977 ( .A(n15162), .B(n15367), .Z(n15166) );
  NAND U15978 ( .A(n15164), .B(n15163), .Z(n15165) );
  NAND U15979 ( .A(n15166), .B(n15165), .Z(n15288) );
  NAND U15980 ( .A(n15168), .B(n15167), .Z(n15172) );
  NAND U15981 ( .A(n15170), .B(n15169), .Z(n15171) );
  AND U15982 ( .A(n15172), .B(n15171), .Z(n15383) );
  AND U15983 ( .A(x[224]), .B(y[1950]), .Z(n15472) );
  AND U15984 ( .A(x[253]), .B(y[1921]), .Z(n15449) );
  XOR U15985 ( .A(o[158]), .B(n15449), .Z(n15474) );
  AND U15986 ( .A(x[254]), .B(y[1920]), .Z(n15473) );
  XOR U15987 ( .A(n15474), .B(n15473), .Z(n15471) );
  XOR U15988 ( .A(n15472), .B(n15471), .Z(n15385) );
  AND U15989 ( .A(x[244]), .B(y[1930]), .Z(n15353) );
  XOR U15990 ( .A(n15354), .B(n15353), .Z(n15352) );
  AND U15991 ( .A(x[232]), .B(y[1942]), .Z(n15351) );
  XNOR U15992 ( .A(n15352), .B(n15351), .Z(n15384) );
  XNOR U15993 ( .A(n15383), .B(n15382), .Z(n15287) );
  XOR U15994 ( .A(n15288), .B(n15287), .Z(n15285) );
  AND U15995 ( .A(x[231]), .B(y[1943]), .Z(n15318) );
  NAND U15996 ( .A(n15173), .B(n15318), .Z(n15177) );
  NAND U15997 ( .A(n15175), .B(n15174), .Z(n15176) );
  AND U15998 ( .A(n15177), .B(n15176), .Z(n15303) );
  AND U15999 ( .A(y[1929]), .B(x[245]), .Z(n15179) );
  AND U16000 ( .A(y[1928]), .B(x[246]), .Z(n15178) );
  XOR U16001 ( .A(n15179), .B(n15178), .Z(n15317) );
  XOR U16002 ( .A(n15318), .B(n15317), .Z(n15306) );
  AND U16003 ( .A(x[241]), .B(y[1933]), .Z(n15346) );
  AND U16004 ( .A(x[226]), .B(y[1948]), .Z(n15348) );
  AND U16005 ( .A(x[250]), .B(y[1924]), .Z(n15347) );
  XOR U16006 ( .A(n15348), .B(n15347), .Z(n15345) );
  XNOR U16007 ( .A(n15346), .B(n15345), .Z(n15305) );
  XNOR U16008 ( .A(n15303), .B(n15304), .Z(n15286) );
  NAND U16009 ( .A(n15181), .B(n15180), .Z(n15185) );
  NAND U16010 ( .A(n15183), .B(n15182), .Z(n15184) );
  NAND U16011 ( .A(n15185), .B(n15184), .Z(n15523) );
  XOR U16012 ( .A(n15524), .B(n15523), .Z(n15521) );
  XOR U16013 ( .A(n15522), .B(n15521), .Z(n15542) );
  NAND U16014 ( .A(n15187), .B(n15186), .Z(n15191) );
  NAND U16015 ( .A(n15189), .B(n15188), .Z(n15190) );
  NAND U16016 ( .A(n15191), .B(n15190), .Z(n15517) );
  NAND U16017 ( .A(n15193), .B(n15192), .Z(n15197) );
  NAND U16018 ( .A(n15195), .B(n15194), .Z(n15196) );
  NAND U16019 ( .A(n15197), .B(n15196), .Z(n15394) );
  NAND U16020 ( .A(n15199), .B(n15198), .Z(n15203) );
  NAND U16021 ( .A(n15201), .B(n15200), .Z(n15202) );
  NAND U16022 ( .A(n15203), .B(n15202), .Z(n15397) );
  AND U16023 ( .A(x[230]), .B(y[1944]), .Z(n15417) );
  AND U16024 ( .A(x[229]), .B(y[1945]), .Z(n15419) );
  AND U16025 ( .A(x[243]), .B(y[1931]), .Z(n15418) );
  XOR U16026 ( .A(n15419), .B(n15418), .Z(n15416) );
  XNOR U16027 ( .A(n15417), .B(n15416), .Z(n15376) );
  AND U16028 ( .A(x[228]), .B(y[1946]), .Z(n15411) );
  AND U16029 ( .A(x[227]), .B(y[1947]), .Z(n15413) );
  AND U16030 ( .A(x[242]), .B(y[1932]), .Z(n15412) );
  XOR U16031 ( .A(n15413), .B(n15412), .Z(n15410) );
  XOR U16032 ( .A(n15411), .B(n15410), .Z(n15379) );
  NANDN U16033 ( .A(n15205), .B(n15204), .Z(n15209) );
  NAND U16034 ( .A(n15207), .B(n15206), .Z(n15208) );
  AND U16035 ( .A(n15209), .B(n15208), .Z(n15378) );
  XOR U16036 ( .A(n15376), .B(n15377), .Z(n15396) );
  XOR U16037 ( .A(n15397), .B(n15396), .Z(n15395) );
  XOR U16038 ( .A(n15394), .B(n15395), .Z(n15518) );
  XOR U16039 ( .A(n15517), .B(n15518), .Z(n15516) );
  NAND U16040 ( .A(n15211), .B(n15210), .Z(n15215) );
  NAND U16041 ( .A(n15213), .B(n15212), .Z(n15214) );
  NAND U16042 ( .A(n15215), .B(n15214), .Z(n15515) );
  XOR U16043 ( .A(n15516), .B(n15515), .Z(n15541) );
  XOR U16044 ( .A(n15542), .B(n15541), .Z(n15539) );
  XOR U16045 ( .A(n15540), .B(n15539), .Z(n15549) );
  NAND U16046 ( .A(n15217), .B(n15216), .Z(n15221) );
  NANDN U16047 ( .A(n15219), .B(n15218), .Z(n15220) );
  AND U16048 ( .A(n15221), .B(n15220), .Z(n15548) );
  NANDN U16049 ( .A(n15223), .B(n15222), .Z(n15227) );
  NANDN U16050 ( .A(n15225), .B(n15224), .Z(n15226) );
  NAND U16051 ( .A(n15227), .B(n15226), .Z(n15535) );
  NANDN U16052 ( .A(n15229), .B(n15228), .Z(n15233) );
  NANDN U16053 ( .A(n15231), .B(n15230), .Z(n15232) );
  AND U16054 ( .A(n15233), .B(n15232), .Z(n15279) );
  NAND U16055 ( .A(n15235), .B(n15234), .Z(n15239) );
  NAND U16056 ( .A(n15237), .B(n15236), .Z(n15238) );
  AND U16057 ( .A(n15239), .B(n15238), .Z(n15506) );
  NAND U16058 ( .A(n15241), .B(n15240), .Z(n15245) );
  NANDN U16059 ( .A(n15243), .B(n15242), .Z(n15244) );
  AND U16060 ( .A(n15245), .B(n15244), .Z(n15505) );
  XOR U16061 ( .A(n15506), .B(n15505), .Z(n15504) );
  NANDN U16062 ( .A(n15247), .B(n15246), .Z(n15251) );
  OR U16063 ( .A(n15249), .B(n15248), .Z(n15250) );
  NAND U16064 ( .A(n15251), .B(n15250), .Z(n15503) );
  XOR U16065 ( .A(n15504), .B(n15503), .Z(n15282) );
  NAND U16066 ( .A(n15252), .B(n15468), .Z(n15256) );
  NAND U16067 ( .A(n15254), .B(n15253), .Z(n15255) );
  AND U16068 ( .A(n15256), .B(n15255), .Z(n15499) );
  NAND U16069 ( .A(n15258), .B(n15257), .Z(n15262) );
  NAND U16070 ( .A(n15260), .B(n15259), .Z(n15261) );
  NAND U16071 ( .A(n15262), .B(n15261), .Z(n15297) );
  AND U16072 ( .A(y[1938]), .B(x[236]), .Z(n15263) );
  XOR U16073 ( .A(n15264), .B(n15263), .Z(n15312) );
  XOR U16074 ( .A(n15313), .B(n15312), .Z(n15466) );
  AND U16075 ( .A(y[1941]), .B(x[233]), .Z(n15266) );
  XOR U16076 ( .A(n15266), .B(n15265), .Z(n15465) );
  XOR U16077 ( .A(n15466), .B(n15465), .Z(n15300) );
  AND U16078 ( .A(x[251]), .B(y[1923]), .Z(n15362) );
  AND U16079 ( .A(x[225]), .B(y[1949]), .Z(n15361) );
  XOR U16080 ( .A(n15362), .B(n15361), .Z(n15359) );
  XOR U16081 ( .A(n15360), .B(n15359), .Z(n15299) );
  XOR U16082 ( .A(n15300), .B(n15299), .Z(n15298) );
  XOR U16083 ( .A(n15297), .B(n15298), .Z(n15500) );
  NAND U16084 ( .A(n15268), .B(n15267), .Z(n15272) );
  NANDN U16085 ( .A(n15270), .B(n15269), .Z(n15271) );
  AND U16086 ( .A(n15272), .B(n15271), .Z(n15497) );
  XNOR U16087 ( .A(n15498), .B(n15497), .Z(n15281) );
  XNOR U16088 ( .A(n15279), .B(n15280), .Z(n15536) );
  XOR U16089 ( .A(n15535), .B(n15536), .Z(n15533) );
  XOR U16090 ( .A(n15534), .B(n15533), .Z(n15560) );
  XOR U16091 ( .A(n15562), .B(n15561), .Z(n15273) );
  XNOR U16092 ( .A(n15274), .B(n15273), .Z(N319) );
  NAND U16093 ( .A(n15274), .B(n15273), .Z(n15278) );
  NANDN U16094 ( .A(n15276), .B(n15275), .Z(n15277) );
  AND U16095 ( .A(n15278), .B(n15277), .Z(n15558) );
  NANDN U16096 ( .A(n15280), .B(n15279), .Z(n15284) );
  NANDN U16097 ( .A(n15282), .B(n15281), .Z(n15283) );
  AND U16098 ( .A(n15284), .B(n15283), .Z(n15532) );
  NANDN U16099 ( .A(n15286), .B(n15285), .Z(n15290) );
  NAND U16100 ( .A(n15288), .B(n15287), .Z(n15289) );
  AND U16101 ( .A(n15290), .B(n15289), .Z(n15514) );
  NAND U16102 ( .A(n15292), .B(n15291), .Z(n15296) );
  NANDN U16103 ( .A(n15294), .B(n15293), .Z(n15295) );
  AND U16104 ( .A(n15296), .B(n15295), .Z(n15496) );
  NAND U16105 ( .A(n15298), .B(n15297), .Z(n15302) );
  NAND U16106 ( .A(n15300), .B(n15299), .Z(n15301) );
  AND U16107 ( .A(n15302), .B(n15301), .Z(n15310) );
  NANDN U16108 ( .A(n15304), .B(n15303), .Z(n15308) );
  NANDN U16109 ( .A(n15306), .B(n15305), .Z(n15307) );
  NAND U16110 ( .A(n15308), .B(n15307), .Z(n15309) );
  XNOR U16111 ( .A(n15310), .B(n15309), .Z(n15494) );
  AND U16112 ( .A(n15311), .B(n15430), .Z(n15315) );
  AND U16113 ( .A(n15313), .B(n15312), .Z(n15314) );
  NOR U16114 ( .A(n15315), .B(n15314), .Z(n15322) );
  AND U16115 ( .A(x[246]), .B(y[1929]), .Z(n15450) );
  NANDN U16116 ( .A(n15316), .B(n15450), .Z(n15320) );
  NAND U16117 ( .A(n15318), .B(n15317), .Z(n15319) );
  AND U16118 ( .A(n15320), .B(n15319), .Z(n15321) );
  XNOR U16119 ( .A(n15322), .B(n15321), .Z(n15393) );
  AND U16120 ( .A(y[1937]), .B(x[238]), .Z(n15324) );
  NAND U16121 ( .A(y[1942]), .B(x[233]), .Z(n15323) );
  XNOR U16122 ( .A(n15324), .B(n15323), .Z(n15344) );
  AND U16123 ( .A(y[1923]), .B(x[252]), .Z(n15342) );
  NAND U16124 ( .A(n15326), .B(n15325), .Z(n15330) );
  NAND U16125 ( .A(n15328), .B(n15327), .Z(n15329) );
  AND U16126 ( .A(n15330), .B(n15329), .Z(n15338) );
  AND U16127 ( .A(y[1940]), .B(x[235]), .Z(n15332) );
  NAND U16128 ( .A(y[1939]), .B(x[236]), .Z(n15331) );
  XNOR U16129 ( .A(n15332), .B(n15331), .Z(n15336) );
  AND U16130 ( .A(y[1921]), .B(x[254]), .Z(n15334) );
  NAND U16131 ( .A(y[1922]), .B(x[253]), .Z(n15333) );
  XNOR U16132 ( .A(n15334), .B(n15333), .Z(n15335) );
  XNOR U16133 ( .A(n15336), .B(n15335), .Z(n15337) );
  XNOR U16134 ( .A(n15338), .B(n15337), .Z(n15339) );
  XNOR U16135 ( .A(n15340), .B(n15339), .Z(n15341) );
  XNOR U16136 ( .A(n15342), .B(n15341), .Z(n15343) );
  XOR U16137 ( .A(n15344), .B(n15343), .Z(n15375) );
  NAND U16138 ( .A(n15346), .B(n15345), .Z(n15350) );
  NAND U16139 ( .A(n15348), .B(n15347), .Z(n15349) );
  AND U16140 ( .A(n15350), .B(n15349), .Z(n15358) );
  NAND U16141 ( .A(n15352), .B(n15351), .Z(n15356) );
  NAND U16142 ( .A(n15354), .B(n15353), .Z(n15355) );
  NAND U16143 ( .A(n15356), .B(n15355), .Z(n15357) );
  XNOR U16144 ( .A(n15358), .B(n15357), .Z(n15373) );
  NAND U16145 ( .A(n15360), .B(n15359), .Z(n15364) );
  NAND U16146 ( .A(n15362), .B(n15361), .Z(n15363) );
  AND U16147 ( .A(n15364), .B(n15363), .Z(n15371) );
  NAND U16148 ( .A(n15366), .B(n15365), .Z(n15369) );
  AND U16149 ( .A(x[249]), .B(y[1926]), .Z(n15451) );
  NAND U16150 ( .A(n15367), .B(n15451), .Z(n15368) );
  NAND U16151 ( .A(n15369), .B(n15368), .Z(n15370) );
  XNOR U16152 ( .A(n15371), .B(n15370), .Z(n15372) );
  XNOR U16153 ( .A(n15373), .B(n15372), .Z(n15374) );
  XNOR U16154 ( .A(n15375), .B(n15374), .Z(n15391) );
  NANDN U16155 ( .A(n15377), .B(n15376), .Z(n15381) );
  NANDN U16156 ( .A(n15379), .B(n15378), .Z(n15380) );
  AND U16157 ( .A(n15381), .B(n15380), .Z(n15389) );
  NAND U16158 ( .A(n15383), .B(n15382), .Z(n15387) );
  NANDN U16159 ( .A(n15385), .B(n15384), .Z(n15386) );
  NAND U16160 ( .A(n15387), .B(n15386), .Z(n15388) );
  XNOR U16161 ( .A(n15389), .B(n15388), .Z(n15390) );
  XOR U16162 ( .A(n15391), .B(n15390), .Z(n15392) );
  XNOR U16163 ( .A(n15393), .B(n15392), .Z(n15409) );
  NAND U16164 ( .A(n15395), .B(n15394), .Z(n15399) );
  NAND U16165 ( .A(n15397), .B(n15396), .Z(n15398) );
  AND U16166 ( .A(n15399), .B(n15398), .Z(n15407) );
  NAND U16167 ( .A(n15401), .B(n15400), .Z(n15405) );
  NAND U16168 ( .A(n15403), .B(n15402), .Z(n15404) );
  NAND U16169 ( .A(n15405), .B(n15404), .Z(n15406) );
  XNOR U16170 ( .A(n15407), .B(n15406), .Z(n15408) );
  XOR U16171 ( .A(n15409), .B(n15408), .Z(n15492) );
  NAND U16172 ( .A(n15411), .B(n15410), .Z(n15415) );
  NAND U16173 ( .A(n15413), .B(n15412), .Z(n15414) );
  AND U16174 ( .A(n15415), .B(n15414), .Z(n15423) );
  NAND U16175 ( .A(n15417), .B(n15416), .Z(n15421) );
  NAND U16176 ( .A(n15419), .B(n15418), .Z(n15420) );
  NAND U16177 ( .A(n15421), .B(n15420), .Z(n15422) );
  XNOR U16178 ( .A(n15423), .B(n15422), .Z(n15490) );
  AND U16179 ( .A(y[1945]), .B(x[230]), .Z(n15425) );
  NAND U16180 ( .A(y[1944]), .B(x[231]), .Z(n15424) );
  XNOR U16181 ( .A(n15425), .B(n15424), .Z(n15429) );
  AND U16182 ( .A(y[1946]), .B(x[229]), .Z(n15427) );
  NAND U16183 ( .A(y[1933]), .B(x[242]), .Z(n15426) );
  XNOR U16184 ( .A(n15427), .B(n15426), .Z(n15428) );
  XOR U16185 ( .A(n15429), .B(n15428), .Z(n15432) );
  AND U16186 ( .A(x[234]), .B(y[1941]), .Z(n15467) );
  XNOR U16187 ( .A(n15430), .B(n15467), .Z(n15431) );
  XNOR U16188 ( .A(n15432), .B(n15431), .Z(n15448) );
  AND U16189 ( .A(y[1928]), .B(x[247]), .Z(n15434) );
  NAND U16190 ( .A(y[1934]), .B(x[241]), .Z(n15433) );
  XNOR U16191 ( .A(n15434), .B(n15433), .Z(n15438) );
  AND U16192 ( .A(y[1924]), .B(x[251]), .Z(n15436) );
  NAND U16193 ( .A(y[1930]), .B(x[245]), .Z(n15435) );
  XNOR U16194 ( .A(n15436), .B(n15435), .Z(n15437) );
  XOR U16195 ( .A(n15438), .B(n15437), .Z(n15446) );
  AND U16196 ( .A(y[1948]), .B(x[227]), .Z(n15440) );
  NAND U16197 ( .A(y[1947]), .B(x[228]), .Z(n15439) );
  XNOR U16198 ( .A(n15440), .B(n15439), .Z(n15444) );
  AND U16199 ( .A(y[1920]), .B(x[255]), .Z(n15442) );
  NAND U16200 ( .A(y[1949]), .B(x[226]), .Z(n15441) );
  XNOR U16201 ( .A(n15442), .B(n15441), .Z(n15443) );
  XNOR U16202 ( .A(n15444), .B(n15443), .Z(n15445) );
  XNOR U16203 ( .A(n15446), .B(n15445), .Z(n15447) );
  XOR U16204 ( .A(n15448), .B(n15447), .Z(n15464) );
  AND U16205 ( .A(y[1931]), .B(x[244]), .Z(n15458) );
  AND U16206 ( .A(n15449), .B(o[158]), .Z(n15456) );
  XOR U16207 ( .A(n15450), .B(o[159]), .Z(n15454) );
  XNOR U16208 ( .A(n15452), .B(n15451), .Z(n15453) );
  XNOR U16209 ( .A(n15454), .B(n15453), .Z(n15455) );
  XNOR U16210 ( .A(n15456), .B(n15455), .Z(n15457) );
  XNOR U16211 ( .A(n15458), .B(n15457), .Z(n15462) );
  AND U16212 ( .A(y[1932]), .B(x[243]), .Z(n15460) );
  NAND U16213 ( .A(y[1943]), .B(x[232]), .Z(n15459) );
  XNOR U16214 ( .A(n15460), .B(n15459), .Z(n15461) );
  XNOR U16215 ( .A(n15462), .B(n15461), .Z(n15463) );
  XNOR U16216 ( .A(n15464), .B(n15463), .Z(n15480) );
  NAND U16217 ( .A(n15466), .B(n15465), .Z(n15470) );
  NAND U16218 ( .A(n15468), .B(n15467), .Z(n15469) );
  AND U16219 ( .A(n15470), .B(n15469), .Z(n15478) );
  NAND U16220 ( .A(n15472), .B(n15471), .Z(n15476) );
  NAND U16221 ( .A(n15474), .B(n15473), .Z(n15475) );
  NAND U16222 ( .A(n15476), .B(n15475), .Z(n15477) );
  XNOR U16223 ( .A(n15478), .B(n15477), .Z(n15479) );
  XOR U16224 ( .A(n15480), .B(n15479), .Z(n15488) );
  AND U16225 ( .A(y[1935]), .B(x[240]), .Z(n15482) );
  NAND U16226 ( .A(y[1951]), .B(x[224]), .Z(n15481) );
  XNOR U16227 ( .A(n15482), .B(n15481), .Z(n15486) );
  AND U16228 ( .A(y[1950]), .B(x[225]), .Z(n15484) );
  NAND U16229 ( .A(y[1925]), .B(x[250]), .Z(n15483) );
  XNOR U16230 ( .A(n15484), .B(n15483), .Z(n15485) );
  XNOR U16231 ( .A(n15486), .B(n15485), .Z(n15487) );
  XNOR U16232 ( .A(n15488), .B(n15487), .Z(n15489) );
  XNOR U16233 ( .A(n15490), .B(n15489), .Z(n15491) );
  XNOR U16234 ( .A(n15492), .B(n15491), .Z(n15493) );
  XNOR U16235 ( .A(n15494), .B(n15493), .Z(n15495) );
  XNOR U16236 ( .A(n15496), .B(n15495), .Z(n15512) );
  NAND U16237 ( .A(n15498), .B(n15497), .Z(n15502) );
  NANDN U16238 ( .A(n15500), .B(n15499), .Z(n15501) );
  AND U16239 ( .A(n15502), .B(n15501), .Z(n15510) );
  NAND U16240 ( .A(n15504), .B(n15503), .Z(n15508) );
  NAND U16241 ( .A(n15506), .B(n15505), .Z(n15507) );
  NAND U16242 ( .A(n15508), .B(n15507), .Z(n15509) );
  XNOR U16243 ( .A(n15510), .B(n15509), .Z(n15511) );
  XNOR U16244 ( .A(n15512), .B(n15511), .Z(n15513) );
  XNOR U16245 ( .A(n15514), .B(n15513), .Z(n15530) );
  NAND U16246 ( .A(n15516), .B(n15515), .Z(n15520) );
  NAND U16247 ( .A(n15518), .B(n15517), .Z(n15519) );
  AND U16248 ( .A(n15520), .B(n15519), .Z(n15528) );
  NAND U16249 ( .A(n15522), .B(n15521), .Z(n15526) );
  NAND U16250 ( .A(n15524), .B(n15523), .Z(n15525) );
  NAND U16251 ( .A(n15526), .B(n15525), .Z(n15527) );
  XNOR U16252 ( .A(n15528), .B(n15527), .Z(n15529) );
  XNOR U16253 ( .A(n15530), .B(n15529), .Z(n15531) );
  XNOR U16254 ( .A(n15532), .B(n15531), .Z(n15556) );
  NAND U16255 ( .A(n15534), .B(n15533), .Z(n15538) );
  NAND U16256 ( .A(n15536), .B(n15535), .Z(n15537) );
  AND U16257 ( .A(n15538), .B(n15537), .Z(n15546) );
  NAND U16258 ( .A(n15540), .B(n15539), .Z(n15544) );
  NAND U16259 ( .A(n15542), .B(n15541), .Z(n15543) );
  NAND U16260 ( .A(n15544), .B(n15543), .Z(n15545) );
  XNOR U16261 ( .A(n15546), .B(n15545), .Z(n15554) );
  ANDN U16262 ( .B(n15548), .A(n15547), .Z(n15550) );
  NANDN U16263 ( .A(n15550), .B(n15549), .Z(n15551) );
  NAND U16264 ( .A(n15552), .B(n15551), .Z(n15553) );
  XNOR U16265 ( .A(n15554), .B(n15553), .Z(n15555) );
  XNOR U16266 ( .A(n15556), .B(n15555), .Z(n15557) );
  XNOR U16267 ( .A(n15558), .B(n15557), .Z(n15574) );
  ANDN U16268 ( .B(n15560), .A(n15559), .Z(n15564) );
  ANDN U16269 ( .B(n15562), .A(n15561), .Z(n15563) );
  NOR U16270 ( .A(n15564), .B(n15563), .Z(n15572) );
  NAND U16271 ( .A(n15566), .B(n15565), .Z(n15570) );
  NAND U16272 ( .A(n15568), .B(n15567), .Z(n15569) );
  AND U16273 ( .A(n15570), .B(n15569), .Z(n15571) );
  XNOR U16274 ( .A(n15572), .B(n15571), .Z(n15573) );
  XNOR U16275 ( .A(n15574), .B(n15573), .Z(N320) );
  AND U16276 ( .A(x[224]), .B(y[1952]), .Z(n16225) );
  XOR U16277 ( .A(n16225), .B(o[160]), .Z(N353) );
  AND U16278 ( .A(x[225]), .B(y[1952]), .Z(n15583) );
  AND U16279 ( .A(x[224]), .B(y[1953]), .Z(n15582) );
  XNOR U16280 ( .A(n15582), .B(o[161]), .Z(n15575) );
  XNOR U16281 ( .A(n15583), .B(n15575), .Z(n15577) );
  NAND U16282 ( .A(n16225), .B(o[160]), .Z(n15576) );
  XNOR U16283 ( .A(n15577), .B(n15576), .Z(N354) );
  NANDN U16284 ( .A(n15583), .B(n15575), .Z(n15579) );
  NAND U16285 ( .A(n15577), .B(n15576), .Z(n15578) );
  AND U16286 ( .A(n15579), .B(n15578), .Z(n15589) );
  AND U16287 ( .A(x[224]), .B(y[1954]), .Z(n15596) );
  XNOR U16288 ( .A(n15596), .B(o[162]), .Z(n15588) );
  XNOR U16289 ( .A(n15589), .B(n15588), .Z(n15591) );
  AND U16290 ( .A(y[1952]), .B(x[226]), .Z(n15581) );
  NAND U16291 ( .A(y[1953]), .B(x[225]), .Z(n15580) );
  XNOR U16292 ( .A(n15581), .B(n15580), .Z(n15585) );
  AND U16293 ( .A(n15582), .B(o[161]), .Z(n15584) );
  XNOR U16294 ( .A(n15585), .B(n15584), .Z(n15590) );
  XNOR U16295 ( .A(n15591), .B(n15590), .Z(N355) );
  NAND U16296 ( .A(x[226]), .B(y[1953]), .Z(n15603) );
  NANDN U16297 ( .A(n15603), .B(n15583), .Z(n15587) );
  NAND U16298 ( .A(n15585), .B(n15584), .Z(n15586) );
  AND U16299 ( .A(n15587), .B(n15586), .Z(n15609) );
  NANDN U16300 ( .A(n15589), .B(n15588), .Z(n15593) );
  NAND U16301 ( .A(n15591), .B(n15590), .Z(n15592) );
  AND U16302 ( .A(n15593), .B(n15592), .Z(n15608) );
  XNOR U16303 ( .A(n15609), .B(n15608), .Z(n15611) );
  AND U16304 ( .A(x[225]), .B(y[1954]), .Z(n15713) );
  XOR U16305 ( .A(n15713), .B(n15605), .Z(n15607) );
  AND U16306 ( .A(y[1952]), .B(x[227]), .Z(n15595) );
  NAND U16307 ( .A(y[1955]), .B(x[224]), .Z(n15594) );
  XNOR U16308 ( .A(n15595), .B(n15594), .Z(n15597) );
  NAND U16309 ( .A(n15596), .B(o[162]), .Z(n15598) );
  XOR U16310 ( .A(n15607), .B(n15606), .Z(n15610) );
  XOR U16311 ( .A(n15611), .B(n15610), .Z(N356) );
  AND U16312 ( .A(y[1955]), .B(x[227]), .Z(n15653) );
  NAND U16313 ( .A(n16225), .B(n15653), .Z(n15600) );
  NANDN U16314 ( .A(n15598), .B(n15597), .Z(n15599) );
  AND U16315 ( .A(n15600), .B(n15599), .Z(n15635) );
  AND U16316 ( .A(y[1956]), .B(x[224]), .Z(n15602) );
  NAND U16317 ( .A(y[1952]), .B(x[228]), .Z(n15601) );
  XNOR U16318 ( .A(n15602), .B(n15601), .Z(n15626) );
  ANDN U16319 ( .B(o[163]), .A(n15603), .Z(n15625) );
  XOR U16320 ( .A(n15626), .B(n15625), .Z(n15633) );
  AND U16321 ( .A(y[1954]), .B(x[226]), .Z(n15748) );
  NAND U16322 ( .A(y[1955]), .B(x[225]), .Z(n15604) );
  XNOR U16323 ( .A(n15748), .B(n15604), .Z(n15622) );
  NAND U16324 ( .A(x[227]), .B(y[1953]), .Z(n15619) );
  XOR U16325 ( .A(n15622), .B(n15621), .Z(n15632) );
  XOR U16326 ( .A(n15633), .B(n15632), .Z(n15634) );
  XOR U16327 ( .A(n15635), .B(n15634), .Z(n15631) );
  NANDN U16328 ( .A(n15609), .B(n15608), .Z(n15613) );
  NAND U16329 ( .A(n15611), .B(n15610), .Z(n15612) );
  NAND U16330 ( .A(n15613), .B(n15612), .Z(n15630) );
  XOR U16331 ( .A(n15629), .B(n15630), .Z(n15614) );
  XNOR U16332 ( .A(n15631), .B(n15614), .Z(N357) );
  AND U16333 ( .A(y[1954]), .B(x[227]), .Z(n15616) );
  NAND U16334 ( .A(y[1956]), .B(x[225]), .Z(n15615) );
  XNOR U16335 ( .A(n15616), .B(n15615), .Z(n15640) );
  AND U16336 ( .A(x[228]), .B(y[1953]), .Z(n15651) );
  XOR U16337 ( .A(n15651), .B(o[165]), .Z(n15639) );
  XNOR U16338 ( .A(n15640), .B(n15639), .Z(n15643) );
  NAND U16339 ( .A(x[226]), .B(y[1955]), .Z(n15721) );
  AND U16340 ( .A(y[1952]), .B(x[229]), .Z(n15618) );
  NAND U16341 ( .A(y[1957]), .B(x[224]), .Z(n15617) );
  XNOR U16342 ( .A(n15618), .B(n15617), .Z(n15646) );
  ANDN U16343 ( .B(o[164]), .A(n15619), .Z(n15645) );
  XOR U16344 ( .A(n15646), .B(n15645), .Z(n15644) );
  XOR U16345 ( .A(n15721), .B(n15644), .Z(n15620) );
  XOR U16346 ( .A(n15643), .B(n15620), .Z(n15665) );
  NANDN U16347 ( .A(n15721), .B(n15713), .Z(n15624) );
  NAND U16348 ( .A(n15622), .B(n15621), .Z(n15623) );
  NAND U16349 ( .A(n15624), .B(n15623), .Z(n15663) );
  AND U16350 ( .A(x[228]), .B(y[1956]), .Z(n16419) );
  NAND U16351 ( .A(n16419), .B(n16225), .Z(n15628) );
  NAND U16352 ( .A(n15626), .B(n15625), .Z(n15627) );
  NAND U16353 ( .A(n15628), .B(n15627), .Z(n15662) );
  XOR U16354 ( .A(n15663), .B(n15662), .Z(n15664) );
  XNOR U16355 ( .A(n15665), .B(n15664), .Z(n15658) );
  NAND U16356 ( .A(n15633), .B(n15632), .Z(n15637) );
  NANDN U16357 ( .A(n15635), .B(n15634), .Z(n15636) );
  NAND U16358 ( .A(n15637), .B(n15636), .Z(n15656) );
  IV U16359 ( .A(n15656), .Z(n15655) );
  XOR U16360 ( .A(n15657), .B(n15655), .Z(n15638) );
  XNOR U16361 ( .A(n15658), .B(n15638), .Z(N358) );
  AND U16362 ( .A(x[227]), .B(y[1956]), .Z(n15722) );
  NAND U16363 ( .A(n15722), .B(n15713), .Z(n15642) );
  NAND U16364 ( .A(n15640), .B(n15639), .Z(n15641) );
  NAND U16365 ( .A(n15642), .B(n15641), .Z(n15700) );
  XOR U16366 ( .A(n15700), .B(n15701), .Z(n15703) );
  AND U16367 ( .A(x[229]), .B(y[1957]), .Z(n15888) );
  NAND U16368 ( .A(n16225), .B(n15888), .Z(n15648) );
  NAND U16369 ( .A(n15646), .B(n15645), .Z(n15647) );
  AND U16370 ( .A(n15648), .B(n15647), .Z(n15670) );
  AND U16371 ( .A(y[1952]), .B(x[230]), .Z(n15650) );
  NAND U16372 ( .A(y[1958]), .B(x[224]), .Z(n15649) );
  XNOR U16373 ( .A(n15650), .B(n15649), .Z(n15676) );
  NAND U16374 ( .A(n15651), .B(o[165]), .Z(n15677) );
  NAND U16375 ( .A(y[1956]), .B(x[226]), .Z(n15652) );
  XNOR U16376 ( .A(n15653), .B(n15652), .Z(n15681) );
  AND U16377 ( .A(y[1957]), .B(x[225]), .Z(n15931) );
  NAND U16378 ( .A(y[1954]), .B(x[228]), .Z(n15654) );
  XNOR U16379 ( .A(n15931), .B(n15654), .Z(n15685) );
  AND U16380 ( .A(x[229]), .B(y[1953]), .Z(n15692) );
  XOR U16381 ( .A(o[166]), .B(n15692), .Z(n15684) );
  XOR U16382 ( .A(n15685), .B(n15684), .Z(n15680) );
  XOR U16383 ( .A(n15681), .B(n15680), .Z(n15671) );
  XOR U16384 ( .A(n15672), .B(n15671), .Z(n15702) );
  XOR U16385 ( .A(n15703), .B(n15702), .Z(n15696) );
  OR U16386 ( .A(n15657), .B(n15655), .Z(n15661) );
  ANDN U16387 ( .B(n15657), .A(n15656), .Z(n15659) );
  OR U16388 ( .A(n15659), .B(n15658), .Z(n15660) );
  AND U16389 ( .A(n15661), .B(n15660), .Z(n15694) );
  NAND U16390 ( .A(n15663), .B(n15662), .Z(n15667) );
  NAND U16391 ( .A(n15665), .B(n15664), .Z(n15666) );
  AND U16392 ( .A(n15667), .B(n15666), .Z(n15695) );
  IV U16393 ( .A(n15695), .Z(n15693) );
  XOR U16394 ( .A(n15694), .B(n15693), .Z(n15668) );
  XNOR U16395 ( .A(n15696), .B(n15668), .Z(N359) );
  NANDN U16396 ( .A(n15670), .B(n15669), .Z(n15674) );
  NAND U16397 ( .A(n15672), .B(n15671), .Z(n15673) );
  AND U16398 ( .A(n15674), .B(n15673), .Z(n15741) );
  AND U16399 ( .A(y[1954]), .B(x[229]), .Z(n15800) );
  NAND U16400 ( .A(y[1958]), .B(x[225]), .Z(n15675) );
  XNOR U16401 ( .A(n15800), .B(n15675), .Z(n15715) );
  NAND U16402 ( .A(x[230]), .B(y[1953]), .Z(n15719) );
  XOR U16403 ( .A(n15715), .B(n15714), .Z(n15733) );
  AND U16404 ( .A(x[230]), .B(y[1958]), .Z(n15951) );
  NAND U16405 ( .A(n16225), .B(n15951), .Z(n15679) );
  NANDN U16406 ( .A(n15677), .B(n15676), .Z(n15678) );
  AND U16407 ( .A(n15679), .B(n15678), .Z(n15732) );
  NANDN U16408 ( .A(n15721), .B(n15722), .Z(n15683) );
  NAND U16409 ( .A(n15681), .B(n15680), .Z(n15682) );
  NAND U16410 ( .A(n15683), .B(n15682), .Z(n15735) );
  AND U16411 ( .A(x[228]), .B(y[1957]), .Z(n16230) );
  NAND U16412 ( .A(n16230), .B(n15713), .Z(n15687) );
  NAND U16413 ( .A(n15685), .B(n15684), .Z(n15686) );
  AND U16414 ( .A(n15687), .B(n15686), .Z(n15710) );
  AND U16415 ( .A(y[1957]), .B(x[226]), .Z(n15689) );
  NAND U16416 ( .A(y[1955]), .B(x[228]), .Z(n15688) );
  XNOR U16417 ( .A(n15689), .B(n15688), .Z(n15723) );
  XNOR U16418 ( .A(n15723), .B(n15722), .Z(n15708) );
  AND U16419 ( .A(y[1952]), .B(x[231]), .Z(n15691) );
  NAND U16420 ( .A(y[1959]), .B(x[224]), .Z(n15690) );
  XNOR U16421 ( .A(n15691), .B(n15690), .Z(n15727) );
  AND U16422 ( .A(o[166]), .B(n15692), .Z(n15726) );
  XNOR U16423 ( .A(n15727), .B(n15726), .Z(n15707) );
  XOR U16424 ( .A(n15708), .B(n15707), .Z(n15709) );
  XOR U16425 ( .A(n15710), .B(n15709), .Z(n15738) );
  XOR U16426 ( .A(n15739), .B(n15738), .Z(n15740) );
  XNOR U16427 ( .A(n15741), .B(n15740), .Z(n15746) );
  NANDN U16428 ( .A(n15693), .B(n15694), .Z(n15699) );
  NOR U16429 ( .A(n15695), .B(n15694), .Z(n15697) );
  OR U16430 ( .A(n15697), .B(n15696), .Z(n15698) );
  AND U16431 ( .A(n15699), .B(n15698), .Z(n15745) );
  NAND U16432 ( .A(n15701), .B(n15700), .Z(n15705) );
  NAND U16433 ( .A(n15703), .B(n15702), .Z(n15704) );
  AND U16434 ( .A(n15705), .B(n15704), .Z(n15744) );
  XOR U16435 ( .A(n15745), .B(n15744), .Z(n15706) );
  XNOR U16436 ( .A(n15746), .B(n15706), .Z(N360) );
  NAND U16437 ( .A(n15708), .B(n15707), .Z(n15712) );
  NAND U16438 ( .A(n15710), .B(n15709), .Z(n15711) );
  AND U16439 ( .A(n15712), .B(n15711), .Z(n15781) );
  AND U16440 ( .A(x[229]), .B(y[1958]), .Z(n15880) );
  NAND U16441 ( .A(n15880), .B(n15713), .Z(n15717) );
  NAND U16442 ( .A(n15715), .B(n15714), .Z(n15716) );
  NAND U16443 ( .A(n15717), .B(n15716), .Z(n15779) );
  AND U16444 ( .A(y[1955]), .B(x[229]), .Z(n16361) );
  NAND U16445 ( .A(y[1959]), .B(x[225]), .Z(n15718) );
  XNOR U16446 ( .A(n16361), .B(n15718), .Z(n15769) );
  ANDN U16447 ( .B(o[167]), .A(n15719), .Z(n15768) );
  XNOR U16448 ( .A(n15769), .B(n15768), .Z(n15753) );
  NAND U16449 ( .A(x[227]), .B(y[1957]), .Z(n16543) );
  AND U16450 ( .A(x[230]), .B(y[1954]), .Z(n15720) );
  AND U16451 ( .A(y[1958]), .B(x[226]), .Z(n16624) );
  XOR U16452 ( .A(n15720), .B(n16624), .Z(n15749) );
  XOR U16453 ( .A(n16419), .B(n15749), .Z(n15752) );
  XOR U16454 ( .A(n15753), .B(n15754), .Z(n15778) );
  XOR U16455 ( .A(n15779), .B(n15778), .Z(n15780) );
  XOR U16456 ( .A(n15781), .B(n15780), .Z(n15787) );
  NANDN U16457 ( .A(n15721), .B(n16230), .Z(n15725) );
  NAND U16458 ( .A(n15723), .B(n15722), .Z(n15724) );
  NAND U16459 ( .A(n15725), .B(n15724), .Z(n15775) );
  AND U16460 ( .A(x[231]), .B(y[1959]), .Z(n16104) );
  NAND U16461 ( .A(n16225), .B(n16104), .Z(n15729) );
  NAND U16462 ( .A(n15727), .B(n15726), .Z(n15728) );
  NAND U16463 ( .A(n15729), .B(n15728), .Z(n15773) );
  AND U16464 ( .A(y[1952]), .B(x[232]), .Z(n15731) );
  NAND U16465 ( .A(y[1960]), .B(x[224]), .Z(n15730) );
  XNOR U16466 ( .A(n15731), .B(n15730), .Z(n15759) );
  AND U16467 ( .A(x[231]), .B(y[1953]), .Z(n15764) );
  XOR U16468 ( .A(o[168]), .B(n15764), .Z(n15758) );
  XOR U16469 ( .A(n15759), .B(n15758), .Z(n15772) );
  XOR U16470 ( .A(n15773), .B(n15772), .Z(n15774) );
  XNOR U16471 ( .A(n15775), .B(n15774), .Z(n15785) );
  NANDN U16472 ( .A(n15733), .B(n15732), .Z(n15737) );
  NANDN U16473 ( .A(n15735), .B(n15734), .Z(n15736) );
  NAND U16474 ( .A(n15737), .B(n15736), .Z(n15784) );
  XOR U16475 ( .A(n15785), .B(n15784), .Z(n15786) );
  XOR U16476 ( .A(n15787), .B(n15786), .Z(n15792) );
  NAND U16477 ( .A(n15739), .B(n15738), .Z(n15743) );
  NAND U16478 ( .A(n15741), .B(n15740), .Z(n15742) );
  NAND U16479 ( .A(n15743), .B(n15742), .Z(n15790) );
  XOR U16480 ( .A(n15790), .B(n15791), .Z(n15747) );
  XNOR U16481 ( .A(n15792), .B(n15747), .Z(N361) );
  NAND U16482 ( .A(n15951), .B(n15748), .Z(n15751) );
  NAND U16483 ( .A(n16419), .B(n15749), .Z(n15750) );
  NAND U16484 ( .A(n15751), .B(n15750), .Z(n15794) );
  NANDN U16485 ( .A(n15752), .B(n16543), .Z(n15756) );
  NANDN U16486 ( .A(n15754), .B(n15753), .Z(n15755) );
  AND U16487 ( .A(n15756), .B(n15755), .Z(n15795) );
  XOR U16488 ( .A(n15794), .B(n15795), .Z(n15796) );
  AND U16489 ( .A(x[232]), .B(y[1960]), .Z(n15757) );
  NAND U16490 ( .A(n16225), .B(n15757), .Z(n15761) );
  NAND U16491 ( .A(n15759), .B(n15758), .Z(n15760) );
  AND U16492 ( .A(n15761), .B(n15760), .Z(n15829) );
  AND U16493 ( .A(y[1956]), .B(x[229]), .Z(n15763) );
  NAND U16494 ( .A(y[1954]), .B(x[231]), .Z(n15762) );
  XNOR U16495 ( .A(n15763), .B(n15762), .Z(n15802) );
  AND U16496 ( .A(o[168]), .B(n15764), .Z(n15801) );
  XOR U16497 ( .A(n15802), .B(n15801), .Z(n15827) );
  AND U16498 ( .A(y[1952]), .B(x[233]), .Z(n15766) );
  NAND U16499 ( .A(y[1961]), .B(x[224]), .Z(n15765) );
  XNOR U16500 ( .A(n15766), .B(n15765), .Z(n15809) );
  AND U16501 ( .A(x[232]), .B(y[1953]), .Z(n15818) );
  XOR U16502 ( .A(o[169]), .B(n15818), .Z(n15808) );
  XNOR U16503 ( .A(n15809), .B(n15808), .Z(n15826) );
  XOR U16504 ( .A(n15829), .B(n15828), .Z(n15823) );
  AND U16505 ( .A(y[1955]), .B(x[230]), .Z(n16182) );
  NAND U16506 ( .A(y[1960]), .B(x[225]), .Z(n15767) );
  XNOR U16507 ( .A(n16182), .B(n15767), .Z(n15813) );
  XOR U16508 ( .A(n16230), .B(n15813), .Z(n15833) );
  NAND U16509 ( .A(x[226]), .B(y[1959]), .Z(n16464) );
  AND U16510 ( .A(x[227]), .B(y[1958]), .Z(n16192) );
  XNOR U16511 ( .A(n16464), .B(n16192), .Z(n15832) );
  NAND U16512 ( .A(x[229]), .B(y[1959]), .Z(n16005) );
  AND U16513 ( .A(x[225]), .B(y[1955]), .Z(n15812) );
  NANDN U16514 ( .A(n16005), .B(n15812), .Z(n15771) );
  NAND U16515 ( .A(n15769), .B(n15768), .Z(n15770) );
  NAND U16516 ( .A(n15771), .B(n15770), .Z(n15820) );
  XOR U16517 ( .A(n15821), .B(n15820), .Z(n15822) );
  XNOR U16518 ( .A(n15796), .B(n15797), .Z(n15839) );
  NAND U16519 ( .A(n15773), .B(n15772), .Z(n15777) );
  NAND U16520 ( .A(n15775), .B(n15774), .Z(n15776) );
  NAND U16521 ( .A(n15777), .B(n15776), .Z(n15837) );
  NAND U16522 ( .A(n15779), .B(n15778), .Z(n15783) );
  NAND U16523 ( .A(n15781), .B(n15780), .Z(n15782) );
  NAND U16524 ( .A(n15783), .B(n15782), .Z(n15836) );
  XOR U16525 ( .A(n15837), .B(n15836), .Z(n15838) );
  XOR U16526 ( .A(n15839), .B(n15838), .Z(n15844) );
  NAND U16527 ( .A(n15785), .B(n15784), .Z(n15789) );
  NANDN U16528 ( .A(n15787), .B(n15786), .Z(n15788) );
  NAND U16529 ( .A(n15789), .B(n15788), .Z(n15842) );
  XOR U16530 ( .A(n15842), .B(n15843), .Z(n15793) );
  XNOR U16531 ( .A(n15844), .B(n15793), .Z(N362) );
  NAND U16532 ( .A(n15795), .B(n15794), .Z(n15799) );
  NANDN U16533 ( .A(n15797), .B(n15796), .Z(n15798) );
  AND U16534 ( .A(n15799), .B(n15798), .Z(n15903) );
  AND U16535 ( .A(x[231]), .B(y[1956]), .Z(n15882) );
  NAND U16536 ( .A(n15882), .B(n15800), .Z(n15804) );
  NAND U16537 ( .A(n15802), .B(n15801), .Z(n15803) );
  AND U16538 ( .A(n15804), .B(n15803), .Z(n15895) );
  AND U16539 ( .A(y[1955]), .B(x[231]), .Z(n15806) );
  NAND U16540 ( .A(y[1958]), .B(x[228]), .Z(n15805) );
  XNOR U16541 ( .A(n15806), .B(n15805), .Z(n15866) );
  AND U16542 ( .A(x[230]), .B(y[1956]), .Z(n15865) );
  XNOR U16543 ( .A(n15866), .B(n15865), .Z(n15893) );
  AND U16544 ( .A(x[232]), .B(y[1954]), .Z(n16078) );
  AND U16545 ( .A(x[233]), .B(y[1953]), .Z(n15876) );
  XOR U16546 ( .A(o[170]), .B(n15876), .Z(n15887) );
  XOR U16547 ( .A(n16078), .B(n15887), .Z(n15889) );
  XNOR U16548 ( .A(n15889), .B(n15888), .Z(n15892) );
  XOR U16549 ( .A(n15893), .B(n15892), .Z(n15894) );
  XOR U16550 ( .A(n15895), .B(n15894), .Z(n15855) );
  AND U16551 ( .A(x[233]), .B(y[1961]), .Z(n15807) );
  NAND U16552 ( .A(n15807), .B(n16225), .Z(n15811) );
  NAND U16553 ( .A(n15809), .B(n15808), .Z(n15810) );
  AND U16554 ( .A(n15811), .B(n15810), .Z(n15853) );
  AND U16555 ( .A(x[230]), .B(y[1960]), .Z(n16114) );
  NAND U16556 ( .A(n16114), .B(n15812), .Z(n15815) );
  NAND U16557 ( .A(n16230), .B(n15813), .Z(n15814) );
  NAND U16558 ( .A(n15815), .B(n15814), .Z(n15861) );
  AND U16559 ( .A(y[1952]), .B(x[234]), .Z(n15817) );
  NAND U16560 ( .A(y[1962]), .B(x[224]), .Z(n15816) );
  XNOR U16561 ( .A(n15817), .B(n15816), .Z(n15871) );
  AND U16562 ( .A(o[169]), .B(n15818), .Z(n15870) );
  XOR U16563 ( .A(n15871), .B(n15870), .Z(n15859) );
  AND U16564 ( .A(y[1959]), .B(x[227]), .Z(n16776) );
  NAND U16565 ( .A(y[1961]), .B(x[225]), .Z(n15819) );
  XNOR U16566 ( .A(n16776), .B(n15819), .Z(n15883) );
  AND U16567 ( .A(x[226]), .B(y[1960]), .Z(n15884) );
  XOR U16568 ( .A(n15883), .B(n15884), .Z(n15858) );
  XOR U16569 ( .A(n15859), .B(n15858), .Z(n15860) );
  XOR U16570 ( .A(n15861), .B(n15860), .Z(n15852) );
  NAND U16571 ( .A(n15821), .B(n15820), .Z(n15825) );
  NANDN U16572 ( .A(n15823), .B(n15822), .Z(n15824) );
  NAND U16573 ( .A(n15825), .B(n15824), .Z(n15849) );
  NANDN U16574 ( .A(n15827), .B(n15826), .Z(n15831) );
  NAND U16575 ( .A(n15829), .B(n15828), .Z(n15830) );
  AND U16576 ( .A(n15831), .B(n15830), .Z(n15846) );
  ANDN U16577 ( .B(n16464), .A(n16192), .Z(n15835) );
  NANDN U16578 ( .A(n15833), .B(n15832), .Z(n15834) );
  NANDN U16579 ( .A(n15835), .B(n15834), .Z(n15847) );
  XNOR U16580 ( .A(n15849), .B(n15848), .Z(n15901) );
  XNOR U16581 ( .A(n15903), .B(n15904), .Z(n15900) );
  NAND U16582 ( .A(n15837), .B(n15836), .Z(n15841) );
  NAND U16583 ( .A(n15839), .B(n15838), .Z(n15840) );
  NAND U16584 ( .A(n15841), .B(n15840), .Z(n15899) );
  XOR U16585 ( .A(n15899), .B(n15898), .Z(n15845) );
  XNOR U16586 ( .A(n15900), .B(n15845), .Z(N363) );
  NANDN U16587 ( .A(n15847), .B(n15846), .Z(n15851) );
  NAND U16588 ( .A(n15849), .B(n15848), .Z(n15850) );
  AND U16589 ( .A(n15851), .B(n15850), .Z(n15911) );
  NANDN U16590 ( .A(n15853), .B(n15852), .Z(n15857) );
  NANDN U16591 ( .A(n15855), .B(n15854), .Z(n15856) );
  AND U16592 ( .A(n15857), .B(n15856), .Z(n15909) );
  NAND U16593 ( .A(n15859), .B(n15858), .Z(n15863) );
  NAND U16594 ( .A(n15861), .B(n15860), .Z(n15862) );
  AND U16595 ( .A(n15863), .B(n15862), .Z(n15973) );
  AND U16596 ( .A(x[231]), .B(y[1958]), .Z(n16000) );
  AND U16597 ( .A(x[228]), .B(y[1955]), .Z(n15864) );
  NAND U16598 ( .A(n16000), .B(n15864), .Z(n15868) );
  NAND U16599 ( .A(n15866), .B(n15865), .Z(n15867) );
  AND U16600 ( .A(n15868), .B(n15867), .Z(n15971) );
  AND U16601 ( .A(x[234]), .B(y[1962]), .Z(n15869) );
  NAND U16602 ( .A(n15869), .B(n16225), .Z(n15873) );
  NAND U16603 ( .A(n15871), .B(n15870), .Z(n15872) );
  AND U16604 ( .A(n15873), .B(n15872), .Z(n15967) );
  AND U16605 ( .A(y[1952]), .B(x[235]), .Z(n15875) );
  NAND U16606 ( .A(y[1963]), .B(x[224]), .Z(n15874) );
  XNOR U16607 ( .A(n15875), .B(n15874), .Z(n15942) );
  AND U16608 ( .A(o[170]), .B(n15876), .Z(n15941) );
  XOR U16609 ( .A(n15942), .B(n15941), .Z(n15965) );
  AND U16610 ( .A(y[1957]), .B(x[230]), .Z(n15878) );
  NAND U16611 ( .A(y[1962]), .B(x[225]), .Z(n15877) );
  XNOR U16612 ( .A(n15878), .B(n15877), .Z(n15933) );
  AND U16613 ( .A(x[234]), .B(y[1953]), .Z(n15952) );
  XOR U16614 ( .A(o[171]), .B(n15952), .Z(n15932) );
  XOR U16615 ( .A(n15933), .B(n15932), .Z(n15964) );
  XOR U16616 ( .A(n15965), .B(n15964), .Z(n15966) );
  AND U16617 ( .A(x[227]), .B(y[1960]), .Z(n16906) );
  NAND U16618 ( .A(y[1961]), .B(x[226]), .Z(n15879) );
  XNOR U16619 ( .A(n15880), .B(n15879), .Z(n15928) );
  AND U16620 ( .A(x[228]), .B(y[1959]), .Z(n15927) );
  XNOR U16621 ( .A(n15928), .B(n15927), .Z(n15959) );
  XNOR U16622 ( .A(n16906), .B(n15959), .Z(n15961) );
  NAND U16623 ( .A(y[1954]), .B(x[233]), .Z(n15881) );
  XNOR U16624 ( .A(n15882), .B(n15881), .Z(n15947) );
  AND U16625 ( .A(x[232]), .B(y[1955]), .Z(n15946) );
  XNOR U16626 ( .A(n15947), .B(n15946), .Z(n15960) );
  XNOR U16627 ( .A(n15961), .B(n15960), .Z(n15924) );
  AND U16628 ( .A(x[227]), .B(y[1961]), .Z(n15996) );
  AND U16629 ( .A(x[225]), .B(y[1959]), .Z(n16220) );
  NAND U16630 ( .A(n15996), .B(n16220), .Z(n15886) );
  NAND U16631 ( .A(n15884), .B(n15883), .Z(n15885) );
  NAND U16632 ( .A(n15886), .B(n15885), .Z(n15922) );
  NAND U16633 ( .A(n16078), .B(n15887), .Z(n15891) );
  NAND U16634 ( .A(n15889), .B(n15888), .Z(n15890) );
  NAND U16635 ( .A(n15891), .B(n15890), .Z(n15921) );
  XOR U16636 ( .A(n15922), .B(n15921), .Z(n15923) );
  XNOR U16637 ( .A(n15924), .B(n15923), .Z(n15954) );
  NAND U16638 ( .A(n15893), .B(n15892), .Z(n15897) );
  NAND U16639 ( .A(n15895), .B(n15894), .Z(n15896) );
  NAND U16640 ( .A(n15897), .B(n15896), .Z(n15953) );
  XOR U16641 ( .A(n15954), .B(n15953), .Z(n15956) );
  XNOR U16642 ( .A(n15955), .B(n15956), .Z(n15908) );
  XOR U16643 ( .A(n15911), .B(n15910), .Z(n15917) );
  NANDN U16644 ( .A(n15902), .B(n15901), .Z(n15906) );
  NANDN U16645 ( .A(n15904), .B(n15903), .Z(n15905) );
  AND U16646 ( .A(n15906), .B(n15905), .Z(n15915) );
  IV U16647 ( .A(n15915), .Z(n15914) );
  XOR U16648 ( .A(n15916), .B(n15914), .Z(n15907) );
  XNOR U16649 ( .A(n15917), .B(n15907), .Z(N364) );
  NANDN U16650 ( .A(n15909), .B(n15908), .Z(n15913) );
  NANDN U16651 ( .A(n15911), .B(n15910), .Z(n15912) );
  NAND U16652 ( .A(n15913), .B(n15912), .Z(n16041) );
  IV U16653 ( .A(n16041), .Z(n16040) );
  OR U16654 ( .A(n15916), .B(n15914), .Z(n15920) );
  ANDN U16655 ( .B(n15916), .A(n15915), .Z(n15918) );
  OR U16656 ( .A(n15918), .B(n15917), .Z(n15919) );
  AND U16657 ( .A(n15920), .B(n15919), .Z(n16042) );
  NAND U16658 ( .A(n15922), .B(n15921), .Z(n15926) );
  NAND U16659 ( .A(n15924), .B(n15923), .Z(n15925) );
  AND U16660 ( .A(n15926), .B(n15925), .Z(n16037) );
  AND U16661 ( .A(x[229]), .B(y[1961]), .Z(n16455) );
  NAND U16662 ( .A(n16624), .B(n16455), .Z(n15930) );
  NAND U16663 ( .A(n15928), .B(n15927), .Z(n15929) );
  NAND U16664 ( .A(n15930), .B(n15929), .Z(n15984) );
  AND U16665 ( .A(x[230]), .B(y[1962]), .Z(n16237) );
  NAND U16666 ( .A(n16237), .B(n15931), .Z(n15935) );
  NAND U16667 ( .A(n15933), .B(n15932), .Z(n15934) );
  NAND U16668 ( .A(n15935), .B(n15934), .Z(n15983) );
  XOR U16669 ( .A(n15984), .B(n15983), .Z(n15985) );
  AND U16670 ( .A(x[233]), .B(y[1955]), .Z(n16619) );
  AND U16671 ( .A(y[1954]), .B(x[234]), .Z(n16662) );
  NAND U16672 ( .A(y[1960]), .B(x[228]), .Z(n15936) );
  XNOR U16673 ( .A(n16662), .B(n15936), .Z(n16027) );
  XOR U16674 ( .A(n16619), .B(n16027), .Z(n16006) );
  NAND U16675 ( .A(x[231]), .B(y[1957]), .Z(n16004) );
  XOR U16676 ( .A(n16005), .B(n16004), .Z(n16007) );
  AND U16677 ( .A(y[1952]), .B(x[236]), .Z(n15938) );
  NAND U16678 ( .A(y[1964]), .B(x[224]), .Z(n15937) );
  XNOR U16679 ( .A(n15938), .B(n15937), .Z(n16021) );
  AND U16680 ( .A(x[235]), .B(y[1953]), .Z(n16001) );
  XOR U16681 ( .A(o[172]), .B(n16001), .Z(n16020) );
  XOR U16682 ( .A(n16021), .B(n16020), .Z(n15990) );
  AND U16683 ( .A(y[1962]), .B(x[226]), .Z(n15940) );
  NAND U16684 ( .A(y[1956]), .B(x[232]), .Z(n15939) );
  XNOR U16685 ( .A(n15940), .B(n15939), .Z(n15995) );
  XOR U16686 ( .A(n15995), .B(n15996), .Z(n15989) );
  XOR U16687 ( .A(n15990), .B(n15989), .Z(n15991) );
  XNOR U16688 ( .A(n15985), .B(n15986), .Z(n16035) );
  AND U16689 ( .A(x[235]), .B(y[1963]), .Z(n17034) );
  NAND U16690 ( .A(n17034), .B(n16225), .Z(n15944) );
  NAND U16691 ( .A(n15942), .B(n15941), .Z(n15943) );
  NAND U16692 ( .A(n15944), .B(n15943), .Z(n16013) );
  AND U16693 ( .A(x[231]), .B(y[1954]), .Z(n16168) );
  AND U16694 ( .A(x[233]), .B(y[1956]), .Z(n15945) );
  NAND U16695 ( .A(n16168), .B(n15945), .Z(n15949) );
  NAND U16696 ( .A(n15947), .B(n15946), .Z(n15948) );
  NAND U16697 ( .A(n15949), .B(n15948), .Z(n16011) );
  NAND U16698 ( .A(y[1963]), .B(x[225]), .Z(n15950) );
  XNOR U16699 ( .A(n15951), .B(n15950), .Z(n16017) );
  AND U16700 ( .A(o[171]), .B(n15952), .Z(n16016) );
  XOR U16701 ( .A(n16017), .B(n16016), .Z(n16010) );
  XOR U16702 ( .A(n16011), .B(n16010), .Z(n16012) );
  XOR U16703 ( .A(n16013), .B(n16012), .Z(n16034) );
  XOR U16704 ( .A(n16035), .B(n16034), .Z(n16036) );
  NAND U16705 ( .A(n15954), .B(n15953), .Z(n15958) );
  NAND U16706 ( .A(n15956), .B(n15955), .Z(n15957) );
  NAND U16707 ( .A(n15958), .B(n15957), .Z(n16047) );
  XOR U16708 ( .A(n16048), .B(n16047), .Z(n16050) );
  NANDN U16709 ( .A(n16906), .B(n15959), .Z(n15963) );
  NAND U16710 ( .A(n15961), .B(n15960), .Z(n15962) );
  AND U16711 ( .A(n15963), .B(n15962), .Z(n15978) );
  NAND U16712 ( .A(n15965), .B(n15964), .Z(n15969) );
  NANDN U16713 ( .A(n15967), .B(n15966), .Z(n15968) );
  AND U16714 ( .A(n15969), .B(n15968), .Z(n15977) );
  NANDN U16715 ( .A(n15971), .B(n15970), .Z(n15975) );
  NANDN U16716 ( .A(n15973), .B(n15972), .Z(n15974) );
  NAND U16717 ( .A(n15975), .B(n15974), .Z(n15980) );
  XOR U16718 ( .A(n16050), .B(n16049), .Z(n16043) );
  XNOR U16719 ( .A(n16042), .B(n16043), .Z(n15976) );
  XOR U16720 ( .A(n16040), .B(n15976), .Z(N365) );
  NANDN U16721 ( .A(n15978), .B(n15977), .Z(n15982) );
  NANDN U16722 ( .A(n15980), .B(n15979), .Z(n15981) );
  AND U16723 ( .A(n15982), .B(n15981), .Z(n16124) );
  NAND U16724 ( .A(n15984), .B(n15983), .Z(n15988) );
  NANDN U16725 ( .A(n15986), .B(n15985), .Z(n15987) );
  NAND U16726 ( .A(n15988), .B(n15987), .Z(n16054) );
  NAND U16727 ( .A(n15990), .B(n15989), .Z(n15994) );
  NANDN U16728 ( .A(n15992), .B(n15991), .Z(n15993) );
  NAND U16729 ( .A(n15994), .B(n15993), .Z(n16062) );
  AND U16730 ( .A(y[1962]), .B(x[232]), .Z(n17272) );
  AND U16731 ( .A(x[226]), .B(y[1956]), .Z(n16178) );
  NAND U16732 ( .A(n17272), .B(n16178), .Z(n15998) );
  NAND U16733 ( .A(n15996), .B(n15995), .Z(n15997) );
  NAND U16734 ( .A(n15998), .B(n15997), .Z(n16093) );
  NAND U16735 ( .A(y[1964]), .B(x[225]), .Z(n15999) );
  XNOR U16736 ( .A(n16000), .B(n15999), .Z(n16084) );
  AND U16737 ( .A(o[172]), .B(n16001), .Z(n16083) );
  XOR U16738 ( .A(n16084), .B(n16083), .Z(n16091) );
  AND U16739 ( .A(x[230]), .B(y[1959]), .Z(n17074) );
  AND U16740 ( .A(y[1963]), .B(x[226]), .Z(n16003) );
  NAND U16741 ( .A(y[1956]), .B(x[233]), .Z(n16002) );
  XNOR U16742 ( .A(n16003), .B(n16002), .Z(n16097) );
  XOR U16743 ( .A(n17074), .B(n16097), .Z(n16090) );
  XOR U16744 ( .A(n16091), .B(n16090), .Z(n16092) );
  XOR U16745 ( .A(n16093), .B(n16092), .Z(n16061) );
  NAND U16746 ( .A(n16005), .B(n16004), .Z(n16009) );
  ANDN U16747 ( .B(n16007), .A(n16006), .Z(n16008) );
  ANDN U16748 ( .B(n16009), .A(n16008), .Z(n16060) );
  XOR U16749 ( .A(n16061), .B(n16060), .Z(n16063) );
  XOR U16750 ( .A(n16062), .B(n16063), .Z(n16055) );
  XOR U16751 ( .A(n16054), .B(n16055), .Z(n16057) );
  NAND U16752 ( .A(n16011), .B(n16010), .Z(n16015) );
  NAND U16753 ( .A(n16013), .B(n16012), .Z(n16014) );
  NAND U16754 ( .A(n16015), .B(n16014), .Z(n16069) );
  AND U16755 ( .A(x[230]), .B(y[1963]), .Z(n16456) );
  AND U16756 ( .A(x[225]), .B(y[1958]), .Z(n16082) );
  NAND U16757 ( .A(n16456), .B(n16082), .Z(n16019) );
  NAND U16758 ( .A(n16017), .B(n16016), .Z(n16018) );
  NAND U16759 ( .A(n16019), .B(n16018), .Z(n16075) );
  AND U16760 ( .A(x[236]), .B(y[1964]), .Z(n17278) );
  NAND U16761 ( .A(n17278), .B(n16225), .Z(n16023) );
  NAND U16762 ( .A(n16021), .B(n16020), .Z(n16022) );
  NAND U16763 ( .A(n16023), .B(n16022), .Z(n16073) );
  AND U16764 ( .A(x[234]), .B(y[1955]), .Z(n16918) );
  AND U16765 ( .A(y[1954]), .B(x[235]), .Z(n16879) );
  NAND U16766 ( .A(y[1957]), .B(x[232]), .Z(n16024) );
  XNOR U16767 ( .A(n16879), .B(n16024), .Z(n16079) );
  XOR U16768 ( .A(n16918), .B(n16079), .Z(n16072) );
  XOR U16769 ( .A(n16073), .B(n16072), .Z(n16074) );
  XOR U16770 ( .A(n16075), .B(n16074), .Z(n16067) );
  AND U16771 ( .A(x[234]), .B(y[1960]), .Z(n16026) );
  AND U16772 ( .A(x[228]), .B(y[1954]), .Z(n16025) );
  NAND U16773 ( .A(n16026), .B(n16025), .Z(n16029) );
  NAND U16774 ( .A(n16027), .B(n16619), .Z(n16028) );
  NAND U16775 ( .A(n16029), .B(n16028), .Z(n16118) );
  AND U16776 ( .A(y[1952]), .B(x[237]), .Z(n16031) );
  NAND U16777 ( .A(y[1965]), .B(x[224]), .Z(n16030) );
  XNOR U16778 ( .A(n16031), .B(n16030), .Z(n16110) );
  AND U16779 ( .A(x[236]), .B(y[1953]), .Z(n16102) );
  XOR U16780 ( .A(o[173]), .B(n16102), .Z(n16109) );
  XOR U16781 ( .A(n16110), .B(n16109), .Z(n16116) );
  AND U16782 ( .A(y[1960]), .B(x[229]), .Z(n16033) );
  NAND U16783 ( .A(y[1962]), .B(x[227]), .Z(n16032) );
  XNOR U16784 ( .A(n16033), .B(n16032), .Z(n16105) );
  AND U16785 ( .A(x[228]), .B(y[1961]), .Z(n16106) );
  XOR U16786 ( .A(n16105), .B(n16106), .Z(n16115) );
  XOR U16787 ( .A(n16116), .B(n16115), .Z(n16117) );
  XOR U16788 ( .A(n16118), .B(n16117), .Z(n16066) );
  XOR U16789 ( .A(n16067), .B(n16066), .Z(n16068) );
  XOR U16790 ( .A(n16069), .B(n16068), .Z(n16056) );
  XOR U16791 ( .A(n16057), .B(n16056), .Z(n16122) );
  NAND U16792 ( .A(n16035), .B(n16034), .Z(n16039) );
  NANDN U16793 ( .A(n16037), .B(n16036), .Z(n16038) );
  AND U16794 ( .A(n16039), .B(n16038), .Z(n16121) );
  XOR U16795 ( .A(n16124), .B(n16123), .Z(n16130) );
  OR U16796 ( .A(n16042), .B(n16040), .Z(n16046) );
  ANDN U16797 ( .B(n16042), .A(n16041), .Z(n16044) );
  OR U16798 ( .A(n16044), .B(n16043), .Z(n16045) );
  AND U16799 ( .A(n16046), .B(n16045), .Z(n16128) );
  NAND U16800 ( .A(n16048), .B(n16047), .Z(n16052) );
  NAND U16801 ( .A(n16050), .B(n16049), .Z(n16051) );
  NAND U16802 ( .A(n16052), .B(n16051), .Z(n16129) );
  IV U16803 ( .A(n16129), .Z(n16127) );
  XOR U16804 ( .A(n16128), .B(n16127), .Z(n16053) );
  XNOR U16805 ( .A(n16130), .B(n16053), .Z(N366) );
  NAND U16806 ( .A(n16055), .B(n16054), .Z(n16059) );
  NAND U16807 ( .A(n16057), .B(n16056), .Z(n16058) );
  NAND U16808 ( .A(n16059), .B(n16058), .Z(n16136) );
  NAND U16809 ( .A(n16061), .B(n16060), .Z(n16065) );
  NAND U16810 ( .A(n16063), .B(n16062), .Z(n16064) );
  NAND U16811 ( .A(n16065), .B(n16064), .Z(n16135) );
  XOR U16812 ( .A(n16136), .B(n16135), .Z(n16137) );
  NAND U16813 ( .A(n16067), .B(n16066), .Z(n16071) );
  NAND U16814 ( .A(n16069), .B(n16068), .Z(n16070) );
  NAND U16815 ( .A(n16071), .B(n16070), .Z(n16147) );
  NAND U16816 ( .A(n16073), .B(n16072), .Z(n16077) );
  NAND U16817 ( .A(n16075), .B(n16074), .Z(n16076) );
  AND U16818 ( .A(n16077), .B(n16076), .Z(n16153) );
  AND U16819 ( .A(x[235]), .B(y[1957]), .Z(n16251) );
  NAND U16820 ( .A(n16251), .B(n16078), .Z(n16081) );
  NAND U16821 ( .A(n16079), .B(n16918), .Z(n16080) );
  NAND U16822 ( .A(n16081), .B(n16080), .Z(n16208) );
  NAND U16823 ( .A(x[231]), .B(y[1964]), .Z(n16634) );
  NANDN U16824 ( .A(n16634), .B(n16082), .Z(n16086) );
  NAND U16825 ( .A(n16084), .B(n16083), .Z(n16085) );
  NAND U16826 ( .A(n16086), .B(n16085), .Z(n16207) );
  XOR U16827 ( .A(n16208), .B(n16207), .Z(n16210) );
  AND U16828 ( .A(x[228]), .B(y[1962]), .Z(n16553) );
  AND U16829 ( .A(y[1963]), .B(x[227]), .Z(n16088) );
  NAND U16830 ( .A(y[1958]), .B(x[232]), .Z(n16087) );
  XNOR U16831 ( .A(n16088), .B(n16087), .Z(n16193) );
  XOR U16832 ( .A(n16455), .B(n16193), .Z(n16202) );
  XOR U16833 ( .A(n16553), .B(n16202), .Z(n16204) );
  AND U16834 ( .A(x[233]), .B(y[1957]), .Z(n16741) );
  AND U16835 ( .A(y[1964]), .B(x[226]), .Z(n16089) );
  AND U16836 ( .A(y[1956]), .B(x[234]), .Z(n16771) );
  XOR U16837 ( .A(n16089), .B(n16771), .Z(n16179) );
  XOR U16838 ( .A(n16741), .B(n16179), .Z(n16203) );
  XOR U16839 ( .A(n16204), .B(n16203), .Z(n16209) );
  XNOR U16840 ( .A(n16210), .B(n16209), .Z(n16151) );
  NAND U16841 ( .A(n16091), .B(n16090), .Z(n16095) );
  NAND U16842 ( .A(n16093), .B(n16092), .Z(n16094) );
  AND U16843 ( .A(n16095), .B(n16094), .Z(n16150) );
  XOR U16844 ( .A(n16151), .B(n16150), .Z(n16152) );
  XNOR U16845 ( .A(n16153), .B(n16152), .Z(n16145) );
  AND U16846 ( .A(x[233]), .B(y[1963]), .Z(n16096) );
  NAND U16847 ( .A(n16096), .B(n16178), .Z(n16099) );
  NAND U16848 ( .A(n16097), .B(n17074), .Z(n16098) );
  NAND U16849 ( .A(n16099), .B(n16098), .Z(n16165) );
  AND U16850 ( .A(y[1952]), .B(x[238]), .Z(n16101) );
  NAND U16851 ( .A(y[1966]), .B(x[224]), .Z(n16100) );
  XNOR U16852 ( .A(n16101), .B(n16100), .Z(n16188) );
  AND U16853 ( .A(o[173]), .B(n16102), .Z(n16187) );
  XOR U16854 ( .A(n16188), .B(n16187), .Z(n16163) );
  NAND U16855 ( .A(y[1954]), .B(x[236]), .Z(n16103) );
  XNOR U16856 ( .A(n16104), .B(n16103), .Z(n16169) );
  NAND U16857 ( .A(x[237]), .B(y[1953]), .Z(n16177) );
  XNOR U16858 ( .A(o[174]), .B(n16177), .Z(n16170) );
  XOR U16859 ( .A(n16169), .B(n16170), .Z(n16162) );
  XOR U16860 ( .A(n16163), .B(n16162), .Z(n16164) );
  XNOR U16861 ( .A(n16165), .B(n16164), .Z(n16214) );
  NAND U16862 ( .A(x[229]), .B(y[1962]), .Z(n16238) );
  NANDN U16863 ( .A(n16238), .B(n16906), .Z(n16108) );
  NAND U16864 ( .A(n16106), .B(n16105), .Z(n16107) );
  AND U16865 ( .A(n16108), .B(n16107), .Z(n16159) );
  AND U16866 ( .A(x[237]), .B(y[1965]), .Z(n17605) );
  NAND U16867 ( .A(n17605), .B(n16225), .Z(n16112) );
  NAND U16868 ( .A(n16110), .B(n16109), .Z(n16111) );
  NAND U16869 ( .A(n16112), .B(n16111), .Z(n16157) );
  NAND U16870 ( .A(y[1955]), .B(x[235]), .Z(n16113) );
  XNOR U16871 ( .A(n16114), .B(n16113), .Z(n16183) );
  NAND U16872 ( .A(x[225]), .B(y[1965]), .Z(n16184) );
  XOR U16873 ( .A(n16157), .B(n16156), .Z(n16158) );
  XOR U16874 ( .A(n16159), .B(n16158), .Z(n16213) );
  XOR U16875 ( .A(n16214), .B(n16213), .Z(n16216) );
  NAND U16876 ( .A(n16116), .B(n16115), .Z(n16120) );
  NAND U16877 ( .A(n16118), .B(n16117), .Z(n16119) );
  AND U16878 ( .A(n16120), .B(n16119), .Z(n16215) );
  XNOR U16879 ( .A(n16216), .B(n16215), .Z(n16144) );
  XOR U16880 ( .A(n16145), .B(n16144), .Z(n16146) );
  XNOR U16881 ( .A(n16147), .B(n16146), .Z(n16138) );
  XNOR U16882 ( .A(n16137), .B(n16138), .Z(n16143) );
  NANDN U16883 ( .A(n16122), .B(n16121), .Z(n16126) );
  NANDN U16884 ( .A(n16124), .B(n16123), .Z(n16125) );
  NAND U16885 ( .A(n16126), .B(n16125), .Z(n16141) );
  NANDN U16886 ( .A(n16127), .B(n16128), .Z(n16133) );
  NOR U16887 ( .A(n16129), .B(n16128), .Z(n16131) );
  OR U16888 ( .A(n16131), .B(n16130), .Z(n16132) );
  AND U16889 ( .A(n16133), .B(n16132), .Z(n16142) );
  XOR U16890 ( .A(n16141), .B(n16142), .Z(n16134) );
  XNOR U16891 ( .A(n16143), .B(n16134), .Z(N367) );
  NAND U16892 ( .A(n16136), .B(n16135), .Z(n16140) );
  NANDN U16893 ( .A(n16138), .B(n16137), .Z(n16139) );
  AND U16894 ( .A(n16140), .B(n16139), .Z(n16308) );
  NAND U16895 ( .A(n16145), .B(n16144), .Z(n16149) );
  NAND U16896 ( .A(n16147), .B(n16146), .Z(n16148) );
  NAND U16897 ( .A(n16149), .B(n16148), .Z(n16305) );
  NAND U16898 ( .A(n16151), .B(n16150), .Z(n16155) );
  NAND U16899 ( .A(n16153), .B(n16152), .Z(n16154) );
  NAND U16900 ( .A(n16155), .B(n16154), .Z(n16280) );
  NAND U16901 ( .A(n16157), .B(n16156), .Z(n16161) );
  NANDN U16902 ( .A(n16159), .B(n16158), .Z(n16160) );
  AND U16903 ( .A(n16161), .B(n16160), .Z(n16287) );
  NAND U16904 ( .A(n16163), .B(n16162), .Z(n16167) );
  NAND U16905 ( .A(n16165), .B(n16164), .Z(n16166) );
  AND U16906 ( .A(n16167), .B(n16166), .Z(n16285) );
  NAND U16907 ( .A(x[236]), .B(y[1959]), .Z(n16626) );
  NANDN U16908 ( .A(n16626), .B(n16168), .Z(n16172) );
  NAND U16909 ( .A(n16170), .B(n16169), .Z(n16171) );
  AND U16910 ( .A(n16172), .B(n16171), .Z(n16261) );
  AND U16911 ( .A(y[1956]), .B(x[235]), .Z(n16174) );
  NAND U16912 ( .A(y[1954]), .B(x[237]), .Z(n16173) );
  XNOR U16913 ( .A(n16174), .B(n16173), .Z(n16265) );
  AND U16914 ( .A(x[236]), .B(y[1955]), .Z(n16264) );
  XNOR U16915 ( .A(n16265), .B(n16264), .Z(n16259) );
  AND U16916 ( .A(y[1952]), .B(x[239]), .Z(n16176) );
  NAND U16917 ( .A(y[1967]), .B(x[224]), .Z(n16175) );
  XNOR U16918 ( .A(n16176), .B(n16175), .Z(n16227) );
  ANDN U16919 ( .B(o[174]), .A(n16177), .Z(n16226) );
  XNOR U16920 ( .A(n16227), .B(n16226), .Z(n16258) );
  XOR U16921 ( .A(n16259), .B(n16258), .Z(n16260) );
  XOR U16922 ( .A(n16261), .B(n16260), .Z(n16293) );
  NAND U16923 ( .A(x[234]), .B(y[1964]), .Z(n17076) );
  NANDN U16924 ( .A(n17076), .B(n16178), .Z(n16181) );
  NAND U16925 ( .A(n16741), .B(n16179), .Z(n16180) );
  AND U16926 ( .A(n16181), .B(n16180), .Z(n16291) );
  AND U16927 ( .A(x[235]), .B(y[1960]), .Z(n16551) );
  NAND U16928 ( .A(n16551), .B(n16182), .Z(n16186) );
  NANDN U16929 ( .A(n16184), .B(n16183), .Z(n16185) );
  NAND U16930 ( .A(n16186), .B(n16185), .Z(n16290) );
  AND U16931 ( .A(x[238]), .B(y[1966]), .Z(n17858) );
  NAND U16932 ( .A(n17858), .B(n16225), .Z(n16190) );
  NAND U16933 ( .A(n16188), .B(n16187), .Z(n16189) );
  NAND U16934 ( .A(n16190), .B(n16189), .Z(n16253) );
  AND U16935 ( .A(x[232]), .B(y[1963]), .Z(n16191) );
  NAND U16936 ( .A(n16192), .B(n16191), .Z(n16195) );
  NAND U16937 ( .A(n16193), .B(n16455), .Z(n16194) );
  NAND U16938 ( .A(n16195), .B(n16194), .Z(n16252) );
  XOR U16939 ( .A(n16253), .B(n16252), .Z(n16255) );
  AND U16940 ( .A(y[1957]), .B(x[234]), .Z(n16197) );
  NAND U16941 ( .A(y[1963]), .B(x[228]), .Z(n16196) );
  XNOR U16942 ( .A(n16197), .B(n16196), .Z(n16233) );
  AND U16943 ( .A(x[231]), .B(y[1960]), .Z(n16232) );
  XNOR U16944 ( .A(n16233), .B(n16232), .Z(n16240) );
  AND U16945 ( .A(x[230]), .B(y[1961]), .Z(n16370) );
  XNOR U16946 ( .A(n16370), .B(n16238), .Z(n16239) );
  XNOR U16947 ( .A(n16240), .B(n16239), .Z(n16275) );
  AND U16948 ( .A(y[1965]), .B(x[226]), .Z(n16199) );
  NAND U16949 ( .A(y[1958]), .B(x[233]), .Z(n16198) );
  XNOR U16950 ( .A(n16199), .B(n16198), .Z(n16243) );
  AND U16951 ( .A(x[227]), .B(y[1964]), .Z(n16244) );
  XOR U16952 ( .A(n16243), .B(n16244), .Z(n16273) );
  AND U16953 ( .A(y[1966]), .B(x[225]), .Z(n16201) );
  NAND U16954 ( .A(y[1959]), .B(x[232]), .Z(n16200) );
  XNOR U16955 ( .A(n16201), .B(n16200), .Z(n16222) );
  NAND U16956 ( .A(x[238]), .B(y[1953]), .Z(n16247) );
  XNOR U16957 ( .A(o[175]), .B(n16247), .Z(n16221) );
  XOR U16958 ( .A(n16222), .B(n16221), .Z(n16272) );
  XOR U16959 ( .A(n16273), .B(n16272), .Z(n16274) );
  XOR U16960 ( .A(n16275), .B(n16274), .Z(n16254) );
  XOR U16961 ( .A(n16255), .B(n16254), .Z(n16297) );
  NAND U16962 ( .A(n16553), .B(n16202), .Z(n16206) );
  NAND U16963 ( .A(n16204), .B(n16203), .Z(n16205) );
  AND U16964 ( .A(n16206), .B(n16205), .Z(n16296) );
  NAND U16965 ( .A(n16208), .B(n16207), .Z(n16212) );
  NAND U16966 ( .A(n16210), .B(n16209), .Z(n16211) );
  AND U16967 ( .A(n16212), .B(n16211), .Z(n16298) );
  XOR U16968 ( .A(n16299), .B(n16298), .Z(n16278) );
  XNOR U16969 ( .A(n16279), .B(n16278), .Z(n16281) );
  XOR U16970 ( .A(n16280), .B(n16281), .Z(n16302) );
  NAND U16971 ( .A(n16214), .B(n16213), .Z(n16218) );
  NAND U16972 ( .A(n16216), .B(n16215), .Z(n16217) );
  AND U16973 ( .A(n16218), .B(n16217), .Z(n16303) );
  XOR U16974 ( .A(n16302), .B(n16303), .Z(n16304) );
  XOR U16975 ( .A(n16305), .B(n16304), .Z(n16310) );
  XNOR U16976 ( .A(n16309), .B(n16310), .Z(n16219) );
  XOR U16977 ( .A(n16308), .B(n16219), .Z(N368) );
  AND U16978 ( .A(x[232]), .B(y[1966]), .Z(n16552) );
  NAND U16979 ( .A(n16552), .B(n16220), .Z(n16224) );
  NAND U16980 ( .A(n16222), .B(n16221), .Z(n16223) );
  NAND U16981 ( .A(n16224), .B(n16223), .Z(n16324) );
  AND U16982 ( .A(x[239]), .B(y[1967]), .Z(n18118) );
  NAND U16983 ( .A(n18118), .B(n16225), .Z(n16229) );
  NAND U16984 ( .A(n16227), .B(n16226), .Z(n16228) );
  NAND U16985 ( .A(n16229), .B(n16228), .Z(n16325) );
  XOR U16986 ( .A(n16324), .B(n16325), .Z(n16326) );
  AND U16987 ( .A(x[234]), .B(y[1963]), .Z(n16231) );
  NAND U16988 ( .A(n16231), .B(n16230), .Z(n16235) );
  NAND U16989 ( .A(n16233), .B(n16232), .Z(n16234) );
  NAND U16990 ( .A(n16235), .B(n16234), .Z(n16357) );
  AND U16991 ( .A(x[224]), .B(y[1968]), .Z(n16379) );
  NAND U16992 ( .A(x[240]), .B(y[1952]), .Z(n16380) );
  XNOR U16993 ( .A(n16379), .B(n16380), .Z(n16381) );
  NAND U16994 ( .A(x[239]), .B(y[1953]), .Z(n16367) );
  XOR U16995 ( .A(o[176]), .B(n16367), .Z(n16382) );
  XNOR U16996 ( .A(n16381), .B(n16382), .Z(n16356) );
  NAND U16997 ( .A(y[1961]), .B(x[231]), .Z(n16236) );
  XNOR U16998 ( .A(n16237), .B(n16236), .Z(n16371) );
  NAND U16999 ( .A(x[234]), .B(y[1958]), .Z(n16372) );
  XNOR U17000 ( .A(n16371), .B(n16372), .Z(n16355) );
  XOR U17001 ( .A(n16356), .B(n16355), .Z(n16358) );
  XNOR U17002 ( .A(n16357), .B(n16358), .Z(n16327) );
  XOR U17003 ( .A(n16326), .B(n16327), .Z(n16351) );
  NANDN U17004 ( .A(n16370), .B(n16238), .Z(n16242) );
  NAND U17005 ( .A(n16240), .B(n16239), .Z(n16241) );
  NAND U17006 ( .A(n16242), .B(n16241), .Z(n16350) );
  NAND U17007 ( .A(x[233]), .B(y[1965]), .Z(n17057) );
  NANDN U17008 ( .A(n17057), .B(n16624), .Z(n16246) );
  NAND U17009 ( .A(n16244), .B(n16243), .Z(n16245) );
  NAND U17010 ( .A(n16246), .B(n16245), .Z(n16389) );
  ANDN U17011 ( .B(o[175]), .A(n16247), .Z(n16375) );
  AND U17012 ( .A(y[1967]), .B(x[225]), .Z(n16249) );
  NAND U17013 ( .A(y[1960]), .B(x[232]), .Z(n16248) );
  XOR U17014 ( .A(n16249), .B(n16248), .Z(n16376) );
  XNOR U17015 ( .A(n16375), .B(n16376), .Z(n16388) );
  NAND U17016 ( .A(y[1954]), .B(x[238]), .Z(n16250) );
  XNOR U17017 ( .A(n16251), .B(n16250), .Z(n16332) );
  NAND U17018 ( .A(x[228]), .B(y[1964]), .Z(n16333) );
  XNOR U17019 ( .A(n16332), .B(n16333), .Z(n16387) );
  XOR U17020 ( .A(n16388), .B(n16387), .Z(n16390) );
  XNOR U17021 ( .A(n16389), .B(n16390), .Z(n16349) );
  XOR U17022 ( .A(n16350), .B(n16349), .Z(n16352) );
  XOR U17023 ( .A(n16351), .B(n16352), .Z(n16318) );
  NAND U17024 ( .A(n16253), .B(n16252), .Z(n16257) );
  NAND U17025 ( .A(n16255), .B(n16254), .Z(n16256) );
  AND U17026 ( .A(n16257), .B(n16256), .Z(n16319) );
  XOR U17027 ( .A(n16318), .B(n16319), .Z(n16321) );
  NAND U17028 ( .A(n16259), .B(n16258), .Z(n16263) );
  NAND U17029 ( .A(n16261), .B(n16260), .Z(n16262) );
  NAND U17030 ( .A(n16263), .B(n16262), .Z(n16345) );
  AND U17031 ( .A(x[237]), .B(y[1956]), .Z(n16342) );
  NAND U17032 ( .A(n16879), .B(n16342), .Z(n16267) );
  NAND U17033 ( .A(n16265), .B(n16264), .Z(n16266) );
  NAND U17034 ( .A(n16267), .B(n16266), .Z(n16330) );
  AND U17035 ( .A(y[1966]), .B(x[226]), .Z(n16269) );
  NAND U17036 ( .A(y[1959]), .B(x[233]), .Z(n16268) );
  XNOR U17037 ( .A(n16269), .B(n16268), .Z(n16336) );
  NAND U17038 ( .A(x[227]), .B(y[1965]), .Z(n16337) );
  XNOR U17039 ( .A(n16336), .B(n16337), .Z(n16329) );
  AND U17040 ( .A(x[236]), .B(y[1956]), .Z(n17045) );
  AND U17041 ( .A(y[1963]), .B(x[229]), .Z(n16271) );
  NAND U17042 ( .A(y[1955]), .B(x[237]), .Z(n16270) );
  XNOR U17043 ( .A(n16271), .B(n16270), .Z(n16362) );
  XOR U17044 ( .A(n17045), .B(n16362), .Z(n16328) );
  XOR U17045 ( .A(n16329), .B(n16328), .Z(n16331) );
  XNOR U17046 ( .A(n16330), .B(n16331), .Z(n16344) );
  NAND U17047 ( .A(n16273), .B(n16272), .Z(n16277) );
  NAND U17048 ( .A(n16275), .B(n16274), .Z(n16276) );
  AND U17049 ( .A(n16277), .B(n16276), .Z(n16343) );
  XOR U17050 ( .A(n16344), .B(n16343), .Z(n16346) );
  XOR U17051 ( .A(n16345), .B(n16346), .Z(n16320) );
  XNOR U17052 ( .A(n16321), .B(n16320), .Z(n16397) );
  NAND U17053 ( .A(n16279), .B(n16278), .Z(n16283) );
  NANDN U17054 ( .A(n16281), .B(n16280), .Z(n16282) );
  AND U17055 ( .A(n16283), .B(n16282), .Z(n16396) );
  XOR U17056 ( .A(n16397), .B(n16396), .Z(n16399) );
  NANDN U17057 ( .A(n16285), .B(n16284), .Z(n16289) );
  NANDN U17058 ( .A(n16287), .B(n16286), .Z(n16288) );
  AND U17059 ( .A(n16289), .B(n16288), .Z(n16315) );
  NANDN U17060 ( .A(n16291), .B(n16290), .Z(n16295) );
  NANDN U17061 ( .A(n16293), .B(n16292), .Z(n16294) );
  AND U17062 ( .A(n16295), .B(n16294), .Z(n16313) );
  NANDN U17063 ( .A(n16297), .B(n16296), .Z(n16301) );
  NAND U17064 ( .A(n16299), .B(n16298), .Z(n16300) );
  AND U17065 ( .A(n16301), .B(n16300), .Z(n16312) );
  XNOR U17066 ( .A(n16399), .B(n16398), .Z(n16395) );
  NAND U17067 ( .A(n16303), .B(n16302), .Z(n16307) );
  NAND U17068 ( .A(n16305), .B(n16304), .Z(n16306) );
  NAND U17069 ( .A(n16307), .B(n16306), .Z(n16394) );
  XOR U17070 ( .A(n16394), .B(n16393), .Z(n16311) );
  XNOR U17071 ( .A(n16395), .B(n16311), .Z(N369) );
  NANDN U17072 ( .A(n16313), .B(n16312), .Z(n16317) );
  NANDN U17073 ( .A(n16315), .B(n16314), .Z(n16316) );
  AND U17074 ( .A(n16317), .B(n16316), .Z(n16492) );
  NAND U17075 ( .A(n16319), .B(n16318), .Z(n16323) );
  NAND U17076 ( .A(n16321), .B(n16320), .Z(n16322) );
  NAND U17077 ( .A(n16323), .B(n16322), .Z(n16405) );
  NAND U17078 ( .A(x[238]), .B(y[1957]), .Z(n16659) );
  NANDN U17079 ( .A(n16659), .B(n16879), .Z(n16335) );
  NANDN U17080 ( .A(n16333), .B(n16332), .Z(n16334) );
  AND U17081 ( .A(n16335), .B(n16334), .Z(n16476) );
  AND U17082 ( .A(x[233]), .B(y[1966]), .Z(n17269) );
  NANDN U17083 ( .A(n16464), .B(n17269), .Z(n16339) );
  NANDN U17084 ( .A(n16337), .B(n16336), .Z(n16338) );
  NAND U17085 ( .A(n16339), .B(n16338), .Z(n16475) );
  XNOR U17086 ( .A(n16476), .B(n16475), .Z(n16477) );
  AND U17087 ( .A(x[229]), .B(y[1964]), .Z(n16513) );
  NAND U17088 ( .A(y[1961]), .B(x[232]), .Z(n16340) );
  XNOR U17089 ( .A(n16513), .B(n16340), .Z(n16457) );
  XOR U17090 ( .A(n16457), .B(n16456), .Z(n16469) );
  AND U17091 ( .A(x[231]), .B(y[1962]), .Z(n16470) );
  XOR U17092 ( .A(n16469), .B(n16470), .Z(n16471) );
  NAND U17093 ( .A(y[1965]), .B(x[228]), .Z(n16341) );
  XNOR U17094 ( .A(n16342), .B(n16341), .Z(n16420) );
  NAND U17095 ( .A(x[235]), .B(y[1958]), .Z(n16421) );
  XOR U17096 ( .A(n16420), .B(n16421), .Z(n16472) );
  XOR U17097 ( .A(n16471), .B(n16472), .Z(n16478) );
  XNOR U17098 ( .A(n16477), .B(n16478), .Z(n16482) );
  XOR U17099 ( .A(n16481), .B(n16482), .Z(n16484) );
  XNOR U17100 ( .A(n16483), .B(n16484), .Z(n16404) );
  NAND U17101 ( .A(n16344), .B(n16343), .Z(n16348) );
  NAND U17102 ( .A(n16346), .B(n16345), .Z(n16347) );
  NAND U17103 ( .A(n16348), .B(n16347), .Z(n16403) );
  XNOR U17104 ( .A(n16404), .B(n16403), .Z(n16406) );
  XOR U17105 ( .A(n16405), .B(n16406), .Z(n16490) );
  NAND U17106 ( .A(n16350), .B(n16349), .Z(n16354) );
  NAND U17107 ( .A(n16352), .B(n16351), .Z(n16353) );
  NAND U17108 ( .A(n16354), .B(n16353), .Z(n16411) );
  NAND U17109 ( .A(n16356), .B(n16355), .Z(n16360) );
  NAND U17110 ( .A(n16358), .B(n16357), .Z(n16359) );
  NAND U17111 ( .A(n16360), .B(n16359), .Z(n16487) );
  AND U17112 ( .A(x[237]), .B(y[1963]), .Z(n17286) );
  NAND U17113 ( .A(n17286), .B(n16361), .Z(n16364) );
  NAND U17114 ( .A(n17045), .B(n16362), .Z(n16363) );
  AND U17115 ( .A(n16364), .B(n16363), .Z(n16442) );
  AND U17116 ( .A(y[1968]), .B(x[225]), .Z(n16366) );
  NAND U17117 ( .A(y[1960]), .B(x[233]), .Z(n16365) );
  XNOR U17118 ( .A(n16366), .B(n16365), .Z(n16460) );
  NANDN U17119 ( .A(n16367), .B(o[176]), .Z(n16461) );
  XNOR U17120 ( .A(n16460), .B(n16461), .Z(n16440) );
  AND U17121 ( .A(y[1954]), .B(x[239]), .Z(n16369) );
  NAND U17122 ( .A(y[1957]), .B(x[236]), .Z(n16368) );
  XNOR U17123 ( .A(n16369), .B(n16368), .Z(n16415) );
  NAND U17124 ( .A(x[238]), .B(y[1955]), .Z(n16416) );
  XOR U17125 ( .A(n16440), .B(n16439), .Z(n16441) );
  XNOR U17126 ( .A(n16442), .B(n16441), .Z(n16486) );
  NAND U17127 ( .A(n16470), .B(n16370), .Z(n16374) );
  NANDN U17128 ( .A(n16372), .B(n16371), .Z(n16373) );
  AND U17129 ( .A(n16374), .B(n16373), .Z(n16450) );
  NAND U17130 ( .A(x[232]), .B(y[1967]), .Z(n17126) );
  AND U17131 ( .A(x[225]), .B(y[1960]), .Z(n16531) );
  NANDN U17132 ( .A(n17126), .B(n16531), .Z(n16378) );
  NANDN U17133 ( .A(n16376), .B(n16375), .Z(n16377) );
  NAND U17134 ( .A(n16378), .B(n16377), .Z(n16449) );
  XNOR U17135 ( .A(n16450), .B(n16449), .Z(n16452) );
  NANDN U17136 ( .A(n16380), .B(n16379), .Z(n16384) );
  NANDN U17137 ( .A(n16382), .B(n16381), .Z(n16383) );
  AND U17138 ( .A(n16384), .B(n16383), .Z(n16446) );
  AND U17139 ( .A(x[224]), .B(y[1969]), .Z(n16429) );
  NAND U17140 ( .A(x[241]), .B(y[1952]), .Z(n16430) );
  NAND U17141 ( .A(x[240]), .B(y[1953]), .Z(n16426) );
  XOR U17142 ( .A(o[177]), .B(n16426), .Z(n16432) );
  AND U17143 ( .A(y[1967]), .B(x[226]), .Z(n16386) );
  NAND U17144 ( .A(y[1959]), .B(x[234]), .Z(n16385) );
  XNOR U17145 ( .A(n16386), .B(n16385), .Z(n16465) );
  NAND U17146 ( .A(x[227]), .B(y[1966]), .Z(n16466) );
  XOR U17147 ( .A(n16465), .B(n16466), .Z(n16444) );
  XNOR U17148 ( .A(n16443), .B(n16444), .Z(n16445) );
  XNOR U17149 ( .A(n16446), .B(n16445), .Z(n16451) );
  XOR U17150 ( .A(n16452), .B(n16451), .Z(n16485) );
  XOR U17151 ( .A(n16486), .B(n16485), .Z(n16488) );
  XNOR U17152 ( .A(n16487), .B(n16488), .Z(n16410) );
  NAND U17153 ( .A(n16388), .B(n16387), .Z(n16392) );
  NAND U17154 ( .A(n16390), .B(n16389), .Z(n16391) );
  AND U17155 ( .A(n16392), .B(n16391), .Z(n16409) );
  XNOR U17156 ( .A(n16410), .B(n16409), .Z(n16412) );
  XOR U17157 ( .A(n16411), .B(n16412), .Z(n16489) );
  XOR U17158 ( .A(n16490), .B(n16489), .Z(n16491) );
  XOR U17159 ( .A(n16492), .B(n16491), .Z(n16497) );
  NAND U17160 ( .A(n16397), .B(n16396), .Z(n16401) );
  NAND U17161 ( .A(n16399), .B(n16398), .Z(n16400) );
  NAND U17162 ( .A(n16401), .B(n16400), .Z(n16495) );
  XNOR U17163 ( .A(n16496), .B(n16495), .Z(n16402) );
  XNOR U17164 ( .A(n16497), .B(n16402), .Z(N370) );
  NAND U17165 ( .A(n16404), .B(n16403), .Z(n16408) );
  NANDN U17166 ( .A(n16406), .B(n16405), .Z(n16407) );
  AND U17167 ( .A(n16408), .B(n16407), .Z(n16603) );
  NAND U17168 ( .A(n16410), .B(n16409), .Z(n16414) );
  NANDN U17169 ( .A(n16412), .B(n16411), .Z(n16413) );
  AND U17170 ( .A(n16414), .B(n16413), .Z(n16601) );
  AND U17171 ( .A(x[236]), .B(y[1954]), .Z(n16731) );
  AND U17172 ( .A(x[239]), .B(y[1957]), .Z(n16632) );
  NAND U17173 ( .A(n16731), .B(n16632), .Z(n16418) );
  NANDN U17174 ( .A(n16416), .B(n16415), .Z(n16417) );
  NAND U17175 ( .A(n16418), .B(n16417), .Z(n16580) );
  NAND U17176 ( .A(n17605), .B(n16419), .Z(n16423) );
  NANDN U17177 ( .A(n16421), .B(n16420), .Z(n16422) );
  AND U17178 ( .A(n16423), .B(n16422), .Z(n16570) );
  AND U17179 ( .A(y[1969]), .B(x[225]), .Z(n16425) );
  NAND U17180 ( .A(y[1960]), .B(x[234]), .Z(n16424) );
  XNOR U17181 ( .A(n16425), .B(n16424), .Z(n16532) );
  NANDN U17182 ( .A(n16426), .B(o[177]), .Z(n16533) );
  XNOR U17183 ( .A(n16532), .B(n16533), .Z(n16567) );
  AND U17184 ( .A(y[1955]), .B(x[239]), .Z(n16428) );
  NAND U17185 ( .A(y[1961]), .B(x[233]), .Z(n16427) );
  XNOR U17186 ( .A(n16428), .B(n16427), .Z(n16523) );
  NAND U17187 ( .A(x[238]), .B(y[1956]), .Z(n16524) );
  XOR U17188 ( .A(n16523), .B(n16524), .Z(n16568) );
  XNOR U17189 ( .A(n16567), .B(n16568), .Z(n16569) );
  XNOR U17190 ( .A(n16570), .B(n16569), .Z(n16579) );
  XOR U17191 ( .A(n16580), .B(n16579), .Z(n16582) );
  NANDN U17192 ( .A(n16430), .B(n16429), .Z(n16434) );
  NANDN U17193 ( .A(n16432), .B(n16431), .Z(n16433) );
  AND U17194 ( .A(n16434), .B(n16433), .Z(n16592) );
  AND U17195 ( .A(y[1954]), .B(x[240]), .Z(n16436) );
  NAND U17196 ( .A(y[1959]), .B(x[235]), .Z(n16435) );
  XNOR U17197 ( .A(n16436), .B(n16435), .Z(n16519) );
  NAND U17198 ( .A(x[226]), .B(y[1968]), .Z(n16520) );
  XNOR U17199 ( .A(n16519), .B(n16520), .Z(n16591) );
  AND U17200 ( .A(x[229]), .B(y[1965]), .Z(n16640) );
  NAND U17201 ( .A(y[1964]), .B(x[230]), .Z(n16437) );
  XNOR U17202 ( .A(n16640), .B(n16437), .Z(n16515) );
  NAND U17203 ( .A(y[1966]), .B(x[228]), .Z(n16438) );
  XNOR U17204 ( .A(n17272), .B(n16438), .Z(n16554) );
  NAND U17205 ( .A(x[231]), .B(y[1963]), .Z(n16555) );
  XNOR U17206 ( .A(n16515), .B(n16516), .Z(n16593) );
  XOR U17207 ( .A(n16594), .B(n16593), .Z(n16581) );
  XOR U17208 ( .A(n16582), .B(n16581), .Z(n16504) );
  NANDN U17209 ( .A(n16444), .B(n16443), .Z(n16448) );
  NANDN U17210 ( .A(n16446), .B(n16445), .Z(n16447) );
  AND U17211 ( .A(n16448), .B(n16447), .Z(n16574) );
  XOR U17212 ( .A(n16573), .B(n16574), .Z(n16575) );
  NANDN U17213 ( .A(n16450), .B(n16449), .Z(n16454) );
  NAND U17214 ( .A(n16452), .B(n16451), .Z(n16453) );
  AND U17215 ( .A(n16454), .B(n16453), .Z(n16576) );
  XOR U17216 ( .A(n16575), .B(n16576), .Z(n16503) );
  XNOR U17217 ( .A(n16504), .B(n16503), .Z(n16506) );
  AND U17218 ( .A(x[232]), .B(y[1964]), .Z(n16777) );
  NAND U17219 ( .A(n16777), .B(n16455), .Z(n16459) );
  NAND U17220 ( .A(n16457), .B(n16456), .Z(n16458) );
  NAND U17221 ( .A(n16459), .B(n16458), .Z(n16586) );
  NAND U17222 ( .A(x[233]), .B(y[1968]), .Z(n17405) );
  NANDN U17223 ( .A(n17405), .B(n16531), .Z(n16463) );
  NANDN U17224 ( .A(n16461), .B(n16460), .Z(n16462) );
  NAND U17225 ( .A(n16463), .B(n16462), .Z(n16585) );
  XOR U17226 ( .A(n16586), .B(n16585), .Z(n16588) );
  NAND U17227 ( .A(x[234]), .B(y[1967]), .Z(n17406) );
  AND U17228 ( .A(x[224]), .B(y[1970]), .Z(n16536) );
  NAND U17229 ( .A(x[242]), .B(y[1952]), .Z(n16537) );
  XNOR U17230 ( .A(n16536), .B(n16537), .Z(n16538) );
  NAND U17231 ( .A(x[241]), .B(y[1953]), .Z(n16558) );
  XOR U17232 ( .A(o[178]), .B(n16558), .Z(n16539) );
  XNOR U17233 ( .A(n16538), .B(n16539), .Z(n16561) );
  AND U17234 ( .A(y[1957]), .B(x[237]), .Z(n16468) );
  NAND U17235 ( .A(y[1967]), .B(x[227]), .Z(n16467) );
  XNOR U17236 ( .A(n16468), .B(n16467), .Z(n16544) );
  NAND U17237 ( .A(x[236]), .B(y[1958]), .Z(n16545) );
  XOR U17238 ( .A(n16544), .B(n16545), .Z(n16562) );
  XNOR U17239 ( .A(n16561), .B(n16562), .Z(n16563) );
  XNOR U17240 ( .A(n16564), .B(n16563), .Z(n16587) );
  XOR U17241 ( .A(n16588), .B(n16587), .Z(n16508) );
  NAND U17242 ( .A(n16470), .B(n16469), .Z(n16474) );
  NANDN U17243 ( .A(n16472), .B(n16471), .Z(n16473) );
  AND U17244 ( .A(n16474), .B(n16473), .Z(n16507) );
  XNOR U17245 ( .A(n16508), .B(n16507), .Z(n16510) );
  NANDN U17246 ( .A(n16476), .B(n16475), .Z(n16480) );
  NANDN U17247 ( .A(n16478), .B(n16477), .Z(n16479) );
  AND U17248 ( .A(n16480), .B(n16479), .Z(n16509) );
  XOR U17249 ( .A(n16510), .B(n16509), .Z(n16505) );
  XOR U17250 ( .A(n16506), .B(n16505), .Z(n16501) );
  XNOR U17251 ( .A(n16499), .B(n16500), .Z(n16502) );
  XOR U17252 ( .A(n16501), .B(n16502), .Z(n16600) );
  XOR U17253 ( .A(n16601), .B(n16600), .Z(n16602) );
  XNOR U17254 ( .A(n16603), .B(n16602), .Z(n16599) );
  NAND U17255 ( .A(n16490), .B(n16489), .Z(n16494) );
  NANDN U17256 ( .A(n16492), .B(n16491), .Z(n16493) );
  NAND U17257 ( .A(n16494), .B(n16493), .Z(n16597) );
  XOR U17258 ( .A(n16597), .B(n16598), .Z(n16498) );
  XNOR U17259 ( .A(n16599), .B(n16498), .Z(N371) );
  NANDN U17260 ( .A(n16508), .B(n16507), .Z(n16512) );
  NAND U17261 ( .A(n16510), .B(n16509), .Z(n16511) );
  AND U17262 ( .A(n16512), .B(n16511), .Z(n16699) );
  AND U17263 ( .A(x[230]), .B(y[1965]), .Z(n16514) );
  NAND U17264 ( .A(n16514), .B(n16513), .Z(n16518) );
  NANDN U17265 ( .A(n16516), .B(n16515), .Z(n16517) );
  AND U17266 ( .A(n16518), .B(n16517), .Z(n16693) );
  AND U17267 ( .A(x[240]), .B(y[1959]), .Z(n17061) );
  NAND U17268 ( .A(n17061), .B(n16879), .Z(n16522) );
  NANDN U17269 ( .A(n16520), .B(n16519), .Z(n16521) );
  AND U17270 ( .A(n16522), .B(n16521), .Z(n16692) );
  AND U17271 ( .A(x[239]), .B(y[1961]), .Z(n17297) );
  NAND U17272 ( .A(n17297), .B(n16619), .Z(n16526) );
  NANDN U17273 ( .A(n16524), .B(n16523), .Z(n16525) );
  AND U17274 ( .A(n16526), .B(n16525), .Z(n16610) );
  AND U17275 ( .A(y[1970]), .B(x[225]), .Z(n16528) );
  NAND U17276 ( .A(y[1963]), .B(x[232]), .Z(n16527) );
  XNOR U17277 ( .A(n16528), .B(n16527), .Z(n16658) );
  AND U17278 ( .A(y[1958]), .B(x[237]), .Z(n16530) );
  NAND U17279 ( .A(y[1969]), .B(x[226]), .Z(n16529) );
  XNOR U17280 ( .A(n16530), .B(n16529), .Z(n16625) );
  XOR U17281 ( .A(n16608), .B(n16607), .Z(n16609) );
  XOR U17282 ( .A(n16692), .B(n16691), .Z(n16694) );
  XOR U17283 ( .A(n16693), .B(n16694), .Z(n16698) );
  NAND U17284 ( .A(x[234]), .B(y[1969]), .Z(n17688) );
  NANDN U17285 ( .A(n17688), .B(n16531), .Z(n16535) );
  NANDN U17286 ( .A(n16533), .B(n16532), .Z(n16534) );
  AND U17287 ( .A(n16535), .B(n16534), .Z(n16670) );
  NANDN U17288 ( .A(n16537), .B(n16536), .Z(n16541) );
  NANDN U17289 ( .A(n16539), .B(n16538), .Z(n16540) );
  AND U17290 ( .A(n16541), .B(n16540), .Z(n16668) );
  AND U17291 ( .A(y[1955]), .B(x[240]), .Z(n17342) );
  NAND U17292 ( .A(y[1962]), .B(x[233]), .Z(n16542) );
  XNOR U17293 ( .A(n17342), .B(n16542), .Z(n16620) );
  NAND U17294 ( .A(x[239]), .B(y[1956]), .Z(n16621) );
  AND U17295 ( .A(x[237]), .B(y[1967]), .Z(n17872) );
  NANDN U17296 ( .A(n16543), .B(n17872), .Z(n16547) );
  NANDN U17297 ( .A(n16545), .B(n16544), .Z(n16546) );
  AND U17298 ( .A(n16547), .B(n16546), .Z(n16676) );
  AND U17299 ( .A(y[1961]), .B(x[234]), .Z(n16549) );
  NAND U17300 ( .A(y[1954]), .B(x[241]), .Z(n16548) );
  XNOR U17301 ( .A(n16549), .B(n16548), .Z(n16664) );
  AND U17302 ( .A(x[242]), .B(y[1953]), .Z(n16639) );
  XOR U17303 ( .A(o[179]), .B(n16639), .Z(n16663) );
  XOR U17304 ( .A(n16664), .B(n16663), .Z(n16674) );
  NAND U17305 ( .A(y[1968]), .B(x[227]), .Z(n16550) );
  XNOR U17306 ( .A(n16551), .B(n16550), .Z(n16633) );
  XOR U17307 ( .A(n16674), .B(n16673), .Z(n16675) );
  NAND U17308 ( .A(n16553), .B(n16552), .Z(n16557) );
  NANDN U17309 ( .A(n16555), .B(n16554), .Z(n16556) );
  AND U17310 ( .A(n16557), .B(n16556), .Z(n16616) );
  AND U17311 ( .A(x[224]), .B(y[1971]), .Z(n16644) );
  NAND U17312 ( .A(x[243]), .B(y[1952]), .Z(n16645) );
  ANDN U17313 ( .B(o[178]), .A(n16558), .Z(n16646) );
  XOR U17314 ( .A(n16647), .B(n16646), .Z(n16614) );
  AND U17315 ( .A(x[228]), .B(y[1967]), .Z(n16791) );
  AND U17316 ( .A(y[1966]), .B(x[229]), .Z(n16560) );
  NAND U17317 ( .A(y[1965]), .B(x[230]), .Z(n16559) );
  XOR U17318 ( .A(n16560), .B(n16559), .Z(n16641) );
  XOR U17319 ( .A(n16614), .B(n16613), .Z(n16615) );
  XOR U17320 ( .A(n16616), .B(n16615), .Z(n16685) );
  XNOR U17321 ( .A(n16686), .B(n16685), .Z(n16688) );
  XOR U17322 ( .A(n16687), .B(n16688), .Z(n16681) );
  NANDN U17323 ( .A(n16562), .B(n16561), .Z(n16566) );
  NANDN U17324 ( .A(n16564), .B(n16563), .Z(n16565) );
  AND U17325 ( .A(n16566), .B(n16565), .Z(n16680) );
  NANDN U17326 ( .A(n16568), .B(n16567), .Z(n16572) );
  NANDN U17327 ( .A(n16570), .B(n16569), .Z(n16571) );
  NAND U17328 ( .A(n16572), .B(n16571), .Z(n16679) );
  XOR U17329 ( .A(n16680), .B(n16679), .Z(n16682) );
  XOR U17330 ( .A(n16681), .B(n16682), .Z(n16697) );
  XOR U17331 ( .A(n16698), .B(n16697), .Z(n16700) );
  XNOR U17332 ( .A(n16699), .B(n16700), .Z(n16712) );
  NAND U17333 ( .A(n16574), .B(n16573), .Z(n16578) );
  NAND U17334 ( .A(n16576), .B(n16575), .Z(n16577) );
  AND U17335 ( .A(n16578), .B(n16577), .Z(n16710) );
  NAND U17336 ( .A(n16580), .B(n16579), .Z(n16584) );
  NAND U17337 ( .A(n16582), .B(n16581), .Z(n16583) );
  AND U17338 ( .A(n16584), .B(n16583), .Z(n16706) );
  NAND U17339 ( .A(n16586), .B(n16585), .Z(n16590) );
  NAND U17340 ( .A(n16588), .B(n16587), .Z(n16589) );
  AND U17341 ( .A(n16590), .B(n16589), .Z(n16704) );
  NANDN U17342 ( .A(n16592), .B(n16591), .Z(n16596) );
  NAND U17343 ( .A(n16594), .B(n16593), .Z(n16595) );
  NAND U17344 ( .A(n16596), .B(n16595), .Z(n16703) );
  XOR U17345 ( .A(n16710), .B(n16709), .Z(n16711) );
  XOR U17346 ( .A(n16712), .B(n16711), .Z(n16718) );
  XNOR U17347 ( .A(n16719), .B(n16718), .Z(n16721) );
  XOR U17348 ( .A(n16720), .B(n16721), .Z(n16717) );
  NAND U17349 ( .A(n16601), .B(n16600), .Z(n16605) );
  NAND U17350 ( .A(n16603), .B(n16602), .Z(n16604) );
  NAND U17351 ( .A(n16605), .B(n16604), .Z(n16715) );
  XNOR U17352 ( .A(n16716), .B(n16715), .Z(n16606) );
  XNOR U17353 ( .A(n16717), .B(n16606), .Z(N372) );
  NAND U17354 ( .A(n16608), .B(n16607), .Z(n16612) );
  NANDN U17355 ( .A(n16610), .B(n16609), .Z(n16611) );
  AND U17356 ( .A(n16612), .B(n16611), .Z(n16726) );
  NAND U17357 ( .A(n16614), .B(n16613), .Z(n16618) );
  NANDN U17358 ( .A(n16616), .B(n16615), .Z(n16617) );
  NAND U17359 ( .A(n16618), .B(n16617), .Z(n16725) );
  AND U17360 ( .A(x[240]), .B(y[1962]), .Z(n17540) );
  NAND U17361 ( .A(n17540), .B(n16619), .Z(n16623) );
  NANDN U17362 ( .A(n16621), .B(n16620), .Z(n16622) );
  AND U17363 ( .A(n16623), .B(n16622), .Z(n16766) );
  AND U17364 ( .A(x[237]), .B(y[1969]), .Z(n18074) );
  NAND U17365 ( .A(n18074), .B(n16624), .Z(n16628) );
  NANDN U17366 ( .A(n16626), .B(n16625), .Z(n16627) );
  AND U17367 ( .A(n16628), .B(n16627), .Z(n16811) );
  AND U17368 ( .A(y[1956]), .B(x[240]), .Z(n16630) );
  NAND U17369 ( .A(y[1962]), .B(x[234]), .Z(n16629) );
  XNOR U17370 ( .A(n16630), .B(n16629), .Z(n16772) );
  AND U17371 ( .A(x[226]), .B(y[1970]), .Z(n16773) );
  XOR U17372 ( .A(n16772), .B(n16773), .Z(n16809) );
  NAND U17373 ( .A(y[1963]), .B(x[233]), .Z(n16631) );
  XNOR U17374 ( .A(n16632), .B(n16631), .Z(n16742) );
  AND U17375 ( .A(x[238]), .B(y[1958]), .Z(n16743) );
  XOR U17376 ( .A(n16742), .B(n16743), .Z(n16808) );
  XOR U17377 ( .A(n16809), .B(n16808), .Z(n16810) );
  NAND U17378 ( .A(x[235]), .B(y[1968]), .Z(n17690) );
  NANDN U17379 ( .A(n17690), .B(n16906), .Z(n16636) );
  NANDN U17380 ( .A(n16634), .B(n16633), .Z(n16635) );
  AND U17381 ( .A(n16636), .B(n16635), .Z(n16817) );
  AND U17382 ( .A(y[1961]), .B(x[235]), .Z(n16638) );
  NAND U17383 ( .A(y[1971]), .B(x[225]), .Z(n16637) );
  XNOR U17384 ( .A(n16638), .B(n16637), .Z(n16738) );
  AND U17385 ( .A(x[243]), .B(y[1953]), .Z(n16746) );
  XOR U17386 ( .A(o[180]), .B(n16746), .Z(n16737) );
  XOR U17387 ( .A(n16738), .B(n16737), .Z(n16815) );
  AND U17388 ( .A(o[179]), .B(n16639), .Z(n16799) );
  AND U17389 ( .A(x[224]), .B(y[1972]), .Z(n16796) );
  AND U17390 ( .A(x[244]), .B(y[1952]), .Z(n16797) );
  XOR U17391 ( .A(n16796), .B(n16797), .Z(n16798) );
  XOR U17392 ( .A(n16799), .B(n16798), .Z(n16814) );
  XOR U17393 ( .A(n16815), .B(n16814), .Z(n16816) );
  XOR U17394 ( .A(n16768), .B(n16767), .Z(n16727) );
  XOR U17395 ( .A(n16728), .B(n16727), .Z(n16823) );
  AND U17396 ( .A(x[230]), .B(y[1966]), .Z(n16748) );
  IV U17397 ( .A(n16748), .Z(n16656) );
  NANDN U17398 ( .A(n16656), .B(n16640), .Z(n16643) );
  NANDN U17399 ( .A(n16641), .B(n16791), .Z(n16642) );
  AND U17400 ( .A(n16643), .B(n16642), .Z(n16756) );
  NANDN U17401 ( .A(n16645), .B(n16644), .Z(n16649) );
  NAND U17402 ( .A(n16647), .B(n16646), .Z(n16648) );
  AND U17403 ( .A(n16649), .B(n16648), .Z(n16754) );
  AND U17404 ( .A(y[1954]), .B(x[242]), .Z(n16651) );
  NAND U17405 ( .A(y[1960]), .B(x[236]), .Z(n16650) );
  XNOR U17406 ( .A(n16651), .B(n16650), .Z(n16732) );
  AND U17407 ( .A(x[241]), .B(y[1955]), .Z(n16733) );
  XOR U17408 ( .A(n16732), .B(n16733), .Z(n16753) );
  AND U17409 ( .A(y[1959]), .B(x[237]), .Z(n16653) );
  NAND U17410 ( .A(y[1969]), .B(x[227]), .Z(n16652) );
  XNOR U17411 ( .A(n16653), .B(n16652), .Z(n16778) );
  XOR U17412 ( .A(n16778), .B(n16777), .Z(n16750) );
  AND U17413 ( .A(y[1967]), .B(x[229]), .Z(n16655) );
  NAND U17414 ( .A(y[1968]), .B(x[228]), .Z(n16654) );
  XNOR U17415 ( .A(n16655), .B(n16654), .Z(n16793) );
  AND U17416 ( .A(x[231]), .B(y[1965]), .Z(n16792) );
  XNOR U17417 ( .A(n16793), .B(n16792), .Z(n16747) );
  XOR U17418 ( .A(n16656), .B(n16747), .Z(n16749) );
  AND U17419 ( .A(x[232]), .B(y[1970]), .Z(n17842) );
  AND U17420 ( .A(x[225]), .B(y[1963]), .Z(n16657) );
  NAND U17421 ( .A(n17842), .B(n16657), .Z(n16661) );
  NANDN U17422 ( .A(n16659), .B(n16658), .Z(n16660) );
  AND U17423 ( .A(n16661), .B(n16660), .Z(n16803) );
  AND U17424 ( .A(x[241]), .B(y[1961]), .Z(n17545) );
  NAND U17425 ( .A(n17545), .B(n16662), .Z(n16666) );
  NAND U17426 ( .A(n16664), .B(n16663), .Z(n16665) );
  NAND U17427 ( .A(n16666), .B(n16665), .Z(n16802) );
  XNOR U17428 ( .A(n16804), .B(n16805), .Z(n16759) );
  XOR U17429 ( .A(n16760), .B(n16759), .Z(n16761) );
  NANDN U17430 ( .A(n16668), .B(n16667), .Z(n16672) );
  NANDN U17431 ( .A(n16670), .B(n16669), .Z(n16671) );
  NAND U17432 ( .A(n16672), .B(n16671), .Z(n16762) );
  NAND U17433 ( .A(n16674), .B(n16673), .Z(n16678) );
  NANDN U17434 ( .A(n16676), .B(n16675), .Z(n16677) );
  NAND U17435 ( .A(n16678), .B(n16677), .Z(n16821) );
  NANDN U17436 ( .A(n16680), .B(n16679), .Z(n16684) );
  NANDN U17437 ( .A(n16682), .B(n16681), .Z(n16683) );
  AND U17438 ( .A(n16684), .B(n16683), .Z(n16835) );
  NAND U17439 ( .A(n16686), .B(n16685), .Z(n16690) );
  NANDN U17440 ( .A(n16688), .B(n16687), .Z(n16689) );
  AND U17441 ( .A(n16690), .B(n16689), .Z(n16833) );
  NANDN U17442 ( .A(n16692), .B(n16691), .Z(n16696) );
  OR U17443 ( .A(n16694), .B(n16693), .Z(n16695) );
  AND U17444 ( .A(n16696), .B(n16695), .Z(n16832) );
  XNOR U17445 ( .A(n16833), .B(n16832), .Z(n16834) );
  XNOR U17446 ( .A(n16835), .B(n16834), .Z(n16826) );
  XOR U17447 ( .A(n16827), .B(n16826), .Z(n16829) );
  NANDN U17448 ( .A(n16698), .B(n16697), .Z(n16702) );
  OR U17449 ( .A(n16700), .B(n16699), .Z(n16701) );
  AND U17450 ( .A(n16702), .B(n16701), .Z(n16828) );
  XOR U17451 ( .A(n16829), .B(n16828), .Z(n16845) );
  NANDN U17452 ( .A(n16704), .B(n16703), .Z(n16708) );
  NANDN U17453 ( .A(n16706), .B(n16705), .Z(n16707) );
  AND U17454 ( .A(n16708), .B(n16707), .Z(n16842) );
  NAND U17455 ( .A(n16710), .B(n16709), .Z(n16714) );
  NAND U17456 ( .A(n16712), .B(n16711), .Z(n16713) );
  AND U17457 ( .A(n16714), .B(n16713), .Z(n16843) );
  XOR U17458 ( .A(n16842), .B(n16843), .Z(n16844) );
  XOR U17459 ( .A(n16845), .B(n16844), .Z(n16841) );
  NAND U17460 ( .A(n16719), .B(n16718), .Z(n16723) );
  NANDN U17461 ( .A(n16721), .B(n16720), .Z(n16722) );
  AND U17462 ( .A(n16723), .B(n16722), .Z(n16840) );
  IV U17463 ( .A(n16840), .Z(n16838) );
  XOR U17464 ( .A(n16839), .B(n16838), .Z(n16724) );
  XNOR U17465 ( .A(n16841), .B(n16724), .Z(N373) );
  NANDN U17466 ( .A(n16726), .B(n16725), .Z(n16730) );
  NAND U17467 ( .A(n16728), .B(n16727), .Z(n16729) );
  AND U17468 ( .A(n16730), .B(n16729), .Z(n16858) );
  AND U17469 ( .A(x[242]), .B(y[1960]), .Z(n17544) );
  NAND U17470 ( .A(n17544), .B(n16731), .Z(n16735) );
  NAND U17471 ( .A(n16733), .B(n16732), .Z(n16734) );
  NAND U17472 ( .A(n16735), .B(n16734), .Z(n16935) );
  NAND U17473 ( .A(x[235]), .B(y[1971]), .Z(n18234) );
  AND U17474 ( .A(x[225]), .B(y[1961]), .Z(n16736) );
  NANDN U17475 ( .A(n18234), .B(n16736), .Z(n16740) );
  NAND U17476 ( .A(n16738), .B(n16737), .Z(n16739) );
  NAND U17477 ( .A(n16740), .B(n16739), .Z(n16934) );
  XOR U17478 ( .A(n16935), .B(n16934), .Z(n16937) );
  AND U17479 ( .A(x[239]), .B(y[1963]), .Z(n17534) );
  NAND U17480 ( .A(n17534), .B(n16741), .Z(n16745) );
  NAND U17481 ( .A(n16743), .B(n16742), .Z(n16744) );
  NAND U17482 ( .A(n16745), .B(n16744), .Z(n16893) );
  AND U17483 ( .A(o[180]), .B(n16746), .Z(n16915) );
  AND U17484 ( .A(x[224]), .B(y[1973]), .Z(n16912) );
  AND U17485 ( .A(x[245]), .B(y[1952]), .Z(n16913) );
  XOR U17486 ( .A(n16912), .B(n16913), .Z(n16914) );
  XOR U17487 ( .A(n16915), .B(n16914), .Z(n16891) );
  AND U17488 ( .A(x[229]), .B(y[1968]), .Z(n16899) );
  AND U17489 ( .A(x[240]), .B(y[1957]), .Z(n16898) );
  XOR U17490 ( .A(n16899), .B(n16898), .Z(n16897) );
  AND U17491 ( .A(x[239]), .B(y[1958]), .Z(n16896) );
  XOR U17492 ( .A(n16897), .B(n16896), .Z(n16890) );
  XOR U17493 ( .A(n16891), .B(n16890), .Z(n16892) );
  XOR U17494 ( .A(n16893), .B(n16892), .Z(n16936) );
  XOR U17495 ( .A(n16937), .B(n16936), .Z(n16929) );
  NANDN U17496 ( .A(n16748), .B(n16747), .Z(n16752) );
  NANDN U17497 ( .A(n16750), .B(n16749), .Z(n16751) );
  NAND U17498 ( .A(n16752), .B(n16751), .Z(n16928) );
  NANDN U17499 ( .A(n16754), .B(n16753), .Z(n16758) );
  NANDN U17500 ( .A(n16756), .B(n16755), .Z(n16757) );
  AND U17501 ( .A(n16758), .B(n16757), .Z(n16930) );
  XOR U17502 ( .A(n16931), .B(n16930), .Z(n16856) );
  NAND U17503 ( .A(n16760), .B(n16759), .Z(n16764) );
  NANDN U17504 ( .A(n16762), .B(n16761), .Z(n16763) );
  AND U17505 ( .A(n16764), .B(n16763), .Z(n16855) );
  NANDN U17506 ( .A(n16766), .B(n16765), .Z(n16770) );
  NAND U17507 ( .A(n16768), .B(n16767), .Z(n16769) );
  AND U17508 ( .A(n16770), .B(n16769), .Z(n16955) );
  NAND U17509 ( .A(n17540), .B(n16771), .Z(n16775) );
  NAND U17510 ( .A(n16773), .B(n16772), .Z(n16774) );
  NAND U17511 ( .A(n16775), .B(n16774), .Z(n16862) );
  NAND U17512 ( .A(n18074), .B(n16776), .Z(n16780) );
  NAND U17513 ( .A(n16778), .B(n16777), .Z(n16779) );
  NAND U17514 ( .A(n16780), .B(n16779), .Z(n16949) );
  AND U17515 ( .A(y[1954]), .B(x[243]), .Z(n16782) );
  NAND U17516 ( .A(y[1962]), .B(x[235]), .Z(n16781) );
  XNOR U17517 ( .A(n16782), .B(n16781), .Z(n16881) );
  AND U17518 ( .A(x[244]), .B(y[1953]), .Z(n16911) );
  XOR U17519 ( .A(o[181]), .B(n16911), .Z(n16880) );
  XOR U17520 ( .A(n16881), .B(n16880), .Z(n16947) );
  AND U17521 ( .A(y[1955]), .B(x[242]), .Z(n16784) );
  NAND U17522 ( .A(y[1963]), .B(x[234]), .Z(n16783) );
  XNOR U17523 ( .A(n16784), .B(n16783), .Z(n16919) );
  AND U17524 ( .A(x[225]), .B(y[1972]), .Z(n16920) );
  XOR U17525 ( .A(n16919), .B(n16920), .Z(n16946) );
  XOR U17526 ( .A(n16947), .B(n16946), .Z(n16948) );
  XOR U17527 ( .A(n16949), .B(n16948), .Z(n16861) );
  XOR U17528 ( .A(n16862), .B(n16861), .Z(n16864) );
  AND U17529 ( .A(x[231]), .B(y[1966]), .Z(n17124) );
  AND U17530 ( .A(y[1967]), .B(x[230]), .Z(n16786) );
  NAND U17531 ( .A(y[1959]), .B(x[238]), .Z(n16785) );
  XNOR U17532 ( .A(n16786), .B(n16785), .Z(n16923) );
  XNOR U17533 ( .A(n17124), .B(n16923), .Z(n16870) );
  NAND U17534 ( .A(x[233]), .B(y[1964]), .Z(n16868) );
  NAND U17535 ( .A(x[232]), .B(y[1965]), .Z(n16867) );
  XOR U17536 ( .A(n16868), .B(n16867), .Z(n16869) );
  XNOR U17537 ( .A(n16870), .B(n16869), .Z(n16886) );
  AND U17538 ( .A(y[1961]), .B(x[236]), .Z(n16788) );
  NAND U17539 ( .A(y[1956]), .B(x[241]), .Z(n16787) );
  XNOR U17540 ( .A(n16788), .B(n16787), .Z(n16873) );
  AND U17541 ( .A(x[226]), .B(y[1971]), .Z(n16874) );
  XOR U17542 ( .A(n16873), .B(n16874), .Z(n16885) );
  AND U17543 ( .A(y[1960]), .B(x[237]), .Z(n16790) );
  NAND U17544 ( .A(y[1970]), .B(x[227]), .Z(n16789) );
  XNOR U17545 ( .A(n16790), .B(n16789), .Z(n16907) );
  AND U17546 ( .A(x[228]), .B(y[1969]), .Z(n16908) );
  XOR U17547 ( .A(n16907), .B(n16908), .Z(n16884) );
  XOR U17548 ( .A(n16885), .B(n16884), .Z(n16887) );
  XOR U17549 ( .A(n16886), .B(n16887), .Z(n16943) );
  NAND U17550 ( .A(n16899), .B(n16791), .Z(n16795) );
  NAND U17551 ( .A(n16793), .B(n16792), .Z(n16794) );
  NAND U17552 ( .A(n16795), .B(n16794), .Z(n16941) );
  NAND U17553 ( .A(n16797), .B(n16796), .Z(n16801) );
  NAND U17554 ( .A(n16799), .B(n16798), .Z(n16800) );
  NAND U17555 ( .A(n16801), .B(n16800), .Z(n16940) );
  XOR U17556 ( .A(n16941), .B(n16940), .Z(n16942) );
  XOR U17557 ( .A(n16943), .B(n16942), .Z(n16863) );
  XOR U17558 ( .A(n16864), .B(n16863), .Z(n16953) );
  NANDN U17559 ( .A(n16803), .B(n16802), .Z(n16807) );
  NAND U17560 ( .A(n16805), .B(n16804), .Z(n16806) );
  NAND U17561 ( .A(n16807), .B(n16806), .Z(n16960) );
  NAND U17562 ( .A(n16809), .B(n16808), .Z(n16813) );
  NANDN U17563 ( .A(n16811), .B(n16810), .Z(n16812) );
  NAND U17564 ( .A(n16813), .B(n16812), .Z(n16959) );
  NAND U17565 ( .A(n16815), .B(n16814), .Z(n16819) );
  NANDN U17566 ( .A(n16817), .B(n16816), .Z(n16818) );
  NAND U17567 ( .A(n16819), .B(n16818), .Z(n16958) );
  XOR U17568 ( .A(n16959), .B(n16958), .Z(n16961) );
  XOR U17569 ( .A(n16960), .B(n16961), .Z(n16952) );
  XOR U17570 ( .A(n16953), .B(n16952), .Z(n16954) );
  NANDN U17571 ( .A(n16821), .B(n16820), .Z(n16825) );
  NANDN U17572 ( .A(n16823), .B(n16822), .Z(n16824) );
  NAND U17573 ( .A(n16825), .B(n16824), .Z(n16849) );
  XOR U17574 ( .A(n16850), .B(n16849), .Z(n16852) );
  XNOR U17575 ( .A(n16851), .B(n16852), .Z(n16969) );
  NAND U17576 ( .A(n16827), .B(n16826), .Z(n16831) );
  NAND U17577 ( .A(n16829), .B(n16828), .Z(n16830) );
  AND U17578 ( .A(n16831), .B(n16830), .Z(n16968) );
  NANDN U17579 ( .A(n16833), .B(n16832), .Z(n16837) );
  NAND U17580 ( .A(n16835), .B(n16834), .Z(n16836) );
  AND U17581 ( .A(n16837), .B(n16836), .Z(n16967) );
  XOR U17582 ( .A(n16968), .B(n16967), .Z(n16970) );
  XOR U17583 ( .A(n16969), .B(n16970), .Z(n16966) );
  NAND U17584 ( .A(n16843), .B(n16842), .Z(n16847) );
  NANDN U17585 ( .A(n16845), .B(n16844), .Z(n16846) );
  AND U17586 ( .A(n16847), .B(n16846), .Z(n16965) );
  XOR U17587 ( .A(n16964), .B(n16965), .Z(n16848) );
  XNOR U17588 ( .A(n16966), .B(n16848), .Z(N374) );
  NAND U17589 ( .A(n16850), .B(n16849), .Z(n16854) );
  NAND U17590 ( .A(n16852), .B(n16851), .Z(n16853) );
  AND U17591 ( .A(n16854), .B(n16853), .Z(n16977) );
  NANDN U17592 ( .A(n16856), .B(n16855), .Z(n16860) );
  NANDN U17593 ( .A(n16858), .B(n16857), .Z(n16859) );
  AND U17594 ( .A(n16860), .B(n16859), .Z(n16975) );
  NAND U17595 ( .A(n16862), .B(n16861), .Z(n16866) );
  NAND U17596 ( .A(n16864), .B(n16863), .Z(n16865) );
  NAND U17597 ( .A(n16866), .B(n16865), .Z(n17100) );
  NAND U17598 ( .A(n16868), .B(n16867), .Z(n16872) );
  NAND U17599 ( .A(n16870), .B(n16869), .Z(n16871) );
  NAND U17600 ( .A(n16872), .B(n16871), .Z(n17094) );
  NAND U17601 ( .A(n17545), .B(n17045), .Z(n16876) );
  NAND U17602 ( .A(n16874), .B(n16873), .Z(n16875) );
  NAND U17603 ( .A(n16876), .B(n16875), .Z(n17021) );
  AND U17604 ( .A(x[229]), .B(y[1969]), .Z(n17067) );
  AND U17605 ( .A(x[241]), .B(y[1957]), .Z(n17068) );
  XOR U17606 ( .A(n17067), .B(n17068), .Z(n17069) );
  AND U17607 ( .A(x[240]), .B(y[1958]), .Z(n17070) );
  XOR U17608 ( .A(n17069), .B(n17070), .Z(n17020) );
  AND U17609 ( .A(y[1956]), .B(x[242]), .Z(n16878) );
  NAND U17610 ( .A(y[1962]), .B(x[236]), .Z(n16877) );
  XNOR U17611 ( .A(n16878), .B(n16877), .Z(n17046) );
  AND U17612 ( .A(x[228]), .B(y[1970]), .Z(n17047) );
  XOR U17613 ( .A(n17046), .B(n17047), .Z(n17019) );
  XOR U17614 ( .A(n17020), .B(n17019), .Z(n17022) );
  XNOR U17615 ( .A(n17021), .B(n17022), .Z(n17091) );
  NAND U17616 ( .A(x[243]), .B(y[1962]), .Z(n17980) );
  NANDN U17617 ( .A(n17980), .B(n16879), .Z(n16883) );
  NAND U17618 ( .A(n16881), .B(n16880), .Z(n16882) );
  AND U17619 ( .A(n16883), .B(n16882), .Z(n17092) );
  XOR U17620 ( .A(n17091), .B(n17092), .Z(n17093) );
  XNOR U17621 ( .A(n17094), .B(n17093), .Z(n17097) );
  NAND U17622 ( .A(n16885), .B(n16884), .Z(n16889) );
  NAND U17623 ( .A(n16887), .B(n16886), .Z(n16888) );
  NAND U17624 ( .A(n16889), .B(n16888), .Z(n17080) );
  NAND U17625 ( .A(n16891), .B(n16890), .Z(n16895) );
  NAND U17626 ( .A(n16893), .B(n16892), .Z(n16894) );
  NAND U17627 ( .A(n16895), .B(n16894), .Z(n17079) );
  XOR U17628 ( .A(n17080), .B(n17079), .Z(n17082) );
  AND U17629 ( .A(n16897), .B(n16896), .Z(n16901) );
  NAND U17630 ( .A(n16899), .B(n16898), .Z(n16900) );
  NANDN U17631 ( .A(n16901), .B(n16900), .Z(n17042) );
  AND U17632 ( .A(y[1961]), .B(x[237]), .Z(n16903) );
  NAND U17633 ( .A(y[1954]), .B(x[244]), .Z(n16902) );
  XNOR U17634 ( .A(n16903), .B(n16902), .Z(n17063) );
  AND U17635 ( .A(x[226]), .B(y[1972]), .Z(n17064) );
  XOR U17636 ( .A(n17063), .B(n17064), .Z(n17040) );
  AND U17637 ( .A(y[1968]), .B(x[230]), .Z(n16905) );
  NAND U17638 ( .A(y[1959]), .B(x[239]), .Z(n16904) );
  XNOR U17639 ( .A(n16905), .B(n16904), .Z(n17075) );
  XOR U17640 ( .A(n17040), .B(n17039), .Z(n17041) );
  XOR U17641 ( .A(n17042), .B(n17041), .Z(n17086) );
  AND U17642 ( .A(x[237]), .B(y[1970]), .Z(n18235) );
  NAND U17643 ( .A(n16906), .B(n18235), .Z(n16910) );
  NAND U17644 ( .A(n16908), .B(n16907), .Z(n16909) );
  NAND U17645 ( .A(n16910), .B(n16909), .Z(n17010) );
  AND U17646 ( .A(x[225]), .B(y[1973]), .Z(n17033) );
  XOR U17647 ( .A(n17034), .B(n17033), .Z(n17032) );
  AND U17648 ( .A(o[181]), .B(n16911), .Z(n17031) );
  XOR U17649 ( .A(n17032), .B(n17031), .Z(n17008) );
  AND U17650 ( .A(x[238]), .B(y[1960]), .Z(n17025) );
  AND U17651 ( .A(x[227]), .B(y[1971]), .Z(n17026) );
  XOR U17652 ( .A(n17025), .B(n17026), .Z(n17027) );
  AND U17653 ( .A(x[243]), .B(y[1955]), .Z(n17028) );
  XOR U17654 ( .A(n17027), .B(n17028), .Z(n17007) );
  XOR U17655 ( .A(n17008), .B(n17007), .Z(n17009) );
  XOR U17656 ( .A(n17010), .B(n17009), .Z(n17085) );
  XOR U17657 ( .A(n17086), .B(n17085), .Z(n17088) );
  NAND U17658 ( .A(n16913), .B(n16912), .Z(n16917) );
  NAND U17659 ( .A(n16915), .B(n16914), .Z(n16916) );
  NAND U17660 ( .A(n16917), .B(n16916), .Z(n17002) );
  AND U17661 ( .A(x[242]), .B(y[1963]), .Z(n17982) );
  NAND U17662 ( .A(n17982), .B(n16918), .Z(n16922) );
  NAND U17663 ( .A(n16920), .B(n16919), .Z(n16921) );
  NAND U17664 ( .A(n16922), .B(n16921), .Z(n17001) );
  XOR U17665 ( .A(n17002), .B(n17001), .Z(n17004) );
  AND U17666 ( .A(x[238]), .B(y[1967]), .Z(n18021) );
  NAND U17667 ( .A(n18021), .B(n17074), .Z(n16925) );
  NAND U17668 ( .A(n17124), .B(n16923), .Z(n16924) );
  NAND U17669 ( .A(n16925), .B(n16924), .Z(n17016) );
  AND U17670 ( .A(x[224]), .B(y[1974]), .Z(n17050) );
  AND U17671 ( .A(x[246]), .B(y[1952]), .Z(n17051) );
  XOR U17672 ( .A(n17050), .B(n17051), .Z(n17053) );
  AND U17673 ( .A(x[245]), .B(y[1953]), .Z(n17073) );
  XOR U17674 ( .A(o[182]), .B(n17073), .Z(n17052) );
  XOR U17675 ( .A(n17053), .B(n17052), .Z(n17014) );
  AND U17676 ( .A(y[1967]), .B(x[231]), .Z(n16927) );
  NAND U17677 ( .A(y[1966]), .B(x[232]), .Z(n16926) );
  XNOR U17678 ( .A(n16927), .B(n16926), .Z(n17056) );
  XOR U17679 ( .A(n17014), .B(n17013), .Z(n17015) );
  XOR U17680 ( .A(n17016), .B(n17015), .Z(n17003) );
  XOR U17681 ( .A(n17004), .B(n17003), .Z(n17087) );
  XOR U17682 ( .A(n17088), .B(n17087), .Z(n17081) );
  XOR U17683 ( .A(n17082), .B(n17081), .Z(n17098) );
  XOR U17684 ( .A(n17097), .B(n17098), .Z(n17099) );
  XOR U17685 ( .A(n17100), .B(n17099), .Z(n16992) );
  NANDN U17686 ( .A(n16929), .B(n16928), .Z(n16933) );
  NAND U17687 ( .A(n16931), .B(n16930), .Z(n16932) );
  NAND U17688 ( .A(n16933), .B(n16932), .Z(n16990) );
  NAND U17689 ( .A(n16935), .B(n16934), .Z(n16939) );
  NAND U17690 ( .A(n16937), .B(n16936), .Z(n16938) );
  AND U17691 ( .A(n16939), .B(n16938), .Z(n16998) );
  NAND U17692 ( .A(n16941), .B(n16940), .Z(n16945) );
  NAND U17693 ( .A(n16943), .B(n16942), .Z(n16944) );
  NAND U17694 ( .A(n16945), .B(n16944), .Z(n16996) );
  NAND U17695 ( .A(n16947), .B(n16946), .Z(n16951) );
  NAND U17696 ( .A(n16949), .B(n16948), .Z(n16950) );
  NAND U17697 ( .A(n16951), .B(n16950), .Z(n16995) );
  XOR U17698 ( .A(n16996), .B(n16995), .Z(n16997) );
  XOR U17699 ( .A(n16998), .B(n16997), .Z(n16989) );
  XOR U17700 ( .A(n16990), .B(n16989), .Z(n16991) );
  NAND U17701 ( .A(n16953), .B(n16952), .Z(n16957) );
  NANDN U17702 ( .A(n16955), .B(n16954), .Z(n16956) );
  NAND U17703 ( .A(n16957), .B(n16956), .Z(n16984) );
  NAND U17704 ( .A(n16959), .B(n16958), .Z(n16963) );
  NAND U17705 ( .A(n16961), .B(n16960), .Z(n16962) );
  NAND U17706 ( .A(n16963), .B(n16962), .Z(n16983) );
  XOR U17707 ( .A(n16984), .B(n16983), .Z(n16985) );
  XNOR U17708 ( .A(n16977), .B(n16976), .Z(n16980) );
  NANDN U17709 ( .A(n16968), .B(n16967), .Z(n16972) );
  NANDN U17710 ( .A(n16970), .B(n16969), .Z(n16971) );
  AND U17711 ( .A(n16972), .B(n16971), .Z(n16982) );
  XOR U17712 ( .A(n16981), .B(n16982), .Z(n16973) );
  XNOR U17713 ( .A(n16980), .B(n16973), .Z(N375) );
  NANDN U17714 ( .A(n16975), .B(n16974), .Z(n16979) );
  NAND U17715 ( .A(n16977), .B(n16976), .Z(n16978) );
  NAND U17716 ( .A(n16979), .B(n16978), .Z(n17237) );
  IV U17717 ( .A(n17237), .Z(n17236) );
  NAND U17718 ( .A(n16984), .B(n16983), .Z(n16988) );
  NANDN U17719 ( .A(n16986), .B(n16985), .Z(n16987) );
  AND U17720 ( .A(n16988), .B(n16987), .Z(n17245) );
  NAND U17721 ( .A(n16990), .B(n16989), .Z(n16994) );
  NANDN U17722 ( .A(n16992), .B(n16991), .Z(n16993) );
  NAND U17723 ( .A(n16994), .B(n16993), .Z(n17243) );
  NAND U17724 ( .A(n16996), .B(n16995), .Z(n17000) );
  NANDN U17725 ( .A(n16998), .B(n16997), .Z(n16999) );
  NAND U17726 ( .A(n17000), .B(n16999), .Z(n17221) );
  NAND U17727 ( .A(n17002), .B(n17001), .Z(n17006) );
  NAND U17728 ( .A(n17004), .B(n17003), .Z(n17005) );
  NAND U17729 ( .A(n17006), .B(n17005), .Z(n17214) );
  NAND U17730 ( .A(n17008), .B(n17007), .Z(n17012) );
  NAND U17731 ( .A(n17010), .B(n17009), .Z(n17011) );
  NAND U17732 ( .A(n17012), .B(n17011), .Z(n17212) );
  NAND U17733 ( .A(n17014), .B(n17013), .Z(n17018) );
  NAND U17734 ( .A(n17016), .B(n17015), .Z(n17017) );
  NAND U17735 ( .A(n17018), .B(n17017), .Z(n17211) );
  XOR U17736 ( .A(n17212), .B(n17211), .Z(n17213) );
  XOR U17737 ( .A(n17214), .B(n17213), .Z(n17233) );
  NAND U17738 ( .A(n17020), .B(n17019), .Z(n17024) );
  NAND U17739 ( .A(n17022), .B(n17021), .Z(n17023) );
  NAND U17740 ( .A(n17024), .B(n17023), .Z(n17231) );
  NAND U17741 ( .A(n17026), .B(n17025), .Z(n17030) );
  NAND U17742 ( .A(n17028), .B(n17027), .Z(n17029) );
  NAND U17743 ( .A(n17030), .B(n17029), .Z(n17158) );
  AND U17744 ( .A(n17032), .B(n17031), .Z(n17036) );
  NAND U17745 ( .A(n17034), .B(n17033), .Z(n17035) );
  NANDN U17746 ( .A(n17036), .B(n17035), .Z(n17157) );
  XOR U17747 ( .A(n17158), .B(n17157), .Z(n17160) );
  AND U17748 ( .A(y[1968]), .B(x[231]), .Z(n17038) );
  NAND U17749 ( .A(y[1966]), .B(x[233]), .Z(n17037) );
  XNOR U17750 ( .A(n17038), .B(n17037), .Z(n17125) );
  NAND U17751 ( .A(x[234]), .B(y[1965]), .Z(n17164) );
  AND U17752 ( .A(x[230]), .B(y[1969]), .Z(n17116) );
  NAND U17753 ( .A(x[239]), .B(y[1960]), .Z(n17117) );
  XNOR U17754 ( .A(n17116), .B(n17117), .Z(n17118) );
  NAND U17755 ( .A(x[235]), .B(y[1964]), .Z(n17119) );
  XOR U17756 ( .A(n17118), .B(n17119), .Z(n17166) );
  XOR U17757 ( .A(n17160), .B(n17159), .Z(n17230) );
  XOR U17758 ( .A(n17231), .B(n17230), .Z(n17232) );
  XOR U17759 ( .A(n17233), .B(n17232), .Z(n17219) );
  NAND U17760 ( .A(n17040), .B(n17039), .Z(n17044) );
  NAND U17761 ( .A(n17042), .B(n17041), .Z(n17043) );
  NAND U17762 ( .A(n17044), .B(n17043), .Z(n17152) );
  AND U17763 ( .A(x[242]), .B(y[1962]), .Z(n17864) );
  NAND U17764 ( .A(n17864), .B(n17045), .Z(n17049) );
  NAND U17765 ( .A(n17047), .B(n17046), .Z(n17048) );
  NAND U17766 ( .A(n17049), .B(n17048), .Z(n17188) );
  NAND U17767 ( .A(n17051), .B(n17050), .Z(n17055) );
  NAND U17768 ( .A(n17053), .B(n17052), .Z(n17054) );
  NAND U17769 ( .A(n17055), .B(n17054), .Z(n17187) );
  XOR U17770 ( .A(n17188), .B(n17187), .Z(n17189) );
  NANDN U17771 ( .A(n17126), .B(n17124), .Z(n17059) );
  NANDN U17772 ( .A(n17057), .B(n17056), .Z(n17058) );
  NAND U17773 ( .A(n17059), .B(n17058), .Z(n17201) );
  AND U17774 ( .A(x[224]), .B(y[1975]), .Z(n17135) );
  NAND U17775 ( .A(x[247]), .B(y[1952]), .Z(n17136) );
  NAND U17776 ( .A(x[246]), .B(y[1953]), .Z(n17115) );
  XOR U17777 ( .A(o[183]), .B(n17115), .Z(n17138) );
  NAND U17778 ( .A(y[1955]), .B(x[244]), .Z(n17060) );
  XNOR U17779 ( .A(n17061), .B(n17060), .Z(n17111) );
  NAND U17780 ( .A(x[243]), .B(y[1956]), .Z(n17112) );
  XNOR U17781 ( .A(n17111), .B(n17112), .Z(n17199) );
  XOR U17782 ( .A(n17200), .B(n17199), .Z(n17202) );
  XOR U17783 ( .A(n17201), .B(n17202), .Z(n17190) );
  XOR U17784 ( .A(n17189), .B(n17190), .Z(n17151) );
  XOR U17785 ( .A(n17152), .B(n17151), .Z(n17154) );
  NAND U17786 ( .A(x[244]), .B(y[1961]), .Z(n18030) );
  AND U17787 ( .A(x[237]), .B(y[1954]), .Z(n17062) );
  NANDN U17788 ( .A(n18030), .B(n17062), .Z(n17066) );
  NAND U17789 ( .A(n17064), .B(n17063), .Z(n17065) );
  NAND U17790 ( .A(n17066), .B(n17065), .Z(n17146) );
  NAND U17791 ( .A(n17068), .B(n17067), .Z(n17072) );
  NAND U17792 ( .A(n17070), .B(n17069), .Z(n17071) );
  NAND U17793 ( .A(n17072), .B(n17071), .Z(n17207) );
  AND U17794 ( .A(x[237]), .B(y[1962]), .Z(n17181) );
  AND U17795 ( .A(x[226]), .B(y[1973]), .Z(n17182) );
  XOR U17796 ( .A(n17181), .B(n17182), .Z(n17183) );
  AND U17797 ( .A(x[245]), .B(y[1954]), .Z(n17184) );
  XOR U17798 ( .A(n17183), .B(n17184), .Z(n17206) );
  AND U17799 ( .A(x[236]), .B(y[1963]), .Z(n17129) );
  AND U17800 ( .A(x[225]), .B(y[1974]), .Z(n17130) );
  XOR U17801 ( .A(n17129), .B(n17130), .Z(n17132) );
  AND U17802 ( .A(o[182]), .B(n17073), .Z(n17131) );
  XOR U17803 ( .A(n17132), .B(n17131), .Z(n17205) );
  XOR U17804 ( .A(n17206), .B(n17205), .Z(n17208) );
  XOR U17805 ( .A(n17207), .B(n17208), .Z(n17145) );
  XOR U17806 ( .A(n17146), .B(n17145), .Z(n17148) );
  AND U17807 ( .A(x[239]), .B(y[1968]), .Z(n18224) );
  NAND U17808 ( .A(n17074), .B(n18224), .Z(n17078) );
  NANDN U17809 ( .A(n17076), .B(n17075), .Z(n17077) );
  NAND U17810 ( .A(n17078), .B(n17077), .Z(n17195) );
  AND U17811 ( .A(x[238]), .B(y[1961]), .Z(n17175) );
  AND U17812 ( .A(x[227]), .B(y[1972]), .Z(n17176) );
  XOR U17813 ( .A(n17175), .B(n17176), .Z(n17177) );
  AND U17814 ( .A(x[228]), .B(y[1971]), .Z(n17178) );
  XOR U17815 ( .A(n17177), .B(n17178), .Z(n17194) );
  AND U17816 ( .A(x[229]), .B(y[1970]), .Z(n17169) );
  NAND U17817 ( .A(x[242]), .B(y[1957]), .Z(n17170) );
  XNOR U17818 ( .A(n17169), .B(n17170), .Z(n17172) );
  AND U17819 ( .A(x[241]), .B(y[1958]), .Z(n17171) );
  XOR U17820 ( .A(n17172), .B(n17171), .Z(n17193) );
  XOR U17821 ( .A(n17194), .B(n17193), .Z(n17196) );
  XOR U17822 ( .A(n17195), .B(n17196), .Z(n17147) );
  XOR U17823 ( .A(n17148), .B(n17147), .Z(n17153) );
  XOR U17824 ( .A(n17154), .B(n17153), .Z(n17218) );
  XOR U17825 ( .A(n17219), .B(n17218), .Z(n17220) );
  XNOR U17826 ( .A(n17221), .B(n17220), .Z(n17106) );
  NAND U17827 ( .A(n17080), .B(n17079), .Z(n17084) );
  NAND U17828 ( .A(n17082), .B(n17081), .Z(n17083) );
  NAND U17829 ( .A(n17084), .B(n17083), .Z(n17227) );
  NAND U17830 ( .A(n17086), .B(n17085), .Z(n17090) );
  NAND U17831 ( .A(n17088), .B(n17087), .Z(n17089) );
  NAND U17832 ( .A(n17090), .B(n17089), .Z(n17225) );
  NAND U17833 ( .A(n17092), .B(n17091), .Z(n17096) );
  NAND U17834 ( .A(n17094), .B(n17093), .Z(n17095) );
  AND U17835 ( .A(n17096), .B(n17095), .Z(n17224) );
  XOR U17836 ( .A(n17225), .B(n17224), .Z(n17226) );
  XNOR U17837 ( .A(n17227), .B(n17226), .Z(n17104) );
  NAND U17838 ( .A(n17098), .B(n17097), .Z(n17102) );
  NAND U17839 ( .A(n17100), .B(n17099), .Z(n17101) );
  AND U17840 ( .A(n17102), .B(n17101), .Z(n17105) );
  XOR U17841 ( .A(n17104), .B(n17105), .Z(n17107) );
  XNOR U17842 ( .A(n17106), .B(n17107), .Z(n17244) );
  XNOR U17843 ( .A(n17245), .B(n17246), .Z(n17239) );
  XNOR U17844 ( .A(n17238), .B(n17239), .Z(n17103) );
  XOR U17845 ( .A(n17236), .B(n17103), .Z(N376) );
  NAND U17846 ( .A(n17105), .B(n17104), .Z(n17109) );
  NAND U17847 ( .A(n17107), .B(n17106), .Z(n17108) );
  AND U17848 ( .A(n17109), .B(n17108), .Z(n17377) );
  AND U17849 ( .A(x[244]), .B(y[1959]), .Z(n17110) );
  NAND U17850 ( .A(n17110), .B(n17342), .Z(n17114) );
  NANDN U17851 ( .A(n17112), .B(n17111), .Z(n17113) );
  NAND U17852 ( .A(n17114), .B(n17113), .Z(n17355) );
  AND U17853 ( .A(x[246]), .B(y[1954]), .Z(n17277) );
  XOR U17854 ( .A(n17278), .B(n17277), .Z(n17279) );
  NAND U17855 ( .A(x[226]), .B(y[1974]), .Z(n17280) );
  XNOR U17856 ( .A(n17279), .B(n17280), .Z(n17354) );
  AND U17857 ( .A(x[225]), .B(y[1975]), .Z(n17285) );
  XOR U17858 ( .A(n17286), .B(n17285), .Z(n17284) );
  ANDN U17859 ( .B(o[183]), .A(n17115), .Z(n17283) );
  XOR U17860 ( .A(n17284), .B(n17283), .Z(n17353) );
  XOR U17861 ( .A(n17354), .B(n17353), .Z(n17356) );
  XOR U17862 ( .A(n17355), .B(n17356), .Z(n17313) );
  NANDN U17863 ( .A(n17117), .B(n17116), .Z(n17121) );
  NANDN U17864 ( .A(n17119), .B(n17118), .Z(n17120) );
  NAND U17865 ( .A(n17121), .B(n17120), .Z(n17359) );
  AND U17866 ( .A(y[1960]), .B(x[240]), .Z(n17123) );
  NAND U17867 ( .A(y[1955]), .B(x[245]), .Z(n17122) );
  XNOR U17868 ( .A(n17123), .B(n17122), .Z(n17344) );
  AND U17869 ( .A(x[229]), .B(y[1971]), .Z(n17343) );
  XOR U17870 ( .A(n17344), .B(n17343), .Z(n17358) );
  AND U17871 ( .A(x[230]), .B(y[1970]), .Z(n17612) );
  AND U17872 ( .A(x[244]), .B(y[1956]), .Z(n17468) );
  XOR U17873 ( .A(n17612), .B(n17468), .Z(n17348) );
  AND U17874 ( .A(x[243]), .B(y[1957]), .Z(n17347) );
  XOR U17875 ( .A(n17348), .B(n17347), .Z(n17357) );
  XOR U17876 ( .A(n17358), .B(n17357), .Z(n17360) );
  XOR U17877 ( .A(n17359), .B(n17360), .Z(n17338) );
  NANDN U17878 ( .A(n17405), .B(n17124), .Z(n17128) );
  NANDN U17879 ( .A(n17126), .B(n17125), .Z(n17127) );
  NAND U17880 ( .A(n17128), .B(n17127), .Z(n17337) );
  NAND U17881 ( .A(n17130), .B(n17129), .Z(n17134) );
  NAND U17882 ( .A(n17132), .B(n17131), .Z(n17133) );
  NAND U17883 ( .A(n17134), .B(n17133), .Z(n17336) );
  XOR U17884 ( .A(n17337), .B(n17336), .Z(n17339) );
  XOR U17885 ( .A(n17338), .B(n17339), .Z(n17312) );
  XOR U17886 ( .A(n17313), .B(n17312), .Z(n17315) );
  NANDN U17887 ( .A(n17136), .B(n17135), .Z(n17140) );
  NANDN U17888 ( .A(n17138), .B(n17137), .Z(n17139) );
  AND U17889 ( .A(n17140), .B(n17139), .Z(n17307) );
  AND U17890 ( .A(x[227]), .B(y[1973]), .Z(n17296) );
  XOR U17891 ( .A(n17297), .B(n17296), .Z(n17298) );
  NAND U17892 ( .A(x[228]), .B(y[1972]), .Z(n17299) );
  XNOR U17893 ( .A(n17298), .B(n17299), .Z(n17306) );
  AND U17894 ( .A(y[1967]), .B(x[233]), .Z(n17142) );
  NAND U17895 ( .A(y[1966]), .B(x[234]), .Z(n17141) );
  XNOR U17896 ( .A(n17142), .B(n17141), .Z(n17271) );
  AND U17897 ( .A(y[1962]), .B(x[238]), .Z(n17144) );
  NAND U17898 ( .A(y[1968]), .B(x[232]), .Z(n17143) );
  XNOR U17899 ( .A(n17144), .B(n17143), .Z(n17273) );
  NAND U17900 ( .A(x[235]), .B(y[1965]), .Z(n17274) );
  XNOR U17901 ( .A(n17273), .B(n17274), .Z(n17270) );
  XOR U17902 ( .A(n17271), .B(n17270), .Z(n17308) );
  XOR U17903 ( .A(n17309), .B(n17308), .Z(n17314) );
  XNOR U17904 ( .A(n17315), .B(n17314), .Z(n17264) );
  NAND U17905 ( .A(n17146), .B(n17145), .Z(n17150) );
  NAND U17906 ( .A(n17148), .B(n17147), .Z(n17149) );
  AND U17907 ( .A(n17150), .B(n17149), .Z(n17263) );
  XOR U17908 ( .A(n17264), .B(n17263), .Z(n17265) );
  NAND U17909 ( .A(n17152), .B(n17151), .Z(n17156) );
  NAND U17910 ( .A(n17154), .B(n17153), .Z(n17155) );
  AND U17911 ( .A(n17156), .B(n17155), .Z(n17266) );
  XOR U17912 ( .A(n17265), .B(n17266), .Z(n17260) );
  NAND U17913 ( .A(n17158), .B(n17157), .Z(n17162) );
  NAND U17914 ( .A(n17160), .B(n17159), .Z(n17161) );
  AND U17915 ( .A(n17162), .B(n17161), .Z(n17321) );
  NANDN U17916 ( .A(n17164), .B(n17163), .Z(n17168) );
  NANDN U17917 ( .A(n17166), .B(n17165), .Z(n17167) );
  AND U17918 ( .A(n17168), .B(n17167), .Z(n17319) );
  NANDN U17919 ( .A(n17170), .B(n17169), .Z(n17174) );
  NAND U17920 ( .A(n17172), .B(n17171), .Z(n17173) );
  NAND U17921 ( .A(n17174), .B(n17173), .Z(n17351) );
  AND U17922 ( .A(x[224]), .B(y[1976]), .Z(n17302) );
  NAND U17923 ( .A(x[248]), .B(y[1952]), .Z(n17303) );
  XNOR U17924 ( .A(n17302), .B(n17303), .Z(n17305) );
  NAND U17925 ( .A(x[247]), .B(y[1953]), .Z(n17295) );
  XOR U17926 ( .A(n17305), .B(n17304), .Z(n17350) );
  AND U17927 ( .A(x[231]), .B(y[1969]), .Z(n17289) );
  NAND U17928 ( .A(x[242]), .B(y[1958]), .Z(n17290) );
  XNOR U17929 ( .A(n17289), .B(n17290), .Z(n17292) );
  AND U17930 ( .A(x[241]), .B(y[1959]), .Z(n17291) );
  XOR U17931 ( .A(n17292), .B(n17291), .Z(n17349) );
  XOR U17932 ( .A(n17350), .B(n17349), .Z(n17352) );
  XOR U17933 ( .A(n17351), .B(n17352), .Z(n17332) );
  NAND U17934 ( .A(n17176), .B(n17175), .Z(n17180) );
  NAND U17935 ( .A(n17178), .B(n17177), .Z(n17179) );
  NAND U17936 ( .A(n17180), .B(n17179), .Z(n17331) );
  NAND U17937 ( .A(n17182), .B(n17181), .Z(n17186) );
  NAND U17938 ( .A(n17184), .B(n17183), .Z(n17185) );
  NAND U17939 ( .A(n17186), .B(n17185), .Z(n17330) );
  XOR U17940 ( .A(n17331), .B(n17330), .Z(n17333) );
  XOR U17941 ( .A(n17332), .B(n17333), .Z(n17318) );
  NAND U17942 ( .A(n17188), .B(n17187), .Z(n17192) );
  NAND U17943 ( .A(n17190), .B(n17189), .Z(n17191) );
  AND U17944 ( .A(n17192), .B(n17191), .Z(n17364) );
  NAND U17945 ( .A(n17194), .B(n17193), .Z(n17198) );
  NAND U17946 ( .A(n17196), .B(n17195), .Z(n17197) );
  AND U17947 ( .A(n17198), .B(n17197), .Z(n17362) );
  NAND U17948 ( .A(n17200), .B(n17199), .Z(n17204) );
  NAND U17949 ( .A(n17202), .B(n17201), .Z(n17203) );
  AND U17950 ( .A(n17204), .B(n17203), .Z(n17361) );
  XOR U17951 ( .A(n17362), .B(n17361), .Z(n17363) );
  XOR U17952 ( .A(n17364), .B(n17363), .Z(n17324) );
  NAND U17953 ( .A(n17206), .B(n17205), .Z(n17210) );
  NAND U17954 ( .A(n17208), .B(n17207), .Z(n17209) );
  AND U17955 ( .A(n17210), .B(n17209), .Z(n17325) );
  XOR U17956 ( .A(n17324), .B(n17325), .Z(n17327) );
  XOR U17957 ( .A(n17326), .B(n17327), .Z(n17257) );
  IV U17958 ( .A(n17257), .Z(n17256) );
  NAND U17959 ( .A(n17212), .B(n17211), .Z(n17216) );
  NAND U17960 ( .A(n17214), .B(n17213), .Z(n17215) );
  AND U17961 ( .A(n17216), .B(n17215), .Z(n17258) );
  XOR U17962 ( .A(n17256), .B(n17258), .Z(n17217) );
  XOR U17963 ( .A(n17260), .B(n17217), .Z(n17374) );
  NAND U17964 ( .A(n17219), .B(n17218), .Z(n17223) );
  NAND U17965 ( .A(n17221), .B(n17220), .Z(n17222) );
  NAND U17966 ( .A(n17223), .B(n17222), .Z(n17253) );
  NAND U17967 ( .A(n17225), .B(n17224), .Z(n17229) );
  NAND U17968 ( .A(n17227), .B(n17226), .Z(n17228) );
  NAND U17969 ( .A(n17229), .B(n17228), .Z(n17251) );
  NAND U17970 ( .A(n17231), .B(n17230), .Z(n17235) );
  NAND U17971 ( .A(n17233), .B(n17232), .Z(n17234) );
  NAND U17972 ( .A(n17235), .B(n17234), .Z(n17250) );
  XOR U17973 ( .A(n17251), .B(n17250), .Z(n17252) );
  XOR U17974 ( .A(n17253), .B(n17252), .Z(n17375) );
  XOR U17975 ( .A(n17374), .B(n17375), .Z(n17376) );
  XNOR U17976 ( .A(n17377), .B(n17376), .Z(n17370) );
  OR U17977 ( .A(n17238), .B(n17236), .Z(n17242) );
  ANDN U17978 ( .B(n17238), .A(n17237), .Z(n17240) );
  OR U17979 ( .A(n17240), .B(n17239), .Z(n17241) );
  AND U17980 ( .A(n17242), .B(n17241), .Z(n17369) );
  NANDN U17981 ( .A(n17244), .B(n17243), .Z(n17248) );
  NANDN U17982 ( .A(n17246), .B(n17245), .Z(n17247) );
  AND U17983 ( .A(n17248), .B(n17247), .Z(n17368) );
  IV U17984 ( .A(n17368), .Z(n17367) );
  XOR U17985 ( .A(n17369), .B(n17367), .Z(n17249) );
  XNOR U17986 ( .A(n17370), .B(n17249), .Z(N377) );
  NAND U17987 ( .A(n17251), .B(n17250), .Z(n17255) );
  NAND U17988 ( .A(n17253), .B(n17252), .Z(n17254) );
  AND U17989 ( .A(n17255), .B(n17254), .Z(n17515) );
  NANDN U17990 ( .A(n17256), .B(n17258), .Z(n17262) );
  OR U17991 ( .A(n17258), .B(n17257), .Z(n17259) );
  NAND U17992 ( .A(n17260), .B(n17259), .Z(n17261) );
  NAND U17993 ( .A(n17262), .B(n17261), .Z(n17513) );
  NAND U17994 ( .A(n17264), .B(n17263), .Z(n17268) );
  NAND U17995 ( .A(n17266), .B(n17265), .Z(n17267) );
  NAND U17996 ( .A(n17268), .B(n17267), .Z(n17382) );
  NAND U17997 ( .A(x[238]), .B(y[1968]), .Z(n18200) );
  NANDN U17998 ( .A(n18200), .B(n17272), .Z(n17276) );
  NANDN U17999 ( .A(n17274), .B(n17273), .Z(n17275) );
  NAND U18000 ( .A(n17276), .B(n17275), .Z(n17445) );
  NAND U18001 ( .A(x[235]), .B(y[1966]), .Z(n17464) );
  NAND U18002 ( .A(x[236]), .B(y[1965]), .Z(n17463) );
  NAND U18003 ( .A(x[231]), .B(y[1970]), .Z(n17462) );
  XOR U18004 ( .A(n17463), .B(n17462), .Z(n17465) );
  XOR U18005 ( .A(n17464), .B(n17465), .Z(n17444) );
  AND U18006 ( .A(x[248]), .B(y[1953]), .Z(n17461) );
  XOR U18007 ( .A(o[185]), .B(n17461), .Z(n17432) );
  AND U18008 ( .A(x[225]), .B(y[1976]), .Z(n17431) );
  XOR U18009 ( .A(n17432), .B(n17431), .Z(n17434) );
  AND U18010 ( .A(x[237]), .B(y[1964]), .Z(n17433) );
  XOR U18011 ( .A(n17434), .B(n17433), .Z(n17443) );
  XOR U18012 ( .A(n17445), .B(n17446), .Z(n17422) );
  XOR U18013 ( .A(n17421), .B(n17422), .Z(n17424) );
  AND U18014 ( .A(n17278), .B(n17277), .Z(n17282) );
  NANDN U18015 ( .A(n17280), .B(n17279), .Z(n17281) );
  NANDN U18016 ( .A(n17282), .B(n17281), .Z(n17413) );
  AND U18017 ( .A(n17284), .B(n17283), .Z(n17288) );
  NAND U18018 ( .A(n17286), .B(n17285), .Z(n17287) );
  NANDN U18019 ( .A(n17288), .B(n17287), .Z(n17414) );
  XOR U18020 ( .A(n17413), .B(n17414), .Z(n17416) );
  NANDN U18021 ( .A(n17290), .B(n17289), .Z(n17294) );
  NAND U18022 ( .A(n17292), .B(n17291), .Z(n17293) );
  NAND U18023 ( .A(n17294), .B(n17293), .Z(n17411) );
  NAND U18024 ( .A(x[232]), .B(y[1969]), .Z(n17407) );
  XOR U18025 ( .A(n17405), .B(n17406), .Z(n17408) );
  XOR U18026 ( .A(n17407), .B(n17408), .Z(n17410) );
  NANDN U18027 ( .A(n17295), .B(o[184]), .Z(n17401) );
  NAND U18028 ( .A(x[249]), .B(y[1952]), .Z(n17400) );
  NAND U18029 ( .A(x[224]), .B(y[1977]), .Z(n17399) );
  XNOR U18030 ( .A(n17400), .B(n17399), .Z(n17402) );
  XOR U18031 ( .A(n17401), .B(n17402), .Z(n17409) );
  XNOR U18032 ( .A(n17410), .B(n17409), .Z(n17412) );
  XOR U18033 ( .A(n17411), .B(n17412), .Z(n17415) );
  XOR U18034 ( .A(n17416), .B(n17415), .Z(n17423) );
  XOR U18035 ( .A(n17424), .B(n17423), .Z(n17496) );
  AND U18036 ( .A(n17297), .B(n17296), .Z(n17301) );
  NANDN U18037 ( .A(n17299), .B(n17298), .Z(n17300) );
  NANDN U18038 ( .A(n17301), .B(n17300), .Z(n17481) );
  AND U18039 ( .A(x[238]), .B(y[1963]), .Z(n17438) );
  AND U18040 ( .A(x[226]), .B(y[1975]), .Z(n17437) );
  XOR U18041 ( .A(n17438), .B(n17437), .Z(n17440) );
  AND U18042 ( .A(x[227]), .B(y[1974]), .Z(n17439) );
  XOR U18043 ( .A(n17440), .B(n17439), .Z(n17480) );
  XOR U18044 ( .A(n17479), .B(n17480), .Z(n17482) );
  XOR U18045 ( .A(n17481), .B(n17482), .Z(n17494) );
  NANDN U18046 ( .A(n17307), .B(n17306), .Z(n17311) );
  NAND U18047 ( .A(n17309), .B(n17308), .Z(n17310) );
  AND U18048 ( .A(n17311), .B(n17310), .Z(n17493) );
  NAND U18049 ( .A(n17313), .B(n17312), .Z(n17317) );
  NAND U18050 ( .A(n17315), .B(n17314), .Z(n17316) );
  AND U18051 ( .A(n17317), .B(n17316), .Z(n17499) );
  XOR U18052 ( .A(n17500), .B(n17499), .Z(n17502) );
  NANDN U18053 ( .A(n17319), .B(n17318), .Z(n17323) );
  NANDN U18054 ( .A(n17321), .B(n17320), .Z(n17322) );
  AND U18055 ( .A(n17323), .B(n17322), .Z(n17501) );
  XOR U18056 ( .A(n17502), .B(n17501), .Z(n17381) );
  XOR U18057 ( .A(n17382), .B(n17381), .Z(n17384) );
  NAND U18058 ( .A(n17325), .B(n17324), .Z(n17329) );
  NAND U18059 ( .A(n17327), .B(n17326), .Z(n17328) );
  NAND U18060 ( .A(n17329), .B(n17328), .Z(n17389) );
  NAND U18061 ( .A(n17331), .B(n17330), .Z(n17335) );
  NAND U18062 ( .A(n17333), .B(n17332), .Z(n17334) );
  NAND U18063 ( .A(n17335), .B(n17334), .Z(n17394) );
  NAND U18064 ( .A(n17337), .B(n17336), .Z(n17341) );
  NAND U18065 ( .A(n17339), .B(n17338), .Z(n17340) );
  NAND U18066 ( .A(n17341), .B(n17340), .Z(n17393) );
  XOR U18067 ( .A(n17394), .B(n17393), .Z(n17396) );
  AND U18068 ( .A(x[245]), .B(y[1960]), .Z(n18242) );
  NAND U18069 ( .A(x[246]), .B(y[1955]), .Z(n17457) );
  NAND U18070 ( .A(x[229]), .B(y[1972]), .Z(n17456) );
  NAND U18071 ( .A(x[241]), .B(y[1960]), .Z(n17455) );
  XOR U18072 ( .A(n17456), .B(n17455), .Z(n17458) );
  XOR U18073 ( .A(n17457), .B(n17458), .Z(n17484) );
  AND U18074 ( .A(y[1957]), .B(x[244]), .Z(n17346) );
  NAND U18075 ( .A(y[1956]), .B(x[245]), .Z(n17345) );
  XNOR U18076 ( .A(n17346), .B(n17345), .Z(n17470) );
  AND U18077 ( .A(x[243]), .B(y[1958]), .Z(n17469) );
  XOR U18078 ( .A(n17470), .B(n17469), .Z(n17483) );
  XNOR U18079 ( .A(n17484), .B(n17483), .Z(n17486) );
  XOR U18080 ( .A(n17485), .B(n17486), .Z(n17418) );
  NAND U18081 ( .A(x[239]), .B(y[1962]), .Z(n17475) );
  NAND U18082 ( .A(x[242]), .B(y[1959]), .Z(n17474) );
  NAND U18083 ( .A(x[230]), .B(y[1971]), .Z(n17473) );
  XOR U18084 ( .A(n17474), .B(n17473), .Z(n17476) );
  XOR U18085 ( .A(n17475), .B(n17476), .Z(n17488) );
  NAND U18086 ( .A(x[247]), .B(y[1954]), .Z(n17451) );
  NAND U18087 ( .A(x[228]), .B(y[1973]), .Z(n17450) );
  NAND U18088 ( .A(x[240]), .B(y[1961]), .Z(n17449) );
  XOR U18089 ( .A(n17450), .B(n17449), .Z(n17452) );
  XOR U18090 ( .A(n17451), .B(n17452), .Z(n17487) );
  XNOR U18091 ( .A(n17488), .B(n17487), .Z(n17490) );
  XOR U18092 ( .A(n17489), .B(n17490), .Z(n17417) );
  XNOR U18093 ( .A(n17418), .B(n17417), .Z(n17420) );
  XOR U18094 ( .A(n17420), .B(n17419), .Z(n17427) );
  XNOR U18095 ( .A(n17425), .B(n17426), .Z(n17428) );
  XOR U18096 ( .A(n17427), .B(n17428), .Z(n17395) );
  XNOR U18097 ( .A(n17396), .B(n17395), .Z(n17388) );
  NAND U18098 ( .A(n17362), .B(n17361), .Z(n17366) );
  NAND U18099 ( .A(n17364), .B(n17363), .Z(n17365) );
  NAND U18100 ( .A(n17366), .B(n17365), .Z(n17387) );
  XOR U18101 ( .A(n17388), .B(n17387), .Z(n17390) );
  XOR U18102 ( .A(n17389), .B(n17390), .Z(n17383) );
  XOR U18103 ( .A(n17384), .B(n17383), .Z(n17512) );
  XOR U18104 ( .A(n17513), .B(n17512), .Z(n17514) );
  XNOR U18105 ( .A(n17515), .B(n17514), .Z(n17508) );
  OR U18106 ( .A(n17369), .B(n17367), .Z(n17373) );
  ANDN U18107 ( .B(n17369), .A(n17368), .Z(n17371) );
  OR U18108 ( .A(n17371), .B(n17370), .Z(n17372) );
  AND U18109 ( .A(n17373), .B(n17372), .Z(n17506) );
  NAND U18110 ( .A(n17375), .B(n17374), .Z(n17379) );
  NAND U18111 ( .A(n17377), .B(n17376), .Z(n17378) );
  AND U18112 ( .A(n17379), .B(n17378), .Z(n17507) );
  IV U18113 ( .A(n17507), .Z(n17505) );
  XOR U18114 ( .A(n17506), .B(n17505), .Z(n17380) );
  XNOR U18115 ( .A(n17508), .B(n17380), .Z(N378) );
  NAND U18116 ( .A(n17382), .B(n17381), .Z(n17386) );
  NAND U18117 ( .A(n17384), .B(n17383), .Z(n17385) );
  AND U18118 ( .A(n17386), .B(n17385), .Z(n17641) );
  NAND U18119 ( .A(n17388), .B(n17387), .Z(n17392) );
  NAND U18120 ( .A(n17390), .B(n17389), .Z(n17391) );
  AND U18121 ( .A(n17392), .B(n17391), .Z(n17642) );
  XOR U18122 ( .A(n17641), .B(n17642), .Z(n17644) );
  NAND U18123 ( .A(n17394), .B(n17393), .Z(n17398) );
  NAND U18124 ( .A(n17396), .B(n17395), .Z(n17397) );
  NAND U18125 ( .A(n17398), .B(n17397), .Z(n17634) );
  AND U18126 ( .A(x[226]), .B(y[1976]), .Z(n17533) );
  XOR U18127 ( .A(n17534), .B(n17533), .Z(n17536) );
  AND U18128 ( .A(x[248]), .B(y[1954]), .Z(n17535) );
  XOR U18129 ( .A(n17536), .B(n17535), .Z(n17564) );
  NAND U18130 ( .A(n17400), .B(n17399), .Z(n17404) );
  NANDN U18131 ( .A(n17402), .B(n17401), .Z(n17403) );
  AND U18132 ( .A(n17404), .B(n17403), .Z(n17563) );
  XOR U18133 ( .A(n17564), .B(n17563), .Z(n17566) );
  XOR U18134 ( .A(n17566), .B(n17565), .Z(n17625) );
  XNOR U18135 ( .A(n17625), .B(n17624), .Z(n17627) );
  XOR U18136 ( .A(n17627), .B(n17626), .Z(n17630) );
  XNOR U18137 ( .A(n17629), .B(n17628), .Z(n17631) );
  XOR U18138 ( .A(n17630), .B(n17631), .Z(n17632) );
  AND U18139 ( .A(x[236]), .B(y[1966]), .Z(n17696) );
  AND U18140 ( .A(x[229]), .B(y[1973]), .Z(n17577) );
  XOR U18141 ( .A(n17696), .B(n17577), .Z(n17579) );
  AND U18142 ( .A(x[234]), .B(y[1968]), .Z(n17578) );
  XOR U18143 ( .A(n17579), .B(n17578), .Z(n17603) );
  AND U18144 ( .A(x[231]), .B(y[1971]), .Z(n17601) );
  AND U18145 ( .A(y[1972]), .B(x[230]), .Z(n17430) );
  NAND U18146 ( .A(y[1970]), .B(x[232]), .Z(n17429) );
  XNOR U18147 ( .A(n17430), .B(n17429), .Z(n17614) );
  AND U18148 ( .A(x[233]), .B(y[1969]), .Z(n17613) );
  XOR U18149 ( .A(n17614), .B(n17613), .Z(n17600) );
  XOR U18150 ( .A(n17601), .B(n17600), .Z(n17602) );
  XOR U18151 ( .A(n17603), .B(n17602), .Z(n17555) );
  NAND U18152 ( .A(n17432), .B(n17431), .Z(n17436) );
  NAND U18153 ( .A(n17434), .B(n17433), .Z(n17435) );
  NAND U18154 ( .A(n17436), .B(n17435), .Z(n17553) );
  NAND U18155 ( .A(n17438), .B(n17437), .Z(n17442) );
  NAND U18156 ( .A(n17440), .B(n17439), .Z(n17441) );
  NAND U18157 ( .A(n17442), .B(n17441), .Z(n17554) );
  XNOR U18158 ( .A(n17553), .B(n17554), .Z(n17556) );
  XOR U18159 ( .A(n17555), .B(n17556), .Z(n17588) );
  NANDN U18160 ( .A(n17444), .B(n17443), .Z(n17448) );
  NAND U18161 ( .A(n17446), .B(n17445), .Z(n17447) );
  AND U18162 ( .A(n17448), .B(n17447), .Z(n17589) );
  XOR U18163 ( .A(n17588), .B(n17589), .Z(n17590) );
  NAND U18164 ( .A(n17450), .B(n17449), .Z(n17454) );
  NAND U18165 ( .A(n17452), .B(n17451), .Z(n17453) );
  AND U18166 ( .A(n17454), .B(n17453), .Z(n17526) );
  NAND U18167 ( .A(n17456), .B(n17455), .Z(n17460) );
  NAND U18168 ( .A(n17458), .B(n17457), .Z(n17459) );
  AND U18169 ( .A(n17460), .B(n17459), .Z(n17525) );
  XOR U18170 ( .A(n17526), .B(n17525), .Z(n17528) );
  AND U18171 ( .A(x[238]), .B(y[1964]), .Z(n17608) );
  XOR U18172 ( .A(n17609), .B(n17608), .Z(n17611) );
  AND U18173 ( .A(x[225]), .B(y[1977]), .Z(n17610) );
  XOR U18174 ( .A(n17611), .B(n17610), .Z(n17570) );
  AND U18175 ( .A(x[249]), .B(y[1953]), .Z(n17617) );
  XOR U18176 ( .A(o[186]), .B(n17617), .Z(n17583) );
  AND U18177 ( .A(x[250]), .B(y[1952]), .Z(n17582) );
  XOR U18178 ( .A(n17583), .B(n17582), .Z(n17585) );
  AND U18179 ( .A(x[224]), .B(y[1978]), .Z(n17584) );
  XOR U18180 ( .A(n17585), .B(n17584), .Z(n17569) );
  XOR U18181 ( .A(n17570), .B(n17569), .Z(n17572) );
  NAND U18182 ( .A(n17463), .B(n17462), .Z(n17467) );
  NAND U18183 ( .A(n17465), .B(n17464), .Z(n17466) );
  AND U18184 ( .A(n17467), .B(n17466), .Z(n17571) );
  XOR U18185 ( .A(n17572), .B(n17571), .Z(n17527) );
  XOR U18186 ( .A(n17528), .B(n17527), .Z(n17560) );
  NAND U18187 ( .A(x[245]), .B(y[1957]), .Z(n17604) );
  NANDN U18188 ( .A(n17604), .B(n17468), .Z(n17472) );
  NAND U18189 ( .A(n17470), .B(n17469), .Z(n17471) );
  NAND U18190 ( .A(n17472), .B(n17471), .Z(n17551) );
  AND U18191 ( .A(x[244]), .B(y[1958]), .Z(n17606) );
  XOR U18192 ( .A(n17607), .B(n17606), .Z(n17550) );
  AND U18193 ( .A(x[247]), .B(y[1955]), .Z(n17539) );
  XOR U18194 ( .A(n17540), .B(n17539), .Z(n17542) );
  AND U18195 ( .A(x[246]), .B(y[1956]), .Z(n17541) );
  XOR U18196 ( .A(n17542), .B(n17541), .Z(n17549) );
  XOR U18197 ( .A(n17550), .B(n17549), .Z(n17552) );
  XOR U18198 ( .A(n17551), .B(n17552), .Z(n17558) );
  AND U18199 ( .A(x[228]), .B(y[1974]), .Z(n17543) );
  XOR U18200 ( .A(n17544), .B(n17543), .Z(n17546) );
  XOR U18201 ( .A(n17546), .B(n17545), .Z(n17530) );
  AND U18202 ( .A(x[243]), .B(y[1959]), .Z(n17619) );
  AND U18203 ( .A(x[227]), .B(y[1975]), .Z(n17618) );
  XOR U18204 ( .A(n17619), .B(n17618), .Z(n17621) );
  AND U18205 ( .A(x[235]), .B(y[1967]), .Z(n17620) );
  XOR U18206 ( .A(n17621), .B(n17620), .Z(n17529) );
  XOR U18207 ( .A(n17530), .B(n17529), .Z(n17532) );
  NAND U18208 ( .A(n17474), .B(n17473), .Z(n17478) );
  NAND U18209 ( .A(n17476), .B(n17475), .Z(n17477) );
  AND U18210 ( .A(n17478), .B(n17477), .Z(n17531) );
  XOR U18211 ( .A(n17532), .B(n17531), .Z(n17557) );
  XOR U18212 ( .A(n17558), .B(n17557), .Z(n17559) );
  XOR U18213 ( .A(n17560), .B(n17559), .Z(n17591) );
  XOR U18214 ( .A(n17590), .B(n17591), .Z(n17592) );
  OR U18215 ( .A(n17488), .B(n17487), .Z(n17492) );
  NANDN U18216 ( .A(n17490), .B(n17489), .Z(n17491) );
  NAND U18217 ( .A(n17492), .B(n17491), .Z(n17597) );
  XOR U18218 ( .A(n17596), .B(n17597), .Z(n17599) );
  XOR U18219 ( .A(n17598), .B(n17599), .Z(n17593) );
  XOR U18220 ( .A(n17592), .B(n17593), .Z(n17595) );
  XOR U18221 ( .A(n17594), .B(n17595), .Z(n17633) );
  XOR U18222 ( .A(n17632), .B(n17633), .Z(n17635) );
  XOR U18223 ( .A(n17634), .B(n17635), .Z(n17522) );
  NANDN U18224 ( .A(n17494), .B(n17493), .Z(n17498) );
  NANDN U18225 ( .A(n17496), .B(n17495), .Z(n17497) );
  AND U18226 ( .A(n17498), .B(n17497), .Z(n17520) );
  NAND U18227 ( .A(n17500), .B(n17499), .Z(n17504) );
  NAND U18228 ( .A(n17502), .B(n17501), .Z(n17503) );
  AND U18229 ( .A(n17504), .B(n17503), .Z(n17519) );
  XOR U18230 ( .A(n17520), .B(n17519), .Z(n17521) );
  XOR U18231 ( .A(n17522), .B(n17521), .Z(n17643) );
  XNOR U18232 ( .A(n17644), .B(n17643), .Z(n17640) );
  NANDN U18233 ( .A(n17505), .B(n17506), .Z(n17511) );
  NOR U18234 ( .A(n17507), .B(n17506), .Z(n17509) );
  OR U18235 ( .A(n17509), .B(n17508), .Z(n17510) );
  AND U18236 ( .A(n17511), .B(n17510), .Z(n17638) );
  NAND U18237 ( .A(n17513), .B(n17512), .Z(n17517) );
  NAND U18238 ( .A(n17515), .B(n17514), .Z(n17516) );
  AND U18239 ( .A(n17517), .B(n17516), .Z(n17639) );
  XOR U18240 ( .A(n17638), .B(n17639), .Z(n17518) );
  XNOR U18241 ( .A(n17640), .B(n17518), .Z(N379) );
  NAND U18242 ( .A(n17520), .B(n17519), .Z(n17524) );
  NAND U18243 ( .A(n17522), .B(n17521), .Z(n17523) );
  AND U18244 ( .A(n17524), .B(n17523), .Z(n17789) );
  AND U18245 ( .A(n17534), .B(n17533), .Z(n17538) );
  NAND U18246 ( .A(n17536), .B(n17535), .Z(n17537) );
  NANDN U18247 ( .A(n17538), .B(n17537), .Z(n17671) );
  XOR U18248 ( .A(n17671), .B(n17670), .Z(n17672) );
  AND U18249 ( .A(n17544), .B(n17543), .Z(n17548) );
  NAND U18250 ( .A(n17546), .B(n17545), .Z(n17547) );
  NANDN U18251 ( .A(n17548), .B(n17547), .Z(n17684) );
  AND U18252 ( .A(x[224]), .B(y[1979]), .Z(n17745) );
  AND U18253 ( .A(x[251]), .B(y[1952]), .Z(n17744) );
  XOR U18254 ( .A(n17745), .B(n17744), .Z(n17747) );
  AND U18255 ( .A(x[250]), .B(y[1953]), .Z(n17737) );
  XOR U18256 ( .A(n17737), .B(o[187]), .Z(n17746) );
  XOR U18257 ( .A(n17747), .B(n17746), .Z(n17683) );
  AND U18258 ( .A(x[233]), .B(y[1970]), .Z(n17734) );
  AND U18259 ( .A(x[245]), .B(y[1958]), .Z(n17733) );
  XOR U18260 ( .A(n17734), .B(n17733), .Z(n17736) );
  AND U18261 ( .A(x[242]), .B(y[1961]), .Z(n17735) );
  XOR U18262 ( .A(n17736), .B(n17735), .Z(n17682) );
  XOR U18263 ( .A(n17683), .B(n17682), .Z(n17685) );
  XNOR U18264 ( .A(n17684), .B(n17685), .Z(n17673) );
  XOR U18265 ( .A(n17755), .B(n17756), .Z(n17758) );
  XOR U18266 ( .A(n17757), .B(n17758), .Z(n17776) );
  XOR U18267 ( .A(n17774), .B(n17773), .Z(n17775) );
  OR U18268 ( .A(n17558), .B(n17557), .Z(n17562) );
  NANDN U18269 ( .A(n17560), .B(n17559), .Z(n17561) );
  AND U18270 ( .A(n17562), .B(n17561), .Z(n17761) );
  NAND U18271 ( .A(n17564), .B(n17563), .Z(n17568) );
  NAND U18272 ( .A(n17566), .B(n17565), .Z(n17567) );
  NAND U18273 ( .A(n17568), .B(n17567), .Z(n17751) );
  NAND U18274 ( .A(n17570), .B(n17569), .Z(n17574) );
  NAND U18275 ( .A(n17572), .B(n17571), .Z(n17573) );
  NAND U18276 ( .A(n17574), .B(n17573), .Z(n17749) );
  AND U18277 ( .A(x[243]), .B(y[1960]), .Z(n17730) );
  AND U18278 ( .A(x[249]), .B(y[1954]), .Z(n17729) );
  XOR U18279 ( .A(n17730), .B(n17729), .Z(n17732) );
  AND U18280 ( .A(x[230]), .B(y[1973]), .Z(n17731) );
  XOR U18281 ( .A(n17732), .B(n17731), .Z(n17722) );
  AND U18282 ( .A(x[239]), .B(y[1964]), .Z(n17702) );
  AND U18283 ( .A(x[226]), .B(y[1977]), .Z(n17701) );
  XOR U18284 ( .A(n17702), .B(n17701), .Z(n17704) );
  AND U18285 ( .A(x[227]), .B(y[1976]), .Z(n17703) );
  XOR U18286 ( .A(n17704), .B(n17703), .Z(n17721) );
  XOR U18287 ( .A(n17722), .B(n17721), .Z(n17723) );
  NAND U18288 ( .A(x[240]), .B(y[1963]), .Z(n17689) );
  XOR U18289 ( .A(n17689), .B(n17688), .Z(n17691) );
  XOR U18290 ( .A(n17690), .B(n17691), .Z(n17698) );
  AND U18291 ( .A(y[1966]), .B(x[237]), .Z(n17576) );
  AND U18292 ( .A(y[1967]), .B(x[236]), .Z(n17575) );
  XOR U18293 ( .A(n17576), .B(n17575), .Z(n17697) );
  XOR U18294 ( .A(n17698), .B(n17697), .Z(n17724) );
  AND U18295 ( .A(n17696), .B(n17577), .Z(n17581) );
  NAND U18296 ( .A(n17579), .B(n17578), .Z(n17580) );
  NANDN U18297 ( .A(n17581), .B(n17580), .Z(n17665) );
  NAND U18298 ( .A(n17583), .B(n17582), .Z(n17587) );
  NAND U18299 ( .A(n17585), .B(n17584), .Z(n17586) );
  NAND U18300 ( .A(n17587), .B(n17586), .Z(n17664) );
  XOR U18301 ( .A(n17665), .B(n17664), .Z(n17666) );
  XOR U18302 ( .A(n17667), .B(n17666), .Z(n17750) );
  XNOR U18303 ( .A(n17749), .B(n17750), .Z(n17752) );
  XNOR U18304 ( .A(n17761), .B(n17762), .Z(n17764) );
  XOR U18305 ( .A(n17764), .B(n17763), .Z(n17652) );
  XOR U18306 ( .A(n17655), .B(n17654), .Z(n17651) );
  XOR U18307 ( .A(n17710), .B(n17709), .Z(n17711) );
  AND U18308 ( .A(x[232]), .B(y[1972]), .Z(n17739) );
  NAND U18309 ( .A(n17612), .B(n17739), .Z(n17616) );
  NAND U18310 ( .A(n17614), .B(n17613), .Z(n17615) );
  NAND U18311 ( .A(n17616), .B(n17615), .Z(n17678) );
  AND U18312 ( .A(x[238]), .B(y[1965]), .Z(n17706) );
  AND U18313 ( .A(x[225]), .B(y[1978]), .Z(n17705) );
  XOR U18314 ( .A(n17706), .B(n17705), .Z(n17707) );
  XOR U18315 ( .A(n17707), .B(n17708), .Z(n17677) );
  AND U18316 ( .A(x[241]), .B(y[1962]), .Z(n17741) );
  AND U18317 ( .A(x[228]), .B(y[1975]), .Z(n17740) );
  XOR U18318 ( .A(n17741), .B(n17740), .Z(n17743) );
  AND U18319 ( .A(x[229]), .B(y[1974]), .Z(n17742) );
  XOR U18320 ( .A(n17743), .B(n17742), .Z(n17676) );
  XOR U18321 ( .A(n17677), .B(n17676), .Z(n17679) );
  XNOR U18322 ( .A(n17678), .B(n17679), .Z(n17712) );
  AND U18323 ( .A(y[1955]), .B(x[248]), .Z(n17623) );
  NAND U18324 ( .A(y[1959]), .B(x[244]), .Z(n17622) );
  XNOR U18325 ( .A(n17623), .B(n17622), .Z(n17728) );
  AND U18326 ( .A(x[231]), .B(y[1972]), .Z(n17727) );
  XOR U18327 ( .A(n17728), .B(n17727), .Z(n17716) );
  AND U18328 ( .A(x[232]), .B(y[1971]), .Z(n17693) );
  AND U18329 ( .A(x[247]), .B(y[1956]), .Z(n17692) );
  XOR U18330 ( .A(n17693), .B(n17692), .Z(n17695) );
  AND U18331 ( .A(x[246]), .B(y[1957]), .Z(n17694) );
  XOR U18332 ( .A(n17695), .B(n17694), .Z(n17715) );
  XOR U18333 ( .A(n17716), .B(n17715), .Z(n17718) );
  XNOR U18334 ( .A(n17717), .B(n17718), .Z(n17768) );
  XOR U18335 ( .A(n17769), .B(n17770), .Z(n17659) );
  XOR U18336 ( .A(n17659), .B(n17658), .Z(n17661) );
  XOR U18337 ( .A(n17660), .B(n17661), .Z(n17649) );
  XOR U18338 ( .A(n17649), .B(n17648), .Z(n17650) );
  XOR U18339 ( .A(n17651), .B(n17650), .Z(n17787) );
  NAND U18340 ( .A(n17633), .B(n17632), .Z(n17637) );
  NAND U18341 ( .A(n17635), .B(n17634), .Z(n17636) );
  AND U18342 ( .A(n17637), .B(n17636), .Z(n17786) );
  XNOR U18343 ( .A(n17789), .B(n17788), .Z(n17782) );
  NAND U18344 ( .A(n17642), .B(n17641), .Z(n17646) );
  NAND U18345 ( .A(n17644), .B(n17643), .Z(n17645) );
  AND U18346 ( .A(n17646), .B(n17645), .Z(n17781) );
  IV U18347 ( .A(n17781), .Z(n17779) );
  XOR U18348 ( .A(n17780), .B(n17779), .Z(n17647) );
  XNOR U18349 ( .A(n17782), .B(n17647), .Z(N380) );
  NANDN U18350 ( .A(n17653), .B(n17652), .Z(n17657) );
  NAND U18351 ( .A(n17655), .B(n17654), .Z(n17656) );
  NAND U18352 ( .A(n17657), .B(n17656), .Z(n17794) );
  XOR U18353 ( .A(n17793), .B(n17794), .Z(n17796) );
  NAND U18354 ( .A(n17659), .B(n17658), .Z(n17663) );
  NAND U18355 ( .A(n17661), .B(n17660), .Z(n17662) );
  NAND U18356 ( .A(n17663), .B(n17662), .Z(n17800) );
  NAND U18357 ( .A(n17665), .B(n17664), .Z(n17669) );
  NAND U18358 ( .A(n17667), .B(n17666), .Z(n17668) );
  NAND U18359 ( .A(n17669), .B(n17668), .Z(n17824) );
  NAND U18360 ( .A(n17671), .B(n17670), .Z(n17675) );
  NANDN U18361 ( .A(n17673), .B(n17672), .Z(n17674) );
  NAND U18362 ( .A(n17675), .B(n17674), .Z(n17903) );
  NAND U18363 ( .A(n17677), .B(n17676), .Z(n17681) );
  NAND U18364 ( .A(n17679), .B(n17678), .Z(n17680) );
  NAND U18365 ( .A(n17681), .B(n17680), .Z(n17902) );
  NAND U18366 ( .A(n17683), .B(n17682), .Z(n17687) );
  NAND U18367 ( .A(n17685), .B(n17684), .Z(n17686) );
  NAND U18368 ( .A(n17687), .B(n17686), .Z(n17901) );
  XOR U18369 ( .A(n17902), .B(n17901), .Z(n17904) );
  XOR U18370 ( .A(n17903), .B(n17904), .Z(n17825) );
  XOR U18371 ( .A(n17824), .B(n17825), .Z(n17827) );
  AND U18372 ( .A(x[231]), .B(y[1973]), .Z(n17860) );
  AND U18373 ( .A(x[236]), .B(y[1968]), .Z(n17859) );
  XOR U18374 ( .A(n17860), .B(n17859), .Z(n17862) );
  AND U18375 ( .A(x[235]), .B(y[1969]), .Z(n17861) );
  XOR U18376 ( .A(n17862), .B(n17861), .Z(n17882) );
  NAND U18377 ( .A(x[251]), .B(y[1953]), .Z(n17870) );
  XNOR U18378 ( .A(o[188]), .B(n17870), .Z(n17876) );
  AND U18379 ( .A(x[250]), .B(y[1954]), .Z(n17875) );
  XOR U18380 ( .A(n17876), .B(n17875), .Z(n17878) );
  AND U18381 ( .A(x[239]), .B(y[1965]), .Z(n17877) );
  XNOR U18382 ( .A(n17878), .B(n17877), .Z(n17881) );
  XNOR U18383 ( .A(n17882), .B(n17881), .Z(n17884) );
  XOR U18384 ( .A(n17883), .B(n17884), .Z(n17920) );
  AND U18385 ( .A(x[241]), .B(y[1963]), .Z(n17835) );
  AND U18386 ( .A(x[246]), .B(y[1958]), .Z(n17834) );
  XOR U18387 ( .A(n17835), .B(n17834), .Z(n17837) );
  AND U18388 ( .A(x[228]), .B(y[1976]), .Z(n17836) );
  XOR U18389 ( .A(n17837), .B(n17836), .Z(n17886) );
  AND U18390 ( .A(x[230]), .B(y[1974]), .Z(n18005) );
  AND U18391 ( .A(x[243]), .B(y[1961]), .Z(n17863) );
  XOR U18392 ( .A(n18005), .B(n17863), .Z(n17865) );
  XOR U18393 ( .A(n17865), .B(n17864), .Z(n17885) );
  XOR U18394 ( .A(n17886), .B(n17885), .Z(n17888) );
  XOR U18395 ( .A(n17887), .B(n17888), .Z(n17919) );
  NAND U18396 ( .A(n17872), .B(n17696), .Z(n17700) );
  NANDN U18397 ( .A(n17698), .B(n17697), .Z(n17699) );
  NAND U18398 ( .A(n17700), .B(n17699), .Z(n17832) );
  XOR U18399 ( .A(n17830), .B(n17831), .Z(n17833) );
  XOR U18400 ( .A(n17832), .B(n17833), .Z(n17921) );
  XOR U18401 ( .A(n17922), .B(n17921), .Z(n17826) );
  XOR U18402 ( .A(n17827), .B(n17826), .Z(n17821) );
  NAND U18403 ( .A(n17710), .B(n17709), .Z(n17714) );
  NANDN U18404 ( .A(n17712), .B(n17711), .Z(n17713) );
  NAND U18405 ( .A(n17714), .B(n17713), .Z(n17891) );
  NAND U18406 ( .A(n17716), .B(n17715), .Z(n17720) );
  NAND U18407 ( .A(n17718), .B(n17717), .Z(n17719) );
  NAND U18408 ( .A(n17720), .B(n17719), .Z(n17890) );
  NAND U18409 ( .A(n17722), .B(n17721), .Z(n17726) );
  NANDN U18410 ( .A(n17724), .B(n17723), .Z(n17725) );
  NAND U18411 ( .A(n17726), .B(n17725), .Z(n17889) );
  XOR U18412 ( .A(n17890), .B(n17889), .Z(n17892) );
  XOR U18413 ( .A(n17891), .B(n17892), .Z(n17819) );
  AND U18414 ( .A(x[248]), .B(y[1959]), .Z(n18157) );
  AND U18415 ( .A(x[249]), .B(y[1955]), .Z(n17857) );
  XOR U18416 ( .A(n17858), .B(n17857), .Z(n17856) );
  AND U18417 ( .A(x[225]), .B(y[1979]), .Z(n17855) );
  XOR U18418 ( .A(n17856), .B(n17855), .Z(n17916) );
  AND U18419 ( .A(x[240]), .B(y[1964]), .Z(n17852) );
  AND U18420 ( .A(x[248]), .B(y[1956]), .Z(n17851) );
  XOR U18421 ( .A(n17852), .B(n17851), .Z(n17854) );
  AND U18422 ( .A(x[226]), .B(y[1978]), .Z(n17853) );
  XOR U18423 ( .A(n17854), .B(n17853), .Z(n17915) );
  XOR U18424 ( .A(n17916), .B(n17915), .Z(n17918) );
  XOR U18425 ( .A(n17917), .B(n17918), .Z(n17898) );
  AND U18426 ( .A(x[227]), .B(y[1977]), .Z(n17871) );
  XOR U18427 ( .A(n17872), .B(n17871), .Z(n17874) );
  AND U18428 ( .A(x[247]), .B(y[1957]), .Z(n17873) );
  XOR U18429 ( .A(n17874), .B(n17873), .Z(n17912) );
  AND U18430 ( .A(x[229]), .B(y[1975]), .Z(n17867) );
  AND U18431 ( .A(x[245]), .B(y[1959]), .Z(n17866) );
  XOR U18432 ( .A(n17867), .B(n17866), .Z(n17869) );
  AND U18433 ( .A(x[244]), .B(y[1960]), .Z(n17868) );
  XOR U18434 ( .A(n17869), .B(n17868), .Z(n17911) );
  XOR U18435 ( .A(n17912), .B(n17911), .Z(n17914) );
  XOR U18436 ( .A(n17913), .B(n17914), .Z(n17896) );
  IV U18437 ( .A(n17896), .Z(n17748) );
  AND U18438 ( .A(x[224]), .B(y[1980]), .Z(n17839) );
  AND U18439 ( .A(x[252]), .B(y[1952]), .Z(n17838) );
  XOR U18440 ( .A(n17839), .B(n17838), .Z(n17841) );
  AND U18441 ( .A(n17737), .B(o[187]), .Z(n17840) );
  XOR U18442 ( .A(n17841), .B(n17840), .Z(n17848) );
  NAND U18443 ( .A(y[1970]), .B(x[234]), .Z(n17738) );
  XNOR U18444 ( .A(n17739), .B(n17738), .Z(n17844) );
  AND U18445 ( .A(x[233]), .B(y[1971]), .Z(n17843) );
  XOR U18446 ( .A(n17844), .B(n17843), .Z(n17847) );
  XOR U18447 ( .A(n17848), .B(n17847), .Z(n17850) );
  XOR U18448 ( .A(n17849), .B(n17850), .Z(n17910) );
  XOR U18449 ( .A(n17907), .B(n17908), .Z(n17909) );
  XNOR U18450 ( .A(n17910), .B(n17909), .Z(n17895) );
  XOR U18451 ( .A(n17748), .B(n17895), .Z(n17897) );
  NAND U18452 ( .A(n17750), .B(n17749), .Z(n17754) );
  NANDN U18453 ( .A(n17752), .B(n17751), .Z(n17753) );
  NAND U18454 ( .A(n17754), .B(n17753), .Z(n17813) );
  NAND U18455 ( .A(n17756), .B(n17755), .Z(n17760) );
  NAND U18456 ( .A(n17758), .B(n17757), .Z(n17759) );
  NAND U18457 ( .A(n17760), .B(n17759), .Z(n17812) );
  XOR U18458 ( .A(n17813), .B(n17812), .Z(n17814) );
  XOR U18459 ( .A(n17800), .B(n17801), .Z(n17802) );
  NANDN U18460 ( .A(n17762), .B(n17761), .Z(n17766) );
  NAND U18461 ( .A(n17764), .B(n17763), .Z(n17765) );
  NAND U18462 ( .A(n17766), .B(n17765), .Z(n17808) );
  NANDN U18463 ( .A(n17768), .B(n17767), .Z(n17772) );
  NAND U18464 ( .A(n17770), .B(n17769), .Z(n17771) );
  NAND U18465 ( .A(n17772), .B(n17771), .Z(n17806) );
  NAND U18466 ( .A(n17774), .B(n17773), .Z(n17778) );
  NANDN U18467 ( .A(n17776), .B(n17775), .Z(n17777) );
  AND U18468 ( .A(n17778), .B(n17777), .Z(n17807) );
  XNOR U18469 ( .A(n17806), .B(n17807), .Z(n17809) );
  XNOR U18470 ( .A(n17802), .B(n17803), .Z(n17795) );
  XNOR U18471 ( .A(n17796), .B(n17795), .Z(n17799) );
  NANDN U18472 ( .A(n17779), .B(n17780), .Z(n17785) );
  NOR U18473 ( .A(n17781), .B(n17780), .Z(n17783) );
  OR U18474 ( .A(n17783), .B(n17782), .Z(n17784) );
  AND U18475 ( .A(n17785), .B(n17784), .Z(n17798) );
  NANDN U18476 ( .A(n17787), .B(n17786), .Z(n17791) );
  NAND U18477 ( .A(n17789), .B(n17788), .Z(n17790) );
  AND U18478 ( .A(n17791), .B(n17790), .Z(n17797) );
  XOR U18479 ( .A(n17798), .B(n17797), .Z(n17792) );
  XNOR U18480 ( .A(n17799), .B(n17792), .Z(N381) );
  NAND U18481 ( .A(n17801), .B(n17800), .Z(n17805) );
  NANDN U18482 ( .A(n17803), .B(n17802), .Z(n17804) );
  NAND U18483 ( .A(n17805), .B(n17804), .Z(n17931) );
  NAND U18484 ( .A(n17807), .B(n17806), .Z(n17811) );
  NANDN U18485 ( .A(n17809), .B(n17808), .Z(n17810) );
  NAND U18486 ( .A(n17811), .B(n17810), .Z(n17929) );
  NAND U18487 ( .A(n17813), .B(n17812), .Z(n17817) );
  NANDN U18488 ( .A(n17815), .B(n17814), .Z(n17816) );
  NAND U18489 ( .A(n17817), .B(n17816), .Z(n17935) );
  NANDN U18490 ( .A(n17819), .B(n17818), .Z(n17823) );
  NANDN U18491 ( .A(n17821), .B(n17820), .Z(n17822) );
  AND U18492 ( .A(n17823), .B(n17822), .Z(n17936) );
  XOR U18493 ( .A(n17935), .B(n17936), .Z(n17938) );
  NAND U18494 ( .A(n17825), .B(n17824), .Z(n17829) );
  NAND U18495 ( .A(n17827), .B(n17826), .Z(n17828) );
  NAND U18496 ( .A(n17829), .B(n17828), .Z(n17947) );
  XOR U18497 ( .A(n18077), .B(n18078), .Z(n18079) );
  AND U18498 ( .A(x[234]), .B(y[1972]), .Z(n18075) );
  NAND U18499 ( .A(n17842), .B(n18075), .Z(n17846) );
  NAND U18500 ( .A(n17844), .B(n17843), .Z(n17845) );
  NAND U18501 ( .A(n17846), .B(n17845), .Z(n18052) );
  AND U18502 ( .A(x[246]), .B(y[1959]), .Z(n18026) );
  AND U18503 ( .A(x[225]), .B(y[1980]), .Z(n18024) );
  AND U18504 ( .A(x[236]), .B(y[1969]), .Z(n18236) );
  XOR U18505 ( .A(n18024), .B(n18236), .Z(n18025) );
  XOR U18506 ( .A(n18026), .B(n18025), .Z(n18051) );
  AND U18507 ( .A(x[239]), .B(y[1966]), .Z(n18027) );
  XOR U18508 ( .A(n18242), .B(n18027), .Z(n18029) );
  XOR U18509 ( .A(n18051), .B(n18050), .Z(n18053) );
  XNOR U18510 ( .A(n18052), .B(n18053), .Z(n18080) );
  XOR U18511 ( .A(n18079), .B(n18080), .Z(n18047) );
  XNOR U18512 ( .A(n18047), .B(n18046), .Z(n18049) );
  XOR U18513 ( .A(n18048), .B(n18049), .Z(n18044) );
  XOR U18514 ( .A(n18056), .B(n18057), .Z(n18058) );
  AND U18515 ( .A(x[235]), .B(y[1970]), .Z(n18002) );
  AND U18516 ( .A(x[227]), .B(y[1978]), .Z(n18000) );
  AND U18517 ( .A(x[241]), .B(y[1964]), .Z(n17999) );
  XOR U18518 ( .A(n18000), .B(n17999), .Z(n18001) );
  XOR U18519 ( .A(n18002), .B(n18001), .Z(n17970) );
  AND U18520 ( .A(x[247]), .B(y[1958]), .Z(n17996) );
  AND U18521 ( .A(x[237]), .B(y[1968]), .Z(n17994) );
  AND U18522 ( .A(x[248]), .B(y[1957]), .Z(n18250) );
  XOR U18523 ( .A(n17994), .B(n18250), .Z(n17995) );
  XOR U18524 ( .A(n17996), .B(n17995), .Z(n17969) );
  XOR U18525 ( .A(n17970), .B(n17969), .Z(n17971) );
  XNOR U18526 ( .A(n17972), .B(n17971), .Z(n18059) );
  XOR U18527 ( .A(n18058), .B(n18059), .Z(n17961) );
  AND U18528 ( .A(x[249]), .B(y[1956]), .Z(n18023) );
  AND U18529 ( .A(x[250]), .B(y[1955]), .Z(n18020) );
  XOR U18530 ( .A(n18021), .B(n18020), .Z(n18022) );
  XOR U18531 ( .A(n18023), .B(n18022), .Z(n18061) );
  AND U18532 ( .A(x[252]), .B(y[1953]), .Z(n18035) );
  XOR U18533 ( .A(o[189]), .B(n18035), .Z(n18072) );
  AND U18534 ( .A(x[224]), .B(y[1981]), .Z(n18070) );
  AND U18535 ( .A(x[253]), .B(y[1952]), .Z(n18069) );
  XOR U18536 ( .A(n18070), .B(n18069), .Z(n18071) );
  XOR U18537 ( .A(n18072), .B(n18071), .Z(n18060) );
  XOR U18538 ( .A(n18061), .B(n18060), .Z(n18062) );
  XOR U18539 ( .A(n18063), .B(n18062), .Z(n17959) );
  ANDN U18540 ( .B(o[188]), .A(n17870), .Z(n17989) );
  AND U18541 ( .A(x[240]), .B(y[1965]), .Z(n17987) );
  AND U18542 ( .A(x[251]), .B(y[1954]), .Z(n17986) );
  XOR U18543 ( .A(n17987), .B(n17986), .Z(n17988) );
  XOR U18544 ( .A(n17989), .B(n17988), .Z(n18013) );
  AND U18545 ( .A(x[226]), .B(y[1979]), .Z(n17979) );
  XOR U18546 ( .A(n17982), .B(n17981), .Z(n18012) );
  XOR U18547 ( .A(n18013), .B(n18012), .Z(n18016) );
  XOR U18548 ( .A(n18015), .B(n18016), .Z(n17960) );
  XNOR U18549 ( .A(n17959), .B(n17960), .Z(n17962) );
  XOR U18550 ( .A(n17961), .B(n17962), .Z(n17965) );
  XOR U18551 ( .A(n17990), .B(n17991), .Z(n17993) );
  AND U18552 ( .A(x[229]), .B(y[1976]), .Z(n17975) );
  AND U18553 ( .A(x[228]), .B(y[1977]), .Z(n17974) );
  AND U18554 ( .A(x[234]), .B(y[1971]), .Z(n17973) );
  XNOR U18555 ( .A(n17974), .B(n17973), .Z(n17976) );
  XNOR U18556 ( .A(n17975), .B(n17976), .Z(n18066) );
  AND U18557 ( .A(x[233]), .B(y[1972]), .Z(n18174) );
  AND U18558 ( .A(x[232]), .B(y[1973]), .Z(n18007) );
  AND U18559 ( .A(y[1975]), .B(x[230]), .Z(n17880) );
  NAND U18560 ( .A(y[1974]), .B(x[231]), .Z(n17879) );
  XNOR U18561 ( .A(n17880), .B(n17879), .Z(n18006) );
  XOR U18562 ( .A(n18007), .B(n18006), .Z(n18064) );
  XOR U18563 ( .A(n18174), .B(n18064), .Z(n18065) );
  XOR U18564 ( .A(n18066), .B(n18065), .Z(n17992) );
  XOR U18565 ( .A(n17993), .B(n17992), .Z(n17964) );
  XOR U18566 ( .A(n17964), .B(n17963), .Z(n17966) );
  XOR U18567 ( .A(n17965), .B(n17966), .Z(n18042) );
  XOR U18568 ( .A(n18042), .B(n18043), .Z(n18045) );
  XOR U18569 ( .A(n18044), .B(n18045), .Z(n17948) );
  XOR U18570 ( .A(n17947), .B(n17948), .Z(n17950) );
  NAND U18571 ( .A(n17890), .B(n17889), .Z(n17894) );
  NAND U18572 ( .A(n17892), .B(n17891), .Z(n17893) );
  NAND U18573 ( .A(n17894), .B(n17893), .Z(n17941) );
  NANDN U18574 ( .A(n17896), .B(n17895), .Z(n17900) );
  NANDN U18575 ( .A(n17898), .B(n17897), .Z(n17899) );
  AND U18576 ( .A(n17900), .B(n17899), .Z(n17942) );
  XOR U18577 ( .A(n17941), .B(n17942), .Z(n17943) );
  NAND U18578 ( .A(n17902), .B(n17901), .Z(n17906) );
  NAND U18579 ( .A(n17904), .B(n17903), .Z(n17905) );
  NAND U18580 ( .A(n17906), .B(n17905), .Z(n17955) );
  XOR U18581 ( .A(n18037), .B(n18038), .Z(n18040) );
  XOR U18582 ( .A(n18039), .B(n18040), .Z(n17954) );
  NANDN U18583 ( .A(n17920), .B(n17919), .Z(n17924) );
  NAND U18584 ( .A(n17922), .B(n17921), .Z(n17923) );
  NAND U18585 ( .A(n17924), .B(n17923), .Z(n17953) );
  XOR U18586 ( .A(n17954), .B(n17953), .Z(n17956) );
  XNOR U18587 ( .A(n17955), .B(n17956), .Z(n17944) );
  XOR U18588 ( .A(n17950), .B(n17949), .Z(n17937) );
  XOR U18589 ( .A(n17938), .B(n17937), .Z(n17930) );
  XOR U18590 ( .A(n17929), .B(n17930), .Z(n17932) );
  XOR U18591 ( .A(n17931), .B(n17932), .Z(n17928) );
  XOR U18592 ( .A(n17926), .B(n17928), .Z(n17925) );
  XOR U18593 ( .A(n17927), .B(n17925), .Z(N382) );
  NAND U18594 ( .A(n17930), .B(n17929), .Z(n17934) );
  NAND U18595 ( .A(n17932), .B(n17931), .Z(n17933) );
  AND U18596 ( .A(n17934), .B(n17933), .Z(n18343) );
  XNOR U18597 ( .A(n18344), .B(n18343), .Z(n18342) );
  NAND U18598 ( .A(n17936), .B(n17935), .Z(n17940) );
  NAND U18599 ( .A(n17938), .B(n17937), .Z(n17939) );
  NAND U18600 ( .A(n17940), .B(n17939), .Z(n18349) );
  NAND U18601 ( .A(n17942), .B(n17941), .Z(n17946) );
  NANDN U18602 ( .A(n17944), .B(n17943), .Z(n17945) );
  AND U18603 ( .A(n17946), .B(n17945), .Z(n18356) );
  NAND U18604 ( .A(n17948), .B(n17947), .Z(n17952) );
  NAND U18605 ( .A(n17950), .B(n17949), .Z(n17951) );
  AND U18606 ( .A(n17952), .B(n17951), .Z(n18355) );
  XOR U18607 ( .A(n18356), .B(n18355), .Z(n18358) );
  NAND U18608 ( .A(n17954), .B(n17953), .Z(n17958) );
  NAND U18609 ( .A(n17956), .B(n17955), .Z(n17957) );
  AND U18610 ( .A(n17958), .B(n17957), .Z(n18357) );
  XOR U18611 ( .A(n18358), .B(n18357), .Z(n18351) );
  NANDN U18612 ( .A(n17964), .B(n17963), .Z(n17968) );
  NANDN U18613 ( .A(n17966), .B(n17965), .Z(n17967) );
  AND U18614 ( .A(n17968), .B(n17967), .Z(n18321) );
  NAND U18615 ( .A(n17974), .B(n17973), .Z(n17978) );
  NANDN U18616 ( .A(n17976), .B(n17975), .Z(n17977) );
  AND U18617 ( .A(n17978), .B(n17977), .Z(n18096) );
  AND U18618 ( .A(x[230]), .B(y[1976]), .Z(n18125) );
  AND U18619 ( .A(x[229]), .B(y[1977]), .Z(n18127) );
  AND U18620 ( .A(x[243]), .B(y[1963]), .Z(n18126) );
  XOR U18621 ( .A(n18127), .B(n18126), .Z(n18124) );
  XOR U18622 ( .A(n18125), .B(n18124), .Z(n18275) );
  IV U18623 ( .A(n18275), .Z(n17985) );
  AND U18624 ( .A(x[228]), .B(y[1978]), .Z(n18204) );
  AND U18625 ( .A(x[227]), .B(y[1979]), .Z(n18206) );
  AND U18626 ( .A(x[242]), .B(y[1964]), .Z(n18205) );
  XOR U18627 ( .A(n18206), .B(n18205), .Z(n18203) );
  XNOR U18628 ( .A(n18204), .B(n18203), .Z(n18273) );
  NANDN U18629 ( .A(n17980), .B(n17979), .Z(n17984) );
  NAND U18630 ( .A(n17982), .B(n17981), .Z(n17983) );
  AND U18631 ( .A(n17984), .B(n17983), .Z(n18274) );
  XOR U18632 ( .A(n18273), .B(n18274), .Z(n18276) );
  XNOR U18633 ( .A(n17985), .B(n18276), .Z(n18097) );
  XNOR U18634 ( .A(n18096), .B(n18097), .Z(n18095) );
  XOR U18635 ( .A(n18095), .B(n18094), .Z(n18084) );
  XOR U18636 ( .A(n18085), .B(n18084), .Z(n18082) );
  XOR U18637 ( .A(n18082), .B(n18081), .Z(n18324) );
  NAND U18638 ( .A(n17994), .B(n18250), .Z(n17998) );
  NAND U18639 ( .A(n17996), .B(n17995), .Z(n17997) );
  NAND U18640 ( .A(n17998), .B(n17997), .Z(n18091) );
  NAND U18641 ( .A(n18000), .B(n17999), .Z(n18004) );
  NAND U18642 ( .A(n18002), .B(n18001), .Z(n18003) );
  AND U18643 ( .A(n18004), .B(n18003), .Z(n18101) );
  AND U18644 ( .A(x[224]), .B(y[1982]), .Z(n18178) );
  AND U18645 ( .A(x[253]), .B(y[1953]), .Z(n18156) );
  XOR U18646 ( .A(o[190]), .B(n18156), .Z(n18180) );
  AND U18647 ( .A(x[254]), .B(y[1952]), .Z(n18179) );
  XOR U18648 ( .A(n18180), .B(n18179), .Z(n18177) );
  XOR U18649 ( .A(n18178), .B(n18177), .Z(n18103) );
  AND U18650 ( .A(x[244]), .B(y[1962]), .Z(n18199) );
  AND U18651 ( .A(x[232]), .B(y[1974]), .Z(n18197) );
  XNOR U18652 ( .A(n18198), .B(n18197), .Z(n18102) );
  XNOR U18653 ( .A(n18101), .B(n18100), .Z(n18090) );
  XOR U18654 ( .A(n18091), .B(n18090), .Z(n18088) );
  AND U18655 ( .A(x[231]), .B(y[1975]), .Z(n18240) );
  NAND U18656 ( .A(n18005), .B(n18240), .Z(n18009) );
  NAND U18657 ( .A(n18007), .B(n18006), .Z(n18008) );
  AND U18658 ( .A(n18009), .B(n18008), .Z(n18110) );
  AND U18659 ( .A(y[1961]), .B(x[245]), .Z(n18011) );
  AND U18660 ( .A(y[1960]), .B(x[246]), .Z(n18010) );
  XOR U18661 ( .A(n18011), .B(n18010), .Z(n18239) );
  XOR U18662 ( .A(n18240), .B(n18239), .Z(n18113) );
  AND U18663 ( .A(x[241]), .B(y[1965]), .Z(n18254) );
  AND U18664 ( .A(x[226]), .B(y[1980]), .Z(n18256) );
  AND U18665 ( .A(x[250]), .B(y[1956]), .Z(n18255) );
  XOR U18666 ( .A(n18256), .B(n18255), .Z(n18253) );
  XNOR U18667 ( .A(n18254), .B(n18253), .Z(n18112) );
  XNOR U18668 ( .A(n18110), .B(n18111), .Z(n18089) );
  XNOR U18669 ( .A(n18088), .B(n18089), .Z(n18306) );
  IV U18670 ( .A(n18012), .Z(n18014) );
  NANDN U18671 ( .A(n18014), .B(n18013), .Z(n18019) );
  IV U18672 ( .A(n18015), .Z(n18017) );
  NANDN U18673 ( .A(n18017), .B(n18016), .Z(n18018) );
  NAND U18674 ( .A(n18019), .B(n18018), .Z(n18305) );
  XOR U18675 ( .A(n18306), .B(n18305), .Z(n18304) );
  IV U18676 ( .A(n18027), .Z(n18028) );
  NANDN U18677 ( .A(n18028), .B(n18242), .Z(n18032) );
  NANDN U18678 ( .A(n18030), .B(n18029), .Z(n18031) );
  AND U18679 ( .A(n18032), .B(n18031), .Z(n18107) );
  AND U18680 ( .A(x[247]), .B(y[1959]), .Z(n18248) );
  AND U18681 ( .A(y[1958]), .B(x[248]), .Z(n18034) );
  AND U18682 ( .A(y[1957]), .B(x[249]), .Z(n18033) );
  XOR U18683 ( .A(n18034), .B(n18033), .Z(n18247) );
  XOR U18684 ( .A(n18248), .B(n18247), .Z(n18109) );
  IV U18685 ( .A(n18109), .Z(n18036) );
  AND U18686 ( .A(x[252]), .B(y[1954]), .Z(n18216) );
  AND U18687 ( .A(x[240]), .B(y[1966]), .Z(n18215) );
  XOR U18688 ( .A(n18216), .B(n18215), .Z(n18213) );
  XNOR U18689 ( .A(n18214), .B(n18213), .Z(n18108) );
  XOR U18690 ( .A(n18036), .B(n18108), .Z(n18106) );
  XNOR U18691 ( .A(n18107), .B(n18106), .Z(n18116) );
  XOR U18692 ( .A(n18117), .B(n18116), .Z(n18115) );
  XOR U18693 ( .A(n18114), .B(n18115), .Z(n18303) );
  XOR U18694 ( .A(n18304), .B(n18303), .Z(n18323) );
  XNOR U18695 ( .A(n18321), .B(n18322), .Z(n18336) );
  XOR U18696 ( .A(n18336), .B(n18333), .Z(n18041) );
  XOR U18697 ( .A(n18334), .B(n18041), .Z(n18316) );
  NAND U18698 ( .A(n18051), .B(n18050), .Z(n18055) );
  NAND U18699 ( .A(n18053), .B(n18052), .Z(n18054) );
  AND U18700 ( .A(n18055), .B(n18054), .Z(n18290) );
  XOR U18701 ( .A(n18290), .B(n18289), .Z(n18288) );
  XOR U18702 ( .A(n18288), .B(n18287), .Z(n18300) );
  NAND U18703 ( .A(n18174), .B(n18064), .Z(n18068) );
  NAND U18704 ( .A(n18066), .B(n18065), .Z(n18067) );
  AND U18705 ( .A(n18068), .B(n18067), .Z(n18283) );
  NAND U18706 ( .A(y[1970]), .B(x[236]), .Z(n18073) );
  XNOR U18707 ( .A(n18074), .B(n18073), .Z(n18233) );
  AND U18708 ( .A(y[1973]), .B(x[233]), .Z(n18076) );
  XOR U18709 ( .A(n18076), .B(n18075), .Z(n18170) );
  XOR U18710 ( .A(n18171), .B(n18170), .Z(n18270) );
  AND U18711 ( .A(x[251]), .B(y[1955]), .Z(n18121) );
  AND U18712 ( .A(x[225]), .B(y[1981]), .Z(n18120) );
  XOR U18713 ( .A(n18121), .B(n18120), .Z(n18119) );
  XOR U18714 ( .A(n18119), .B(n18118), .Z(n18269) );
  XOR U18715 ( .A(n18270), .B(n18269), .Z(n18268) );
  XOR U18716 ( .A(n18267), .B(n18268), .Z(n18284) );
  XNOR U18717 ( .A(n18281), .B(n18282), .Z(n18299) );
  XNOR U18718 ( .A(n18297), .B(n18298), .Z(n18318) );
  XOR U18719 ( .A(n18317), .B(n18318), .Z(n18315) );
  XOR U18720 ( .A(n18316), .B(n18315), .Z(n18352) );
  XOR U18721 ( .A(n18349), .B(n18350), .Z(n18341) );
  XNOR U18722 ( .A(n18342), .B(n18341), .Z(N383) );
  IV U18723 ( .A(n18081), .Z(n18083) );
  NANDN U18724 ( .A(n18083), .B(n18082), .Z(n18087) );
  NAND U18725 ( .A(n18085), .B(n18084), .Z(n18086) );
  AND U18726 ( .A(n18087), .B(n18086), .Z(n18332) );
  NANDN U18727 ( .A(n18089), .B(n18088), .Z(n18093) );
  NAND U18728 ( .A(n18091), .B(n18090), .Z(n18092) );
  AND U18729 ( .A(n18093), .B(n18092), .Z(n18314) );
  NAND U18730 ( .A(n18095), .B(n18094), .Z(n18099) );
  NANDN U18731 ( .A(n18097), .B(n18096), .Z(n18098) );
  AND U18732 ( .A(n18099), .B(n18098), .Z(n18296) );
  NAND U18733 ( .A(n18101), .B(n18100), .Z(n18105) );
  NANDN U18734 ( .A(n18103), .B(n18102), .Z(n18104) );
  AND U18735 ( .A(n18105), .B(n18104), .Z(n18280) );
  NAND U18736 ( .A(n18119), .B(n18118), .Z(n18123) );
  NAND U18737 ( .A(n18121), .B(n18120), .Z(n18122) );
  AND U18738 ( .A(n18123), .B(n18122), .Z(n18131) );
  NAND U18739 ( .A(n18125), .B(n18124), .Z(n18129) );
  NAND U18740 ( .A(n18127), .B(n18126), .Z(n18128) );
  NAND U18741 ( .A(n18129), .B(n18128), .Z(n18130) );
  XNOR U18742 ( .A(n18131), .B(n18130), .Z(n18196) );
  AND U18743 ( .A(y[1967]), .B(x[240]), .Z(n18133) );
  NAND U18744 ( .A(y[1963]), .B(x[244]), .Z(n18132) );
  XNOR U18745 ( .A(n18133), .B(n18132), .Z(n18137) );
  AND U18746 ( .A(y[1953]), .B(x[254]), .Z(n18135) );
  NAND U18747 ( .A(y[1954]), .B(x[253]), .Z(n18134) );
  XNOR U18748 ( .A(n18135), .B(n18134), .Z(n18136) );
  XOR U18749 ( .A(n18137), .B(n18136), .Z(n18139) );
  AND U18750 ( .A(x[234]), .B(y[1973]), .Z(n18173) );
  XNOR U18751 ( .A(n18235), .B(n18173), .Z(n18138) );
  XNOR U18752 ( .A(n18139), .B(n18138), .Z(n18155) );
  AND U18753 ( .A(y[1978]), .B(x[229]), .Z(n18141) );
  NAND U18754 ( .A(y[1977]), .B(x[230]), .Z(n18140) );
  XNOR U18755 ( .A(n18141), .B(n18140), .Z(n18145) );
  AND U18756 ( .A(y[1976]), .B(x[231]), .Z(n18143) );
  NAND U18757 ( .A(y[1981]), .B(x[226]), .Z(n18142) );
  XNOR U18758 ( .A(n18143), .B(n18142), .Z(n18144) );
  XOR U18759 ( .A(n18145), .B(n18144), .Z(n18153) );
  AND U18760 ( .A(y[1980]), .B(x[227]), .Z(n18147) );
  NAND U18761 ( .A(y[1965]), .B(x[242]), .Z(n18146) );
  XNOR U18762 ( .A(n18147), .B(n18146), .Z(n18151) );
  AND U18763 ( .A(y[1952]), .B(x[255]), .Z(n18149) );
  NAND U18764 ( .A(y[1979]), .B(x[228]), .Z(n18148) );
  XNOR U18765 ( .A(n18149), .B(n18148), .Z(n18150) );
  XNOR U18766 ( .A(n18151), .B(n18150), .Z(n18152) );
  XNOR U18767 ( .A(n18153), .B(n18152), .Z(n18154) );
  XOR U18768 ( .A(n18155), .B(n18154), .Z(n18169) );
  AND U18769 ( .A(y[1975]), .B(x[232]), .Z(n18163) );
  AND U18770 ( .A(n18156), .B(o[190]), .Z(n18161) );
  AND U18771 ( .A(x[249]), .B(y[1958]), .Z(n18249) );
  XOR U18772 ( .A(n18249), .B(o[191]), .Z(n18159) );
  AND U18773 ( .A(x[246]), .B(y[1961]), .Z(n18241) );
  XNOR U18774 ( .A(n18157), .B(n18241), .Z(n18158) );
  XNOR U18775 ( .A(n18159), .B(n18158), .Z(n18160) );
  XNOR U18776 ( .A(n18161), .B(n18160), .Z(n18162) );
  XNOR U18777 ( .A(n18163), .B(n18162), .Z(n18167) );
  AND U18778 ( .A(y[1969]), .B(x[238]), .Z(n18165) );
  NAND U18779 ( .A(y[1974]), .B(x[233]), .Z(n18164) );
  XNOR U18780 ( .A(n18165), .B(n18164), .Z(n18166) );
  XNOR U18781 ( .A(n18167), .B(n18166), .Z(n18168) );
  XNOR U18782 ( .A(n18169), .B(n18168), .Z(n18186) );
  IV U18783 ( .A(n18170), .Z(n18172) );
  NANDN U18784 ( .A(n18172), .B(n18171), .Z(n18176) );
  NAND U18785 ( .A(n18174), .B(n18173), .Z(n18175) );
  AND U18786 ( .A(n18176), .B(n18175), .Z(n18184) );
  NAND U18787 ( .A(n18178), .B(n18177), .Z(n18182) );
  NAND U18788 ( .A(n18180), .B(n18179), .Z(n18181) );
  NAND U18789 ( .A(n18182), .B(n18181), .Z(n18183) );
  XNOR U18790 ( .A(n18184), .B(n18183), .Z(n18185) );
  XOR U18791 ( .A(n18186), .B(n18185), .Z(n18194) );
  AND U18792 ( .A(y[1964]), .B(x[243]), .Z(n18188) );
  NAND U18793 ( .A(y[1962]), .B(x[245]), .Z(n18187) );
  XNOR U18794 ( .A(n18188), .B(n18187), .Z(n18192) );
  AND U18795 ( .A(y[1982]), .B(x[225]), .Z(n18190) );
  NAND U18796 ( .A(y[1983]), .B(x[224]), .Z(n18189) );
  XNOR U18797 ( .A(n18190), .B(n18189), .Z(n18191) );
  XNOR U18798 ( .A(n18192), .B(n18191), .Z(n18193) );
  XNOR U18799 ( .A(n18194), .B(n18193), .Z(n18195) );
  NAND U18800 ( .A(n18198), .B(n18197), .Z(n18202) );
  NANDN U18801 ( .A(n18200), .B(n18199), .Z(n18201) );
  AND U18802 ( .A(n18202), .B(n18201), .Z(n18210) );
  NAND U18803 ( .A(n18204), .B(n18203), .Z(n18208) );
  NAND U18804 ( .A(n18206), .B(n18205), .Z(n18207) );
  NAND U18805 ( .A(n18208), .B(n18207), .Z(n18209) );
  XNOR U18806 ( .A(n18210), .B(n18209), .Z(n18266) );
  AND U18807 ( .A(y[1972]), .B(x[235]), .Z(n18212) );
  NAND U18808 ( .A(y[1957]), .B(x[250]), .Z(n18211) );
  XNOR U18809 ( .A(n18212), .B(n18211), .Z(n18232) );
  NAND U18810 ( .A(n18214), .B(n18213), .Z(n18218) );
  NAND U18811 ( .A(n18216), .B(n18215), .Z(n18217) );
  AND U18812 ( .A(n18218), .B(n18217), .Z(n18230) );
  AND U18813 ( .A(y[1971]), .B(x[236]), .Z(n18220) );
  NAND U18814 ( .A(y[1955]), .B(x[252]), .Z(n18219) );
  XNOR U18815 ( .A(n18220), .B(n18219), .Z(n18228) );
  AND U18816 ( .A(y[1966]), .B(x[241]), .Z(n18226) );
  AND U18817 ( .A(y[1956]), .B(x[251]), .Z(n18222) );
  NAND U18818 ( .A(y[1960]), .B(x[247]), .Z(n18221) );
  XNOR U18819 ( .A(n18222), .B(n18221), .Z(n18223) );
  XNOR U18820 ( .A(n18224), .B(n18223), .Z(n18225) );
  XNOR U18821 ( .A(n18226), .B(n18225), .Z(n18227) );
  XNOR U18822 ( .A(n18228), .B(n18227), .Z(n18229) );
  XNOR U18823 ( .A(n18230), .B(n18229), .Z(n18231) );
  XOR U18824 ( .A(n18232), .B(n18231), .Z(n18264) );
  NANDN U18825 ( .A(n18234), .B(n18233), .Z(n18238) );
  NAND U18826 ( .A(n18236), .B(n18235), .Z(n18237) );
  AND U18827 ( .A(n18238), .B(n18237), .Z(n18246) );
  NAND U18828 ( .A(n18240), .B(n18239), .Z(n18244) );
  NAND U18829 ( .A(n18242), .B(n18241), .Z(n18243) );
  NAND U18830 ( .A(n18244), .B(n18243), .Z(n18245) );
  XNOR U18831 ( .A(n18246), .B(n18245), .Z(n18262) );
  NAND U18832 ( .A(n18248), .B(n18247), .Z(n18252) );
  NAND U18833 ( .A(n18250), .B(n18249), .Z(n18251) );
  AND U18834 ( .A(n18252), .B(n18251), .Z(n18260) );
  NAND U18835 ( .A(n18254), .B(n18253), .Z(n18258) );
  NAND U18836 ( .A(n18256), .B(n18255), .Z(n18257) );
  NAND U18837 ( .A(n18258), .B(n18257), .Z(n18259) );
  XNOR U18838 ( .A(n18260), .B(n18259), .Z(n18261) );
  XNOR U18839 ( .A(n18262), .B(n18261), .Z(n18263) );
  XNOR U18840 ( .A(n18264), .B(n18263), .Z(n18265) );
  AND U18841 ( .A(n18270), .B(n18269), .Z(n18271) );
  AND U18842 ( .A(n18274), .B(n18273), .Z(n18278) );
  ANDN U18843 ( .B(n18276), .A(n18275), .Z(n18277) );
  XNOR U18844 ( .A(n18280), .B(n18279), .Z(n18294) );
  NAND U18845 ( .A(n18282), .B(n18281), .Z(n18286) );
  NANDN U18846 ( .A(n18284), .B(n18283), .Z(n18285) );
  AND U18847 ( .A(n18286), .B(n18285), .Z(n18292) );
  XNOR U18848 ( .A(n18292), .B(n18291), .Z(n18293) );
  XNOR U18849 ( .A(n18294), .B(n18293), .Z(n18295) );
  XNOR U18850 ( .A(n18296), .B(n18295), .Z(n18312) );
  NANDN U18851 ( .A(n18298), .B(n18297), .Z(n18302) );
  NANDN U18852 ( .A(n18300), .B(n18299), .Z(n18301) );
  AND U18853 ( .A(n18302), .B(n18301), .Z(n18310) );
  NAND U18854 ( .A(n18304), .B(n18303), .Z(n18308) );
  NAND U18855 ( .A(n18306), .B(n18305), .Z(n18307) );
  NAND U18856 ( .A(n18308), .B(n18307), .Z(n18309) );
  XNOR U18857 ( .A(n18310), .B(n18309), .Z(n18311) );
  XNOR U18858 ( .A(n18312), .B(n18311), .Z(n18313) );
  XNOR U18859 ( .A(n18314), .B(n18313), .Z(n18330) );
  NAND U18860 ( .A(n18316), .B(n18315), .Z(n18320) );
  NAND U18861 ( .A(n18318), .B(n18317), .Z(n18319) );
  AND U18862 ( .A(n18320), .B(n18319), .Z(n18328) );
  NANDN U18863 ( .A(n18322), .B(n18321), .Z(n18326) );
  NANDN U18864 ( .A(n18324), .B(n18323), .Z(n18325) );
  NAND U18865 ( .A(n18326), .B(n18325), .Z(n18327) );
  XNOR U18866 ( .A(n18328), .B(n18327), .Z(n18329) );
  XNOR U18867 ( .A(n18330), .B(n18329), .Z(n18331) );
  XNOR U18868 ( .A(n18332), .B(n18331), .Z(n18340) );
  OR U18869 ( .A(n18333), .B(n18334), .Z(n18338) );
  AND U18870 ( .A(n18334), .B(n18333), .Z(n18335) );
  OR U18871 ( .A(n18336), .B(n18335), .Z(n18337) );
  NAND U18872 ( .A(n18338), .B(n18337), .Z(n18339) );
  XNOR U18873 ( .A(n18340), .B(n18339), .Z(n18348) );
  NAND U18874 ( .A(n18342), .B(n18341), .Z(n18346) );
  NANDN U18875 ( .A(n18344), .B(n18343), .Z(n18345) );
  NAND U18876 ( .A(n18346), .B(n18345), .Z(n18347) );
  XNOR U18877 ( .A(n18348), .B(n18347), .Z(n18364) );
  NANDN U18878 ( .A(n18350), .B(n18349), .Z(n18354) );
  ANDN U18879 ( .B(n18352), .A(n18351), .Z(n18353) );
  ANDN U18880 ( .B(n18354), .A(n18353), .Z(n18362) );
  AND U18881 ( .A(n18356), .B(n18355), .Z(n18360) );
  AND U18882 ( .A(n18358), .B(n18357), .Z(n18359) );
  OR U18883 ( .A(n18360), .B(n18359), .Z(n18361) );
  XNOR U18884 ( .A(n18362), .B(n18361), .Z(n18363) );
  XNOR U18885 ( .A(n18364), .B(n18363), .Z(N384) );
  AND U18886 ( .A(x[224]), .B(y[1984]), .Z(n19017) );
  XOR U18887 ( .A(n19017), .B(o[192]), .Z(N417) );
  AND U18888 ( .A(x[225]), .B(y[1984]), .Z(n18373) );
  AND U18889 ( .A(x[224]), .B(y[1985]), .Z(n18372) );
  XNOR U18890 ( .A(n18372), .B(o[193]), .Z(n18365) );
  XNOR U18891 ( .A(n18373), .B(n18365), .Z(n18367) );
  NAND U18892 ( .A(n19017), .B(o[192]), .Z(n18366) );
  XNOR U18893 ( .A(n18367), .B(n18366), .Z(N418) );
  NANDN U18894 ( .A(n18373), .B(n18365), .Z(n18369) );
  NAND U18895 ( .A(n18367), .B(n18366), .Z(n18368) );
  AND U18896 ( .A(n18369), .B(n18368), .Z(n18379) );
  AND U18897 ( .A(x[224]), .B(y[1986]), .Z(n18386) );
  XNOR U18898 ( .A(n18386), .B(o[194]), .Z(n18378) );
  XNOR U18899 ( .A(n18379), .B(n18378), .Z(n18381) );
  AND U18900 ( .A(y[1984]), .B(x[226]), .Z(n18371) );
  NAND U18901 ( .A(y[1985]), .B(x[225]), .Z(n18370) );
  XNOR U18902 ( .A(n18371), .B(n18370), .Z(n18375) );
  AND U18903 ( .A(n18372), .B(o[193]), .Z(n18374) );
  XNOR U18904 ( .A(n18375), .B(n18374), .Z(n18380) );
  XNOR U18905 ( .A(n18381), .B(n18380), .Z(N419) );
  NAND U18906 ( .A(x[226]), .B(y[1985]), .Z(n18393) );
  NANDN U18907 ( .A(n18393), .B(n18373), .Z(n18377) );
  NAND U18908 ( .A(n18375), .B(n18374), .Z(n18376) );
  AND U18909 ( .A(n18377), .B(n18376), .Z(n18399) );
  NANDN U18910 ( .A(n18379), .B(n18378), .Z(n18383) );
  NAND U18911 ( .A(n18381), .B(n18380), .Z(n18382) );
  AND U18912 ( .A(n18383), .B(n18382), .Z(n18398) );
  XNOR U18913 ( .A(n18399), .B(n18398), .Z(n18401) );
  AND U18914 ( .A(x[225]), .B(y[1986]), .Z(n18505) );
  XOR U18915 ( .A(n18505), .B(n18395), .Z(n18397) );
  AND U18916 ( .A(y[1984]), .B(x[227]), .Z(n18385) );
  NAND U18917 ( .A(y[1987]), .B(x[224]), .Z(n18384) );
  XNOR U18918 ( .A(n18385), .B(n18384), .Z(n18387) );
  NAND U18919 ( .A(n18386), .B(o[194]), .Z(n18388) );
  XOR U18920 ( .A(n18397), .B(n18396), .Z(n18400) );
  XOR U18921 ( .A(n18401), .B(n18400), .Z(N420) );
  AND U18922 ( .A(x[227]), .B(y[1987]), .Z(n18445) );
  NAND U18923 ( .A(n19017), .B(n18445), .Z(n18390) );
  NANDN U18924 ( .A(n18388), .B(n18387), .Z(n18389) );
  AND U18925 ( .A(n18390), .B(n18389), .Z(n18424) );
  AND U18926 ( .A(y[1988]), .B(x[224]), .Z(n18392) );
  NAND U18927 ( .A(y[1984]), .B(x[228]), .Z(n18391) );
  XNOR U18928 ( .A(n18392), .B(n18391), .Z(n18415) );
  ANDN U18929 ( .B(o[195]), .A(n18393), .Z(n18414) );
  XOR U18930 ( .A(n18415), .B(n18414), .Z(n18422) );
  AND U18931 ( .A(y[1986]), .B(x[226]), .Z(n18540) );
  NAND U18932 ( .A(y[1987]), .B(x[225]), .Z(n18394) );
  XNOR U18933 ( .A(n18540), .B(n18394), .Z(n18411) );
  AND U18934 ( .A(x[227]), .B(y[1985]), .Z(n18409) );
  XOR U18935 ( .A(o[196]), .B(n18409), .Z(n18410) );
  XOR U18936 ( .A(n18411), .B(n18410), .Z(n18421) );
  XOR U18937 ( .A(n18422), .B(n18421), .Z(n18423) );
  XOR U18938 ( .A(n18424), .B(n18423), .Z(n18420) );
  NANDN U18939 ( .A(n18399), .B(n18398), .Z(n18403) );
  NAND U18940 ( .A(n18401), .B(n18400), .Z(n18402) );
  NAND U18941 ( .A(n18403), .B(n18402), .Z(n18419) );
  XOR U18942 ( .A(n18418), .B(n18419), .Z(n18404) );
  XNOR U18943 ( .A(n18420), .B(n18404), .Z(N421) );
  AND U18944 ( .A(x[226]), .B(y[1987]), .Z(n18513) );
  AND U18945 ( .A(y[1986]), .B(x[227]), .Z(n18406) );
  NAND U18946 ( .A(y[1988]), .B(x[225]), .Z(n18405) );
  XNOR U18947 ( .A(n18406), .B(n18405), .Z(n18429) );
  AND U18948 ( .A(x[228]), .B(y[1985]), .Z(n18443) );
  XOR U18949 ( .A(o[197]), .B(n18443), .Z(n18428) );
  XOR U18950 ( .A(n18429), .B(n18428), .Z(n18432) );
  XOR U18951 ( .A(n18513), .B(n18432), .Z(n18434) );
  AND U18952 ( .A(y[1984]), .B(x[229]), .Z(n18408) );
  NAND U18953 ( .A(y[1989]), .B(x[224]), .Z(n18407) );
  XNOR U18954 ( .A(n18408), .B(n18407), .Z(n18438) );
  AND U18955 ( .A(o[196]), .B(n18409), .Z(n18437) );
  XOR U18956 ( .A(n18438), .B(n18437), .Z(n18433) );
  XOR U18957 ( .A(n18434), .B(n18433), .Z(n18457) );
  NAND U18958 ( .A(n18513), .B(n18505), .Z(n18413) );
  NAND U18959 ( .A(n18411), .B(n18410), .Z(n18412) );
  NAND U18960 ( .A(n18413), .B(n18412), .Z(n18455) );
  AND U18961 ( .A(x[228]), .B(y[1988]), .Z(n19205) );
  NAND U18962 ( .A(n19205), .B(n19017), .Z(n18417) );
  NAND U18963 ( .A(n18415), .B(n18414), .Z(n18416) );
  NAND U18964 ( .A(n18417), .B(n18416), .Z(n18454) );
  XOR U18965 ( .A(n18455), .B(n18454), .Z(n18456) );
  XNOR U18966 ( .A(n18457), .B(n18456), .Z(n18450) );
  NAND U18967 ( .A(n18422), .B(n18421), .Z(n18426) );
  NANDN U18968 ( .A(n18424), .B(n18423), .Z(n18425) );
  NAND U18969 ( .A(n18426), .B(n18425), .Z(n18448) );
  IV U18970 ( .A(n18448), .Z(n18447) );
  XOR U18971 ( .A(n18449), .B(n18447), .Z(n18427) );
  XNOR U18972 ( .A(n18450), .B(n18427), .Z(N422) );
  AND U18973 ( .A(x[227]), .B(y[1988]), .Z(n18514) );
  NAND U18974 ( .A(n18514), .B(n18505), .Z(n18431) );
  NAND U18975 ( .A(n18429), .B(n18428), .Z(n18430) );
  NAND U18976 ( .A(n18431), .B(n18430), .Z(n18486) );
  NAND U18977 ( .A(n18513), .B(n18432), .Z(n18436) );
  NAND U18978 ( .A(n18434), .B(n18433), .Z(n18435) );
  NAND U18979 ( .A(n18436), .B(n18435), .Z(n18485) );
  XOR U18980 ( .A(n18486), .B(n18485), .Z(n18488) );
  AND U18981 ( .A(x[229]), .B(y[1989]), .Z(n18684) );
  NAND U18982 ( .A(n19017), .B(n18684), .Z(n18440) );
  NAND U18983 ( .A(n18438), .B(n18437), .Z(n18439) );
  NAND U18984 ( .A(n18440), .B(n18439), .Z(n18462) );
  AND U18985 ( .A(y[1984]), .B(x[230]), .Z(n18442) );
  NAND U18986 ( .A(y[1990]), .B(x[224]), .Z(n18441) );
  XNOR U18987 ( .A(n18442), .B(n18441), .Z(n18469) );
  AND U18988 ( .A(o[197]), .B(n18443), .Z(n18468) );
  XOR U18989 ( .A(n18469), .B(n18468), .Z(n18461) );
  XOR U18990 ( .A(n18462), .B(n18461), .Z(n18464) );
  NAND U18991 ( .A(y[1988]), .B(x[226]), .Z(n18444) );
  XNOR U18992 ( .A(n18445), .B(n18444), .Z(n18473) );
  AND U18993 ( .A(y[1989]), .B(x[225]), .Z(n18731) );
  NAND U18994 ( .A(y[1986]), .B(x[228]), .Z(n18446) );
  XNOR U18995 ( .A(n18731), .B(n18446), .Z(n18477) );
  AND U18996 ( .A(x[229]), .B(y[1985]), .Z(n18484) );
  XOR U18997 ( .A(o[198]), .B(n18484), .Z(n18476) );
  XOR U18998 ( .A(n18477), .B(n18476), .Z(n18472) );
  XOR U18999 ( .A(n18473), .B(n18472), .Z(n18463) );
  XOR U19000 ( .A(n18464), .B(n18463), .Z(n18487) );
  XOR U19001 ( .A(n18488), .B(n18487), .Z(n18494) );
  OR U19002 ( .A(n18449), .B(n18447), .Z(n18453) );
  ANDN U19003 ( .B(n18449), .A(n18448), .Z(n18451) );
  OR U19004 ( .A(n18451), .B(n18450), .Z(n18452) );
  AND U19005 ( .A(n18453), .B(n18452), .Z(n18492) );
  NAND U19006 ( .A(n18455), .B(n18454), .Z(n18459) );
  NAND U19007 ( .A(n18457), .B(n18456), .Z(n18458) );
  AND U19008 ( .A(n18459), .B(n18458), .Z(n18493) );
  IV U19009 ( .A(n18493), .Z(n18491) );
  XOR U19010 ( .A(n18492), .B(n18491), .Z(n18460) );
  XNOR U19011 ( .A(n18494), .B(n18460), .Z(N423) );
  NAND U19012 ( .A(n18462), .B(n18461), .Z(n18466) );
  NAND U19013 ( .A(n18464), .B(n18463), .Z(n18465) );
  AND U19014 ( .A(n18466), .B(n18465), .Z(n18536) );
  AND U19015 ( .A(y[1986]), .B(x[229]), .Z(n18596) );
  NAND U19016 ( .A(y[1990]), .B(x[225]), .Z(n18467) );
  XNOR U19017 ( .A(n18596), .B(n18467), .Z(n18507) );
  AND U19018 ( .A(x[230]), .B(y[1985]), .Z(n18510) );
  XOR U19019 ( .A(o[199]), .B(n18510), .Z(n18506) );
  XOR U19020 ( .A(n18507), .B(n18506), .Z(n18525) );
  AND U19021 ( .A(x[230]), .B(y[1990]), .Z(n18752) );
  NAND U19022 ( .A(n19017), .B(n18752), .Z(n18471) );
  NAND U19023 ( .A(n18469), .B(n18468), .Z(n18470) );
  AND U19024 ( .A(n18471), .B(n18470), .Z(n18524) );
  NAND U19025 ( .A(n18513), .B(n18514), .Z(n18475) );
  NAND U19026 ( .A(n18473), .B(n18472), .Z(n18474) );
  NAND U19027 ( .A(n18475), .B(n18474), .Z(n18527) );
  AND U19028 ( .A(x[228]), .B(y[1989]), .Z(n19022) );
  NAND U19029 ( .A(n19022), .B(n18505), .Z(n18479) );
  NAND U19030 ( .A(n18477), .B(n18476), .Z(n18478) );
  AND U19031 ( .A(n18479), .B(n18478), .Z(n18502) );
  AND U19032 ( .A(y[1989]), .B(x[226]), .Z(n18481) );
  NAND U19033 ( .A(y[1987]), .B(x[228]), .Z(n18480) );
  XNOR U19034 ( .A(n18481), .B(n18480), .Z(n18515) );
  XNOR U19035 ( .A(n18515), .B(n18514), .Z(n18500) );
  AND U19036 ( .A(y[1984]), .B(x[231]), .Z(n18483) );
  NAND U19037 ( .A(y[1991]), .B(x[224]), .Z(n18482) );
  XNOR U19038 ( .A(n18483), .B(n18482), .Z(n18519) );
  AND U19039 ( .A(o[198]), .B(n18484), .Z(n18518) );
  XNOR U19040 ( .A(n18519), .B(n18518), .Z(n18499) );
  XOR U19041 ( .A(n18500), .B(n18499), .Z(n18501) );
  XOR U19042 ( .A(n18502), .B(n18501), .Z(n18533) );
  XOR U19043 ( .A(n18534), .B(n18533), .Z(n18535) );
  XOR U19044 ( .A(n18536), .B(n18535), .Z(n18532) );
  NAND U19045 ( .A(n18486), .B(n18485), .Z(n18490) );
  NAND U19046 ( .A(n18488), .B(n18487), .Z(n18489) );
  NAND U19047 ( .A(n18490), .B(n18489), .Z(n18531) );
  NANDN U19048 ( .A(n18491), .B(n18492), .Z(n18497) );
  NOR U19049 ( .A(n18493), .B(n18492), .Z(n18495) );
  OR U19050 ( .A(n18495), .B(n18494), .Z(n18496) );
  AND U19051 ( .A(n18497), .B(n18496), .Z(n18530) );
  XOR U19052 ( .A(n18531), .B(n18530), .Z(n18498) );
  XNOR U19053 ( .A(n18532), .B(n18498), .Z(N424) );
  NAND U19054 ( .A(n18500), .B(n18499), .Z(n18504) );
  NAND U19055 ( .A(n18502), .B(n18501), .Z(n18503) );
  AND U19056 ( .A(n18504), .B(n18503), .Z(n18573) );
  AND U19057 ( .A(x[229]), .B(y[1990]), .Z(n18676) );
  NAND U19058 ( .A(n18676), .B(n18505), .Z(n18509) );
  NAND U19059 ( .A(n18507), .B(n18506), .Z(n18508) );
  NAND U19060 ( .A(n18509), .B(n18508), .Z(n18571) );
  AND U19061 ( .A(o[199]), .B(n18510), .Z(n18560) );
  AND U19062 ( .A(y[1987]), .B(x[229]), .Z(n19146) );
  NAND U19063 ( .A(y[1991]), .B(x[225]), .Z(n18511) );
  XNOR U19064 ( .A(n19146), .B(n18511), .Z(n18561) );
  XNOR U19065 ( .A(n18560), .B(n18561), .Z(n18545) );
  AND U19066 ( .A(x[227]), .B(y[1989]), .Z(n19332) );
  AND U19067 ( .A(x[230]), .B(y[1986]), .Z(n18512) );
  AND U19068 ( .A(y[1990]), .B(x[226]), .Z(n19419) );
  XOR U19069 ( .A(n18512), .B(n19419), .Z(n18541) );
  XNOR U19070 ( .A(n19205), .B(n18541), .Z(n18544) );
  XOR U19071 ( .A(n19332), .B(n18544), .Z(n18546) );
  XOR U19072 ( .A(n18545), .B(n18546), .Z(n18570) );
  XOR U19073 ( .A(n18571), .B(n18570), .Z(n18572) );
  XOR U19074 ( .A(n18573), .B(n18572), .Z(n18579) );
  NAND U19075 ( .A(n19022), .B(n18513), .Z(n18517) );
  NAND U19076 ( .A(n18515), .B(n18514), .Z(n18516) );
  NAND U19077 ( .A(n18517), .B(n18516), .Z(n18567) );
  AND U19078 ( .A(x[231]), .B(y[1991]), .Z(n18897) );
  NAND U19079 ( .A(n19017), .B(n18897), .Z(n18521) );
  NAND U19080 ( .A(n18519), .B(n18518), .Z(n18520) );
  NAND U19081 ( .A(n18521), .B(n18520), .Z(n18565) );
  AND U19082 ( .A(y[1984]), .B(x[232]), .Z(n18523) );
  NAND U19083 ( .A(y[1992]), .B(x[224]), .Z(n18522) );
  XNOR U19084 ( .A(n18523), .B(n18522), .Z(n18551) );
  AND U19085 ( .A(x[231]), .B(y[1985]), .Z(n18554) );
  XOR U19086 ( .A(o[200]), .B(n18554), .Z(n18550) );
  XOR U19087 ( .A(n18551), .B(n18550), .Z(n18564) );
  XOR U19088 ( .A(n18565), .B(n18564), .Z(n18566) );
  XNOR U19089 ( .A(n18567), .B(n18566), .Z(n18577) );
  NANDN U19090 ( .A(n18525), .B(n18524), .Z(n18529) );
  NANDN U19091 ( .A(n18527), .B(n18526), .Z(n18528) );
  NAND U19092 ( .A(n18529), .B(n18528), .Z(n18576) );
  XOR U19093 ( .A(n18577), .B(n18576), .Z(n18578) );
  XOR U19094 ( .A(n18579), .B(n18578), .Z(n18585) );
  NAND U19095 ( .A(n18534), .B(n18533), .Z(n18538) );
  NAND U19096 ( .A(n18536), .B(n18535), .Z(n18537) );
  NAND U19097 ( .A(n18538), .B(n18537), .Z(n18584) );
  IV U19098 ( .A(n18584), .Z(n18582) );
  XOR U19099 ( .A(n18583), .B(n18582), .Z(n18539) );
  XNOR U19100 ( .A(n18585), .B(n18539), .Z(N425) );
  NAND U19101 ( .A(n18752), .B(n18540), .Z(n18543) );
  NAND U19102 ( .A(n19205), .B(n18541), .Z(n18542) );
  NAND U19103 ( .A(n18543), .B(n18542), .Z(n18590) );
  NANDN U19104 ( .A(n19332), .B(n18544), .Z(n18548) );
  NANDN U19105 ( .A(n18546), .B(n18545), .Z(n18547) );
  AND U19106 ( .A(n18548), .B(n18547), .Z(n18591) );
  XOR U19107 ( .A(n18590), .B(n18591), .Z(n18592) );
  AND U19108 ( .A(x[232]), .B(y[1992]), .Z(n18549) );
  NAND U19109 ( .A(n18549), .B(n19017), .Z(n18553) );
  NAND U19110 ( .A(n18551), .B(n18550), .Z(n18552) );
  AND U19111 ( .A(n18553), .B(n18552), .Z(n18625) );
  AND U19112 ( .A(o[200]), .B(n18554), .Z(n18598) );
  AND U19113 ( .A(y[1988]), .B(x[229]), .Z(n18556) );
  NAND U19114 ( .A(y[1986]), .B(x[231]), .Z(n18555) );
  XNOR U19115 ( .A(n18556), .B(n18555), .Z(n18597) );
  XNOR U19116 ( .A(n18598), .B(n18597), .Z(n18623) );
  AND U19117 ( .A(y[1984]), .B(x[233]), .Z(n18558) );
  NAND U19118 ( .A(y[1993]), .B(x[224]), .Z(n18557) );
  XNOR U19119 ( .A(n18558), .B(n18557), .Z(n18605) );
  AND U19120 ( .A(x[232]), .B(y[1985]), .Z(n18614) );
  XOR U19121 ( .A(o[201]), .B(n18614), .Z(n18604) );
  XNOR U19122 ( .A(n18605), .B(n18604), .Z(n18622) );
  XOR U19123 ( .A(n18623), .B(n18622), .Z(n18624) );
  XNOR U19124 ( .A(n18625), .B(n18624), .Z(n18619) );
  AND U19125 ( .A(y[1987]), .B(x[230]), .Z(n18945) );
  NAND U19126 ( .A(y[1992]), .B(x[225]), .Z(n18559) );
  XNOR U19127 ( .A(n18945), .B(n18559), .Z(n18609) );
  XNOR U19128 ( .A(n19022), .B(n18609), .Z(n18629) );
  NAND U19129 ( .A(x[226]), .B(y[1991]), .Z(n19119) );
  NAND U19130 ( .A(x[227]), .B(y[1990]), .Z(n18955) );
  XOR U19131 ( .A(n19119), .B(n18955), .Z(n18628) );
  XNOR U19132 ( .A(n18629), .B(n18628), .Z(n18617) );
  NAND U19133 ( .A(x[229]), .B(y[1991]), .Z(n18814) );
  AND U19134 ( .A(x[225]), .B(y[1987]), .Z(n18608) );
  NANDN U19135 ( .A(n18814), .B(n18608), .Z(n18563) );
  NAND U19136 ( .A(n18561), .B(n18560), .Z(n18562) );
  NAND U19137 ( .A(n18563), .B(n18562), .Z(n18616) );
  XOR U19138 ( .A(n18617), .B(n18616), .Z(n18618) );
  XNOR U19139 ( .A(n18619), .B(n18618), .Z(n18593) );
  XNOR U19140 ( .A(n18592), .B(n18593), .Z(n18635) );
  NAND U19141 ( .A(n18565), .B(n18564), .Z(n18569) );
  NAND U19142 ( .A(n18567), .B(n18566), .Z(n18568) );
  NAND U19143 ( .A(n18569), .B(n18568), .Z(n18633) );
  NAND U19144 ( .A(n18571), .B(n18570), .Z(n18575) );
  NAND U19145 ( .A(n18573), .B(n18572), .Z(n18574) );
  NAND U19146 ( .A(n18575), .B(n18574), .Z(n18632) );
  XOR U19147 ( .A(n18633), .B(n18632), .Z(n18634) );
  XOR U19148 ( .A(n18635), .B(n18634), .Z(n18640) );
  NAND U19149 ( .A(n18577), .B(n18576), .Z(n18581) );
  NANDN U19150 ( .A(n18579), .B(n18578), .Z(n18580) );
  NAND U19151 ( .A(n18581), .B(n18580), .Z(n18638) );
  NANDN U19152 ( .A(n18582), .B(n18583), .Z(n18588) );
  NOR U19153 ( .A(n18584), .B(n18583), .Z(n18586) );
  OR U19154 ( .A(n18586), .B(n18585), .Z(n18587) );
  AND U19155 ( .A(n18588), .B(n18587), .Z(n18639) );
  XOR U19156 ( .A(n18638), .B(n18639), .Z(n18589) );
  XNOR U19157 ( .A(n18640), .B(n18589), .Z(N426) );
  NAND U19158 ( .A(n18591), .B(n18590), .Z(n18595) );
  NANDN U19159 ( .A(n18593), .B(n18592), .Z(n18594) );
  AND U19160 ( .A(n18595), .B(n18594), .Z(n18699) );
  AND U19161 ( .A(x[231]), .B(y[1988]), .Z(n18678) );
  NAND U19162 ( .A(n18678), .B(n18596), .Z(n18600) );
  NAND U19163 ( .A(n18598), .B(n18597), .Z(n18599) );
  AND U19164 ( .A(n18600), .B(n18599), .Z(n18691) );
  AND U19165 ( .A(y[1987]), .B(x[231]), .Z(n18602) );
  NAND U19166 ( .A(y[1990]), .B(x[228]), .Z(n18601) );
  XNOR U19167 ( .A(n18602), .B(n18601), .Z(n18662) );
  AND U19168 ( .A(x[230]), .B(y[1988]), .Z(n18661) );
  XNOR U19169 ( .A(n18662), .B(n18661), .Z(n18689) );
  AND U19170 ( .A(x[232]), .B(y[1986]), .Z(n18877) );
  AND U19171 ( .A(x[233]), .B(y[1985]), .Z(n18672) );
  XOR U19172 ( .A(o[202]), .B(n18672), .Z(n18683) );
  XOR U19173 ( .A(n18877), .B(n18683), .Z(n18685) );
  XNOR U19174 ( .A(n18685), .B(n18684), .Z(n18688) );
  XOR U19175 ( .A(n18689), .B(n18688), .Z(n18690) );
  XNOR U19176 ( .A(n18691), .B(n18690), .Z(n18651) );
  AND U19177 ( .A(x[233]), .B(y[1993]), .Z(n18603) );
  NAND U19178 ( .A(n18603), .B(n19017), .Z(n18607) );
  NAND U19179 ( .A(n18605), .B(n18604), .Z(n18606) );
  NAND U19180 ( .A(n18607), .B(n18606), .Z(n18649) );
  AND U19181 ( .A(x[230]), .B(y[1992]), .Z(n18903) );
  NAND U19182 ( .A(n18903), .B(n18608), .Z(n18611) );
  NAND U19183 ( .A(n19022), .B(n18609), .Z(n18610) );
  NAND U19184 ( .A(n18611), .B(n18610), .Z(n18657) );
  AND U19185 ( .A(y[1984]), .B(x[234]), .Z(n18613) );
  NAND U19186 ( .A(y[1994]), .B(x[224]), .Z(n18612) );
  XNOR U19187 ( .A(n18613), .B(n18612), .Z(n18667) );
  AND U19188 ( .A(o[201]), .B(n18614), .Z(n18666) );
  XOR U19189 ( .A(n18667), .B(n18666), .Z(n18655) );
  AND U19190 ( .A(y[1991]), .B(x[227]), .Z(n19564) );
  NAND U19191 ( .A(y[1993]), .B(x[225]), .Z(n18615) );
  XNOR U19192 ( .A(n19564), .B(n18615), .Z(n18679) );
  AND U19193 ( .A(x[226]), .B(y[1992]), .Z(n18680) );
  XOR U19194 ( .A(n18679), .B(n18680), .Z(n18654) );
  XOR U19195 ( .A(n18655), .B(n18654), .Z(n18656) );
  XOR U19196 ( .A(n18657), .B(n18656), .Z(n18648) );
  XOR U19197 ( .A(n18649), .B(n18648), .Z(n18650) );
  XOR U19198 ( .A(n18651), .B(n18650), .Z(n18698) );
  NAND U19199 ( .A(n18617), .B(n18616), .Z(n18621) );
  NAND U19200 ( .A(n18619), .B(n18618), .Z(n18620) );
  NAND U19201 ( .A(n18621), .B(n18620), .Z(n18645) );
  NAND U19202 ( .A(n18623), .B(n18622), .Z(n18627) );
  NAND U19203 ( .A(n18625), .B(n18624), .Z(n18626) );
  AND U19204 ( .A(n18627), .B(n18626), .Z(n18642) );
  NAND U19205 ( .A(n18629), .B(n18628), .Z(n18631) );
  IV U19206 ( .A(n19119), .Z(n19252) );
  ANDN U19207 ( .B(n18955), .A(n19252), .Z(n18630) );
  ANDN U19208 ( .B(n18631), .A(n18630), .Z(n18643) );
  XOR U19209 ( .A(n18642), .B(n18643), .Z(n18644) );
  XNOR U19210 ( .A(n18645), .B(n18644), .Z(n18697) );
  XNOR U19211 ( .A(n18699), .B(n18700), .Z(n18696) );
  NAND U19212 ( .A(n18633), .B(n18632), .Z(n18637) );
  NAND U19213 ( .A(n18635), .B(n18634), .Z(n18636) );
  NAND U19214 ( .A(n18637), .B(n18636), .Z(n18695) );
  XOR U19215 ( .A(n18695), .B(n18694), .Z(n18641) );
  XNOR U19216 ( .A(n18696), .B(n18641), .Z(N427) );
  NAND U19217 ( .A(n18643), .B(n18642), .Z(n18647) );
  NAND U19218 ( .A(n18645), .B(n18644), .Z(n18646) );
  AND U19219 ( .A(n18647), .B(n18646), .Z(n18769) );
  NAND U19220 ( .A(n18649), .B(n18648), .Z(n18653) );
  NAND U19221 ( .A(n18651), .B(n18650), .Z(n18652) );
  NAND U19222 ( .A(n18653), .B(n18652), .Z(n18767) );
  NAND U19223 ( .A(n18655), .B(n18654), .Z(n18659) );
  NAND U19224 ( .A(n18657), .B(n18656), .Z(n18658) );
  NAND U19225 ( .A(n18659), .B(n18658), .Z(n18718) );
  AND U19226 ( .A(x[231]), .B(y[1990]), .Z(n18810) );
  AND U19227 ( .A(x[228]), .B(y[1987]), .Z(n18660) );
  NAND U19228 ( .A(n18810), .B(n18660), .Z(n18664) );
  NAND U19229 ( .A(n18662), .B(n18661), .Z(n18663) );
  NAND U19230 ( .A(n18664), .B(n18663), .Z(n18716) );
  AND U19231 ( .A(x[234]), .B(y[1994]), .Z(n18665) );
  NAND U19232 ( .A(n18665), .B(n19017), .Z(n18669) );
  NAND U19233 ( .A(n18667), .B(n18666), .Z(n18668) );
  NAND U19234 ( .A(n18669), .B(n18668), .Z(n18712) );
  AND U19235 ( .A(y[1984]), .B(x[235]), .Z(n18671) );
  NAND U19236 ( .A(y[1995]), .B(x[224]), .Z(n18670) );
  XNOR U19237 ( .A(n18671), .B(n18670), .Z(n18743) );
  AND U19238 ( .A(o[202]), .B(n18672), .Z(n18742) );
  XOR U19239 ( .A(n18743), .B(n18742), .Z(n18710) );
  AND U19240 ( .A(y[1989]), .B(x[230]), .Z(n18674) );
  NAND U19241 ( .A(y[1994]), .B(x[225]), .Z(n18673) );
  XNOR U19242 ( .A(n18674), .B(n18673), .Z(n18733) );
  AND U19243 ( .A(x[234]), .B(y[1985]), .Z(n18751) );
  XOR U19244 ( .A(o[203]), .B(n18751), .Z(n18732) );
  XOR U19245 ( .A(n18733), .B(n18732), .Z(n18709) );
  XOR U19246 ( .A(n18710), .B(n18709), .Z(n18711) );
  XOR U19247 ( .A(n18712), .B(n18711), .Z(n18715) );
  XOR U19248 ( .A(n18716), .B(n18715), .Z(n18717) );
  XNOR U19249 ( .A(n18718), .B(n18717), .Z(n18755) );
  AND U19250 ( .A(x[227]), .B(y[1992]), .Z(n19697) );
  NAND U19251 ( .A(y[1993]), .B(x[226]), .Z(n18675) );
  XNOR U19252 ( .A(n18676), .B(n18675), .Z(n18728) );
  AND U19253 ( .A(x[228]), .B(y[1991]), .Z(n18727) );
  XNOR U19254 ( .A(n18728), .B(n18727), .Z(n18704) );
  XNOR U19255 ( .A(n19697), .B(n18704), .Z(n18706) );
  NAND U19256 ( .A(y[1986]), .B(x[233]), .Z(n18677) );
  XNOR U19257 ( .A(n18678), .B(n18677), .Z(n18748) );
  AND U19258 ( .A(x[232]), .B(y[1987]), .Z(n18747) );
  XNOR U19259 ( .A(n18748), .B(n18747), .Z(n18705) );
  XNOR U19260 ( .A(n18706), .B(n18705), .Z(n18724) );
  AND U19261 ( .A(x[227]), .B(y[1993]), .Z(n18741) );
  IV U19262 ( .A(n18741), .Z(n18805) );
  AND U19263 ( .A(x[225]), .B(y[1991]), .Z(n19012) );
  NANDN U19264 ( .A(n18805), .B(n19012), .Z(n18682) );
  NAND U19265 ( .A(n18680), .B(n18679), .Z(n18681) );
  NAND U19266 ( .A(n18682), .B(n18681), .Z(n18722) );
  NAND U19267 ( .A(n18877), .B(n18683), .Z(n18687) );
  NAND U19268 ( .A(n18685), .B(n18684), .Z(n18686) );
  NAND U19269 ( .A(n18687), .B(n18686), .Z(n18721) );
  XOR U19270 ( .A(n18722), .B(n18721), .Z(n18723) );
  XNOR U19271 ( .A(n18724), .B(n18723), .Z(n18754) );
  NAND U19272 ( .A(n18689), .B(n18688), .Z(n18693) );
  NAND U19273 ( .A(n18691), .B(n18690), .Z(n18692) );
  NAND U19274 ( .A(n18693), .B(n18692), .Z(n18753) );
  XOR U19275 ( .A(n18754), .B(n18753), .Z(n18756) );
  XNOR U19276 ( .A(n18755), .B(n18756), .Z(n18766) );
  XOR U19277 ( .A(n18767), .B(n18766), .Z(n18768) );
  XOR U19278 ( .A(n18769), .B(n18768), .Z(n18762) );
  NANDN U19279 ( .A(n18698), .B(n18697), .Z(n18702) );
  NANDN U19280 ( .A(n18700), .B(n18699), .Z(n18701) );
  AND U19281 ( .A(n18702), .B(n18701), .Z(n18760) );
  IV U19282 ( .A(n18760), .Z(n18759) );
  XOR U19283 ( .A(n18761), .B(n18759), .Z(n18703) );
  XNOR U19284 ( .A(n18762), .B(n18703), .Z(N428) );
  NANDN U19285 ( .A(n19697), .B(n18704), .Z(n18708) );
  NAND U19286 ( .A(n18706), .B(n18705), .Z(n18707) );
  NAND U19287 ( .A(n18708), .B(n18707), .Z(n18787) );
  NAND U19288 ( .A(n18710), .B(n18709), .Z(n18714) );
  NAND U19289 ( .A(n18712), .B(n18711), .Z(n18713) );
  AND U19290 ( .A(n18714), .B(n18713), .Z(n18786) );
  XOR U19291 ( .A(n18787), .B(n18786), .Z(n18788) );
  NAND U19292 ( .A(n18716), .B(n18715), .Z(n18720) );
  NAND U19293 ( .A(n18718), .B(n18717), .Z(n18719) );
  AND U19294 ( .A(n18720), .B(n18719), .Z(n18789) );
  XOR U19295 ( .A(n18788), .B(n18789), .Z(n18776) );
  NAND U19296 ( .A(n18722), .B(n18721), .Z(n18726) );
  NAND U19297 ( .A(n18724), .B(n18723), .Z(n18725) );
  NAND U19298 ( .A(n18726), .B(n18725), .Z(n18842) );
  AND U19299 ( .A(x[229]), .B(y[1993]), .Z(n19243) );
  NAND U19300 ( .A(n19419), .B(n19243), .Z(n18730) );
  NAND U19301 ( .A(n18728), .B(n18727), .Z(n18729) );
  NAND U19302 ( .A(n18730), .B(n18729), .Z(n18793) );
  AND U19303 ( .A(x[230]), .B(y[1994]), .Z(n19029) );
  NAND U19304 ( .A(n19029), .B(n18731), .Z(n18735) );
  NAND U19305 ( .A(n18733), .B(n18732), .Z(n18734) );
  NAND U19306 ( .A(n18735), .B(n18734), .Z(n18792) );
  XOR U19307 ( .A(n18793), .B(n18792), .Z(n18795) );
  AND U19308 ( .A(x[233]), .B(y[1987]), .Z(n19414) );
  AND U19309 ( .A(x[234]), .B(y[1986]), .Z(n19468) );
  AND U19310 ( .A(y[1992]), .B(x[228]), .Z(n18736) );
  XOR U19311 ( .A(n19468), .B(n18736), .Z(n18832) );
  XOR U19312 ( .A(n19414), .B(n18832), .Z(n18815) );
  NAND U19313 ( .A(x[231]), .B(y[1989]), .Z(n18813) );
  XOR U19314 ( .A(n18814), .B(n18813), .Z(n18816) );
  AND U19315 ( .A(y[1984]), .B(x[236]), .Z(n18738) );
  NAND U19316 ( .A(y[1996]), .B(x[224]), .Z(n18737) );
  XNOR U19317 ( .A(n18738), .B(n18737), .Z(n18828) );
  AND U19318 ( .A(x[235]), .B(y[1985]), .Z(n18808) );
  XOR U19319 ( .A(n18808), .B(o[204]), .Z(n18827) );
  XOR U19320 ( .A(n18828), .B(n18827), .Z(n18799) );
  AND U19321 ( .A(y[1994]), .B(x[226]), .Z(n18740) );
  NAND U19322 ( .A(y[1988]), .B(x[232]), .Z(n18739) );
  XNOR U19323 ( .A(n18740), .B(n18739), .Z(n18804) );
  XOR U19324 ( .A(n18804), .B(n18741), .Z(n18798) );
  XOR U19325 ( .A(n18799), .B(n18798), .Z(n18801) );
  XOR U19326 ( .A(n18800), .B(n18801), .Z(n18794) );
  XOR U19327 ( .A(n18795), .B(n18794), .Z(n18840) );
  AND U19328 ( .A(x[235]), .B(y[1995]), .Z(n19810) );
  NAND U19329 ( .A(n19810), .B(n19017), .Z(n18745) );
  NAND U19330 ( .A(n18743), .B(n18742), .Z(n18744) );
  NAND U19331 ( .A(n18745), .B(n18744), .Z(n18822) );
  AND U19332 ( .A(x[231]), .B(y[1986]), .Z(n18931) );
  AND U19333 ( .A(x[233]), .B(y[1988]), .Z(n18746) );
  NAND U19334 ( .A(n18931), .B(n18746), .Z(n18750) );
  NAND U19335 ( .A(n18748), .B(n18747), .Z(n18749) );
  NAND U19336 ( .A(n18750), .B(n18749), .Z(n18820) );
  AND U19337 ( .A(y[1995]), .B(x[225]), .Z(n19463) );
  XOR U19338 ( .A(n18752), .B(n19463), .Z(n18825) );
  XOR U19339 ( .A(n18826), .B(n18825), .Z(n18819) );
  XOR U19340 ( .A(n18820), .B(n18819), .Z(n18821) );
  XOR U19341 ( .A(n18822), .B(n18821), .Z(n18839) );
  XOR U19342 ( .A(n18840), .B(n18839), .Z(n18841) );
  XNOR U19343 ( .A(n18842), .B(n18841), .Z(n18774) );
  NAND U19344 ( .A(n18754), .B(n18753), .Z(n18758) );
  NAND U19345 ( .A(n18756), .B(n18755), .Z(n18757) );
  NAND U19346 ( .A(n18758), .B(n18757), .Z(n18773) );
  XOR U19347 ( .A(n18774), .B(n18773), .Z(n18775) );
  XNOR U19348 ( .A(n18776), .B(n18775), .Z(n18782) );
  OR U19349 ( .A(n18761), .B(n18759), .Z(n18765) );
  ANDN U19350 ( .B(n18761), .A(n18760), .Z(n18763) );
  OR U19351 ( .A(n18763), .B(n18762), .Z(n18764) );
  AND U19352 ( .A(n18765), .B(n18764), .Z(n18780) );
  NAND U19353 ( .A(n18767), .B(n18766), .Z(n18771) );
  NANDN U19354 ( .A(n18769), .B(n18768), .Z(n18770) );
  AND U19355 ( .A(n18771), .B(n18770), .Z(n18781) );
  IV U19356 ( .A(n18781), .Z(n18779) );
  XOR U19357 ( .A(n18780), .B(n18779), .Z(n18772) );
  XNOR U19358 ( .A(n18782), .B(n18772), .Z(N429) );
  NAND U19359 ( .A(n18774), .B(n18773), .Z(n18778) );
  NAND U19360 ( .A(n18776), .B(n18775), .Z(n18777) );
  AND U19361 ( .A(n18778), .B(n18777), .Z(n18853) );
  NANDN U19362 ( .A(n18779), .B(n18780), .Z(n18785) );
  NOR U19363 ( .A(n18781), .B(n18780), .Z(n18783) );
  OR U19364 ( .A(n18783), .B(n18782), .Z(n18784) );
  AND U19365 ( .A(n18785), .B(n18784), .Z(n18852) );
  NAND U19366 ( .A(n18787), .B(n18786), .Z(n18791) );
  NAND U19367 ( .A(n18789), .B(n18788), .Z(n18790) );
  NAND U19368 ( .A(n18791), .B(n18790), .Z(n18849) );
  NAND U19369 ( .A(n18793), .B(n18792), .Z(n18797) );
  NAND U19370 ( .A(n18795), .B(n18794), .Z(n18796) );
  NAND U19371 ( .A(n18797), .B(n18796), .Z(n18856) );
  NAND U19372 ( .A(n18799), .B(n18798), .Z(n18803) );
  NAND U19373 ( .A(n18801), .B(n18800), .Z(n18802) );
  NAND U19374 ( .A(n18803), .B(n18802), .Z(n18863) );
  AND U19375 ( .A(y[1994]), .B(x[232]), .Z(n20066) );
  AND U19376 ( .A(x[226]), .B(y[1988]), .Z(n18941) );
  NAND U19377 ( .A(n20066), .B(n18941), .Z(n18807) );
  NANDN U19378 ( .A(n18805), .B(n18804), .Z(n18806) );
  NAND U19379 ( .A(n18807), .B(n18806), .Z(n18887) );
  AND U19380 ( .A(n18808), .B(o[204]), .Z(n18881) );
  AND U19381 ( .A(y[1996]), .B(x[225]), .Z(n18809) );
  XOR U19382 ( .A(n18810), .B(n18809), .Z(n18880) );
  XOR U19383 ( .A(n18881), .B(n18880), .Z(n18886) );
  AND U19384 ( .A(x[230]), .B(y[1991]), .Z(n19850) );
  AND U19385 ( .A(y[1995]), .B(x[226]), .Z(n18812) );
  NAND U19386 ( .A(y[1988]), .B(x[233]), .Z(n18811) );
  XNOR U19387 ( .A(n18812), .B(n18811), .Z(n18890) );
  XOR U19388 ( .A(n19850), .B(n18890), .Z(n18885) );
  XOR U19389 ( .A(n18886), .B(n18885), .Z(n18888) );
  XOR U19390 ( .A(n18887), .B(n18888), .Z(n18862) );
  NAND U19391 ( .A(n18814), .B(n18813), .Z(n18818) );
  ANDN U19392 ( .B(n18816), .A(n18815), .Z(n18817) );
  ANDN U19393 ( .B(n18818), .A(n18817), .Z(n18861) );
  XOR U19394 ( .A(n18862), .B(n18861), .Z(n18864) );
  XOR U19395 ( .A(n18863), .B(n18864), .Z(n18855) );
  XOR U19396 ( .A(n18856), .B(n18855), .Z(n18858) );
  NAND U19397 ( .A(n18820), .B(n18819), .Z(n18824) );
  NAND U19398 ( .A(n18822), .B(n18821), .Z(n18823) );
  NAND U19399 ( .A(n18824), .B(n18823), .Z(n18869) );
  AND U19400 ( .A(x[230]), .B(y[1995]), .Z(n19125) );
  IV U19401 ( .A(n19125), .Z(n19245) );
  AND U19402 ( .A(x[225]), .B(y[1990]), .Z(n18879) );
  AND U19403 ( .A(x[236]), .B(y[1996]), .Z(n20072) );
  AND U19404 ( .A(x[234]), .B(y[1987]), .Z(n19709) );
  AND U19405 ( .A(y[1986]), .B(x[235]), .Z(n19670) );
  AND U19406 ( .A(y[1989]), .B(x[232]), .Z(n18829) );
  XOR U19407 ( .A(n19670), .B(n18829), .Z(n18878) );
  XOR U19408 ( .A(n19709), .B(n18878), .Z(n18874) );
  XOR U19409 ( .A(n18873), .B(n18874), .Z(n18876) );
  XOR U19410 ( .A(n18875), .B(n18876), .Z(n18867) );
  AND U19411 ( .A(x[234]), .B(y[1992]), .Z(n18831) );
  AND U19412 ( .A(x[228]), .B(y[1986]), .Z(n18830) );
  NAND U19413 ( .A(n18831), .B(n18830), .Z(n18834) );
  NAND U19414 ( .A(n19414), .B(n18832), .Z(n18833) );
  NAND U19415 ( .A(n18834), .B(n18833), .Z(n18906) );
  AND U19416 ( .A(y[1984]), .B(x[237]), .Z(n18836) );
  NAND U19417 ( .A(y[1997]), .B(x[224]), .Z(n18835) );
  XNOR U19418 ( .A(n18836), .B(n18835), .Z(n18901) );
  AND U19419 ( .A(x[236]), .B(y[1985]), .Z(n18895) );
  XOR U19420 ( .A(n18895), .B(o[205]), .Z(n18900) );
  XOR U19421 ( .A(n18901), .B(n18900), .Z(n18905) );
  AND U19422 ( .A(y[1992]), .B(x[229]), .Z(n18838) );
  NAND U19423 ( .A(y[1994]), .B(x[227]), .Z(n18837) );
  XNOR U19424 ( .A(n18838), .B(n18837), .Z(n18899) );
  AND U19425 ( .A(x[228]), .B(y[1993]), .Z(n18898) );
  XOR U19426 ( .A(n18899), .B(n18898), .Z(n18904) );
  XOR U19427 ( .A(n18905), .B(n18904), .Z(n18907) );
  XOR U19428 ( .A(n18906), .B(n18907), .Z(n18868) );
  XOR U19429 ( .A(n18867), .B(n18868), .Z(n18870) );
  XOR U19430 ( .A(n18869), .B(n18870), .Z(n18857) );
  XNOR U19431 ( .A(n18858), .B(n18857), .Z(n18847) );
  NAND U19432 ( .A(n18840), .B(n18839), .Z(n18844) );
  NAND U19433 ( .A(n18842), .B(n18841), .Z(n18843) );
  AND U19434 ( .A(n18844), .B(n18843), .Z(n18846) );
  XOR U19435 ( .A(n18847), .B(n18846), .Z(n18848) );
  XOR U19436 ( .A(n18849), .B(n18848), .Z(n18854) );
  XNOR U19437 ( .A(n18852), .B(n18854), .Z(n18845) );
  XOR U19438 ( .A(n18853), .B(n18845), .Z(N430) );
  NAND U19439 ( .A(n18847), .B(n18846), .Z(n18851) );
  NAND U19440 ( .A(n18849), .B(n18848), .Z(n18850) );
  NAND U19441 ( .A(n18851), .B(n18850), .Z(n18986) );
  IV U19442 ( .A(n18986), .Z(n18984) );
  NAND U19443 ( .A(n18856), .B(n18855), .Z(n18860) );
  NAND U19444 ( .A(n18858), .B(n18857), .Z(n18859) );
  NAND U19445 ( .A(n18860), .B(n18859), .Z(n18979) );
  NAND U19446 ( .A(n18862), .B(n18861), .Z(n18866) );
  NAND U19447 ( .A(n18864), .B(n18863), .Z(n18865) );
  NAND U19448 ( .A(n18866), .B(n18865), .Z(n18978) );
  XOR U19449 ( .A(n18979), .B(n18978), .Z(n18981) );
  NAND U19450 ( .A(n18868), .B(n18867), .Z(n18872) );
  NAND U19451 ( .A(n18870), .B(n18869), .Z(n18871) );
  NAND U19452 ( .A(n18872), .B(n18871), .Z(n18913) );
  AND U19453 ( .A(x[235]), .B(y[1989]), .Z(n19043) );
  NAND U19454 ( .A(x[231]), .B(y[1996]), .Z(n19429) );
  XOR U19455 ( .A(n18968), .B(n18969), .Z(n18971) );
  AND U19456 ( .A(x[228]), .B(y[1994]), .Z(n19341) );
  AND U19457 ( .A(y[1995]), .B(x[227]), .Z(n18883) );
  NAND U19458 ( .A(y[1990]), .B(x[232]), .Z(n18882) );
  XNOR U19459 ( .A(n18883), .B(n18882), .Z(n18956) );
  XOR U19460 ( .A(n19243), .B(n18956), .Z(n18965) );
  XOR U19461 ( .A(n19341), .B(n18965), .Z(n18967) );
  AND U19462 ( .A(x[233]), .B(y[1989]), .Z(n19529) );
  AND U19463 ( .A(y[1996]), .B(x[226]), .Z(n18884) );
  AND U19464 ( .A(y[1988]), .B(x[234]), .Z(n19559) );
  XOR U19465 ( .A(n18884), .B(n19559), .Z(n18942) );
  XOR U19466 ( .A(n19529), .B(n18942), .Z(n18966) );
  XOR U19467 ( .A(n18967), .B(n18966), .Z(n18970) );
  XOR U19468 ( .A(n18971), .B(n18970), .Z(n18918) );
  XOR U19469 ( .A(n18918), .B(n18917), .Z(n18920) );
  XOR U19470 ( .A(n18919), .B(n18920), .Z(n18912) );
  AND U19471 ( .A(x[233]), .B(y[1995]), .Z(n18889) );
  NAND U19472 ( .A(n18889), .B(n18941), .Z(n18892) );
  NAND U19473 ( .A(n19850), .B(n18890), .Z(n18891) );
  NAND U19474 ( .A(n18892), .B(n18891), .Z(n18929) );
  AND U19475 ( .A(y[1984]), .B(x[238]), .Z(n18894) );
  NAND U19476 ( .A(y[1998]), .B(x[224]), .Z(n18893) );
  XNOR U19477 ( .A(n18894), .B(n18893), .Z(n18950) );
  NAND U19478 ( .A(n18895), .B(o[205]), .Z(n18951) );
  XNOR U19479 ( .A(n18950), .B(n18951), .Z(n18928) );
  NAND U19480 ( .A(y[1986]), .B(x[236]), .Z(n18896) );
  XNOR U19481 ( .A(n18897), .B(n18896), .Z(n18933) );
  AND U19482 ( .A(x[237]), .B(y[1985]), .Z(n18940) );
  XOR U19483 ( .A(o[206]), .B(n18940), .Z(n18932) );
  XOR U19484 ( .A(n18933), .B(n18932), .Z(n18927) );
  XOR U19485 ( .A(n18928), .B(n18927), .Z(n18930) );
  XNOR U19486 ( .A(n18929), .B(n18930), .Z(n18973) );
  AND U19487 ( .A(x[229]), .B(y[1994]), .Z(n19030) );
  AND U19488 ( .A(x[237]), .B(y[1997]), .Z(n20453) );
  NAND U19489 ( .A(y[1987]), .B(x[235]), .Z(n18902) );
  XNOR U19490 ( .A(n18903), .B(n18902), .Z(n18947) );
  AND U19491 ( .A(x[225]), .B(y[1997]), .Z(n18946) );
  XOR U19492 ( .A(n18947), .B(n18946), .Z(n18923) );
  XNOR U19493 ( .A(n18924), .B(n18923), .Z(n18926) );
  XOR U19494 ( .A(n18925), .B(n18926), .Z(n18972) );
  XOR U19495 ( .A(n18973), .B(n18972), .Z(n18975) );
  NAND U19496 ( .A(n18905), .B(n18904), .Z(n18909) );
  NAND U19497 ( .A(n18907), .B(n18906), .Z(n18908) );
  AND U19498 ( .A(n18909), .B(n18908), .Z(n18974) );
  XNOR U19499 ( .A(n18975), .B(n18974), .Z(n18911) );
  XOR U19500 ( .A(n18912), .B(n18911), .Z(n18914) );
  XOR U19501 ( .A(n18913), .B(n18914), .Z(n18980) );
  XOR U19502 ( .A(n18981), .B(n18980), .Z(n18987) );
  XNOR U19503 ( .A(n18985), .B(n18987), .Z(n18910) );
  XOR U19504 ( .A(n18984), .B(n18910), .Z(N431) );
  NAND U19505 ( .A(n18912), .B(n18911), .Z(n18916) );
  NAND U19506 ( .A(n18914), .B(n18913), .Z(n18915) );
  NAND U19507 ( .A(n18916), .B(n18915), .Z(n19077) );
  NANDN U19508 ( .A(n18918), .B(n18917), .Z(n18922) );
  NANDN U19509 ( .A(n18920), .B(n18919), .Z(n18921) );
  NAND U19510 ( .A(n18922), .B(n18921), .Z(n19052) );
  NAND U19511 ( .A(x[236]), .B(y[1991]), .Z(n19421) );
  NANDN U19512 ( .A(n19421), .B(n18931), .Z(n18935) );
  NAND U19513 ( .A(n18933), .B(n18932), .Z(n18934) );
  AND U19514 ( .A(n18935), .B(n18934), .Z(n18995) );
  AND U19515 ( .A(y[1988]), .B(x[235]), .Z(n18937) );
  NAND U19516 ( .A(y[1986]), .B(x[237]), .Z(n18936) );
  XNOR U19517 ( .A(n18937), .B(n18936), .Z(n18999) );
  AND U19518 ( .A(x[236]), .B(y[1987]), .Z(n18998) );
  XNOR U19519 ( .A(n18999), .B(n18998), .Z(n18993) );
  AND U19520 ( .A(y[1984]), .B(x[239]), .Z(n18939) );
  NAND U19521 ( .A(y[1999]), .B(x[224]), .Z(n18938) );
  XNOR U19522 ( .A(n18939), .B(n18938), .Z(n19019) );
  AND U19523 ( .A(o[206]), .B(n18940), .Z(n19018) );
  XNOR U19524 ( .A(n19019), .B(n19018), .Z(n18992) );
  XOR U19525 ( .A(n18993), .B(n18992), .Z(n18994) );
  XOR U19526 ( .A(n18995), .B(n18994), .Z(n19063) );
  NAND U19527 ( .A(x[234]), .B(y[1996]), .Z(n19852) );
  NANDN U19528 ( .A(n19852), .B(n18941), .Z(n18944) );
  NAND U19529 ( .A(n19529), .B(n18942), .Z(n18943) );
  NAND U19530 ( .A(n18944), .B(n18943), .Z(n19061) );
  AND U19531 ( .A(x[235]), .B(y[1992]), .Z(n19340) );
  NAND U19532 ( .A(n19340), .B(n18945), .Z(n18949) );
  NAND U19533 ( .A(n18947), .B(n18946), .Z(n18948) );
  NAND U19534 ( .A(n18949), .B(n18948), .Z(n19060) );
  XOR U19535 ( .A(n19061), .B(n19060), .Z(n19062) );
  XOR U19536 ( .A(n19054), .B(n19055), .Z(n19057) );
  XOR U19537 ( .A(n19056), .B(n19057), .Z(n19051) );
  AND U19538 ( .A(x[238]), .B(y[1998]), .Z(n20695) );
  NAND U19539 ( .A(n20695), .B(n19017), .Z(n18953) );
  NANDN U19540 ( .A(n18951), .B(n18950), .Z(n18952) );
  NAND U19541 ( .A(n18953), .B(n18952), .Z(n19045) );
  AND U19542 ( .A(x[232]), .B(y[1995]), .Z(n18954) );
  NANDN U19543 ( .A(n18955), .B(n18954), .Z(n18958) );
  NAND U19544 ( .A(n19243), .B(n18956), .Z(n18957) );
  NAND U19545 ( .A(n18958), .B(n18957), .Z(n19044) );
  XOR U19546 ( .A(n19045), .B(n19044), .Z(n19047) );
  AND U19547 ( .A(y[1989]), .B(x[234]), .Z(n18960) );
  NAND U19548 ( .A(y[1995]), .B(x[228]), .Z(n18959) );
  XNOR U19549 ( .A(n18960), .B(n18959), .Z(n19025) );
  AND U19550 ( .A(x[231]), .B(y[1992]), .Z(n19024) );
  XNOR U19551 ( .A(n19025), .B(n19024), .Z(n19032) );
  NAND U19552 ( .A(x[230]), .B(y[1993]), .Z(n19156) );
  XNOR U19553 ( .A(n19156), .B(n19030), .Z(n19031) );
  XNOR U19554 ( .A(n19032), .B(n19031), .Z(n19008) );
  AND U19555 ( .A(y[1997]), .B(x[226]), .Z(n18962) );
  NAND U19556 ( .A(y[1990]), .B(x[233]), .Z(n18961) );
  XNOR U19557 ( .A(n18962), .B(n18961), .Z(n19035) );
  AND U19558 ( .A(x[227]), .B(y[1996]), .Z(n19036) );
  XOR U19559 ( .A(n19035), .B(n19036), .Z(n19007) );
  AND U19560 ( .A(y[1998]), .B(x[225]), .Z(n18964) );
  NAND U19561 ( .A(y[1991]), .B(x[232]), .Z(n18963) );
  XNOR U19562 ( .A(n18964), .B(n18963), .Z(n19014) );
  AND U19563 ( .A(x[238]), .B(y[1985]), .Z(n19041) );
  XOR U19564 ( .A(o[207]), .B(n19041), .Z(n19013) );
  XOR U19565 ( .A(n19014), .B(n19013), .Z(n19006) );
  XOR U19566 ( .A(n19007), .B(n19006), .Z(n19009) );
  XOR U19567 ( .A(n19008), .B(n19009), .Z(n19046) );
  XOR U19568 ( .A(n19047), .B(n19046), .Z(n19067) );
  XOR U19569 ( .A(n19069), .B(n19068), .Z(n19050) );
  XNOR U19570 ( .A(n19051), .B(n19050), .Z(n19053) );
  XNOR U19571 ( .A(n19052), .B(n19053), .Z(n19076) );
  NAND U19572 ( .A(n18973), .B(n18972), .Z(n18977) );
  NAND U19573 ( .A(n18975), .B(n18974), .Z(n18976) );
  AND U19574 ( .A(n18977), .B(n18976), .Z(n19075) );
  XNOR U19575 ( .A(n19076), .B(n19075), .Z(n19078) );
  XOR U19576 ( .A(n19077), .B(n19078), .Z(n19074) );
  NAND U19577 ( .A(n18979), .B(n18978), .Z(n18983) );
  NAND U19578 ( .A(n18981), .B(n18980), .Z(n18982) );
  NAND U19579 ( .A(n18983), .B(n18982), .Z(n19073) );
  NANDN U19580 ( .A(n18984), .B(n18985), .Z(n18990) );
  NOR U19581 ( .A(n18986), .B(n18985), .Z(n18988) );
  OR U19582 ( .A(n18988), .B(n18987), .Z(n18989) );
  AND U19583 ( .A(n18990), .B(n18989), .Z(n19072) );
  XOR U19584 ( .A(n19073), .B(n19072), .Z(n18991) );
  XNOR U19585 ( .A(n19074), .B(n18991), .Z(N432) );
  NAND U19586 ( .A(n18993), .B(n18992), .Z(n18997) );
  NAND U19587 ( .A(n18995), .B(n18994), .Z(n18996) );
  NAND U19588 ( .A(n18997), .B(n18996), .Z(n19131) );
  AND U19589 ( .A(x[237]), .B(y[1988]), .Z(n19127) );
  NAND U19590 ( .A(n19670), .B(n19127), .Z(n19001) );
  NAND U19591 ( .A(n18999), .B(n18998), .Z(n19000) );
  NAND U19592 ( .A(n19001), .B(n19000), .Z(n19112) );
  AND U19593 ( .A(y[1998]), .B(x[226]), .Z(n19003) );
  NAND U19594 ( .A(y[1991]), .B(x[233]), .Z(n19002) );
  XNOR U19595 ( .A(n19003), .B(n19002), .Z(n19120) );
  AND U19596 ( .A(x[227]), .B(y[1997]), .Z(n19121) );
  XOR U19597 ( .A(n19120), .B(n19121), .Z(n19110) );
  AND U19598 ( .A(x[236]), .B(y[1988]), .Z(n19821) );
  AND U19599 ( .A(y[1995]), .B(x[229]), .Z(n19005) );
  NAND U19600 ( .A(y[1987]), .B(x[237]), .Z(n19004) );
  XNOR U19601 ( .A(n19005), .B(n19004), .Z(n19147) );
  XOR U19602 ( .A(n19821), .B(n19147), .Z(n19109) );
  XOR U19603 ( .A(n19110), .B(n19109), .Z(n19111) );
  XNOR U19604 ( .A(n19112), .B(n19111), .Z(n19128) );
  NAND U19605 ( .A(n19007), .B(n19006), .Z(n19011) );
  NAND U19606 ( .A(n19009), .B(n19008), .Z(n19010) );
  AND U19607 ( .A(n19011), .B(n19010), .Z(n19129) );
  XOR U19608 ( .A(n19128), .B(n19129), .Z(n19130) );
  XOR U19609 ( .A(n19131), .B(n19130), .Z(n19100) );
  AND U19610 ( .A(x[232]), .B(y[1998]), .Z(n19342) );
  NAND U19611 ( .A(n19342), .B(n19012), .Z(n19016) );
  NAND U19612 ( .A(n19014), .B(n19013), .Z(n19015) );
  NAND U19613 ( .A(n19016), .B(n19015), .Z(n19104) );
  AND U19614 ( .A(x[239]), .B(y[1999]), .Z(n21055) );
  NAND U19615 ( .A(n21055), .B(n19017), .Z(n19021) );
  NAND U19616 ( .A(n19019), .B(n19018), .Z(n19020) );
  NAND U19617 ( .A(n19021), .B(n19020), .Z(n19103) );
  XOR U19618 ( .A(n19104), .B(n19103), .Z(n19106) );
  AND U19619 ( .A(x[234]), .B(y[1995]), .Z(n19023) );
  NAND U19620 ( .A(n19023), .B(n19022), .Z(n19027) );
  NAND U19621 ( .A(n19025), .B(n19024), .Z(n19026) );
  NAND U19622 ( .A(n19027), .B(n19026), .Z(n19142) );
  AND U19623 ( .A(x[224]), .B(y[2000]), .Z(n19165) );
  AND U19624 ( .A(x[240]), .B(y[1984]), .Z(n19166) );
  XOR U19625 ( .A(n19165), .B(n19166), .Z(n19168) );
  NAND U19626 ( .A(x[239]), .B(y[1985]), .Z(n19152) );
  XOR U19627 ( .A(n19168), .B(n19167), .Z(n19141) );
  NAND U19628 ( .A(y[1993]), .B(x[231]), .Z(n19028) );
  XNOR U19629 ( .A(n19029), .B(n19028), .Z(n19158) );
  AND U19630 ( .A(x[234]), .B(y[1990]), .Z(n19157) );
  XOR U19631 ( .A(n19158), .B(n19157), .Z(n19140) );
  XOR U19632 ( .A(n19141), .B(n19140), .Z(n19143) );
  XOR U19633 ( .A(n19142), .B(n19143), .Z(n19105) );
  XNOR U19634 ( .A(n19106), .B(n19105), .Z(n19137) );
  NANDN U19635 ( .A(n19030), .B(n19156), .Z(n19034) );
  NAND U19636 ( .A(n19032), .B(n19031), .Z(n19033) );
  NAND U19637 ( .A(n19034), .B(n19033), .Z(n19135) );
  NAND U19638 ( .A(x[233]), .B(y[1997]), .Z(n19833) );
  NANDN U19639 ( .A(n19833), .B(n19419), .Z(n19038) );
  NAND U19640 ( .A(n19036), .B(n19035), .Z(n19037) );
  AND U19641 ( .A(n19038), .B(n19037), .Z(n19176) );
  AND U19642 ( .A(y[1999]), .B(x[225]), .Z(n19040) );
  NAND U19643 ( .A(y[1992]), .B(x[232]), .Z(n19039) );
  XNOR U19644 ( .A(n19040), .B(n19039), .Z(n19162) );
  AND U19645 ( .A(o[207]), .B(n19041), .Z(n19161) );
  XOR U19646 ( .A(n19162), .B(n19161), .Z(n19174) );
  NAND U19647 ( .A(y[1986]), .B(x[238]), .Z(n19042) );
  XNOR U19648 ( .A(n19043), .B(n19042), .Z(n19115) );
  AND U19649 ( .A(x[228]), .B(y[1996]), .Z(n19116) );
  XOR U19650 ( .A(n19115), .B(n19116), .Z(n19173) );
  XOR U19651 ( .A(n19174), .B(n19173), .Z(n19175) );
  XOR U19652 ( .A(n19176), .B(n19175), .Z(n19134) );
  XOR U19653 ( .A(n19135), .B(n19134), .Z(n19136) );
  XOR U19654 ( .A(n19137), .B(n19136), .Z(n19097) );
  NAND U19655 ( .A(n19045), .B(n19044), .Z(n19049) );
  NAND U19656 ( .A(n19047), .B(n19046), .Z(n19048) );
  AND U19657 ( .A(n19049), .B(n19048), .Z(n19098) );
  XOR U19658 ( .A(n19097), .B(n19098), .Z(n19099) );
  XOR U19659 ( .A(n19100), .B(n19099), .Z(n19083) );
  XNOR U19660 ( .A(n19083), .B(n19082), .Z(n19085) );
  NAND U19661 ( .A(n19055), .B(n19054), .Z(n19059) );
  NAND U19662 ( .A(n19057), .B(n19056), .Z(n19058) );
  NAND U19663 ( .A(n19059), .B(n19058), .Z(n19093) );
  NAND U19664 ( .A(n19061), .B(n19060), .Z(n19065) );
  NANDN U19665 ( .A(n19063), .B(n19062), .Z(n19064) );
  NAND U19666 ( .A(n19065), .B(n19064), .Z(n19091) );
  NANDN U19667 ( .A(n19067), .B(n19066), .Z(n19071) );
  NAND U19668 ( .A(n19069), .B(n19068), .Z(n19070) );
  AND U19669 ( .A(n19071), .B(n19070), .Z(n19092) );
  XOR U19670 ( .A(n19091), .B(n19092), .Z(n19094) );
  XOR U19671 ( .A(n19093), .B(n19094), .Z(n19084) );
  XNOR U19672 ( .A(n19085), .B(n19084), .Z(n19090) );
  NAND U19673 ( .A(n19076), .B(n19075), .Z(n19080) );
  NANDN U19674 ( .A(n19078), .B(n19077), .Z(n19079) );
  NAND U19675 ( .A(n19080), .B(n19079), .Z(n19088) );
  XNOR U19676 ( .A(n19089), .B(n19088), .Z(n19081) );
  XNOR U19677 ( .A(n19090), .B(n19081), .Z(N433) );
  NANDN U19678 ( .A(n19083), .B(n19082), .Z(n19087) );
  NAND U19679 ( .A(n19085), .B(n19084), .Z(n19086) );
  AND U19680 ( .A(n19087), .B(n19086), .Z(n19187) );
  NAND U19681 ( .A(n19092), .B(n19091), .Z(n19096) );
  NAND U19682 ( .A(n19094), .B(n19093), .Z(n19095) );
  NAND U19683 ( .A(n19096), .B(n19095), .Z(n19182) );
  NAND U19684 ( .A(n19098), .B(n19097), .Z(n19102) );
  NAND U19685 ( .A(n19100), .B(n19099), .Z(n19101) );
  NAND U19686 ( .A(n19102), .B(n19101), .Z(n19192) );
  NAND U19687 ( .A(n19104), .B(n19103), .Z(n19108) );
  NAND U19688 ( .A(n19106), .B(n19105), .Z(n19107) );
  NAND U19689 ( .A(n19108), .B(n19107), .Z(n19274) );
  NAND U19690 ( .A(n19110), .B(n19109), .Z(n19114) );
  NAND U19691 ( .A(n19112), .B(n19111), .Z(n19113) );
  NAND U19692 ( .A(n19114), .B(n19113), .Z(n19272) );
  NAND U19693 ( .A(x[238]), .B(y[1989]), .Z(n19465) );
  NANDN U19694 ( .A(n19465), .B(n19670), .Z(n19118) );
  NAND U19695 ( .A(n19116), .B(n19115), .Z(n19117) );
  NAND U19696 ( .A(n19118), .B(n19117), .Z(n19266) );
  AND U19697 ( .A(x[233]), .B(y[1998]), .Z(n20061) );
  NANDN U19698 ( .A(n19119), .B(n20061), .Z(n19123) );
  NAND U19699 ( .A(n19121), .B(n19120), .Z(n19122) );
  NAND U19700 ( .A(n19123), .B(n19122), .Z(n19265) );
  XOR U19701 ( .A(n19266), .B(n19265), .Z(n19268) );
  AND U19702 ( .A(x[229]), .B(y[1996]), .Z(n19302) );
  NAND U19703 ( .A(y[1993]), .B(x[232]), .Z(n19124) );
  XNOR U19704 ( .A(n19302), .B(n19124), .Z(n19244) );
  XOR U19705 ( .A(n19244), .B(n19125), .Z(n19259) );
  NAND U19706 ( .A(x[231]), .B(y[1994]), .Z(n19260) );
  IV U19707 ( .A(n19260), .Z(n19155) );
  XOR U19708 ( .A(n19259), .B(n19155), .Z(n19262) );
  NAND U19709 ( .A(y[1997]), .B(x[228]), .Z(n19126) );
  XNOR U19710 ( .A(n19127), .B(n19126), .Z(n19206) );
  AND U19711 ( .A(x[235]), .B(y[1990]), .Z(n19207) );
  XOR U19712 ( .A(n19206), .B(n19207), .Z(n19261) );
  XOR U19713 ( .A(n19262), .B(n19261), .Z(n19267) );
  XOR U19714 ( .A(n19268), .B(n19267), .Z(n19271) );
  XOR U19715 ( .A(n19272), .B(n19271), .Z(n19273) );
  XNOR U19716 ( .A(n19274), .B(n19273), .Z(n19190) );
  NAND U19717 ( .A(n19129), .B(n19128), .Z(n19133) );
  NAND U19718 ( .A(n19131), .B(n19130), .Z(n19132) );
  NAND U19719 ( .A(n19133), .B(n19132), .Z(n19189) );
  XOR U19720 ( .A(n19190), .B(n19189), .Z(n19191) );
  XOR U19721 ( .A(n19192), .B(n19191), .Z(n19181) );
  NAND U19722 ( .A(n19135), .B(n19134), .Z(n19139) );
  NAND U19723 ( .A(n19137), .B(n19136), .Z(n19138) );
  AND U19724 ( .A(n19139), .B(n19138), .Z(n19198) );
  NAND U19725 ( .A(n19141), .B(n19140), .Z(n19145) );
  NAND U19726 ( .A(n19143), .B(n19142), .Z(n19144) );
  NAND U19727 ( .A(n19145), .B(n19144), .Z(n19280) );
  AND U19728 ( .A(x[237]), .B(y[1995]), .Z(n20080) );
  NAND U19729 ( .A(n20080), .B(n19146), .Z(n19149) );
  NAND U19730 ( .A(n19147), .B(n19821), .Z(n19148) );
  NAND U19731 ( .A(n19149), .B(n19148), .Z(n19228) );
  AND U19732 ( .A(y[2000]), .B(x[225]), .Z(n19151) );
  NAND U19733 ( .A(y[1992]), .B(x[233]), .Z(n19150) );
  XNOR U19734 ( .A(n19151), .B(n19150), .Z(n19249) );
  ANDN U19735 ( .B(o[208]), .A(n19152), .Z(n19248) );
  XOR U19736 ( .A(n19249), .B(n19248), .Z(n19226) );
  AND U19737 ( .A(y[1986]), .B(x[239]), .Z(n19154) );
  NAND U19738 ( .A(y[1989]), .B(x[236]), .Z(n19153) );
  XNOR U19739 ( .A(n19154), .B(n19153), .Z(n19201) );
  NAND U19740 ( .A(x[238]), .B(y[1987]), .Z(n19202) );
  XOR U19741 ( .A(n19226), .B(n19225), .Z(n19227) );
  XOR U19742 ( .A(n19228), .B(n19227), .Z(n19278) );
  NANDN U19743 ( .A(n19156), .B(n19155), .Z(n19160) );
  NAND U19744 ( .A(n19158), .B(n19157), .Z(n19159) );
  NAND U19745 ( .A(n19160), .B(n19159), .Z(n19238) );
  NAND U19746 ( .A(x[232]), .B(y[1999]), .Z(n19920) );
  AND U19747 ( .A(x[225]), .B(y[1992]), .Z(n19320) );
  NANDN U19748 ( .A(n19920), .B(n19320), .Z(n19164) );
  NAND U19749 ( .A(n19162), .B(n19161), .Z(n19163) );
  NAND U19750 ( .A(n19164), .B(n19163), .Z(n19237) );
  XOR U19751 ( .A(n19238), .B(n19237), .Z(n19240) );
  NAND U19752 ( .A(n19166), .B(n19165), .Z(n19170) );
  NAND U19753 ( .A(n19168), .B(n19167), .Z(n19169) );
  NAND U19754 ( .A(n19170), .B(n19169), .Z(n19234) );
  AND U19755 ( .A(x[224]), .B(y[2001]), .Z(n19215) );
  NAND U19756 ( .A(x[241]), .B(y[1984]), .Z(n19216) );
  AND U19757 ( .A(x[240]), .B(y[1985]), .Z(n19212) );
  XOR U19758 ( .A(o[209]), .B(n19212), .Z(n19217) );
  XOR U19759 ( .A(n19218), .B(n19217), .Z(n19232) );
  AND U19760 ( .A(y[1999]), .B(x[226]), .Z(n19172) );
  NAND U19761 ( .A(y[1991]), .B(x[234]), .Z(n19171) );
  XNOR U19762 ( .A(n19172), .B(n19171), .Z(n19253) );
  NAND U19763 ( .A(x[227]), .B(y[1998]), .Z(n19254) );
  XOR U19764 ( .A(n19232), .B(n19231), .Z(n19233) );
  XOR U19765 ( .A(n19234), .B(n19233), .Z(n19239) );
  XOR U19766 ( .A(n19240), .B(n19239), .Z(n19277) );
  XOR U19767 ( .A(n19278), .B(n19277), .Z(n19279) );
  XNOR U19768 ( .A(n19280), .B(n19279), .Z(n19195) );
  NAND U19769 ( .A(n19174), .B(n19173), .Z(n19178) );
  NANDN U19770 ( .A(n19176), .B(n19175), .Z(n19177) );
  AND U19771 ( .A(n19178), .B(n19177), .Z(n19196) );
  XOR U19772 ( .A(n19195), .B(n19196), .Z(n19197) );
  XOR U19773 ( .A(n19198), .B(n19197), .Z(n19180) );
  XOR U19774 ( .A(n19182), .B(n19183), .Z(n19188) );
  XOR U19775 ( .A(n19186), .B(n19188), .Z(n19179) );
  XOR U19776 ( .A(n19187), .B(n19179), .Z(N434) );
  NANDN U19777 ( .A(n19181), .B(n19180), .Z(n19185) );
  NAND U19778 ( .A(n19183), .B(n19182), .Z(n19184) );
  AND U19779 ( .A(n19185), .B(n19184), .Z(n19392) );
  NAND U19780 ( .A(n19190), .B(n19189), .Z(n19194) );
  NAND U19781 ( .A(n19192), .B(n19191), .Z(n19193) );
  AND U19782 ( .A(n19194), .B(n19193), .Z(n19389) );
  NAND U19783 ( .A(n19196), .B(n19195), .Z(n19200) );
  NANDN U19784 ( .A(n19198), .B(n19197), .Z(n19199) );
  AND U19785 ( .A(n19200), .B(n19199), .Z(n19387) );
  AND U19786 ( .A(x[239]), .B(y[1989]), .Z(n19427) );
  AND U19787 ( .A(x[236]), .B(y[1986]), .Z(n19519) );
  NAND U19788 ( .A(n19427), .B(n19519), .Z(n19204) );
  NANDN U19789 ( .A(n19202), .B(n19201), .Z(n19203) );
  NAND U19790 ( .A(n19204), .B(n19203), .Z(n19369) );
  NAND U19791 ( .A(n20453), .B(n19205), .Z(n19209) );
  NAND U19792 ( .A(n19207), .B(n19206), .Z(n19208) );
  AND U19793 ( .A(n19209), .B(n19208), .Z(n19359) );
  AND U19794 ( .A(y[2001]), .B(x[225]), .Z(n19211) );
  NAND U19795 ( .A(y[1992]), .B(x[234]), .Z(n19210) );
  XNOR U19796 ( .A(n19211), .B(n19210), .Z(n19322) );
  AND U19797 ( .A(o[209]), .B(n19212), .Z(n19321) );
  XOR U19798 ( .A(n19322), .B(n19321), .Z(n19357) );
  AND U19799 ( .A(y[1987]), .B(x[239]), .Z(n19214) );
  NAND U19800 ( .A(y[1993]), .B(x[233]), .Z(n19213) );
  XNOR U19801 ( .A(n19214), .B(n19213), .Z(n19312) );
  AND U19802 ( .A(x[238]), .B(y[1988]), .Z(n19313) );
  XOR U19803 ( .A(n19312), .B(n19313), .Z(n19356) );
  XOR U19804 ( .A(n19357), .B(n19356), .Z(n19358) );
  XOR U19805 ( .A(n19369), .B(n19368), .Z(n19371) );
  NANDN U19806 ( .A(n19216), .B(n19215), .Z(n19220) );
  NAND U19807 ( .A(n19218), .B(n19217), .Z(n19219) );
  AND U19808 ( .A(n19220), .B(n19219), .Z(n19381) );
  AND U19809 ( .A(y[1986]), .B(x[240]), .Z(n19222) );
  NAND U19810 ( .A(y[1991]), .B(x[235]), .Z(n19221) );
  XNOR U19811 ( .A(n19222), .B(n19221), .Z(n19308) );
  NAND U19812 ( .A(x[226]), .B(y[2000]), .Z(n19309) );
  AND U19813 ( .A(y[1997]), .B(x[229]), .Z(n19447) );
  NAND U19814 ( .A(y[1996]), .B(x[230]), .Z(n19223) );
  XNOR U19815 ( .A(n19447), .B(n19223), .Z(n19305) );
  NAND U19816 ( .A(y[1998]), .B(x[228]), .Z(n19224) );
  XNOR U19817 ( .A(n20066), .B(n19224), .Z(n19343) );
  AND U19818 ( .A(x[231]), .B(y[1995]), .Z(n19344) );
  XOR U19819 ( .A(n19343), .B(n19344), .Z(n19304) );
  XOR U19820 ( .A(n19305), .B(n19304), .Z(n19382) );
  XOR U19821 ( .A(n19383), .B(n19382), .Z(n19370) );
  XNOR U19822 ( .A(n19371), .B(n19370), .Z(n19291) );
  NAND U19823 ( .A(n19226), .B(n19225), .Z(n19230) );
  NAND U19824 ( .A(n19228), .B(n19227), .Z(n19229) );
  AND U19825 ( .A(n19230), .B(n19229), .Z(n19362) );
  NAND U19826 ( .A(n19232), .B(n19231), .Z(n19236) );
  NAND U19827 ( .A(n19234), .B(n19233), .Z(n19235) );
  AND U19828 ( .A(n19236), .B(n19235), .Z(n19363) );
  XOR U19829 ( .A(n19362), .B(n19363), .Z(n19364) );
  NAND U19830 ( .A(n19238), .B(n19237), .Z(n19242) );
  NAND U19831 ( .A(n19240), .B(n19239), .Z(n19241) );
  AND U19832 ( .A(n19242), .B(n19241), .Z(n19365) );
  XOR U19833 ( .A(n19364), .B(n19365), .Z(n19290) );
  XOR U19834 ( .A(n19291), .B(n19290), .Z(n19293) );
  AND U19835 ( .A(x[232]), .B(y[1996]), .Z(n19565) );
  NAND U19836 ( .A(n19565), .B(n19243), .Z(n19247) );
  NANDN U19837 ( .A(n19245), .B(n19244), .Z(n19246) );
  NAND U19838 ( .A(n19247), .B(n19246), .Z(n19375) );
  AND U19839 ( .A(x[233]), .B(y[2000]), .Z(n20219) );
  IV U19840 ( .A(n20219), .Z(n20090) );
  NANDN U19841 ( .A(n20090), .B(n19320), .Z(n19251) );
  NAND U19842 ( .A(n19249), .B(n19248), .Z(n19250) );
  NAND U19843 ( .A(n19251), .B(n19250), .Z(n19374) );
  XOR U19844 ( .A(n19375), .B(n19374), .Z(n19377) );
  AND U19845 ( .A(x[234]), .B(y[1999]), .Z(n20089) );
  IV U19846 ( .A(n20089), .Z(n20218) );
  NANDN U19847 ( .A(n20218), .B(n19252), .Z(n19256) );
  NANDN U19848 ( .A(n19254), .B(n19253), .Z(n19255) );
  AND U19849 ( .A(n19256), .B(n19255), .Z(n19353) );
  AND U19850 ( .A(x[224]), .B(y[2002]), .Z(n19325) );
  AND U19851 ( .A(x[242]), .B(y[1984]), .Z(n19326) );
  XOR U19852 ( .A(n19325), .B(n19326), .Z(n19328) );
  AND U19853 ( .A(x[241]), .B(y[1985]), .Z(n19347) );
  XOR U19854 ( .A(o[210]), .B(n19347), .Z(n19327) );
  XOR U19855 ( .A(n19328), .B(n19327), .Z(n19351) );
  AND U19856 ( .A(y[1989]), .B(x[237]), .Z(n19258) );
  NAND U19857 ( .A(y[1999]), .B(x[227]), .Z(n19257) );
  XNOR U19858 ( .A(n19258), .B(n19257), .Z(n19333) );
  AND U19859 ( .A(x[236]), .B(y[1990]), .Z(n19334) );
  XOR U19860 ( .A(n19333), .B(n19334), .Z(n19350) );
  XOR U19861 ( .A(n19351), .B(n19350), .Z(n19352) );
  XNOR U19862 ( .A(n19377), .B(n19376), .Z(n19297) );
  NANDN U19863 ( .A(n19260), .B(n19259), .Z(n19264) );
  NAND U19864 ( .A(n19262), .B(n19261), .Z(n19263) );
  AND U19865 ( .A(n19264), .B(n19263), .Z(n19296) );
  XOR U19866 ( .A(n19297), .B(n19296), .Z(n19298) );
  NAND U19867 ( .A(n19266), .B(n19265), .Z(n19270) );
  NAND U19868 ( .A(n19268), .B(n19267), .Z(n19269) );
  AND U19869 ( .A(n19270), .B(n19269), .Z(n19299) );
  XOR U19870 ( .A(n19298), .B(n19299), .Z(n19292) );
  XNOR U19871 ( .A(n19293), .B(n19292), .Z(n19287) );
  NAND U19872 ( .A(n19272), .B(n19271), .Z(n19276) );
  NAND U19873 ( .A(n19274), .B(n19273), .Z(n19275) );
  NAND U19874 ( .A(n19276), .B(n19275), .Z(n19285) );
  NAND U19875 ( .A(n19278), .B(n19277), .Z(n19282) );
  NAND U19876 ( .A(n19280), .B(n19279), .Z(n19281) );
  NAND U19877 ( .A(n19282), .B(n19281), .Z(n19284) );
  XOR U19878 ( .A(n19285), .B(n19284), .Z(n19286) );
  XOR U19879 ( .A(n19287), .B(n19286), .Z(n19386) );
  XOR U19880 ( .A(n19387), .B(n19386), .Z(n19388) );
  XOR U19881 ( .A(n19389), .B(n19388), .Z(n19394) );
  XNOR U19882 ( .A(n19393), .B(n19394), .Z(n19283) );
  XOR U19883 ( .A(n19392), .B(n19283), .Z(N435) );
  NAND U19884 ( .A(n19285), .B(n19284), .Z(n19289) );
  NAND U19885 ( .A(n19287), .B(n19286), .Z(n19288) );
  AND U19886 ( .A(n19289), .B(n19288), .Z(n19509) );
  NAND U19887 ( .A(n19291), .B(n19290), .Z(n19295) );
  NAND U19888 ( .A(n19293), .B(n19292), .Z(n19294) );
  AND U19889 ( .A(n19295), .B(n19294), .Z(n19507) );
  NAND U19890 ( .A(n19297), .B(n19296), .Z(n19301) );
  NAND U19891 ( .A(n19299), .B(n19298), .Z(n19300) );
  AND U19892 ( .A(n19301), .B(n19300), .Z(n19399) );
  AND U19893 ( .A(x[230]), .B(y[1997]), .Z(n19303) );
  NAND U19894 ( .A(n19303), .B(n19302), .Z(n19307) );
  NAND U19895 ( .A(n19305), .B(n19304), .Z(n19306) );
  AND U19896 ( .A(n19307), .B(n19306), .Z(n19488) );
  AND U19897 ( .A(x[240]), .B(y[1991]), .Z(n19837) );
  NAND U19898 ( .A(n19837), .B(n19670), .Z(n19311) );
  NANDN U19899 ( .A(n19309), .B(n19308), .Z(n19310) );
  AND U19900 ( .A(n19311), .B(n19310), .Z(n19486) );
  AND U19901 ( .A(x[239]), .B(y[1993]), .Z(n20093) );
  NAND U19902 ( .A(n20093), .B(n19414), .Z(n19315) );
  NAND U19903 ( .A(n19313), .B(n19312), .Z(n19314) );
  NAND U19904 ( .A(n19315), .B(n19314), .Z(n19405) );
  AND U19905 ( .A(y[2002]), .B(x[225]), .Z(n19317) );
  NAND U19906 ( .A(y[1995]), .B(x[232]), .Z(n19316) );
  XNOR U19907 ( .A(n19317), .B(n19316), .Z(n19464) );
  AND U19908 ( .A(y[1990]), .B(x[237]), .Z(n19319) );
  NAND U19909 ( .A(y[2001]), .B(x[226]), .Z(n19318) );
  XNOR U19910 ( .A(n19319), .B(n19318), .Z(n19420) );
  XOR U19911 ( .A(n19403), .B(n19402), .Z(n19404) );
  XOR U19912 ( .A(n19405), .B(n19404), .Z(n19485) );
  AND U19913 ( .A(x[234]), .B(y[2001]), .Z(n20541) );
  IV U19914 ( .A(n20541), .Z(n20408) );
  NANDN U19915 ( .A(n20408), .B(n19320), .Z(n19324) );
  NAND U19916 ( .A(n19322), .B(n19321), .Z(n19323) );
  NAND U19917 ( .A(n19324), .B(n19323), .Z(n19444) );
  NAND U19918 ( .A(n19326), .B(n19325), .Z(n19330) );
  NAND U19919 ( .A(n19328), .B(n19327), .Z(n19329) );
  NAND U19920 ( .A(n19330), .B(n19329), .Z(n19442) );
  AND U19921 ( .A(y[1987]), .B(x[240]), .Z(n20146) );
  NAND U19922 ( .A(y[1994]), .B(x[233]), .Z(n19331) );
  XNOR U19923 ( .A(n20146), .B(n19331), .Z(n19415) );
  NAND U19924 ( .A(x[239]), .B(y[1988]), .Z(n19416) );
  XOR U19925 ( .A(n19442), .B(n19441), .Z(n19443) );
  XNOR U19926 ( .A(n19444), .B(n19443), .Z(n19481) );
  AND U19927 ( .A(x[237]), .B(y[1999]), .Z(n20714) );
  NAND U19928 ( .A(n19332), .B(n20714), .Z(n19336) );
  NAND U19929 ( .A(n19334), .B(n19333), .Z(n19335) );
  NAND U19930 ( .A(n19336), .B(n19335), .Z(n19438) );
  AND U19931 ( .A(y[1993]), .B(x[234]), .Z(n19338) );
  NAND U19932 ( .A(y[1986]), .B(x[241]), .Z(n19337) );
  XNOR U19933 ( .A(n19338), .B(n19337), .Z(n19470) );
  AND U19934 ( .A(x[242]), .B(y[1985]), .Z(n19434) );
  XOR U19935 ( .A(o[211]), .B(n19434), .Z(n19469) );
  XOR U19936 ( .A(n19470), .B(n19469), .Z(n19436) );
  NAND U19937 ( .A(y[2000]), .B(x[227]), .Z(n19339) );
  XNOR U19938 ( .A(n19340), .B(n19339), .Z(n19428) );
  XOR U19939 ( .A(n19436), .B(n19435), .Z(n19437) );
  XNOR U19940 ( .A(n19438), .B(n19437), .Z(n19480) );
  NAND U19941 ( .A(n19342), .B(n19341), .Z(n19346) );
  NAND U19942 ( .A(n19344), .B(n19343), .Z(n19345) );
  AND U19943 ( .A(n19346), .B(n19345), .Z(n19411) );
  AND U19944 ( .A(x[224]), .B(y[2003]), .Z(n19451) );
  AND U19945 ( .A(x[243]), .B(y[1984]), .Z(n19452) );
  XOR U19946 ( .A(n19451), .B(n19452), .Z(n19454) );
  AND U19947 ( .A(o[210]), .B(n19347), .Z(n19453) );
  XOR U19948 ( .A(n19454), .B(n19453), .Z(n19409) );
  AND U19949 ( .A(x[228]), .B(y[1999]), .Z(n19579) );
  AND U19950 ( .A(y[1998]), .B(x[229]), .Z(n19349) );
  NAND U19951 ( .A(y[1997]), .B(x[230]), .Z(n19348) );
  XNOR U19952 ( .A(n19349), .B(n19348), .Z(n19448) );
  XOR U19953 ( .A(n19579), .B(n19448), .Z(n19408) );
  XOR U19954 ( .A(n19409), .B(n19408), .Z(n19410) );
  XOR U19955 ( .A(n19411), .B(n19410), .Z(n19479) );
  XOR U19956 ( .A(n19480), .B(n19479), .Z(n19482) );
  XNOR U19957 ( .A(n19481), .B(n19482), .Z(n19475) );
  NAND U19958 ( .A(n19351), .B(n19350), .Z(n19355) );
  NANDN U19959 ( .A(n19353), .B(n19352), .Z(n19354) );
  AND U19960 ( .A(n19355), .B(n19354), .Z(n19474) );
  NAND U19961 ( .A(n19357), .B(n19356), .Z(n19361) );
  NANDN U19962 ( .A(n19359), .B(n19358), .Z(n19360) );
  NAND U19963 ( .A(n19361), .B(n19360), .Z(n19473) );
  XNOR U19964 ( .A(n19475), .B(n19476), .Z(n19396) );
  XOR U19965 ( .A(n19397), .B(n19396), .Z(n19398) );
  NAND U19966 ( .A(n19363), .B(n19362), .Z(n19367) );
  NAND U19967 ( .A(n19365), .B(n19364), .Z(n19366) );
  AND U19968 ( .A(n19367), .B(n19366), .Z(n19498) );
  NAND U19969 ( .A(n19369), .B(n19368), .Z(n19373) );
  NAND U19970 ( .A(n19371), .B(n19370), .Z(n19372) );
  AND U19971 ( .A(n19373), .B(n19372), .Z(n19494) );
  NAND U19972 ( .A(n19375), .B(n19374), .Z(n19379) );
  NAND U19973 ( .A(n19377), .B(n19376), .Z(n19378) );
  AND U19974 ( .A(n19379), .B(n19378), .Z(n19492) );
  NANDN U19975 ( .A(n19381), .B(n19380), .Z(n19385) );
  NAND U19976 ( .A(n19383), .B(n19382), .Z(n19384) );
  NAND U19977 ( .A(n19385), .B(n19384), .Z(n19491) );
  XOR U19978 ( .A(n19498), .B(n19497), .Z(n19500) );
  XOR U19979 ( .A(n19499), .B(n19500), .Z(n19506) );
  XOR U19980 ( .A(n19507), .B(n19506), .Z(n19508) );
  XOR U19981 ( .A(n19509), .B(n19508), .Z(n19505) );
  NAND U19982 ( .A(n19387), .B(n19386), .Z(n19391) );
  NAND U19983 ( .A(n19389), .B(n19388), .Z(n19390) );
  NAND U19984 ( .A(n19391), .B(n19390), .Z(n19504) );
  XOR U19985 ( .A(n19504), .B(n19503), .Z(n19395) );
  XNOR U19986 ( .A(n19505), .B(n19395), .Z(N436) );
  NAND U19987 ( .A(n19397), .B(n19396), .Z(n19401) );
  NANDN U19988 ( .A(n19399), .B(n19398), .Z(n19400) );
  AND U19989 ( .A(n19401), .B(n19400), .Z(n19617) );
  NAND U19990 ( .A(n19403), .B(n19402), .Z(n19407) );
  NAND U19991 ( .A(n19405), .B(n19404), .Z(n19406) );
  NAND U19992 ( .A(n19407), .B(n19406), .Z(n19514) );
  NAND U19993 ( .A(n19409), .B(n19408), .Z(n19413) );
  NANDN U19994 ( .A(n19411), .B(n19410), .Z(n19412) );
  NAND U19995 ( .A(n19413), .B(n19412), .Z(n19513) );
  XOR U19996 ( .A(n19514), .B(n19513), .Z(n19516) );
  AND U19997 ( .A(x[240]), .B(y[1994]), .Z(n20367) );
  NAND U19998 ( .A(n20367), .B(n19414), .Z(n19418) );
  NANDN U19999 ( .A(n19416), .B(n19415), .Z(n19417) );
  AND U20000 ( .A(n19418), .B(n19417), .Z(n19554) );
  AND U20001 ( .A(x[237]), .B(y[2001]), .Z(n20932) );
  NAND U20002 ( .A(n20932), .B(n19419), .Z(n19423) );
  NANDN U20003 ( .A(n19421), .B(n19420), .Z(n19422) );
  AND U20004 ( .A(n19423), .B(n19422), .Z(n19599) );
  AND U20005 ( .A(y[1988]), .B(x[240]), .Z(n19425) );
  NAND U20006 ( .A(y[1994]), .B(x[234]), .Z(n19424) );
  XNOR U20007 ( .A(n19425), .B(n19424), .Z(n19560) );
  AND U20008 ( .A(x[226]), .B(y[2002]), .Z(n19561) );
  XOR U20009 ( .A(n19560), .B(n19561), .Z(n19597) );
  NAND U20010 ( .A(y[1995]), .B(x[233]), .Z(n19426) );
  XNOR U20011 ( .A(n19427), .B(n19426), .Z(n19530) );
  AND U20012 ( .A(x[238]), .B(y[1990]), .Z(n19531) );
  XOR U20013 ( .A(n19530), .B(n19531), .Z(n19596) );
  XOR U20014 ( .A(n19597), .B(n19596), .Z(n19598) );
  NAND U20015 ( .A(x[235]), .B(y[2000]), .Z(n20542) );
  NANDN U20016 ( .A(n20542), .B(n19697), .Z(n19431) );
  NANDN U20017 ( .A(n19429), .B(n19428), .Z(n19430) );
  AND U20018 ( .A(n19431), .B(n19430), .Z(n19605) );
  AND U20019 ( .A(y[1993]), .B(x[235]), .Z(n19433) );
  NAND U20020 ( .A(y[2003]), .B(x[225]), .Z(n19432) );
  XNOR U20021 ( .A(n19433), .B(n19432), .Z(n19526) );
  AND U20022 ( .A(x[243]), .B(y[1985]), .Z(n19534) );
  XOR U20023 ( .A(o[212]), .B(n19534), .Z(n19525) );
  XOR U20024 ( .A(n19526), .B(n19525), .Z(n19603) );
  AND U20025 ( .A(x[224]), .B(y[2004]), .Z(n19584) );
  AND U20026 ( .A(x[244]), .B(y[1984]), .Z(n19585) );
  XOR U20027 ( .A(n19584), .B(n19585), .Z(n19587) );
  AND U20028 ( .A(o[211]), .B(n19434), .Z(n19586) );
  XOR U20029 ( .A(n19587), .B(n19586), .Z(n19602) );
  XOR U20030 ( .A(n19603), .B(n19602), .Z(n19604) );
  XOR U20031 ( .A(n19556), .B(n19555), .Z(n19515) );
  XNOR U20032 ( .A(n19516), .B(n19515), .Z(n19611) );
  NAND U20033 ( .A(n19436), .B(n19435), .Z(n19440) );
  NAND U20034 ( .A(n19438), .B(n19437), .Z(n19439) );
  AND U20035 ( .A(n19440), .B(n19439), .Z(n19609) );
  NAND U20036 ( .A(n19442), .B(n19441), .Z(n19446) );
  NAND U20037 ( .A(n19444), .B(n19443), .Z(n19445) );
  AND U20038 ( .A(n19446), .B(n19445), .Z(n19550) );
  NAND U20039 ( .A(x[230]), .B(y[1998]), .Z(n19536) );
  NANDN U20040 ( .A(n19536), .B(n19447), .Z(n19450) );
  NAND U20041 ( .A(n19448), .B(n19579), .Z(n19449) );
  NAND U20042 ( .A(n19450), .B(n19449), .Z(n19544) );
  NAND U20043 ( .A(n19452), .B(n19451), .Z(n19456) );
  NAND U20044 ( .A(n19454), .B(n19453), .Z(n19455) );
  NAND U20045 ( .A(n19456), .B(n19455), .Z(n19542) );
  AND U20046 ( .A(y[1986]), .B(x[242]), .Z(n19458) );
  NAND U20047 ( .A(y[1992]), .B(x[236]), .Z(n19457) );
  XNOR U20048 ( .A(n19458), .B(n19457), .Z(n19520) );
  AND U20049 ( .A(x[241]), .B(y[1987]), .Z(n19521) );
  XOR U20050 ( .A(n19520), .B(n19521), .Z(n19541) );
  XOR U20051 ( .A(n19542), .B(n19541), .Z(n19543) );
  XNOR U20052 ( .A(n19544), .B(n19543), .Z(n19548) );
  AND U20053 ( .A(y[1991]), .B(x[237]), .Z(n19460) );
  NAND U20054 ( .A(y[2001]), .B(x[227]), .Z(n19459) );
  XNOR U20055 ( .A(n19460), .B(n19459), .Z(n19566) );
  XNOR U20056 ( .A(n19566), .B(n19565), .Z(n19538) );
  AND U20057 ( .A(y[1999]), .B(x[229]), .Z(n19462) );
  NAND U20058 ( .A(y[2000]), .B(x[228]), .Z(n19461) );
  XNOR U20059 ( .A(n19462), .B(n19461), .Z(n19581) );
  AND U20060 ( .A(x[231]), .B(y[1997]), .Z(n19580) );
  XNOR U20061 ( .A(n19581), .B(n19580), .Z(n19535) );
  XOR U20062 ( .A(n19536), .B(n19535), .Z(n19537) );
  XNOR U20063 ( .A(n19538), .B(n19537), .Z(n19592) );
  AND U20064 ( .A(x[232]), .B(y[2002]), .Z(n20679) );
  NAND U20065 ( .A(n20679), .B(n19463), .Z(n19467) );
  NANDN U20066 ( .A(n19465), .B(n19464), .Z(n19466) );
  AND U20067 ( .A(n19467), .B(n19466), .Z(n19591) );
  AND U20068 ( .A(x[241]), .B(y[1993]), .Z(n20298) );
  IV U20069 ( .A(n20298), .Z(n20375) );
  NANDN U20070 ( .A(n20375), .B(n19468), .Z(n19472) );
  NAND U20071 ( .A(n19470), .B(n19469), .Z(n19471) );
  NAND U20072 ( .A(n19472), .B(n19471), .Z(n19590) );
  XNOR U20073 ( .A(n19592), .B(n19593), .Z(n19547) );
  XOR U20074 ( .A(n19548), .B(n19547), .Z(n19549) );
  XOR U20075 ( .A(n19550), .B(n19549), .Z(n19608) );
  XOR U20076 ( .A(n19609), .B(n19608), .Z(n19610) );
  XNOR U20077 ( .A(n19611), .B(n19610), .Z(n19615) );
  NANDN U20078 ( .A(n19474), .B(n19473), .Z(n19478) );
  NAND U20079 ( .A(n19476), .B(n19475), .Z(n19477) );
  AND U20080 ( .A(n19478), .B(n19477), .Z(n19623) );
  NAND U20081 ( .A(n19480), .B(n19479), .Z(n19484) );
  NAND U20082 ( .A(n19482), .B(n19481), .Z(n19483) );
  AND U20083 ( .A(n19484), .B(n19483), .Z(n19621) );
  NANDN U20084 ( .A(n19486), .B(n19485), .Z(n19490) );
  NANDN U20085 ( .A(n19488), .B(n19487), .Z(n19489) );
  AND U20086 ( .A(n19490), .B(n19489), .Z(n19620) );
  XNOR U20087 ( .A(n19623), .B(n19622), .Z(n19614) );
  XOR U20088 ( .A(n19615), .B(n19614), .Z(n19616) );
  XOR U20089 ( .A(n19617), .B(n19616), .Z(n19636) );
  NANDN U20090 ( .A(n19492), .B(n19491), .Z(n19496) );
  NANDN U20091 ( .A(n19494), .B(n19493), .Z(n19495) );
  AND U20092 ( .A(n19496), .B(n19495), .Z(n19633) );
  NAND U20093 ( .A(n19498), .B(n19497), .Z(n19502) );
  NAND U20094 ( .A(n19500), .B(n19499), .Z(n19501) );
  AND U20095 ( .A(n19502), .B(n19501), .Z(n19634) );
  XOR U20096 ( .A(n19633), .B(n19634), .Z(n19635) );
  XOR U20097 ( .A(n19636), .B(n19635), .Z(n19629) );
  NAND U20098 ( .A(n19507), .B(n19506), .Z(n19511) );
  NANDN U20099 ( .A(n19509), .B(n19508), .Z(n19510) );
  AND U20100 ( .A(n19511), .B(n19510), .Z(n19628) );
  IV U20101 ( .A(n19628), .Z(n19626) );
  XOR U20102 ( .A(n19627), .B(n19626), .Z(n19512) );
  XNOR U20103 ( .A(n19629), .B(n19512), .Z(N437) );
  NAND U20104 ( .A(n19514), .B(n19513), .Z(n19518) );
  NAND U20105 ( .A(n19516), .B(n19515), .Z(n19517) );
  NAND U20106 ( .A(n19518), .B(n19517), .Z(n19649) );
  AND U20107 ( .A(x[242]), .B(y[1992]), .Z(n20373) );
  NAND U20108 ( .A(n20373), .B(n19519), .Z(n19523) );
  NAND U20109 ( .A(n19521), .B(n19520), .Z(n19522) );
  NAND U20110 ( .A(n19523), .B(n19522), .Z(n19726) );
  AND U20111 ( .A(x[235]), .B(y[2003]), .Z(n20985) );
  AND U20112 ( .A(x[225]), .B(y[1993]), .Z(n19524) );
  NAND U20113 ( .A(n20985), .B(n19524), .Z(n19528) );
  NAND U20114 ( .A(n19526), .B(n19525), .Z(n19527) );
  NAND U20115 ( .A(n19528), .B(n19527), .Z(n19725) );
  XOR U20116 ( .A(n19726), .B(n19725), .Z(n19728) );
  AND U20117 ( .A(x[239]), .B(y[1995]), .Z(n20361) );
  NAND U20118 ( .A(n20361), .B(n19529), .Z(n19533) );
  NAND U20119 ( .A(n19531), .B(n19530), .Z(n19532) );
  NAND U20120 ( .A(n19533), .B(n19532), .Z(n19684) );
  AND U20121 ( .A(x[224]), .B(y[2005]), .Z(n19703) );
  AND U20122 ( .A(x[245]), .B(y[1984]), .Z(n19704) );
  XOR U20123 ( .A(n19703), .B(n19704), .Z(n19706) );
  AND U20124 ( .A(o[212]), .B(n19534), .Z(n19705) );
  XOR U20125 ( .A(n19706), .B(n19705), .Z(n19682) );
  AND U20126 ( .A(x[229]), .B(y[2000]), .Z(n19690) );
  AND U20127 ( .A(x[240]), .B(y[1989]), .Z(n19689) );
  XOR U20128 ( .A(n19690), .B(n19689), .Z(n19688) );
  AND U20129 ( .A(x[239]), .B(y[1990]), .Z(n19687) );
  XOR U20130 ( .A(n19688), .B(n19687), .Z(n19681) );
  XOR U20131 ( .A(n19682), .B(n19681), .Z(n19683) );
  XOR U20132 ( .A(n19684), .B(n19683), .Z(n19727) );
  XOR U20133 ( .A(n19728), .B(n19727), .Z(n19720) );
  NAND U20134 ( .A(n19536), .B(n19535), .Z(n19540) );
  NAND U20135 ( .A(n19538), .B(n19537), .Z(n19539) );
  NAND U20136 ( .A(n19540), .B(n19539), .Z(n19719) );
  NAND U20137 ( .A(n19542), .B(n19541), .Z(n19546) );
  NAND U20138 ( .A(n19544), .B(n19543), .Z(n19545) );
  AND U20139 ( .A(n19546), .B(n19545), .Z(n19721) );
  XNOR U20140 ( .A(n19722), .B(n19721), .Z(n19647) );
  NAND U20141 ( .A(n19548), .B(n19547), .Z(n19552) );
  NAND U20142 ( .A(n19550), .B(n19549), .Z(n19551) );
  AND U20143 ( .A(n19552), .B(n19551), .Z(n19646) );
  XOR U20144 ( .A(n19647), .B(n19646), .Z(n19648) );
  XNOR U20145 ( .A(n19649), .B(n19648), .Z(n19642) );
  NANDN U20146 ( .A(n19554), .B(n19553), .Z(n19558) );
  NAND U20147 ( .A(n19556), .B(n19555), .Z(n19557) );
  NAND U20148 ( .A(n19558), .B(n19557), .Z(n19746) );
  NAND U20149 ( .A(n20367), .B(n19559), .Z(n19563) );
  NAND U20150 ( .A(n19561), .B(n19560), .Z(n19562) );
  NAND U20151 ( .A(n19563), .B(n19562), .Z(n19653) );
  NAND U20152 ( .A(n20932), .B(n19564), .Z(n19568) );
  NAND U20153 ( .A(n19566), .B(n19565), .Z(n19567) );
  NAND U20154 ( .A(n19568), .B(n19567), .Z(n19740) );
  AND U20155 ( .A(y[1986]), .B(x[243]), .Z(n19570) );
  NAND U20156 ( .A(y[1994]), .B(x[235]), .Z(n19569) );
  XNOR U20157 ( .A(n19570), .B(n19569), .Z(n19672) );
  AND U20158 ( .A(x[244]), .B(y[1985]), .Z(n19702) );
  XOR U20159 ( .A(o[213]), .B(n19702), .Z(n19671) );
  XOR U20160 ( .A(n19672), .B(n19671), .Z(n19738) );
  AND U20161 ( .A(y[1987]), .B(x[242]), .Z(n19572) );
  NAND U20162 ( .A(y[1995]), .B(x[234]), .Z(n19571) );
  XNOR U20163 ( .A(n19572), .B(n19571), .Z(n19710) );
  AND U20164 ( .A(x[225]), .B(y[2004]), .Z(n19711) );
  XOR U20165 ( .A(n19710), .B(n19711), .Z(n19737) );
  XOR U20166 ( .A(n19738), .B(n19737), .Z(n19739) );
  XOR U20167 ( .A(n19740), .B(n19739), .Z(n19652) );
  XOR U20168 ( .A(n19653), .B(n19652), .Z(n19655) );
  AND U20169 ( .A(x[231]), .B(y[1998]), .Z(n19918) );
  AND U20170 ( .A(y[1999]), .B(x[230]), .Z(n19574) );
  NAND U20171 ( .A(y[1991]), .B(x[238]), .Z(n19573) );
  XNOR U20172 ( .A(n19574), .B(n19573), .Z(n19714) );
  XNOR U20173 ( .A(n19918), .B(n19714), .Z(n19661) );
  NAND U20174 ( .A(x[233]), .B(y[1996]), .Z(n19659) );
  NAND U20175 ( .A(x[232]), .B(y[1997]), .Z(n19658) );
  XOR U20176 ( .A(n19659), .B(n19658), .Z(n19660) );
  XNOR U20177 ( .A(n19661), .B(n19660), .Z(n19677) );
  AND U20178 ( .A(y[1993]), .B(x[236]), .Z(n19576) );
  NAND U20179 ( .A(y[1988]), .B(x[241]), .Z(n19575) );
  XNOR U20180 ( .A(n19576), .B(n19575), .Z(n19664) );
  AND U20181 ( .A(x[226]), .B(y[2003]), .Z(n19665) );
  XOR U20182 ( .A(n19664), .B(n19665), .Z(n19676) );
  AND U20183 ( .A(y[1992]), .B(x[237]), .Z(n19578) );
  NAND U20184 ( .A(y[2002]), .B(x[227]), .Z(n19577) );
  XNOR U20185 ( .A(n19578), .B(n19577), .Z(n19698) );
  AND U20186 ( .A(x[228]), .B(y[2001]), .Z(n19699) );
  XOR U20187 ( .A(n19698), .B(n19699), .Z(n19675) );
  XOR U20188 ( .A(n19676), .B(n19675), .Z(n19678) );
  XOR U20189 ( .A(n19677), .B(n19678), .Z(n19734) );
  NAND U20190 ( .A(n19690), .B(n19579), .Z(n19583) );
  NAND U20191 ( .A(n19581), .B(n19580), .Z(n19582) );
  NAND U20192 ( .A(n19583), .B(n19582), .Z(n19732) );
  NAND U20193 ( .A(n19585), .B(n19584), .Z(n19589) );
  NAND U20194 ( .A(n19587), .B(n19586), .Z(n19588) );
  NAND U20195 ( .A(n19589), .B(n19588), .Z(n19731) );
  XOR U20196 ( .A(n19732), .B(n19731), .Z(n19733) );
  XOR U20197 ( .A(n19734), .B(n19733), .Z(n19654) );
  XOR U20198 ( .A(n19655), .B(n19654), .Z(n19744) );
  NANDN U20199 ( .A(n19591), .B(n19590), .Z(n19595) );
  NAND U20200 ( .A(n19593), .B(n19592), .Z(n19594) );
  NAND U20201 ( .A(n19595), .B(n19594), .Z(n19751) );
  NAND U20202 ( .A(n19597), .B(n19596), .Z(n19601) );
  NANDN U20203 ( .A(n19599), .B(n19598), .Z(n19600) );
  NAND U20204 ( .A(n19601), .B(n19600), .Z(n19750) );
  NAND U20205 ( .A(n19603), .B(n19602), .Z(n19607) );
  NANDN U20206 ( .A(n19605), .B(n19604), .Z(n19606) );
  NAND U20207 ( .A(n19607), .B(n19606), .Z(n19749) );
  XOR U20208 ( .A(n19750), .B(n19749), .Z(n19752) );
  XOR U20209 ( .A(n19751), .B(n19752), .Z(n19743) );
  XOR U20210 ( .A(n19744), .B(n19743), .Z(n19745) );
  XNOR U20211 ( .A(n19746), .B(n19745), .Z(n19641) );
  NAND U20212 ( .A(n19609), .B(n19608), .Z(n19613) );
  NAND U20213 ( .A(n19611), .B(n19610), .Z(n19612) );
  NAND U20214 ( .A(n19613), .B(n19612), .Z(n19640) );
  XOR U20215 ( .A(n19641), .B(n19640), .Z(n19643) );
  XNOR U20216 ( .A(n19642), .B(n19643), .Z(n19760) );
  NAND U20217 ( .A(n19615), .B(n19614), .Z(n19619) );
  NAND U20218 ( .A(n19617), .B(n19616), .Z(n19618) );
  AND U20219 ( .A(n19619), .B(n19618), .Z(n19759) );
  NANDN U20220 ( .A(n19621), .B(n19620), .Z(n19625) );
  NAND U20221 ( .A(n19623), .B(n19622), .Z(n19624) );
  AND U20222 ( .A(n19625), .B(n19624), .Z(n19758) );
  XNOR U20223 ( .A(n19760), .B(n19761), .Z(n19757) );
  NANDN U20224 ( .A(n19626), .B(n19627), .Z(n19632) );
  NOR U20225 ( .A(n19628), .B(n19627), .Z(n19630) );
  OR U20226 ( .A(n19630), .B(n19629), .Z(n19631) );
  AND U20227 ( .A(n19632), .B(n19631), .Z(n19755) );
  NAND U20228 ( .A(n19634), .B(n19633), .Z(n19638) );
  NANDN U20229 ( .A(n19636), .B(n19635), .Z(n19637) );
  AND U20230 ( .A(n19638), .B(n19637), .Z(n19756) );
  XOR U20231 ( .A(n19755), .B(n19756), .Z(n19639) );
  XNOR U20232 ( .A(n19757), .B(n19639), .Z(N438) );
  NAND U20233 ( .A(n19641), .B(n19640), .Z(n19645) );
  NAND U20234 ( .A(n19643), .B(n19642), .Z(n19644) );
  AND U20235 ( .A(n19645), .B(n19644), .Z(n19895) );
  NAND U20236 ( .A(n19647), .B(n19646), .Z(n19651) );
  NAND U20237 ( .A(n19649), .B(n19648), .Z(n19650) );
  NAND U20238 ( .A(n19651), .B(n19650), .Z(n19893) );
  NAND U20239 ( .A(n19653), .B(n19652), .Z(n19657) );
  NAND U20240 ( .A(n19655), .B(n19654), .Z(n19656) );
  NAND U20241 ( .A(n19657), .B(n19656), .Z(n19876) );
  NAND U20242 ( .A(n19659), .B(n19658), .Z(n19663) );
  NAND U20243 ( .A(n19661), .B(n19660), .Z(n19662) );
  NAND U20244 ( .A(n19663), .B(n19662), .Z(n19870) );
  NANDN U20245 ( .A(n20375), .B(n19821), .Z(n19667) );
  NAND U20246 ( .A(n19665), .B(n19664), .Z(n19666) );
  NAND U20247 ( .A(n19667), .B(n19666), .Z(n19797) );
  AND U20248 ( .A(x[229]), .B(y[2001]), .Z(n19843) );
  AND U20249 ( .A(x[241]), .B(y[1989]), .Z(n19844) );
  XOR U20250 ( .A(n19843), .B(n19844), .Z(n19845) );
  AND U20251 ( .A(x[240]), .B(y[1990]), .Z(n19846) );
  XOR U20252 ( .A(n19845), .B(n19846), .Z(n19796) );
  AND U20253 ( .A(y[1988]), .B(x[242]), .Z(n19669) );
  NAND U20254 ( .A(y[1994]), .B(x[236]), .Z(n19668) );
  XNOR U20255 ( .A(n19669), .B(n19668), .Z(n19822) );
  AND U20256 ( .A(x[228]), .B(y[2002]), .Z(n19823) );
  XOR U20257 ( .A(n19822), .B(n19823), .Z(n19795) );
  XOR U20258 ( .A(n19796), .B(n19795), .Z(n19798) );
  XNOR U20259 ( .A(n19797), .B(n19798), .Z(n19867) );
  NAND U20260 ( .A(x[243]), .B(y[1994]), .Z(n20841) );
  NANDN U20261 ( .A(n20841), .B(n19670), .Z(n19674) );
  NAND U20262 ( .A(n19672), .B(n19671), .Z(n19673) );
  AND U20263 ( .A(n19674), .B(n19673), .Z(n19868) );
  XOR U20264 ( .A(n19867), .B(n19868), .Z(n19869) );
  XNOR U20265 ( .A(n19870), .B(n19869), .Z(n19873) );
  NAND U20266 ( .A(n19676), .B(n19675), .Z(n19680) );
  NAND U20267 ( .A(n19678), .B(n19677), .Z(n19679) );
  NAND U20268 ( .A(n19680), .B(n19679), .Z(n19856) );
  NAND U20269 ( .A(n19682), .B(n19681), .Z(n19686) );
  NAND U20270 ( .A(n19684), .B(n19683), .Z(n19685) );
  NAND U20271 ( .A(n19686), .B(n19685), .Z(n19855) );
  XOR U20272 ( .A(n19856), .B(n19855), .Z(n19858) );
  AND U20273 ( .A(n19688), .B(n19687), .Z(n19692) );
  NAND U20274 ( .A(n19690), .B(n19689), .Z(n19691) );
  NANDN U20275 ( .A(n19692), .B(n19691), .Z(n19818) );
  AND U20276 ( .A(y[1993]), .B(x[237]), .Z(n19694) );
  NAND U20277 ( .A(y[1986]), .B(x[244]), .Z(n19693) );
  XNOR U20278 ( .A(n19694), .B(n19693), .Z(n19839) );
  AND U20279 ( .A(x[226]), .B(y[2004]), .Z(n19840) );
  XOR U20280 ( .A(n19839), .B(n19840), .Z(n19816) );
  AND U20281 ( .A(y[2000]), .B(x[230]), .Z(n19696) );
  NAND U20282 ( .A(y[1991]), .B(x[239]), .Z(n19695) );
  XNOR U20283 ( .A(n19696), .B(n19695), .Z(n19851) );
  XOR U20284 ( .A(n19816), .B(n19815), .Z(n19817) );
  XOR U20285 ( .A(n19818), .B(n19817), .Z(n19862) );
  AND U20286 ( .A(x[237]), .B(y[2002]), .Z(n21017) );
  NAND U20287 ( .A(n19697), .B(n21017), .Z(n19701) );
  NAND U20288 ( .A(n19699), .B(n19698), .Z(n19700) );
  NAND U20289 ( .A(n19701), .B(n19700), .Z(n19786) );
  AND U20290 ( .A(x[225]), .B(y[2005]), .Z(n19809) );
  XOR U20291 ( .A(n19810), .B(n19809), .Z(n19808) );
  AND U20292 ( .A(o[213]), .B(n19702), .Z(n19807) );
  XOR U20293 ( .A(n19808), .B(n19807), .Z(n19784) );
  AND U20294 ( .A(x[238]), .B(y[1992]), .Z(n19801) );
  NAND U20295 ( .A(x[227]), .B(y[2003]), .Z(n19802) );
  NAND U20296 ( .A(x[243]), .B(y[1987]), .Z(n19804) );
  XOR U20297 ( .A(n19784), .B(n19783), .Z(n19785) );
  XOR U20298 ( .A(n19786), .B(n19785), .Z(n19861) );
  XOR U20299 ( .A(n19862), .B(n19861), .Z(n19864) );
  NAND U20300 ( .A(n19704), .B(n19703), .Z(n19708) );
  NAND U20301 ( .A(n19706), .B(n19705), .Z(n19707) );
  NAND U20302 ( .A(n19708), .B(n19707), .Z(n19778) );
  AND U20303 ( .A(x[242]), .B(y[1995]), .Z(n20843) );
  NAND U20304 ( .A(n20843), .B(n19709), .Z(n19713) );
  NAND U20305 ( .A(n19711), .B(n19710), .Z(n19712) );
  NAND U20306 ( .A(n19713), .B(n19712), .Z(n19777) );
  XOR U20307 ( .A(n19778), .B(n19777), .Z(n19780) );
  AND U20308 ( .A(x[238]), .B(y[1999]), .Z(n20881) );
  NAND U20309 ( .A(n20881), .B(n19850), .Z(n19716) );
  NAND U20310 ( .A(n19918), .B(n19714), .Z(n19715) );
  NAND U20311 ( .A(n19716), .B(n19715), .Z(n19792) );
  AND U20312 ( .A(x[224]), .B(y[2006]), .Z(n19826) );
  NAND U20313 ( .A(x[246]), .B(y[1984]), .Z(n19827) );
  NAND U20314 ( .A(x[245]), .B(y[1985]), .Z(n19849) );
  XOR U20315 ( .A(n19829), .B(n19828), .Z(n19790) );
  AND U20316 ( .A(y[1999]), .B(x[231]), .Z(n19718) );
  NAND U20317 ( .A(y[1998]), .B(x[232]), .Z(n19717) );
  XNOR U20318 ( .A(n19718), .B(n19717), .Z(n19832) );
  XOR U20319 ( .A(n19790), .B(n19789), .Z(n19791) );
  XOR U20320 ( .A(n19792), .B(n19791), .Z(n19779) );
  XOR U20321 ( .A(n19780), .B(n19779), .Z(n19863) );
  XOR U20322 ( .A(n19864), .B(n19863), .Z(n19857) );
  XOR U20323 ( .A(n19858), .B(n19857), .Z(n19874) );
  XOR U20324 ( .A(n19873), .B(n19874), .Z(n19875) );
  XNOR U20325 ( .A(n19876), .B(n19875), .Z(n19767) );
  NANDN U20326 ( .A(n19720), .B(n19719), .Z(n19724) );
  NAND U20327 ( .A(n19722), .B(n19721), .Z(n19723) );
  AND U20328 ( .A(n19724), .B(n19723), .Z(n19766) );
  NAND U20329 ( .A(n19726), .B(n19725), .Z(n19730) );
  NAND U20330 ( .A(n19728), .B(n19727), .Z(n19729) );
  AND U20331 ( .A(n19730), .B(n19729), .Z(n19774) );
  NAND U20332 ( .A(n19732), .B(n19731), .Z(n19736) );
  NAND U20333 ( .A(n19734), .B(n19733), .Z(n19735) );
  NAND U20334 ( .A(n19736), .B(n19735), .Z(n19772) );
  NAND U20335 ( .A(n19738), .B(n19737), .Z(n19742) );
  NAND U20336 ( .A(n19740), .B(n19739), .Z(n19741) );
  NAND U20337 ( .A(n19742), .B(n19741), .Z(n19771) );
  XOR U20338 ( .A(n19772), .B(n19771), .Z(n19773) );
  XOR U20339 ( .A(n19774), .B(n19773), .Z(n19765) );
  XNOR U20340 ( .A(n19767), .B(n19768), .Z(n19881) );
  NAND U20341 ( .A(n19744), .B(n19743), .Z(n19748) );
  NAND U20342 ( .A(n19746), .B(n19745), .Z(n19747) );
  AND U20343 ( .A(n19748), .B(n19747), .Z(n19880) );
  NAND U20344 ( .A(n19750), .B(n19749), .Z(n19754) );
  NAND U20345 ( .A(n19752), .B(n19751), .Z(n19753) );
  NAND U20346 ( .A(n19754), .B(n19753), .Z(n19879) );
  XOR U20347 ( .A(n19881), .B(n19882), .Z(n19892) );
  XOR U20348 ( .A(n19893), .B(n19892), .Z(n19894) );
  XNOR U20349 ( .A(n19895), .B(n19894), .Z(n19888) );
  NANDN U20350 ( .A(n19759), .B(n19758), .Z(n19763) );
  NAND U20351 ( .A(n19761), .B(n19760), .Z(n19762) );
  NAND U20352 ( .A(n19763), .B(n19762), .Z(n19886) );
  IV U20353 ( .A(n19886), .Z(n19885) );
  XOR U20354 ( .A(n19887), .B(n19885), .Z(n19764) );
  XNOR U20355 ( .A(n19888), .B(n19764), .Z(N439) );
  NANDN U20356 ( .A(n19766), .B(n19765), .Z(n19770) );
  NAND U20357 ( .A(n19768), .B(n19767), .Z(n19769) );
  AND U20358 ( .A(n19770), .B(n19769), .Z(n20030) );
  NAND U20359 ( .A(n19772), .B(n19771), .Z(n19776) );
  NANDN U20360 ( .A(n19774), .B(n19773), .Z(n19775) );
  NAND U20361 ( .A(n19776), .B(n19775), .Z(n20014) );
  NAND U20362 ( .A(n19778), .B(n19777), .Z(n19782) );
  NAND U20363 ( .A(n19780), .B(n19779), .Z(n19781) );
  NAND U20364 ( .A(n19782), .B(n19781), .Z(n20008) );
  NAND U20365 ( .A(n19784), .B(n19783), .Z(n19788) );
  NAND U20366 ( .A(n19786), .B(n19785), .Z(n19787) );
  NAND U20367 ( .A(n19788), .B(n19787), .Z(n20006) );
  NAND U20368 ( .A(n19790), .B(n19789), .Z(n19794) );
  NAND U20369 ( .A(n19792), .B(n19791), .Z(n19793) );
  NAND U20370 ( .A(n19794), .B(n19793), .Z(n20005) );
  XOR U20371 ( .A(n20006), .B(n20005), .Z(n20007) );
  XOR U20372 ( .A(n20008), .B(n20007), .Z(n20026) );
  NAND U20373 ( .A(n19796), .B(n19795), .Z(n19800) );
  NAND U20374 ( .A(n19798), .B(n19797), .Z(n19799) );
  NAND U20375 ( .A(n19800), .B(n19799), .Z(n20024) );
  NANDN U20376 ( .A(n19802), .B(n19801), .Z(n19806) );
  NANDN U20377 ( .A(n19804), .B(n19803), .Z(n19805) );
  NAND U20378 ( .A(n19806), .B(n19805), .Z(n19952) );
  AND U20379 ( .A(n19808), .B(n19807), .Z(n19812) );
  NAND U20380 ( .A(n19810), .B(n19809), .Z(n19811) );
  NANDN U20381 ( .A(n19812), .B(n19811), .Z(n19951) );
  XOR U20382 ( .A(n19952), .B(n19951), .Z(n19954) );
  AND U20383 ( .A(y[2000]), .B(x[231]), .Z(n19814) );
  NAND U20384 ( .A(y[1998]), .B(x[233]), .Z(n19813) );
  XNOR U20385 ( .A(n19814), .B(n19813), .Z(n19919) );
  NAND U20386 ( .A(x[234]), .B(y[1997]), .Z(n19958) );
  AND U20387 ( .A(x[230]), .B(y[2001]), .Z(n19910) );
  NAND U20388 ( .A(x[239]), .B(y[1992]), .Z(n19911) );
  NAND U20389 ( .A(x[235]), .B(y[1996]), .Z(n19913) );
  XOR U20390 ( .A(n19960), .B(n19959), .Z(n19953) );
  XOR U20391 ( .A(n19954), .B(n19953), .Z(n20023) );
  XOR U20392 ( .A(n20024), .B(n20023), .Z(n20025) );
  XOR U20393 ( .A(n20026), .B(n20025), .Z(n20012) );
  NAND U20394 ( .A(n19816), .B(n19815), .Z(n19820) );
  NAND U20395 ( .A(n19818), .B(n19817), .Z(n19819) );
  NAND U20396 ( .A(n19820), .B(n19819), .Z(n19946) );
  AND U20397 ( .A(x[242]), .B(y[1994]), .Z(n20701) );
  NAND U20398 ( .A(n20701), .B(n19821), .Z(n19825) );
  NAND U20399 ( .A(n19823), .B(n19822), .Z(n19824) );
  NAND U20400 ( .A(n19825), .B(n19824), .Z(n19982) );
  NANDN U20401 ( .A(n19827), .B(n19826), .Z(n19831) );
  NAND U20402 ( .A(n19829), .B(n19828), .Z(n19830) );
  NAND U20403 ( .A(n19831), .B(n19830), .Z(n19981) );
  XOR U20404 ( .A(n19982), .B(n19981), .Z(n19983) );
  NANDN U20405 ( .A(n19920), .B(n19918), .Z(n19835) );
  NANDN U20406 ( .A(n19833), .B(n19832), .Z(n19834) );
  NAND U20407 ( .A(n19835), .B(n19834), .Z(n19995) );
  AND U20408 ( .A(x[224]), .B(y[2007]), .Z(n19929) );
  NAND U20409 ( .A(x[247]), .B(y[1984]), .Z(n19930) );
  NAND U20410 ( .A(x[246]), .B(y[1985]), .Z(n19909) );
  XOR U20411 ( .A(n19932), .B(n19931), .Z(n19994) );
  NAND U20412 ( .A(y[1987]), .B(x[244]), .Z(n19836) );
  XNOR U20413 ( .A(n19837), .B(n19836), .Z(n19905) );
  NAND U20414 ( .A(x[243]), .B(y[1988]), .Z(n19906) );
  XOR U20415 ( .A(n19994), .B(n19993), .Z(n19996) );
  XOR U20416 ( .A(n19995), .B(n19996), .Z(n19984) );
  XOR U20417 ( .A(n19983), .B(n19984), .Z(n19945) );
  XOR U20418 ( .A(n19946), .B(n19945), .Z(n19948) );
  NAND U20419 ( .A(x[244]), .B(y[1993]), .Z(n20889) );
  AND U20420 ( .A(x[237]), .B(y[1986]), .Z(n19838) );
  NANDN U20421 ( .A(n20889), .B(n19838), .Z(n19842) );
  NAND U20422 ( .A(n19840), .B(n19839), .Z(n19841) );
  NAND U20423 ( .A(n19842), .B(n19841), .Z(n19940) );
  NAND U20424 ( .A(n19844), .B(n19843), .Z(n19848) );
  NAND U20425 ( .A(n19846), .B(n19845), .Z(n19847) );
  NAND U20426 ( .A(n19848), .B(n19847), .Z(n20001) );
  AND U20427 ( .A(x[237]), .B(y[1994]), .Z(n19975) );
  AND U20428 ( .A(x[226]), .B(y[2005]), .Z(n19976) );
  XOR U20429 ( .A(n19975), .B(n19976), .Z(n19977) );
  AND U20430 ( .A(x[245]), .B(y[1986]), .Z(n19978) );
  XOR U20431 ( .A(n19977), .B(n19978), .Z(n20000) );
  AND U20432 ( .A(x[236]), .B(y[1995]), .Z(n19923) );
  NAND U20433 ( .A(x[225]), .B(y[2006]), .Z(n19924) );
  ANDN U20434 ( .B(o[214]), .A(n19849), .Z(n19925) );
  XOR U20435 ( .A(n19926), .B(n19925), .Z(n19999) );
  XOR U20436 ( .A(n20000), .B(n19999), .Z(n20002) );
  XOR U20437 ( .A(n20001), .B(n20002), .Z(n19939) );
  XOR U20438 ( .A(n19940), .B(n19939), .Z(n19942) );
  AND U20439 ( .A(x[239]), .B(y[2000]), .Z(n21011) );
  NAND U20440 ( .A(n21011), .B(n19850), .Z(n19854) );
  NANDN U20441 ( .A(n19852), .B(n19851), .Z(n19853) );
  NAND U20442 ( .A(n19854), .B(n19853), .Z(n19989) );
  AND U20443 ( .A(x[238]), .B(y[1993]), .Z(n19969) );
  AND U20444 ( .A(x[227]), .B(y[2004]), .Z(n19970) );
  XOR U20445 ( .A(n19969), .B(n19970), .Z(n19971) );
  AND U20446 ( .A(x[228]), .B(y[2003]), .Z(n19972) );
  XOR U20447 ( .A(n19971), .B(n19972), .Z(n19988) );
  AND U20448 ( .A(x[229]), .B(y[2002]), .Z(n19963) );
  AND U20449 ( .A(x[242]), .B(y[1989]), .Z(n19964) );
  XOR U20450 ( .A(n19963), .B(n19964), .Z(n19966) );
  AND U20451 ( .A(x[241]), .B(y[1990]), .Z(n19965) );
  XOR U20452 ( .A(n19966), .B(n19965), .Z(n19987) );
  XOR U20453 ( .A(n19988), .B(n19987), .Z(n19990) );
  XOR U20454 ( .A(n19989), .B(n19990), .Z(n19941) );
  XOR U20455 ( .A(n19942), .B(n19941), .Z(n19947) );
  XOR U20456 ( .A(n19948), .B(n19947), .Z(n20011) );
  XOR U20457 ( .A(n20012), .B(n20011), .Z(n20013) );
  XNOR U20458 ( .A(n20014), .B(n20013), .Z(n19901) );
  NAND U20459 ( .A(n19856), .B(n19855), .Z(n19860) );
  NAND U20460 ( .A(n19858), .B(n19857), .Z(n19859) );
  NAND U20461 ( .A(n19860), .B(n19859), .Z(n20020) );
  NAND U20462 ( .A(n19862), .B(n19861), .Z(n19866) );
  NAND U20463 ( .A(n19864), .B(n19863), .Z(n19865) );
  NAND U20464 ( .A(n19866), .B(n19865), .Z(n20018) );
  NAND U20465 ( .A(n19868), .B(n19867), .Z(n19872) );
  NAND U20466 ( .A(n19870), .B(n19869), .Z(n19871) );
  AND U20467 ( .A(n19872), .B(n19871), .Z(n20017) );
  XOR U20468 ( .A(n20018), .B(n20017), .Z(n20019) );
  XNOR U20469 ( .A(n20020), .B(n20019), .Z(n19899) );
  NAND U20470 ( .A(n19874), .B(n19873), .Z(n19878) );
  NAND U20471 ( .A(n19876), .B(n19875), .Z(n19877) );
  AND U20472 ( .A(n19878), .B(n19877), .Z(n19900) );
  XOR U20473 ( .A(n19899), .B(n19900), .Z(n19902) );
  XOR U20474 ( .A(n19901), .B(n19902), .Z(n20029) );
  NANDN U20475 ( .A(n19880), .B(n19879), .Z(n19884) );
  NAND U20476 ( .A(n19882), .B(n19881), .Z(n19883) );
  AND U20477 ( .A(n19884), .B(n19883), .Z(n20031) );
  XNOR U20478 ( .A(n20032), .B(n20031), .Z(n20038) );
  OR U20479 ( .A(n19887), .B(n19885), .Z(n19891) );
  ANDN U20480 ( .B(n19887), .A(n19886), .Z(n19889) );
  OR U20481 ( .A(n19889), .B(n19888), .Z(n19890) );
  AND U20482 ( .A(n19891), .B(n19890), .Z(n20036) );
  NAND U20483 ( .A(n19893), .B(n19892), .Z(n19897) );
  NAND U20484 ( .A(n19895), .B(n19894), .Z(n19896) );
  AND U20485 ( .A(n19897), .B(n19896), .Z(n20037) );
  IV U20486 ( .A(n20037), .Z(n20035) );
  XOR U20487 ( .A(n20036), .B(n20035), .Z(n19898) );
  XNOR U20488 ( .A(n20038), .B(n19898), .Z(N440) );
  NAND U20489 ( .A(n19900), .B(n19899), .Z(n19904) );
  NAND U20490 ( .A(n19902), .B(n19901), .Z(n19903) );
  AND U20491 ( .A(n19904), .B(n19903), .Z(n20178) );
  AND U20492 ( .A(x[244]), .B(y[1991]), .Z(n20476) );
  NAND U20493 ( .A(n20476), .B(n20146), .Z(n19908) );
  NANDN U20494 ( .A(n19906), .B(n19905), .Z(n19907) );
  AND U20495 ( .A(n19908), .B(n19907), .Z(n20160) );
  AND U20496 ( .A(x[246]), .B(y[1986]), .Z(n20071) );
  XOR U20497 ( .A(n20072), .B(n20071), .Z(n20074) );
  AND U20498 ( .A(x[226]), .B(y[2006]), .Z(n20073) );
  XOR U20499 ( .A(n20074), .B(n20073), .Z(n20158) );
  AND U20500 ( .A(x[225]), .B(y[2007]), .Z(n20079) );
  XOR U20501 ( .A(n20080), .B(n20079), .Z(n20078) );
  ANDN U20502 ( .B(o[215]), .A(n19909), .Z(n20077) );
  XOR U20503 ( .A(n20078), .B(n20077), .Z(n20157) );
  XOR U20504 ( .A(n20158), .B(n20157), .Z(n20159) );
  NANDN U20505 ( .A(n19911), .B(n19910), .Z(n19915) );
  NANDN U20506 ( .A(n19913), .B(n19912), .Z(n19914) );
  AND U20507 ( .A(n19915), .B(n19914), .Z(n20166) );
  AND U20508 ( .A(y[1992]), .B(x[240]), .Z(n19917) );
  NAND U20509 ( .A(y[1987]), .B(x[245]), .Z(n19916) );
  XNOR U20510 ( .A(n19917), .B(n19916), .Z(n20148) );
  AND U20511 ( .A(x[229]), .B(y[2003]), .Z(n20147) );
  XOR U20512 ( .A(n20148), .B(n20147), .Z(n20164) );
  AND U20513 ( .A(x[230]), .B(y[2002]), .Z(n20464) );
  AND U20514 ( .A(x[244]), .B(y[1988]), .Z(n20293) );
  XOR U20515 ( .A(n20464), .B(n20293), .Z(n20154) );
  AND U20516 ( .A(x[243]), .B(y[1989]), .Z(n20153) );
  XOR U20517 ( .A(n20154), .B(n20153), .Z(n20163) );
  XOR U20518 ( .A(n20164), .B(n20163), .Z(n20165) );
  NANDN U20519 ( .A(n20090), .B(n19918), .Z(n19922) );
  NANDN U20520 ( .A(n19920), .B(n19919), .Z(n19921) );
  AND U20521 ( .A(n19922), .B(n19921), .Z(n20135) );
  NANDN U20522 ( .A(n19924), .B(n19923), .Z(n19928) );
  NAND U20523 ( .A(n19926), .B(n19925), .Z(n19927) );
  NAND U20524 ( .A(n19928), .B(n19927), .Z(n20134) );
  XOR U20525 ( .A(n20137), .B(n20136), .Z(n20110) );
  XOR U20526 ( .A(n20111), .B(n20110), .Z(n20113) );
  NANDN U20527 ( .A(n19930), .B(n19929), .Z(n19934) );
  NAND U20528 ( .A(n19932), .B(n19931), .Z(n19933) );
  AND U20529 ( .A(n19934), .B(n19933), .Z(n20105) );
  AND U20530 ( .A(x[227]), .B(y[2005]), .Z(n20092) );
  XOR U20531 ( .A(n20093), .B(n20092), .Z(n20095) );
  NAND U20532 ( .A(x[228]), .B(y[2004]), .Z(n20094) );
  AND U20533 ( .A(y[1999]), .B(x[233]), .Z(n19936) );
  NAND U20534 ( .A(y[1998]), .B(x[234]), .Z(n19935) );
  XNOR U20535 ( .A(n19936), .B(n19935), .Z(n20063) );
  AND U20536 ( .A(y[1994]), .B(x[238]), .Z(n19938) );
  NAND U20537 ( .A(y[2000]), .B(x[232]), .Z(n19937) );
  XNOR U20538 ( .A(n19938), .B(n19937), .Z(n20067) );
  NAND U20539 ( .A(x[235]), .B(y[1997]), .Z(n20068) );
  XOR U20540 ( .A(n20063), .B(n20062), .Z(n20106) );
  XOR U20541 ( .A(n20107), .B(n20106), .Z(n20112) );
  XOR U20542 ( .A(n20113), .B(n20112), .Z(n20056) );
  NAND U20543 ( .A(n19940), .B(n19939), .Z(n19944) );
  NAND U20544 ( .A(n19942), .B(n19941), .Z(n19943) );
  AND U20545 ( .A(n19944), .B(n19943), .Z(n20055) );
  NAND U20546 ( .A(n19946), .B(n19945), .Z(n19950) );
  NAND U20547 ( .A(n19948), .B(n19947), .Z(n19949) );
  NAND U20548 ( .A(n19950), .B(n19949), .Z(n20058) );
  NAND U20549 ( .A(n19952), .B(n19951), .Z(n19956) );
  NAND U20550 ( .A(n19954), .B(n19953), .Z(n19955) );
  AND U20551 ( .A(n19956), .B(n19955), .Z(n20119) );
  NANDN U20552 ( .A(n19958), .B(n19957), .Z(n19962) );
  NAND U20553 ( .A(n19960), .B(n19959), .Z(n19961) );
  AND U20554 ( .A(n19962), .B(n19961), .Z(n20117) );
  NAND U20555 ( .A(n19964), .B(n19963), .Z(n19968) );
  NAND U20556 ( .A(n19966), .B(n19965), .Z(n19967) );
  AND U20557 ( .A(n19968), .B(n19967), .Z(n20143) );
  AND U20558 ( .A(x[224]), .B(y[2008]), .Z(n20099) );
  AND U20559 ( .A(x[248]), .B(y[1984]), .Z(n20098) );
  XOR U20560 ( .A(n20099), .B(n20098), .Z(n20101) );
  AND U20561 ( .A(x[247]), .B(y[1985]), .Z(n20091) );
  XOR U20562 ( .A(n20091), .B(o[216]), .Z(n20100) );
  XOR U20563 ( .A(n20101), .B(n20100), .Z(n20141) );
  AND U20564 ( .A(x[231]), .B(y[2001]), .Z(n20084) );
  AND U20565 ( .A(x[242]), .B(y[1990]), .Z(n20083) );
  XOR U20566 ( .A(n20084), .B(n20083), .Z(n20086) );
  AND U20567 ( .A(x[241]), .B(y[1991]), .Z(n20085) );
  XOR U20568 ( .A(n20086), .B(n20085), .Z(n20140) );
  XOR U20569 ( .A(n20141), .B(n20140), .Z(n20142) );
  NAND U20570 ( .A(n19970), .B(n19969), .Z(n19974) );
  NAND U20571 ( .A(n19972), .B(n19971), .Z(n19973) );
  AND U20572 ( .A(n19974), .B(n19973), .Z(n20129) );
  NAND U20573 ( .A(n19976), .B(n19975), .Z(n19980) );
  NAND U20574 ( .A(n19978), .B(n19977), .Z(n19979) );
  NAND U20575 ( .A(n19980), .B(n19979), .Z(n20128) );
  XOR U20576 ( .A(n20131), .B(n20130), .Z(n20116) );
  NAND U20577 ( .A(n19982), .B(n19981), .Z(n19986) );
  NAND U20578 ( .A(n19984), .B(n19983), .Z(n19985) );
  AND U20579 ( .A(n19986), .B(n19985), .Z(n20172) );
  NAND U20580 ( .A(n19988), .B(n19987), .Z(n19992) );
  NAND U20581 ( .A(n19990), .B(n19989), .Z(n19991) );
  AND U20582 ( .A(n19992), .B(n19991), .Z(n20170) );
  NAND U20583 ( .A(n19994), .B(n19993), .Z(n19998) );
  NAND U20584 ( .A(n19996), .B(n19995), .Z(n19997) );
  AND U20585 ( .A(n19998), .B(n19997), .Z(n20169) );
  XOR U20586 ( .A(n20170), .B(n20169), .Z(n20171) );
  XOR U20587 ( .A(n20172), .B(n20171), .Z(n20122) );
  NAND U20588 ( .A(n20000), .B(n19999), .Z(n20004) );
  NAND U20589 ( .A(n20002), .B(n20001), .Z(n20003) );
  NAND U20590 ( .A(n20004), .B(n20003), .Z(n20123) );
  XOR U20591 ( .A(n20124), .B(n20125), .Z(n20049) );
  NAND U20592 ( .A(n20006), .B(n20005), .Z(n20010) );
  NAND U20593 ( .A(n20008), .B(n20007), .Z(n20009) );
  AND U20594 ( .A(n20010), .B(n20009), .Z(n20050) );
  XOR U20595 ( .A(n20049), .B(n20050), .Z(n20051) );
  XNOR U20596 ( .A(n20052), .B(n20051), .Z(n20176) );
  NAND U20597 ( .A(n20012), .B(n20011), .Z(n20016) );
  NAND U20598 ( .A(n20014), .B(n20013), .Z(n20015) );
  NAND U20599 ( .A(n20016), .B(n20015), .Z(n20046) );
  NAND U20600 ( .A(n20018), .B(n20017), .Z(n20022) );
  NAND U20601 ( .A(n20020), .B(n20019), .Z(n20021) );
  NAND U20602 ( .A(n20022), .B(n20021), .Z(n20044) );
  NAND U20603 ( .A(n20024), .B(n20023), .Z(n20028) );
  NAND U20604 ( .A(n20026), .B(n20025), .Z(n20027) );
  NAND U20605 ( .A(n20028), .B(n20027), .Z(n20043) );
  XOR U20606 ( .A(n20044), .B(n20043), .Z(n20045) );
  XOR U20607 ( .A(n20046), .B(n20045), .Z(n20175) );
  XOR U20608 ( .A(n20176), .B(n20175), .Z(n20177) );
  XOR U20609 ( .A(n20178), .B(n20177), .Z(n20183) );
  NANDN U20610 ( .A(n20030), .B(n20029), .Z(n20034) );
  NAND U20611 ( .A(n20032), .B(n20031), .Z(n20033) );
  NAND U20612 ( .A(n20034), .B(n20033), .Z(n20181) );
  NANDN U20613 ( .A(n20035), .B(n20036), .Z(n20041) );
  NOR U20614 ( .A(n20037), .B(n20036), .Z(n20039) );
  OR U20615 ( .A(n20039), .B(n20038), .Z(n20040) );
  AND U20616 ( .A(n20041), .B(n20040), .Z(n20182) );
  XOR U20617 ( .A(n20181), .B(n20182), .Z(n20042) );
  XNOR U20618 ( .A(n20183), .B(n20042), .Z(N441) );
  NAND U20619 ( .A(n20044), .B(n20043), .Z(n20048) );
  NAND U20620 ( .A(n20046), .B(n20045), .Z(n20047) );
  AND U20621 ( .A(n20048), .B(n20047), .Z(n20188) );
  NAND U20622 ( .A(n20050), .B(n20049), .Z(n20054) );
  NAND U20623 ( .A(n20052), .B(n20051), .Z(n20053) );
  NAND U20624 ( .A(n20054), .B(n20053), .Z(n20186) );
  NANDN U20625 ( .A(n20056), .B(n20055), .Z(n20060) );
  NANDN U20626 ( .A(n20058), .B(n20057), .Z(n20059) );
  NAND U20627 ( .A(n20060), .B(n20059), .Z(n20194) );
  NANDN U20628 ( .A(n20218), .B(n20061), .Z(n20065) );
  NAND U20629 ( .A(n20063), .B(n20062), .Z(n20064) );
  AND U20630 ( .A(n20065), .B(n20064), .Z(n20243) );
  AND U20631 ( .A(x[238]), .B(y[2000]), .Z(n21051) );
  NAND U20632 ( .A(n21051), .B(n20066), .Z(n20070) );
  NANDN U20633 ( .A(n20068), .B(n20067), .Z(n20069) );
  AND U20634 ( .A(n20070), .B(n20069), .Z(n20271) );
  NAND U20635 ( .A(x[235]), .B(y[1998]), .Z(n20289) );
  NAND U20636 ( .A(x[236]), .B(y[1997]), .Z(n20288) );
  NAND U20637 ( .A(x[231]), .B(y[2002]), .Z(n20287) );
  XNOR U20638 ( .A(n20288), .B(n20287), .Z(n20290) );
  AND U20639 ( .A(x[248]), .B(y[1985]), .Z(n20286) );
  XOR U20640 ( .A(o[217]), .B(n20286), .Z(n20256) );
  NAND U20641 ( .A(x[225]), .B(y[2008]), .Z(n20257) );
  NAND U20642 ( .A(x[237]), .B(y[1996]), .Z(n20259) );
  XOR U20643 ( .A(n20268), .B(n20269), .Z(n20270) );
  NAND U20644 ( .A(n20072), .B(n20071), .Z(n20076) );
  AND U20645 ( .A(n20074), .B(n20073), .Z(n20075) );
  ANDN U20646 ( .B(n20076), .A(n20075), .Z(n20231) );
  AND U20647 ( .A(n20078), .B(n20077), .Z(n20082) );
  NAND U20648 ( .A(n20080), .B(n20079), .Z(n20081) );
  NANDN U20649 ( .A(n20082), .B(n20081), .Z(n20230) );
  NAND U20650 ( .A(n20084), .B(n20083), .Z(n20088) );
  NAND U20651 ( .A(n20086), .B(n20085), .Z(n20087) );
  AND U20652 ( .A(n20088), .B(n20087), .Z(n20227) );
  AND U20653 ( .A(x[232]), .B(y[2001]), .Z(n20221) );
  XNOR U20654 ( .A(n20090), .B(n20089), .Z(n20220) );
  AND U20655 ( .A(n20091), .B(o[216]), .Z(n20215) );
  AND U20656 ( .A(x[249]), .B(y[1984]), .Z(n20213) );
  NAND U20657 ( .A(x[224]), .B(y[2009]), .Z(n20212) );
  XOR U20658 ( .A(n20215), .B(n20214), .Z(n20224) );
  XOR U20659 ( .A(n20225), .B(n20224), .Z(n20226) );
  XOR U20660 ( .A(n20233), .B(n20232), .Z(n20244) );
  XOR U20661 ( .A(n20245), .B(n20244), .Z(n20332) );
  NAND U20662 ( .A(n20093), .B(n20092), .Z(n20097) );
  ANDN U20663 ( .B(n20095), .A(n20094), .Z(n20096) );
  ANDN U20664 ( .B(n20097), .A(n20096), .Z(n20308) );
  NAND U20665 ( .A(n20099), .B(n20098), .Z(n20103) );
  NAND U20666 ( .A(n20101), .B(n20100), .Z(n20102) );
  AND U20667 ( .A(n20103), .B(n20102), .Z(n20306) );
  AND U20668 ( .A(x[238]), .B(y[1995]), .Z(n20262) );
  NAND U20669 ( .A(x[226]), .B(y[2007]), .Z(n20263) );
  NAND U20670 ( .A(x[227]), .B(y[2006]), .Z(n20265) );
  NANDN U20671 ( .A(n20105), .B(n20104), .Z(n20109) );
  NAND U20672 ( .A(n20107), .B(n20106), .Z(n20108) );
  AND U20673 ( .A(n20109), .B(n20108), .Z(n20329) );
  NAND U20674 ( .A(n20111), .B(n20110), .Z(n20115) );
  NAND U20675 ( .A(n20113), .B(n20112), .Z(n20114) );
  NAND U20676 ( .A(n20115), .B(n20114), .Z(n20324) );
  NANDN U20677 ( .A(n20117), .B(n20116), .Z(n20121) );
  NANDN U20678 ( .A(n20119), .B(n20118), .Z(n20120) );
  NAND U20679 ( .A(n20121), .B(n20120), .Z(n20326) );
  XOR U20680 ( .A(n20194), .B(n20195), .Z(n20196) );
  NANDN U20681 ( .A(n20123), .B(n20122), .Z(n20127) );
  NAND U20682 ( .A(n20125), .B(n20124), .Z(n20126) );
  NAND U20683 ( .A(n20127), .B(n20126), .Z(n20202) );
  NANDN U20684 ( .A(n20129), .B(n20128), .Z(n20133) );
  NAND U20685 ( .A(n20131), .B(n20130), .Z(n20132) );
  AND U20686 ( .A(n20133), .B(n20132), .Z(n20207) );
  NANDN U20687 ( .A(n20135), .B(n20134), .Z(n20139) );
  NAND U20688 ( .A(n20137), .B(n20136), .Z(n20138) );
  NAND U20689 ( .A(n20139), .B(n20138), .Z(n20206) );
  NAND U20690 ( .A(n20141), .B(n20140), .Z(n20145) );
  NANDN U20691 ( .A(n20143), .B(n20142), .Z(n20144) );
  AND U20692 ( .A(n20145), .B(n20144), .Z(n20239) );
  NAND U20693 ( .A(x[245]), .B(y[1992]), .Z(n20989) );
  NANDN U20694 ( .A(n20989), .B(n20146), .Z(n20150) );
  NAND U20695 ( .A(n20148), .B(n20147), .Z(n20149) );
  NAND U20696 ( .A(n20150), .B(n20149), .Z(n20313) );
  NAND U20697 ( .A(x[246]), .B(y[1987]), .Z(n20282) );
  NAND U20698 ( .A(x[229]), .B(y[2004]), .Z(n20281) );
  NAND U20699 ( .A(x[241]), .B(y[1992]), .Z(n20280) );
  XOR U20700 ( .A(n20281), .B(n20280), .Z(n20283) );
  XOR U20701 ( .A(n20282), .B(n20283), .Z(n20312) );
  AND U20702 ( .A(y[1989]), .B(x[244]), .Z(n20152) );
  NAND U20703 ( .A(y[1988]), .B(x[245]), .Z(n20151) );
  XNOR U20704 ( .A(n20152), .B(n20151), .Z(n20295) );
  AND U20705 ( .A(x[243]), .B(y[1990]), .Z(n20294) );
  XOR U20706 ( .A(n20295), .B(n20294), .Z(n20311) );
  XOR U20707 ( .A(n20313), .B(n20314), .Z(n20237) );
  NAND U20708 ( .A(n20464), .B(n20293), .Z(n20156) );
  NAND U20709 ( .A(n20154), .B(n20153), .Z(n20155) );
  NAND U20710 ( .A(n20156), .B(n20155), .Z(n20319) );
  NAND U20711 ( .A(x[239]), .B(y[1994]), .Z(n20301) );
  NAND U20712 ( .A(x[242]), .B(y[1991]), .Z(n20300) );
  NAND U20713 ( .A(x[230]), .B(y[2003]), .Z(n20299) );
  XOR U20714 ( .A(n20300), .B(n20299), .Z(n20302) );
  XOR U20715 ( .A(n20301), .B(n20302), .Z(n20318) );
  NAND U20716 ( .A(x[247]), .B(y[1986]), .Z(n20276) );
  NAND U20717 ( .A(x[228]), .B(y[2005]), .Z(n20275) );
  NAND U20718 ( .A(x[240]), .B(y[1993]), .Z(n20274) );
  XOR U20719 ( .A(n20275), .B(n20274), .Z(n20277) );
  XNOR U20720 ( .A(n20276), .B(n20277), .Z(n20317) );
  XOR U20721 ( .A(n20319), .B(n20320), .Z(n20236) );
  XOR U20722 ( .A(n20239), .B(n20238), .Z(n20251) );
  NAND U20723 ( .A(n20158), .B(n20157), .Z(n20162) );
  NANDN U20724 ( .A(n20160), .B(n20159), .Z(n20161) );
  AND U20725 ( .A(n20162), .B(n20161), .Z(n20249) );
  NAND U20726 ( .A(n20164), .B(n20163), .Z(n20168) );
  NANDN U20727 ( .A(n20166), .B(n20165), .Z(n20167) );
  NAND U20728 ( .A(n20168), .B(n20167), .Z(n20248) );
  XOR U20729 ( .A(n20209), .B(n20208), .Z(n20201) );
  NAND U20730 ( .A(n20170), .B(n20169), .Z(n20174) );
  NAND U20731 ( .A(n20172), .B(n20171), .Z(n20173) );
  NAND U20732 ( .A(n20174), .B(n20173), .Z(n20200) );
  XOR U20733 ( .A(n20202), .B(n20203), .Z(n20197) );
  XNOR U20734 ( .A(n20196), .B(n20197), .Z(n20185) );
  XOR U20735 ( .A(n20186), .B(n20185), .Z(n20187) );
  XOR U20736 ( .A(n20188), .B(n20187), .Z(n20193) );
  NAND U20737 ( .A(n20176), .B(n20175), .Z(n20180) );
  NAND U20738 ( .A(n20178), .B(n20177), .Z(n20179) );
  NAND U20739 ( .A(n20180), .B(n20179), .Z(n20192) );
  XOR U20740 ( .A(n20192), .B(n20191), .Z(n20184) );
  XNOR U20741 ( .A(n20193), .B(n20184), .Z(N442) );
  NAND U20742 ( .A(n20186), .B(n20185), .Z(n20190) );
  NAND U20743 ( .A(n20188), .B(n20187), .Z(n20189) );
  NAND U20744 ( .A(n20190), .B(n20189), .Z(n20486) );
  IV U20745 ( .A(n20486), .Z(n20484) );
  NAND U20746 ( .A(n20195), .B(n20194), .Z(n20199) );
  NANDN U20747 ( .A(n20197), .B(n20196), .Z(n20198) );
  AND U20748 ( .A(n20199), .B(n20198), .Z(n20492) );
  NANDN U20749 ( .A(n20201), .B(n20200), .Z(n20205) );
  NANDN U20750 ( .A(n20203), .B(n20202), .Z(n20204) );
  AND U20751 ( .A(n20205), .B(n20204), .Z(n20491) );
  XOR U20752 ( .A(n20492), .B(n20491), .Z(n20494) );
  NANDN U20753 ( .A(n20207), .B(n20206), .Z(n20211) );
  NAND U20754 ( .A(n20209), .B(n20208), .Z(n20210) );
  AND U20755 ( .A(n20211), .B(n20210), .Z(n20345) );
  AND U20756 ( .A(x[226]), .B(y[2008]), .Z(n20360) );
  XOR U20757 ( .A(n20361), .B(n20360), .Z(n20363) );
  AND U20758 ( .A(x[248]), .B(y[1986]), .Z(n20362) );
  XOR U20759 ( .A(n20363), .B(n20362), .Z(n20397) );
  NANDN U20760 ( .A(n20213), .B(n20212), .Z(n20217) );
  NANDN U20761 ( .A(n20215), .B(n20214), .Z(n20216) );
  AND U20762 ( .A(n20217), .B(n20216), .Z(n20396) );
  XOR U20763 ( .A(n20397), .B(n20396), .Z(n20399) );
  NANDN U20764 ( .A(n20219), .B(n20218), .Z(n20223) );
  NANDN U20765 ( .A(n20221), .B(n20220), .Z(n20222) );
  AND U20766 ( .A(n20223), .B(n20222), .Z(n20398) );
  XOR U20767 ( .A(n20399), .B(n20398), .Z(n20441) );
  NAND U20768 ( .A(n20225), .B(n20224), .Z(n20229) );
  NANDN U20769 ( .A(n20227), .B(n20226), .Z(n20228) );
  AND U20770 ( .A(n20229), .B(n20228), .Z(n20440) );
  NANDN U20771 ( .A(n20231), .B(n20230), .Z(n20235) );
  NAND U20772 ( .A(n20233), .B(n20232), .Z(n20234) );
  AND U20773 ( .A(n20235), .B(n20234), .Z(n20442) );
  XOR U20774 ( .A(n20443), .B(n20442), .Z(n20437) );
  NANDN U20775 ( .A(n20237), .B(n20236), .Z(n20241) );
  NAND U20776 ( .A(n20239), .B(n20238), .Z(n20240) );
  NAND U20777 ( .A(n20241), .B(n20240), .Z(n20434) );
  NANDN U20778 ( .A(n20243), .B(n20242), .Z(n20247) );
  NAND U20779 ( .A(n20245), .B(n20244), .Z(n20246) );
  AND U20780 ( .A(n20247), .B(n20246), .Z(n20435) );
  XOR U20781 ( .A(n20434), .B(n20435), .Z(n20436) );
  XOR U20782 ( .A(n20437), .B(n20436), .Z(n20343) );
  NANDN U20783 ( .A(n20249), .B(n20248), .Z(n20253) );
  NANDN U20784 ( .A(n20251), .B(n20250), .Z(n20252) );
  NAND U20785 ( .A(n20253), .B(n20252), .Z(n20430) );
  AND U20786 ( .A(x[236]), .B(y[1998]), .Z(n20548) );
  AND U20787 ( .A(x[229]), .B(y[2005]), .Z(n20411) );
  XOR U20788 ( .A(n20548), .B(n20411), .Z(n20413) );
  AND U20789 ( .A(x[234]), .B(y[2000]), .Z(n20412) );
  XOR U20790 ( .A(n20413), .B(n20412), .Z(n20449) );
  AND U20791 ( .A(x[231]), .B(y[2003]), .Z(n20447) );
  AND U20792 ( .A(y[2004]), .B(x[230]), .Z(n20255) );
  NAND U20793 ( .A(y[2002]), .B(x[232]), .Z(n20254) );
  XNOR U20794 ( .A(n20255), .B(n20254), .Z(n20466) );
  AND U20795 ( .A(x[233]), .B(y[2001]), .Z(n20465) );
  XOR U20796 ( .A(n20466), .B(n20465), .Z(n20446) );
  XOR U20797 ( .A(n20447), .B(n20446), .Z(n20448) );
  XOR U20798 ( .A(n20449), .B(n20448), .Z(n20386) );
  NANDN U20799 ( .A(n20257), .B(n20256), .Z(n20261) );
  NANDN U20800 ( .A(n20259), .B(n20258), .Z(n20260) );
  NAND U20801 ( .A(n20261), .B(n20260), .Z(n20385) );
  NANDN U20802 ( .A(n20263), .B(n20262), .Z(n20267) );
  NANDN U20803 ( .A(n20265), .B(n20264), .Z(n20266) );
  NAND U20804 ( .A(n20267), .B(n20266), .Z(n20384) );
  XNOR U20805 ( .A(n20385), .B(n20384), .Z(n20387) );
  NAND U20806 ( .A(n20269), .B(n20268), .Z(n20273) );
  NANDN U20807 ( .A(n20271), .B(n20270), .Z(n20272) );
  AND U20808 ( .A(n20273), .B(n20272), .Z(n20422) );
  NAND U20809 ( .A(n20275), .B(n20274), .Z(n20279) );
  NAND U20810 ( .A(n20277), .B(n20276), .Z(n20278) );
  AND U20811 ( .A(n20279), .B(n20278), .Z(n20349) );
  NAND U20812 ( .A(n20281), .B(n20280), .Z(n20285) );
  NAND U20813 ( .A(n20283), .B(n20282), .Z(n20284) );
  AND U20814 ( .A(n20285), .B(n20284), .Z(n20348) );
  XOR U20815 ( .A(n20349), .B(n20348), .Z(n20351) );
  AND U20816 ( .A(n20286), .B(o[217]), .Z(n20459) );
  AND U20817 ( .A(x[238]), .B(y[1996]), .Z(n20458) );
  XOR U20818 ( .A(n20459), .B(n20458), .Z(n20461) );
  AND U20819 ( .A(x[225]), .B(y[2009]), .Z(n20460) );
  XOR U20820 ( .A(n20461), .B(n20460), .Z(n20403) );
  AND U20821 ( .A(x[249]), .B(y[1985]), .Z(n20469) );
  XOR U20822 ( .A(o[218]), .B(n20469), .Z(n20417) );
  AND U20823 ( .A(x[250]), .B(y[1984]), .Z(n20416) );
  XOR U20824 ( .A(n20417), .B(n20416), .Z(n20419) );
  AND U20825 ( .A(x[224]), .B(y[2010]), .Z(n20418) );
  XOR U20826 ( .A(n20419), .B(n20418), .Z(n20402) );
  XOR U20827 ( .A(n20403), .B(n20402), .Z(n20405) );
  NAND U20828 ( .A(n20288), .B(n20287), .Z(n20292) );
  NANDN U20829 ( .A(n20290), .B(n20289), .Z(n20291) );
  AND U20830 ( .A(n20292), .B(n20291), .Z(n20404) );
  XOR U20831 ( .A(n20405), .B(n20404), .Z(n20350) );
  XNOR U20832 ( .A(n20351), .B(n20350), .Z(n20392) );
  NAND U20833 ( .A(x[245]), .B(y[1989]), .Z(n20452) );
  NANDN U20834 ( .A(n20452), .B(n20293), .Z(n20297) );
  NAND U20835 ( .A(n20295), .B(n20294), .Z(n20296) );
  NAND U20836 ( .A(n20297), .B(n20296), .Z(n20380) );
  AND U20837 ( .A(x[244]), .B(y[1990]), .Z(n20454) );
  XOR U20838 ( .A(n20455), .B(n20454), .Z(n20379) );
  AND U20839 ( .A(x[247]), .B(y[1987]), .Z(n20366) );
  XOR U20840 ( .A(n20367), .B(n20366), .Z(n20369) );
  AND U20841 ( .A(x[246]), .B(y[1988]), .Z(n20368) );
  XOR U20842 ( .A(n20369), .B(n20368), .Z(n20378) );
  XOR U20843 ( .A(n20379), .B(n20378), .Z(n20381) );
  XOR U20844 ( .A(n20380), .B(n20381), .Z(n20391) );
  AND U20845 ( .A(x[228]), .B(y[2006]), .Z(n20372) );
  XOR U20846 ( .A(n20373), .B(n20372), .Z(n20374) );
  XOR U20847 ( .A(n20374), .B(n20298), .Z(n20355) );
  AND U20848 ( .A(x[243]), .B(y[1991]), .Z(n20471) );
  AND U20849 ( .A(x[227]), .B(y[2007]), .Z(n20470) );
  XOR U20850 ( .A(n20471), .B(n20470), .Z(n20473) );
  AND U20851 ( .A(x[235]), .B(y[1999]), .Z(n20472) );
  XOR U20852 ( .A(n20473), .B(n20472), .Z(n20354) );
  XOR U20853 ( .A(n20355), .B(n20354), .Z(n20357) );
  NAND U20854 ( .A(n20300), .B(n20299), .Z(n20304) );
  NAND U20855 ( .A(n20302), .B(n20301), .Z(n20303) );
  AND U20856 ( .A(n20304), .B(n20303), .Z(n20356) );
  XNOR U20857 ( .A(n20357), .B(n20356), .Z(n20390) );
  XOR U20858 ( .A(n20392), .B(n20393), .Z(n20425) );
  XNOR U20859 ( .A(n20424), .B(n20425), .Z(n20429) );
  NANDN U20860 ( .A(n20306), .B(n20305), .Z(n20310) );
  NANDN U20861 ( .A(n20308), .B(n20307), .Z(n20309) );
  NAND U20862 ( .A(n20310), .B(n20309), .Z(n20480) );
  NANDN U20863 ( .A(n20312), .B(n20311), .Z(n20316) );
  NAND U20864 ( .A(n20314), .B(n20313), .Z(n20315) );
  NAND U20865 ( .A(n20316), .B(n20315), .Z(n20479) );
  NANDN U20866 ( .A(n20318), .B(n20317), .Z(n20322) );
  NANDN U20867 ( .A(n20320), .B(n20319), .Z(n20321) );
  NAND U20868 ( .A(n20322), .B(n20321), .Z(n20478) );
  XOR U20869 ( .A(n20479), .B(n20478), .Z(n20481) );
  XOR U20870 ( .A(n20480), .B(n20481), .Z(n20428) );
  XOR U20871 ( .A(n20430), .B(n20431), .Z(n20342) );
  NANDN U20872 ( .A(n20324), .B(n20323), .Z(n20328) );
  NANDN U20873 ( .A(n20326), .B(n20325), .Z(n20327) );
  AND U20874 ( .A(n20328), .B(n20327), .Z(n20336) );
  NANDN U20875 ( .A(n20330), .B(n20329), .Z(n20334) );
  NANDN U20876 ( .A(n20332), .B(n20331), .Z(n20333) );
  NAND U20877 ( .A(n20334), .B(n20333), .Z(n20337) );
  XOR U20878 ( .A(n20339), .B(n20338), .Z(n20493) );
  XOR U20879 ( .A(n20494), .B(n20493), .Z(n20487) );
  XNOR U20880 ( .A(n20485), .B(n20487), .Z(n20335) );
  XOR U20881 ( .A(n20484), .B(n20335), .Z(N443) );
  NANDN U20882 ( .A(n20337), .B(n20336), .Z(n20341) );
  NAND U20883 ( .A(n20339), .B(n20338), .Z(n20340) );
  AND U20884 ( .A(n20341), .B(n20340), .Z(n20633) );
  NANDN U20885 ( .A(n20343), .B(n20342), .Z(n20347) );
  NANDN U20886 ( .A(n20345), .B(n20344), .Z(n20346) );
  AND U20887 ( .A(n20347), .B(n20346), .Z(n20631) );
  NAND U20888 ( .A(n20349), .B(n20348), .Z(n20353) );
  NAND U20889 ( .A(n20351), .B(n20350), .Z(n20352) );
  NAND U20890 ( .A(n20353), .B(n20352), .Z(n20608) );
  NAND U20891 ( .A(n20355), .B(n20354), .Z(n20359) );
  NAND U20892 ( .A(n20357), .B(n20356), .Z(n20358) );
  NAND U20893 ( .A(n20359), .B(n20358), .Z(n20606) );
  AND U20894 ( .A(n20361), .B(n20360), .Z(n20365) );
  NAND U20895 ( .A(n20363), .B(n20362), .Z(n20364) );
  NANDN U20896 ( .A(n20365), .B(n20364), .Z(n20523) );
  NAND U20897 ( .A(n20367), .B(n20366), .Z(n20371) );
  NAND U20898 ( .A(n20369), .B(n20368), .Z(n20370) );
  NAND U20899 ( .A(n20371), .B(n20370), .Z(n20522) );
  XOR U20900 ( .A(n20523), .B(n20522), .Z(n20524) );
  AND U20901 ( .A(n20373), .B(n20372), .Z(n20377) );
  NANDN U20902 ( .A(n20375), .B(n20374), .Z(n20376) );
  NANDN U20903 ( .A(n20377), .B(n20376), .Z(n20536) );
  AND U20904 ( .A(x[224]), .B(y[2011]), .Z(n20590) );
  AND U20905 ( .A(x[251]), .B(y[1984]), .Z(n20589) );
  XOR U20906 ( .A(n20590), .B(n20589), .Z(n20592) );
  AND U20907 ( .A(x[250]), .B(y[1985]), .Z(n20593) );
  XOR U20908 ( .A(n20593), .B(o[219]), .Z(n20591) );
  XOR U20909 ( .A(n20592), .B(n20591), .Z(n20535) );
  AND U20910 ( .A(x[233]), .B(y[2002]), .Z(n20597) );
  AND U20911 ( .A(x[245]), .B(y[1990]), .Z(n20596) );
  XOR U20912 ( .A(n20597), .B(n20596), .Z(n20599) );
  AND U20913 ( .A(x[242]), .B(y[1993]), .Z(n20598) );
  XOR U20914 ( .A(n20599), .B(n20598), .Z(n20534) );
  XOR U20915 ( .A(n20535), .B(n20534), .Z(n20537) );
  XNOR U20916 ( .A(n20536), .B(n20537), .Z(n20525) );
  XOR U20917 ( .A(n20606), .B(n20607), .Z(n20609) );
  XOR U20918 ( .A(n20608), .B(n20609), .Z(n20627) );
  NAND U20919 ( .A(n20379), .B(n20378), .Z(n20383) );
  NAND U20920 ( .A(n20381), .B(n20380), .Z(n20382) );
  AND U20921 ( .A(n20383), .B(n20382), .Z(n20625) );
  NAND U20922 ( .A(n20385), .B(n20384), .Z(n20389) );
  NANDN U20923 ( .A(n20387), .B(n20386), .Z(n20388) );
  AND U20924 ( .A(n20389), .B(n20388), .Z(n20624) );
  XOR U20925 ( .A(n20625), .B(n20624), .Z(n20626) );
  NANDN U20926 ( .A(n20391), .B(n20390), .Z(n20395) );
  NANDN U20927 ( .A(n20393), .B(n20392), .Z(n20394) );
  AND U20928 ( .A(n20395), .B(n20394), .Z(n20612) );
  NAND U20929 ( .A(n20397), .B(n20396), .Z(n20401) );
  NAND U20930 ( .A(n20399), .B(n20398), .Z(n20400) );
  NAND U20931 ( .A(n20401), .B(n20400), .Z(n20602) );
  NAND U20932 ( .A(n20403), .B(n20402), .Z(n20407) );
  NAND U20933 ( .A(n20405), .B(n20404), .Z(n20406) );
  NAND U20934 ( .A(n20407), .B(n20406), .Z(n20600) );
  AND U20935 ( .A(x[230]), .B(y[2005]), .Z(n20584) );
  AND U20936 ( .A(x[249]), .B(y[1986]), .Z(n20582) );
  AND U20937 ( .A(x[243]), .B(y[1992]), .Z(n20581) );
  XOR U20938 ( .A(n20582), .B(n20581), .Z(n20583) );
  XOR U20939 ( .A(n20584), .B(n20583), .Z(n20574) );
  AND U20940 ( .A(x[239]), .B(y[1996]), .Z(n20554) );
  AND U20941 ( .A(x[226]), .B(y[2009]), .Z(n20553) );
  XOR U20942 ( .A(n20554), .B(n20553), .Z(n20556) );
  AND U20943 ( .A(x[227]), .B(y[2008]), .Z(n20555) );
  XOR U20944 ( .A(n20556), .B(n20555), .Z(n20573) );
  XOR U20945 ( .A(n20574), .B(n20573), .Z(n20575) );
  NAND U20946 ( .A(x[240]), .B(y[1995]), .Z(n20540) );
  XOR U20947 ( .A(n20540), .B(n20408), .Z(n20543) );
  XOR U20948 ( .A(n20542), .B(n20543), .Z(n20550) );
  AND U20949 ( .A(y[1998]), .B(x[237]), .Z(n20410) );
  AND U20950 ( .A(y[1999]), .B(x[236]), .Z(n20409) );
  XOR U20951 ( .A(n20410), .B(n20409), .Z(n20549) );
  XOR U20952 ( .A(n20550), .B(n20549), .Z(n20576) );
  AND U20953 ( .A(n20548), .B(n20411), .Z(n20415) );
  NAND U20954 ( .A(n20413), .B(n20412), .Z(n20414) );
  NANDN U20955 ( .A(n20415), .B(n20414), .Z(n20517) );
  NAND U20956 ( .A(n20417), .B(n20416), .Z(n20421) );
  NAND U20957 ( .A(n20419), .B(n20418), .Z(n20420) );
  NAND U20958 ( .A(n20421), .B(n20420), .Z(n20516) );
  XOR U20959 ( .A(n20517), .B(n20516), .Z(n20518) );
  XOR U20960 ( .A(n20519), .B(n20518), .Z(n20601) );
  XNOR U20961 ( .A(n20600), .B(n20601), .Z(n20603) );
  XNOR U20962 ( .A(n20612), .B(n20613), .Z(n20615) );
  NANDN U20963 ( .A(n20423), .B(n20422), .Z(n20427) );
  NANDN U20964 ( .A(n20425), .B(n20424), .Z(n20426) );
  AND U20965 ( .A(n20427), .B(n20426), .Z(n20614) );
  XOR U20966 ( .A(n20615), .B(n20614), .Z(n20498) );
  NANDN U20967 ( .A(n20429), .B(n20428), .Z(n20433) );
  NAND U20968 ( .A(n20431), .B(n20430), .Z(n20432) );
  NAND U20969 ( .A(n20433), .B(n20432), .Z(n20500) );
  XOR U20970 ( .A(n20501), .B(n20500), .Z(n20507) );
  NAND U20971 ( .A(n20435), .B(n20434), .Z(n20439) );
  NAND U20972 ( .A(n20437), .B(n20436), .Z(n20438) );
  NAND U20973 ( .A(n20439), .B(n20438), .Z(n20504) );
  NANDN U20974 ( .A(n20441), .B(n20440), .Z(n20445) );
  NAND U20975 ( .A(n20443), .B(n20442), .Z(n20444) );
  NAND U20976 ( .A(n20445), .B(n20444), .Z(n20511) );
  NAND U20977 ( .A(n20447), .B(n20446), .Z(n20451) );
  NAND U20978 ( .A(n20449), .B(n20448), .Z(n20450) );
  NAND U20979 ( .A(n20451), .B(n20450), .Z(n20620) );
  ANDN U20980 ( .B(n20453), .A(n20452), .Z(n20457) );
  NAND U20981 ( .A(n20455), .B(n20454), .Z(n20456) );
  NANDN U20982 ( .A(n20457), .B(n20456), .Z(n20562) );
  NAND U20983 ( .A(n20459), .B(n20458), .Z(n20463) );
  NAND U20984 ( .A(n20461), .B(n20460), .Z(n20462) );
  NAND U20985 ( .A(n20463), .B(n20462), .Z(n20561) );
  XOR U20986 ( .A(n20562), .B(n20561), .Z(n20563) );
  AND U20987 ( .A(x[232]), .B(y[2004]), .Z(n20595) );
  NAND U20988 ( .A(n20464), .B(n20595), .Z(n20468) );
  NAND U20989 ( .A(n20466), .B(n20465), .Z(n20467) );
  NAND U20990 ( .A(n20468), .B(n20467), .Z(n20530) );
  AND U20991 ( .A(x[225]), .B(y[2010]), .Z(n20558) );
  AND U20992 ( .A(x[238]), .B(y[1997]), .Z(n20557) );
  XOR U20993 ( .A(n20558), .B(n20557), .Z(n20559) );
  XOR U20994 ( .A(n20560), .B(n20559), .Z(n20529) );
  AND U20995 ( .A(x[241]), .B(y[1994]), .Z(n20586) );
  AND U20996 ( .A(x[228]), .B(y[2007]), .Z(n20585) );
  XOR U20997 ( .A(n20586), .B(n20585), .Z(n20588) );
  AND U20998 ( .A(x[229]), .B(y[2006]), .Z(n20587) );
  XOR U20999 ( .A(n20588), .B(n20587), .Z(n20528) );
  XOR U21000 ( .A(n20529), .B(n20528), .Z(n20531) );
  XNOR U21001 ( .A(n20530), .B(n20531), .Z(n20564) );
  NAND U21002 ( .A(n20471), .B(n20470), .Z(n20475) );
  NAND U21003 ( .A(n20473), .B(n20472), .Z(n20474) );
  NAND U21004 ( .A(n20475), .B(n20474), .Z(n20569) );
  AND U21005 ( .A(x[231]), .B(y[2004]), .Z(n20580) );
  AND U21006 ( .A(y[1987]), .B(x[248]), .Z(n20477) );
  XOR U21007 ( .A(n20477), .B(n20476), .Z(n20579) );
  XOR U21008 ( .A(n20580), .B(n20579), .Z(n20568) );
  AND U21009 ( .A(x[246]), .B(y[1989]), .Z(n20547) );
  AND U21010 ( .A(x[232]), .B(y[2003]), .Z(n20545) );
  AND U21011 ( .A(x[247]), .B(y[1988]), .Z(n20544) );
  XOR U21012 ( .A(n20545), .B(n20544), .Z(n20546) );
  XOR U21013 ( .A(n20547), .B(n20546), .Z(n20567) );
  XOR U21014 ( .A(n20568), .B(n20567), .Z(n20570) );
  XOR U21015 ( .A(n20569), .B(n20570), .Z(n20618) );
  XOR U21016 ( .A(n20619), .B(n20618), .Z(n20621) );
  XNOR U21017 ( .A(n20620), .B(n20621), .Z(n20510) );
  XOR U21018 ( .A(n20511), .B(n20510), .Z(n20513) );
  NAND U21019 ( .A(n20479), .B(n20478), .Z(n20483) );
  NAND U21020 ( .A(n20481), .B(n20480), .Z(n20482) );
  AND U21021 ( .A(n20483), .B(n20482), .Z(n20512) );
  XOR U21022 ( .A(n20513), .B(n20512), .Z(n20505) );
  XOR U21023 ( .A(n20504), .B(n20505), .Z(n20506) );
  XOR U21024 ( .A(n20631), .B(n20630), .Z(n20632) );
  XNOR U21025 ( .A(n20633), .B(n20632), .Z(n20638) );
  NANDN U21026 ( .A(n20484), .B(n20485), .Z(n20490) );
  NOR U21027 ( .A(n20486), .B(n20485), .Z(n20488) );
  OR U21028 ( .A(n20488), .B(n20487), .Z(n20489) );
  AND U21029 ( .A(n20490), .B(n20489), .Z(n20637) );
  NAND U21030 ( .A(n20492), .B(n20491), .Z(n20496) );
  NAND U21031 ( .A(n20494), .B(n20493), .Z(n20495) );
  AND U21032 ( .A(n20496), .B(n20495), .Z(n20636) );
  XOR U21033 ( .A(n20637), .B(n20636), .Z(n20497) );
  XNOR U21034 ( .A(n20638), .B(n20497), .Z(N444) );
  NANDN U21035 ( .A(n20499), .B(n20498), .Z(n20503) );
  NAND U21036 ( .A(n20501), .B(n20500), .Z(n20502) );
  NAND U21037 ( .A(n20503), .B(n20502), .Z(n20640) );
  NAND U21038 ( .A(n20505), .B(n20504), .Z(n20509) );
  NANDN U21039 ( .A(n20507), .B(n20506), .Z(n20508) );
  AND U21040 ( .A(n20509), .B(n20508), .Z(n20641) );
  XOR U21041 ( .A(n20640), .B(n20641), .Z(n20643) );
  NAND U21042 ( .A(n20511), .B(n20510), .Z(n20515) );
  NAND U21043 ( .A(n20513), .B(n20512), .Z(n20514) );
  AND U21044 ( .A(n20515), .B(n20514), .Z(n20649) );
  NAND U21045 ( .A(n20517), .B(n20516), .Z(n20521) );
  NAND U21046 ( .A(n20519), .B(n20518), .Z(n20520) );
  NAND U21047 ( .A(n20521), .B(n20520), .Z(n20661) );
  NAND U21048 ( .A(n20523), .B(n20522), .Z(n20527) );
  NANDN U21049 ( .A(n20525), .B(n20524), .Z(n20526) );
  NAND U21050 ( .A(n20527), .B(n20526), .Z(n20744) );
  NAND U21051 ( .A(n20529), .B(n20528), .Z(n20533) );
  NAND U21052 ( .A(n20531), .B(n20530), .Z(n20532) );
  NAND U21053 ( .A(n20533), .B(n20532), .Z(n20743) );
  NAND U21054 ( .A(n20535), .B(n20534), .Z(n20539) );
  NAND U21055 ( .A(n20537), .B(n20536), .Z(n20538) );
  NAND U21056 ( .A(n20539), .B(n20538), .Z(n20742) );
  XOR U21057 ( .A(n20743), .B(n20742), .Z(n20745) );
  XOR U21058 ( .A(n20744), .B(n20745), .Z(n20662) );
  XOR U21059 ( .A(n20661), .B(n20662), .Z(n20664) );
  AND U21060 ( .A(x[239]), .B(y[1997]), .Z(n20720) );
  NAND U21061 ( .A(x[251]), .B(y[1985]), .Z(n20707) );
  XNOR U21062 ( .A(o[220]), .B(n20707), .Z(n20718) );
  AND U21063 ( .A(x[250]), .B(y[1986]), .Z(n20717) );
  XOR U21064 ( .A(n20718), .B(n20717), .Z(n20719) );
  XOR U21065 ( .A(n20720), .B(n20719), .Z(n20710) );
  AND U21066 ( .A(x[231]), .B(y[2005]), .Z(n20697) );
  AND U21067 ( .A(x[236]), .B(y[2000]), .Z(n20696) );
  XOR U21068 ( .A(n20697), .B(n20696), .Z(n20699) );
  AND U21069 ( .A(x[235]), .B(y[2001]), .Z(n20698) );
  XNOR U21070 ( .A(n20699), .B(n20698), .Z(n20709) );
  XNOR U21071 ( .A(n20710), .B(n20709), .Z(n20712) );
  XOR U21072 ( .A(n20711), .B(n20712), .Z(n20749) );
  AND U21073 ( .A(x[241]), .B(y[1995]), .Z(n20672) );
  AND U21074 ( .A(x[246]), .B(y[1990]), .Z(n20671) );
  XOR U21075 ( .A(n20672), .B(n20671), .Z(n20674) );
  AND U21076 ( .A(x[228]), .B(y[2008]), .Z(n20673) );
  XOR U21077 ( .A(n20674), .B(n20673), .Z(n20727) );
  AND U21078 ( .A(x[230]), .B(y[2006]), .Z(n20865) );
  AND U21079 ( .A(x[243]), .B(y[1993]), .Z(n20700) );
  XOR U21080 ( .A(n20865), .B(n20700), .Z(n20702) );
  XOR U21081 ( .A(n20702), .B(n20701), .Z(n20726) );
  XOR U21082 ( .A(n20727), .B(n20726), .Z(n20729) );
  XOR U21083 ( .A(n20728), .B(n20729), .Z(n20748) );
  NAND U21084 ( .A(n20548), .B(n20714), .Z(n20552) );
  NANDN U21085 ( .A(n20550), .B(n20549), .Z(n20551) );
  NAND U21086 ( .A(n20552), .B(n20551), .Z(n20686) );
  XOR U21087 ( .A(n20684), .B(n20685), .Z(n20687) );
  XOR U21088 ( .A(n20686), .B(n20687), .Z(n20750) );
  XOR U21089 ( .A(n20751), .B(n20750), .Z(n20663) );
  XNOR U21090 ( .A(n20664), .B(n20663), .Z(n20769) );
  NAND U21091 ( .A(n20562), .B(n20561), .Z(n20566) );
  NANDN U21092 ( .A(n20564), .B(n20563), .Z(n20565) );
  NAND U21093 ( .A(n20566), .B(n20565), .Z(n20732) );
  NAND U21094 ( .A(n20568), .B(n20567), .Z(n20572) );
  NAND U21095 ( .A(n20570), .B(n20569), .Z(n20571) );
  NAND U21096 ( .A(n20572), .B(n20571), .Z(n20731) );
  NAND U21097 ( .A(n20574), .B(n20573), .Z(n20578) );
  NANDN U21098 ( .A(n20576), .B(n20575), .Z(n20577) );
  NAND U21099 ( .A(n20578), .B(n20577), .Z(n20730) );
  XOR U21100 ( .A(n20731), .B(n20730), .Z(n20733) );
  XOR U21101 ( .A(n20732), .B(n20733), .Z(n20767) );
  AND U21102 ( .A(x[248]), .B(y[1991]), .Z(n20999) );
  AND U21103 ( .A(x[249]), .B(y[1987]), .Z(n20694) );
  XOR U21104 ( .A(n20695), .B(n20694), .Z(n20693) );
  AND U21105 ( .A(x[225]), .B(y[2011]), .Z(n20692) );
  XOR U21106 ( .A(n20693), .B(n20692), .Z(n20763) );
  AND U21107 ( .A(x[240]), .B(y[1996]), .Z(n20689) );
  AND U21108 ( .A(x[248]), .B(y[1988]), .Z(n20688) );
  XOR U21109 ( .A(n20689), .B(n20688), .Z(n20691) );
  AND U21110 ( .A(x[226]), .B(y[2010]), .Z(n20690) );
  XOR U21111 ( .A(n20691), .B(n20690), .Z(n20762) );
  XOR U21112 ( .A(n20763), .B(n20762), .Z(n20765) );
  XOR U21113 ( .A(n20764), .B(n20765), .Z(n20739) );
  AND U21114 ( .A(x[227]), .B(y[2009]), .Z(n20713) );
  XOR U21115 ( .A(n20714), .B(n20713), .Z(n20716) );
  AND U21116 ( .A(x[247]), .B(y[1989]), .Z(n20715) );
  XOR U21117 ( .A(n20716), .B(n20715), .Z(n20759) );
  AND U21118 ( .A(x[229]), .B(y[2007]), .Z(n20704) );
  AND U21119 ( .A(x[245]), .B(y[1991]), .Z(n20703) );
  XOR U21120 ( .A(n20704), .B(n20703), .Z(n20706) );
  AND U21121 ( .A(x[244]), .B(y[1992]), .Z(n20705) );
  XOR U21122 ( .A(n20706), .B(n20705), .Z(n20758) );
  XOR U21123 ( .A(n20759), .B(n20758), .Z(n20761) );
  XOR U21124 ( .A(n20760), .B(n20761), .Z(n20737) );
  XOR U21125 ( .A(n20754), .B(n20755), .Z(n20757) );
  AND U21126 ( .A(n20593), .B(o[219]), .Z(n20678) );
  AND U21127 ( .A(x[224]), .B(y[2012]), .Z(n20676) );
  AND U21128 ( .A(x[252]), .B(y[1984]), .Z(n20675) );
  XOR U21129 ( .A(n20676), .B(n20675), .Z(n20677) );
  XOR U21130 ( .A(n20678), .B(n20677), .Z(n20668) );
  NAND U21131 ( .A(y[2002]), .B(x[234]), .Z(n20594) );
  XNOR U21132 ( .A(n20595), .B(n20594), .Z(n20681) );
  AND U21133 ( .A(x[233]), .B(y[2003]), .Z(n20680) );
  XOR U21134 ( .A(n20681), .B(n20680), .Z(n20667) );
  XOR U21135 ( .A(n20668), .B(n20667), .Z(n20670) );
  XOR U21136 ( .A(n20670), .B(n20669), .Z(n20756) );
  XNOR U21137 ( .A(n20757), .B(n20756), .Z(n20736) );
  XNOR U21138 ( .A(n20769), .B(n20768), .Z(n20774) );
  NAND U21139 ( .A(n20601), .B(n20600), .Z(n20605) );
  NANDN U21140 ( .A(n20603), .B(n20602), .Z(n20604) );
  NAND U21141 ( .A(n20605), .B(n20604), .Z(n20773) );
  NAND U21142 ( .A(n20607), .B(n20606), .Z(n20611) );
  NAND U21143 ( .A(n20609), .B(n20608), .Z(n20610) );
  NAND U21144 ( .A(n20611), .B(n20610), .Z(n20772) );
  XNOR U21145 ( .A(n20773), .B(n20772), .Z(n20775) );
  XNOR U21146 ( .A(n20649), .B(n20650), .Z(n20652) );
  NANDN U21147 ( .A(n20613), .B(n20612), .Z(n20617) );
  NAND U21148 ( .A(n20615), .B(n20614), .Z(n20616) );
  NAND U21149 ( .A(n20617), .B(n20616), .Z(n20657) );
  NAND U21150 ( .A(n20619), .B(n20618), .Z(n20623) );
  NAND U21151 ( .A(n20621), .B(n20620), .Z(n20622) );
  NAND U21152 ( .A(n20623), .B(n20622), .Z(n20655) );
  NAND U21153 ( .A(n20625), .B(n20624), .Z(n20629) );
  NANDN U21154 ( .A(n20627), .B(n20626), .Z(n20628) );
  AND U21155 ( .A(n20629), .B(n20628), .Z(n20656) );
  XOR U21156 ( .A(n20655), .B(n20656), .Z(n20658) );
  XOR U21157 ( .A(n20657), .B(n20658), .Z(n20651) );
  XOR U21158 ( .A(n20652), .B(n20651), .Z(n20642) );
  XOR U21159 ( .A(n20643), .B(n20642), .Z(n20648) );
  NAND U21160 ( .A(n20631), .B(n20630), .Z(n20635) );
  NAND U21161 ( .A(n20633), .B(n20632), .Z(n20634) );
  NAND U21162 ( .A(n20635), .B(n20634), .Z(n20646) );
  XOR U21163 ( .A(n20646), .B(n20647), .Z(n20639) );
  XNOR U21164 ( .A(n20648), .B(n20639), .Z(N445) );
  NAND U21165 ( .A(n20641), .B(n20640), .Z(n20645) );
  NAND U21166 ( .A(n20643), .B(n20642), .Z(n20644) );
  AND U21167 ( .A(n20645), .B(n20644), .Z(n20780) );
  NANDN U21168 ( .A(n20650), .B(n20649), .Z(n20654) );
  NAND U21169 ( .A(n20652), .B(n20651), .Z(n20653) );
  NAND U21170 ( .A(n20654), .B(n20653), .Z(n20788) );
  NAND U21171 ( .A(n20656), .B(n20655), .Z(n20660) );
  NAND U21172 ( .A(n20658), .B(n20657), .Z(n20659) );
  NAND U21173 ( .A(n20660), .B(n20659), .Z(n20787) );
  NAND U21174 ( .A(n20662), .B(n20661), .Z(n20666) );
  NAND U21175 ( .A(n20664), .B(n20663), .Z(n20665) );
  NAND U21176 ( .A(n20666), .B(n20665), .Z(n20804) );
  XOR U21177 ( .A(n20935), .B(n20936), .Z(n20937) );
  AND U21178 ( .A(x[234]), .B(y[2004]), .Z(n20933) );
  NAND U21179 ( .A(n20679), .B(n20933), .Z(n20683) );
  NAND U21180 ( .A(n20681), .B(n20680), .Z(n20682) );
  NAND U21181 ( .A(n20683), .B(n20682), .Z(n20911) );
  AND U21182 ( .A(x[246]), .B(y[1991]), .Z(n20886) );
  AND U21183 ( .A(x[236]), .B(y[2001]), .Z(n20986) );
  AND U21184 ( .A(x[225]), .B(y[2012]), .Z(n20884) );
  XOR U21185 ( .A(n20986), .B(n20884), .Z(n20885) );
  XOR U21186 ( .A(n20886), .B(n20885), .Z(n20910) );
  AND U21187 ( .A(x[239]), .B(y[1998]), .Z(n20887) );
  XOR U21188 ( .A(n20910), .B(n20909), .Z(n20912) );
  XNOR U21189 ( .A(n20911), .B(n20912), .Z(n20938) );
  XOR U21190 ( .A(n20937), .B(n20938), .Z(n20905) );
  XOR U21191 ( .A(n20906), .B(n20905), .Z(n20908) );
  XOR U21192 ( .A(n20908), .B(n20907), .Z(n20904) );
  XOR U21193 ( .A(n20915), .B(n20916), .Z(n20917) );
  AND U21194 ( .A(x[235]), .B(y[2002]), .Z(n20861) );
  AND U21195 ( .A(x[227]), .B(y[2010]), .Z(n20859) );
  AND U21196 ( .A(x[241]), .B(y[1996]), .Z(n20858) );
  XOR U21197 ( .A(n20859), .B(n20858), .Z(n20860) );
  XOR U21198 ( .A(n20861), .B(n20860), .Z(n20827) );
  AND U21199 ( .A(x[247]), .B(y[1990]), .Z(n20855) );
  AND U21200 ( .A(x[237]), .B(y[2000]), .Z(n20853) );
  AND U21201 ( .A(x[248]), .B(y[1989]), .Z(n21124) );
  XOR U21202 ( .A(n20853), .B(n21124), .Z(n20854) );
  XOR U21203 ( .A(n20855), .B(n20854), .Z(n20826) );
  XOR U21204 ( .A(n20827), .B(n20826), .Z(n20828) );
  XNOR U21205 ( .A(n20829), .B(n20828), .Z(n20918) );
  XOR U21206 ( .A(n20917), .B(n20918), .Z(n20818) );
  AND U21207 ( .A(x[249]), .B(y[1988]), .Z(n20883) );
  AND U21208 ( .A(x[250]), .B(y[1987]), .Z(n20880) );
  XOR U21209 ( .A(n20881), .B(n20880), .Z(n20882) );
  XOR U21210 ( .A(n20883), .B(n20882), .Z(n20920) );
  AND U21211 ( .A(x[252]), .B(y[1985]), .Z(n20894) );
  XOR U21212 ( .A(o[221]), .B(n20894), .Z(n20930) );
  AND U21213 ( .A(x[224]), .B(y[2013]), .Z(n20928) );
  AND U21214 ( .A(x[253]), .B(y[1984]), .Z(n20927) );
  XOR U21215 ( .A(n20928), .B(n20927), .Z(n20929) );
  XOR U21216 ( .A(n20930), .B(n20929), .Z(n20919) );
  XOR U21217 ( .A(n20920), .B(n20919), .Z(n20921) );
  XOR U21218 ( .A(n20922), .B(n20921), .Z(n20816) );
  ANDN U21219 ( .B(o[220]), .A(n20707), .Z(n20833) );
  AND U21220 ( .A(x[240]), .B(y[1997]), .Z(n20831) );
  AND U21221 ( .A(x[251]), .B(y[1986]), .Z(n20830) );
  XOR U21222 ( .A(n20831), .B(n20830), .Z(n20832) );
  XOR U21223 ( .A(n20833), .B(n20832), .Z(n20873) );
  AND U21224 ( .A(x[226]), .B(y[2011]), .Z(n20840) );
  XOR U21225 ( .A(n20843), .B(n20842), .Z(n20872) );
  XOR U21226 ( .A(n20873), .B(n20872), .Z(n20876) );
  XOR U21227 ( .A(n20875), .B(n20876), .Z(n20817) );
  IV U21228 ( .A(n20817), .Z(n20708) );
  XOR U21229 ( .A(n20816), .B(n20708), .Z(n20819) );
  XOR U21230 ( .A(n20818), .B(n20819), .Z(n20824) );
  NAND U21231 ( .A(n20718), .B(n20717), .Z(n20723) );
  IV U21232 ( .A(n20719), .Z(n20721) );
  NANDN U21233 ( .A(n20721), .B(n20720), .Z(n20722) );
  NAND U21234 ( .A(n20723), .B(n20722), .Z(n20847) );
  XOR U21235 ( .A(n20846), .B(n20847), .Z(n20849) );
  AND U21236 ( .A(x[232]), .B(y[2005]), .Z(n20867) );
  AND U21237 ( .A(y[2007]), .B(x[230]), .Z(n20725) );
  NAND U21238 ( .A(y[2006]), .B(x[231]), .Z(n20724) );
  XNOR U21239 ( .A(n20725), .B(n20724), .Z(n20866) );
  XNOR U21240 ( .A(n20867), .B(n20866), .Z(n20925) );
  AND U21241 ( .A(x[229]), .B(y[2008]), .Z(n20836) );
  AND U21242 ( .A(x[228]), .B(y[2009]), .Z(n20835) );
  AND U21243 ( .A(x[234]), .B(y[2003]), .Z(n20834) );
  XNOR U21244 ( .A(n20835), .B(n20834), .Z(n20837) );
  XNOR U21245 ( .A(n20836), .B(n20837), .Z(n20926) );
  AND U21246 ( .A(x[233]), .B(y[2004]), .Z(n20996) );
  XOR U21247 ( .A(n20849), .B(n20850), .Z(n20823) );
  XNOR U21248 ( .A(n20822), .B(n20823), .Z(n20825) );
  XOR U21249 ( .A(n20824), .B(n20825), .Z(n20901) );
  XOR U21250 ( .A(n20901), .B(n20902), .Z(n20903) );
  XNOR U21251 ( .A(n20904), .B(n20903), .Z(n20805) );
  XOR U21252 ( .A(n20804), .B(n20805), .Z(n20807) );
  NAND U21253 ( .A(n20731), .B(n20730), .Z(n20735) );
  NAND U21254 ( .A(n20733), .B(n20732), .Z(n20734) );
  NAND U21255 ( .A(n20735), .B(n20734), .Z(n20798) );
  NANDN U21256 ( .A(n20737), .B(n20736), .Z(n20741) );
  NANDN U21257 ( .A(n20739), .B(n20738), .Z(n20740) );
  AND U21258 ( .A(n20741), .B(n20740), .Z(n20799) );
  XOR U21259 ( .A(n20798), .B(n20799), .Z(n20801) );
  NAND U21260 ( .A(n20743), .B(n20742), .Z(n20747) );
  NAND U21261 ( .A(n20745), .B(n20744), .Z(n20746) );
  NAND U21262 ( .A(n20747), .B(n20746), .Z(n20812) );
  NANDN U21263 ( .A(n20749), .B(n20748), .Z(n20753) );
  NAND U21264 ( .A(n20751), .B(n20750), .Z(n20752) );
  NAND U21265 ( .A(n20753), .B(n20752), .Z(n20810) );
  XOR U21266 ( .A(n20896), .B(n20897), .Z(n20899) );
  XOR U21267 ( .A(n20898), .B(n20899), .Z(n20811) );
  XOR U21268 ( .A(n20810), .B(n20811), .Z(n20813) );
  XOR U21269 ( .A(n20812), .B(n20813), .Z(n20800) );
  XOR U21270 ( .A(n20801), .B(n20800), .Z(n20806) );
  XNOR U21271 ( .A(n20807), .B(n20806), .Z(n20794) );
  NANDN U21272 ( .A(n20767), .B(n20766), .Z(n20771) );
  NAND U21273 ( .A(n20769), .B(n20768), .Z(n20770) );
  NAND U21274 ( .A(n20771), .B(n20770), .Z(n20792) );
  NAND U21275 ( .A(n20773), .B(n20772), .Z(n20777) );
  NANDN U21276 ( .A(n20775), .B(n20774), .Z(n20776) );
  AND U21277 ( .A(n20777), .B(n20776), .Z(n20793) );
  XNOR U21278 ( .A(n20792), .B(n20793), .Z(n20795) );
  XOR U21279 ( .A(n20794), .B(n20795), .Z(n20786) );
  XOR U21280 ( .A(n20787), .B(n20786), .Z(n20789) );
  XOR U21281 ( .A(n20788), .B(n20789), .Z(n20782) );
  XNOR U21282 ( .A(n20781), .B(n20782), .Z(n20778) );
  XOR U21283 ( .A(n20780), .B(n20778), .Z(N446) );
  IV U21284 ( .A(n20780), .Z(n20779) );
  OR U21285 ( .A(n20781), .B(n20779), .Z(n20785) );
  ANDN U21286 ( .B(n20781), .A(n20780), .Z(n20783) );
  OR U21287 ( .A(n20783), .B(n20782), .Z(n20784) );
  AND U21288 ( .A(n20785), .B(n20784), .Z(n21186) );
  NAND U21289 ( .A(n20787), .B(n20786), .Z(n20791) );
  NAND U21290 ( .A(n20789), .B(n20788), .Z(n20790) );
  AND U21291 ( .A(n20791), .B(n20790), .Z(n21185) );
  XNOR U21292 ( .A(n21186), .B(n21185), .Z(n21184) );
  NAND U21293 ( .A(n20793), .B(n20792), .Z(n20797) );
  NANDN U21294 ( .A(n20795), .B(n20794), .Z(n20796) );
  AND U21295 ( .A(n20797), .B(n20796), .Z(n21188) );
  NAND U21296 ( .A(n20799), .B(n20798), .Z(n20803) );
  NAND U21297 ( .A(n20801), .B(n20800), .Z(n20802) );
  AND U21298 ( .A(n20803), .B(n20802), .Z(n21192) );
  NAND U21299 ( .A(n20805), .B(n20804), .Z(n20809) );
  NAND U21300 ( .A(n20807), .B(n20806), .Z(n20808) );
  AND U21301 ( .A(n20809), .B(n20808), .Z(n21191) );
  XOR U21302 ( .A(n21192), .B(n21191), .Z(n21194) );
  NAND U21303 ( .A(n20811), .B(n20810), .Z(n20815) );
  NAND U21304 ( .A(n20813), .B(n20812), .Z(n20814) );
  AND U21305 ( .A(n20815), .B(n20814), .Z(n21193) );
  XOR U21306 ( .A(n21194), .B(n21193), .Z(n21189) );
  IV U21307 ( .A(n21189), .Z(n20939) );
  NANDN U21308 ( .A(n20817), .B(n20816), .Z(n20821) );
  NAND U21309 ( .A(n20819), .B(n20818), .Z(n20820) );
  AND U21310 ( .A(n20821), .B(n20820), .Z(n21180) );
  NAND U21311 ( .A(n20835), .B(n20834), .Z(n20839) );
  NANDN U21312 ( .A(n20837), .B(n20836), .Z(n20838) );
  NAND U21313 ( .A(n20839), .B(n20838), .Z(n20953) );
  AND U21314 ( .A(x[230]), .B(y[2008]), .Z(n21108) );
  AND U21315 ( .A(x[229]), .B(y[2009]), .Z(n21110) );
  AND U21316 ( .A(x[243]), .B(y[1995]), .Z(n21109) );
  XOR U21317 ( .A(n21110), .B(n21109), .Z(n21107) );
  XNOR U21318 ( .A(n21108), .B(n21107), .Z(n21096) );
  AND U21319 ( .A(x[228]), .B(y[2010]), .Z(n21061) );
  AND U21320 ( .A(x[227]), .B(y[2011]), .Z(n21063) );
  AND U21321 ( .A(x[242]), .B(y[1996]), .Z(n21062) );
  XOR U21322 ( .A(n21063), .B(n21062), .Z(n21060) );
  XOR U21323 ( .A(n21061), .B(n21060), .Z(n21093) );
  NANDN U21324 ( .A(n20841), .B(n20840), .Z(n20845) );
  NAND U21325 ( .A(n20843), .B(n20842), .Z(n20844) );
  AND U21326 ( .A(n20845), .B(n20844), .Z(n21094) );
  XOR U21327 ( .A(n21096), .B(n21095), .Z(n20952) );
  XOR U21328 ( .A(n20953), .B(n20952), .Z(n20951) );
  XOR U21329 ( .A(n20950), .B(n20951), .Z(n20942) );
  IV U21330 ( .A(n20846), .Z(n20848) );
  NANDN U21331 ( .A(n20848), .B(n20847), .Z(n20852) );
  NANDN U21332 ( .A(n20850), .B(n20849), .Z(n20851) );
  AND U21333 ( .A(n20852), .B(n20851), .Z(n20940) );
  XOR U21334 ( .A(n20941), .B(n20940), .Z(n21173) );
  IV U21335 ( .A(n21173), .Z(n20895) );
  NAND U21336 ( .A(n20853), .B(n21124), .Z(n20857) );
  NAND U21337 ( .A(n20855), .B(n20854), .Z(n20856) );
  NAND U21338 ( .A(n20857), .B(n20856), .Z(n20947) );
  NAND U21339 ( .A(n20859), .B(n20858), .Z(n20863) );
  NAND U21340 ( .A(n20861), .B(n20860), .Z(n20862) );
  AND U21341 ( .A(n20863), .B(n20862), .Z(n20957) );
  AND U21342 ( .A(x[224]), .B(y[2014]), .Z(n20981) );
  AND U21343 ( .A(x[253]), .B(y[1985]), .Z(n20997) );
  XOR U21344 ( .A(o[222]), .B(n20997), .Z(n20983) );
  AND U21345 ( .A(x[254]), .B(y[1984]), .Z(n20982) );
  XOR U21346 ( .A(n20983), .B(n20982), .Z(n20980) );
  XOR U21347 ( .A(n20981), .B(n20980), .Z(n20959) );
  IV U21348 ( .A(n20959), .Z(n20864) );
  AND U21349 ( .A(x[244]), .B(y[1994]), .Z(n21050) );
  XOR U21350 ( .A(n21051), .B(n21050), .Z(n21049) );
  AND U21351 ( .A(x[232]), .B(y[2006]), .Z(n21048) );
  XNOR U21352 ( .A(n21049), .B(n21048), .Z(n20958) );
  XOR U21353 ( .A(n20864), .B(n20958), .Z(n20956) );
  XNOR U21354 ( .A(n20957), .B(n20956), .Z(n20946) );
  XOR U21355 ( .A(n20947), .B(n20946), .Z(n20944) );
  AND U21356 ( .A(x[231]), .B(y[2007]), .Z(n20988) );
  NAND U21357 ( .A(n20865), .B(n20988), .Z(n20869) );
  NAND U21358 ( .A(n20867), .B(n20866), .Z(n20868) );
  AND U21359 ( .A(n20869), .B(n20868), .Z(n20968) );
  AND U21360 ( .A(y[1993]), .B(x[245]), .Z(n20871) );
  AND U21361 ( .A(y[1992]), .B(x[246]), .Z(n20870) );
  XOR U21362 ( .A(n20871), .B(n20870), .Z(n20987) );
  XOR U21363 ( .A(n20988), .B(n20987), .Z(n20971) );
  AND U21364 ( .A(x[241]), .B(y[1997]), .Z(n21102) );
  AND U21365 ( .A(x[226]), .B(y[2012]), .Z(n21104) );
  AND U21366 ( .A(x[250]), .B(y[1988]), .Z(n21103) );
  XOR U21367 ( .A(n21104), .B(n21103), .Z(n21101) );
  XNOR U21368 ( .A(n21102), .B(n21101), .Z(n20970) );
  XNOR U21369 ( .A(n20968), .B(n20969), .Z(n20945) );
  XNOR U21370 ( .A(n20944), .B(n20945), .Z(n21161) );
  IV U21371 ( .A(n20872), .Z(n20874) );
  NANDN U21372 ( .A(n20874), .B(n20873), .Z(n20879) );
  IV U21373 ( .A(n20875), .Z(n20877) );
  NANDN U21374 ( .A(n20877), .B(n20876), .Z(n20878) );
  NAND U21375 ( .A(n20879), .B(n20878), .Z(n21160) );
  XOR U21376 ( .A(n21161), .B(n21160), .Z(n21159) );
  NANDN U21377 ( .A(n20989), .B(n20887), .Z(n20891) );
  NANDN U21378 ( .A(n20889), .B(n20888), .Z(n20890) );
  AND U21379 ( .A(n20891), .B(n20890), .Z(n20963) );
  AND U21380 ( .A(x[247]), .B(y[1991]), .Z(n21122) );
  AND U21381 ( .A(y[1990]), .B(x[248]), .Z(n20893) );
  AND U21382 ( .A(y[1989]), .B(x[249]), .Z(n20892) );
  XOR U21383 ( .A(n20893), .B(n20892), .Z(n21121) );
  XOR U21384 ( .A(n21122), .B(n21121), .Z(n20965) );
  AND U21385 ( .A(x[252]), .B(y[1986]), .Z(n21118) );
  AND U21386 ( .A(x[240]), .B(y[1998]), .Z(n21117) );
  XOR U21387 ( .A(n21118), .B(n21117), .Z(n21115) );
  XNOR U21388 ( .A(n21116), .B(n21115), .Z(n20964) );
  XNOR U21389 ( .A(n20963), .B(n20962), .Z(n20978) );
  XOR U21390 ( .A(n20979), .B(n20978), .Z(n20977) );
  XOR U21391 ( .A(n20976), .B(n20977), .Z(n21158) );
  XOR U21392 ( .A(n21159), .B(n21158), .Z(n21172) );
  XNOR U21393 ( .A(n20895), .B(n21172), .Z(n21171) );
  XNOR U21394 ( .A(n21170), .B(n21171), .Z(n21178) );
  XOR U21395 ( .A(n21178), .B(n21179), .Z(n20900) );
  XOR U21396 ( .A(n21180), .B(n20900), .Z(n21176) );
  NAND U21397 ( .A(n20910), .B(n20909), .Z(n20914) );
  NAND U21398 ( .A(n20912), .B(n20911), .Z(n20913) );
  AND U21399 ( .A(n20914), .B(n20913), .Z(n21143) );
  XOR U21400 ( .A(n21143), .B(n21142), .Z(n21140) );
  OR U21401 ( .A(n20920), .B(n20919), .Z(n20924) );
  NAND U21402 ( .A(n20922), .B(n20921), .Z(n20923) );
  NAND U21403 ( .A(n20924), .B(n20923), .Z(n21139) );
  XOR U21404 ( .A(n21140), .B(n21139), .Z(n21155) );
  AND U21405 ( .A(y[2002]), .B(x[236]), .Z(n20931) );
  XOR U21406 ( .A(n20932), .B(n20931), .Z(n20984) );
  XOR U21407 ( .A(n20985), .B(n20984), .Z(n20995) );
  AND U21408 ( .A(y[2005]), .B(x[233]), .Z(n20934) );
  XOR U21409 ( .A(n20934), .B(n20933), .Z(n20994) );
  XOR U21410 ( .A(n20995), .B(n20994), .Z(n21090) );
  AND U21411 ( .A(x[251]), .B(y[1987]), .Z(n21057) );
  AND U21412 ( .A(x[225]), .B(y[2013]), .Z(n21056) );
  XOR U21413 ( .A(n21057), .B(n21056), .Z(n21054) );
  XOR U21414 ( .A(n21055), .B(n21054), .Z(n21089) );
  XOR U21415 ( .A(n21090), .B(n21089), .Z(n21087) );
  XOR U21416 ( .A(n21086), .B(n21087), .Z(n21136) );
  XNOR U21417 ( .A(n21134), .B(n21133), .Z(n21154) );
  XOR U21418 ( .A(n21153), .B(n21152), .Z(n21174) );
  XNOR U21419 ( .A(n21175), .B(n21174), .Z(n21177) );
  XNOR U21420 ( .A(n21176), .B(n21177), .Z(n21190) );
  XOR U21421 ( .A(n20939), .B(n21190), .Z(n21187) );
  XNOR U21422 ( .A(n21188), .B(n21187), .Z(n21183) );
  XNOR U21423 ( .A(n21184), .B(n21183), .Z(N447) );
  NANDN U21424 ( .A(n20945), .B(n20944), .Z(n20949) );
  NAND U21425 ( .A(n20947), .B(n20946), .Z(n20948) );
  AND U21426 ( .A(n20949), .B(n20948), .Z(n21169) );
  NAND U21427 ( .A(n20951), .B(n20950), .Z(n20955) );
  NAND U21428 ( .A(n20953), .B(n20952), .Z(n20954) );
  AND U21429 ( .A(n20955), .B(n20954), .Z(n21151) );
  NAND U21430 ( .A(n20957), .B(n20956), .Z(n20961) );
  NANDN U21431 ( .A(n20959), .B(n20958), .Z(n20960) );
  AND U21432 ( .A(n20961), .B(n20960), .Z(n21132) );
  NAND U21433 ( .A(n20963), .B(n20962), .Z(n20967) );
  NANDN U21434 ( .A(n20965), .B(n20964), .Z(n20966) );
  AND U21435 ( .A(n20967), .B(n20966), .Z(n20975) );
  NANDN U21436 ( .A(n20969), .B(n20968), .Z(n20973) );
  NANDN U21437 ( .A(n20971), .B(n20970), .Z(n20972) );
  NAND U21438 ( .A(n20973), .B(n20972), .Z(n20974) );
  XNOR U21439 ( .A(n20975), .B(n20974), .Z(n21130) );
  NAND U21440 ( .A(n20988), .B(n20987), .Z(n20991) );
  AND U21441 ( .A(x[246]), .B(y[1993]), .Z(n20998) );
  NANDN U21442 ( .A(n20989), .B(n20998), .Z(n20990) );
  NAND U21443 ( .A(n20991), .B(n20990), .Z(n20992) );
  AND U21444 ( .A(x[234]), .B(y[2005]), .Z(n21016) );
  AND U21445 ( .A(y[1988]), .B(x[251]), .Z(n21005) );
  AND U21446 ( .A(n20997), .B(o[222]), .Z(n21003) );
  AND U21447 ( .A(x[249]), .B(y[1990]), .Z(n21123) );
  XOR U21448 ( .A(n21123), .B(o[223]), .Z(n21001) );
  XNOR U21449 ( .A(n20999), .B(n20998), .Z(n21000) );
  XNOR U21450 ( .A(n21001), .B(n21000), .Z(n21002) );
  XNOR U21451 ( .A(n21003), .B(n21002), .Z(n21004) );
  XNOR U21452 ( .A(n21005), .B(n21004), .Z(n21045) );
  AND U21453 ( .A(y[1996]), .B(x[243]), .Z(n21007) );
  NAND U21454 ( .A(y[1994]), .B(x[245]), .Z(n21006) );
  XNOR U21455 ( .A(n21007), .B(n21006), .Z(n21015) );
  AND U21456 ( .A(y[1995]), .B(x[244]), .Z(n21013) );
  AND U21457 ( .A(y[1992]), .B(x[247]), .Z(n21009) );
  NAND U21458 ( .A(y[2007]), .B(x[232]), .Z(n21008) );
  XNOR U21459 ( .A(n21009), .B(n21008), .Z(n21010) );
  XNOR U21460 ( .A(n21011), .B(n21010), .Z(n21012) );
  XNOR U21461 ( .A(n21013), .B(n21012), .Z(n21014) );
  XOR U21462 ( .A(n21015), .B(n21014), .Z(n21019) );
  XNOR U21463 ( .A(n21017), .B(n21016), .Z(n21018) );
  XNOR U21464 ( .A(n21019), .B(n21018), .Z(n21035) );
  AND U21465 ( .A(y[2010]), .B(x[229]), .Z(n21021) );
  NAND U21466 ( .A(y[2009]), .B(x[230]), .Z(n21020) );
  XNOR U21467 ( .A(n21021), .B(n21020), .Z(n21025) );
  AND U21468 ( .A(y[2004]), .B(x[235]), .Z(n21023) );
  NAND U21469 ( .A(y[1989]), .B(x[250]), .Z(n21022) );
  XNOR U21470 ( .A(n21023), .B(n21022), .Z(n21024) );
  XOR U21471 ( .A(n21025), .B(n21024), .Z(n21033) );
  AND U21472 ( .A(y[1987]), .B(x[252]), .Z(n21027) );
  NAND U21473 ( .A(y[2015]), .B(x[224]), .Z(n21026) );
  XNOR U21474 ( .A(n21027), .B(n21026), .Z(n21031) );
  AND U21475 ( .A(y[2008]), .B(x[231]), .Z(n21029) );
  NAND U21476 ( .A(y[2014]), .B(x[225]), .Z(n21028) );
  XNOR U21477 ( .A(n21029), .B(n21028), .Z(n21030) );
  XNOR U21478 ( .A(n21031), .B(n21030), .Z(n21032) );
  XNOR U21479 ( .A(n21033), .B(n21032), .Z(n21034) );
  XOR U21480 ( .A(n21035), .B(n21034), .Z(n21043) );
  AND U21481 ( .A(y[2012]), .B(x[227]), .Z(n21037) );
  NAND U21482 ( .A(y[2013]), .B(x[226]), .Z(n21036) );
  XNOR U21483 ( .A(n21037), .B(n21036), .Z(n21041) );
  AND U21484 ( .A(y[1997]), .B(x[242]), .Z(n21039) );
  NAND U21485 ( .A(y[1998]), .B(x[241]), .Z(n21038) );
  XNOR U21486 ( .A(n21039), .B(n21038), .Z(n21040) );
  XNOR U21487 ( .A(n21041), .B(n21040), .Z(n21042) );
  XNOR U21488 ( .A(n21043), .B(n21042), .Z(n21044) );
  XNOR U21489 ( .A(n21045), .B(n21044), .Z(n21046) );
  NAND U21490 ( .A(n21049), .B(n21048), .Z(n21053) );
  NAND U21491 ( .A(n21051), .B(n21050), .Z(n21052) );
  AND U21492 ( .A(n21053), .B(n21052), .Z(n21085) );
  NAND U21493 ( .A(n21055), .B(n21054), .Z(n21059) );
  NAND U21494 ( .A(n21057), .B(n21056), .Z(n21058) );
  AND U21495 ( .A(n21059), .B(n21058), .Z(n21067) );
  NAND U21496 ( .A(n21061), .B(n21060), .Z(n21065) );
  NAND U21497 ( .A(n21063), .B(n21062), .Z(n21064) );
  NAND U21498 ( .A(n21065), .B(n21064), .Z(n21066) );
  XNOR U21499 ( .A(n21067), .B(n21066), .Z(n21083) );
  AND U21500 ( .A(y[1985]), .B(x[254]), .Z(n21069) );
  NAND U21501 ( .A(y[2006]), .B(x[233]), .Z(n21068) );
  XNOR U21502 ( .A(n21069), .B(n21068), .Z(n21073) );
  AND U21503 ( .A(y[2001]), .B(x[238]), .Z(n21071) );
  NAND U21504 ( .A(y[2003]), .B(x[236]), .Z(n21070) );
  XNOR U21505 ( .A(n21071), .B(n21070), .Z(n21072) );
  XOR U21506 ( .A(n21073), .B(n21072), .Z(n21081) );
  AND U21507 ( .A(y[1986]), .B(x[253]), .Z(n21075) );
  NAND U21508 ( .A(y[1999]), .B(x[240]), .Z(n21074) );
  XNOR U21509 ( .A(n21075), .B(n21074), .Z(n21079) );
  AND U21510 ( .A(y[1984]), .B(x[255]), .Z(n21077) );
  NAND U21511 ( .A(y[2011]), .B(x[228]), .Z(n21076) );
  XNOR U21512 ( .A(n21077), .B(n21076), .Z(n21078) );
  XNOR U21513 ( .A(n21079), .B(n21078), .Z(n21080) );
  XNOR U21514 ( .A(n21081), .B(n21080), .Z(n21082) );
  XNOR U21515 ( .A(n21083), .B(n21082), .Z(n21084) );
  IV U21516 ( .A(n21086), .Z(n21088) );
  NANDN U21517 ( .A(n21088), .B(n21087), .Z(n21092) );
  AND U21518 ( .A(n21090), .B(n21089), .Z(n21091) );
  ANDN U21519 ( .B(n21092), .A(n21091), .Z(n21100) );
  ANDN U21520 ( .B(n21094), .A(n21093), .Z(n21098) );
  ANDN U21521 ( .B(n21096), .A(n21095), .Z(n21097) );
  OR U21522 ( .A(n21098), .B(n21097), .Z(n21099) );
  NAND U21523 ( .A(n21102), .B(n21101), .Z(n21106) );
  NAND U21524 ( .A(n21104), .B(n21103), .Z(n21105) );
  AND U21525 ( .A(n21106), .B(n21105), .Z(n21114) );
  NAND U21526 ( .A(n21108), .B(n21107), .Z(n21112) );
  NAND U21527 ( .A(n21110), .B(n21109), .Z(n21111) );
  NAND U21528 ( .A(n21112), .B(n21111), .Z(n21113) );
  NAND U21529 ( .A(n21116), .B(n21115), .Z(n21120) );
  NAND U21530 ( .A(n21118), .B(n21117), .Z(n21119) );
  AND U21531 ( .A(n21120), .B(n21119), .Z(n21128) );
  NAND U21532 ( .A(n21122), .B(n21121), .Z(n21126) );
  NAND U21533 ( .A(n21124), .B(n21123), .Z(n21125) );
  NAND U21534 ( .A(n21126), .B(n21125), .Z(n21127) );
  XNOR U21535 ( .A(n21130), .B(n21129), .Z(n21131) );
  XNOR U21536 ( .A(n21132), .B(n21131), .Z(n21149) );
  NAND U21537 ( .A(n21134), .B(n21133), .Z(n21138) );
  NANDN U21538 ( .A(n21136), .B(n21135), .Z(n21137) );
  AND U21539 ( .A(n21138), .B(n21137), .Z(n21147) );
  IV U21540 ( .A(n21139), .Z(n21141) );
  NANDN U21541 ( .A(n21141), .B(n21140), .Z(n21145) );
  NAND U21542 ( .A(n21143), .B(n21142), .Z(n21144) );
  NAND U21543 ( .A(n21145), .B(n21144), .Z(n21146) );
  XNOR U21544 ( .A(n21147), .B(n21146), .Z(n21148) );
  XNOR U21545 ( .A(n21149), .B(n21148), .Z(n21150) );
  XNOR U21546 ( .A(n21151), .B(n21150), .Z(n21167) );
  NAND U21547 ( .A(n21153), .B(n21152), .Z(n21157) );
  NANDN U21548 ( .A(n21155), .B(n21154), .Z(n21156) );
  AND U21549 ( .A(n21157), .B(n21156), .Z(n21165) );
  NAND U21550 ( .A(n21159), .B(n21158), .Z(n21163) );
  NAND U21551 ( .A(n21161), .B(n21160), .Z(n21162) );
  NAND U21552 ( .A(n21163), .B(n21162), .Z(n21164) );
  XNOR U21553 ( .A(n21165), .B(n21164), .Z(n21166) );
  XNOR U21554 ( .A(n21167), .B(n21166), .Z(n21168) );
  AND U21555 ( .A(x[224]), .B(y[2016]), .Z(n21844) );
  XOR U21556 ( .A(n21844), .B(o[224]), .Z(N481) );
  AND U21557 ( .A(x[225]), .B(y[2016]), .Z(n21203) );
  AND U21558 ( .A(x[224]), .B(y[2017]), .Z(n21202) );
  XNOR U21559 ( .A(n21202), .B(o[225]), .Z(n21195) );
  XNOR U21560 ( .A(n21203), .B(n21195), .Z(n21197) );
  NAND U21561 ( .A(n21844), .B(o[224]), .Z(n21196) );
  XNOR U21562 ( .A(n21197), .B(n21196), .Z(N482) );
  NANDN U21563 ( .A(n21203), .B(n21195), .Z(n21199) );
  NAND U21564 ( .A(n21197), .B(n21196), .Z(n21198) );
  AND U21565 ( .A(n21199), .B(n21198), .Z(n21209) );
  AND U21566 ( .A(x[224]), .B(y[2018]), .Z(n21216) );
  XNOR U21567 ( .A(n21216), .B(o[226]), .Z(n21208) );
  XNOR U21568 ( .A(n21209), .B(n21208), .Z(n21211) );
  AND U21569 ( .A(y[2016]), .B(x[226]), .Z(n21201) );
  NAND U21570 ( .A(y[2017]), .B(x[225]), .Z(n21200) );
  XNOR U21571 ( .A(n21201), .B(n21200), .Z(n21205) );
  AND U21572 ( .A(n21202), .B(o[225]), .Z(n21204) );
  XNOR U21573 ( .A(n21205), .B(n21204), .Z(n21210) );
  XNOR U21574 ( .A(n21211), .B(n21210), .Z(N483) );
  AND U21575 ( .A(x[226]), .B(y[2017]), .Z(n21223) );
  NAND U21576 ( .A(n21223), .B(n21203), .Z(n21207) );
  NAND U21577 ( .A(n21205), .B(n21204), .Z(n21206) );
  AND U21578 ( .A(n21207), .B(n21206), .Z(n21226) );
  NANDN U21579 ( .A(n21209), .B(n21208), .Z(n21213) );
  NAND U21580 ( .A(n21211), .B(n21210), .Z(n21212) );
  AND U21581 ( .A(n21213), .B(n21212), .Z(n21225) );
  XNOR U21582 ( .A(n21226), .B(n21225), .Z(n21228) );
  AND U21583 ( .A(x[225]), .B(y[2018]), .Z(n21331) );
  XOR U21584 ( .A(n21223), .B(o[227]), .Z(n21231) );
  XOR U21585 ( .A(n21331), .B(n21231), .Z(n21233) );
  AND U21586 ( .A(y[2016]), .B(x[227]), .Z(n21215) );
  NAND U21587 ( .A(y[2019]), .B(x[224]), .Z(n21214) );
  XNOR U21588 ( .A(n21215), .B(n21214), .Z(n21218) );
  AND U21589 ( .A(n21216), .B(o[226]), .Z(n21217) );
  XOR U21590 ( .A(n21218), .B(n21217), .Z(n21232) );
  XOR U21591 ( .A(n21233), .B(n21232), .Z(n21227) );
  XOR U21592 ( .A(n21228), .B(n21227), .Z(N484) );
  AND U21593 ( .A(x[227]), .B(y[2019]), .Z(n21275) );
  NAND U21594 ( .A(n21844), .B(n21275), .Z(n21220) );
  NAND U21595 ( .A(n21218), .B(n21217), .Z(n21219) );
  AND U21596 ( .A(n21220), .B(n21219), .Z(n21254) );
  AND U21597 ( .A(y[2020]), .B(x[224]), .Z(n21222) );
  NAND U21598 ( .A(y[2016]), .B(x[228]), .Z(n21221) );
  XNOR U21599 ( .A(n21222), .B(n21221), .Z(n21247) );
  NAND U21600 ( .A(n21223), .B(o[227]), .Z(n21248) );
  AND U21601 ( .A(y[2018]), .B(x[226]), .Z(n21391) );
  NAND U21602 ( .A(y[2019]), .B(x[225]), .Z(n21224) );
  XNOR U21603 ( .A(n21391), .B(n21224), .Z(n21244) );
  AND U21604 ( .A(x[227]), .B(y[2017]), .Z(n21241) );
  XOR U21605 ( .A(o[228]), .B(n21241), .Z(n21243) );
  XOR U21606 ( .A(n21244), .B(n21243), .Z(n21251) );
  XOR U21607 ( .A(n21252), .B(n21251), .Z(n21253) );
  XOR U21608 ( .A(n21254), .B(n21253), .Z(n21259) );
  NANDN U21609 ( .A(n21226), .B(n21225), .Z(n21230) );
  NAND U21610 ( .A(n21228), .B(n21227), .Z(n21229) );
  NAND U21611 ( .A(n21230), .B(n21229), .Z(n21257) );
  NAND U21612 ( .A(n21331), .B(n21231), .Z(n21235) );
  NAND U21613 ( .A(n21233), .B(n21232), .Z(n21234) );
  NAND U21614 ( .A(n21235), .B(n21234), .Z(n21258) );
  XOR U21615 ( .A(n21257), .B(n21258), .Z(n21236) );
  XNOR U21616 ( .A(n21259), .B(n21236), .Z(N485) );
  AND U21617 ( .A(y[2018]), .B(x[227]), .Z(n21238) );
  NAND U21618 ( .A(y[2020]), .B(x[225]), .Z(n21237) );
  XNOR U21619 ( .A(n21238), .B(n21237), .Z(n21262) );
  AND U21620 ( .A(x[228]), .B(y[2017]), .Z(n21273) );
  XOR U21621 ( .A(n21273), .B(o[229]), .Z(n21261) );
  XNOR U21622 ( .A(n21262), .B(n21261), .Z(n21265) );
  NAND U21623 ( .A(x[226]), .B(y[2019]), .Z(n21340) );
  AND U21624 ( .A(y[2016]), .B(x[229]), .Z(n21240) );
  NAND U21625 ( .A(y[2021]), .B(x[224]), .Z(n21239) );
  XNOR U21626 ( .A(n21240), .B(n21239), .Z(n21268) );
  AND U21627 ( .A(o[228]), .B(n21241), .Z(n21267) );
  XOR U21628 ( .A(n21268), .B(n21267), .Z(n21266) );
  XOR U21629 ( .A(n21340), .B(n21266), .Z(n21242) );
  XOR U21630 ( .A(n21265), .B(n21242), .Z(n21283) );
  NANDN U21631 ( .A(n21340), .B(n21331), .Z(n21246) );
  NAND U21632 ( .A(n21244), .B(n21243), .Z(n21245) );
  AND U21633 ( .A(n21246), .B(n21245), .Z(n21281) );
  AND U21634 ( .A(x[228]), .B(y[2020]), .Z(n22051) );
  NAND U21635 ( .A(n22051), .B(n21844), .Z(n21250) );
  NANDN U21636 ( .A(n21248), .B(n21247), .Z(n21249) );
  NAND U21637 ( .A(n21250), .B(n21249), .Z(n21280) );
  XNOR U21638 ( .A(n21283), .B(n21282), .Z(n21279) );
  NAND U21639 ( .A(n21252), .B(n21251), .Z(n21256) );
  NANDN U21640 ( .A(n21254), .B(n21253), .Z(n21255) );
  NAND U21641 ( .A(n21256), .B(n21255), .Z(n21277) );
  XOR U21642 ( .A(n21277), .B(n21278), .Z(n21260) );
  XNOR U21643 ( .A(n21279), .B(n21260), .Z(N486) );
  AND U21644 ( .A(x[227]), .B(y[2020]), .Z(n21342) );
  NAND U21645 ( .A(n21331), .B(n21342), .Z(n21264) );
  NAND U21646 ( .A(n21262), .B(n21261), .Z(n21263) );
  NAND U21647 ( .A(n21264), .B(n21263), .Z(n21319) );
  XOR U21648 ( .A(n21319), .B(n21318), .Z(n21321) );
  AND U21649 ( .A(x[229]), .B(y[2021]), .Z(n21511) );
  NAND U21650 ( .A(n21844), .B(n21511), .Z(n21270) );
  NAND U21651 ( .A(n21268), .B(n21267), .Z(n21269) );
  AND U21652 ( .A(n21270), .B(n21269), .Z(n21288) );
  AND U21653 ( .A(y[2016]), .B(x[230]), .Z(n21272) );
  NAND U21654 ( .A(y[2022]), .B(x[224]), .Z(n21271) );
  XNOR U21655 ( .A(n21272), .B(n21271), .Z(n21294) );
  AND U21656 ( .A(n21273), .B(o[229]), .Z(n21295) );
  XOR U21657 ( .A(n21294), .B(n21295), .Z(n21287) );
  NAND U21658 ( .A(y[2020]), .B(x[226]), .Z(n21274) );
  XNOR U21659 ( .A(n21275), .B(n21274), .Z(n21299) );
  AND U21660 ( .A(y[2021]), .B(x[225]), .Z(n21562) );
  NAND U21661 ( .A(y[2018]), .B(x[228]), .Z(n21276) );
  XNOR U21662 ( .A(n21562), .B(n21276), .Z(n21303) );
  AND U21663 ( .A(x[229]), .B(y[2017]), .Z(n21308) );
  XOR U21664 ( .A(o[230]), .B(n21308), .Z(n21302) );
  XOR U21665 ( .A(n21303), .B(n21302), .Z(n21298) );
  XOR U21666 ( .A(n21299), .B(n21298), .Z(n21289) );
  XOR U21667 ( .A(n21290), .B(n21289), .Z(n21320) );
  XNOR U21668 ( .A(n21321), .B(n21320), .Z(n21314) );
  NANDN U21669 ( .A(n21281), .B(n21280), .Z(n21285) );
  NAND U21670 ( .A(n21283), .B(n21282), .Z(n21284) );
  NAND U21671 ( .A(n21285), .B(n21284), .Z(n21312) );
  IV U21672 ( .A(n21312), .Z(n21311) );
  XOR U21673 ( .A(n21313), .B(n21311), .Z(n21286) );
  XNOR U21674 ( .A(n21314), .B(n21286), .Z(N487) );
  NANDN U21675 ( .A(n21288), .B(n21287), .Z(n21292) );
  NAND U21676 ( .A(n21290), .B(n21289), .Z(n21291) );
  AND U21677 ( .A(n21292), .B(n21291), .Z(n21360) );
  AND U21678 ( .A(y[2018]), .B(x[229]), .Z(n21423) );
  NAND U21679 ( .A(y[2022]), .B(x[225]), .Z(n21293) );
  XNOR U21680 ( .A(n21423), .B(n21293), .Z(n21333) );
  NAND U21681 ( .A(x[230]), .B(y[2017]), .Z(n21337) );
  XNOR U21682 ( .A(n21333), .B(n21332), .Z(n21352) );
  AND U21683 ( .A(x[230]), .B(y[2022]), .Z(n21582) );
  NAND U21684 ( .A(n21844), .B(n21582), .Z(n21297) );
  NAND U21685 ( .A(n21295), .B(n21294), .Z(n21296) );
  AND U21686 ( .A(n21297), .B(n21296), .Z(n21351) );
  XOR U21687 ( .A(n21352), .B(n21351), .Z(n21353) );
  NANDN U21688 ( .A(n21340), .B(n21342), .Z(n21301) );
  NAND U21689 ( .A(n21299), .B(n21298), .Z(n21300) );
  AND U21690 ( .A(n21301), .B(n21300), .Z(n21354) );
  XOR U21691 ( .A(n21353), .B(n21354), .Z(n21358) );
  AND U21692 ( .A(x[228]), .B(y[2021]), .Z(n21849) );
  NAND U21693 ( .A(n21849), .B(n21331), .Z(n21305) );
  NAND U21694 ( .A(n21303), .B(n21302), .Z(n21304) );
  AND U21695 ( .A(n21305), .B(n21304), .Z(n21328) );
  AND U21696 ( .A(y[2021]), .B(x[226]), .Z(n21307) );
  NAND U21697 ( .A(y[2019]), .B(x[228]), .Z(n21306) );
  XNOR U21698 ( .A(n21307), .B(n21306), .Z(n21341) );
  XNOR U21699 ( .A(n21342), .B(n21341), .Z(n21326) );
  AND U21700 ( .A(o[230]), .B(n21308), .Z(n21346) );
  AND U21701 ( .A(y[2016]), .B(x[231]), .Z(n21310) );
  NAND U21702 ( .A(y[2023]), .B(x[224]), .Z(n21309) );
  XNOR U21703 ( .A(n21310), .B(n21309), .Z(n21345) );
  XNOR U21704 ( .A(n21346), .B(n21345), .Z(n21325) );
  XOR U21705 ( .A(n21326), .B(n21325), .Z(n21327) );
  XOR U21706 ( .A(n21328), .B(n21327), .Z(n21357) );
  XOR U21707 ( .A(n21358), .B(n21357), .Z(n21359) );
  XNOR U21708 ( .A(n21360), .B(n21359), .Z(n21366) );
  OR U21709 ( .A(n21313), .B(n21311), .Z(n21317) );
  ANDN U21710 ( .B(n21313), .A(n21312), .Z(n21315) );
  OR U21711 ( .A(n21315), .B(n21314), .Z(n21316) );
  AND U21712 ( .A(n21317), .B(n21316), .Z(n21364) );
  NAND U21713 ( .A(n21319), .B(n21318), .Z(n21323) );
  NAND U21714 ( .A(n21321), .B(n21320), .Z(n21322) );
  AND U21715 ( .A(n21323), .B(n21322), .Z(n21365) );
  IV U21716 ( .A(n21365), .Z(n21363) );
  XOR U21717 ( .A(n21364), .B(n21363), .Z(n21324) );
  XNOR U21718 ( .A(n21366), .B(n21324), .Z(N488) );
  NAND U21719 ( .A(n21326), .B(n21325), .Z(n21330) );
  NAND U21720 ( .A(n21328), .B(n21327), .Z(n21329) );
  AND U21721 ( .A(n21330), .B(n21329), .Z(n21404) );
  AND U21722 ( .A(x[229]), .B(y[2022]), .Z(n21503) );
  NAND U21723 ( .A(n21503), .B(n21331), .Z(n21335) );
  NAND U21724 ( .A(n21333), .B(n21332), .Z(n21334) );
  NAND U21725 ( .A(n21335), .B(n21334), .Z(n21402) );
  AND U21726 ( .A(y[2019]), .B(x[229]), .Z(n21953) );
  NAND U21727 ( .A(y[2023]), .B(x[225]), .Z(n21336) );
  XNOR U21728 ( .A(n21953), .B(n21336), .Z(n21383) );
  ANDN U21729 ( .B(o[231]), .A(n21337), .Z(n21382) );
  XOR U21730 ( .A(n21383), .B(n21382), .Z(n21388) );
  AND U21731 ( .A(x[227]), .B(y[2021]), .Z(n22191) );
  AND U21732 ( .A(y[2018]), .B(x[230]), .Z(n21339) );
  NAND U21733 ( .A(y[2022]), .B(x[226]), .Z(n21338) );
  XNOR U21734 ( .A(n21339), .B(n21338), .Z(n21392) );
  XNOR U21735 ( .A(n22051), .B(n21392), .Z(n21386) );
  XNOR U21736 ( .A(n22191), .B(n21386), .Z(n21387) );
  XOR U21737 ( .A(n21388), .B(n21387), .Z(n21401) );
  XOR U21738 ( .A(n21402), .B(n21401), .Z(n21403) );
  XOR U21739 ( .A(n21404), .B(n21403), .Z(n21413) );
  NANDN U21740 ( .A(n21340), .B(n21849), .Z(n21344) );
  NAND U21741 ( .A(n21342), .B(n21341), .Z(n21343) );
  NAND U21742 ( .A(n21344), .B(n21343), .Z(n21398) );
  AND U21743 ( .A(x[231]), .B(y[2023]), .Z(n21723) );
  NAND U21744 ( .A(n21844), .B(n21723), .Z(n21348) );
  NAND U21745 ( .A(n21346), .B(n21345), .Z(n21347) );
  NAND U21746 ( .A(n21348), .B(n21347), .Z(n21396) );
  AND U21747 ( .A(y[2016]), .B(x[232]), .Z(n21350) );
  NAND U21748 ( .A(y[2024]), .B(x[224]), .Z(n21349) );
  XNOR U21749 ( .A(n21350), .B(n21349), .Z(n21373) );
  AND U21750 ( .A(x[231]), .B(y[2017]), .Z(n21378) );
  XOR U21751 ( .A(o[232]), .B(n21378), .Z(n21372) );
  XOR U21752 ( .A(n21373), .B(n21372), .Z(n21395) );
  XOR U21753 ( .A(n21396), .B(n21395), .Z(n21397) );
  XNOR U21754 ( .A(n21398), .B(n21397), .Z(n21411) );
  NAND U21755 ( .A(n21352), .B(n21351), .Z(n21356) );
  NAND U21756 ( .A(n21354), .B(n21353), .Z(n21355) );
  NAND U21757 ( .A(n21356), .B(n21355), .Z(n21410) );
  XOR U21758 ( .A(n21411), .B(n21410), .Z(n21412) );
  XOR U21759 ( .A(n21413), .B(n21412), .Z(n21409) );
  NAND U21760 ( .A(n21358), .B(n21357), .Z(n21362) );
  NAND U21761 ( .A(n21360), .B(n21359), .Z(n21361) );
  NAND U21762 ( .A(n21362), .B(n21361), .Z(n21407) );
  NANDN U21763 ( .A(n21363), .B(n21364), .Z(n21369) );
  NOR U21764 ( .A(n21365), .B(n21364), .Z(n21367) );
  OR U21765 ( .A(n21367), .B(n21366), .Z(n21368) );
  AND U21766 ( .A(n21369), .B(n21368), .Z(n21408) );
  XOR U21767 ( .A(n21407), .B(n21408), .Z(n21370) );
  XNOR U21768 ( .A(n21409), .B(n21370), .Z(N489) );
  AND U21769 ( .A(x[232]), .B(y[2024]), .Z(n21371) );
  NAND U21770 ( .A(n21371), .B(n21844), .Z(n21375) );
  NAND U21771 ( .A(n21373), .B(n21372), .Z(n21374) );
  AND U21772 ( .A(n21375), .B(n21374), .Z(n21452) );
  AND U21773 ( .A(y[2020]), .B(x[229]), .Z(n21377) );
  NAND U21774 ( .A(y[2018]), .B(x[231]), .Z(n21376) );
  XNOR U21775 ( .A(n21377), .B(n21376), .Z(n21425) );
  AND U21776 ( .A(o[232]), .B(n21378), .Z(n21424) );
  XOR U21777 ( .A(n21425), .B(n21424), .Z(n21450) );
  AND U21778 ( .A(y[2016]), .B(x[233]), .Z(n21380) );
  NAND U21779 ( .A(y[2025]), .B(x[224]), .Z(n21379) );
  XNOR U21780 ( .A(n21380), .B(n21379), .Z(n21432) );
  AND U21781 ( .A(x[232]), .B(y[2017]), .Z(n21439) );
  XOR U21782 ( .A(o[233]), .B(n21439), .Z(n21431) );
  XNOR U21783 ( .A(n21432), .B(n21431), .Z(n21449) );
  XOR U21784 ( .A(n21452), .B(n21451), .Z(n21446) );
  AND U21785 ( .A(y[2019]), .B(x[230]), .Z(n21788) );
  NAND U21786 ( .A(y[2024]), .B(x[225]), .Z(n21381) );
  XNOR U21787 ( .A(n21788), .B(n21381), .Z(n21436) );
  XNOR U21788 ( .A(n21849), .B(n21436), .Z(n21455) );
  NAND U21789 ( .A(x[226]), .B(y[2023]), .Z(n22098) );
  AND U21790 ( .A(x[227]), .B(y[2022]), .Z(n21798) );
  XOR U21791 ( .A(n22098), .B(n21798), .Z(n21456) );
  XOR U21792 ( .A(n21455), .B(n21456), .Z(n21444) );
  NAND U21793 ( .A(x[229]), .B(y[2023]), .Z(n21637) );
  AND U21794 ( .A(x[225]), .B(y[2019]), .Z(n21435) );
  NANDN U21795 ( .A(n21637), .B(n21435), .Z(n21385) );
  NAND U21796 ( .A(n21383), .B(n21382), .Z(n21384) );
  NAND U21797 ( .A(n21385), .B(n21384), .Z(n21443) );
  XOR U21798 ( .A(n21444), .B(n21443), .Z(n21445) );
  NANDN U21799 ( .A(n22191), .B(n21386), .Z(n21390) );
  NANDN U21800 ( .A(n21388), .B(n21387), .Z(n21389) );
  AND U21801 ( .A(n21390), .B(n21389), .Z(n21418) );
  NAND U21802 ( .A(n21582), .B(n21391), .Z(n21394) );
  NAND U21803 ( .A(n22051), .B(n21392), .Z(n21393) );
  AND U21804 ( .A(n21394), .B(n21393), .Z(n21417) );
  XNOR U21805 ( .A(n21419), .B(n21420), .Z(n21464) );
  NAND U21806 ( .A(n21396), .B(n21395), .Z(n21400) );
  NAND U21807 ( .A(n21398), .B(n21397), .Z(n21399) );
  NAND U21808 ( .A(n21400), .B(n21399), .Z(n21463) );
  NAND U21809 ( .A(n21402), .B(n21401), .Z(n21406) );
  NAND U21810 ( .A(n21404), .B(n21403), .Z(n21405) );
  NAND U21811 ( .A(n21406), .B(n21405), .Z(n21462) );
  XOR U21812 ( .A(n21463), .B(n21462), .Z(n21465) );
  XNOR U21813 ( .A(n21464), .B(n21465), .Z(n21461) );
  NAND U21814 ( .A(n21411), .B(n21410), .Z(n21415) );
  NANDN U21815 ( .A(n21413), .B(n21412), .Z(n21414) );
  AND U21816 ( .A(n21415), .B(n21414), .Z(n21460) );
  XOR U21817 ( .A(n21459), .B(n21460), .Z(n21416) );
  XNOR U21818 ( .A(n21461), .B(n21416), .Z(N490) );
  NANDN U21819 ( .A(n21418), .B(n21417), .Z(n21422) );
  NAND U21820 ( .A(n21420), .B(n21419), .Z(n21421) );
  AND U21821 ( .A(n21422), .B(n21421), .Z(n21524) );
  AND U21822 ( .A(x[231]), .B(y[2020]), .Z(n21505) );
  NAND U21823 ( .A(n21505), .B(n21423), .Z(n21427) );
  NAND U21824 ( .A(n21425), .B(n21424), .Z(n21426) );
  AND U21825 ( .A(n21427), .B(n21426), .Z(n21518) );
  AND U21826 ( .A(y[2019]), .B(x[231]), .Z(n21429) );
  NAND U21827 ( .A(y[2022]), .B(x[228]), .Z(n21428) );
  XNOR U21828 ( .A(n21429), .B(n21428), .Z(n21489) );
  AND U21829 ( .A(x[230]), .B(y[2020]), .Z(n21488) );
  XNOR U21830 ( .A(n21489), .B(n21488), .Z(n21516) );
  AND U21831 ( .A(x[232]), .B(y[2018]), .Z(n21697) );
  NAND U21832 ( .A(x[233]), .B(y[2017]), .Z(n21499) );
  XOR U21833 ( .A(n21697), .B(n21510), .Z(n21512) );
  XNOR U21834 ( .A(n21512), .B(n21511), .Z(n21515) );
  XOR U21835 ( .A(n21516), .B(n21515), .Z(n21517) );
  XNOR U21836 ( .A(n21518), .B(n21517), .Z(n21477) );
  AND U21837 ( .A(x[233]), .B(y[2025]), .Z(n21430) );
  NAND U21838 ( .A(n21430), .B(n21844), .Z(n21434) );
  NAND U21839 ( .A(n21432), .B(n21431), .Z(n21433) );
  NAND U21840 ( .A(n21434), .B(n21433), .Z(n21475) );
  AND U21841 ( .A(x[230]), .B(y[2024]), .Z(n21733) );
  NAND U21842 ( .A(n21733), .B(n21435), .Z(n21438) );
  NAND U21843 ( .A(n21436), .B(n21849), .Z(n21437) );
  NAND U21844 ( .A(n21438), .B(n21437), .Z(n21484) );
  AND U21845 ( .A(o[233]), .B(n21439), .Z(n21494) );
  AND U21846 ( .A(y[2016]), .B(x[234]), .Z(n21441) );
  AND U21847 ( .A(y[2026]), .B(x[224]), .Z(n21440) );
  XOR U21848 ( .A(n21441), .B(n21440), .Z(n21493) );
  XOR U21849 ( .A(n21494), .B(n21493), .Z(n21482) );
  AND U21850 ( .A(y[2023]), .B(x[227]), .Z(n22427) );
  NAND U21851 ( .A(y[2025]), .B(x[225]), .Z(n21442) );
  XNOR U21852 ( .A(n22427), .B(n21442), .Z(n21506) );
  AND U21853 ( .A(x[226]), .B(y[2024]), .Z(n21507) );
  XOR U21854 ( .A(n21506), .B(n21507), .Z(n21481) );
  XOR U21855 ( .A(n21482), .B(n21481), .Z(n21483) );
  XNOR U21856 ( .A(n21484), .B(n21483), .Z(n21476) );
  XOR U21857 ( .A(n21475), .B(n21476), .Z(n21478) );
  XOR U21858 ( .A(n21477), .B(n21478), .Z(n21522) );
  NAND U21859 ( .A(n21444), .B(n21443), .Z(n21448) );
  NANDN U21860 ( .A(n21446), .B(n21445), .Z(n21447) );
  NAND U21861 ( .A(n21448), .B(n21447), .Z(n21471) );
  NANDN U21862 ( .A(n21450), .B(n21449), .Z(n21454) );
  NAND U21863 ( .A(n21452), .B(n21451), .Z(n21453) );
  AND U21864 ( .A(n21454), .B(n21453), .Z(n21470) );
  NANDN U21865 ( .A(n21456), .B(n21455), .Z(n21458) );
  ANDN U21866 ( .B(n22098), .A(n21798), .Z(n21457) );
  ANDN U21867 ( .B(n21458), .A(n21457), .Z(n21469) );
  XOR U21868 ( .A(n21470), .B(n21469), .Z(n21472) );
  XNOR U21869 ( .A(n21471), .B(n21472), .Z(n21521) );
  XOR U21870 ( .A(n21522), .B(n21521), .Z(n21523) );
  XOR U21871 ( .A(n21524), .B(n21523), .Z(n21530) );
  NAND U21872 ( .A(n21463), .B(n21462), .Z(n21467) );
  NAND U21873 ( .A(n21465), .B(n21464), .Z(n21466) );
  AND U21874 ( .A(n21467), .B(n21466), .Z(n21529) );
  IV U21875 ( .A(n21529), .Z(n21527) );
  XOR U21876 ( .A(n21528), .B(n21527), .Z(n21468) );
  XNOR U21877 ( .A(n21530), .B(n21468), .Z(N491) );
  NAND U21878 ( .A(n21470), .B(n21469), .Z(n21474) );
  NAND U21879 ( .A(n21472), .B(n21471), .Z(n21473) );
  NAND U21880 ( .A(n21474), .B(n21473), .Z(n21595) );
  NANDN U21881 ( .A(n21476), .B(n21475), .Z(n21480) );
  NANDN U21882 ( .A(n21478), .B(n21477), .Z(n21479) );
  NAND U21883 ( .A(n21480), .B(n21479), .Z(n21594) );
  NAND U21884 ( .A(n21482), .B(n21481), .Z(n21486) );
  NAND U21885 ( .A(n21484), .B(n21483), .Z(n21485) );
  NAND U21886 ( .A(n21486), .B(n21485), .Z(n21548) );
  AND U21887 ( .A(x[231]), .B(y[2022]), .Z(n21632) );
  AND U21888 ( .A(x[228]), .B(y[2019]), .Z(n21487) );
  NAND U21889 ( .A(n21632), .B(n21487), .Z(n21491) );
  NAND U21890 ( .A(n21489), .B(n21488), .Z(n21490) );
  NAND U21891 ( .A(n21491), .B(n21490), .Z(n21546) );
  AND U21892 ( .A(x[234]), .B(y[2026]), .Z(n21492) );
  NAND U21893 ( .A(n21492), .B(n21844), .Z(n21496) );
  NAND U21894 ( .A(n21494), .B(n21493), .Z(n21495) );
  NAND U21895 ( .A(n21496), .B(n21495), .Z(n21542) );
  AND U21896 ( .A(y[2016]), .B(x[235]), .Z(n21498) );
  NAND U21897 ( .A(y[2027]), .B(x[224]), .Z(n21497) );
  XNOR U21898 ( .A(n21498), .B(n21497), .Z(n21573) );
  ANDN U21899 ( .B(o[234]), .A(n21499), .Z(n21572) );
  XOR U21900 ( .A(n21573), .B(n21572), .Z(n21541) );
  AND U21901 ( .A(y[2021]), .B(x[230]), .Z(n21501) );
  NAND U21902 ( .A(y[2026]), .B(x[225]), .Z(n21500) );
  XNOR U21903 ( .A(n21501), .B(n21500), .Z(n21564) );
  AND U21904 ( .A(x[234]), .B(y[2017]), .Z(n21583) );
  XOR U21905 ( .A(o[235]), .B(n21583), .Z(n21563) );
  XOR U21906 ( .A(n21564), .B(n21563), .Z(n21540) );
  XOR U21907 ( .A(n21541), .B(n21540), .Z(n21543) );
  XNOR U21908 ( .A(n21542), .B(n21543), .Z(n21547) );
  XOR U21909 ( .A(n21548), .B(n21549), .Z(n21586) );
  AND U21910 ( .A(x[227]), .B(y[2024]), .Z(n22568) );
  NAND U21911 ( .A(y[2025]), .B(x[226]), .Z(n21502) );
  XNOR U21912 ( .A(n21503), .B(n21502), .Z(n21559) );
  AND U21913 ( .A(x[228]), .B(y[2023]), .Z(n21558) );
  XNOR U21914 ( .A(n21559), .B(n21558), .Z(n21535) );
  XNOR U21915 ( .A(n22568), .B(n21535), .Z(n21537) );
  NAND U21916 ( .A(y[2018]), .B(x[233]), .Z(n21504) );
  XNOR U21917 ( .A(n21505), .B(n21504), .Z(n21578) );
  AND U21918 ( .A(x[232]), .B(y[2019]), .Z(n21577) );
  XNOR U21919 ( .A(n21578), .B(n21577), .Z(n21536) );
  XNOR U21920 ( .A(n21537), .B(n21536), .Z(n21555) );
  AND U21921 ( .A(x[227]), .B(y[2025]), .Z(n21628) );
  AND U21922 ( .A(x[225]), .B(y[2023]), .Z(n21839) );
  NAND U21923 ( .A(n21628), .B(n21839), .Z(n21509) );
  NAND U21924 ( .A(n21507), .B(n21506), .Z(n21508) );
  NAND U21925 ( .A(n21509), .B(n21508), .Z(n21553) );
  NAND U21926 ( .A(n21697), .B(n21510), .Z(n21514) );
  NAND U21927 ( .A(n21512), .B(n21511), .Z(n21513) );
  NAND U21928 ( .A(n21514), .B(n21513), .Z(n21552) );
  XOR U21929 ( .A(n21553), .B(n21552), .Z(n21554) );
  XNOR U21930 ( .A(n21555), .B(n21554), .Z(n21585) );
  NAND U21931 ( .A(n21516), .B(n21515), .Z(n21520) );
  NAND U21932 ( .A(n21518), .B(n21517), .Z(n21519) );
  NAND U21933 ( .A(n21520), .B(n21519), .Z(n21584) );
  XOR U21934 ( .A(n21585), .B(n21584), .Z(n21587) );
  XNOR U21935 ( .A(n21586), .B(n21587), .Z(n21593) );
  XOR U21936 ( .A(n21594), .B(n21593), .Z(n21596) );
  XOR U21937 ( .A(n21595), .B(n21596), .Z(n21592) );
  NAND U21938 ( .A(n21522), .B(n21521), .Z(n21526) );
  NANDN U21939 ( .A(n21524), .B(n21523), .Z(n21525) );
  NAND U21940 ( .A(n21526), .B(n21525), .Z(n21590) );
  NANDN U21941 ( .A(n21527), .B(n21528), .Z(n21533) );
  NOR U21942 ( .A(n21529), .B(n21528), .Z(n21531) );
  OR U21943 ( .A(n21531), .B(n21530), .Z(n21532) );
  AND U21944 ( .A(n21533), .B(n21532), .Z(n21591) );
  XOR U21945 ( .A(n21590), .B(n21591), .Z(n21534) );
  XNOR U21946 ( .A(n21592), .B(n21534), .Z(N492) );
  NANDN U21947 ( .A(n22568), .B(n21535), .Z(n21539) );
  NAND U21948 ( .A(n21537), .B(n21536), .Z(n21538) );
  NAND U21949 ( .A(n21539), .B(n21538), .Z(n21609) );
  NAND U21950 ( .A(n21541), .B(n21540), .Z(n21545) );
  NAND U21951 ( .A(n21543), .B(n21542), .Z(n21544) );
  AND U21952 ( .A(n21545), .B(n21544), .Z(n21610) );
  XOR U21953 ( .A(n21609), .B(n21610), .Z(n21612) );
  NANDN U21954 ( .A(n21547), .B(n21546), .Z(n21551) );
  NANDN U21955 ( .A(n21549), .B(n21548), .Z(n21550) );
  AND U21956 ( .A(n21551), .B(n21550), .Z(n21611) );
  XOR U21957 ( .A(n21612), .B(n21611), .Z(n21603) );
  NAND U21958 ( .A(n21553), .B(n21552), .Z(n21557) );
  NAND U21959 ( .A(n21555), .B(n21554), .Z(n21556) );
  NAND U21960 ( .A(n21557), .B(n21556), .Z(n21668) );
  AND U21961 ( .A(x[229]), .B(y[2025]), .Z(n22089) );
  AND U21962 ( .A(x[226]), .B(y[2022]), .Z(n22278) );
  NAND U21963 ( .A(n22089), .B(n22278), .Z(n21561) );
  NAND U21964 ( .A(n21559), .B(n21558), .Z(n21560) );
  AND U21965 ( .A(n21561), .B(n21560), .Z(n21616) );
  AND U21966 ( .A(x[230]), .B(y[2026]), .Z(n21856) );
  NAND U21967 ( .A(n21856), .B(n21562), .Z(n21566) );
  NAND U21968 ( .A(n21564), .B(n21563), .Z(n21565) );
  NAND U21969 ( .A(n21566), .B(n21565), .Z(n21615) );
  AND U21970 ( .A(x[233]), .B(y[2019]), .Z(n22273) );
  AND U21971 ( .A(y[2018]), .B(x[234]), .Z(n22315) );
  NAND U21972 ( .A(y[2024]), .B(x[228]), .Z(n21567) );
  XOR U21973 ( .A(n22315), .B(n21567), .Z(n21659) );
  NAND U21974 ( .A(x[231]), .B(y[2021]), .Z(n21636) );
  XOR U21975 ( .A(n21637), .B(n21636), .Z(n21639) );
  AND U21976 ( .A(y[2016]), .B(x[236]), .Z(n21569) );
  NAND U21977 ( .A(y[2028]), .B(x[224]), .Z(n21568) );
  XNOR U21978 ( .A(n21569), .B(n21568), .Z(n21653) );
  AND U21979 ( .A(x[235]), .B(y[2017]), .Z(n21633) );
  XOR U21980 ( .A(o[236]), .B(n21633), .Z(n21652) );
  XOR U21981 ( .A(n21653), .B(n21652), .Z(n21622) );
  AND U21982 ( .A(y[2026]), .B(x[226]), .Z(n21571) );
  NAND U21983 ( .A(y[2020]), .B(x[232]), .Z(n21570) );
  XNOR U21984 ( .A(n21571), .B(n21570), .Z(n21627) );
  XOR U21985 ( .A(n21627), .B(n21628), .Z(n21621) );
  XOR U21986 ( .A(n21622), .B(n21621), .Z(n21624) );
  XOR U21987 ( .A(n21623), .B(n21624), .Z(n21617) );
  XOR U21988 ( .A(n21618), .B(n21617), .Z(n21667) );
  AND U21989 ( .A(x[235]), .B(y[2027]), .Z(n22679) );
  NAND U21990 ( .A(n22679), .B(n21844), .Z(n21575) );
  NAND U21991 ( .A(n21573), .B(n21572), .Z(n21574) );
  AND U21992 ( .A(n21575), .B(n21574), .Z(n21645) );
  AND U21993 ( .A(x[231]), .B(y[2018]), .Z(n21774) );
  AND U21994 ( .A(x[233]), .B(y[2020]), .Z(n21576) );
  NAND U21995 ( .A(n21774), .B(n21576), .Z(n21580) );
  NAND U21996 ( .A(n21578), .B(n21577), .Z(n21579) );
  AND U21997 ( .A(n21580), .B(n21579), .Z(n21643) );
  NAND U21998 ( .A(y[2027]), .B(x[225]), .Z(n21581) );
  XNOR U21999 ( .A(n21582), .B(n21581), .Z(n21649) );
  AND U22000 ( .A(o[235]), .B(n21583), .Z(n21648) );
  XOR U22001 ( .A(n21649), .B(n21648), .Z(n21642) );
  XOR U22002 ( .A(n21667), .B(n21666), .Z(n21669) );
  XNOR U22003 ( .A(n21668), .B(n21669), .Z(n21601) );
  NAND U22004 ( .A(n21585), .B(n21584), .Z(n21589) );
  NAND U22005 ( .A(n21587), .B(n21586), .Z(n21588) );
  NAND U22006 ( .A(n21589), .B(n21588), .Z(n21600) );
  XOR U22007 ( .A(n21601), .B(n21600), .Z(n21602) );
  XNOR U22008 ( .A(n21603), .B(n21602), .Z(n21608) );
  NAND U22009 ( .A(n21594), .B(n21593), .Z(n21598) );
  NAND U22010 ( .A(n21596), .B(n21595), .Z(n21597) );
  AND U22011 ( .A(n21598), .B(n21597), .Z(n21606) );
  XOR U22012 ( .A(n21607), .B(n21606), .Z(n21599) );
  XNOR U22013 ( .A(n21608), .B(n21599), .Z(N493) );
  NAND U22014 ( .A(n21601), .B(n21600), .Z(n21605) );
  NAND U22015 ( .A(n21603), .B(n21602), .Z(n21604) );
  AND U22016 ( .A(n21605), .B(n21604), .Z(n21741) );
  NAND U22017 ( .A(n21610), .B(n21609), .Z(n21614) );
  NAND U22018 ( .A(n21612), .B(n21611), .Z(n21613) );
  NAND U22019 ( .A(n21614), .B(n21613), .Z(n21745) );
  NANDN U22020 ( .A(n21616), .B(n21615), .Z(n21620) );
  NAND U22021 ( .A(n21618), .B(n21617), .Z(n21619) );
  AND U22022 ( .A(n21620), .B(n21619), .Z(n21674) );
  NAND U22023 ( .A(n21622), .B(n21621), .Z(n21626) );
  NAND U22024 ( .A(n21624), .B(n21623), .Z(n21625) );
  NAND U22025 ( .A(n21626), .B(n21625), .Z(n21681) );
  AND U22026 ( .A(y[2026]), .B(x[232]), .Z(n22920) );
  AND U22027 ( .A(x[226]), .B(y[2020]), .Z(n21784) );
  NAND U22028 ( .A(n22920), .B(n21784), .Z(n21630) );
  NAND U22029 ( .A(n21628), .B(n21627), .Z(n21629) );
  NAND U22030 ( .A(n21630), .B(n21629), .Z(n21712) );
  NAND U22031 ( .A(y[2028]), .B(x[225]), .Z(n21631) );
  XNOR U22032 ( .A(n21632), .B(n21631), .Z(n21703) );
  AND U22033 ( .A(o[236]), .B(n21633), .Z(n21702) );
  XOR U22034 ( .A(n21703), .B(n21702), .Z(n21710) );
  AND U22035 ( .A(x[230]), .B(y[2023]), .Z(n22719) );
  AND U22036 ( .A(y[2027]), .B(x[226]), .Z(n21635) );
  NAND U22037 ( .A(y[2020]), .B(x[233]), .Z(n21634) );
  XNOR U22038 ( .A(n21635), .B(n21634), .Z(n21716) );
  XOR U22039 ( .A(n22719), .B(n21716), .Z(n21709) );
  XOR U22040 ( .A(n21710), .B(n21709), .Z(n21711) );
  XOR U22041 ( .A(n21712), .B(n21711), .Z(n21680) );
  NAND U22042 ( .A(n21637), .B(n21636), .Z(n21641) );
  ANDN U22043 ( .B(n21639), .A(n21638), .Z(n21640) );
  ANDN U22044 ( .B(n21641), .A(n21640), .Z(n21679) );
  XOR U22045 ( .A(n21680), .B(n21679), .Z(n21682) );
  XOR U22046 ( .A(n21681), .B(n21682), .Z(n21673) );
  NANDN U22047 ( .A(n21643), .B(n21642), .Z(n21647) );
  NANDN U22048 ( .A(n21645), .B(n21644), .Z(n21646) );
  AND U22049 ( .A(n21647), .B(n21646), .Z(n21688) );
  AND U22050 ( .A(x[230]), .B(y[2027]), .Z(n22012) );
  IV U22051 ( .A(n22012), .Z(n22091) );
  AND U22052 ( .A(x[225]), .B(y[2022]), .Z(n21701) );
  NANDN U22053 ( .A(n22091), .B(n21701), .Z(n21651) );
  NAND U22054 ( .A(n21649), .B(n21648), .Z(n21650) );
  NAND U22055 ( .A(n21651), .B(n21650), .Z(n21694) );
  AND U22056 ( .A(x[236]), .B(y[2028]), .Z(n22928) );
  NAND U22057 ( .A(n22928), .B(n21844), .Z(n21655) );
  NAND U22058 ( .A(n21653), .B(n21652), .Z(n21654) );
  NAND U22059 ( .A(n21655), .B(n21654), .Z(n21692) );
  AND U22060 ( .A(x[234]), .B(y[2019]), .Z(n22580) );
  AND U22061 ( .A(y[2018]), .B(x[235]), .Z(n22541) );
  NAND U22062 ( .A(y[2021]), .B(x[232]), .Z(n21656) );
  XNOR U22063 ( .A(n22541), .B(n21656), .Z(n21698) );
  XOR U22064 ( .A(n22580), .B(n21698), .Z(n21691) );
  XOR U22065 ( .A(n21692), .B(n21691), .Z(n21693) );
  XOR U22066 ( .A(n21694), .B(n21693), .Z(n21686) );
  AND U22067 ( .A(x[234]), .B(y[2024]), .Z(n21658) );
  AND U22068 ( .A(x[228]), .B(y[2018]), .Z(n21657) );
  NAND U22069 ( .A(n21658), .B(n21657), .Z(n21661) );
  NANDN U22070 ( .A(n21659), .B(n22273), .Z(n21660) );
  AND U22071 ( .A(n21661), .B(n21660), .Z(n21737) );
  AND U22072 ( .A(y[2016]), .B(x[237]), .Z(n21663) );
  NAND U22073 ( .A(y[2029]), .B(x[224]), .Z(n21662) );
  XNOR U22074 ( .A(n21663), .B(n21662), .Z(n21729) );
  AND U22075 ( .A(x[236]), .B(y[2017]), .Z(n21721) );
  XOR U22076 ( .A(o[237]), .B(n21721), .Z(n21728) );
  XOR U22077 ( .A(n21729), .B(n21728), .Z(n21735) );
  AND U22078 ( .A(y[2024]), .B(x[229]), .Z(n21665) );
  NAND U22079 ( .A(y[2026]), .B(x[227]), .Z(n21664) );
  XNOR U22080 ( .A(n21665), .B(n21664), .Z(n21724) );
  AND U22081 ( .A(x[228]), .B(y[2025]), .Z(n21725) );
  XOR U22082 ( .A(n21724), .B(n21725), .Z(n21734) );
  XOR U22083 ( .A(n21735), .B(n21734), .Z(n21736) );
  XOR U22084 ( .A(n21686), .B(n21685), .Z(n21687) );
  XOR U22085 ( .A(n21676), .B(n21675), .Z(n21744) );
  NAND U22086 ( .A(n21667), .B(n21666), .Z(n21671) );
  NAND U22087 ( .A(n21669), .B(n21668), .Z(n21670) );
  AND U22088 ( .A(n21671), .B(n21670), .Z(n21743) );
  XOR U22089 ( .A(n21745), .B(n21746), .Z(n21742) );
  XNOR U22090 ( .A(n21740), .B(n21742), .Z(n21672) );
  XOR U22091 ( .A(n21741), .B(n21672), .Z(N494) );
  NANDN U22092 ( .A(n21674), .B(n21673), .Z(n21678) );
  NAND U22093 ( .A(n21676), .B(n21675), .Z(n21677) );
  AND U22094 ( .A(n21678), .B(n21677), .Z(n21833) );
  NAND U22095 ( .A(n21680), .B(n21679), .Z(n21684) );
  NAND U22096 ( .A(n21682), .B(n21681), .Z(n21683) );
  NAND U22097 ( .A(n21684), .B(n21683), .Z(n21832) );
  NAND U22098 ( .A(n21686), .B(n21685), .Z(n21690) );
  NANDN U22099 ( .A(n21688), .B(n21687), .Z(n21689) );
  AND U22100 ( .A(n21690), .B(n21689), .Z(n21753) );
  NAND U22101 ( .A(n21692), .B(n21691), .Z(n21696) );
  NAND U22102 ( .A(n21694), .B(n21693), .Z(n21695) );
  AND U22103 ( .A(n21696), .B(n21695), .Z(n21759) );
  AND U22104 ( .A(x[235]), .B(y[2021]), .Z(n21870) );
  NAND U22105 ( .A(n21870), .B(n21697), .Z(n21700) );
  NAND U22106 ( .A(n21698), .B(n22580), .Z(n21699) );
  NAND U22107 ( .A(n21700), .B(n21699), .Z(n21814) );
  NAND U22108 ( .A(x[231]), .B(y[2028]), .Z(n22288) );
  NANDN U22109 ( .A(n22288), .B(n21701), .Z(n21705) );
  NAND U22110 ( .A(n21703), .B(n21702), .Z(n21704) );
  NAND U22111 ( .A(n21705), .B(n21704), .Z(n21813) );
  XOR U22112 ( .A(n21814), .B(n21813), .Z(n21816) );
  AND U22113 ( .A(x[228]), .B(y[2026]), .Z(n22200) );
  AND U22114 ( .A(y[2027]), .B(x[227]), .Z(n21707) );
  NAND U22115 ( .A(y[2022]), .B(x[232]), .Z(n21706) );
  XNOR U22116 ( .A(n21707), .B(n21706), .Z(n21799) );
  XOR U22117 ( .A(n22089), .B(n21799), .Z(n21808) );
  XOR U22118 ( .A(n22200), .B(n21808), .Z(n21810) );
  AND U22119 ( .A(x[233]), .B(y[2021]), .Z(n22398) );
  AND U22120 ( .A(y[2028]), .B(x[226]), .Z(n21708) );
  AND U22121 ( .A(y[2020]), .B(x[234]), .Z(n22422) );
  XOR U22122 ( .A(n21708), .B(n22422), .Z(n21785) );
  XOR U22123 ( .A(n22398), .B(n21785), .Z(n21809) );
  XOR U22124 ( .A(n21810), .B(n21809), .Z(n21815) );
  XNOR U22125 ( .A(n21816), .B(n21815), .Z(n21757) );
  NAND U22126 ( .A(n21710), .B(n21709), .Z(n21714) );
  NAND U22127 ( .A(n21712), .B(n21711), .Z(n21713) );
  AND U22128 ( .A(n21714), .B(n21713), .Z(n21756) );
  XOR U22129 ( .A(n21757), .B(n21756), .Z(n21758) );
  XOR U22130 ( .A(n21759), .B(n21758), .Z(n21751) );
  AND U22131 ( .A(x[233]), .B(y[2027]), .Z(n21715) );
  NAND U22132 ( .A(n21715), .B(n21784), .Z(n21718) );
  NAND U22133 ( .A(n21716), .B(n22719), .Z(n21717) );
  NAND U22134 ( .A(n21718), .B(n21717), .Z(n21771) );
  AND U22135 ( .A(y[2016]), .B(x[238]), .Z(n21720) );
  NAND U22136 ( .A(y[2030]), .B(x[224]), .Z(n21719) );
  XNOR U22137 ( .A(n21720), .B(n21719), .Z(n21794) );
  AND U22138 ( .A(o[237]), .B(n21721), .Z(n21793) );
  XOR U22139 ( .A(n21794), .B(n21793), .Z(n21769) );
  NAND U22140 ( .A(y[2018]), .B(x[236]), .Z(n21722) );
  XNOR U22141 ( .A(n21723), .B(n21722), .Z(n21776) );
  AND U22142 ( .A(x[237]), .B(y[2017]), .Z(n21783) );
  XOR U22143 ( .A(o[238]), .B(n21783), .Z(n21775) );
  XOR U22144 ( .A(n21776), .B(n21775), .Z(n21768) );
  XOR U22145 ( .A(n21769), .B(n21768), .Z(n21770) );
  XNOR U22146 ( .A(n21771), .B(n21770), .Z(n21820) );
  AND U22147 ( .A(x[229]), .B(y[2026]), .Z(n21857) );
  NAND U22148 ( .A(n22568), .B(n21857), .Z(n21727) );
  NAND U22149 ( .A(n21725), .B(n21724), .Z(n21726) );
  AND U22150 ( .A(n21727), .B(n21726), .Z(n21765) );
  AND U22151 ( .A(x[237]), .B(y[2029]), .Z(n23307) );
  NAND U22152 ( .A(n23307), .B(n21844), .Z(n21731) );
  NAND U22153 ( .A(n21729), .B(n21728), .Z(n21730) );
  NAND U22154 ( .A(n21731), .B(n21730), .Z(n21763) );
  NAND U22155 ( .A(y[2019]), .B(x[235]), .Z(n21732) );
  XNOR U22156 ( .A(n21733), .B(n21732), .Z(n21789) );
  AND U22157 ( .A(x[225]), .B(y[2029]), .Z(n21790) );
  XOR U22158 ( .A(n21789), .B(n21790), .Z(n21762) );
  XOR U22159 ( .A(n21763), .B(n21762), .Z(n21764) );
  XOR U22160 ( .A(n21765), .B(n21764), .Z(n21819) );
  XOR U22161 ( .A(n21820), .B(n21819), .Z(n21822) );
  NAND U22162 ( .A(n21735), .B(n21734), .Z(n21739) );
  NANDN U22163 ( .A(n21737), .B(n21736), .Z(n21738) );
  AND U22164 ( .A(n21739), .B(n21738), .Z(n21821) );
  XNOR U22165 ( .A(n21822), .B(n21821), .Z(n21750) );
  XNOR U22166 ( .A(n21835), .B(n21834), .Z(n21828) );
  NANDN U22167 ( .A(n21744), .B(n21743), .Z(n21748) );
  NAND U22168 ( .A(n21746), .B(n21745), .Z(n21747) );
  AND U22169 ( .A(n21748), .B(n21747), .Z(n21826) );
  IV U22170 ( .A(n21826), .Z(n21825) );
  XOR U22171 ( .A(n21827), .B(n21825), .Z(n21749) );
  XNOR U22172 ( .A(n21828), .B(n21749), .Z(N495) );
  NANDN U22173 ( .A(n21751), .B(n21750), .Z(n21755) );
  NANDN U22174 ( .A(n21753), .B(n21752), .Z(n21754) );
  AND U22175 ( .A(n21755), .B(n21754), .Z(n21931) );
  NAND U22176 ( .A(n21757), .B(n21756), .Z(n21761) );
  NAND U22177 ( .A(n21759), .B(n21758), .Z(n21760) );
  NAND U22178 ( .A(n21761), .B(n21760), .Z(n21900) );
  NAND U22179 ( .A(n21763), .B(n21762), .Z(n21767) );
  NANDN U22180 ( .A(n21765), .B(n21764), .Z(n21766) );
  NAND U22181 ( .A(n21767), .B(n21766), .Z(n21906) );
  NAND U22182 ( .A(n21769), .B(n21768), .Z(n21773) );
  NAND U22183 ( .A(n21771), .B(n21770), .Z(n21772) );
  NAND U22184 ( .A(n21773), .B(n21772), .Z(n21904) );
  AND U22185 ( .A(x[236]), .B(y[2023]), .Z(n22279) );
  NAND U22186 ( .A(n22279), .B(n21774), .Z(n21778) );
  NAND U22187 ( .A(n21776), .B(n21775), .Z(n21777) );
  AND U22188 ( .A(n21778), .B(n21777), .Z(n21880) );
  AND U22189 ( .A(y[2020]), .B(x[235]), .Z(n21780) );
  NAND U22190 ( .A(y[2018]), .B(x[237]), .Z(n21779) );
  XNOR U22191 ( .A(n21780), .B(n21779), .Z(n21884) );
  AND U22192 ( .A(x[236]), .B(y[2019]), .Z(n21883) );
  XNOR U22193 ( .A(n21884), .B(n21883), .Z(n21878) );
  AND U22194 ( .A(y[2016]), .B(x[239]), .Z(n21782) );
  NAND U22195 ( .A(y[2031]), .B(x[224]), .Z(n21781) );
  XNOR U22196 ( .A(n21782), .B(n21781), .Z(n21846) );
  AND U22197 ( .A(o[238]), .B(n21783), .Z(n21845) );
  XNOR U22198 ( .A(n21846), .B(n21845), .Z(n21877) );
  XOR U22199 ( .A(n21878), .B(n21877), .Z(n21879) );
  XNOR U22200 ( .A(n21880), .B(n21879), .Z(n21912) );
  NAND U22201 ( .A(x[234]), .B(y[2028]), .Z(n22721) );
  NANDN U22202 ( .A(n22721), .B(n21784), .Z(n21787) );
  NAND U22203 ( .A(n22398), .B(n21785), .Z(n21786) );
  NAND U22204 ( .A(n21787), .B(n21786), .Z(n21910) );
  AND U22205 ( .A(x[235]), .B(y[2024]), .Z(n22199) );
  NAND U22206 ( .A(n22199), .B(n21788), .Z(n21792) );
  NAND U22207 ( .A(n21790), .B(n21789), .Z(n21791) );
  NAND U22208 ( .A(n21792), .B(n21791), .Z(n21909) );
  XOR U22209 ( .A(n21910), .B(n21909), .Z(n21911) );
  XOR U22210 ( .A(n21912), .B(n21911), .Z(n21903) );
  XOR U22211 ( .A(n21904), .B(n21903), .Z(n21905) );
  XNOR U22212 ( .A(n21906), .B(n21905), .Z(n21897) );
  AND U22213 ( .A(x[238]), .B(y[2030]), .Z(n23573) );
  NAND U22214 ( .A(n23573), .B(n21844), .Z(n21796) );
  NAND U22215 ( .A(n21794), .B(n21793), .Z(n21795) );
  NAND U22216 ( .A(n21796), .B(n21795), .Z(n21872) );
  AND U22217 ( .A(x[232]), .B(y[2027]), .Z(n21797) );
  NAND U22218 ( .A(n21798), .B(n21797), .Z(n21801) );
  NAND U22219 ( .A(n21799), .B(n22089), .Z(n21800) );
  NAND U22220 ( .A(n21801), .B(n21800), .Z(n21871) );
  XOR U22221 ( .A(n21872), .B(n21871), .Z(n21874) );
  AND U22222 ( .A(y[2021]), .B(x[234]), .Z(n21803) );
  NAND U22223 ( .A(y[2027]), .B(x[228]), .Z(n21802) );
  XNOR U22224 ( .A(n21803), .B(n21802), .Z(n21852) );
  AND U22225 ( .A(x[231]), .B(y[2024]), .Z(n21851) );
  XNOR U22226 ( .A(n21852), .B(n21851), .Z(n21859) );
  NAND U22227 ( .A(x[230]), .B(y[2025]), .Z(n21962) );
  XNOR U22228 ( .A(n21962), .B(n21857), .Z(n21858) );
  XNOR U22229 ( .A(n21859), .B(n21858), .Z(n21893) );
  AND U22230 ( .A(y[2029]), .B(x[226]), .Z(n21805) );
  NAND U22231 ( .A(y[2022]), .B(x[233]), .Z(n21804) );
  XNOR U22232 ( .A(n21805), .B(n21804), .Z(n21862) );
  AND U22233 ( .A(x[227]), .B(y[2028]), .Z(n21863) );
  XOR U22234 ( .A(n21862), .B(n21863), .Z(n21892) );
  AND U22235 ( .A(y[2030]), .B(x[225]), .Z(n21807) );
  NAND U22236 ( .A(y[2023]), .B(x[232]), .Z(n21806) );
  XNOR U22237 ( .A(n21807), .B(n21806), .Z(n21841) );
  AND U22238 ( .A(x[238]), .B(y[2017]), .Z(n21868) );
  XOR U22239 ( .A(o[239]), .B(n21868), .Z(n21840) );
  XOR U22240 ( .A(n21841), .B(n21840), .Z(n21891) );
  XOR U22241 ( .A(n21892), .B(n21891), .Z(n21894) );
  XOR U22242 ( .A(n21893), .B(n21894), .Z(n21873) );
  XNOR U22243 ( .A(n21874), .B(n21873), .Z(n21916) );
  NAND U22244 ( .A(n22200), .B(n21808), .Z(n21812) );
  NAND U22245 ( .A(n21810), .B(n21809), .Z(n21811) );
  AND U22246 ( .A(n21812), .B(n21811), .Z(n21915) );
  XOR U22247 ( .A(n21916), .B(n21915), .Z(n21917) );
  NAND U22248 ( .A(n21814), .B(n21813), .Z(n21818) );
  NAND U22249 ( .A(n21816), .B(n21815), .Z(n21817) );
  AND U22250 ( .A(n21818), .B(n21817), .Z(n21918) );
  XOR U22251 ( .A(n21917), .B(n21918), .Z(n21898) );
  XOR U22252 ( .A(n21897), .B(n21898), .Z(n21899) );
  XNOR U22253 ( .A(n21900), .B(n21899), .Z(n21928) );
  NAND U22254 ( .A(n21820), .B(n21819), .Z(n21824) );
  NAND U22255 ( .A(n21822), .B(n21821), .Z(n21823) );
  AND U22256 ( .A(n21824), .B(n21823), .Z(n21929) );
  XOR U22257 ( .A(n21928), .B(n21929), .Z(n21930) );
  XOR U22258 ( .A(n21931), .B(n21930), .Z(n21924) );
  OR U22259 ( .A(n21827), .B(n21825), .Z(n21831) );
  ANDN U22260 ( .B(n21827), .A(n21826), .Z(n21829) );
  OR U22261 ( .A(n21829), .B(n21828), .Z(n21830) );
  AND U22262 ( .A(n21831), .B(n21830), .Z(n21923) );
  NANDN U22263 ( .A(n21833), .B(n21832), .Z(n21837) );
  NAND U22264 ( .A(n21835), .B(n21834), .Z(n21836) );
  NAND U22265 ( .A(n21837), .B(n21836), .Z(n21922) );
  IV U22266 ( .A(n21922), .Z(n21921) );
  XOR U22267 ( .A(n21923), .B(n21921), .Z(n21838) );
  XNOR U22268 ( .A(n21924), .B(n21838), .Z(N496) );
  AND U22269 ( .A(x[232]), .B(y[2030]), .Z(n22201) );
  NAND U22270 ( .A(n22201), .B(n21839), .Z(n21843) );
  NAND U22271 ( .A(n21841), .B(n21840), .Z(n21842) );
  NAND U22272 ( .A(n21843), .B(n21842), .Z(n21992) );
  AND U22273 ( .A(x[239]), .B(y[2031]), .Z(n23962) );
  NAND U22274 ( .A(n23962), .B(n21844), .Z(n21848) );
  NAND U22275 ( .A(n21846), .B(n21845), .Z(n21847) );
  NAND U22276 ( .A(n21848), .B(n21847), .Z(n21991) );
  XOR U22277 ( .A(n21992), .B(n21991), .Z(n21994) );
  AND U22278 ( .A(x[234]), .B(y[2027]), .Z(n21850) );
  NAND U22279 ( .A(n21850), .B(n21849), .Z(n21854) );
  NAND U22280 ( .A(n21852), .B(n21851), .Z(n21853) );
  NAND U22281 ( .A(n21854), .B(n21853), .Z(n21949) );
  AND U22282 ( .A(x[224]), .B(y[2032]), .Z(n21971) );
  AND U22283 ( .A(x[240]), .B(y[2016]), .Z(n21972) );
  XOR U22284 ( .A(n21971), .B(n21972), .Z(n21974) );
  AND U22285 ( .A(x[239]), .B(y[2017]), .Z(n21959) );
  XOR U22286 ( .A(o[240]), .B(n21959), .Z(n21973) );
  XOR U22287 ( .A(n21974), .B(n21973), .Z(n21948) );
  NAND U22288 ( .A(y[2025]), .B(x[231]), .Z(n21855) );
  XNOR U22289 ( .A(n21856), .B(n21855), .Z(n21964) );
  AND U22290 ( .A(x[234]), .B(y[2022]), .Z(n21963) );
  XOR U22291 ( .A(n21964), .B(n21963), .Z(n21947) );
  XOR U22292 ( .A(n21948), .B(n21947), .Z(n21950) );
  XOR U22293 ( .A(n21949), .B(n21950), .Z(n21993) );
  XNOR U22294 ( .A(n21994), .B(n21993), .Z(n21944) );
  NANDN U22295 ( .A(n21857), .B(n21962), .Z(n21861) );
  NAND U22296 ( .A(n21859), .B(n21858), .Z(n21860) );
  NAND U22297 ( .A(n21861), .B(n21860), .Z(n21942) );
  NAND U22298 ( .A(x[233]), .B(y[2029]), .Z(n22702) );
  NANDN U22299 ( .A(n22702), .B(n22278), .Z(n21865) );
  NAND U22300 ( .A(n21863), .B(n21862), .Z(n21864) );
  AND U22301 ( .A(n21865), .B(n21864), .Z(n21982) );
  AND U22302 ( .A(y[2031]), .B(x[225]), .Z(n21867) );
  NAND U22303 ( .A(y[2024]), .B(x[232]), .Z(n21866) );
  XNOR U22304 ( .A(n21867), .B(n21866), .Z(n21968) );
  AND U22305 ( .A(o[239]), .B(n21868), .Z(n21967) );
  XOR U22306 ( .A(n21968), .B(n21967), .Z(n21980) );
  NAND U22307 ( .A(y[2018]), .B(x[238]), .Z(n21869) );
  XNOR U22308 ( .A(n21870), .B(n21869), .Z(n22003) );
  AND U22309 ( .A(x[228]), .B(y[2028]), .Z(n22004) );
  XOR U22310 ( .A(n22003), .B(n22004), .Z(n21979) );
  XOR U22311 ( .A(n21980), .B(n21979), .Z(n21981) );
  XOR U22312 ( .A(n21982), .B(n21981), .Z(n21941) );
  XOR U22313 ( .A(n21942), .B(n21941), .Z(n21943) );
  XOR U22314 ( .A(n21944), .B(n21943), .Z(n21985) );
  NAND U22315 ( .A(n21872), .B(n21871), .Z(n21876) );
  NAND U22316 ( .A(n21874), .B(n21873), .Z(n21875) );
  AND U22317 ( .A(n21876), .B(n21875), .Z(n21986) );
  XOR U22318 ( .A(n21985), .B(n21986), .Z(n21988) );
  NAND U22319 ( .A(n21878), .B(n21877), .Z(n21882) );
  NAND U22320 ( .A(n21880), .B(n21879), .Z(n21881) );
  NAND U22321 ( .A(n21882), .B(n21881), .Z(n22018) );
  AND U22322 ( .A(x[237]), .B(y[2020]), .Z(n22014) );
  NAND U22323 ( .A(n22541), .B(n22014), .Z(n21886) );
  NAND U22324 ( .A(n21884), .B(n21883), .Z(n21885) );
  NAND U22325 ( .A(n21886), .B(n21885), .Z(n22000) );
  AND U22326 ( .A(y[2030]), .B(x[226]), .Z(n21888) );
  NAND U22327 ( .A(y[2023]), .B(x[233]), .Z(n21887) );
  XNOR U22328 ( .A(n21888), .B(n21887), .Z(n22007) );
  AND U22329 ( .A(x[227]), .B(y[2029]), .Z(n22008) );
  XOR U22330 ( .A(n22007), .B(n22008), .Z(n21998) );
  AND U22331 ( .A(x[236]), .B(y[2020]), .Z(n22690) );
  AND U22332 ( .A(y[2027]), .B(x[229]), .Z(n21890) );
  NAND U22333 ( .A(y[2019]), .B(x[237]), .Z(n21889) );
  XNOR U22334 ( .A(n21890), .B(n21889), .Z(n21954) );
  XOR U22335 ( .A(n22690), .B(n21954), .Z(n21997) );
  XOR U22336 ( .A(n21998), .B(n21997), .Z(n21999) );
  XNOR U22337 ( .A(n22000), .B(n21999), .Z(n22015) );
  NAND U22338 ( .A(n21892), .B(n21891), .Z(n21896) );
  NAND U22339 ( .A(n21894), .B(n21893), .Z(n21895) );
  AND U22340 ( .A(n21896), .B(n21895), .Z(n22016) );
  XOR U22341 ( .A(n22015), .B(n22016), .Z(n22017) );
  XOR U22342 ( .A(n22018), .B(n22017), .Z(n21987) );
  XNOR U22343 ( .A(n21988), .B(n21987), .Z(n22029) );
  NAND U22344 ( .A(n21898), .B(n21897), .Z(n21902) );
  NAND U22345 ( .A(n21900), .B(n21899), .Z(n21901) );
  AND U22346 ( .A(n21902), .B(n21901), .Z(n22028) );
  XOR U22347 ( .A(n22029), .B(n22028), .Z(n22031) );
  NAND U22348 ( .A(n21904), .B(n21903), .Z(n21908) );
  NAND U22349 ( .A(n21906), .B(n21905), .Z(n21907) );
  NAND U22350 ( .A(n21908), .B(n21907), .Z(n21938) );
  NAND U22351 ( .A(n21910), .B(n21909), .Z(n21914) );
  NAND U22352 ( .A(n21912), .B(n21911), .Z(n21913) );
  NAND U22353 ( .A(n21914), .B(n21913), .Z(n21936) );
  NAND U22354 ( .A(n21916), .B(n21915), .Z(n21920) );
  NAND U22355 ( .A(n21918), .B(n21917), .Z(n21919) );
  AND U22356 ( .A(n21920), .B(n21919), .Z(n21935) );
  XOR U22357 ( .A(n21936), .B(n21935), .Z(n21937) );
  XOR U22358 ( .A(n21938), .B(n21937), .Z(n22030) );
  XNOR U22359 ( .A(n22031), .B(n22030), .Z(n22024) );
  OR U22360 ( .A(n21923), .B(n21921), .Z(n21927) );
  ANDN U22361 ( .B(n21923), .A(n21922), .Z(n21925) );
  OR U22362 ( .A(n21925), .B(n21924), .Z(n21926) );
  AND U22363 ( .A(n21927), .B(n21926), .Z(n22023) );
  NAND U22364 ( .A(n21929), .B(n21928), .Z(n21933) );
  NANDN U22365 ( .A(n21931), .B(n21930), .Z(n21932) );
  NAND U22366 ( .A(n21933), .B(n21932), .Z(n22022) );
  IV U22367 ( .A(n22022), .Z(n22021) );
  XOR U22368 ( .A(n22023), .B(n22021), .Z(n21934) );
  XNOR U22369 ( .A(n22024), .B(n21934), .Z(N497) );
  NAND U22370 ( .A(n21936), .B(n21935), .Z(n21940) );
  NAND U22371 ( .A(n21938), .B(n21937), .Z(n21939) );
  NAND U22372 ( .A(n21940), .B(n21939), .Z(n22132) );
  NAND U22373 ( .A(n21942), .B(n21941), .Z(n21946) );
  NAND U22374 ( .A(n21944), .B(n21943), .Z(n21945) );
  NAND U22375 ( .A(n21946), .B(n21945), .Z(n22044) );
  NAND U22376 ( .A(n21948), .B(n21947), .Z(n21952) );
  NAND U22377 ( .A(n21950), .B(n21949), .Z(n21951) );
  NAND U22378 ( .A(n21952), .B(n21951), .Z(n22126) );
  AND U22379 ( .A(x[237]), .B(y[2027]), .Z(n22934) );
  NAND U22380 ( .A(n22934), .B(n21953), .Z(n21956) );
  NAND U22381 ( .A(n21954), .B(n22690), .Z(n21955) );
  NAND U22382 ( .A(n21956), .B(n21955), .Z(n22074) );
  AND U22383 ( .A(y[2032]), .B(x[225]), .Z(n21958) );
  NAND U22384 ( .A(y[2024]), .B(x[233]), .Z(n21957) );
  XNOR U22385 ( .A(n21958), .B(n21957), .Z(n22095) );
  AND U22386 ( .A(o[240]), .B(n21959), .Z(n22094) );
  XOR U22387 ( .A(n22095), .B(n22094), .Z(n22072) );
  AND U22388 ( .A(y[2018]), .B(x[239]), .Z(n21961) );
  NAND U22389 ( .A(y[2021]), .B(x[236]), .Z(n21960) );
  XNOR U22390 ( .A(n21961), .B(n21960), .Z(n22048) );
  AND U22391 ( .A(x[238]), .B(y[2019]), .Z(n22047) );
  XOR U22392 ( .A(n22048), .B(n22047), .Z(n22071) );
  XOR U22393 ( .A(n22072), .B(n22071), .Z(n22073) );
  XOR U22394 ( .A(n22074), .B(n22073), .Z(n22124) );
  AND U22395 ( .A(x[231]), .B(y[2026]), .Z(n22106) );
  NANDN U22396 ( .A(n21962), .B(n22106), .Z(n21966) );
  NAND U22397 ( .A(n21964), .B(n21963), .Z(n21965) );
  NAND U22398 ( .A(n21966), .B(n21965), .Z(n22084) );
  NAND U22399 ( .A(x[232]), .B(y[2031]), .Z(n22784) );
  AND U22400 ( .A(x[225]), .B(y[2024]), .Z(n22179) );
  NANDN U22401 ( .A(n22784), .B(n22179), .Z(n21970) );
  NAND U22402 ( .A(n21968), .B(n21967), .Z(n21969) );
  NAND U22403 ( .A(n21970), .B(n21969), .Z(n22083) );
  XOR U22404 ( .A(n22084), .B(n22083), .Z(n22086) );
  NAND U22405 ( .A(n21972), .B(n21971), .Z(n21976) );
  NAND U22406 ( .A(n21974), .B(n21973), .Z(n21975) );
  NAND U22407 ( .A(n21976), .B(n21975), .Z(n22080) );
  AND U22408 ( .A(x[224]), .B(y[2033]), .Z(n22062) );
  AND U22409 ( .A(x[241]), .B(y[2016]), .Z(n22061) );
  XOR U22410 ( .A(n22062), .B(n22061), .Z(n22064) );
  AND U22411 ( .A(x[240]), .B(y[2017]), .Z(n22058) );
  XOR U22412 ( .A(n22058), .B(o[241]), .Z(n22063) );
  XOR U22413 ( .A(n22064), .B(n22063), .Z(n22078) );
  AND U22414 ( .A(y[2031]), .B(x[226]), .Z(n21978) );
  NAND U22415 ( .A(y[2023]), .B(x[234]), .Z(n21977) );
  XNOR U22416 ( .A(n21978), .B(n21977), .Z(n22099) );
  AND U22417 ( .A(x[227]), .B(y[2030]), .Z(n22100) );
  XOR U22418 ( .A(n22099), .B(n22100), .Z(n22077) );
  XOR U22419 ( .A(n22078), .B(n22077), .Z(n22079) );
  XOR U22420 ( .A(n22080), .B(n22079), .Z(n22085) );
  XOR U22421 ( .A(n22086), .B(n22085), .Z(n22123) );
  XOR U22422 ( .A(n22124), .B(n22123), .Z(n22125) );
  XNOR U22423 ( .A(n22126), .B(n22125), .Z(n22041) );
  NAND U22424 ( .A(n21980), .B(n21979), .Z(n21984) );
  NANDN U22425 ( .A(n21982), .B(n21981), .Z(n21983) );
  AND U22426 ( .A(n21984), .B(n21983), .Z(n22042) );
  XOR U22427 ( .A(n22041), .B(n22042), .Z(n22043) );
  XNOR U22428 ( .A(n22044), .B(n22043), .Z(n22130) );
  NAND U22429 ( .A(n21986), .B(n21985), .Z(n21990) );
  NAND U22430 ( .A(n21988), .B(n21987), .Z(n21989) );
  AND U22431 ( .A(n21990), .B(n21989), .Z(n22038) );
  NAND U22432 ( .A(n21992), .B(n21991), .Z(n21996) );
  NAND U22433 ( .A(n21994), .B(n21993), .Z(n21995) );
  NAND U22434 ( .A(n21996), .B(n21995), .Z(n22120) );
  NAND U22435 ( .A(n21998), .B(n21997), .Z(n22002) );
  NAND U22436 ( .A(n22000), .B(n21999), .Z(n22001) );
  NAND U22437 ( .A(n22002), .B(n22001), .Z(n22118) );
  AND U22438 ( .A(x[238]), .B(y[2021]), .Z(n22311) );
  NAND U22439 ( .A(n22541), .B(n22311), .Z(n22006) );
  NAND U22440 ( .A(n22004), .B(n22003), .Z(n22005) );
  NAND U22441 ( .A(n22006), .B(n22005), .Z(n22112) );
  AND U22442 ( .A(x[233]), .B(y[2030]), .Z(n22915) );
  NANDN U22443 ( .A(n22098), .B(n22915), .Z(n22010) );
  NAND U22444 ( .A(n22008), .B(n22007), .Z(n22009) );
  NAND U22445 ( .A(n22010), .B(n22009), .Z(n22111) );
  XOR U22446 ( .A(n22112), .B(n22111), .Z(n22114) );
  AND U22447 ( .A(y[2028]), .B(x[229]), .Z(n22162) );
  NAND U22448 ( .A(y[2025]), .B(x[232]), .Z(n22011) );
  XNOR U22449 ( .A(n22162), .B(n22011), .Z(n22090) );
  XOR U22450 ( .A(n22090), .B(n22012), .Z(n22105) );
  XOR U22451 ( .A(n22106), .B(n22105), .Z(n22108) );
  NAND U22452 ( .A(y[2029]), .B(x[228]), .Z(n22013) );
  XNOR U22453 ( .A(n22014), .B(n22013), .Z(n22052) );
  AND U22454 ( .A(x[235]), .B(y[2022]), .Z(n22053) );
  XOR U22455 ( .A(n22052), .B(n22053), .Z(n22107) );
  XOR U22456 ( .A(n22108), .B(n22107), .Z(n22113) );
  XOR U22457 ( .A(n22114), .B(n22113), .Z(n22117) );
  XOR U22458 ( .A(n22118), .B(n22117), .Z(n22119) );
  XNOR U22459 ( .A(n22120), .B(n22119), .Z(n22036) );
  NAND U22460 ( .A(n22016), .B(n22015), .Z(n22020) );
  NAND U22461 ( .A(n22018), .B(n22017), .Z(n22019) );
  NAND U22462 ( .A(n22020), .B(n22019), .Z(n22035) );
  XOR U22463 ( .A(n22036), .B(n22035), .Z(n22037) );
  XOR U22464 ( .A(n22038), .B(n22037), .Z(n22129) );
  XOR U22465 ( .A(n22130), .B(n22129), .Z(n22131) );
  XOR U22466 ( .A(n22132), .B(n22131), .Z(n22138) );
  OR U22467 ( .A(n22023), .B(n22021), .Z(n22027) );
  ANDN U22468 ( .B(n22023), .A(n22022), .Z(n22025) );
  OR U22469 ( .A(n22025), .B(n22024), .Z(n22026) );
  AND U22470 ( .A(n22027), .B(n22026), .Z(n22136) );
  NAND U22471 ( .A(n22029), .B(n22028), .Z(n22033) );
  NAND U22472 ( .A(n22031), .B(n22030), .Z(n22032) );
  AND U22473 ( .A(n22033), .B(n22032), .Z(n22137) );
  IV U22474 ( .A(n22137), .Z(n22135) );
  XOR U22475 ( .A(n22136), .B(n22135), .Z(n22034) );
  XNOR U22476 ( .A(n22138), .B(n22034), .Z(N498) );
  NAND U22477 ( .A(n22036), .B(n22035), .Z(n22040) );
  NANDN U22478 ( .A(n22038), .B(n22037), .Z(n22039) );
  AND U22479 ( .A(n22040), .B(n22039), .Z(n22251) );
  NAND U22480 ( .A(n22042), .B(n22041), .Z(n22046) );
  NAND U22481 ( .A(n22044), .B(n22043), .Z(n22045) );
  AND U22482 ( .A(n22046), .B(n22045), .Z(n22249) );
  AND U22483 ( .A(x[236]), .B(y[2018]), .Z(n22388) );
  AND U22484 ( .A(x[239]), .B(y[2021]), .Z(n22286) );
  NAND U22485 ( .A(n22388), .B(n22286), .Z(n22050) );
  NAND U22486 ( .A(n22048), .B(n22047), .Z(n22049) );
  NAND U22487 ( .A(n22050), .B(n22049), .Z(n22227) );
  NAND U22488 ( .A(n23307), .B(n22051), .Z(n22055) );
  NAND U22489 ( .A(n22053), .B(n22052), .Z(n22054) );
  NAND U22490 ( .A(n22055), .B(n22054), .Z(n22218) );
  AND U22491 ( .A(y[2033]), .B(x[225]), .Z(n22057) );
  NAND U22492 ( .A(y[2024]), .B(x[234]), .Z(n22056) );
  XNOR U22493 ( .A(n22057), .B(n22056), .Z(n22180) );
  AND U22494 ( .A(n22058), .B(o[241]), .Z(n22181) );
  XOR U22495 ( .A(n22180), .B(n22181), .Z(n22216) );
  AND U22496 ( .A(y[2019]), .B(x[239]), .Z(n22060) );
  NAND U22497 ( .A(y[2025]), .B(x[233]), .Z(n22059) );
  XNOR U22498 ( .A(n22060), .B(n22059), .Z(n22171) );
  AND U22499 ( .A(x[238]), .B(y[2020]), .Z(n22172) );
  XOR U22500 ( .A(n22171), .B(n22172), .Z(n22215) );
  XOR U22501 ( .A(n22216), .B(n22215), .Z(n22217) );
  XOR U22502 ( .A(n22218), .B(n22217), .Z(n22228) );
  XOR U22503 ( .A(n22227), .B(n22228), .Z(n22230) );
  NAND U22504 ( .A(n22062), .B(n22061), .Z(n22066) );
  NAND U22505 ( .A(n22064), .B(n22063), .Z(n22065) );
  NAND U22506 ( .A(n22066), .B(n22065), .Z(n22239) );
  AND U22507 ( .A(y[2018]), .B(x[240]), .Z(n22068) );
  NAND U22508 ( .A(y[2023]), .B(x[235]), .Z(n22067) );
  XNOR U22509 ( .A(n22068), .B(n22067), .Z(n22167) );
  AND U22510 ( .A(x[226]), .B(y[2032]), .Z(n22168) );
  XOR U22511 ( .A(n22167), .B(n22168), .Z(n22240) );
  XOR U22512 ( .A(n22239), .B(n22240), .Z(n22242) );
  AND U22513 ( .A(y[2029]), .B(x[229]), .Z(n22294) );
  NAND U22514 ( .A(y[2028]), .B(x[230]), .Z(n22069) );
  XNOR U22515 ( .A(n22294), .B(n22069), .Z(n22164) );
  NAND U22516 ( .A(y[2030]), .B(x[228]), .Z(n22070) );
  XNOR U22517 ( .A(n22920), .B(n22070), .Z(n22203) );
  AND U22518 ( .A(x[231]), .B(y[2027]), .Z(n22202) );
  XOR U22519 ( .A(n22203), .B(n22202), .Z(n22163) );
  XOR U22520 ( .A(n22164), .B(n22163), .Z(n22241) );
  XOR U22521 ( .A(n22242), .B(n22241), .Z(n22229) );
  XNOR U22522 ( .A(n22230), .B(n22229), .Z(n22150) );
  NAND U22523 ( .A(n22072), .B(n22071), .Z(n22076) );
  NAND U22524 ( .A(n22074), .B(n22073), .Z(n22075) );
  AND U22525 ( .A(n22076), .B(n22075), .Z(n22222) );
  NAND U22526 ( .A(n22078), .B(n22077), .Z(n22082) );
  NAND U22527 ( .A(n22080), .B(n22079), .Z(n22081) );
  AND U22528 ( .A(n22082), .B(n22081), .Z(n22221) );
  XOR U22529 ( .A(n22222), .B(n22221), .Z(n22224) );
  NAND U22530 ( .A(n22084), .B(n22083), .Z(n22088) );
  NAND U22531 ( .A(n22086), .B(n22085), .Z(n22087) );
  AND U22532 ( .A(n22088), .B(n22087), .Z(n22223) );
  XOR U22533 ( .A(n22224), .B(n22223), .Z(n22149) );
  XOR U22534 ( .A(n22150), .B(n22149), .Z(n22152) );
  AND U22535 ( .A(x[232]), .B(y[2028]), .Z(n22428) );
  NAND U22536 ( .A(n22428), .B(n22089), .Z(n22093) );
  NANDN U22537 ( .A(n22091), .B(n22090), .Z(n22092) );
  NAND U22538 ( .A(n22093), .B(n22092), .Z(n22234) );
  AND U22539 ( .A(x[233]), .B(y[2032]), .Z(n23081) );
  NAND U22540 ( .A(n23081), .B(n22179), .Z(n22097) );
  NAND U22541 ( .A(n22095), .B(n22094), .Z(n22096) );
  NAND U22542 ( .A(n22097), .B(n22096), .Z(n22233) );
  XOR U22543 ( .A(n22234), .B(n22233), .Z(n22236) );
  AND U22544 ( .A(x[234]), .B(y[2031]), .Z(n22943) );
  NANDN U22545 ( .A(n22098), .B(n22943), .Z(n22102) );
  NAND U22546 ( .A(n22100), .B(n22099), .Z(n22101) );
  NAND U22547 ( .A(n22102), .B(n22101), .Z(n22212) );
  AND U22548 ( .A(x[224]), .B(y[2034]), .Z(n22184) );
  AND U22549 ( .A(x[242]), .B(y[2016]), .Z(n22185) );
  XOR U22550 ( .A(n22184), .B(n22185), .Z(n22187) );
  AND U22551 ( .A(x[241]), .B(y[2017]), .Z(n22206) );
  XOR U22552 ( .A(o[242]), .B(n22206), .Z(n22186) );
  XOR U22553 ( .A(n22187), .B(n22186), .Z(n22210) );
  AND U22554 ( .A(y[2021]), .B(x[237]), .Z(n22104) );
  NAND U22555 ( .A(y[2031]), .B(x[227]), .Z(n22103) );
  XNOR U22556 ( .A(n22104), .B(n22103), .Z(n22192) );
  AND U22557 ( .A(x[236]), .B(y[2022]), .Z(n22193) );
  XOR U22558 ( .A(n22192), .B(n22193), .Z(n22209) );
  XOR U22559 ( .A(n22210), .B(n22209), .Z(n22211) );
  XOR U22560 ( .A(n22212), .B(n22211), .Z(n22235) );
  XNOR U22561 ( .A(n22236), .B(n22235), .Z(n22156) );
  NAND U22562 ( .A(n22106), .B(n22105), .Z(n22110) );
  NAND U22563 ( .A(n22108), .B(n22107), .Z(n22109) );
  AND U22564 ( .A(n22110), .B(n22109), .Z(n22155) );
  XOR U22565 ( .A(n22156), .B(n22155), .Z(n22157) );
  NAND U22566 ( .A(n22112), .B(n22111), .Z(n22116) );
  NAND U22567 ( .A(n22114), .B(n22113), .Z(n22115) );
  AND U22568 ( .A(n22116), .B(n22115), .Z(n22158) );
  XOR U22569 ( .A(n22157), .B(n22158), .Z(n22151) );
  XNOR U22570 ( .A(n22152), .B(n22151), .Z(n22146) );
  NAND U22571 ( .A(n22118), .B(n22117), .Z(n22122) );
  NAND U22572 ( .A(n22120), .B(n22119), .Z(n22121) );
  NAND U22573 ( .A(n22122), .B(n22121), .Z(n22144) );
  NAND U22574 ( .A(n22124), .B(n22123), .Z(n22128) );
  NAND U22575 ( .A(n22126), .B(n22125), .Z(n22127) );
  NAND U22576 ( .A(n22128), .B(n22127), .Z(n22143) );
  XOR U22577 ( .A(n22144), .B(n22143), .Z(n22145) );
  XOR U22578 ( .A(n22146), .B(n22145), .Z(n22248) );
  XOR U22579 ( .A(n22249), .B(n22248), .Z(n22250) );
  XNOR U22580 ( .A(n22251), .B(n22250), .Z(n22247) );
  NAND U22581 ( .A(n22130), .B(n22129), .Z(n22134) );
  NAND U22582 ( .A(n22132), .B(n22131), .Z(n22133) );
  NAND U22583 ( .A(n22134), .B(n22133), .Z(n22246) );
  NANDN U22584 ( .A(n22135), .B(n22136), .Z(n22141) );
  NOR U22585 ( .A(n22137), .B(n22136), .Z(n22139) );
  OR U22586 ( .A(n22139), .B(n22138), .Z(n22140) );
  AND U22587 ( .A(n22141), .B(n22140), .Z(n22245) );
  XOR U22588 ( .A(n22246), .B(n22245), .Z(n22142) );
  XNOR U22589 ( .A(n22247), .B(n22142), .Z(N499) );
  NAND U22590 ( .A(n22144), .B(n22143), .Z(n22148) );
  NAND U22591 ( .A(n22146), .B(n22145), .Z(n22147) );
  NAND U22592 ( .A(n22148), .B(n22147), .Z(n22365) );
  NAND U22593 ( .A(n22150), .B(n22149), .Z(n22154) );
  NAND U22594 ( .A(n22152), .B(n22151), .Z(n22153) );
  AND U22595 ( .A(n22154), .B(n22153), .Z(n22363) );
  NAND U22596 ( .A(n22156), .B(n22155), .Z(n22160) );
  NAND U22597 ( .A(n22158), .B(n22157), .Z(n22159) );
  NAND U22598 ( .A(n22160), .B(n22159), .Z(n22258) );
  AND U22599 ( .A(x[230]), .B(y[2029]), .Z(n22161) );
  NAND U22600 ( .A(n22162), .B(n22161), .Z(n22166) );
  NAND U22601 ( .A(n22164), .B(n22163), .Z(n22165) );
  NAND U22602 ( .A(n22166), .B(n22165), .Z(n22347) );
  AND U22603 ( .A(x[240]), .B(y[2023]), .Z(n22706) );
  NAND U22604 ( .A(n22706), .B(n22541), .Z(n22170) );
  NAND U22605 ( .A(n22168), .B(n22167), .Z(n22169) );
  NAND U22606 ( .A(n22170), .B(n22169), .Z(n22345) );
  AND U22607 ( .A(x[239]), .B(y[2025]), .Z(n22948) );
  NAND U22608 ( .A(n22948), .B(n22273), .Z(n22174) );
  NAND U22609 ( .A(n22172), .B(n22171), .Z(n22173) );
  NAND U22610 ( .A(n22174), .B(n22173), .Z(n22263) );
  AND U22611 ( .A(y[2034]), .B(x[225]), .Z(n22176) );
  NAND U22612 ( .A(y[2027]), .B(x[232]), .Z(n22175) );
  XNOR U22613 ( .A(n22176), .B(n22175), .Z(n22312) );
  XOR U22614 ( .A(n22311), .B(n22312), .Z(n22262) );
  AND U22615 ( .A(y[2022]), .B(x[237]), .Z(n22178) );
  NAND U22616 ( .A(y[2033]), .B(x[226]), .Z(n22177) );
  XNOR U22617 ( .A(n22178), .B(n22177), .Z(n22280) );
  XOR U22618 ( .A(n22280), .B(n22279), .Z(n22261) );
  XOR U22619 ( .A(n22262), .B(n22261), .Z(n22264) );
  XOR U22620 ( .A(n22263), .B(n22264), .Z(n22344) );
  XOR U22621 ( .A(n22345), .B(n22344), .Z(n22346) );
  XNOR U22622 ( .A(n22347), .B(n22346), .Z(n22256) );
  AND U22623 ( .A(x[234]), .B(y[2033]), .Z(n23399) );
  NAND U22624 ( .A(n23399), .B(n22179), .Z(n22183) );
  NAND U22625 ( .A(n22181), .B(n22180), .Z(n22182) );
  NAND U22626 ( .A(n22183), .B(n22182), .Z(n22322) );
  NAND U22627 ( .A(n22185), .B(n22184), .Z(n22189) );
  NAND U22628 ( .A(n22187), .B(n22186), .Z(n22188) );
  NAND U22629 ( .A(n22189), .B(n22188), .Z(n22320) );
  AND U22630 ( .A(y[2019]), .B(x[240]), .Z(n22999) );
  NAND U22631 ( .A(y[2026]), .B(x[233]), .Z(n22190) );
  XNOR U22632 ( .A(n22999), .B(n22190), .Z(n22275) );
  AND U22633 ( .A(x[239]), .B(y[2020]), .Z(n22274) );
  XOR U22634 ( .A(n22275), .B(n22274), .Z(n22321) );
  XOR U22635 ( .A(n22320), .B(n22321), .Z(n22323) );
  XNOR U22636 ( .A(n22322), .B(n22323), .Z(n22340) );
  AND U22637 ( .A(x[237]), .B(y[2031]), .Z(n23594) );
  NAND U22638 ( .A(n22191), .B(n23594), .Z(n22195) );
  NAND U22639 ( .A(n22193), .B(n22192), .Z(n22194) );
  NAND U22640 ( .A(n22195), .B(n22194), .Z(n22328) );
  AND U22641 ( .A(y[2025]), .B(x[234]), .Z(n22197) );
  NAND U22642 ( .A(y[2018]), .B(x[241]), .Z(n22196) );
  XNOR U22643 ( .A(n22197), .B(n22196), .Z(n22317) );
  AND U22644 ( .A(x[242]), .B(y[2017]), .Z(n22293) );
  XOR U22645 ( .A(o[243]), .B(n22293), .Z(n22316) );
  XOR U22646 ( .A(n22317), .B(n22316), .Z(n22327) );
  NAND U22647 ( .A(y[2032]), .B(x[227]), .Z(n22198) );
  XNOR U22648 ( .A(n22199), .B(n22198), .Z(n22287) );
  XOR U22649 ( .A(n22327), .B(n22326), .Z(n22329) );
  XNOR U22650 ( .A(n22328), .B(n22329), .Z(n22339) );
  NAND U22651 ( .A(n22201), .B(n22200), .Z(n22205) );
  NAND U22652 ( .A(n22203), .B(n22202), .Z(n22204) );
  NAND U22653 ( .A(n22205), .B(n22204), .Z(n22269) );
  AND U22654 ( .A(o[242]), .B(n22206), .Z(n22301) );
  AND U22655 ( .A(x[224]), .B(y[2035]), .Z(n22298) );
  AND U22656 ( .A(x[243]), .B(y[2016]), .Z(n22299) );
  XOR U22657 ( .A(n22298), .B(n22299), .Z(n22300) );
  XOR U22658 ( .A(n22301), .B(n22300), .Z(n22268) );
  AND U22659 ( .A(x[228]), .B(y[2031]), .Z(n22442) );
  AND U22660 ( .A(y[2030]), .B(x[229]), .Z(n22208) );
  NAND U22661 ( .A(y[2029]), .B(x[230]), .Z(n22207) );
  XNOR U22662 ( .A(n22208), .B(n22207), .Z(n22295) );
  XOR U22663 ( .A(n22442), .B(n22295), .Z(n22267) );
  XOR U22664 ( .A(n22268), .B(n22267), .Z(n22270) );
  XNOR U22665 ( .A(n22269), .B(n22270), .Z(n22338) );
  XOR U22666 ( .A(n22339), .B(n22338), .Z(n22341) );
  XNOR U22667 ( .A(n22340), .B(n22341), .Z(n22334) );
  NAND U22668 ( .A(n22210), .B(n22209), .Z(n22214) );
  NAND U22669 ( .A(n22212), .B(n22211), .Z(n22213) );
  NAND U22670 ( .A(n22214), .B(n22213), .Z(n22333) );
  NAND U22671 ( .A(n22216), .B(n22215), .Z(n22220) );
  NAND U22672 ( .A(n22218), .B(n22217), .Z(n22219) );
  NAND U22673 ( .A(n22220), .B(n22219), .Z(n22332) );
  XOR U22674 ( .A(n22333), .B(n22332), .Z(n22335) );
  XNOR U22675 ( .A(n22334), .B(n22335), .Z(n22255) );
  XOR U22676 ( .A(n22256), .B(n22255), .Z(n22257) );
  XOR U22677 ( .A(n22258), .B(n22257), .Z(n22359) );
  NAND U22678 ( .A(n22222), .B(n22221), .Z(n22226) );
  NAND U22679 ( .A(n22224), .B(n22223), .Z(n22225) );
  AND U22680 ( .A(n22226), .B(n22225), .Z(n22356) );
  NAND U22681 ( .A(n22228), .B(n22227), .Z(n22232) );
  NAND U22682 ( .A(n22230), .B(n22229), .Z(n22231) );
  NAND U22683 ( .A(n22232), .B(n22231), .Z(n22352) );
  NAND U22684 ( .A(n22234), .B(n22233), .Z(n22238) );
  NAND U22685 ( .A(n22236), .B(n22235), .Z(n22237) );
  NAND U22686 ( .A(n22238), .B(n22237), .Z(n22351) );
  NAND U22687 ( .A(n22240), .B(n22239), .Z(n22244) );
  NAND U22688 ( .A(n22242), .B(n22241), .Z(n22243) );
  NAND U22689 ( .A(n22244), .B(n22243), .Z(n22350) );
  XNOR U22690 ( .A(n22351), .B(n22350), .Z(n22353) );
  XNOR U22691 ( .A(n22356), .B(n22357), .Z(n22358) );
  XOR U22692 ( .A(n22363), .B(n22362), .Z(n22364) );
  XOR U22693 ( .A(n22365), .B(n22364), .Z(n22371) );
  NAND U22694 ( .A(n22249), .B(n22248), .Z(n22253) );
  NAND U22695 ( .A(n22251), .B(n22250), .Z(n22252) );
  AND U22696 ( .A(n22253), .B(n22252), .Z(n22370) );
  IV U22697 ( .A(n22370), .Z(n22368) );
  XOR U22698 ( .A(n22369), .B(n22368), .Z(n22254) );
  XNOR U22699 ( .A(n22371), .B(n22254), .Z(N500) );
  NAND U22700 ( .A(n22256), .B(n22255), .Z(n22260) );
  NAND U22701 ( .A(n22258), .B(n22257), .Z(n22259) );
  AND U22702 ( .A(n22260), .B(n22259), .Z(n22480) );
  NAND U22703 ( .A(n22262), .B(n22261), .Z(n22266) );
  NAND U22704 ( .A(n22264), .B(n22263), .Z(n22265) );
  NAND U22705 ( .A(n22266), .B(n22265), .Z(n22377) );
  NAND U22706 ( .A(n22268), .B(n22267), .Z(n22272) );
  NAND U22707 ( .A(n22270), .B(n22269), .Z(n22271) );
  NAND U22708 ( .A(n22272), .B(n22271), .Z(n22376) );
  XOR U22709 ( .A(n22377), .B(n22376), .Z(n22379) );
  AND U22710 ( .A(x[240]), .B(y[2026]), .Z(n23221) );
  NAND U22711 ( .A(n23221), .B(n22273), .Z(n22277) );
  NAND U22712 ( .A(n22275), .B(n22274), .Z(n22276) );
  NAND U22713 ( .A(n22277), .B(n22276), .Z(n22417) );
  AND U22714 ( .A(x[237]), .B(y[2033]), .Z(n23850) );
  NAND U22715 ( .A(n23850), .B(n22278), .Z(n22282) );
  NAND U22716 ( .A(n22280), .B(n22279), .Z(n22281) );
  NAND U22717 ( .A(n22282), .B(n22281), .Z(n22462) );
  AND U22718 ( .A(y[2020]), .B(x[240]), .Z(n22284) );
  NAND U22719 ( .A(y[2026]), .B(x[234]), .Z(n22283) );
  XNOR U22720 ( .A(n22284), .B(n22283), .Z(n22423) );
  AND U22721 ( .A(x[226]), .B(y[2034]), .Z(n22424) );
  XOR U22722 ( .A(n22423), .B(n22424), .Z(n22460) );
  NAND U22723 ( .A(y[2027]), .B(x[233]), .Z(n22285) );
  XNOR U22724 ( .A(n22286), .B(n22285), .Z(n22399) );
  AND U22725 ( .A(x[238]), .B(y[2022]), .Z(n22400) );
  XOR U22726 ( .A(n22399), .B(n22400), .Z(n22459) );
  XOR U22727 ( .A(n22460), .B(n22459), .Z(n22461) );
  XOR U22728 ( .A(n22462), .B(n22461), .Z(n22416) );
  XOR U22729 ( .A(n22417), .B(n22416), .Z(n22419) );
  AND U22730 ( .A(x[235]), .B(y[2032]), .Z(n23401) );
  IV U22731 ( .A(n23401), .Z(n23263) );
  NANDN U22732 ( .A(n23263), .B(n22568), .Z(n22290) );
  NANDN U22733 ( .A(n22288), .B(n22287), .Z(n22289) );
  NAND U22734 ( .A(n22290), .B(n22289), .Z(n22468) );
  AND U22735 ( .A(y[2025]), .B(x[235]), .Z(n22292) );
  NAND U22736 ( .A(y[2035]), .B(x[225]), .Z(n22291) );
  XNOR U22737 ( .A(n22292), .B(n22291), .Z(n22395) );
  AND U22738 ( .A(x[243]), .B(y[2017]), .Z(n22403) );
  XOR U22739 ( .A(o[244]), .B(n22403), .Z(n22394) );
  XOR U22740 ( .A(n22395), .B(n22394), .Z(n22466) );
  AND U22741 ( .A(x[224]), .B(y[2036]), .Z(n22447) );
  AND U22742 ( .A(x[244]), .B(y[2016]), .Z(n22448) );
  XOR U22743 ( .A(n22447), .B(n22448), .Z(n22450) );
  AND U22744 ( .A(o[243]), .B(n22293), .Z(n22449) );
  XOR U22745 ( .A(n22450), .B(n22449), .Z(n22465) );
  XOR U22746 ( .A(n22466), .B(n22465), .Z(n22467) );
  XOR U22747 ( .A(n22468), .B(n22467), .Z(n22418) );
  XOR U22748 ( .A(n22419), .B(n22418), .Z(n22378) );
  XOR U22749 ( .A(n22379), .B(n22378), .Z(n22474) );
  NAND U22750 ( .A(x[230]), .B(y[2030]), .Z(n22383) );
  NANDN U22751 ( .A(n22383), .B(n22294), .Z(n22297) );
  NAND U22752 ( .A(n22295), .B(n22442), .Z(n22296) );
  NAND U22753 ( .A(n22297), .B(n22296), .Z(n22407) );
  NAND U22754 ( .A(n22299), .B(n22298), .Z(n22303) );
  NAND U22755 ( .A(n22301), .B(n22300), .Z(n22302) );
  NAND U22756 ( .A(n22303), .B(n22302), .Z(n22405) );
  AND U22757 ( .A(y[2018]), .B(x[242]), .Z(n22305) );
  NAND U22758 ( .A(y[2024]), .B(x[236]), .Z(n22304) );
  XNOR U22759 ( .A(n22305), .B(n22304), .Z(n22389) );
  AND U22760 ( .A(x[241]), .B(y[2019]), .Z(n22390) );
  XOR U22761 ( .A(n22389), .B(n22390), .Z(n22404) );
  XOR U22762 ( .A(n22405), .B(n22404), .Z(n22406) );
  XOR U22763 ( .A(n22407), .B(n22406), .Z(n22411) );
  AND U22764 ( .A(y[2023]), .B(x[237]), .Z(n22307) );
  NAND U22765 ( .A(y[2033]), .B(x[227]), .Z(n22306) );
  XNOR U22766 ( .A(n22307), .B(n22306), .Z(n22429) );
  XNOR U22767 ( .A(n22429), .B(n22428), .Z(n22385) );
  AND U22768 ( .A(y[2031]), .B(x[229]), .Z(n22309) );
  NAND U22769 ( .A(y[2032]), .B(x[228]), .Z(n22308) );
  XNOR U22770 ( .A(n22309), .B(n22308), .Z(n22444) );
  AND U22771 ( .A(x[231]), .B(y[2029]), .Z(n22443) );
  XNOR U22772 ( .A(n22444), .B(n22443), .Z(n22382) );
  XOR U22773 ( .A(n22383), .B(n22382), .Z(n22384) );
  XNOR U22774 ( .A(n22385), .B(n22384), .Z(n22455) );
  AND U22775 ( .A(x[232]), .B(y[2034]), .Z(n23553) );
  AND U22776 ( .A(x[225]), .B(y[2027]), .Z(n22310) );
  NAND U22777 ( .A(n23553), .B(n22310), .Z(n22314) );
  NAND U22778 ( .A(n22312), .B(n22311), .Z(n22313) );
  NAND U22779 ( .A(n22314), .B(n22313), .Z(n22454) );
  NAND U22780 ( .A(x[241]), .B(y[2025]), .Z(n23229) );
  NANDN U22781 ( .A(n23229), .B(n22315), .Z(n22319) );
  NAND U22782 ( .A(n22317), .B(n22316), .Z(n22318) );
  NAND U22783 ( .A(n22319), .B(n22318), .Z(n22453) );
  XOR U22784 ( .A(n22454), .B(n22453), .Z(n22456) );
  XNOR U22785 ( .A(n22455), .B(n22456), .Z(n22410) );
  NAND U22786 ( .A(n22321), .B(n22320), .Z(n22325) );
  NAND U22787 ( .A(n22323), .B(n22322), .Z(n22324) );
  AND U22788 ( .A(n22325), .B(n22324), .Z(n22412) );
  XOR U22789 ( .A(n22413), .B(n22412), .Z(n22472) );
  NAND U22790 ( .A(n22327), .B(n22326), .Z(n22331) );
  NAND U22791 ( .A(n22329), .B(n22328), .Z(n22330) );
  AND U22792 ( .A(n22331), .B(n22330), .Z(n22471) );
  XOR U22793 ( .A(n22472), .B(n22471), .Z(n22473) );
  NAND U22794 ( .A(n22333), .B(n22332), .Z(n22337) );
  NAND U22795 ( .A(n22335), .B(n22334), .Z(n22336) );
  AND U22796 ( .A(n22337), .B(n22336), .Z(n22486) );
  NAND U22797 ( .A(n22339), .B(n22338), .Z(n22343) );
  NAND U22798 ( .A(n22341), .B(n22340), .Z(n22342) );
  AND U22799 ( .A(n22343), .B(n22342), .Z(n22484) );
  NAND U22800 ( .A(n22345), .B(n22344), .Z(n22349) );
  NAND U22801 ( .A(n22347), .B(n22346), .Z(n22348) );
  AND U22802 ( .A(n22349), .B(n22348), .Z(n22483) );
  XNOR U22803 ( .A(n22486), .B(n22485), .Z(n22477) );
  XOR U22804 ( .A(n22478), .B(n22477), .Z(n22479) );
  XOR U22805 ( .A(n22480), .B(n22479), .Z(n22495) );
  NAND U22806 ( .A(n22351), .B(n22350), .Z(n22355) );
  NANDN U22807 ( .A(n22353), .B(n22352), .Z(n22354) );
  AND U22808 ( .A(n22355), .B(n22354), .Z(n22493) );
  NANDN U22809 ( .A(n22357), .B(n22356), .Z(n22361) );
  NANDN U22810 ( .A(n22359), .B(n22358), .Z(n22360) );
  AND U22811 ( .A(n22361), .B(n22360), .Z(n22492) );
  XOR U22812 ( .A(n22493), .B(n22492), .Z(n22494) );
  NAND U22813 ( .A(n22363), .B(n22362), .Z(n22367) );
  NAND U22814 ( .A(n22365), .B(n22364), .Z(n22366) );
  NAND U22815 ( .A(n22367), .B(n22366), .Z(n22490) );
  NANDN U22816 ( .A(n22368), .B(n22369), .Z(n22374) );
  NOR U22817 ( .A(n22370), .B(n22369), .Z(n22372) );
  OR U22818 ( .A(n22372), .B(n22371), .Z(n22373) );
  AND U22819 ( .A(n22374), .B(n22373), .Z(n22489) );
  XOR U22820 ( .A(n22490), .B(n22489), .Z(n22375) );
  XNOR U22821 ( .A(n22491), .B(n22375), .Z(N501) );
  NAND U22822 ( .A(n22377), .B(n22376), .Z(n22381) );
  NAND U22823 ( .A(n22379), .B(n22378), .Z(n22380) );
  NAND U22824 ( .A(n22381), .B(n22380), .Z(n22507) );
  NAND U22825 ( .A(n22383), .B(n22382), .Z(n22387) );
  NAND U22826 ( .A(n22385), .B(n22384), .Z(n22386) );
  NAND U22827 ( .A(n22387), .B(n22386), .Z(n22609) );
  AND U22828 ( .A(x[242]), .B(y[2024]), .Z(n23228) );
  NAND U22829 ( .A(n23228), .B(n22388), .Z(n22392) );
  NAND U22830 ( .A(n22390), .B(n22389), .Z(n22391) );
  NAND U22831 ( .A(n22392), .B(n22391), .Z(n22591) );
  AND U22832 ( .A(x[235]), .B(y[2035]), .Z(n23988) );
  AND U22833 ( .A(x[225]), .B(y[2025]), .Z(n22393) );
  NAND U22834 ( .A(n23988), .B(n22393), .Z(n22397) );
  NAND U22835 ( .A(n22395), .B(n22394), .Z(n22396) );
  NAND U22836 ( .A(n22397), .B(n22396), .Z(n22590) );
  XOR U22837 ( .A(n22591), .B(n22590), .Z(n22593) );
  AND U22838 ( .A(x[239]), .B(y[2027]), .Z(n23218) );
  NAND U22839 ( .A(n23218), .B(n22398), .Z(n22402) );
  NAND U22840 ( .A(n22400), .B(n22399), .Z(n22401) );
  NAND U22841 ( .A(n22402), .B(n22401), .Z(n22555) );
  AND U22842 ( .A(x[224]), .B(y[2037]), .Z(n22574) );
  AND U22843 ( .A(x[245]), .B(y[2016]), .Z(n22575) );
  XOR U22844 ( .A(n22574), .B(n22575), .Z(n22577) );
  AND U22845 ( .A(o[244]), .B(n22403), .Z(n22576) );
  XOR U22846 ( .A(n22577), .B(n22576), .Z(n22553) );
  AND U22847 ( .A(x[229]), .B(y[2032]), .Z(n22561) );
  AND U22848 ( .A(x[240]), .B(y[2021]), .Z(n22560) );
  XOR U22849 ( .A(n22561), .B(n22560), .Z(n22559) );
  AND U22850 ( .A(x[239]), .B(y[2022]), .Z(n22558) );
  XOR U22851 ( .A(n22559), .B(n22558), .Z(n22552) );
  XOR U22852 ( .A(n22553), .B(n22552), .Z(n22554) );
  XOR U22853 ( .A(n22555), .B(n22554), .Z(n22592) );
  XNOR U22854 ( .A(n22593), .B(n22592), .Z(n22608) );
  XOR U22855 ( .A(n22609), .B(n22608), .Z(n22610) );
  NAND U22856 ( .A(n22405), .B(n22404), .Z(n22409) );
  NAND U22857 ( .A(n22407), .B(n22406), .Z(n22408) );
  AND U22858 ( .A(n22409), .B(n22408), .Z(n22611) );
  XOR U22859 ( .A(n22610), .B(n22611), .Z(n22506) );
  NANDN U22860 ( .A(n22411), .B(n22410), .Z(n22415) );
  NAND U22861 ( .A(n22413), .B(n22412), .Z(n22414) );
  AND U22862 ( .A(n22415), .B(n22414), .Z(n22505) );
  XNOR U22863 ( .A(n22507), .B(n22508), .Z(n22501) );
  NAND U22864 ( .A(n22417), .B(n22416), .Z(n22421) );
  NAND U22865 ( .A(n22419), .B(n22418), .Z(n22420) );
  NAND U22866 ( .A(n22421), .B(n22420), .Z(n22514) );
  NAND U22867 ( .A(n23221), .B(n22422), .Z(n22426) );
  NAND U22868 ( .A(n22424), .B(n22423), .Z(n22425) );
  NAND U22869 ( .A(n22426), .B(n22425), .Z(n22524) );
  NAND U22870 ( .A(n23850), .B(n22427), .Z(n22431) );
  NAND U22871 ( .A(n22429), .B(n22428), .Z(n22430) );
  NAND U22872 ( .A(n22431), .B(n22430), .Z(n22605) );
  AND U22873 ( .A(y[2018]), .B(x[243]), .Z(n22433) );
  NAND U22874 ( .A(y[2026]), .B(x[235]), .Z(n22432) );
  XNOR U22875 ( .A(n22433), .B(n22432), .Z(n22543) );
  AND U22876 ( .A(x[244]), .B(y[2017]), .Z(n22573) );
  XOR U22877 ( .A(o[245]), .B(n22573), .Z(n22542) );
  XOR U22878 ( .A(n22543), .B(n22542), .Z(n22603) );
  AND U22879 ( .A(y[2019]), .B(x[242]), .Z(n22435) );
  NAND U22880 ( .A(y[2027]), .B(x[234]), .Z(n22434) );
  XNOR U22881 ( .A(n22435), .B(n22434), .Z(n22581) );
  AND U22882 ( .A(x[225]), .B(y[2036]), .Z(n22582) );
  XOR U22883 ( .A(n22581), .B(n22582), .Z(n22602) );
  XOR U22884 ( .A(n22603), .B(n22602), .Z(n22604) );
  XOR U22885 ( .A(n22605), .B(n22604), .Z(n22523) );
  XOR U22886 ( .A(n22524), .B(n22523), .Z(n22526) );
  AND U22887 ( .A(x[231]), .B(y[2030]), .Z(n22782) );
  AND U22888 ( .A(y[2031]), .B(x[230]), .Z(n22437) );
  NAND U22889 ( .A(y[2023]), .B(x[238]), .Z(n22436) );
  XNOR U22890 ( .A(n22437), .B(n22436), .Z(n22585) );
  XNOR U22891 ( .A(n22782), .B(n22585), .Z(n22532) );
  NAND U22892 ( .A(x[233]), .B(y[2028]), .Z(n22530) );
  NAND U22893 ( .A(x[232]), .B(y[2029]), .Z(n22529) );
  XOR U22894 ( .A(n22530), .B(n22529), .Z(n22531) );
  XNOR U22895 ( .A(n22532), .B(n22531), .Z(n22548) );
  AND U22896 ( .A(y[2025]), .B(x[236]), .Z(n22439) );
  NAND U22897 ( .A(y[2020]), .B(x[241]), .Z(n22438) );
  XNOR U22898 ( .A(n22439), .B(n22438), .Z(n22535) );
  AND U22899 ( .A(x[226]), .B(y[2035]), .Z(n22536) );
  XOR U22900 ( .A(n22535), .B(n22536), .Z(n22547) );
  AND U22901 ( .A(y[2024]), .B(x[237]), .Z(n22441) );
  NAND U22902 ( .A(y[2034]), .B(x[227]), .Z(n22440) );
  XNOR U22903 ( .A(n22441), .B(n22440), .Z(n22569) );
  AND U22904 ( .A(x[228]), .B(y[2033]), .Z(n22570) );
  XOR U22905 ( .A(n22569), .B(n22570), .Z(n22546) );
  XOR U22906 ( .A(n22547), .B(n22546), .Z(n22549) );
  XOR U22907 ( .A(n22548), .B(n22549), .Z(n22599) );
  NAND U22908 ( .A(n22561), .B(n22442), .Z(n22446) );
  NAND U22909 ( .A(n22444), .B(n22443), .Z(n22445) );
  NAND U22910 ( .A(n22446), .B(n22445), .Z(n22597) );
  NAND U22911 ( .A(n22448), .B(n22447), .Z(n22452) );
  NAND U22912 ( .A(n22450), .B(n22449), .Z(n22451) );
  NAND U22913 ( .A(n22452), .B(n22451), .Z(n22596) );
  XOR U22914 ( .A(n22597), .B(n22596), .Z(n22598) );
  XOR U22915 ( .A(n22599), .B(n22598), .Z(n22525) );
  XOR U22916 ( .A(n22526), .B(n22525), .Z(n22512) );
  NAND U22917 ( .A(n22454), .B(n22453), .Z(n22458) );
  NAND U22918 ( .A(n22456), .B(n22455), .Z(n22457) );
  NAND U22919 ( .A(n22458), .B(n22457), .Z(n22519) );
  NAND U22920 ( .A(n22460), .B(n22459), .Z(n22464) );
  NAND U22921 ( .A(n22462), .B(n22461), .Z(n22463) );
  NAND U22922 ( .A(n22464), .B(n22463), .Z(n22518) );
  NAND U22923 ( .A(n22466), .B(n22465), .Z(n22470) );
  NAND U22924 ( .A(n22468), .B(n22467), .Z(n22469) );
  NAND U22925 ( .A(n22470), .B(n22469), .Z(n22517) );
  XOR U22926 ( .A(n22518), .B(n22517), .Z(n22520) );
  XOR U22927 ( .A(n22519), .B(n22520), .Z(n22511) );
  XOR U22928 ( .A(n22512), .B(n22511), .Z(n22513) );
  XOR U22929 ( .A(n22514), .B(n22513), .Z(n22500) );
  NAND U22930 ( .A(n22472), .B(n22471), .Z(n22476) );
  NANDN U22931 ( .A(n22474), .B(n22473), .Z(n22475) );
  NAND U22932 ( .A(n22476), .B(n22475), .Z(n22499) );
  XOR U22933 ( .A(n22501), .B(n22502), .Z(n22623) );
  NAND U22934 ( .A(n22478), .B(n22477), .Z(n22482) );
  NAND U22935 ( .A(n22480), .B(n22479), .Z(n22481) );
  NAND U22936 ( .A(n22482), .B(n22481), .Z(n22622) );
  NANDN U22937 ( .A(n22484), .B(n22483), .Z(n22488) );
  NAND U22938 ( .A(n22486), .B(n22485), .Z(n22487) );
  AND U22939 ( .A(n22488), .B(n22487), .Z(n22621) );
  XOR U22940 ( .A(n22622), .B(n22621), .Z(n22624) );
  XNOR U22941 ( .A(n22623), .B(n22624), .Z(n22617) );
  NAND U22942 ( .A(n22493), .B(n22492), .Z(n22497) );
  NANDN U22943 ( .A(n22495), .B(n22494), .Z(n22496) );
  AND U22944 ( .A(n22497), .B(n22496), .Z(n22615) );
  IV U22945 ( .A(n22615), .Z(n22614) );
  XOR U22946 ( .A(n22616), .B(n22614), .Z(n22498) );
  XNOR U22947 ( .A(n22617), .B(n22498), .Z(N502) );
  NANDN U22948 ( .A(n22500), .B(n22499), .Z(n22504) );
  NANDN U22949 ( .A(n22502), .B(n22501), .Z(n22503) );
  AND U22950 ( .A(n22504), .B(n22503), .Z(n22757) );
  NANDN U22951 ( .A(n22506), .B(n22505), .Z(n22510) );
  NAND U22952 ( .A(n22508), .B(n22507), .Z(n22509) );
  NAND U22953 ( .A(n22510), .B(n22509), .Z(n22755) );
  NAND U22954 ( .A(n22512), .B(n22511), .Z(n22516) );
  NAND U22955 ( .A(n22514), .B(n22513), .Z(n22515) );
  NAND U22956 ( .A(n22516), .B(n22515), .Z(n22629) );
  NAND U22957 ( .A(n22518), .B(n22517), .Z(n22522) );
  NAND U22958 ( .A(n22520), .B(n22519), .Z(n22521) );
  NAND U22959 ( .A(n22522), .B(n22521), .Z(n22628) );
  XOR U22960 ( .A(n22629), .B(n22628), .Z(n22631) );
  NAND U22961 ( .A(n22524), .B(n22523), .Z(n22528) );
  NAND U22962 ( .A(n22526), .B(n22525), .Z(n22527) );
  AND U22963 ( .A(n22528), .B(n22527), .Z(n22745) );
  NAND U22964 ( .A(n22530), .B(n22529), .Z(n22534) );
  NAND U22965 ( .A(n22532), .B(n22531), .Z(n22533) );
  NAND U22966 ( .A(n22534), .B(n22533), .Z(n22739) );
  NANDN U22967 ( .A(n23229), .B(n22690), .Z(n22538) );
  NAND U22968 ( .A(n22536), .B(n22535), .Z(n22537) );
  NAND U22969 ( .A(n22538), .B(n22537), .Z(n22666) );
  AND U22970 ( .A(x[229]), .B(y[2033]), .Z(n22712) );
  AND U22971 ( .A(x[241]), .B(y[2021]), .Z(n22713) );
  XOR U22972 ( .A(n22712), .B(n22713), .Z(n22714) );
  AND U22973 ( .A(x[240]), .B(y[2022]), .Z(n22715) );
  XOR U22974 ( .A(n22714), .B(n22715), .Z(n22665) );
  AND U22975 ( .A(y[2020]), .B(x[242]), .Z(n22540) );
  NAND U22976 ( .A(y[2026]), .B(x[236]), .Z(n22539) );
  XNOR U22977 ( .A(n22540), .B(n22539), .Z(n22691) );
  AND U22978 ( .A(x[228]), .B(y[2034]), .Z(n22692) );
  XOR U22979 ( .A(n22691), .B(n22692), .Z(n22664) );
  XOR U22980 ( .A(n22665), .B(n22664), .Z(n22667) );
  XNOR U22981 ( .A(n22666), .B(n22667), .Z(n22736) );
  AND U22982 ( .A(x[243]), .B(y[2026]), .Z(n23741) );
  NAND U22983 ( .A(n23741), .B(n22541), .Z(n22545) );
  NAND U22984 ( .A(n22543), .B(n22542), .Z(n22544) );
  AND U22985 ( .A(n22545), .B(n22544), .Z(n22737) );
  XOR U22986 ( .A(n22736), .B(n22737), .Z(n22738) );
  XNOR U22987 ( .A(n22739), .B(n22738), .Z(n22742) );
  NAND U22988 ( .A(n22547), .B(n22546), .Z(n22551) );
  NAND U22989 ( .A(n22549), .B(n22548), .Z(n22550) );
  NAND U22990 ( .A(n22551), .B(n22550), .Z(n22725) );
  NAND U22991 ( .A(n22553), .B(n22552), .Z(n22557) );
  NAND U22992 ( .A(n22555), .B(n22554), .Z(n22556) );
  NAND U22993 ( .A(n22557), .B(n22556), .Z(n22724) );
  XOR U22994 ( .A(n22725), .B(n22724), .Z(n22727) );
  AND U22995 ( .A(n22559), .B(n22558), .Z(n22563) );
  NAND U22996 ( .A(n22561), .B(n22560), .Z(n22562) );
  NANDN U22997 ( .A(n22563), .B(n22562), .Z(n22687) );
  AND U22998 ( .A(y[2025]), .B(x[237]), .Z(n22565) );
  NAND U22999 ( .A(y[2018]), .B(x[244]), .Z(n22564) );
  XNOR U23000 ( .A(n22565), .B(n22564), .Z(n22708) );
  AND U23001 ( .A(x[226]), .B(y[2036]), .Z(n22709) );
  XOR U23002 ( .A(n22708), .B(n22709), .Z(n22685) );
  AND U23003 ( .A(y[2032]), .B(x[230]), .Z(n22567) );
  NAND U23004 ( .A(y[2023]), .B(x[239]), .Z(n22566) );
  XNOR U23005 ( .A(n22567), .B(n22566), .Z(n22720) );
  XOR U23006 ( .A(n22685), .B(n22684), .Z(n22686) );
  XOR U23007 ( .A(n22687), .B(n22686), .Z(n22731) );
  AND U23008 ( .A(x[237]), .B(y[2034]), .Z(n24032) );
  NAND U23009 ( .A(n22568), .B(n24032), .Z(n22572) );
  NAND U23010 ( .A(n22570), .B(n22569), .Z(n22571) );
  NAND U23011 ( .A(n22572), .B(n22571), .Z(n22655) );
  AND U23012 ( .A(x[225]), .B(y[2037]), .Z(n22678) );
  XOR U23013 ( .A(n22679), .B(n22678), .Z(n22677) );
  AND U23014 ( .A(o[245]), .B(n22573), .Z(n22676) );
  XOR U23015 ( .A(n22677), .B(n22676), .Z(n22653) );
  AND U23016 ( .A(x[238]), .B(y[2024]), .Z(n22670) );
  AND U23017 ( .A(x[227]), .B(y[2035]), .Z(n22671) );
  XOR U23018 ( .A(n22670), .B(n22671), .Z(n22672) );
  AND U23019 ( .A(x[243]), .B(y[2019]), .Z(n22673) );
  XOR U23020 ( .A(n22672), .B(n22673), .Z(n22652) );
  XOR U23021 ( .A(n22653), .B(n22652), .Z(n22654) );
  XOR U23022 ( .A(n22655), .B(n22654), .Z(n22730) );
  XOR U23023 ( .A(n22731), .B(n22730), .Z(n22733) );
  NAND U23024 ( .A(n22575), .B(n22574), .Z(n22579) );
  NAND U23025 ( .A(n22577), .B(n22576), .Z(n22578) );
  NAND U23026 ( .A(n22579), .B(n22578), .Z(n22647) );
  AND U23027 ( .A(x[242]), .B(y[2027]), .Z(n23744) );
  NAND U23028 ( .A(n23744), .B(n22580), .Z(n22584) );
  NAND U23029 ( .A(n22582), .B(n22581), .Z(n22583) );
  NAND U23030 ( .A(n22584), .B(n22583), .Z(n22646) );
  XOR U23031 ( .A(n22647), .B(n22646), .Z(n22649) );
  AND U23032 ( .A(x[238]), .B(y[2031]), .Z(n23754) );
  NAND U23033 ( .A(n23754), .B(n22719), .Z(n22587) );
  NAND U23034 ( .A(n22782), .B(n22585), .Z(n22586) );
  NAND U23035 ( .A(n22587), .B(n22586), .Z(n22661) );
  AND U23036 ( .A(x[224]), .B(y[2038]), .Z(n22695) );
  AND U23037 ( .A(x[246]), .B(y[2016]), .Z(n22696) );
  XOR U23038 ( .A(n22695), .B(n22696), .Z(n22698) );
  AND U23039 ( .A(x[245]), .B(y[2017]), .Z(n22718) );
  XOR U23040 ( .A(o[246]), .B(n22718), .Z(n22697) );
  XOR U23041 ( .A(n22698), .B(n22697), .Z(n22659) );
  AND U23042 ( .A(y[2031]), .B(x[231]), .Z(n22589) );
  NAND U23043 ( .A(y[2030]), .B(x[232]), .Z(n22588) );
  XNOR U23044 ( .A(n22589), .B(n22588), .Z(n22701) );
  XOR U23045 ( .A(n22659), .B(n22658), .Z(n22660) );
  XOR U23046 ( .A(n22661), .B(n22660), .Z(n22648) );
  XOR U23047 ( .A(n22649), .B(n22648), .Z(n22732) );
  XOR U23048 ( .A(n22733), .B(n22732), .Z(n22726) );
  XOR U23049 ( .A(n22727), .B(n22726), .Z(n22743) );
  XOR U23050 ( .A(n22742), .B(n22743), .Z(n22744) );
  NAND U23051 ( .A(n22591), .B(n22590), .Z(n22595) );
  NAND U23052 ( .A(n22593), .B(n22592), .Z(n22594) );
  NAND U23053 ( .A(n22595), .B(n22594), .Z(n22643) );
  NAND U23054 ( .A(n22597), .B(n22596), .Z(n22601) );
  NAND U23055 ( .A(n22599), .B(n22598), .Z(n22600) );
  NAND U23056 ( .A(n22601), .B(n22600), .Z(n22641) );
  NAND U23057 ( .A(n22603), .B(n22602), .Z(n22607) );
  NAND U23058 ( .A(n22605), .B(n22604), .Z(n22606) );
  NAND U23059 ( .A(n22607), .B(n22606), .Z(n22640) );
  XOR U23060 ( .A(n22641), .B(n22640), .Z(n22642) );
  XOR U23061 ( .A(n22643), .B(n22642), .Z(n22634) );
  NAND U23062 ( .A(n22609), .B(n22608), .Z(n22613) );
  NAND U23063 ( .A(n22611), .B(n22610), .Z(n22612) );
  AND U23064 ( .A(n22613), .B(n22612), .Z(n22635) );
  XOR U23065 ( .A(n22634), .B(n22635), .Z(n22636) );
  XOR U23066 ( .A(n22637), .B(n22636), .Z(n22630) );
  XOR U23067 ( .A(n22631), .B(n22630), .Z(n22756) );
  XNOR U23068 ( .A(n22755), .B(n22756), .Z(n22758) );
  OR U23069 ( .A(n22616), .B(n22614), .Z(n22620) );
  ANDN U23070 ( .B(n22616), .A(n22615), .Z(n22618) );
  OR U23071 ( .A(n22618), .B(n22617), .Z(n22619) );
  AND U23072 ( .A(n22620), .B(n22619), .Z(n22749) );
  NAND U23073 ( .A(n22622), .B(n22621), .Z(n22626) );
  NAND U23074 ( .A(n22624), .B(n22623), .Z(n22625) );
  AND U23075 ( .A(n22626), .B(n22625), .Z(n22750) );
  IV U23076 ( .A(n22750), .Z(n22748) );
  XOR U23077 ( .A(n22749), .B(n22748), .Z(n22627) );
  XNOR U23078 ( .A(n22751), .B(n22627), .Z(N503) );
  NAND U23079 ( .A(n22629), .B(n22628), .Z(n22633) );
  NAND U23080 ( .A(n22631), .B(n22630), .Z(n22632) );
  AND U23081 ( .A(n22633), .B(n22632), .Z(n22899) );
  NAND U23082 ( .A(n22635), .B(n22634), .Z(n22639) );
  NAND U23083 ( .A(n22637), .B(n22636), .Z(n22638) );
  AND U23084 ( .A(n22639), .B(n22638), .Z(n22897) );
  NAND U23085 ( .A(n22641), .B(n22640), .Z(n22645) );
  NAND U23086 ( .A(n22643), .B(n22642), .Z(n22644) );
  NAND U23087 ( .A(n22645), .B(n22644), .Z(n22878) );
  NAND U23088 ( .A(n22647), .B(n22646), .Z(n22651) );
  NAND U23089 ( .A(n22649), .B(n22648), .Z(n22650) );
  NAND U23090 ( .A(n22651), .B(n22650), .Z(n22872) );
  NAND U23091 ( .A(n22653), .B(n22652), .Z(n22657) );
  NAND U23092 ( .A(n22655), .B(n22654), .Z(n22656) );
  NAND U23093 ( .A(n22657), .B(n22656), .Z(n22870) );
  NAND U23094 ( .A(n22659), .B(n22658), .Z(n22663) );
  NAND U23095 ( .A(n22661), .B(n22660), .Z(n22662) );
  NAND U23096 ( .A(n22663), .B(n22662), .Z(n22869) );
  XOR U23097 ( .A(n22870), .B(n22869), .Z(n22871) );
  XOR U23098 ( .A(n22872), .B(n22871), .Z(n22890) );
  NAND U23099 ( .A(n22665), .B(n22664), .Z(n22669) );
  NAND U23100 ( .A(n22667), .B(n22666), .Z(n22668) );
  NAND U23101 ( .A(n22669), .B(n22668), .Z(n22888) );
  NAND U23102 ( .A(n22671), .B(n22670), .Z(n22675) );
  NAND U23103 ( .A(n22673), .B(n22672), .Z(n22674) );
  NAND U23104 ( .A(n22675), .B(n22674), .Z(n22816) );
  AND U23105 ( .A(n22677), .B(n22676), .Z(n22681) );
  NAND U23106 ( .A(n22679), .B(n22678), .Z(n22680) );
  NANDN U23107 ( .A(n22681), .B(n22680), .Z(n22815) );
  XOR U23108 ( .A(n22816), .B(n22815), .Z(n22818) );
  AND U23109 ( .A(y[2032]), .B(x[231]), .Z(n22683) );
  NAND U23110 ( .A(y[2030]), .B(x[233]), .Z(n22682) );
  XNOR U23111 ( .A(n22683), .B(n22682), .Z(n22783) );
  AND U23112 ( .A(x[234]), .B(y[2029]), .Z(n22822) );
  XOR U23113 ( .A(n22821), .B(n22822), .Z(n22824) );
  AND U23114 ( .A(x[230]), .B(y[2033]), .Z(n22774) );
  AND U23115 ( .A(x[239]), .B(y[2024]), .Z(n22775) );
  XOR U23116 ( .A(n22774), .B(n22775), .Z(n22776) );
  AND U23117 ( .A(x[235]), .B(y[2028]), .Z(n22777) );
  XOR U23118 ( .A(n22776), .B(n22777), .Z(n22823) );
  XOR U23119 ( .A(n22824), .B(n22823), .Z(n22817) );
  XOR U23120 ( .A(n22818), .B(n22817), .Z(n22887) );
  XOR U23121 ( .A(n22888), .B(n22887), .Z(n22889) );
  XOR U23122 ( .A(n22890), .B(n22889), .Z(n22876) );
  NAND U23123 ( .A(n22685), .B(n22684), .Z(n22689) );
  NAND U23124 ( .A(n22687), .B(n22686), .Z(n22688) );
  NAND U23125 ( .A(n22689), .B(n22688), .Z(n22810) );
  NAND U23126 ( .A(x[242]), .B(y[2026]), .Z(n23584) );
  NANDN U23127 ( .A(n23584), .B(n22690), .Z(n22694) );
  NAND U23128 ( .A(n22692), .B(n22691), .Z(n22693) );
  AND U23129 ( .A(n22694), .B(n22693), .Z(n22858) );
  NAND U23130 ( .A(n22696), .B(n22695), .Z(n22700) );
  NAND U23131 ( .A(n22698), .B(n22697), .Z(n22699) );
  NAND U23132 ( .A(n22700), .B(n22699), .Z(n22857) );
  NANDN U23133 ( .A(n22784), .B(n22782), .Z(n22704) );
  NANDN U23134 ( .A(n22702), .B(n22701), .Z(n22703) );
  AND U23135 ( .A(n22704), .B(n22703), .Z(n22854) );
  AND U23136 ( .A(x[224]), .B(y[2039]), .Z(n22793) );
  AND U23137 ( .A(x[247]), .B(y[2016]), .Z(n22794) );
  XOR U23138 ( .A(n22793), .B(n22794), .Z(n22796) );
  AND U23139 ( .A(x[246]), .B(y[2017]), .Z(n22773) );
  XOR U23140 ( .A(o[247]), .B(n22773), .Z(n22795) );
  XOR U23141 ( .A(n22796), .B(n22795), .Z(n22852) );
  NAND U23142 ( .A(y[2019]), .B(x[244]), .Z(n22705) );
  XNOR U23143 ( .A(n22706), .B(n22705), .Z(n22769) );
  AND U23144 ( .A(x[243]), .B(y[2020]), .Z(n22770) );
  XOR U23145 ( .A(n22769), .B(n22770), .Z(n22851) );
  XOR U23146 ( .A(n22852), .B(n22851), .Z(n22853) );
  XOR U23147 ( .A(n22860), .B(n22859), .Z(n22809) );
  XOR U23148 ( .A(n22810), .B(n22809), .Z(n22812) );
  NAND U23149 ( .A(x[244]), .B(y[2025]), .Z(n23766) );
  AND U23150 ( .A(x[237]), .B(y[2018]), .Z(n22707) );
  NANDN U23151 ( .A(n23766), .B(n22707), .Z(n22711) );
  NAND U23152 ( .A(n22709), .B(n22708), .Z(n22710) );
  NAND U23153 ( .A(n22711), .B(n22710), .Z(n22804) );
  NAND U23154 ( .A(n22713), .B(n22712), .Z(n22717) );
  NAND U23155 ( .A(n22715), .B(n22714), .Z(n22716) );
  AND U23156 ( .A(n22717), .B(n22716), .Z(n22866) );
  AND U23157 ( .A(x[237]), .B(y[2026]), .Z(n22839) );
  AND U23158 ( .A(x[226]), .B(y[2037]), .Z(n22840) );
  XOR U23159 ( .A(n22839), .B(n22840), .Z(n22841) );
  AND U23160 ( .A(x[245]), .B(y[2018]), .Z(n22842) );
  XOR U23161 ( .A(n22841), .B(n22842), .Z(n22864) );
  AND U23162 ( .A(x[236]), .B(y[2027]), .Z(n22787) );
  AND U23163 ( .A(x[225]), .B(y[2038]), .Z(n22788) );
  XOR U23164 ( .A(n22787), .B(n22788), .Z(n22790) );
  AND U23165 ( .A(o[246]), .B(n22718), .Z(n22789) );
  XOR U23166 ( .A(n22790), .B(n22789), .Z(n22863) );
  XOR U23167 ( .A(n22864), .B(n22863), .Z(n22865) );
  XOR U23168 ( .A(n22804), .B(n22803), .Z(n22806) );
  AND U23169 ( .A(x[239]), .B(y[2032]), .Z(n24020) );
  NAND U23170 ( .A(n24020), .B(n22719), .Z(n22723) );
  NANDN U23171 ( .A(n22721), .B(n22720), .Z(n22722) );
  AND U23172 ( .A(n22723), .B(n22722), .Z(n22848) );
  AND U23173 ( .A(x[238]), .B(y[2025]), .Z(n22833) );
  AND U23174 ( .A(x[227]), .B(y[2036]), .Z(n22834) );
  XOR U23175 ( .A(n22833), .B(n22834), .Z(n22835) );
  AND U23176 ( .A(x[228]), .B(y[2035]), .Z(n22836) );
  XOR U23177 ( .A(n22835), .B(n22836), .Z(n22846) );
  AND U23178 ( .A(x[229]), .B(y[2034]), .Z(n22827) );
  AND U23179 ( .A(x[242]), .B(y[2021]), .Z(n22828) );
  XOR U23180 ( .A(n22827), .B(n22828), .Z(n22829) );
  AND U23181 ( .A(x[241]), .B(y[2022]), .Z(n22830) );
  XOR U23182 ( .A(n22829), .B(n22830), .Z(n22845) );
  XOR U23183 ( .A(n22846), .B(n22845), .Z(n22847) );
  XOR U23184 ( .A(n22806), .B(n22805), .Z(n22811) );
  XOR U23185 ( .A(n22812), .B(n22811), .Z(n22875) );
  XOR U23186 ( .A(n22876), .B(n22875), .Z(n22877) );
  XNOR U23187 ( .A(n22878), .B(n22877), .Z(n22764) );
  NAND U23188 ( .A(n22725), .B(n22724), .Z(n22729) );
  NAND U23189 ( .A(n22727), .B(n22726), .Z(n22728) );
  NAND U23190 ( .A(n22729), .B(n22728), .Z(n22884) );
  NAND U23191 ( .A(n22731), .B(n22730), .Z(n22735) );
  NAND U23192 ( .A(n22733), .B(n22732), .Z(n22734) );
  NAND U23193 ( .A(n22735), .B(n22734), .Z(n22882) );
  NAND U23194 ( .A(n22737), .B(n22736), .Z(n22741) );
  NAND U23195 ( .A(n22739), .B(n22738), .Z(n22740) );
  AND U23196 ( .A(n22741), .B(n22740), .Z(n22881) );
  XOR U23197 ( .A(n22882), .B(n22881), .Z(n22883) );
  XNOR U23198 ( .A(n22884), .B(n22883), .Z(n22762) );
  NAND U23199 ( .A(n22743), .B(n22742), .Z(n22747) );
  NANDN U23200 ( .A(n22745), .B(n22744), .Z(n22746) );
  AND U23201 ( .A(n22747), .B(n22746), .Z(n22763) );
  XOR U23202 ( .A(n22762), .B(n22763), .Z(n22765) );
  XOR U23203 ( .A(n22764), .B(n22765), .Z(n22896) );
  XOR U23204 ( .A(n22897), .B(n22896), .Z(n22898) );
  XNOR U23205 ( .A(n22899), .B(n22898), .Z(n22895) );
  NANDN U23206 ( .A(n22748), .B(n22749), .Z(n22754) );
  NOR U23207 ( .A(n22750), .B(n22749), .Z(n22752) );
  OR U23208 ( .A(n22752), .B(n22751), .Z(n22753) );
  AND U23209 ( .A(n22754), .B(n22753), .Z(n22894) );
  NAND U23210 ( .A(n22756), .B(n22755), .Z(n22760) );
  NANDN U23211 ( .A(n22758), .B(n22757), .Z(n22759) );
  AND U23212 ( .A(n22760), .B(n22759), .Z(n22893) );
  XOR U23213 ( .A(n22894), .B(n22893), .Z(n22761) );
  XNOR U23214 ( .A(n22895), .B(n22761), .Z(N504) );
  NAND U23215 ( .A(n22763), .B(n22762), .Z(n22767) );
  NAND U23216 ( .A(n22765), .B(n22764), .Z(n22766) );
  AND U23217 ( .A(n22767), .B(n22766), .Z(n23040) );
  AND U23218 ( .A(x[244]), .B(y[2023]), .Z(n22768) );
  NAND U23219 ( .A(n22768), .B(n22999), .Z(n22772) );
  NAND U23220 ( .A(n22770), .B(n22769), .Z(n22771) );
  NAND U23221 ( .A(n22772), .B(n22771), .Z(n23019) );
  AND U23222 ( .A(x[246]), .B(y[2018]), .Z(n22927) );
  XOR U23223 ( .A(n22928), .B(n22927), .Z(n22926) );
  AND U23224 ( .A(x[226]), .B(y[2038]), .Z(n22925) );
  XOR U23225 ( .A(n22926), .B(n22925), .Z(n23017) );
  AND U23226 ( .A(x[225]), .B(y[2039]), .Z(n22933) );
  XOR U23227 ( .A(n22934), .B(n22933), .Z(n22932) );
  AND U23228 ( .A(o[247]), .B(n22773), .Z(n22931) );
  XOR U23229 ( .A(n22932), .B(n22931), .Z(n23016) );
  XOR U23230 ( .A(n23017), .B(n23016), .Z(n23018) );
  XOR U23231 ( .A(n23019), .B(n23018), .Z(n22964) );
  NAND U23232 ( .A(n22775), .B(n22774), .Z(n22779) );
  NAND U23233 ( .A(n22777), .B(n22776), .Z(n22778) );
  NAND U23234 ( .A(n22779), .B(n22778), .Z(n23013) );
  AND U23235 ( .A(y[2024]), .B(x[240]), .Z(n22781) );
  NAND U23236 ( .A(y[2019]), .B(x[245]), .Z(n22780) );
  XNOR U23237 ( .A(n22781), .B(n22780), .Z(n23000) );
  AND U23238 ( .A(x[229]), .B(y[2035]), .Z(n23001) );
  XOR U23239 ( .A(n23000), .B(n23001), .Z(n23011) );
  AND U23240 ( .A(x[230]), .B(y[2034]), .Z(n23318) );
  NAND U23241 ( .A(x[244]), .B(y[2020]), .Z(n23156) );
  AND U23242 ( .A(x[243]), .B(y[2021]), .Z(n23007) );
  XOR U23243 ( .A(n23006), .B(n23007), .Z(n23010) );
  XOR U23244 ( .A(n23011), .B(n23010), .Z(n23012) );
  XOR U23245 ( .A(n23013), .B(n23012), .Z(n22990) );
  NAND U23246 ( .A(n23081), .B(n22782), .Z(n22786) );
  NANDN U23247 ( .A(n22784), .B(n22783), .Z(n22785) );
  NAND U23248 ( .A(n22786), .B(n22785), .Z(n22988) );
  NAND U23249 ( .A(n22788), .B(n22787), .Z(n22792) );
  NAND U23250 ( .A(n22790), .B(n22789), .Z(n22791) );
  NAND U23251 ( .A(n22792), .B(n22791), .Z(n22987) );
  XOR U23252 ( .A(n22988), .B(n22987), .Z(n22989) );
  XOR U23253 ( .A(n22990), .B(n22989), .Z(n22963) );
  XOR U23254 ( .A(n22964), .B(n22963), .Z(n22966) );
  NAND U23255 ( .A(n22794), .B(n22793), .Z(n22798) );
  NAND U23256 ( .A(n22796), .B(n22795), .Z(n22797) );
  NAND U23257 ( .A(n22798), .B(n22797), .Z(n22958) );
  AND U23258 ( .A(x[227]), .B(y[2037]), .Z(n22947) );
  XOR U23259 ( .A(n22948), .B(n22947), .Z(n22946) );
  AND U23260 ( .A(x[228]), .B(y[2036]), .Z(n22945) );
  XOR U23261 ( .A(n22946), .B(n22945), .Z(n22957) );
  XOR U23262 ( .A(n22958), .B(n22957), .Z(n22960) );
  AND U23263 ( .A(y[2031]), .B(x[233]), .Z(n22800) );
  NAND U23264 ( .A(y[2030]), .B(x[234]), .Z(n22799) );
  XNOR U23265 ( .A(n22800), .B(n22799), .Z(n22917) );
  AND U23266 ( .A(y[2026]), .B(x[238]), .Z(n22802) );
  NAND U23267 ( .A(y[2032]), .B(x[232]), .Z(n22801) );
  XNOR U23268 ( .A(n22802), .B(n22801), .Z(n22921) );
  NAND U23269 ( .A(x[235]), .B(y[2029]), .Z(n22922) );
  XOR U23270 ( .A(n22917), .B(n22916), .Z(n22959) );
  XOR U23271 ( .A(n22960), .B(n22959), .Z(n22965) );
  XNOR U23272 ( .A(n22966), .B(n22965), .Z(n22910) );
  NAND U23273 ( .A(n22804), .B(n22803), .Z(n22808) );
  NAND U23274 ( .A(n22806), .B(n22805), .Z(n22807) );
  AND U23275 ( .A(n22808), .B(n22807), .Z(n22909) );
  XOR U23276 ( .A(n22910), .B(n22909), .Z(n22912) );
  NAND U23277 ( .A(n22810), .B(n22809), .Z(n22814) );
  NAND U23278 ( .A(n22812), .B(n22811), .Z(n22813) );
  AND U23279 ( .A(n22814), .B(n22813), .Z(n22911) );
  XOR U23280 ( .A(n22912), .B(n22911), .Z(n23031) );
  NAND U23281 ( .A(n22816), .B(n22815), .Z(n22820) );
  NAND U23282 ( .A(n22818), .B(n22817), .Z(n22819) );
  NAND U23283 ( .A(n22820), .B(n22819), .Z(n22972) );
  NAND U23284 ( .A(n22822), .B(n22821), .Z(n22826) );
  NAND U23285 ( .A(n22824), .B(n22823), .Z(n22825) );
  NAND U23286 ( .A(n22826), .B(n22825), .Z(n22970) );
  NAND U23287 ( .A(n22828), .B(n22827), .Z(n22832) );
  NAND U23288 ( .A(n22830), .B(n22829), .Z(n22831) );
  NAND U23289 ( .A(n22832), .B(n22831), .Z(n22996) );
  AND U23290 ( .A(x[224]), .B(y[2040]), .Z(n22951) );
  AND U23291 ( .A(x[248]), .B(y[2016]), .Z(n22952) );
  XOR U23292 ( .A(n22951), .B(n22952), .Z(n22953) );
  NAND U23293 ( .A(x[247]), .B(y[2017]), .Z(n22944) );
  XNOR U23294 ( .A(o[248]), .B(n22944), .Z(n22954) );
  XOR U23295 ( .A(n22953), .B(n22954), .Z(n22994) );
  AND U23296 ( .A(x[231]), .B(y[2033]), .Z(n22937) );
  AND U23297 ( .A(x[242]), .B(y[2022]), .Z(n22938) );
  XOR U23298 ( .A(n22937), .B(n22938), .Z(n22939) );
  AND U23299 ( .A(x[241]), .B(y[2023]), .Z(n22940) );
  XOR U23300 ( .A(n22939), .B(n22940), .Z(n22993) );
  XOR U23301 ( .A(n22994), .B(n22993), .Z(n22995) );
  XOR U23302 ( .A(n22996), .B(n22995), .Z(n22984) );
  NAND U23303 ( .A(n22834), .B(n22833), .Z(n22838) );
  NAND U23304 ( .A(n22836), .B(n22835), .Z(n22837) );
  NAND U23305 ( .A(n22838), .B(n22837), .Z(n22982) );
  NAND U23306 ( .A(n22840), .B(n22839), .Z(n22844) );
  NAND U23307 ( .A(n22842), .B(n22841), .Z(n22843) );
  NAND U23308 ( .A(n22844), .B(n22843), .Z(n22981) );
  XOR U23309 ( .A(n22982), .B(n22981), .Z(n22983) );
  XOR U23310 ( .A(n22984), .B(n22983), .Z(n22969) );
  XOR U23311 ( .A(n22970), .B(n22969), .Z(n22971) );
  XNOR U23312 ( .A(n22972), .B(n22971), .Z(n22978) );
  NAND U23313 ( .A(n22846), .B(n22845), .Z(n22850) );
  NANDN U23314 ( .A(n22848), .B(n22847), .Z(n22849) );
  AND U23315 ( .A(n22850), .B(n22849), .Z(n23023) );
  NAND U23316 ( .A(n22852), .B(n22851), .Z(n22856) );
  NANDN U23317 ( .A(n22854), .B(n22853), .Z(n22855) );
  AND U23318 ( .A(n22856), .B(n22855), .Z(n23022) );
  XOR U23319 ( .A(n23023), .B(n23022), .Z(n23025) );
  NANDN U23320 ( .A(n22858), .B(n22857), .Z(n22862) );
  NAND U23321 ( .A(n22860), .B(n22859), .Z(n22861) );
  AND U23322 ( .A(n22862), .B(n22861), .Z(n23024) );
  XOR U23323 ( .A(n23025), .B(n23024), .Z(n22976) );
  NAND U23324 ( .A(n22864), .B(n22863), .Z(n22868) );
  NANDN U23325 ( .A(n22866), .B(n22865), .Z(n22867) );
  AND U23326 ( .A(n22868), .B(n22867), .Z(n22975) );
  XOR U23327 ( .A(n22976), .B(n22975), .Z(n22977) );
  XOR U23328 ( .A(n22978), .B(n22977), .Z(n23028) );
  NAND U23329 ( .A(n22870), .B(n22869), .Z(n22874) );
  NAND U23330 ( .A(n22872), .B(n22871), .Z(n22873) );
  AND U23331 ( .A(n22874), .B(n22873), .Z(n23029) );
  XOR U23332 ( .A(n23028), .B(n23029), .Z(n23030) );
  XOR U23333 ( .A(n23031), .B(n23030), .Z(n23038) );
  NAND U23334 ( .A(n22876), .B(n22875), .Z(n22880) );
  NAND U23335 ( .A(n22878), .B(n22877), .Z(n22879) );
  NAND U23336 ( .A(n22880), .B(n22879), .Z(n22906) );
  NAND U23337 ( .A(n22882), .B(n22881), .Z(n22886) );
  NAND U23338 ( .A(n22884), .B(n22883), .Z(n22885) );
  NAND U23339 ( .A(n22886), .B(n22885), .Z(n22904) );
  NAND U23340 ( .A(n22888), .B(n22887), .Z(n22892) );
  NAND U23341 ( .A(n22890), .B(n22889), .Z(n22891) );
  NAND U23342 ( .A(n22892), .B(n22891), .Z(n22903) );
  XOR U23343 ( .A(n22904), .B(n22903), .Z(n22905) );
  XOR U23344 ( .A(n22906), .B(n22905), .Z(n23037) );
  XNOR U23345 ( .A(n23040), .B(n23039), .Z(n23036) );
  NAND U23346 ( .A(n22897), .B(n22896), .Z(n22901) );
  NAND U23347 ( .A(n22899), .B(n22898), .Z(n22900) );
  AND U23348 ( .A(n22901), .B(n22900), .Z(n23035) );
  XOR U23349 ( .A(n23034), .B(n23035), .Z(n22902) );
  XNOR U23350 ( .A(n23036), .B(n22902), .Z(N505) );
  NAND U23351 ( .A(n22904), .B(n22903), .Z(n22908) );
  NAND U23352 ( .A(n22906), .B(n22905), .Z(n22907) );
  AND U23353 ( .A(n22908), .B(n22907), .Z(n23195) );
  NAND U23354 ( .A(n22910), .B(n22909), .Z(n22914) );
  NAND U23355 ( .A(n22912), .B(n22911), .Z(n22913) );
  NAND U23356 ( .A(n22914), .B(n22913), .Z(n23044) );
  IV U23357 ( .A(n22943), .Z(n23080) );
  NANDN U23358 ( .A(n23080), .B(n22915), .Z(n22919) );
  NAND U23359 ( .A(n22917), .B(n22916), .Z(n22918) );
  NAND U23360 ( .A(n22919), .B(n22918), .Z(n23105) );
  AND U23361 ( .A(x[238]), .B(y[2032]), .Z(n23942) );
  NAND U23362 ( .A(n23942), .B(n22920), .Z(n22924) );
  NANDN U23363 ( .A(n22922), .B(n22921), .Z(n22923) );
  AND U23364 ( .A(n22924), .B(n22923), .Z(n23134) );
  AND U23365 ( .A(x[235]), .B(y[2030]), .Z(n23152) );
  AND U23366 ( .A(x[236]), .B(y[2029]), .Z(n23151) );
  NAND U23367 ( .A(x[231]), .B(y[2034]), .Z(n23150) );
  XOR U23368 ( .A(n23151), .B(n23150), .Z(n23153) );
  XOR U23369 ( .A(n23152), .B(n23153), .Z(n23132) );
  NAND U23370 ( .A(x[248]), .B(y[2017]), .Z(n23149) );
  XNOR U23371 ( .A(o[249]), .B(n23149), .Z(n23119) );
  NAND U23372 ( .A(x[225]), .B(y[2040]), .Z(n23120) );
  NAND U23373 ( .A(x[237]), .B(y[2028]), .Z(n23122) );
  XOR U23374 ( .A(n23105), .B(n23104), .Z(n23107) );
  AND U23375 ( .A(n22926), .B(n22925), .Z(n22930) );
  NAND U23376 ( .A(n22928), .B(n22927), .Z(n22929) );
  NANDN U23377 ( .A(n22930), .B(n22929), .Z(n23093) );
  AND U23378 ( .A(n22932), .B(n22931), .Z(n22936) );
  NAND U23379 ( .A(n22934), .B(n22933), .Z(n22935) );
  NANDN U23380 ( .A(n22936), .B(n22935), .Z(n23092) );
  XOR U23381 ( .A(n23093), .B(n23092), .Z(n23095) );
  NAND U23382 ( .A(n22938), .B(n22937), .Z(n22942) );
  NAND U23383 ( .A(n22940), .B(n22939), .Z(n22941) );
  NAND U23384 ( .A(n22942), .B(n22941), .Z(n23089) );
  AND U23385 ( .A(x[232]), .B(y[2033]), .Z(n23083) );
  XOR U23386 ( .A(n23081), .B(n22943), .Z(n23082) );
  XOR U23387 ( .A(n23083), .B(n23082), .Z(n23087) );
  ANDN U23388 ( .B(o[248]), .A(n22944), .Z(n23076) );
  AND U23389 ( .A(x[249]), .B(y[2016]), .Z(n23075) );
  NAND U23390 ( .A(x[224]), .B(y[2041]), .Z(n23074) );
  XOR U23391 ( .A(n23075), .B(n23074), .Z(n23077) );
  XNOR U23392 ( .A(n23076), .B(n23077), .Z(n23086) );
  XOR U23393 ( .A(n23087), .B(n23086), .Z(n23088) );
  XOR U23394 ( .A(n23089), .B(n23088), .Z(n23094) );
  XOR U23395 ( .A(n23095), .B(n23094), .Z(n23106) );
  XNOR U23396 ( .A(n23107), .B(n23106), .Z(n23065) );
  AND U23397 ( .A(n22946), .B(n22945), .Z(n22950) );
  NAND U23398 ( .A(n22948), .B(n22947), .Z(n22949) );
  NANDN U23399 ( .A(n22950), .B(n22949), .Z(n23170) );
  NAND U23400 ( .A(n22952), .B(n22951), .Z(n22956) );
  NAND U23401 ( .A(n22954), .B(n22953), .Z(n22955) );
  NAND U23402 ( .A(n22956), .B(n22955), .Z(n23168) );
  AND U23403 ( .A(x[238]), .B(y[2027]), .Z(n23125) );
  NAND U23404 ( .A(x[226]), .B(y[2039]), .Z(n23126) );
  NAND U23405 ( .A(x[227]), .B(y[2038]), .Z(n23128) );
  XOR U23406 ( .A(n23168), .B(n23167), .Z(n23169) );
  XNOR U23407 ( .A(n23170), .B(n23169), .Z(n23063) );
  NAND U23408 ( .A(n22958), .B(n22957), .Z(n22962) );
  NAND U23409 ( .A(n22960), .B(n22959), .Z(n22961) );
  AND U23410 ( .A(n22962), .B(n22961), .Z(n23062) );
  XOR U23411 ( .A(n23063), .B(n23062), .Z(n23064) );
  XOR U23412 ( .A(n23065), .B(n23064), .Z(n23056) );
  NAND U23413 ( .A(n22964), .B(n22963), .Z(n22968) );
  NAND U23414 ( .A(n22966), .B(n22965), .Z(n22967) );
  AND U23415 ( .A(n22968), .B(n22967), .Z(n23057) );
  XOR U23416 ( .A(n23056), .B(n23057), .Z(n23058) );
  NAND U23417 ( .A(n22970), .B(n22969), .Z(n22974) );
  NAND U23418 ( .A(n22972), .B(n22971), .Z(n22973) );
  AND U23419 ( .A(n22974), .B(n22973), .Z(n23059) );
  XOR U23420 ( .A(n23058), .B(n23059), .Z(n23045) );
  XOR U23421 ( .A(n23044), .B(n23045), .Z(n23047) );
  NAND U23422 ( .A(n22976), .B(n22975), .Z(n22980) );
  NAND U23423 ( .A(n22978), .B(n22977), .Z(n22979) );
  NAND U23424 ( .A(n22980), .B(n22979), .Z(n23052) );
  NAND U23425 ( .A(n22982), .B(n22981), .Z(n22986) );
  NAND U23426 ( .A(n22984), .B(n22983), .Z(n22985) );
  NAND U23427 ( .A(n22986), .B(n22985), .Z(n23069) );
  NAND U23428 ( .A(n22988), .B(n22987), .Z(n22992) );
  NAND U23429 ( .A(n22990), .B(n22989), .Z(n22991) );
  NAND U23430 ( .A(n22992), .B(n22991), .Z(n23068) );
  XOR U23431 ( .A(n23069), .B(n23068), .Z(n23071) );
  NAND U23432 ( .A(n22994), .B(n22993), .Z(n22998) );
  NAND U23433 ( .A(n22996), .B(n22995), .Z(n22997) );
  AND U23434 ( .A(n22998), .B(n22997), .Z(n23101) );
  AND U23435 ( .A(x[245]), .B(y[2024]), .Z(n23917) );
  NAND U23436 ( .A(n23917), .B(n22999), .Z(n23003) );
  NAND U23437 ( .A(n23001), .B(n23000), .Z(n23002) );
  NAND U23438 ( .A(n23003), .B(n23002), .Z(n23176) );
  AND U23439 ( .A(x[246]), .B(y[2019]), .Z(n23145) );
  AND U23440 ( .A(x[229]), .B(y[2036]), .Z(n23144) );
  NAND U23441 ( .A(x[241]), .B(y[2024]), .Z(n23143) );
  XOR U23442 ( .A(n23144), .B(n23143), .Z(n23146) );
  XNOR U23443 ( .A(n23145), .B(n23146), .Z(n23174) );
  AND U23444 ( .A(y[2021]), .B(x[244]), .Z(n23005) );
  NAND U23445 ( .A(y[2020]), .B(x[245]), .Z(n23004) );
  XNOR U23446 ( .A(n23005), .B(n23004), .Z(n23157) );
  NAND U23447 ( .A(x[243]), .B(y[2022]), .Z(n23158) );
  XOR U23448 ( .A(n23174), .B(n23173), .Z(n23175) );
  XNOR U23449 ( .A(n23176), .B(n23175), .Z(n23099) );
  NANDN U23450 ( .A(n23156), .B(n23318), .Z(n23009) );
  NAND U23451 ( .A(n23007), .B(n23006), .Z(n23008) );
  AND U23452 ( .A(n23009), .B(n23008), .Z(n23182) );
  AND U23453 ( .A(x[239]), .B(y[2026]), .Z(n23163) );
  AND U23454 ( .A(x[242]), .B(y[2023]), .Z(n23162) );
  NAND U23455 ( .A(x[230]), .B(y[2035]), .Z(n23161) );
  XOR U23456 ( .A(n23162), .B(n23161), .Z(n23164) );
  XNOR U23457 ( .A(n23163), .B(n23164), .Z(n23180) );
  AND U23458 ( .A(x[247]), .B(y[2018]), .Z(n23139) );
  AND U23459 ( .A(x[228]), .B(y[2037]), .Z(n23138) );
  NAND U23460 ( .A(x[240]), .B(y[2025]), .Z(n23137) );
  XOR U23461 ( .A(n23138), .B(n23137), .Z(n23140) );
  XNOR U23462 ( .A(n23139), .B(n23140), .Z(n23179) );
  XOR U23463 ( .A(n23180), .B(n23179), .Z(n23181) );
  XOR U23464 ( .A(n23182), .B(n23181), .Z(n23098) );
  XOR U23465 ( .A(n23099), .B(n23098), .Z(n23100) );
  XNOR U23466 ( .A(n23101), .B(n23100), .Z(n23113) );
  NAND U23467 ( .A(n23011), .B(n23010), .Z(n23015) );
  NAND U23468 ( .A(n23013), .B(n23012), .Z(n23014) );
  NAND U23469 ( .A(n23015), .B(n23014), .Z(n23111) );
  NAND U23470 ( .A(n23017), .B(n23016), .Z(n23021) );
  NAND U23471 ( .A(n23019), .B(n23018), .Z(n23020) );
  NAND U23472 ( .A(n23021), .B(n23020), .Z(n23110) );
  XOR U23473 ( .A(n23111), .B(n23110), .Z(n23112) );
  XOR U23474 ( .A(n23113), .B(n23112), .Z(n23070) );
  XOR U23475 ( .A(n23071), .B(n23070), .Z(n23051) );
  NAND U23476 ( .A(n23023), .B(n23022), .Z(n23027) );
  NAND U23477 ( .A(n23025), .B(n23024), .Z(n23026) );
  NAND U23478 ( .A(n23027), .B(n23026), .Z(n23050) );
  XOR U23479 ( .A(n23052), .B(n23053), .Z(n23046) );
  XNOR U23480 ( .A(n23047), .B(n23046), .Z(n23193) );
  NAND U23481 ( .A(n23029), .B(n23028), .Z(n23033) );
  NAND U23482 ( .A(n23031), .B(n23030), .Z(n23032) );
  AND U23483 ( .A(n23033), .B(n23032), .Z(n23192) );
  XOR U23484 ( .A(n23193), .B(n23192), .Z(n23194) );
  XOR U23485 ( .A(n23195), .B(n23194), .Z(n23188) );
  NANDN U23486 ( .A(n23038), .B(n23037), .Z(n23042) );
  NAND U23487 ( .A(n23040), .B(n23039), .Z(n23041) );
  NAND U23488 ( .A(n23042), .B(n23041), .Z(n23186) );
  IV U23489 ( .A(n23186), .Z(n23185) );
  XOR U23490 ( .A(n23187), .B(n23185), .Z(n23043) );
  XNOR U23491 ( .A(n23188), .B(n23043), .Z(N506) );
  NAND U23492 ( .A(n23045), .B(n23044), .Z(n23049) );
  NAND U23493 ( .A(n23047), .B(n23046), .Z(n23048) );
  AND U23494 ( .A(n23049), .B(n23048), .Z(n23350) );
  NANDN U23495 ( .A(n23051), .B(n23050), .Z(n23055) );
  NAND U23496 ( .A(n23053), .B(n23052), .Z(n23054) );
  AND U23497 ( .A(n23055), .B(n23054), .Z(n23349) );
  XOR U23498 ( .A(n23350), .B(n23349), .Z(n23352) );
  NAND U23499 ( .A(n23057), .B(n23056), .Z(n23061) );
  NAND U23500 ( .A(n23059), .B(n23058), .Z(n23060) );
  AND U23501 ( .A(n23061), .B(n23060), .Z(n23199) );
  NAND U23502 ( .A(n23063), .B(n23062), .Z(n23067) );
  NAND U23503 ( .A(n23065), .B(n23064), .Z(n23066) );
  AND U23504 ( .A(n23067), .B(n23066), .Z(n23200) );
  XOR U23505 ( .A(n23199), .B(n23200), .Z(n23202) );
  NAND U23506 ( .A(n23069), .B(n23068), .Z(n23073) );
  NAND U23507 ( .A(n23071), .B(n23070), .Z(n23072) );
  NAND U23508 ( .A(n23073), .B(n23072), .Z(n23339) );
  AND U23509 ( .A(x[226]), .B(y[2040]), .Z(n23217) );
  XOR U23510 ( .A(n23218), .B(n23217), .Z(n23216) );
  AND U23511 ( .A(x[248]), .B(y[2018]), .Z(n23215) );
  XOR U23512 ( .A(n23216), .B(n23215), .Z(n23251) );
  NANDN U23513 ( .A(n23075), .B(n23074), .Z(n23079) );
  OR U23514 ( .A(n23077), .B(n23076), .Z(n23078) );
  NAND U23515 ( .A(n23079), .B(n23078), .Z(n23252) );
  XNOR U23516 ( .A(n23251), .B(n23252), .Z(n23254) );
  NANDN U23517 ( .A(n23081), .B(n23080), .Z(n23085) );
  NANDN U23518 ( .A(n23083), .B(n23082), .Z(n23084) );
  AND U23519 ( .A(n23085), .B(n23084), .Z(n23253) );
  XNOR U23520 ( .A(n23254), .B(n23253), .Z(n23290) );
  NAND U23521 ( .A(n23087), .B(n23086), .Z(n23091) );
  NAND U23522 ( .A(n23089), .B(n23088), .Z(n23090) );
  AND U23523 ( .A(n23091), .B(n23090), .Z(n23289) );
  XOR U23524 ( .A(n23290), .B(n23289), .Z(n23291) );
  NAND U23525 ( .A(n23093), .B(n23092), .Z(n23097) );
  NAND U23526 ( .A(n23095), .B(n23094), .Z(n23096) );
  AND U23527 ( .A(n23097), .B(n23096), .Z(n23292) );
  XOR U23528 ( .A(n23291), .B(n23292), .Z(n23333) );
  NAND U23529 ( .A(n23099), .B(n23098), .Z(n23103) );
  NAND U23530 ( .A(n23101), .B(n23100), .Z(n23102) );
  NAND U23531 ( .A(n23103), .B(n23102), .Z(n23330) );
  NAND U23532 ( .A(n23105), .B(n23104), .Z(n23109) );
  NAND U23533 ( .A(n23107), .B(n23106), .Z(n23108) );
  AND U23534 ( .A(n23109), .B(n23108), .Z(n23331) );
  XOR U23535 ( .A(n23330), .B(n23331), .Z(n23332) );
  XNOR U23536 ( .A(n23333), .B(n23332), .Z(n23337) );
  NAND U23537 ( .A(n23111), .B(n23110), .Z(n23115) );
  NAND U23538 ( .A(n23113), .B(n23112), .Z(n23114) );
  NAND U23539 ( .A(n23115), .B(n23114), .Z(n23285) );
  NAND U23540 ( .A(x[231]), .B(y[2035]), .Z(n23295) );
  AND U23541 ( .A(x[236]), .B(y[2030]), .Z(n23410) );
  AND U23542 ( .A(x[229]), .B(y[2037]), .Z(n23268) );
  XOR U23543 ( .A(n23410), .B(n23268), .Z(n23267) );
  AND U23544 ( .A(x[234]), .B(y[2032]), .Z(n23266) );
  XNOR U23545 ( .A(n23267), .B(n23266), .Z(n23297) );
  AND U23546 ( .A(y[2036]), .B(x[230]), .Z(n23117) );
  NAND U23547 ( .A(y[2034]), .B(x[232]), .Z(n23116) );
  XNOR U23548 ( .A(n23117), .B(n23116), .Z(n23320) );
  AND U23549 ( .A(x[233]), .B(y[2033]), .Z(n23319) );
  XNOR U23550 ( .A(n23320), .B(n23319), .Z(n23296) );
  XNOR U23551 ( .A(n23297), .B(n23296), .Z(n23118) );
  XOR U23552 ( .A(n23295), .B(n23118), .Z(n23242) );
  NANDN U23553 ( .A(n23120), .B(n23119), .Z(n23124) );
  NANDN U23554 ( .A(n23122), .B(n23121), .Z(n23123) );
  NAND U23555 ( .A(n23124), .B(n23123), .Z(n23240) );
  NANDN U23556 ( .A(n23126), .B(n23125), .Z(n23130) );
  NANDN U23557 ( .A(n23128), .B(n23127), .Z(n23129) );
  NAND U23558 ( .A(n23130), .B(n23129), .Z(n23239) );
  XOR U23559 ( .A(n23240), .B(n23239), .Z(n23241) );
  XNOR U23560 ( .A(n23242), .B(n23241), .Z(n23278) );
  NANDN U23561 ( .A(n23132), .B(n23131), .Z(n23136) );
  NANDN U23562 ( .A(n23134), .B(n23133), .Z(n23135) );
  AND U23563 ( .A(n23136), .B(n23135), .Z(n23277) );
  XOR U23564 ( .A(n23278), .B(n23277), .Z(n23280) );
  NANDN U23565 ( .A(n23138), .B(n23137), .Z(n23142) );
  OR U23566 ( .A(n23140), .B(n23139), .Z(n23141) );
  AND U23567 ( .A(n23142), .B(n23141), .Z(n23205) );
  NANDN U23568 ( .A(n23144), .B(n23143), .Z(n23148) );
  OR U23569 ( .A(n23146), .B(n23145), .Z(n23147) );
  NAND U23570 ( .A(n23148), .B(n23147), .Z(n23206) );
  XNOR U23571 ( .A(n23205), .B(n23206), .Z(n23208) );
  ANDN U23572 ( .B(o[249]), .A(n23149), .Z(n23312) );
  AND U23573 ( .A(x[238]), .B(y[2028]), .Z(n23313) );
  XOR U23574 ( .A(n23312), .B(n23313), .Z(n23314) );
  AND U23575 ( .A(x[225]), .B(y[2041]), .Z(n23315) );
  XOR U23576 ( .A(n23314), .B(n23315), .Z(n23257) );
  AND U23577 ( .A(x[249]), .B(y[2017]), .Z(n23323) );
  XOR U23578 ( .A(o[250]), .B(n23323), .Z(n23271) );
  NAND U23579 ( .A(x[250]), .B(y[2016]), .Z(n23272) );
  XNOR U23580 ( .A(n23271), .B(n23272), .Z(n23273) );
  NAND U23581 ( .A(x[224]), .B(y[2042]), .Z(n23274) );
  XOR U23582 ( .A(n23273), .B(n23274), .Z(n23258) );
  XNOR U23583 ( .A(n23257), .B(n23258), .Z(n23259) );
  NANDN U23584 ( .A(n23151), .B(n23150), .Z(n23155) );
  OR U23585 ( .A(n23153), .B(n23152), .Z(n23154) );
  NAND U23586 ( .A(n23155), .B(n23154), .Z(n23260) );
  XNOR U23587 ( .A(n23259), .B(n23260), .Z(n23207) );
  XNOR U23588 ( .A(n23208), .B(n23207), .Z(n23248) );
  AND U23589 ( .A(x[245]), .B(y[2021]), .Z(n23306) );
  NANDN U23590 ( .A(n23156), .B(n23306), .Z(n23160) );
  NANDN U23591 ( .A(n23158), .B(n23157), .Z(n23159) );
  NAND U23592 ( .A(n23160), .B(n23159), .Z(n23236) );
  XOR U23593 ( .A(n23307), .B(n23306), .Z(n23309) );
  NAND U23594 ( .A(x[244]), .B(y[2022]), .Z(n23308) );
  XNOR U23595 ( .A(n23309), .B(n23308), .Z(n23233) );
  NAND U23596 ( .A(x[247]), .B(y[2019]), .Z(n23222) );
  XNOR U23597 ( .A(n23221), .B(n23222), .Z(n23223) );
  NAND U23598 ( .A(x[246]), .B(y[2020]), .Z(n23224) );
  XNOR U23599 ( .A(n23223), .B(n23224), .Z(n23234) );
  XOR U23600 ( .A(n23233), .B(n23234), .Z(n23235) );
  XNOR U23601 ( .A(n23236), .B(n23235), .Z(n23246) );
  AND U23602 ( .A(x[228]), .B(y[2038]), .Z(n23227) );
  XOR U23603 ( .A(n23228), .B(n23227), .Z(n23230) );
  AND U23604 ( .A(x[227]), .B(y[2039]), .Z(n23298) );
  AND U23605 ( .A(x[235]), .B(y[2031]), .Z(n23299) );
  XOR U23606 ( .A(n23298), .B(n23299), .Z(n23300) );
  AND U23607 ( .A(x[243]), .B(y[2023]), .Z(n23301) );
  XOR U23608 ( .A(n23300), .B(n23301), .Z(n23211) );
  XOR U23609 ( .A(n23212), .B(n23211), .Z(n23214) );
  NANDN U23610 ( .A(n23162), .B(n23161), .Z(n23166) );
  OR U23611 ( .A(n23164), .B(n23163), .Z(n23165) );
  AND U23612 ( .A(n23166), .B(n23165), .Z(n23213) );
  XNOR U23613 ( .A(n23214), .B(n23213), .Z(n23245) );
  XOR U23614 ( .A(n23246), .B(n23245), .Z(n23247) );
  XOR U23615 ( .A(n23248), .B(n23247), .Z(n23279) );
  XNOR U23616 ( .A(n23280), .B(n23279), .Z(n23284) );
  NAND U23617 ( .A(n23168), .B(n23167), .Z(n23172) );
  NAND U23618 ( .A(n23170), .B(n23169), .Z(n23171) );
  NAND U23619 ( .A(n23172), .B(n23171), .Z(n23327) );
  NAND U23620 ( .A(n23174), .B(n23173), .Z(n23178) );
  NAND U23621 ( .A(n23176), .B(n23175), .Z(n23177) );
  NAND U23622 ( .A(n23178), .B(n23177), .Z(n23325) );
  NAND U23623 ( .A(n23180), .B(n23179), .Z(n23184) );
  NANDN U23624 ( .A(n23182), .B(n23181), .Z(n23183) );
  NAND U23625 ( .A(n23184), .B(n23183), .Z(n23324) );
  XOR U23626 ( .A(n23325), .B(n23324), .Z(n23326) );
  XOR U23627 ( .A(n23327), .B(n23326), .Z(n23283) );
  XOR U23628 ( .A(n23284), .B(n23283), .Z(n23286) );
  XOR U23629 ( .A(n23285), .B(n23286), .Z(n23336) );
  XOR U23630 ( .A(n23337), .B(n23336), .Z(n23338) );
  XOR U23631 ( .A(n23339), .B(n23338), .Z(n23201) );
  XOR U23632 ( .A(n23202), .B(n23201), .Z(n23351) );
  XOR U23633 ( .A(n23352), .B(n23351), .Z(n23345) );
  OR U23634 ( .A(n23187), .B(n23185), .Z(n23191) );
  ANDN U23635 ( .B(n23187), .A(n23186), .Z(n23189) );
  OR U23636 ( .A(n23189), .B(n23188), .Z(n23190) );
  AND U23637 ( .A(n23191), .B(n23190), .Z(n23343) );
  NAND U23638 ( .A(n23193), .B(n23192), .Z(n23197) );
  NANDN U23639 ( .A(n23195), .B(n23194), .Z(n23196) );
  AND U23640 ( .A(n23197), .B(n23196), .Z(n23344) );
  IV U23641 ( .A(n23344), .Z(n23342) );
  XOR U23642 ( .A(n23343), .B(n23342), .Z(n23198) );
  XNOR U23643 ( .A(n23345), .B(n23198), .Z(N507) );
  NAND U23644 ( .A(n23200), .B(n23199), .Z(n23204) );
  NAND U23645 ( .A(n23202), .B(n23201), .Z(n23203) );
  AND U23646 ( .A(n23204), .B(n23203), .Z(n23513) );
  NANDN U23647 ( .A(n23206), .B(n23205), .Z(n23210) );
  NAND U23648 ( .A(n23208), .B(n23207), .Z(n23209) );
  AND U23649 ( .A(n23210), .B(n23209), .Z(n23485) );
  AND U23650 ( .A(n23216), .B(n23215), .Z(n23220) );
  NAND U23651 ( .A(n23218), .B(n23217), .Z(n23219) );
  NANDN U23652 ( .A(n23220), .B(n23219), .Z(n23381) );
  NANDN U23653 ( .A(n23222), .B(n23221), .Z(n23226) );
  NANDN U23654 ( .A(n23224), .B(n23223), .Z(n23225) );
  NAND U23655 ( .A(n23226), .B(n23225), .Z(n23380) );
  XOR U23656 ( .A(n23381), .B(n23380), .Z(n23383) );
  NAND U23657 ( .A(n23228), .B(n23227), .Z(n23232) );
  ANDN U23658 ( .B(n23230), .A(n23229), .Z(n23231) );
  ANDN U23659 ( .B(n23232), .A(n23231), .Z(n23395) );
  AND U23660 ( .A(x[224]), .B(y[2043]), .Z(n23471) );
  AND U23661 ( .A(x[251]), .B(y[2016]), .Z(n23472) );
  XOR U23662 ( .A(n23471), .B(n23472), .Z(n23474) );
  AND U23663 ( .A(x[250]), .B(y[2017]), .Z(n23462) );
  XOR U23664 ( .A(o[251]), .B(n23462), .Z(n23473) );
  XOR U23665 ( .A(n23474), .B(n23473), .Z(n23393) );
  AND U23666 ( .A(x[233]), .B(y[2034]), .Z(n23456) );
  AND U23667 ( .A(x[245]), .B(y[2022]), .Z(n23457) );
  XOR U23668 ( .A(n23456), .B(n23457), .Z(n23458) );
  AND U23669 ( .A(x[242]), .B(y[2025]), .Z(n23459) );
  XOR U23670 ( .A(n23458), .B(n23459), .Z(n23392) );
  XOR U23671 ( .A(n23393), .B(n23392), .Z(n23394) );
  XOR U23672 ( .A(n23383), .B(n23382), .Z(n23483) );
  XOR U23673 ( .A(n23484), .B(n23483), .Z(n23486) );
  XOR U23674 ( .A(n23485), .B(n23486), .Z(n23504) );
  NAND U23675 ( .A(n23234), .B(n23233), .Z(n23238) );
  NAND U23676 ( .A(n23236), .B(n23235), .Z(n23237) );
  AND U23677 ( .A(n23238), .B(n23237), .Z(n23501) );
  NAND U23678 ( .A(n23240), .B(n23239), .Z(n23244) );
  NAND U23679 ( .A(n23242), .B(n23241), .Z(n23243) );
  NAND U23680 ( .A(n23244), .B(n23243), .Z(n23502) );
  NAND U23681 ( .A(n23246), .B(n23245), .Z(n23250) );
  NAND U23682 ( .A(n23248), .B(n23247), .Z(n23249) );
  AND U23683 ( .A(n23250), .B(n23249), .Z(n23489) );
  NANDN U23684 ( .A(n23252), .B(n23251), .Z(n23256) );
  NAND U23685 ( .A(n23254), .B(n23253), .Z(n23255) );
  AND U23686 ( .A(n23256), .B(n23255), .Z(n23480) );
  NANDN U23687 ( .A(n23258), .B(n23257), .Z(n23262) );
  NANDN U23688 ( .A(n23260), .B(n23259), .Z(n23261) );
  AND U23689 ( .A(n23262), .B(n23261), .Z(n23478) );
  AND U23690 ( .A(x[243]), .B(y[2024]), .Z(n23450) );
  AND U23691 ( .A(x[249]), .B(y[2018]), .Z(n23451) );
  XOR U23692 ( .A(n23450), .B(n23451), .Z(n23452) );
  AND U23693 ( .A(x[230]), .B(y[2037]), .Z(n23453) );
  XOR U23694 ( .A(n23452), .B(n23453), .Z(n23440) );
  AND U23695 ( .A(x[239]), .B(y[2028]), .Z(n23415) );
  NAND U23696 ( .A(x[226]), .B(y[2041]), .Z(n23416) );
  NAND U23697 ( .A(x[227]), .B(y[2040]), .Z(n23418) );
  XOR U23698 ( .A(n23440), .B(n23439), .Z(n23442) );
  NAND U23699 ( .A(x[240]), .B(y[2027]), .Z(n23398) );
  XNOR U23700 ( .A(n23398), .B(n23399), .Z(n23400) );
  XNOR U23701 ( .A(n23263), .B(n23400), .Z(n23411) );
  AND U23702 ( .A(y[2030]), .B(x[237]), .Z(n23265) );
  NAND U23703 ( .A(y[2031]), .B(x[236]), .Z(n23264) );
  XNOR U23704 ( .A(n23265), .B(n23264), .Z(n23412) );
  XOR U23705 ( .A(n23411), .B(n23412), .Z(n23441) );
  XOR U23706 ( .A(n23442), .B(n23441), .Z(n23377) );
  AND U23707 ( .A(n23267), .B(n23266), .Z(n23270) );
  NAND U23708 ( .A(n23410), .B(n23268), .Z(n23269) );
  NANDN U23709 ( .A(n23270), .B(n23269), .Z(n23375) );
  NANDN U23710 ( .A(n23272), .B(n23271), .Z(n23276) );
  NANDN U23711 ( .A(n23274), .B(n23273), .Z(n23275) );
  NAND U23712 ( .A(n23276), .B(n23275), .Z(n23374) );
  XOR U23713 ( .A(n23375), .B(n23374), .Z(n23376) );
  XOR U23714 ( .A(n23377), .B(n23376), .Z(n23477) );
  XNOR U23715 ( .A(n23478), .B(n23477), .Z(n23479) );
  XOR U23716 ( .A(n23480), .B(n23479), .Z(n23490) );
  NAND U23717 ( .A(n23278), .B(n23277), .Z(n23282) );
  NAND U23718 ( .A(n23280), .B(n23279), .Z(n23281) );
  NAND U23719 ( .A(n23282), .B(n23281), .Z(n23492) );
  NAND U23720 ( .A(n23284), .B(n23283), .Z(n23288) );
  NAND U23721 ( .A(n23286), .B(n23285), .Z(n23287) );
  NAND U23722 ( .A(n23288), .B(n23287), .Z(n23364) );
  XOR U23723 ( .A(n23365), .B(n23364), .Z(n23359) );
  NAND U23724 ( .A(n23290), .B(n23289), .Z(n23294) );
  NAND U23725 ( .A(n23292), .B(n23291), .Z(n23293) );
  AND U23726 ( .A(n23294), .B(n23293), .Z(n23369) );
  NAND U23727 ( .A(n23299), .B(n23298), .Z(n23303) );
  NAND U23728 ( .A(n23301), .B(n23300), .Z(n23302) );
  AND U23729 ( .A(n23303), .B(n23302), .Z(n23435) );
  AND U23730 ( .A(y[2019]), .B(x[248]), .Z(n23305) );
  NAND U23731 ( .A(y[2023]), .B(x[244]), .Z(n23304) );
  XNOR U23732 ( .A(n23305), .B(n23304), .Z(n23446) );
  AND U23733 ( .A(x[231]), .B(y[2036]), .Z(n23447) );
  XOR U23734 ( .A(n23446), .B(n23447), .Z(n23433) );
  AND U23735 ( .A(x[232]), .B(y[2035]), .Z(n23404) );
  NAND U23736 ( .A(x[247]), .B(y[2020]), .Z(n23405) );
  XNOR U23737 ( .A(n23404), .B(n23405), .Z(n23406) );
  NAND U23738 ( .A(x[246]), .B(y[2021]), .Z(n23407) );
  XOR U23739 ( .A(n23406), .B(n23407), .Z(n23434) );
  XOR U23740 ( .A(n23433), .B(n23434), .Z(n23436) );
  XOR U23741 ( .A(n23435), .B(n23436), .Z(n23496) );
  NAND U23742 ( .A(n23307), .B(n23306), .Z(n23311) );
  ANDN U23743 ( .B(n23309), .A(n23308), .Z(n23310) );
  ANDN U23744 ( .B(n23311), .A(n23310), .Z(n23428) );
  NAND U23745 ( .A(n23313), .B(n23312), .Z(n23317) );
  NAND U23746 ( .A(n23315), .B(n23314), .Z(n23316) );
  NAND U23747 ( .A(n23317), .B(n23316), .Z(n23427) );
  XNOR U23748 ( .A(n23428), .B(n23427), .Z(n23430) );
  AND U23749 ( .A(x[232]), .B(y[2036]), .Z(n23464) );
  NAND U23750 ( .A(n23318), .B(n23464), .Z(n23322) );
  NAND U23751 ( .A(n23320), .B(n23319), .Z(n23321) );
  AND U23752 ( .A(n23322), .B(n23321), .Z(n23389) );
  AND U23753 ( .A(x[238]), .B(y[2029]), .Z(n23421) );
  NAND U23754 ( .A(x[225]), .B(y[2042]), .Z(n23422) );
  AND U23755 ( .A(o[250]), .B(n23323), .Z(n23423) );
  XOR U23756 ( .A(n23424), .B(n23423), .Z(n23386) );
  AND U23757 ( .A(x[241]), .B(y[2026]), .Z(n23465) );
  AND U23758 ( .A(x[228]), .B(y[2039]), .Z(n23466) );
  XOR U23759 ( .A(n23465), .B(n23466), .Z(n23468) );
  AND U23760 ( .A(x[229]), .B(y[2038]), .Z(n23467) );
  XNOR U23761 ( .A(n23468), .B(n23467), .Z(n23387) );
  XNOR U23762 ( .A(n23386), .B(n23387), .Z(n23388) );
  XNOR U23763 ( .A(n23389), .B(n23388), .Z(n23429) );
  XNOR U23764 ( .A(n23430), .B(n23429), .Z(n23495) );
  XOR U23765 ( .A(n23498), .B(n23497), .Z(n23368) );
  NAND U23766 ( .A(n23325), .B(n23324), .Z(n23329) );
  NAND U23767 ( .A(n23327), .B(n23326), .Z(n23328) );
  NAND U23768 ( .A(n23329), .B(n23328), .Z(n23371) );
  NAND U23769 ( .A(n23331), .B(n23330), .Z(n23335) );
  NAND U23770 ( .A(n23333), .B(n23332), .Z(n23334) );
  AND U23771 ( .A(n23335), .B(n23334), .Z(n23356) );
  XOR U23772 ( .A(n23357), .B(n23356), .Z(n23358) );
  XNOR U23773 ( .A(n23359), .B(n23358), .Z(n23511) );
  NAND U23774 ( .A(n23337), .B(n23336), .Z(n23341) );
  NAND U23775 ( .A(n23339), .B(n23338), .Z(n23340) );
  AND U23776 ( .A(n23341), .B(n23340), .Z(n23510) );
  XOR U23777 ( .A(n23511), .B(n23510), .Z(n23512) );
  XNOR U23778 ( .A(n23513), .B(n23512), .Z(n23509) );
  NANDN U23779 ( .A(n23342), .B(n23343), .Z(n23348) );
  NOR U23780 ( .A(n23344), .B(n23343), .Z(n23346) );
  OR U23781 ( .A(n23346), .B(n23345), .Z(n23347) );
  AND U23782 ( .A(n23348), .B(n23347), .Z(n23508) );
  NAND U23783 ( .A(n23350), .B(n23349), .Z(n23354) );
  NAND U23784 ( .A(n23352), .B(n23351), .Z(n23353) );
  AND U23785 ( .A(n23354), .B(n23353), .Z(n23507) );
  XOR U23786 ( .A(n23508), .B(n23507), .Z(n23355) );
  XNOR U23787 ( .A(n23509), .B(n23355), .Z(N508) );
  NAND U23788 ( .A(n23357), .B(n23356), .Z(n23361) );
  NAND U23789 ( .A(n23359), .B(n23358), .Z(n23360) );
  NAND U23790 ( .A(n23361), .B(n23360), .Z(n23678) );
  NANDN U23791 ( .A(n23363), .B(n23362), .Z(n23367) );
  NAND U23792 ( .A(n23365), .B(n23364), .Z(n23366) );
  NAND U23793 ( .A(n23367), .B(n23366), .Z(n23677) );
  XOR U23794 ( .A(n23678), .B(n23677), .Z(n23680) );
  NANDN U23795 ( .A(n23369), .B(n23368), .Z(n23373) );
  NANDN U23796 ( .A(n23371), .B(n23370), .Z(n23372) );
  AND U23797 ( .A(n23373), .B(n23372), .Z(n23518) );
  NAND U23798 ( .A(n23375), .B(n23374), .Z(n23379) );
  NAND U23799 ( .A(n23377), .B(n23376), .Z(n23378) );
  AND U23800 ( .A(n23379), .B(n23378), .Z(n23530) );
  NAND U23801 ( .A(n23381), .B(n23380), .Z(n23385) );
  NAND U23802 ( .A(n23383), .B(n23382), .Z(n23384) );
  AND U23803 ( .A(n23385), .B(n23384), .Z(n23635) );
  NANDN U23804 ( .A(n23387), .B(n23386), .Z(n23391) );
  NANDN U23805 ( .A(n23389), .B(n23388), .Z(n23390) );
  AND U23806 ( .A(n23391), .B(n23390), .Z(n23633) );
  NAND U23807 ( .A(n23393), .B(n23392), .Z(n23397) );
  NANDN U23808 ( .A(n23395), .B(n23394), .Z(n23396) );
  NAND U23809 ( .A(n23397), .B(n23396), .Z(n23632) );
  NANDN U23810 ( .A(n23399), .B(n23398), .Z(n23403) );
  NANDN U23811 ( .A(n23401), .B(n23400), .Z(n23402) );
  AND U23812 ( .A(n23403), .B(n23402), .Z(n23611) );
  AND U23813 ( .A(x[231]), .B(y[2037]), .Z(n23577) );
  AND U23814 ( .A(x[236]), .B(y[2032]), .Z(n23576) );
  XOR U23815 ( .A(n23577), .B(n23576), .Z(n23579) );
  AND U23816 ( .A(x[235]), .B(y[2033]), .Z(n23578) );
  XOR U23817 ( .A(n23579), .B(n23578), .Z(n23609) );
  AND U23818 ( .A(x[251]), .B(y[2017]), .Z(n23593) );
  XOR U23819 ( .A(o[252]), .B(n23593), .Z(n23600) );
  NAND U23820 ( .A(x[250]), .B(y[2018]), .Z(n23601) );
  AND U23821 ( .A(x[239]), .B(y[2029]), .Z(n23602) );
  XNOR U23822 ( .A(n23603), .B(n23602), .Z(n23608) );
  NANDN U23823 ( .A(n23405), .B(n23404), .Z(n23409) );
  NANDN U23824 ( .A(n23407), .B(n23406), .Z(n23408) );
  AND U23825 ( .A(n23409), .B(n23408), .Z(n23617) );
  AND U23826 ( .A(x[241]), .B(y[2027]), .Z(n23542) );
  AND U23827 ( .A(x[246]), .B(y[2022]), .Z(n23541) );
  XOR U23828 ( .A(n23542), .B(n23541), .Z(n23544) );
  AND U23829 ( .A(x[228]), .B(y[2040]), .Z(n23543) );
  XOR U23830 ( .A(n23544), .B(n23543), .Z(n23615) );
  AND U23831 ( .A(x[230]), .B(y[2038]), .Z(n23783) );
  NAND U23832 ( .A(x[243]), .B(y[2025]), .Z(n23582) );
  XOR U23833 ( .A(n23615), .B(n23614), .Z(n23616) );
  XOR U23834 ( .A(n23656), .B(n23657), .Z(n23659) );
  NAND U23835 ( .A(n23594), .B(n23410), .Z(n23414) );
  NAND U23836 ( .A(n23412), .B(n23411), .Z(n23413) );
  AND U23837 ( .A(n23414), .B(n23413), .Z(n23538) );
  NANDN U23838 ( .A(n23416), .B(n23415), .Z(n23420) );
  NANDN U23839 ( .A(n23418), .B(n23417), .Z(n23419) );
  AND U23840 ( .A(n23420), .B(n23419), .Z(n23536) );
  NANDN U23841 ( .A(n23422), .B(n23421), .Z(n23426) );
  NAND U23842 ( .A(n23424), .B(n23423), .Z(n23425) );
  NAND U23843 ( .A(n23426), .B(n23425), .Z(n23535) );
  XOR U23844 ( .A(n23659), .B(n23658), .Z(n23531) );
  XNOR U23845 ( .A(n23532), .B(n23531), .Z(n23664) );
  NANDN U23846 ( .A(n23428), .B(n23427), .Z(n23432) );
  NAND U23847 ( .A(n23430), .B(n23429), .Z(n23431) );
  NAND U23848 ( .A(n23432), .B(n23431), .Z(n23623) );
  NANDN U23849 ( .A(n23434), .B(n23433), .Z(n23438) );
  OR U23850 ( .A(n23436), .B(n23435), .Z(n23437) );
  AND U23851 ( .A(n23438), .B(n23437), .Z(n23621) );
  NAND U23852 ( .A(n23440), .B(n23439), .Z(n23444) );
  NAND U23853 ( .A(n23442), .B(n23441), .Z(n23443) );
  NAND U23854 ( .A(n23444), .B(n23443), .Z(n23620) );
  XNOR U23855 ( .A(n23623), .B(n23622), .Z(n23662) );
  AND U23856 ( .A(x[248]), .B(y[2023]), .Z(n24010) );
  AND U23857 ( .A(x[244]), .B(y[2019]), .Z(n23445) );
  NAND U23858 ( .A(n24010), .B(n23445), .Z(n23449) );
  NAND U23859 ( .A(n23447), .B(n23446), .Z(n23448) );
  AND U23860 ( .A(n23449), .B(n23448), .Z(n23653) );
  AND U23861 ( .A(x[249]), .B(y[2019]), .Z(n23572) );
  XOR U23862 ( .A(n23573), .B(n23572), .Z(n23571) );
  NAND U23863 ( .A(x[225]), .B(y[2043]), .Z(n23570) );
  AND U23864 ( .A(x[240]), .B(y[2028]), .Z(n23564) );
  NAND U23865 ( .A(x[248]), .B(y[2020]), .Z(n23565) );
  NAND U23866 ( .A(x[226]), .B(y[2042]), .Z(n23567) );
  XOR U23867 ( .A(n23651), .B(n23650), .Z(n23652) );
  NAND U23868 ( .A(n23451), .B(n23450), .Z(n23455) );
  NAND U23869 ( .A(n23453), .B(n23452), .Z(n23454) );
  AND U23870 ( .A(n23455), .B(n23454), .Z(n23647) );
  NAND U23871 ( .A(x[227]), .B(y[2041]), .Z(n23595) );
  NAND U23872 ( .A(x[247]), .B(y[2021]), .Z(n23597) );
  AND U23873 ( .A(x[229]), .B(y[2039]), .Z(n23587) );
  NAND U23874 ( .A(x[245]), .B(y[2023]), .Z(n23588) );
  NAND U23875 ( .A(x[244]), .B(y[2024]), .Z(n23590) );
  XOR U23876 ( .A(n23645), .B(n23644), .Z(n23646) );
  NAND U23877 ( .A(n23457), .B(n23456), .Z(n23461) );
  NAND U23878 ( .A(n23459), .B(n23458), .Z(n23460) );
  NAND U23879 ( .A(n23461), .B(n23460), .Z(n23560) );
  AND U23880 ( .A(x[224]), .B(y[2044]), .Z(n23548) );
  AND U23881 ( .A(x[252]), .B(y[2016]), .Z(n23547) );
  XOR U23882 ( .A(n23548), .B(n23547), .Z(n23550) );
  AND U23883 ( .A(n23462), .B(o[251]), .Z(n23549) );
  XOR U23884 ( .A(n23550), .B(n23549), .Z(n23559) );
  NAND U23885 ( .A(y[2034]), .B(x[234]), .Z(n23463) );
  XNOR U23886 ( .A(n23464), .B(n23463), .Z(n23555) );
  AND U23887 ( .A(x[233]), .B(y[2035]), .Z(n23554) );
  XOR U23888 ( .A(n23555), .B(n23554), .Z(n23558) );
  XOR U23889 ( .A(n23559), .B(n23558), .Z(n23561) );
  XOR U23890 ( .A(n23560), .B(n23561), .Z(n23641) );
  NAND U23891 ( .A(n23466), .B(n23465), .Z(n23470) );
  NAND U23892 ( .A(n23468), .B(n23467), .Z(n23469) );
  AND U23893 ( .A(n23470), .B(n23469), .Z(n23639) );
  NAND U23894 ( .A(n23472), .B(n23471), .Z(n23476) );
  NAND U23895 ( .A(n23474), .B(n23473), .Z(n23475) );
  NAND U23896 ( .A(n23476), .B(n23475), .Z(n23638) );
  XNOR U23897 ( .A(n23641), .B(n23640), .Z(n23626) );
  XOR U23898 ( .A(n23627), .B(n23626), .Z(n23629) );
  XOR U23899 ( .A(n23628), .B(n23629), .Z(n23663) );
  XNOR U23900 ( .A(n23662), .B(n23663), .Z(n23665) );
  XOR U23901 ( .A(n23664), .B(n23665), .Z(n23671) );
  NANDN U23902 ( .A(n23478), .B(n23477), .Z(n23482) );
  NANDN U23903 ( .A(n23480), .B(n23479), .Z(n23481) );
  AND U23904 ( .A(n23482), .B(n23481), .Z(n23669) );
  NANDN U23905 ( .A(n23484), .B(n23483), .Z(n23488) );
  OR U23906 ( .A(n23486), .B(n23485), .Z(n23487) );
  NAND U23907 ( .A(n23488), .B(n23487), .Z(n23668) );
  XNOR U23908 ( .A(n23669), .B(n23668), .Z(n23670) );
  XOR U23909 ( .A(n23671), .B(n23670), .Z(n23517) );
  XOR U23910 ( .A(n23518), .B(n23517), .Z(n23520) );
  NANDN U23911 ( .A(n23490), .B(n23489), .Z(n23494) );
  NANDN U23912 ( .A(n23492), .B(n23491), .Z(n23493) );
  AND U23913 ( .A(n23494), .B(n23493), .Z(n23526) );
  NANDN U23914 ( .A(n23496), .B(n23495), .Z(n23500) );
  NAND U23915 ( .A(n23498), .B(n23497), .Z(n23499) );
  AND U23916 ( .A(n23500), .B(n23499), .Z(n23523) );
  NANDN U23917 ( .A(n23502), .B(n23501), .Z(n23506) );
  NANDN U23918 ( .A(n23504), .B(n23503), .Z(n23505) );
  NAND U23919 ( .A(n23506), .B(n23505), .Z(n23524) );
  XOR U23920 ( .A(n23520), .B(n23519), .Z(n23679) );
  XNOR U23921 ( .A(n23680), .B(n23679), .Z(n23676) );
  NAND U23922 ( .A(n23511), .B(n23510), .Z(n23515) );
  NAND U23923 ( .A(n23513), .B(n23512), .Z(n23514) );
  AND U23924 ( .A(n23515), .B(n23514), .Z(n23675) );
  XOR U23925 ( .A(n23674), .B(n23675), .Z(n23516) );
  XNOR U23926 ( .A(n23676), .B(n23516), .Z(N509) );
  NAND U23927 ( .A(n23518), .B(n23517), .Z(n23522) );
  NAND U23928 ( .A(n23520), .B(n23519), .Z(n23521) );
  AND U23929 ( .A(n23522), .B(n23521), .Z(n23690) );
  NANDN U23930 ( .A(n23524), .B(n23523), .Z(n23528) );
  NANDN U23931 ( .A(n23526), .B(n23525), .Z(n23527) );
  AND U23932 ( .A(n23528), .B(n23527), .Z(n23688) );
  NANDN U23933 ( .A(n23530), .B(n23529), .Z(n23534) );
  NAND U23934 ( .A(n23532), .B(n23531), .Z(n23533) );
  AND U23935 ( .A(n23534), .B(n23533), .Z(n23706) );
  NANDN U23936 ( .A(n23536), .B(n23535), .Z(n23540) );
  NANDN U23937 ( .A(n23538), .B(n23537), .Z(n23539) );
  AND U23938 ( .A(n23540), .B(n23539), .Z(n23817) );
  NAND U23939 ( .A(n23542), .B(n23541), .Z(n23546) );
  NAND U23940 ( .A(n23544), .B(n23543), .Z(n23545) );
  NAND U23941 ( .A(n23546), .B(n23545), .Z(n23854) );
  NAND U23942 ( .A(n23548), .B(n23547), .Z(n23552) );
  NAND U23943 ( .A(n23550), .B(n23549), .Z(n23551) );
  NAND U23944 ( .A(n23552), .B(n23551), .Z(n23853) );
  XOR U23945 ( .A(n23854), .B(n23853), .Z(n23855) );
  AND U23946 ( .A(y[2036]), .B(x[234]), .Z(n23851) );
  NAND U23947 ( .A(n23553), .B(n23851), .Z(n23557) );
  NAND U23948 ( .A(n23555), .B(n23554), .Z(n23556) );
  NAND U23949 ( .A(n23557), .B(n23556), .Z(n23822) );
  AND U23950 ( .A(x[246]), .B(y[2023]), .Z(n23761) );
  AND U23951 ( .A(x[225]), .B(y[2044]), .Z(n23759) );
  NAND U23952 ( .A(x[236]), .B(y[2033]), .Z(n23990) );
  XOR U23953 ( .A(n23761), .B(n23760), .Z(n23821) );
  NAND U23954 ( .A(x[239]), .B(y[2030]), .Z(n23764) );
  XOR U23955 ( .A(n23821), .B(n23820), .Z(n23823) );
  XNOR U23956 ( .A(n23822), .B(n23823), .Z(n23856) );
  NAND U23957 ( .A(n23559), .B(n23558), .Z(n23563) );
  NAND U23958 ( .A(n23561), .B(n23560), .Z(n23562) );
  AND U23959 ( .A(n23563), .B(n23562), .Z(n23814) );
  XOR U23960 ( .A(n23817), .B(n23816), .Z(n23811) );
  NANDN U23961 ( .A(n23565), .B(n23564), .Z(n23569) );
  NANDN U23962 ( .A(n23567), .B(n23566), .Z(n23568) );
  NAND U23963 ( .A(n23569), .B(n23568), .Z(n23827) );
  ANDN U23964 ( .B(n23571), .A(n23570), .Z(n23575) );
  NAND U23965 ( .A(n23573), .B(n23572), .Z(n23574) );
  NANDN U23966 ( .A(n23575), .B(n23574), .Z(n23826) );
  XOR U23967 ( .A(n23827), .B(n23826), .Z(n23828) );
  NAND U23968 ( .A(n23577), .B(n23576), .Z(n23581) );
  NAND U23969 ( .A(n23579), .B(n23578), .Z(n23580) );
  NAND U23970 ( .A(n23581), .B(n23580), .Z(n23725) );
  AND U23971 ( .A(x[235]), .B(y[2034]), .Z(n23780) );
  AND U23972 ( .A(x[227]), .B(y[2042]), .Z(n23778) );
  AND U23973 ( .A(x[241]), .B(y[2028]), .Z(n23777) );
  XOR U23974 ( .A(n23778), .B(n23777), .Z(n23779) );
  XOR U23975 ( .A(n23780), .B(n23779), .Z(n23724) );
  AND U23976 ( .A(x[247]), .B(y[2022]), .Z(n23774) );
  AND U23977 ( .A(x[237]), .B(y[2032]), .Z(n23772) );
  AND U23978 ( .A(x[248]), .B(y[2021]), .Z(n23970) );
  XOR U23979 ( .A(n23772), .B(n23970), .Z(n23773) );
  XOR U23980 ( .A(n23774), .B(n23773), .Z(n23723) );
  XOR U23981 ( .A(n23724), .B(n23723), .Z(n23726) );
  XNOR U23982 ( .A(n23725), .B(n23726), .Z(n23829) );
  NANDN U23983 ( .A(n23582), .B(n23783), .Z(n23586) );
  NANDN U23984 ( .A(n23584), .B(n23583), .Z(n23585) );
  AND U23985 ( .A(n23586), .B(n23585), .Z(n23834) );
  AND U23986 ( .A(x[249]), .B(y[2020]), .Z(n23756) );
  AND U23987 ( .A(x[250]), .B(y[2019]), .Z(n23753) );
  XOR U23988 ( .A(n23754), .B(n23753), .Z(n23755) );
  XOR U23989 ( .A(n23756), .B(n23755), .Z(n23833) );
  AND U23990 ( .A(x[252]), .B(y[2017]), .Z(n23771) );
  XOR U23991 ( .A(o[253]), .B(n23771), .Z(n23846) );
  AND U23992 ( .A(x[224]), .B(y[2045]), .Z(n23844) );
  AND U23993 ( .A(x[253]), .B(y[2016]), .Z(n23843) );
  XOR U23994 ( .A(n23844), .B(n23843), .Z(n23845) );
  XNOR U23995 ( .A(n23846), .B(n23845), .Z(n23832) );
  XNOR U23996 ( .A(n23834), .B(n23835), .Z(n23802) );
  NANDN U23997 ( .A(n23588), .B(n23587), .Z(n23592) );
  NANDN U23998 ( .A(n23590), .B(n23589), .Z(n23591) );
  NAND U23999 ( .A(n23592), .B(n23591), .Z(n23792) );
  AND U24000 ( .A(o[252]), .B(n23593), .Z(n23732) );
  AND U24001 ( .A(x[240]), .B(y[2029]), .Z(n23730) );
  AND U24002 ( .A(x[251]), .B(y[2018]), .Z(n23729) );
  XOR U24003 ( .A(n23730), .B(n23729), .Z(n23731) );
  XOR U24004 ( .A(n23732), .B(n23731), .Z(n23791) );
  AND U24005 ( .A(x[226]), .B(y[2043]), .Z(n23742) );
  XOR U24006 ( .A(n23742), .B(n23741), .Z(n23743) );
  XOR U24007 ( .A(n23744), .B(n23743), .Z(n23790) );
  XOR U24008 ( .A(n23791), .B(n23790), .Z(n23793) );
  XOR U24009 ( .A(n23792), .B(n23793), .Z(n23803) );
  NANDN U24010 ( .A(n23595), .B(n23594), .Z(n23599) );
  NANDN U24011 ( .A(n23597), .B(n23596), .Z(n23598) );
  NAND U24012 ( .A(n23599), .B(n23598), .Z(n23748) );
  NANDN U24013 ( .A(n23601), .B(n23600), .Z(n23605) );
  NAND U24014 ( .A(n23603), .B(n23602), .Z(n23604) );
  NAND U24015 ( .A(n23605), .B(n23604), .Z(n23747) );
  XOR U24016 ( .A(n23748), .B(n23747), .Z(n23750) );
  AND U24017 ( .A(x[233]), .B(y[2036]), .Z(n23985) );
  AND U24018 ( .A(x[232]), .B(y[2037]), .Z(n23785) );
  AND U24019 ( .A(y[2039]), .B(x[230]), .Z(n23607) );
  NAND U24020 ( .A(y[2038]), .B(x[231]), .Z(n23606) );
  XNOR U24021 ( .A(n23607), .B(n23606), .Z(n23784) );
  XOR U24022 ( .A(n23785), .B(n23784), .Z(n23838) );
  XOR U24023 ( .A(n23985), .B(n23838), .Z(n23840) );
  AND U24024 ( .A(x[229]), .B(y[2040]), .Z(n23738) );
  AND U24025 ( .A(x[228]), .B(y[2041]), .Z(n23736) );
  AND U24026 ( .A(x[234]), .B(y[2035]), .Z(n23735) );
  XOR U24027 ( .A(n23736), .B(n23735), .Z(n23737) );
  XOR U24028 ( .A(n23738), .B(n23737), .Z(n23839) );
  XOR U24029 ( .A(n23840), .B(n23839), .Z(n23749) );
  XOR U24030 ( .A(n23750), .B(n23749), .Z(n23718) );
  NANDN U24031 ( .A(n23609), .B(n23608), .Z(n23613) );
  NANDN U24032 ( .A(n23611), .B(n23610), .Z(n23612) );
  NAND U24033 ( .A(n23613), .B(n23612), .Z(n23717) );
  XOR U24034 ( .A(n23720), .B(n23719), .Z(n23809) );
  NAND U24035 ( .A(n23615), .B(n23614), .Z(n23619) );
  NANDN U24036 ( .A(n23617), .B(n23616), .Z(n23618) );
  NAND U24037 ( .A(n23619), .B(n23618), .Z(n23808) );
  NANDN U24038 ( .A(n23621), .B(n23620), .Z(n23625) );
  NAND U24039 ( .A(n23623), .B(n23622), .Z(n23624) );
  AND U24040 ( .A(n23625), .B(n23624), .Z(n23700) );
  NAND U24041 ( .A(n23627), .B(n23626), .Z(n23631) );
  NAND U24042 ( .A(n23629), .B(n23628), .Z(n23630) );
  AND U24043 ( .A(n23631), .B(n23630), .Z(n23699) );
  NANDN U24044 ( .A(n23633), .B(n23632), .Z(n23637) );
  NANDN U24045 ( .A(n23635), .B(n23634), .Z(n23636) );
  NAND U24046 ( .A(n23637), .B(n23636), .Z(n23713) );
  NANDN U24047 ( .A(n23639), .B(n23638), .Z(n23643) );
  NAND U24048 ( .A(n23641), .B(n23640), .Z(n23642) );
  AND U24049 ( .A(n23643), .B(n23642), .Z(n23799) );
  NAND U24050 ( .A(n23645), .B(n23644), .Z(n23649) );
  NANDN U24051 ( .A(n23647), .B(n23646), .Z(n23648) );
  AND U24052 ( .A(n23649), .B(n23648), .Z(n23797) );
  NAND U24053 ( .A(n23651), .B(n23650), .Z(n23655) );
  NANDN U24054 ( .A(n23653), .B(n23652), .Z(n23654) );
  NAND U24055 ( .A(n23655), .B(n23654), .Z(n23796) );
  NAND U24056 ( .A(n23657), .B(n23656), .Z(n23661) );
  NAND U24057 ( .A(n23659), .B(n23658), .Z(n23660) );
  NAND U24058 ( .A(n23661), .B(n23660), .Z(n23711) );
  XOR U24059 ( .A(n23712), .B(n23711), .Z(n23714) );
  XOR U24060 ( .A(n23713), .B(n23714), .Z(n23701) );
  XOR U24061 ( .A(n23702), .B(n23701), .Z(n23707) );
  XOR U24062 ( .A(n23708), .B(n23707), .Z(n23695) );
  NAND U24063 ( .A(n23663), .B(n23662), .Z(n23667) );
  NANDN U24064 ( .A(n23665), .B(n23664), .Z(n23666) );
  AND U24065 ( .A(n23667), .B(n23666), .Z(n23694) );
  NANDN U24066 ( .A(n23669), .B(n23668), .Z(n23673) );
  NAND U24067 ( .A(n23671), .B(n23670), .Z(n23672) );
  AND U24068 ( .A(n23673), .B(n23672), .Z(n23693) );
  XOR U24069 ( .A(n23694), .B(n23693), .Z(n23696) );
  XNOR U24070 ( .A(n23695), .B(n23696), .Z(n23687) );
  XOR U24071 ( .A(n23690), .B(n23689), .Z(n23686) );
  NAND U24072 ( .A(n23678), .B(n23677), .Z(n23682) );
  NAND U24073 ( .A(n23680), .B(n23679), .Z(n23681) );
  NAND U24074 ( .A(n23682), .B(n23681), .Z(n23684) );
  XNOR U24075 ( .A(n23685), .B(n23684), .Z(n23683) );
  XNOR U24076 ( .A(n23686), .B(n23683), .Z(N510) );
  NANDN U24077 ( .A(n23688), .B(n23687), .Z(n23692) );
  NANDN U24078 ( .A(n23690), .B(n23689), .Z(n23691) );
  AND U24079 ( .A(n23692), .B(n23691), .Z(n24145) );
  NANDN U24080 ( .A(n23694), .B(n23693), .Z(n23698) );
  OR U24081 ( .A(n23696), .B(n23695), .Z(n23697) );
  AND U24082 ( .A(n23698), .B(n23697), .Z(n23860) );
  NANDN U24083 ( .A(n23700), .B(n23699), .Z(n23704) );
  NAND U24084 ( .A(n23702), .B(n23701), .Z(n23703) );
  AND U24085 ( .A(n23704), .B(n23703), .Z(n24152) );
  NANDN U24086 ( .A(n23706), .B(n23705), .Z(n23710) );
  NAND U24087 ( .A(n23708), .B(n23707), .Z(n23709) );
  AND U24088 ( .A(n23710), .B(n23709), .Z(n24151) );
  XOR U24089 ( .A(n24152), .B(n24151), .Z(n24150) );
  NAND U24090 ( .A(n23712), .B(n23711), .Z(n23716) );
  NAND U24091 ( .A(n23714), .B(n23713), .Z(n23715) );
  AND U24092 ( .A(n23716), .B(n23715), .Z(n24149) );
  XOR U24093 ( .A(n24150), .B(n24149), .Z(n23862) );
  NANDN U24094 ( .A(n23718), .B(n23717), .Z(n23722) );
  NAND U24095 ( .A(n23720), .B(n23719), .Z(n23721) );
  AND U24096 ( .A(n23722), .B(n23721), .Z(n24131) );
  NAND U24097 ( .A(n23724), .B(n23723), .Z(n23728) );
  NAND U24098 ( .A(n23726), .B(n23725), .Z(n23727) );
  AND U24099 ( .A(n23728), .B(n23727), .Z(n23873) );
  NAND U24100 ( .A(n23730), .B(n23729), .Z(n23734) );
  NAND U24101 ( .A(n23732), .B(n23731), .Z(n23733) );
  NAND U24102 ( .A(n23734), .B(n23733), .Z(n24073) );
  NAND U24103 ( .A(n23736), .B(n23735), .Z(n23740) );
  NAND U24104 ( .A(n23738), .B(n23737), .Z(n23739) );
  NAND U24105 ( .A(n23740), .B(n23739), .Z(n24076) );
  AND U24106 ( .A(x[230]), .B(y[2040]), .Z(n23955) );
  AND U24107 ( .A(x[229]), .B(y[2041]), .Z(n23957) );
  AND U24108 ( .A(x[243]), .B(y[2027]), .Z(n23956) );
  XOR U24109 ( .A(n23957), .B(n23956), .Z(n23954) );
  XNOR U24110 ( .A(n23955), .B(n23954), .Z(n23903) );
  AND U24111 ( .A(x[228]), .B(y[2042]), .Z(n23949) );
  AND U24112 ( .A(x[227]), .B(y[2043]), .Z(n23951) );
  AND U24113 ( .A(x[242]), .B(y[2028]), .Z(n23950) );
  XOR U24114 ( .A(n23951), .B(n23950), .Z(n23948) );
  XOR U24115 ( .A(n23949), .B(n23948), .Z(n23906) );
  NAND U24116 ( .A(n23742), .B(n23741), .Z(n23746) );
  NAND U24117 ( .A(n23744), .B(n23743), .Z(n23745) );
  AND U24118 ( .A(n23746), .B(n23745), .Z(n23905) );
  XOR U24119 ( .A(n23903), .B(n23904), .Z(n24075) );
  XOR U24120 ( .A(n24076), .B(n24075), .Z(n24074) );
  XOR U24121 ( .A(n24073), .B(n24074), .Z(n23874) );
  NAND U24122 ( .A(n23748), .B(n23747), .Z(n23752) );
  NAND U24123 ( .A(n23750), .B(n23749), .Z(n23751) );
  AND U24124 ( .A(n23752), .B(n23751), .Z(n23871) );
  XOR U24125 ( .A(n23872), .B(n23871), .Z(n24134) );
  AND U24126 ( .A(n23754), .B(n23753), .Z(n23758) );
  NAND U24127 ( .A(n23756), .B(n23755), .Z(n23757) );
  NANDN U24128 ( .A(n23758), .B(n23757), .Z(n24067) );
  NANDN U24129 ( .A(n23990), .B(n23759), .Z(n23763) );
  NAND U24130 ( .A(n23761), .B(n23760), .Z(n23762) );
  NAND U24131 ( .A(n23763), .B(n23762), .Z(n24070) );
  NANDN U24132 ( .A(n23764), .B(n23917), .Z(n23768) );
  NANDN U24133 ( .A(n23766), .B(n23765), .Z(n23767) );
  AND U24134 ( .A(n23768), .B(n23767), .Z(n23884) );
  AND U24135 ( .A(x[247]), .B(y[2023]), .Z(n23969) );
  AND U24136 ( .A(y[2022]), .B(x[248]), .Z(n23770) );
  AND U24137 ( .A(y[2021]), .B(x[249]), .Z(n23769) );
  XOR U24138 ( .A(n23770), .B(n23769), .Z(n23968) );
  XOR U24139 ( .A(n23969), .B(n23968), .Z(n23886) );
  AND U24140 ( .A(n23771), .B(o[253]), .Z(n23994) );
  AND U24141 ( .A(x[252]), .B(y[2018]), .Z(n23996) );
  AND U24142 ( .A(x[240]), .B(y[2030]), .Z(n23995) );
  XOR U24143 ( .A(n23996), .B(n23995), .Z(n23993) );
  XNOR U24144 ( .A(n23994), .B(n23993), .Z(n23885) );
  XNOR U24145 ( .A(n23884), .B(n23883), .Z(n24069) );
  XOR U24146 ( .A(n24070), .B(n24069), .Z(n24068) );
  XOR U24147 ( .A(n24067), .B(n24068), .Z(n24114) );
  NAND U24148 ( .A(n23772), .B(n23970), .Z(n23776) );
  NAND U24149 ( .A(n23774), .B(n23773), .Z(n23775) );
  NAND U24150 ( .A(n23776), .B(n23775), .Z(n24098) );
  NAND U24151 ( .A(n23778), .B(n23777), .Z(n23782) );
  NAND U24152 ( .A(n23780), .B(n23779), .Z(n23781) );
  AND U24153 ( .A(n23782), .B(n23781), .Z(n23910) );
  AND U24154 ( .A(x[224]), .B(y[2046]), .Z(n24002) );
  AND U24155 ( .A(x[253]), .B(y[2017]), .Z(n24007) );
  XOR U24156 ( .A(o[254]), .B(n24007), .Z(n24004) );
  AND U24157 ( .A(x[254]), .B(y[2016]), .Z(n24003) );
  XOR U24158 ( .A(n24004), .B(n24003), .Z(n24001) );
  XOR U24159 ( .A(n24002), .B(n24001), .Z(n23912) );
  AND U24160 ( .A(x[244]), .B(y[2026]), .Z(n23943) );
  XOR U24161 ( .A(n23943), .B(n23942), .Z(n23941) );
  AND U24162 ( .A(x[232]), .B(y[2038]), .Z(n23940) );
  XNOR U24163 ( .A(n23941), .B(n23940), .Z(n23911) );
  XNOR U24164 ( .A(n23910), .B(n23909), .Z(n24097) );
  XOR U24165 ( .A(n24098), .B(n24097), .Z(n24095) );
  AND U24166 ( .A(x[231]), .B(y[2039]), .Z(n23916) );
  NAND U24167 ( .A(n23783), .B(n23916), .Z(n23787) );
  NAND U24168 ( .A(n23785), .B(n23784), .Z(n23786) );
  AND U24169 ( .A(n23787), .B(n23786), .Z(n23895) );
  AND U24170 ( .A(y[2025]), .B(x[245]), .Z(n23789) );
  AND U24171 ( .A(y[2024]), .B(x[246]), .Z(n23788) );
  XOR U24172 ( .A(n23789), .B(n23788), .Z(n23915) );
  XOR U24173 ( .A(n23916), .B(n23915), .Z(n23898) );
  AND U24174 ( .A(x[241]), .B(y[2029]), .Z(n23935) );
  AND U24175 ( .A(x[226]), .B(y[2044]), .Z(n23937) );
  AND U24176 ( .A(x[250]), .B(y[2020]), .Z(n23936) );
  XOR U24177 ( .A(n23937), .B(n23936), .Z(n23934) );
  XNOR U24178 ( .A(n23935), .B(n23934), .Z(n23897) );
  XNOR U24179 ( .A(n23895), .B(n23896), .Z(n24096) );
  NAND U24180 ( .A(n23791), .B(n23790), .Z(n23795) );
  NAND U24181 ( .A(n23793), .B(n23792), .Z(n23794) );
  NAND U24182 ( .A(n23795), .B(n23794), .Z(n24115) );
  XOR U24183 ( .A(n24116), .B(n24115), .Z(n24113) );
  XOR U24184 ( .A(n24114), .B(n24113), .Z(n24133) );
  XNOR U24185 ( .A(n24131), .B(n24132), .Z(n24126) );
  NANDN U24186 ( .A(n23797), .B(n23796), .Z(n23801) );
  NANDN U24187 ( .A(n23799), .B(n23798), .Z(n23800) );
  AND U24188 ( .A(n23801), .B(n23800), .Z(n24128) );
  NANDN U24189 ( .A(n23803), .B(n23802), .Z(n23807) );
  NANDN U24190 ( .A(n23805), .B(n23804), .Z(n23806) );
  NAND U24191 ( .A(n23807), .B(n23806), .Z(n24127) );
  XOR U24192 ( .A(n24128), .B(n24127), .Z(n24125) );
  NANDN U24193 ( .A(n23809), .B(n23808), .Z(n23813) );
  NANDN U24194 ( .A(n23811), .B(n23810), .Z(n23812) );
  NAND U24195 ( .A(n23813), .B(n23812), .Z(n23867) );
  NANDN U24196 ( .A(n23815), .B(n23814), .Z(n23819) );
  NAND U24197 ( .A(n23817), .B(n23816), .Z(n23818) );
  AND U24198 ( .A(n23819), .B(n23818), .Z(n24107) );
  NAND U24199 ( .A(n23821), .B(n23820), .Z(n23825) );
  NAND U24200 ( .A(n23823), .B(n23822), .Z(n23824) );
  AND U24201 ( .A(n23825), .B(n23824), .Z(n23880) );
  NAND U24202 ( .A(n23827), .B(n23826), .Z(n23831) );
  NANDN U24203 ( .A(n23829), .B(n23828), .Z(n23830) );
  AND U24204 ( .A(n23831), .B(n23830), .Z(n23879) );
  XOR U24205 ( .A(n23880), .B(n23879), .Z(n23878) );
  NANDN U24206 ( .A(n23833), .B(n23832), .Z(n23837) );
  NANDN U24207 ( .A(n23835), .B(n23834), .Z(n23836) );
  NAND U24208 ( .A(n23837), .B(n23836), .Z(n23877) );
  XOR U24209 ( .A(n23878), .B(n23877), .Z(n24110) );
  NAND U24210 ( .A(n23985), .B(n23838), .Z(n23842) );
  NAND U24211 ( .A(n23840), .B(n23839), .Z(n23841) );
  AND U24212 ( .A(n23842), .B(n23841), .Z(n24091) );
  NAND U24213 ( .A(n23844), .B(n23843), .Z(n23848) );
  NAND U24214 ( .A(n23846), .B(n23845), .Z(n23847) );
  NAND U24215 ( .A(n23848), .B(n23847), .Z(n23889) );
  NAND U24216 ( .A(y[2034]), .B(x[236]), .Z(n23849) );
  XNOR U24217 ( .A(n23850), .B(n23849), .Z(n23989) );
  XOR U24218 ( .A(n23989), .B(n23988), .Z(n23984) );
  AND U24219 ( .A(y[2037]), .B(x[233]), .Z(n23852) );
  XOR U24220 ( .A(n23852), .B(n23851), .Z(n23983) );
  XOR U24221 ( .A(n23984), .B(n23983), .Z(n23892) );
  AND U24222 ( .A(x[251]), .B(y[2019]), .Z(n23965) );
  AND U24223 ( .A(x[225]), .B(y[2045]), .Z(n23964) );
  XOR U24224 ( .A(n23965), .B(n23964), .Z(n23963) );
  XOR U24225 ( .A(n23963), .B(n23962), .Z(n23891) );
  XOR U24226 ( .A(n23892), .B(n23891), .Z(n23890) );
  XOR U24227 ( .A(n23889), .B(n23890), .Z(n24092) );
  NAND U24228 ( .A(n23854), .B(n23853), .Z(n23858) );
  NANDN U24229 ( .A(n23856), .B(n23855), .Z(n23857) );
  AND U24230 ( .A(n23858), .B(n23857), .Z(n24089) );
  XNOR U24231 ( .A(n24090), .B(n24089), .Z(n24109) );
  XNOR U24232 ( .A(n24107), .B(n24108), .Z(n23868) );
  XOR U24233 ( .A(n23867), .B(n23868), .Z(n23865) );
  XNOR U24234 ( .A(n23860), .B(n23859), .Z(n24143) );
  XNOR U24235 ( .A(n24144), .B(n24143), .Z(N511) );
  NAND U24236 ( .A(n23860), .B(n23859), .Z(n23864) );
  NANDN U24237 ( .A(n23862), .B(n23861), .Z(n23863) );
  AND U24238 ( .A(n23864), .B(n23863), .Z(n24160) );
  NANDN U24239 ( .A(n23866), .B(n23865), .Z(n23870) );
  NAND U24240 ( .A(n23868), .B(n23867), .Z(n23869) );
  AND U24241 ( .A(n23870), .B(n23869), .Z(n24142) );
  NAND U24242 ( .A(n23872), .B(n23871), .Z(n23876) );
  NANDN U24243 ( .A(n23874), .B(n23873), .Z(n23875) );
  AND U24244 ( .A(n23876), .B(n23875), .Z(n24124) );
  NAND U24245 ( .A(n23878), .B(n23877), .Z(n23882) );
  NAND U24246 ( .A(n23880), .B(n23879), .Z(n23881) );
  AND U24247 ( .A(n23882), .B(n23881), .Z(n24106) );
  NAND U24248 ( .A(n23884), .B(n23883), .Z(n23888) );
  NANDN U24249 ( .A(n23886), .B(n23885), .Z(n23887) );
  AND U24250 ( .A(n23888), .B(n23887), .Z(n24088) );
  NAND U24251 ( .A(n23890), .B(n23889), .Z(n23894) );
  NAND U24252 ( .A(n23892), .B(n23891), .Z(n23893) );
  AND U24253 ( .A(n23894), .B(n23893), .Z(n23902) );
  NANDN U24254 ( .A(n23896), .B(n23895), .Z(n23900) );
  NANDN U24255 ( .A(n23898), .B(n23897), .Z(n23899) );
  NAND U24256 ( .A(n23900), .B(n23899), .Z(n23901) );
  XNOR U24257 ( .A(n23902), .B(n23901), .Z(n24086) );
  NANDN U24258 ( .A(n23904), .B(n23903), .Z(n23908) );
  NANDN U24259 ( .A(n23906), .B(n23905), .Z(n23907) );
  AND U24260 ( .A(n23908), .B(n23907), .Z(n24084) );
  NAND U24261 ( .A(n23910), .B(n23909), .Z(n23914) );
  NANDN U24262 ( .A(n23912), .B(n23911), .Z(n23913) );
  AND U24263 ( .A(n23914), .B(n23913), .Z(n24066) );
  NAND U24264 ( .A(n23916), .B(n23915), .Z(n23919) );
  AND U24265 ( .A(x[246]), .B(y[2025]), .Z(n24008) );
  AND U24266 ( .A(n23917), .B(n24008), .Z(n23918) );
  ANDN U24267 ( .B(n23919), .A(n23918), .Z(n23982) );
  AND U24268 ( .A(y[2033]), .B(x[238]), .Z(n23921) );
  NAND U24269 ( .A(y[2038]), .B(x[233]), .Z(n23920) );
  XNOR U24270 ( .A(n23921), .B(n23920), .Z(n23925) );
  AND U24271 ( .A(y[2046]), .B(x[225]), .Z(n23923) );
  NAND U24272 ( .A(y[2047]), .B(x[224]), .Z(n23922) );
  XNOR U24273 ( .A(n23923), .B(n23922), .Z(n23924) );
  XOR U24274 ( .A(n23925), .B(n23924), .Z(n23933) );
  AND U24275 ( .A(y[2036]), .B(x[235]), .Z(n23927) );
  NAND U24276 ( .A(y[2021]), .B(x[250]), .Z(n23926) );
  XNOR U24277 ( .A(n23927), .B(n23926), .Z(n23931) );
  AND U24278 ( .A(y[2031]), .B(x[240]), .Z(n23929) );
  NAND U24279 ( .A(y[2035]), .B(x[236]), .Z(n23928) );
  XNOR U24280 ( .A(n23929), .B(n23928), .Z(n23930) );
  XNOR U24281 ( .A(n23931), .B(n23930), .Z(n23932) );
  XNOR U24282 ( .A(n23933), .B(n23932), .Z(n23980) );
  NAND U24283 ( .A(n23935), .B(n23934), .Z(n23939) );
  NAND U24284 ( .A(n23937), .B(n23936), .Z(n23938) );
  AND U24285 ( .A(n23939), .B(n23938), .Z(n23947) );
  NAND U24286 ( .A(n23941), .B(n23940), .Z(n23945) );
  NAND U24287 ( .A(n23943), .B(n23942), .Z(n23944) );
  NAND U24288 ( .A(n23945), .B(n23944), .Z(n23946) );
  XNOR U24289 ( .A(n23947), .B(n23946), .Z(n23978) );
  NAND U24290 ( .A(n23949), .B(n23948), .Z(n23953) );
  NAND U24291 ( .A(n23951), .B(n23950), .Z(n23952) );
  AND U24292 ( .A(n23953), .B(n23952), .Z(n23961) );
  NAND U24293 ( .A(n23955), .B(n23954), .Z(n23959) );
  NAND U24294 ( .A(n23957), .B(n23956), .Z(n23958) );
  NAND U24295 ( .A(n23959), .B(n23958), .Z(n23960) );
  XNOR U24296 ( .A(n23961), .B(n23960), .Z(n23976) );
  NAND U24297 ( .A(n23963), .B(n23962), .Z(n23967) );
  NAND U24298 ( .A(n23965), .B(n23964), .Z(n23966) );
  AND U24299 ( .A(n23967), .B(n23966), .Z(n23974) );
  NAND U24300 ( .A(n23969), .B(n23968), .Z(n23972) );
  AND U24301 ( .A(x[249]), .B(y[2022]), .Z(n24009) );
  NAND U24302 ( .A(n23970), .B(n24009), .Z(n23971) );
  NAND U24303 ( .A(n23972), .B(n23971), .Z(n23973) );
  XNOR U24304 ( .A(n23974), .B(n23973), .Z(n23975) );
  XNOR U24305 ( .A(n23976), .B(n23975), .Z(n23977) );
  XNOR U24306 ( .A(n23978), .B(n23977), .Z(n23979) );
  XNOR U24307 ( .A(n23980), .B(n23979), .Z(n23981) );
  XNOR U24308 ( .A(n23982), .B(n23981), .Z(n24064) );
  NAND U24309 ( .A(n23984), .B(n23983), .Z(n23987) );
  AND U24310 ( .A(x[234]), .B(y[2037]), .Z(n24031) );
  NAND U24311 ( .A(n23985), .B(n24031), .Z(n23986) );
  AND U24312 ( .A(n23987), .B(n23986), .Z(n24062) );
  NAND U24313 ( .A(n23989), .B(n23988), .Z(n23992) );
  NANDN U24314 ( .A(n23990), .B(n24032), .Z(n23991) );
  AND U24315 ( .A(n23992), .B(n23991), .Z(n24000) );
  NAND U24316 ( .A(n23994), .B(n23993), .Z(n23998) );
  NAND U24317 ( .A(n23996), .B(n23995), .Z(n23997) );
  NAND U24318 ( .A(n23998), .B(n23997), .Z(n23999) );
  XNOR U24319 ( .A(n24000), .B(n23999), .Z(n24060) );
  NAND U24320 ( .A(n24002), .B(n24001), .Z(n24006) );
  NAND U24321 ( .A(n24004), .B(n24003), .Z(n24005) );
  AND U24322 ( .A(n24006), .B(n24005), .Z(n24058) );
  AND U24323 ( .A(y[2044]), .B(x[227]), .Z(n24016) );
  AND U24324 ( .A(n24007), .B(o[254]), .Z(n24014) );
  XOR U24325 ( .A(n24008), .B(o[255]), .Z(n24012) );
  XNOR U24326 ( .A(n24010), .B(n24009), .Z(n24011) );
  XNOR U24327 ( .A(n24012), .B(n24011), .Z(n24013) );
  XNOR U24328 ( .A(n24014), .B(n24013), .Z(n24015) );
  XNOR U24329 ( .A(n24016), .B(n24015), .Z(n24056) );
  AND U24330 ( .A(y[2019]), .B(x[252]), .Z(n24022) );
  AND U24331 ( .A(y[2020]), .B(x[251]), .Z(n24018) );
  NAND U24332 ( .A(y[2024]), .B(x[247]), .Z(n24017) );
  XNOR U24333 ( .A(n24018), .B(n24017), .Z(n24019) );
  XNOR U24334 ( .A(n24020), .B(n24019), .Z(n24021) );
  XNOR U24335 ( .A(n24022), .B(n24021), .Z(n24046) );
  AND U24336 ( .A(y[2028]), .B(x[243]), .Z(n24024) );
  NAND U24337 ( .A(y[2026]), .B(x[245]), .Z(n24023) );
  XNOR U24338 ( .A(n24024), .B(n24023), .Z(n24036) );
  AND U24339 ( .A(y[2039]), .B(x[232]), .Z(n24026) );
  NAND U24340 ( .A(y[2043]), .B(x[228]), .Z(n24025) );
  XNOR U24341 ( .A(n24026), .B(n24025), .Z(n24030) );
  AND U24342 ( .A(y[2016]), .B(x[255]), .Z(n24028) );
  NAND U24343 ( .A(y[2041]), .B(x[230]), .Z(n24027) );
  XNOR U24344 ( .A(n24028), .B(n24027), .Z(n24029) );
  XOR U24345 ( .A(n24030), .B(n24029), .Z(n24034) );
  XNOR U24346 ( .A(n24032), .B(n24031), .Z(n24033) );
  XNOR U24347 ( .A(n24034), .B(n24033), .Z(n24035) );
  XOR U24348 ( .A(n24036), .B(n24035), .Z(n24044) );
  AND U24349 ( .A(y[2017]), .B(x[254]), .Z(n24038) );
  NAND U24350 ( .A(y[2029]), .B(x[242]), .Z(n24037) );
  XNOR U24351 ( .A(n24038), .B(n24037), .Z(n24042) );
  AND U24352 ( .A(y[2018]), .B(x[253]), .Z(n24040) );
  NAND U24353 ( .A(y[2027]), .B(x[244]), .Z(n24039) );
  XNOR U24354 ( .A(n24040), .B(n24039), .Z(n24041) );
  XNOR U24355 ( .A(n24042), .B(n24041), .Z(n24043) );
  XNOR U24356 ( .A(n24044), .B(n24043), .Z(n24045) );
  XOR U24357 ( .A(n24046), .B(n24045), .Z(n24054) );
  AND U24358 ( .A(y[2042]), .B(x[229]), .Z(n24048) );
  NAND U24359 ( .A(y[2040]), .B(x[231]), .Z(n24047) );
  XNOR U24360 ( .A(n24048), .B(n24047), .Z(n24052) );
  AND U24361 ( .A(y[2045]), .B(x[226]), .Z(n24050) );
  NAND U24362 ( .A(y[2030]), .B(x[241]), .Z(n24049) );
  XNOR U24363 ( .A(n24050), .B(n24049), .Z(n24051) );
  XNOR U24364 ( .A(n24052), .B(n24051), .Z(n24053) );
  XNOR U24365 ( .A(n24054), .B(n24053), .Z(n24055) );
  XNOR U24366 ( .A(n24056), .B(n24055), .Z(n24057) );
  XNOR U24367 ( .A(n24058), .B(n24057), .Z(n24059) );
  XNOR U24368 ( .A(n24060), .B(n24059), .Z(n24061) );
  XNOR U24369 ( .A(n24062), .B(n24061), .Z(n24063) );
  XNOR U24370 ( .A(n24064), .B(n24063), .Z(n24065) );
  XNOR U24371 ( .A(n24066), .B(n24065), .Z(n24082) );
  NAND U24372 ( .A(n24068), .B(n24067), .Z(n24072) );
  NAND U24373 ( .A(n24070), .B(n24069), .Z(n24071) );
  AND U24374 ( .A(n24072), .B(n24071), .Z(n24080) );
  NAND U24375 ( .A(n24074), .B(n24073), .Z(n24078) );
  NAND U24376 ( .A(n24076), .B(n24075), .Z(n24077) );
  NAND U24377 ( .A(n24078), .B(n24077), .Z(n24079) );
  XNOR U24378 ( .A(n24080), .B(n24079), .Z(n24081) );
  XNOR U24379 ( .A(n24082), .B(n24081), .Z(n24083) );
  XNOR U24380 ( .A(n24084), .B(n24083), .Z(n24085) );
  XNOR U24381 ( .A(n24086), .B(n24085), .Z(n24087) );
  XNOR U24382 ( .A(n24088), .B(n24087), .Z(n24104) );
  NAND U24383 ( .A(n24090), .B(n24089), .Z(n24094) );
  NANDN U24384 ( .A(n24092), .B(n24091), .Z(n24093) );
  AND U24385 ( .A(n24094), .B(n24093), .Z(n24102) );
  NANDN U24386 ( .A(n24096), .B(n24095), .Z(n24100) );
  NAND U24387 ( .A(n24098), .B(n24097), .Z(n24099) );
  NAND U24388 ( .A(n24100), .B(n24099), .Z(n24101) );
  XNOR U24389 ( .A(n24102), .B(n24101), .Z(n24103) );
  XNOR U24390 ( .A(n24104), .B(n24103), .Z(n24105) );
  XNOR U24391 ( .A(n24106), .B(n24105), .Z(n24122) );
  NANDN U24392 ( .A(n24108), .B(n24107), .Z(n24112) );
  NANDN U24393 ( .A(n24110), .B(n24109), .Z(n24111) );
  AND U24394 ( .A(n24112), .B(n24111), .Z(n24120) );
  NAND U24395 ( .A(n24114), .B(n24113), .Z(n24118) );
  NAND U24396 ( .A(n24116), .B(n24115), .Z(n24117) );
  NAND U24397 ( .A(n24118), .B(n24117), .Z(n24119) );
  XNOR U24398 ( .A(n24120), .B(n24119), .Z(n24121) );
  XNOR U24399 ( .A(n24122), .B(n24121), .Z(n24123) );
  XNOR U24400 ( .A(n24124), .B(n24123), .Z(n24140) );
  NANDN U24401 ( .A(n24126), .B(n24125), .Z(n24130) );
  NAND U24402 ( .A(n24128), .B(n24127), .Z(n24129) );
  AND U24403 ( .A(n24130), .B(n24129), .Z(n24138) );
  NANDN U24404 ( .A(n24132), .B(n24131), .Z(n24136) );
  NANDN U24405 ( .A(n24134), .B(n24133), .Z(n24135) );
  NAND U24406 ( .A(n24136), .B(n24135), .Z(n24137) );
  XNOR U24407 ( .A(n24138), .B(n24137), .Z(n24139) );
  XNOR U24408 ( .A(n24140), .B(n24139), .Z(n24141) );
  XNOR U24409 ( .A(n24142), .B(n24141), .Z(n24158) );
  NAND U24410 ( .A(n24144), .B(n24143), .Z(n24148) );
  NANDN U24411 ( .A(n24146), .B(n24145), .Z(n24147) );
  AND U24412 ( .A(n24148), .B(n24147), .Z(n24156) );
  NAND U24413 ( .A(n24150), .B(n24149), .Z(n24154) );
  NAND U24414 ( .A(n24152), .B(n24151), .Z(n24153) );
  NAND U24415 ( .A(n24154), .B(n24153), .Z(n24155) );
  XNOR U24416 ( .A(n24156), .B(n24155), .Z(n24157) );
  XNOR U24417 ( .A(n24158), .B(n24157), .Z(n24159) );
  XNOR U24418 ( .A(n24160), .B(n24159), .Z(N512) );
endmodule

