
module mult_N128_CC16 ( clk, rst, a, b, c );
  input [127:0] a;
  input [7:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320;
  wire   [255:0] sreg;

  DFF \sreg_reg[247]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[122]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[121]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[120]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[119]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NANDN U11 ( .A(b[0]), .B(a[127]), .Z(n1) );
  NAND U12 ( .A(b[1]), .B(n1), .Z(n5141) );
  XNOR U13 ( .A(n5145), .B(n5144), .Z(n5146) );
  XNOR U14 ( .A(n5170), .B(b[1]), .Z(n5172) );
  NAND U15 ( .A(n83), .B(n82), .Z(n2) );
  NANDN U16 ( .A(n85), .B(n84), .Z(n3) );
  AND U17 ( .A(n2), .B(n3), .Z(n106) );
  XNOR U18 ( .A(n5053), .B(n5052), .Z(n5055) );
  XNOR U19 ( .A(n5099), .B(n5098), .Z(n5100) );
  XNOR U20 ( .A(n5114), .B(n5113), .Z(n5115) );
  XNOR U21 ( .A(n5147), .B(n5146), .Z(n5150) );
  XNOR U22 ( .A(n5165), .B(n5164), .Z(n5166) );
  XNOR U23 ( .A(n5201), .B(n5200), .Z(n5202) );
  XNOR U24 ( .A(n5235), .B(n5234), .Z(n5237) );
  XNOR U25 ( .A(n5270), .B(n5269), .Z(n5279) );
  XOR U26 ( .A(n67), .B(n65), .Z(n4) );
  NANDN U27 ( .A(n66), .B(n4), .Z(n5) );
  NAND U28 ( .A(n67), .B(n65), .Z(n6) );
  AND U29 ( .A(n5), .B(n6), .Z(n85) );
  XNOR U30 ( .A(n5299), .B(n5298), .Z(n5300) );
  XNOR U31 ( .A(n5059), .B(n5058), .Z(n5060) );
  XNOR U32 ( .A(n5093), .B(n5092), .Z(n5094) );
  XNOR U33 ( .A(n5139), .B(n5138), .Z(n5140) );
  XNOR U34 ( .A(n5207), .B(n5206), .Z(n5208) );
  XNOR U35 ( .A(n5049), .B(n5048), .Z(n5040) );
  XNOR U36 ( .A(n5151), .B(n5150), .Z(n5152) );
  XNOR U37 ( .A(n5255), .B(n5254), .Z(n5256) );
  XNOR U38 ( .A(n5087), .B(n5086), .Z(n5088) );
  XNOR U39 ( .A(n5167), .B(n5166), .Z(n5158) );
  XNOR U40 ( .A(n5203), .B(n5202), .Z(n5194) );
  XNOR U41 ( .A(n5280), .B(n5279), .Z(n5281) );
  XOR U42 ( .A(n5301), .B(n5300), .Z(n5304) );
  NAND U43 ( .A(sreg[123]), .B(n78), .Z(n7) );
  XOR U44 ( .A(sreg[123]), .B(n78), .Z(n8) );
  NANDN U45 ( .A(n77), .B(n8), .Z(n9) );
  NAND U46 ( .A(n7), .B(n9), .Z(n80) );
  XOR U47 ( .A(n133), .B(sreg[126]), .Z(n10) );
  NANDN U48 ( .A(n134), .B(n10), .Z(n11) );
  NAND U49 ( .A(n133), .B(sreg[126]), .Z(n12) );
  AND U50 ( .A(n11), .B(n12), .Z(n169) );
  XOR U51 ( .A(n5318), .B(n5319), .Z(n5314) );
  XNOR U52 ( .A(n5141), .B(n5140), .Z(n5144) );
  XOR U53 ( .A(n5189), .B(n5188), .Z(n5171) );
  XNOR U54 ( .A(n5221), .B(n5220), .Z(n5222) );
  XNOR U55 ( .A(n5047), .B(n5046), .Z(n5048) );
  XNOR U56 ( .A(n5095), .B(n5094), .Z(n5113) );
  XOR U57 ( .A(n5153), .B(n5152), .Z(n5121) );
  XOR U58 ( .A(n5282), .B(n5281), .Z(n5263) );
  XNOR U59 ( .A(n5089), .B(n5088), .Z(n5081) );
  XNOR U60 ( .A(n5159), .B(n5158), .Z(n5160) );
  XNOR U61 ( .A(n5195), .B(n5194), .Z(n5196) );
  XNOR U62 ( .A(n5229), .B(n5228), .Z(n5230) );
  XOR U63 ( .A(sreg[124]), .B(n80), .Z(n13) );
  NANDN U64 ( .A(n81), .B(n13), .Z(n14) );
  NAND U65 ( .A(sreg[124]), .B(n80), .Z(n15) );
  AND U66 ( .A(n14), .B(n15), .Z(n129) );
  NAND U67 ( .A(sreg[128]), .B(n206), .Z(n16) );
  XOR U68 ( .A(sreg[128]), .B(n206), .Z(n17) );
  NANDN U69 ( .A(n205), .B(n17), .Z(n18) );
  NAND U70 ( .A(n16), .B(n18), .Z(n281) );
  XNOR U71 ( .A(n5313), .B(n5314), .Z(n19) );
  XNOR U72 ( .A(n5312), .B(n19), .Z(n20) );
  NAND U73 ( .A(n5315), .B(n20), .Z(n21) );
  NANDN U74 ( .A(n5313), .B(n5314), .Z(n22) );
  NAND U75 ( .A(n5312), .B(n19), .Z(n23) );
  NAND U76 ( .A(n22), .B(n23), .Z(n24) );
  NAND U77 ( .A(n21), .B(n24), .Z(n25) );
  NAND U78 ( .A(n5317), .B(n5316), .Z(n26) );
  NANDN U79 ( .A(n5318), .B(n5319), .Z(n27) );
  AND U80 ( .A(n26), .B(n27), .Z(n28) );
  XNOR U81 ( .A(a[127]), .B(a[126]), .Z(n29) );
  XNOR U82 ( .A(n5320), .B(n29), .Z(n30) );
  AND U83 ( .A(n30), .B(b[7]), .Z(n31) );
  XNOR U84 ( .A(n25), .B(n28), .Z(n32) );
  XNOR U85 ( .A(n31), .B(n32), .Z(c[255]) );
  AND U86 ( .A(b[0]), .B(a[0]), .Z(n34) );
  XOR U87 ( .A(n34), .B(sreg[120]), .Z(c[120]) );
  AND U88 ( .A(b[0]), .B(a[1]), .Z(n44) );
  NAND U89 ( .A(a[0]), .B(b[1]), .Z(n33) );
  XOR U90 ( .A(n44), .B(n33), .Z(n35) );
  XNOR U91 ( .A(sreg[121]), .B(n35), .Z(n37) );
  AND U92 ( .A(n34), .B(sreg[120]), .Z(n36) );
  XOR U93 ( .A(n37), .B(n36), .Z(c[121]) );
  NANDN U94 ( .A(n35), .B(sreg[121]), .Z(n39) );
  NAND U95 ( .A(n37), .B(n36), .Z(n38) );
  AND U96 ( .A(n39), .B(n38), .Z(n47) );
  XNOR U97 ( .A(n47), .B(sreg[122]), .Z(n49) );
  NAND U98 ( .A(b[0]), .B(a[2]), .Z(n40) );
  XNOR U99 ( .A(b[1]), .B(n40), .Z(n42) );
  NANDN U100 ( .A(b[0]), .B(a[1]), .Z(n41) );
  NAND U101 ( .A(n42), .B(n41), .Z(n53) );
  NAND U102 ( .A(a[0]), .B(b[2]), .Z(n43) );
  XNOR U103 ( .A(b[1]), .B(n43), .Z(n46) );
  NANDN U104 ( .A(a[0]), .B(n44), .Z(n45) );
  NAND U105 ( .A(n46), .B(n45), .Z(n52) );
  XOR U106 ( .A(n53), .B(n52), .Z(n48) );
  XOR U107 ( .A(n49), .B(n48), .Z(c[122]) );
  NANDN U108 ( .A(n47), .B(sreg[122]), .Z(n51) );
  NAND U109 ( .A(n49), .B(n48), .Z(n50) );
  NAND U110 ( .A(n51), .B(n50), .Z(n78) );
  NOR U111 ( .A(n53), .B(n52), .Z(n67) );
  NAND U112 ( .A(b[0]), .B(a[3]), .Z(n54) );
  XNOR U113 ( .A(b[1]), .B(n54), .Z(n56) );
  NANDN U114 ( .A(b[0]), .B(a[2]), .Z(n55) );
  NAND U115 ( .A(n56), .B(n55), .Z(n75) );
  XOR U116 ( .A(b[3]), .B(b[2]), .Z(n68) );
  XOR U117 ( .A(b[3]), .B(a[0]), .Z(n57) );
  NAND U118 ( .A(n68), .B(n57), .Z(n58) );
  XOR U119 ( .A(b[1]), .B(b[2]), .Z(n5135) );
  OR U120 ( .A(n58), .B(n5135), .Z(n60) );
  XOR U121 ( .A(b[3]), .B(a[1]), .Z(n69) );
  NAND U122 ( .A(n5135), .B(n69), .Z(n59) );
  AND U123 ( .A(n60), .B(n59), .Z(n76) );
  XNOR U124 ( .A(n75), .B(n76), .Z(n66) );
  IV U125 ( .A(n5135), .Z(n5177) );
  NANDN U126 ( .A(n5177), .B(a[0]), .Z(n62) );
  NAND U127 ( .A(b[1]), .B(b[2]), .Z(n61) );
  AND U128 ( .A(b[3]), .B(n61), .Z(n5241) );
  IV U129 ( .A(n5241), .Z(n5219) );
  ANDN U130 ( .B(n62), .A(n5219), .Z(n65) );
  XOR U131 ( .A(n66), .B(n65), .Z(n63) );
  XOR U132 ( .A(n67), .B(n63), .Z(n77) );
  XOR U133 ( .A(sreg[123]), .B(n77), .Z(n64) );
  XNOR U134 ( .A(n78), .B(n64), .Z(c[123]) );
  ANDN U135 ( .B(n68), .A(n5135), .Z(n5134) );
  IV U136 ( .A(n5134), .Z(n5176) );
  NANDN U137 ( .A(n5176), .B(n69), .Z(n71) );
  XOR U138 ( .A(b[3]), .B(a[2]), .Z(n86) );
  NANDN U139 ( .A(n5177), .B(n86), .Z(n70) );
  AND U140 ( .A(n71), .B(n70), .Z(n100) );
  XOR U141 ( .A(b[4]), .B(b[3]), .Z(n5251) );
  IV U142 ( .A(n5251), .Z(n5184) );
  ANDN U143 ( .B(a[0]), .A(n5184), .Z(n97) );
  NAND U144 ( .A(b[0]), .B(a[4]), .Z(n72) );
  XNOR U145 ( .A(b[1]), .B(n72), .Z(n74) );
  NANDN U146 ( .A(b[0]), .B(a[3]), .Z(n73) );
  NAND U147 ( .A(n74), .B(n73), .Z(n98) );
  XNOR U148 ( .A(n97), .B(n98), .Z(n99) );
  XNOR U149 ( .A(n100), .B(n99), .Z(n83) );
  NOR U150 ( .A(n76), .B(n75), .Z(n82) );
  XOR U151 ( .A(n83), .B(n82), .Z(n84) );
  XOR U152 ( .A(n85), .B(n84), .Z(n81) );
  XOR U153 ( .A(n80), .B(sreg[124]), .Z(n79) );
  XNOR U154 ( .A(n81), .B(n79), .Z(c[124]) );
  NANDN U155 ( .A(n5176), .B(n86), .Z(n88) );
  XOR U156 ( .A(b[3]), .B(a[3]), .Z(n115) );
  NANDN U157 ( .A(n5177), .B(n115), .Z(n87) );
  AND U158 ( .A(n88), .B(n87), .Z(n122) );
  NAND U159 ( .A(b[3]), .B(b[4]), .Z(n89) );
  AND U160 ( .A(b[5]), .B(n89), .Z(n5285) );
  ANDN U161 ( .B(n5285), .A(n97), .Z(n121) );
  XNOR U162 ( .A(n122), .B(n121), .Z(n124) );
  XOR U163 ( .A(b[5]), .B(b[4]), .Z(n109) );
  XOR U164 ( .A(b[5]), .B(a[0]), .Z(n90) );
  NAND U165 ( .A(n109), .B(n90), .Z(n91) );
  OR U166 ( .A(n91), .B(n5251), .Z(n93) );
  XOR U167 ( .A(b[5]), .B(a[1]), .Z(n110) );
  NAND U168 ( .A(n5251), .B(n110), .Z(n92) );
  NAND U169 ( .A(n93), .B(n92), .Z(n114) );
  NAND U170 ( .A(b[0]), .B(a[5]), .Z(n94) );
  XNOR U171 ( .A(b[1]), .B(n94), .Z(n96) );
  NANDN U172 ( .A(b[0]), .B(a[4]), .Z(n95) );
  NAND U173 ( .A(n96), .B(n95), .Z(n113) );
  XNOR U174 ( .A(n114), .B(n113), .Z(n123) );
  XOR U175 ( .A(n124), .B(n123), .Z(n104) );
  NANDN U176 ( .A(n98), .B(n97), .Z(n102) );
  NANDN U177 ( .A(n100), .B(n99), .Z(n101) );
  AND U178 ( .A(n102), .B(n101), .Z(n103) );
  XNOR U179 ( .A(n104), .B(n103), .Z(n105) );
  XOR U180 ( .A(n106), .B(n105), .Z(n127) );
  XNOR U181 ( .A(n127), .B(sreg[125]), .Z(n128) );
  XNOR U182 ( .A(n129), .B(n128), .Z(c[125]) );
  NANDN U183 ( .A(n104), .B(n103), .Z(n108) );
  NAND U184 ( .A(n106), .B(n105), .Z(n107) );
  AND U185 ( .A(n108), .B(n107), .Z(n138) );
  ANDN U186 ( .B(n109), .A(n5251), .Z(n5216) );
  IV U187 ( .A(n5216), .Z(n5249) );
  NANDN U188 ( .A(n5249), .B(n110), .Z(n112) );
  XOR U189 ( .A(b[5]), .B(a[2]), .Z(n141) );
  NANDN U190 ( .A(n5184), .B(n141), .Z(n111) );
  AND U191 ( .A(n112), .B(n111), .Z(n162) );
  ANDN U192 ( .B(n114), .A(n113), .Z(n161) );
  XNOR U193 ( .A(n162), .B(n161), .Z(n164) );
  NANDN U194 ( .A(n5176), .B(n115), .Z(n117) );
  XOR U195 ( .A(b[3]), .B(a[4]), .Z(n152) );
  NANDN U196 ( .A(n5177), .B(n152), .Z(n116) );
  AND U197 ( .A(n117), .B(n116), .Z(n158) );
  XOR U198 ( .A(b[5]), .B(b[6]), .Z(n5291) );
  IV U199 ( .A(n5291), .Z(n5275) );
  ANDN U200 ( .B(a[0]), .A(n5275), .Z(n155) );
  NAND U201 ( .A(b[0]), .B(a[6]), .Z(n118) );
  XNOR U202 ( .A(b[1]), .B(n118), .Z(n120) );
  NANDN U203 ( .A(b[0]), .B(a[5]), .Z(n119) );
  NAND U204 ( .A(n120), .B(n119), .Z(n156) );
  XNOR U205 ( .A(n155), .B(n156), .Z(n157) );
  XNOR U206 ( .A(n158), .B(n157), .Z(n163) );
  XOR U207 ( .A(n164), .B(n163), .Z(n136) );
  NANDN U208 ( .A(n122), .B(n121), .Z(n126) );
  NAND U209 ( .A(n124), .B(n123), .Z(n125) );
  AND U210 ( .A(n126), .B(n125), .Z(n135) );
  XNOR U211 ( .A(n136), .B(n135), .Z(n137) );
  XNOR U212 ( .A(n138), .B(n137), .Z(n134) );
  NANDN U213 ( .A(n127), .B(sreg[125]), .Z(n131) );
  NANDN U214 ( .A(n129), .B(n128), .Z(n130) );
  NAND U215 ( .A(n131), .B(n130), .Z(n133) );
  XOR U216 ( .A(n133), .B(sreg[126]), .Z(n132) );
  XNOR U217 ( .A(n134), .B(n132), .Z(c[126]) );
  NANDN U218 ( .A(n136), .B(n135), .Z(n140) );
  NANDN U219 ( .A(n138), .B(n137), .Z(n139) );
  AND U220 ( .A(n140), .B(n139), .Z(n200) );
  NANDN U221 ( .A(n5249), .B(n141), .Z(n143) );
  XOR U222 ( .A(b[5]), .B(a[3]), .Z(n189) );
  NANDN U223 ( .A(n5184), .B(n189), .Z(n142) );
  AND U224 ( .A(n143), .B(n142), .Z(n179) );
  XOR U225 ( .A(b[6]), .B(b[7]), .Z(n144) );
  ANDN U226 ( .B(n144), .A(n5291), .Z(n5293) );
  IV U227 ( .A(n5293), .Z(n5274) );
  XOR U228 ( .A(a[0]), .B(b[7]), .Z(n145) );
  NANDN U229 ( .A(n5274), .B(n145), .Z(n147) );
  XOR U230 ( .A(b[7]), .B(a[1]), .Z(n180) );
  ANDN U231 ( .B(n180), .A(n5275), .Z(n146) );
  ANDN U232 ( .B(n147), .A(n146), .Z(n178) );
  XOR U233 ( .A(n179), .B(n178), .Z(n195) );
  NAND U234 ( .A(b[5]), .B(b[6]), .Z(n5320) );
  AND U235 ( .A(b[7]), .B(n5320), .Z(n148) );
  ANDN U236 ( .B(n148), .A(n155), .Z(n193) );
  NAND U237 ( .A(b[0]), .B(a[7]), .Z(n149) );
  XNOR U238 ( .A(b[1]), .B(n149), .Z(n151) );
  NANDN U239 ( .A(b[0]), .B(a[6]), .Z(n150) );
  NAND U240 ( .A(n151), .B(n150), .Z(n192) );
  XNOR U241 ( .A(n193), .B(n192), .Z(n194) );
  XNOR U242 ( .A(n195), .B(n194), .Z(n172) );
  NAND U243 ( .A(n5134), .B(n152), .Z(n154) );
  XNOR U244 ( .A(b[3]), .B(a[5]), .Z(n183) );
  NANDN U245 ( .A(n183), .B(n5135), .Z(n153) );
  NAND U246 ( .A(n154), .B(n153), .Z(n173) );
  XNOR U247 ( .A(n172), .B(n173), .Z(n174) );
  NANDN U248 ( .A(n156), .B(n155), .Z(n160) );
  NANDN U249 ( .A(n158), .B(n157), .Z(n159) );
  NAND U250 ( .A(n160), .B(n159), .Z(n175) );
  XNOR U251 ( .A(n174), .B(n175), .Z(n198) );
  NANDN U252 ( .A(n162), .B(n161), .Z(n166) );
  NAND U253 ( .A(n164), .B(n163), .Z(n165) );
  NAND U254 ( .A(n166), .B(n165), .Z(n199) );
  XOR U255 ( .A(n198), .B(n199), .Z(n201) );
  XOR U256 ( .A(n200), .B(n201), .Z(n167) );
  XNOR U257 ( .A(n167), .B(sreg[127]), .Z(n168) );
  XNOR U258 ( .A(n169), .B(n168), .Z(c[127]) );
  NANDN U259 ( .A(n167), .B(sreg[127]), .Z(n171) );
  NANDN U260 ( .A(n169), .B(n168), .Z(n170) );
  AND U261 ( .A(n171), .B(n170), .Z(n205) );
  NANDN U262 ( .A(n173), .B(n172), .Z(n177) );
  NANDN U263 ( .A(n175), .B(n174), .Z(n176) );
  AND U264 ( .A(n177), .B(n176), .Z(n237) );
  NOR U265 ( .A(n179), .B(n178), .Z(n227) );
  NAND U266 ( .A(n5293), .B(n180), .Z(n182) );
  XNOR U267 ( .A(b[7]), .B(a[2]), .Z(n213) );
  NANDN U268 ( .A(n213), .B(n5291), .Z(n181) );
  AND U269 ( .A(n182), .B(n181), .Z(n225) );
  NANDN U270 ( .A(n183), .B(n5134), .Z(n185) );
  XNOR U271 ( .A(b[3]), .B(a[6]), .Z(n216) );
  NANDN U272 ( .A(n216), .B(n5135), .Z(n184) );
  NAND U273 ( .A(n185), .B(n184), .Z(n226) );
  XOR U274 ( .A(n225), .B(n226), .Z(n228) );
  XOR U275 ( .A(n227), .B(n228), .Z(n232) );
  NAND U276 ( .A(b[0]), .B(a[8]), .Z(n186) );
  XNOR U277 ( .A(b[1]), .B(n186), .Z(n188) );
  NANDN U278 ( .A(b[0]), .B(a[7]), .Z(n187) );
  NAND U279 ( .A(n188), .B(n187), .Z(n210) );
  NANDN U280 ( .A(n5249), .B(n189), .Z(n191) );
  XOR U281 ( .A(b[5]), .B(a[4]), .Z(n222) );
  NANDN U282 ( .A(n5184), .B(n222), .Z(n190) );
  AND U283 ( .A(n191), .B(n190), .Z(n208) );
  AND U284 ( .A(b[7]), .B(a[0]), .Z(n207) );
  XNOR U285 ( .A(n208), .B(n207), .Z(n209) );
  XNOR U286 ( .A(n210), .B(n209), .Z(n231) );
  XNOR U287 ( .A(n232), .B(n231), .Z(n233) );
  NANDN U288 ( .A(n193), .B(n192), .Z(n197) );
  NANDN U289 ( .A(n195), .B(n194), .Z(n196) );
  NAND U290 ( .A(n197), .B(n196), .Z(n234) );
  XOR U291 ( .A(n233), .B(n234), .Z(n238) );
  XNOR U292 ( .A(n237), .B(n238), .Z(n239) );
  NANDN U293 ( .A(n199), .B(n198), .Z(n203) );
  OR U294 ( .A(n201), .B(n200), .Z(n202) );
  NAND U295 ( .A(n203), .B(n202), .Z(n240) );
  XNOR U296 ( .A(n239), .B(n240), .Z(n206) );
  XNOR U297 ( .A(sreg[128]), .B(n206), .Z(n204) );
  XOR U298 ( .A(n205), .B(n204), .Z(c[128]) );
  NANDN U299 ( .A(n208), .B(n207), .Z(n212) );
  NANDN U300 ( .A(n210), .B(n209), .Z(n211) );
  AND U301 ( .A(n212), .B(n211), .Z(n274) );
  NANDN U302 ( .A(n213), .B(n5293), .Z(n215) );
  XOR U303 ( .A(b[7]), .B(a[3]), .Z(n249) );
  NANDN U304 ( .A(n5275), .B(n249), .Z(n214) );
  AND U305 ( .A(n215), .B(n214), .Z(n268) );
  NANDN U306 ( .A(n216), .B(n5134), .Z(n218) );
  XOR U307 ( .A(b[3]), .B(a[7]), .Z(n252) );
  NANDN U308 ( .A(n5177), .B(n252), .Z(n217) );
  NAND U309 ( .A(n218), .B(n217), .Z(n267) );
  XNOR U310 ( .A(n268), .B(n267), .Z(n269) );
  NAND U311 ( .A(b[0]), .B(a[9]), .Z(n219) );
  XNOR U312 ( .A(b[1]), .B(n219), .Z(n221) );
  NANDN U313 ( .A(b[0]), .B(a[8]), .Z(n220) );
  NAND U314 ( .A(n221), .B(n220), .Z(n264) );
  NANDN U315 ( .A(n5249), .B(n222), .Z(n224) );
  XOR U316 ( .A(b[5]), .B(a[5]), .Z(n258) );
  NANDN U317 ( .A(n5184), .B(n258), .Z(n223) );
  AND U318 ( .A(n224), .B(n223), .Z(n262) );
  AND U319 ( .A(b[7]), .B(a[1]), .Z(n261) );
  XNOR U320 ( .A(n262), .B(n261), .Z(n263) );
  XOR U321 ( .A(n264), .B(n263), .Z(n270) );
  XNOR U322 ( .A(n269), .B(n270), .Z(n273) );
  XNOR U323 ( .A(n274), .B(n273), .Z(n276) );
  NANDN U324 ( .A(n226), .B(n225), .Z(n230) );
  OR U325 ( .A(n228), .B(n227), .Z(n229) );
  AND U326 ( .A(n230), .B(n229), .Z(n275) );
  XOR U327 ( .A(n276), .B(n275), .Z(n244) );
  NANDN U328 ( .A(n232), .B(n231), .Z(n236) );
  NANDN U329 ( .A(n234), .B(n233), .Z(n235) );
  AND U330 ( .A(n236), .B(n235), .Z(n243) );
  XNOR U331 ( .A(n244), .B(n243), .Z(n246) );
  NANDN U332 ( .A(n238), .B(n237), .Z(n242) );
  NANDN U333 ( .A(n240), .B(n239), .Z(n241) );
  AND U334 ( .A(n242), .B(n241), .Z(n245) );
  XOR U335 ( .A(n246), .B(n245), .Z(n279) );
  XNOR U336 ( .A(n279), .B(sreg[129]), .Z(n280) );
  XOR U337 ( .A(n281), .B(n280), .Z(c[129]) );
  NANDN U338 ( .A(n244), .B(n243), .Z(n248) );
  NAND U339 ( .A(n246), .B(n245), .Z(n247) );
  AND U340 ( .A(n248), .B(n247), .Z(n291) );
  NANDN U341 ( .A(n5274), .B(n249), .Z(n251) );
  XOR U342 ( .A(b[7]), .B(a[4]), .Z(n301) );
  NANDN U343 ( .A(n5275), .B(n301), .Z(n250) );
  AND U344 ( .A(n251), .B(n250), .Z(n320) );
  NANDN U345 ( .A(n5176), .B(n252), .Z(n254) );
  XOR U346 ( .A(b[3]), .B(a[8]), .Z(n304) );
  NANDN U347 ( .A(n5177), .B(n304), .Z(n253) );
  NAND U348 ( .A(n254), .B(n253), .Z(n319) );
  XNOR U349 ( .A(n320), .B(n319), .Z(n322) );
  NAND U350 ( .A(b[0]), .B(a[10]), .Z(n255) );
  XNOR U351 ( .A(b[1]), .B(n255), .Z(n257) );
  NANDN U352 ( .A(b[0]), .B(a[9]), .Z(n256) );
  NAND U353 ( .A(n257), .B(n256), .Z(n316) );
  NANDN U354 ( .A(n5249), .B(n258), .Z(n260) );
  XOR U355 ( .A(b[5]), .B(a[6]), .Z(n310) );
  NANDN U356 ( .A(n5184), .B(n310), .Z(n259) );
  AND U357 ( .A(n260), .B(n259), .Z(n314) );
  AND U358 ( .A(b[7]), .B(a[2]), .Z(n313) );
  XNOR U359 ( .A(n314), .B(n313), .Z(n315) );
  XNOR U360 ( .A(n316), .B(n315), .Z(n321) );
  XOR U361 ( .A(n322), .B(n321), .Z(n296) );
  NANDN U362 ( .A(n262), .B(n261), .Z(n266) );
  NANDN U363 ( .A(n264), .B(n263), .Z(n265) );
  AND U364 ( .A(n266), .B(n265), .Z(n295) );
  XNOR U365 ( .A(n296), .B(n295), .Z(n297) );
  NANDN U366 ( .A(n268), .B(n267), .Z(n272) );
  NANDN U367 ( .A(n270), .B(n269), .Z(n271) );
  NAND U368 ( .A(n272), .B(n271), .Z(n298) );
  XNOR U369 ( .A(n297), .B(n298), .Z(n289) );
  NANDN U370 ( .A(n274), .B(n273), .Z(n278) );
  NAND U371 ( .A(n276), .B(n275), .Z(n277) );
  NAND U372 ( .A(n278), .B(n277), .Z(n290) );
  XOR U373 ( .A(n289), .B(n290), .Z(n292) );
  XOR U374 ( .A(n291), .B(n292), .Z(n284) );
  XNOR U375 ( .A(n284), .B(sreg[130]), .Z(n286) );
  NANDN U376 ( .A(n279), .B(sreg[129]), .Z(n283) );
  NAND U377 ( .A(n281), .B(n280), .Z(n282) );
  NAND U378 ( .A(n283), .B(n282), .Z(n285) );
  XOR U379 ( .A(n286), .B(n285), .Z(c[130]) );
  NANDN U380 ( .A(n284), .B(sreg[130]), .Z(n288) );
  NAND U381 ( .A(n286), .B(n285), .Z(n287) );
  AND U382 ( .A(n288), .B(n287), .Z(n363) );
  NANDN U383 ( .A(n290), .B(n289), .Z(n294) );
  OR U384 ( .A(n292), .B(n291), .Z(n293) );
  AND U385 ( .A(n294), .B(n293), .Z(n328) );
  NANDN U386 ( .A(n296), .B(n295), .Z(n300) );
  NANDN U387 ( .A(n298), .B(n297), .Z(n299) );
  AND U388 ( .A(n300), .B(n299), .Z(n326) );
  NANDN U389 ( .A(n5274), .B(n301), .Z(n303) );
  XOR U390 ( .A(b[7]), .B(a[5]), .Z(n337) );
  NANDN U391 ( .A(n5275), .B(n337), .Z(n302) );
  AND U392 ( .A(n303), .B(n302), .Z(n356) );
  NANDN U393 ( .A(n5176), .B(n304), .Z(n306) );
  XOR U394 ( .A(b[3]), .B(a[9]), .Z(n340) );
  NANDN U395 ( .A(n5177), .B(n340), .Z(n305) );
  NAND U396 ( .A(n306), .B(n305), .Z(n355) );
  XNOR U397 ( .A(n356), .B(n355), .Z(n358) );
  NAND U398 ( .A(b[0]), .B(a[11]), .Z(n307) );
  XNOR U399 ( .A(b[1]), .B(n307), .Z(n309) );
  NANDN U400 ( .A(b[0]), .B(a[10]), .Z(n308) );
  NAND U401 ( .A(n309), .B(n308), .Z(n352) );
  NANDN U402 ( .A(n5249), .B(n310), .Z(n312) );
  XOR U403 ( .A(b[5]), .B(a[7]), .Z(n346) );
  NANDN U404 ( .A(n5184), .B(n346), .Z(n311) );
  AND U405 ( .A(n312), .B(n311), .Z(n350) );
  AND U406 ( .A(b[7]), .B(a[3]), .Z(n349) );
  XNOR U407 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U408 ( .A(n352), .B(n351), .Z(n357) );
  XOR U409 ( .A(n358), .B(n357), .Z(n332) );
  NANDN U410 ( .A(n314), .B(n313), .Z(n318) );
  NANDN U411 ( .A(n316), .B(n315), .Z(n317) );
  AND U412 ( .A(n318), .B(n317), .Z(n331) );
  XNOR U413 ( .A(n332), .B(n331), .Z(n333) );
  NANDN U414 ( .A(n320), .B(n319), .Z(n324) );
  NAND U415 ( .A(n322), .B(n321), .Z(n323) );
  NAND U416 ( .A(n324), .B(n323), .Z(n334) );
  XNOR U417 ( .A(n333), .B(n334), .Z(n325) );
  XNOR U418 ( .A(n326), .B(n325), .Z(n327) );
  XNOR U419 ( .A(n328), .B(n327), .Z(n361) );
  XNOR U420 ( .A(sreg[131]), .B(n361), .Z(n362) );
  XNOR U421 ( .A(n363), .B(n362), .Z(c[131]) );
  NANDN U422 ( .A(n326), .B(n325), .Z(n330) );
  NANDN U423 ( .A(n328), .B(n327), .Z(n329) );
  AND U424 ( .A(n330), .B(n329), .Z(n373) );
  NANDN U425 ( .A(n332), .B(n331), .Z(n336) );
  NANDN U426 ( .A(n334), .B(n333), .Z(n335) );
  AND U427 ( .A(n336), .B(n335), .Z(n372) );
  NANDN U428 ( .A(n5274), .B(n337), .Z(n339) );
  XOR U429 ( .A(b[7]), .B(a[6]), .Z(n383) );
  NANDN U430 ( .A(n5275), .B(n383), .Z(n338) );
  AND U431 ( .A(n339), .B(n338), .Z(n402) );
  NANDN U432 ( .A(n5176), .B(n340), .Z(n342) );
  XOR U433 ( .A(b[3]), .B(a[10]), .Z(n386) );
  NANDN U434 ( .A(n5177), .B(n386), .Z(n341) );
  NAND U435 ( .A(n342), .B(n341), .Z(n401) );
  XNOR U436 ( .A(n402), .B(n401), .Z(n404) );
  NAND U437 ( .A(b[0]), .B(a[12]), .Z(n343) );
  XNOR U438 ( .A(b[1]), .B(n343), .Z(n345) );
  NANDN U439 ( .A(b[0]), .B(a[11]), .Z(n344) );
  NAND U440 ( .A(n345), .B(n344), .Z(n398) );
  NANDN U441 ( .A(n5249), .B(n346), .Z(n348) );
  XOR U442 ( .A(b[5]), .B(a[8]), .Z(n389) );
  NANDN U443 ( .A(n5184), .B(n389), .Z(n347) );
  AND U444 ( .A(n348), .B(n347), .Z(n396) );
  AND U445 ( .A(b[7]), .B(a[4]), .Z(n395) );
  XNOR U446 ( .A(n396), .B(n395), .Z(n397) );
  XNOR U447 ( .A(n398), .B(n397), .Z(n403) );
  XOR U448 ( .A(n404), .B(n403), .Z(n378) );
  NANDN U449 ( .A(n350), .B(n349), .Z(n354) );
  NANDN U450 ( .A(n352), .B(n351), .Z(n353) );
  AND U451 ( .A(n354), .B(n353), .Z(n377) );
  XNOR U452 ( .A(n378), .B(n377), .Z(n379) );
  NANDN U453 ( .A(n356), .B(n355), .Z(n360) );
  NAND U454 ( .A(n358), .B(n357), .Z(n359) );
  NAND U455 ( .A(n360), .B(n359), .Z(n380) );
  XNOR U456 ( .A(n379), .B(n380), .Z(n371) );
  XOR U457 ( .A(n372), .B(n371), .Z(n374) );
  XOR U458 ( .A(n373), .B(n374), .Z(n366) );
  XNOR U459 ( .A(n366), .B(sreg[132]), .Z(n368) );
  NANDN U460 ( .A(sreg[131]), .B(n361), .Z(n365) );
  NAND U461 ( .A(n363), .B(n362), .Z(n364) );
  AND U462 ( .A(n365), .B(n364), .Z(n367) );
  XOR U463 ( .A(n368), .B(n367), .Z(c[132]) );
  NANDN U464 ( .A(n366), .B(sreg[132]), .Z(n370) );
  NAND U465 ( .A(n368), .B(n367), .Z(n369) );
  AND U466 ( .A(n370), .B(n369), .Z(n445) );
  NANDN U467 ( .A(n372), .B(n371), .Z(n376) );
  OR U468 ( .A(n374), .B(n373), .Z(n375) );
  AND U469 ( .A(n376), .B(n375), .Z(n410) );
  NANDN U470 ( .A(n378), .B(n377), .Z(n382) );
  NANDN U471 ( .A(n380), .B(n379), .Z(n381) );
  AND U472 ( .A(n382), .B(n381), .Z(n408) );
  NANDN U473 ( .A(n5274), .B(n383), .Z(n385) );
  XOR U474 ( .A(b[7]), .B(a[7]), .Z(n419) );
  NANDN U475 ( .A(n5275), .B(n419), .Z(n384) );
  AND U476 ( .A(n385), .B(n384), .Z(n438) );
  NANDN U477 ( .A(n5176), .B(n386), .Z(n388) );
  XOR U478 ( .A(b[3]), .B(a[11]), .Z(n422) );
  NANDN U479 ( .A(n5177), .B(n422), .Z(n387) );
  NAND U480 ( .A(n388), .B(n387), .Z(n437) );
  XNOR U481 ( .A(n438), .B(n437), .Z(n440) );
  NANDN U482 ( .A(n5249), .B(n389), .Z(n391) );
  XOR U483 ( .A(b[5]), .B(a[9]), .Z(n428) );
  NANDN U484 ( .A(n5184), .B(n428), .Z(n390) );
  AND U485 ( .A(n391), .B(n390), .Z(n432) );
  AND U486 ( .A(b[7]), .B(a[5]), .Z(n431) );
  XNOR U487 ( .A(n432), .B(n431), .Z(n433) );
  NAND U488 ( .A(b[0]), .B(a[13]), .Z(n392) );
  XNOR U489 ( .A(b[1]), .B(n392), .Z(n394) );
  NANDN U490 ( .A(b[0]), .B(a[12]), .Z(n393) );
  NAND U491 ( .A(n394), .B(n393), .Z(n434) );
  XNOR U492 ( .A(n433), .B(n434), .Z(n439) );
  XOR U493 ( .A(n440), .B(n439), .Z(n414) );
  NANDN U494 ( .A(n396), .B(n395), .Z(n400) );
  NANDN U495 ( .A(n398), .B(n397), .Z(n399) );
  AND U496 ( .A(n400), .B(n399), .Z(n413) );
  XNOR U497 ( .A(n414), .B(n413), .Z(n415) );
  NANDN U498 ( .A(n402), .B(n401), .Z(n406) );
  NAND U499 ( .A(n404), .B(n403), .Z(n405) );
  NAND U500 ( .A(n406), .B(n405), .Z(n416) );
  XNOR U501 ( .A(n415), .B(n416), .Z(n407) );
  XNOR U502 ( .A(n408), .B(n407), .Z(n409) );
  XNOR U503 ( .A(n410), .B(n409), .Z(n443) );
  XNOR U504 ( .A(sreg[133]), .B(n443), .Z(n444) );
  XNOR U505 ( .A(n445), .B(n444), .Z(c[133]) );
  NANDN U506 ( .A(n408), .B(n407), .Z(n412) );
  NANDN U507 ( .A(n410), .B(n409), .Z(n411) );
  AND U508 ( .A(n412), .B(n411), .Z(n451) );
  NANDN U509 ( .A(n414), .B(n413), .Z(n418) );
  NANDN U510 ( .A(n416), .B(n415), .Z(n417) );
  AND U511 ( .A(n418), .B(n417), .Z(n449) );
  NANDN U512 ( .A(n5274), .B(n419), .Z(n421) );
  XOR U513 ( .A(b[7]), .B(a[8]), .Z(n460) );
  NANDN U514 ( .A(n5275), .B(n460), .Z(n420) );
  AND U515 ( .A(n421), .B(n420), .Z(n479) );
  NANDN U516 ( .A(n5176), .B(n422), .Z(n424) );
  XOR U517 ( .A(b[3]), .B(a[12]), .Z(n463) );
  NANDN U518 ( .A(n5177), .B(n463), .Z(n423) );
  NAND U519 ( .A(n424), .B(n423), .Z(n478) );
  XNOR U520 ( .A(n479), .B(n478), .Z(n481) );
  NAND U521 ( .A(b[0]), .B(a[14]), .Z(n425) );
  XNOR U522 ( .A(b[1]), .B(n425), .Z(n427) );
  NANDN U523 ( .A(b[0]), .B(a[13]), .Z(n426) );
  NAND U524 ( .A(n427), .B(n426), .Z(n475) );
  NANDN U525 ( .A(n5249), .B(n428), .Z(n430) );
  XOR U526 ( .A(b[5]), .B(a[10]), .Z(n469) );
  NANDN U527 ( .A(n5184), .B(n469), .Z(n429) );
  AND U528 ( .A(n430), .B(n429), .Z(n473) );
  AND U529 ( .A(b[7]), .B(a[6]), .Z(n472) );
  XNOR U530 ( .A(n473), .B(n472), .Z(n474) );
  XNOR U531 ( .A(n475), .B(n474), .Z(n480) );
  XOR U532 ( .A(n481), .B(n480), .Z(n455) );
  NANDN U533 ( .A(n432), .B(n431), .Z(n436) );
  NANDN U534 ( .A(n434), .B(n433), .Z(n435) );
  AND U535 ( .A(n436), .B(n435), .Z(n454) );
  XNOR U536 ( .A(n455), .B(n454), .Z(n456) );
  NANDN U537 ( .A(n438), .B(n437), .Z(n442) );
  NAND U538 ( .A(n440), .B(n439), .Z(n441) );
  NAND U539 ( .A(n442), .B(n441), .Z(n457) );
  XNOR U540 ( .A(n456), .B(n457), .Z(n448) );
  XNOR U541 ( .A(n449), .B(n448), .Z(n450) );
  XNOR U542 ( .A(n451), .B(n450), .Z(n484) );
  XNOR U543 ( .A(sreg[134]), .B(n484), .Z(n486) );
  NANDN U544 ( .A(sreg[133]), .B(n443), .Z(n447) );
  NAND U545 ( .A(n445), .B(n444), .Z(n446) );
  NAND U546 ( .A(n447), .B(n446), .Z(n485) );
  XNOR U547 ( .A(n486), .B(n485), .Z(c[134]) );
  NANDN U548 ( .A(n449), .B(n448), .Z(n453) );
  NANDN U549 ( .A(n451), .B(n450), .Z(n452) );
  AND U550 ( .A(n453), .B(n452), .Z(n492) );
  NANDN U551 ( .A(n455), .B(n454), .Z(n459) );
  NANDN U552 ( .A(n457), .B(n456), .Z(n458) );
  AND U553 ( .A(n459), .B(n458), .Z(n490) );
  NANDN U554 ( .A(n5274), .B(n460), .Z(n462) );
  XOR U555 ( .A(b[7]), .B(a[9]), .Z(n501) );
  NANDN U556 ( .A(n5275), .B(n501), .Z(n461) );
  AND U557 ( .A(n462), .B(n461), .Z(n520) );
  NANDN U558 ( .A(n5176), .B(n463), .Z(n465) );
  XOR U559 ( .A(b[3]), .B(a[13]), .Z(n504) );
  NANDN U560 ( .A(n5177), .B(n504), .Z(n464) );
  NAND U561 ( .A(n465), .B(n464), .Z(n519) );
  XNOR U562 ( .A(n520), .B(n519), .Z(n522) );
  AND U563 ( .A(b[0]), .B(a[15]), .Z(n466) );
  XOR U564 ( .A(b[1]), .B(n466), .Z(n468) );
  NANDN U565 ( .A(b[0]), .B(a[14]), .Z(n467) );
  AND U566 ( .A(n468), .B(n467), .Z(n515) );
  NANDN U567 ( .A(n5249), .B(n469), .Z(n471) );
  XOR U568 ( .A(b[5]), .B(a[11]), .Z(n510) );
  NANDN U569 ( .A(n5184), .B(n510), .Z(n470) );
  AND U570 ( .A(n471), .B(n470), .Z(n514) );
  AND U571 ( .A(b[7]), .B(a[7]), .Z(n513) );
  XOR U572 ( .A(n514), .B(n513), .Z(n516) );
  XNOR U573 ( .A(n515), .B(n516), .Z(n521) );
  XOR U574 ( .A(n522), .B(n521), .Z(n496) );
  NANDN U575 ( .A(n473), .B(n472), .Z(n477) );
  NANDN U576 ( .A(n475), .B(n474), .Z(n476) );
  AND U577 ( .A(n477), .B(n476), .Z(n495) );
  XNOR U578 ( .A(n496), .B(n495), .Z(n497) );
  NANDN U579 ( .A(n479), .B(n478), .Z(n483) );
  NAND U580 ( .A(n481), .B(n480), .Z(n482) );
  NAND U581 ( .A(n483), .B(n482), .Z(n498) );
  XNOR U582 ( .A(n497), .B(n498), .Z(n489) );
  XNOR U583 ( .A(n490), .B(n489), .Z(n491) );
  XNOR U584 ( .A(n492), .B(n491), .Z(n525) );
  XNOR U585 ( .A(sreg[135]), .B(n525), .Z(n527) );
  NANDN U586 ( .A(sreg[134]), .B(n484), .Z(n488) );
  NAND U587 ( .A(n486), .B(n485), .Z(n487) );
  NAND U588 ( .A(n488), .B(n487), .Z(n526) );
  XNOR U589 ( .A(n527), .B(n526), .Z(c[135]) );
  NANDN U590 ( .A(n490), .B(n489), .Z(n494) );
  NANDN U591 ( .A(n492), .B(n491), .Z(n493) );
  AND U592 ( .A(n494), .B(n493), .Z(n533) );
  NANDN U593 ( .A(n496), .B(n495), .Z(n500) );
  NANDN U594 ( .A(n498), .B(n497), .Z(n499) );
  AND U595 ( .A(n500), .B(n499), .Z(n531) );
  NANDN U596 ( .A(n5274), .B(n501), .Z(n503) );
  XOR U597 ( .A(b[7]), .B(a[10]), .Z(n542) );
  NANDN U598 ( .A(n5275), .B(n542), .Z(n502) );
  AND U599 ( .A(n503), .B(n502), .Z(n561) );
  NANDN U600 ( .A(n5176), .B(n504), .Z(n506) );
  XOR U601 ( .A(b[3]), .B(a[14]), .Z(n545) );
  NANDN U602 ( .A(n5177), .B(n545), .Z(n505) );
  NAND U603 ( .A(n506), .B(n505), .Z(n560) );
  XNOR U604 ( .A(n561), .B(n560), .Z(n563) );
  NAND U605 ( .A(b[0]), .B(a[16]), .Z(n507) );
  XNOR U606 ( .A(b[1]), .B(n507), .Z(n509) );
  NANDN U607 ( .A(b[0]), .B(a[15]), .Z(n508) );
  NAND U608 ( .A(n509), .B(n508), .Z(n557) );
  NANDN U609 ( .A(n5249), .B(n510), .Z(n512) );
  XOR U610 ( .A(b[5]), .B(a[12]), .Z(n551) );
  NANDN U611 ( .A(n5184), .B(n551), .Z(n511) );
  AND U612 ( .A(n512), .B(n511), .Z(n555) );
  AND U613 ( .A(b[7]), .B(a[8]), .Z(n554) );
  XNOR U614 ( .A(n555), .B(n554), .Z(n556) );
  XNOR U615 ( .A(n557), .B(n556), .Z(n562) );
  XOR U616 ( .A(n563), .B(n562), .Z(n537) );
  NANDN U617 ( .A(n514), .B(n513), .Z(n518) );
  NANDN U618 ( .A(n516), .B(n515), .Z(n517) );
  AND U619 ( .A(n518), .B(n517), .Z(n536) );
  XNOR U620 ( .A(n537), .B(n536), .Z(n538) );
  NANDN U621 ( .A(n520), .B(n519), .Z(n524) );
  NAND U622 ( .A(n522), .B(n521), .Z(n523) );
  NAND U623 ( .A(n524), .B(n523), .Z(n539) );
  XNOR U624 ( .A(n538), .B(n539), .Z(n530) );
  XNOR U625 ( .A(n531), .B(n530), .Z(n532) );
  XNOR U626 ( .A(n533), .B(n532), .Z(n566) );
  XNOR U627 ( .A(sreg[136]), .B(n566), .Z(n568) );
  NANDN U628 ( .A(sreg[135]), .B(n525), .Z(n529) );
  NAND U629 ( .A(n527), .B(n526), .Z(n528) );
  NAND U630 ( .A(n529), .B(n528), .Z(n567) );
  XNOR U631 ( .A(n568), .B(n567), .Z(c[136]) );
  NANDN U632 ( .A(n531), .B(n530), .Z(n535) );
  NANDN U633 ( .A(n533), .B(n532), .Z(n534) );
  AND U634 ( .A(n535), .B(n534), .Z(n574) );
  NANDN U635 ( .A(n537), .B(n536), .Z(n541) );
  NANDN U636 ( .A(n539), .B(n538), .Z(n540) );
  AND U637 ( .A(n541), .B(n540), .Z(n572) );
  NANDN U638 ( .A(n5274), .B(n542), .Z(n544) );
  XOR U639 ( .A(b[7]), .B(a[11]), .Z(n583) );
  NANDN U640 ( .A(n5275), .B(n583), .Z(n543) );
  AND U641 ( .A(n544), .B(n543), .Z(n602) );
  NANDN U642 ( .A(n5176), .B(n545), .Z(n547) );
  XOR U643 ( .A(b[3]), .B(a[15]), .Z(n586) );
  NANDN U644 ( .A(n5177), .B(n586), .Z(n546) );
  NAND U645 ( .A(n547), .B(n546), .Z(n601) );
  XNOR U646 ( .A(n602), .B(n601), .Z(n604) );
  NAND U647 ( .A(b[0]), .B(a[17]), .Z(n548) );
  XNOR U648 ( .A(b[1]), .B(n548), .Z(n550) );
  NANDN U649 ( .A(b[0]), .B(a[16]), .Z(n549) );
  NAND U650 ( .A(n550), .B(n549), .Z(n598) );
  NANDN U651 ( .A(n5249), .B(n551), .Z(n553) );
  XOR U652 ( .A(b[5]), .B(a[13]), .Z(n592) );
  NANDN U653 ( .A(n5184), .B(n592), .Z(n552) );
  AND U654 ( .A(n553), .B(n552), .Z(n596) );
  AND U655 ( .A(b[7]), .B(a[9]), .Z(n595) );
  XNOR U656 ( .A(n596), .B(n595), .Z(n597) );
  XNOR U657 ( .A(n598), .B(n597), .Z(n603) );
  XOR U658 ( .A(n604), .B(n603), .Z(n578) );
  NANDN U659 ( .A(n555), .B(n554), .Z(n559) );
  NANDN U660 ( .A(n557), .B(n556), .Z(n558) );
  AND U661 ( .A(n559), .B(n558), .Z(n577) );
  XNOR U662 ( .A(n578), .B(n577), .Z(n579) );
  NANDN U663 ( .A(n561), .B(n560), .Z(n565) );
  NAND U664 ( .A(n563), .B(n562), .Z(n564) );
  NAND U665 ( .A(n565), .B(n564), .Z(n580) );
  XNOR U666 ( .A(n579), .B(n580), .Z(n571) );
  XNOR U667 ( .A(n572), .B(n571), .Z(n573) );
  XNOR U668 ( .A(n574), .B(n573), .Z(n607) );
  XNOR U669 ( .A(sreg[137]), .B(n607), .Z(n609) );
  NANDN U670 ( .A(sreg[136]), .B(n566), .Z(n570) );
  NAND U671 ( .A(n568), .B(n567), .Z(n569) );
  NAND U672 ( .A(n570), .B(n569), .Z(n608) );
  XNOR U673 ( .A(n609), .B(n608), .Z(c[137]) );
  NANDN U674 ( .A(n572), .B(n571), .Z(n576) );
  NANDN U675 ( .A(n574), .B(n573), .Z(n575) );
  AND U676 ( .A(n576), .B(n575), .Z(n615) );
  NANDN U677 ( .A(n578), .B(n577), .Z(n582) );
  NANDN U678 ( .A(n580), .B(n579), .Z(n581) );
  AND U679 ( .A(n582), .B(n581), .Z(n613) );
  NANDN U680 ( .A(n5274), .B(n583), .Z(n585) );
  XOR U681 ( .A(b[7]), .B(a[12]), .Z(n624) );
  NANDN U682 ( .A(n5275), .B(n624), .Z(n584) );
  AND U683 ( .A(n585), .B(n584), .Z(n643) );
  NANDN U684 ( .A(n5176), .B(n586), .Z(n588) );
  XOR U685 ( .A(b[3]), .B(a[16]), .Z(n627) );
  NANDN U686 ( .A(n5177), .B(n627), .Z(n587) );
  NAND U687 ( .A(n588), .B(n587), .Z(n642) );
  XNOR U688 ( .A(n643), .B(n642), .Z(n645) );
  NAND U689 ( .A(b[0]), .B(a[18]), .Z(n589) );
  XNOR U690 ( .A(b[1]), .B(n589), .Z(n591) );
  NANDN U691 ( .A(b[0]), .B(a[17]), .Z(n590) );
  NAND U692 ( .A(n591), .B(n590), .Z(n639) );
  NANDN U693 ( .A(n5249), .B(n592), .Z(n594) );
  XOR U694 ( .A(b[5]), .B(a[14]), .Z(n633) );
  NANDN U695 ( .A(n5184), .B(n633), .Z(n593) );
  AND U696 ( .A(n594), .B(n593), .Z(n637) );
  AND U697 ( .A(b[7]), .B(a[10]), .Z(n636) );
  XNOR U698 ( .A(n637), .B(n636), .Z(n638) );
  XNOR U699 ( .A(n639), .B(n638), .Z(n644) );
  XOR U700 ( .A(n645), .B(n644), .Z(n619) );
  NANDN U701 ( .A(n596), .B(n595), .Z(n600) );
  NANDN U702 ( .A(n598), .B(n597), .Z(n599) );
  AND U703 ( .A(n600), .B(n599), .Z(n618) );
  XNOR U704 ( .A(n619), .B(n618), .Z(n620) );
  NANDN U705 ( .A(n602), .B(n601), .Z(n606) );
  NAND U706 ( .A(n604), .B(n603), .Z(n605) );
  NAND U707 ( .A(n606), .B(n605), .Z(n621) );
  XNOR U708 ( .A(n620), .B(n621), .Z(n612) );
  XNOR U709 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U710 ( .A(n615), .B(n614), .Z(n648) );
  XNOR U711 ( .A(sreg[138]), .B(n648), .Z(n650) );
  NANDN U712 ( .A(sreg[137]), .B(n607), .Z(n611) );
  NAND U713 ( .A(n609), .B(n608), .Z(n610) );
  NAND U714 ( .A(n611), .B(n610), .Z(n649) );
  XNOR U715 ( .A(n650), .B(n649), .Z(c[138]) );
  NANDN U716 ( .A(n613), .B(n612), .Z(n617) );
  NANDN U717 ( .A(n615), .B(n614), .Z(n616) );
  AND U718 ( .A(n617), .B(n616), .Z(n656) );
  NANDN U719 ( .A(n619), .B(n618), .Z(n623) );
  NANDN U720 ( .A(n621), .B(n620), .Z(n622) );
  AND U721 ( .A(n623), .B(n622), .Z(n654) );
  NANDN U722 ( .A(n5274), .B(n624), .Z(n626) );
  XOR U723 ( .A(b[7]), .B(a[13]), .Z(n665) );
  NANDN U724 ( .A(n5275), .B(n665), .Z(n625) );
  AND U725 ( .A(n626), .B(n625), .Z(n684) );
  NANDN U726 ( .A(n5176), .B(n627), .Z(n629) );
  XOR U727 ( .A(b[3]), .B(a[17]), .Z(n668) );
  NANDN U728 ( .A(n5177), .B(n668), .Z(n628) );
  NAND U729 ( .A(n629), .B(n628), .Z(n683) );
  XNOR U730 ( .A(n684), .B(n683), .Z(n686) );
  NAND U731 ( .A(b[0]), .B(a[19]), .Z(n630) );
  XNOR U732 ( .A(b[1]), .B(n630), .Z(n632) );
  NANDN U733 ( .A(b[0]), .B(a[18]), .Z(n631) );
  NAND U734 ( .A(n632), .B(n631), .Z(n680) );
  NANDN U735 ( .A(n5249), .B(n633), .Z(n635) );
  XOR U736 ( .A(b[5]), .B(a[15]), .Z(n674) );
  NANDN U737 ( .A(n5184), .B(n674), .Z(n634) );
  AND U738 ( .A(n635), .B(n634), .Z(n678) );
  AND U739 ( .A(b[7]), .B(a[11]), .Z(n677) );
  XNOR U740 ( .A(n678), .B(n677), .Z(n679) );
  XNOR U741 ( .A(n680), .B(n679), .Z(n685) );
  XOR U742 ( .A(n686), .B(n685), .Z(n660) );
  NANDN U743 ( .A(n637), .B(n636), .Z(n641) );
  NANDN U744 ( .A(n639), .B(n638), .Z(n640) );
  AND U745 ( .A(n641), .B(n640), .Z(n659) );
  XNOR U746 ( .A(n660), .B(n659), .Z(n661) );
  NANDN U747 ( .A(n643), .B(n642), .Z(n647) );
  NAND U748 ( .A(n645), .B(n644), .Z(n646) );
  NAND U749 ( .A(n647), .B(n646), .Z(n662) );
  XNOR U750 ( .A(n661), .B(n662), .Z(n653) );
  XNOR U751 ( .A(n654), .B(n653), .Z(n655) );
  XNOR U752 ( .A(n656), .B(n655), .Z(n689) );
  XNOR U753 ( .A(sreg[139]), .B(n689), .Z(n691) );
  NANDN U754 ( .A(sreg[138]), .B(n648), .Z(n652) );
  NAND U755 ( .A(n650), .B(n649), .Z(n651) );
  NAND U756 ( .A(n652), .B(n651), .Z(n690) );
  XNOR U757 ( .A(n691), .B(n690), .Z(c[139]) );
  NANDN U758 ( .A(n654), .B(n653), .Z(n658) );
  NANDN U759 ( .A(n656), .B(n655), .Z(n657) );
  AND U760 ( .A(n658), .B(n657), .Z(n697) );
  NANDN U761 ( .A(n660), .B(n659), .Z(n664) );
  NANDN U762 ( .A(n662), .B(n661), .Z(n663) );
  AND U763 ( .A(n664), .B(n663), .Z(n695) );
  NANDN U764 ( .A(n5274), .B(n665), .Z(n667) );
  XOR U765 ( .A(b[7]), .B(a[14]), .Z(n706) );
  NANDN U766 ( .A(n5275), .B(n706), .Z(n666) );
  AND U767 ( .A(n667), .B(n666), .Z(n725) );
  NANDN U768 ( .A(n5176), .B(n668), .Z(n670) );
  XOR U769 ( .A(b[3]), .B(a[18]), .Z(n709) );
  NANDN U770 ( .A(n5177), .B(n709), .Z(n669) );
  NAND U771 ( .A(n670), .B(n669), .Z(n724) );
  XNOR U772 ( .A(n725), .B(n724), .Z(n727) );
  NAND U773 ( .A(b[0]), .B(a[20]), .Z(n671) );
  XNOR U774 ( .A(b[1]), .B(n671), .Z(n673) );
  NANDN U775 ( .A(b[0]), .B(a[19]), .Z(n672) );
  NAND U776 ( .A(n673), .B(n672), .Z(n721) );
  NANDN U777 ( .A(n5249), .B(n674), .Z(n676) );
  XOR U778 ( .A(b[5]), .B(a[16]), .Z(n715) );
  NANDN U779 ( .A(n5184), .B(n715), .Z(n675) );
  AND U780 ( .A(n676), .B(n675), .Z(n719) );
  AND U781 ( .A(b[7]), .B(a[12]), .Z(n718) );
  XNOR U782 ( .A(n719), .B(n718), .Z(n720) );
  XNOR U783 ( .A(n721), .B(n720), .Z(n726) );
  XOR U784 ( .A(n727), .B(n726), .Z(n701) );
  NANDN U785 ( .A(n678), .B(n677), .Z(n682) );
  NANDN U786 ( .A(n680), .B(n679), .Z(n681) );
  AND U787 ( .A(n682), .B(n681), .Z(n700) );
  XNOR U788 ( .A(n701), .B(n700), .Z(n702) );
  NANDN U789 ( .A(n684), .B(n683), .Z(n688) );
  NAND U790 ( .A(n686), .B(n685), .Z(n687) );
  NAND U791 ( .A(n688), .B(n687), .Z(n703) );
  XNOR U792 ( .A(n702), .B(n703), .Z(n694) );
  XNOR U793 ( .A(n695), .B(n694), .Z(n696) );
  XNOR U794 ( .A(n697), .B(n696), .Z(n730) );
  XNOR U795 ( .A(sreg[140]), .B(n730), .Z(n732) );
  NANDN U796 ( .A(sreg[139]), .B(n689), .Z(n693) );
  NAND U797 ( .A(n691), .B(n690), .Z(n692) );
  NAND U798 ( .A(n693), .B(n692), .Z(n731) );
  XNOR U799 ( .A(n732), .B(n731), .Z(c[140]) );
  NANDN U800 ( .A(n695), .B(n694), .Z(n699) );
  NANDN U801 ( .A(n697), .B(n696), .Z(n698) );
  AND U802 ( .A(n699), .B(n698), .Z(n738) );
  NANDN U803 ( .A(n701), .B(n700), .Z(n705) );
  NANDN U804 ( .A(n703), .B(n702), .Z(n704) );
  AND U805 ( .A(n705), .B(n704), .Z(n736) );
  NANDN U806 ( .A(n5274), .B(n706), .Z(n708) );
  XOR U807 ( .A(b[7]), .B(a[15]), .Z(n747) );
  NANDN U808 ( .A(n5275), .B(n747), .Z(n707) );
  AND U809 ( .A(n708), .B(n707), .Z(n766) );
  NANDN U810 ( .A(n5176), .B(n709), .Z(n711) );
  XOR U811 ( .A(b[3]), .B(a[19]), .Z(n750) );
  NANDN U812 ( .A(n5177), .B(n750), .Z(n710) );
  NAND U813 ( .A(n711), .B(n710), .Z(n765) );
  XNOR U814 ( .A(n766), .B(n765), .Z(n768) );
  NAND U815 ( .A(b[0]), .B(a[21]), .Z(n712) );
  XNOR U816 ( .A(b[1]), .B(n712), .Z(n714) );
  NANDN U817 ( .A(b[0]), .B(a[20]), .Z(n713) );
  NAND U818 ( .A(n714), .B(n713), .Z(n762) );
  NANDN U819 ( .A(n5249), .B(n715), .Z(n717) );
  XOR U820 ( .A(b[5]), .B(a[17]), .Z(n756) );
  NANDN U821 ( .A(n5184), .B(n756), .Z(n716) );
  AND U822 ( .A(n717), .B(n716), .Z(n760) );
  AND U823 ( .A(b[7]), .B(a[13]), .Z(n759) );
  XNOR U824 ( .A(n760), .B(n759), .Z(n761) );
  XNOR U825 ( .A(n762), .B(n761), .Z(n767) );
  XOR U826 ( .A(n768), .B(n767), .Z(n742) );
  NANDN U827 ( .A(n719), .B(n718), .Z(n723) );
  NANDN U828 ( .A(n721), .B(n720), .Z(n722) );
  AND U829 ( .A(n723), .B(n722), .Z(n741) );
  XNOR U830 ( .A(n742), .B(n741), .Z(n743) );
  NANDN U831 ( .A(n725), .B(n724), .Z(n729) );
  NAND U832 ( .A(n727), .B(n726), .Z(n728) );
  NAND U833 ( .A(n729), .B(n728), .Z(n744) );
  XNOR U834 ( .A(n743), .B(n744), .Z(n735) );
  XNOR U835 ( .A(n736), .B(n735), .Z(n737) );
  XNOR U836 ( .A(n738), .B(n737), .Z(n771) );
  XNOR U837 ( .A(sreg[141]), .B(n771), .Z(n773) );
  NANDN U838 ( .A(sreg[140]), .B(n730), .Z(n734) );
  NAND U839 ( .A(n732), .B(n731), .Z(n733) );
  NAND U840 ( .A(n734), .B(n733), .Z(n772) );
  XNOR U841 ( .A(n773), .B(n772), .Z(c[141]) );
  NANDN U842 ( .A(n736), .B(n735), .Z(n740) );
  NANDN U843 ( .A(n738), .B(n737), .Z(n739) );
  AND U844 ( .A(n740), .B(n739), .Z(n779) );
  NANDN U845 ( .A(n742), .B(n741), .Z(n746) );
  NANDN U846 ( .A(n744), .B(n743), .Z(n745) );
  AND U847 ( .A(n746), .B(n745), .Z(n777) );
  NANDN U848 ( .A(n5274), .B(n747), .Z(n749) );
  XOR U849 ( .A(b[7]), .B(a[16]), .Z(n788) );
  NANDN U850 ( .A(n5275), .B(n788), .Z(n748) );
  AND U851 ( .A(n749), .B(n748), .Z(n807) );
  NANDN U852 ( .A(n5176), .B(n750), .Z(n752) );
  XOR U853 ( .A(b[3]), .B(a[20]), .Z(n791) );
  NANDN U854 ( .A(n5177), .B(n791), .Z(n751) );
  NAND U855 ( .A(n752), .B(n751), .Z(n806) );
  XNOR U856 ( .A(n807), .B(n806), .Z(n809) );
  NAND U857 ( .A(b[0]), .B(a[22]), .Z(n753) );
  XNOR U858 ( .A(b[1]), .B(n753), .Z(n755) );
  NANDN U859 ( .A(b[0]), .B(a[21]), .Z(n754) );
  NAND U860 ( .A(n755), .B(n754), .Z(n803) );
  NANDN U861 ( .A(n5249), .B(n756), .Z(n758) );
  XOR U862 ( .A(b[5]), .B(a[18]), .Z(n794) );
  NANDN U863 ( .A(n5184), .B(n794), .Z(n757) );
  AND U864 ( .A(n758), .B(n757), .Z(n801) );
  AND U865 ( .A(b[7]), .B(a[14]), .Z(n800) );
  XNOR U866 ( .A(n801), .B(n800), .Z(n802) );
  XNOR U867 ( .A(n803), .B(n802), .Z(n808) );
  XOR U868 ( .A(n809), .B(n808), .Z(n783) );
  NANDN U869 ( .A(n760), .B(n759), .Z(n764) );
  NANDN U870 ( .A(n762), .B(n761), .Z(n763) );
  AND U871 ( .A(n764), .B(n763), .Z(n782) );
  XNOR U872 ( .A(n783), .B(n782), .Z(n784) );
  NANDN U873 ( .A(n766), .B(n765), .Z(n770) );
  NAND U874 ( .A(n768), .B(n767), .Z(n769) );
  NAND U875 ( .A(n770), .B(n769), .Z(n785) );
  XNOR U876 ( .A(n784), .B(n785), .Z(n776) );
  XNOR U877 ( .A(n777), .B(n776), .Z(n778) );
  XNOR U878 ( .A(n779), .B(n778), .Z(n812) );
  XNOR U879 ( .A(sreg[142]), .B(n812), .Z(n814) );
  NANDN U880 ( .A(sreg[141]), .B(n771), .Z(n775) );
  NAND U881 ( .A(n773), .B(n772), .Z(n774) );
  NAND U882 ( .A(n775), .B(n774), .Z(n813) );
  XNOR U883 ( .A(n814), .B(n813), .Z(c[142]) );
  NANDN U884 ( .A(n777), .B(n776), .Z(n781) );
  NANDN U885 ( .A(n779), .B(n778), .Z(n780) );
  AND U886 ( .A(n781), .B(n780), .Z(n820) );
  NANDN U887 ( .A(n783), .B(n782), .Z(n787) );
  NANDN U888 ( .A(n785), .B(n784), .Z(n786) );
  AND U889 ( .A(n787), .B(n786), .Z(n818) );
  NANDN U890 ( .A(n5274), .B(n788), .Z(n790) );
  XOR U891 ( .A(b[7]), .B(a[17]), .Z(n829) );
  NANDN U892 ( .A(n5275), .B(n829), .Z(n789) );
  AND U893 ( .A(n790), .B(n789), .Z(n848) );
  NANDN U894 ( .A(n5176), .B(n791), .Z(n793) );
  XOR U895 ( .A(b[3]), .B(a[21]), .Z(n832) );
  NANDN U896 ( .A(n5177), .B(n832), .Z(n792) );
  NAND U897 ( .A(n793), .B(n792), .Z(n847) );
  XNOR U898 ( .A(n848), .B(n847), .Z(n850) );
  NANDN U899 ( .A(n5249), .B(n794), .Z(n796) );
  XOR U900 ( .A(b[5]), .B(a[19]), .Z(n838) );
  NANDN U901 ( .A(n5184), .B(n838), .Z(n795) );
  AND U902 ( .A(n796), .B(n795), .Z(n842) );
  AND U903 ( .A(b[7]), .B(a[15]), .Z(n841) );
  XNOR U904 ( .A(n842), .B(n841), .Z(n843) );
  NAND U905 ( .A(b[0]), .B(a[23]), .Z(n797) );
  XNOR U906 ( .A(b[1]), .B(n797), .Z(n799) );
  NANDN U907 ( .A(b[0]), .B(a[22]), .Z(n798) );
  NAND U908 ( .A(n799), .B(n798), .Z(n844) );
  XNOR U909 ( .A(n843), .B(n844), .Z(n849) );
  XOR U910 ( .A(n850), .B(n849), .Z(n824) );
  NANDN U911 ( .A(n801), .B(n800), .Z(n805) );
  NANDN U912 ( .A(n803), .B(n802), .Z(n804) );
  AND U913 ( .A(n805), .B(n804), .Z(n823) );
  XNOR U914 ( .A(n824), .B(n823), .Z(n825) );
  NANDN U915 ( .A(n807), .B(n806), .Z(n811) );
  NAND U916 ( .A(n809), .B(n808), .Z(n810) );
  NAND U917 ( .A(n811), .B(n810), .Z(n826) );
  XNOR U918 ( .A(n825), .B(n826), .Z(n817) );
  XNOR U919 ( .A(n818), .B(n817), .Z(n819) );
  XNOR U920 ( .A(n820), .B(n819), .Z(n853) );
  XNOR U921 ( .A(sreg[143]), .B(n853), .Z(n855) );
  NANDN U922 ( .A(sreg[142]), .B(n812), .Z(n816) );
  NAND U923 ( .A(n814), .B(n813), .Z(n815) );
  NAND U924 ( .A(n816), .B(n815), .Z(n854) );
  XNOR U925 ( .A(n855), .B(n854), .Z(c[143]) );
  NANDN U926 ( .A(n818), .B(n817), .Z(n822) );
  NANDN U927 ( .A(n820), .B(n819), .Z(n821) );
  AND U928 ( .A(n822), .B(n821), .Z(n861) );
  NANDN U929 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U930 ( .A(n826), .B(n825), .Z(n827) );
  AND U931 ( .A(n828), .B(n827), .Z(n859) );
  NANDN U932 ( .A(n5274), .B(n829), .Z(n831) );
  XOR U933 ( .A(b[7]), .B(a[18]), .Z(n870) );
  NANDN U934 ( .A(n5275), .B(n870), .Z(n830) );
  AND U935 ( .A(n831), .B(n830), .Z(n889) );
  NANDN U936 ( .A(n5176), .B(n832), .Z(n834) );
  XOR U937 ( .A(b[3]), .B(a[22]), .Z(n873) );
  NANDN U938 ( .A(n5177), .B(n873), .Z(n833) );
  NAND U939 ( .A(n834), .B(n833), .Z(n888) );
  XNOR U940 ( .A(n889), .B(n888), .Z(n891) );
  NAND U941 ( .A(b[0]), .B(a[24]), .Z(n835) );
  XNOR U942 ( .A(b[1]), .B(n835), .Z(n837) );
  NANDN U943 ( .A(b[0]), .B(a[23]), .Z(n836) );
  NAND U944 ( .A(n837), .B(n836), .Z(n885) );
  NANDN U945 ( .A(n5249), .B(n838), .Z(n840) );
  XOR U946 ( .A(b[5]), .B(a[20]), .Z(n879) );
  NANDN U947 ( .A(n5184), .B(n879), .Z(n839) );
  AND U948 ( .A(n840), .B(n839), .Z(n883) );
  AND U949 ( .A(b[7]), .B(a[16]), .Z(n882) );
  XNOR U950 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U951 ( .A(n885), .B(n884), .Z(n890) );
  XOR U952 ( .A(n891), .B(n890), .Z(n865) );
  NANDN U953 ( .A(n842), .B(n841), .Z(n846) );
  NANDN U954 ( .A(n844), .B(n843), .Z(n845) );
  AND U955 ( .A(n846), .B(n845), .Z(n864) );
  XNOR U956 ( .A(n865), .B(n864), .Z(n866) );
  NANDN U957 ( .A(n848), .B(n847), .Z(n852) );
  NAND U958 ( .A(n850), .B(n849), .Z(n851) );
  NAND U959 ( .A(n852), .B(n851), .Z(n867) );
  XNOR U960 ( .A(n866), .B(n867), .Z(n858) );
  XNOR U961 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U962 ( .A(n861), .B(n860), .Z(n894) );
  XNOR U963 ( .A(sreg[144]), .B(n894), .Z(n896) );
  NANDN U964 ( .A(sreg[143]), .B(n853), .Z(n857) );
  NAND U965 ( .A(n855), .B(n854), .Z(n856) );
  NAND U966 ( .A(n857), .B(n856), .Z(n895) );
  XNOR U967 ( .A(n896), .B(n895), .Z(c[144]) );
  NANDN U968 ( .A(n859), .B(n858), .Z(n863) );
  NANDN U969 ( .A(n861), .B(n860), .Z(n862) );
  AND U970 ( .A(n863), .B(n862), .Z(n902) );
  NANDN U971 ( .A(n865), .B(n864), .Z(n869) );
  NANDN U972 ( .A(n867), .B(n866), .Z(n868) );
  AND U973 ( .A(n869), .B(n868), .Z(n900) );
  NANDN U974 ( .A(n5274), .B(n870), .Z(n872) );
  XOR U975 ( .A(b[7]), .B(a[19]), .Z(n911) );
  NANDN U976 ( .A(n5275), .B(n911), .Z(n871) );
  AND U977 ( .A(n872), .B(n871), .Z(n930) );
  NANDN U978 ( .A(n5176), .B(n873), .Z(n875) );
  XOR U979 ( .A(b[3]), .B(a[23]), .Z(n914) );
  NANDN U980 ( .A(n5177), .B(n914), .Z(n874) );
  NAND U981 ( .A(n875), .B(n874), .Z(n929) );
  XNOR U982 ( .A(n930), .B(n929), .Z(n932) );
  NAND U983 ( .A(b[0]), .B(a[25]), .Z(n876) );
  XNOR U984 ( .A(b[1]), .B(n876), .Z(n878) );
  NANDN U985 ( .A(b[0]), .B(a[24]), .Z(n877) );
  NAND U986 ( .A(n878), .B(n877), .Z(n926) );
  NANDN U987 ( .A(n5249), .B(n879), .Z(n881) );
  XOR U988 ( .A(b[5]), .B(a[21]), .Z(n917) );
  NANDN U989 ( .A(n5184), .B(n917), .Z(n880) );
  AND U990 ( .A(n881), .B(n880), .Z(n924) );
  AND U991 ( .A(b[7]), .B(a[17]), .Z(n923) );
  XNOR U992 ( .A(n924), .B(n923), .Z(n925) );
  XNOR U993 ( .A(n926), .B(n925), .Z(n931) );
  XOR U994 ( .A(n932), .B(n931), .Z(n906) );
  NANDN U995 ( .A(n883), .B(n882), .Z(n887) );
  NANDN U996 ( .A(n885), .B(n884), .Z(n886) );
  AND U997 ( .A(n887), .B(n886), .Z(n905) );
  XNOR U998 ( .A(n906), .B(n905), .Z(n907) );
  NANDN U999 ( .A(n889), .B(n888), .Z(n893) );
  NAND U1000 ( .A(n891), .B(n890), .Z(n892) );
  NAND U1001 ( .A(n893), .B(n892), .Z(n908) );
  XNOR U1002 ( .A(n907), .B(n908), .Z(n899) );
  XNOR U1003 ( .A(n900), .B(n899), .Z(n901) );
  XNOR U1004 ( .A(n902), .B(n901), .Z(n935) );
  XNOR U1005 ( .A(sreg[145]), .B(n935), .Z(n937) );
  NANDN U1006 ( .A(sreg[144]), .B(n894), .Z(n898) );
  NAND U1007 ( .A(n896), .B(n895), .Z(n897) );
  NAND U1008 ( .A(n898), .B(n897), .Z(n936) );
  XNOR U1009 ( .A(n937), .B(n936), .Z(c[145]) );
  NANDN U1010 ( .A(n900), .B(n899), .Z(n904) );
  NANDN U1011 ( .A(n902), .B(n901), .Z(n903) );
  AND U1012 ( .A(n904), .B(n903), .Z(n943) );
  NANDN U1013 ( .A(n906), .B(n905), .Z(n910) );
  NANDN U1014 ( .A(n908), .B(n907), .Z(n909) );
  AND U1015 ( .A(n910), .B(n909), .Z(n941) );
  NANDN U1016 ( .A(n5274), .B(n911), .Z(n913) );
  XOR U1017 ( .A(b[7]), .B(a[20]), .Z(n952) );
  NANDN U1018 ( .A(n5275), .B(n952), .Z(n912) );
  AND U1019 ( .A(n913), .B(n912), .Z(n971) );
  NANDN U1020 ( .A(n5176), .B(n914), .Z(n916) );
  XOR U1021 ( .A(b[3]), .B(a[24]), .Z(n955) );
  NANDN U1022 ( .A(n5177), .B(n955), .Z(n915) );
  NAND U1023 ( .A(n916), .B(n915), .Z(n970) );
  XNOR U1024 ( .A(n971), .B(n970), .Z(n973) );
  NANDN U1025 ( .A(n5249), .B(n917), .Z(n919) );
  XOR U1026 ( .A(b[5]), .B(a[22]), .Z(n961) );
  NANDN U1027 ( .A(n5184), .B(n961), .Z(n918) );
  AND U1028 ( .A(n919), .B(n918), .Z(n965) );
  AND U1029 ( .A(b[7]), .B(a[18]), .Z(n964) );
  XNOR U1030 ( .A(n965), .B(n964), .Z(n966) );
  NAND U1031 ( .A(b[0]), .B(a[26]), .Z(n920) );
  XNOR U1032 ( .A(b[1]), .B(n920), .Z(n922) );
  NANDN U1033 ( .A(b[0]), .B(a[25]), .Z(n921) );
  NAND U1034 ( .A(n922), .B(n921), .Z(n967) );
  XNOR U1035 ( .A(n966), .B(n967), .Z(n972) );
  XOR U1036 ( .A(n973), .B(n972), .Z(n947) );
  NANDN U1037 ( .A(n924), .B(n923), .Z(n928) );
  NANDN U1038 ( .A(n926), .B(n925), .Z(n927) );
  AND U1039 ( .A(n928), .B(n927), .Z(n946) );
  XNOR U1040 ( .A(n947), .B(n946), .Z(n948) );
  NANDN U1041 ( .A(n930), .B(n929), .Z(n934) );
  NAND U1042 ( .A(n932), .B(n931), .Z(n933) );
  NAND U1043 ( .A(n934), .B(n933), .Z(n949) );
  XNOR U1044 ( .A(n948), .B(n949), .Z(n940) );
  XNOR U1045 ( .A(n941), .B(n940), .Z(n942) );
  XNOR U1046 ( .A(n943), .B(n942), .Z(n976) );
  XNOR U1047 ( .A(sreg[146]), .B(n976), .Z(n978) );
  NANDN U1048 ( .A(sreg[145]), .B(n935), .Z(n939) );
  NAND U1049 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1050 ( .A(n939), .B(n938), .Z(n977) );
  XNOR U1051 ( .A(n978), .B(n977), .Z(c[146]) );
  NANDN U1052 ( .A(n941), .B(n940), .Z(n945) );
  NANDN U1053 ( .A(n943), .B(n942), .Z(n944) );
  AND U1054 ( .A(n945), .B(n944), .Z(n984) );
  NANDN U1055 ( .A(n947), .B(n946), .Z(n951) );
  NANDN U1056 ( .A(n949), .B(n948), .Z(n950) );
  AND U1057 ( .A(n951), .B(n950), .Z(n982) );
  NANDN U1058 ( .A(n5274), .B(n952), .Z(n954) );
  XOR U1059 ( .A(b[7]), .B(a[21]), .Z(n993) );
  NANDN U1060 ( .A(n5275), .B(n993), .Z(n953) );
  AND U1061 ( .A(n954), .B(n953), .Z(n1012) );
  NANDN U1062 ( .A(n5176), .B(n955), .Z(n957) );
  XOR U1063 ( .A(b[3]), .B(a[25]), .Z(n996) );
  NANDN U1064 ( .A(n5177), .B(n996), .Z(n956) );
  NAND U1065 ( .A(n957), .B(n956), .Z(n1011) );
  XNOR U1066 ( .A(n1012), .B(n1011), .Z(n1014) );
  NAND U1067 ( .A(b[0]), .B(a[27]), .Z(n958) );
  XNOR U1068 ( .A(b[1]), .B(n958), .Z(n960) );
  NANDN U1069 ( .A(b[0]), .B(a[26]), .Z(n959) );
  NAND U1070 ( .A(n960), .B(n959), .Z(n1008) );
  NANDN U1071 ( .A(n5249), .B(n961), .Z(n963) );
  XOR U1072 ( .A(b[5]), .B(a[23]), .Z(n1002) );
  NANDN U1073 ( .A(n5184), .B(n1002), .Z(n962) );
  AND U1074 ( .A(n963), .B(n962), .Z(n1006) );
  AND U1075 ( .A(b[7]), .B(a[19]), .Z(n1005) );
  XNOR U1076 ( .A(n1006), .B(n1005), .Z(n1007) );
  XNOR U1077 ( .A(n1008), .B(n1007), .Z(n1013) );
  XOR U1078 ( .A(n1014), .B(n1013), .Z(n988) );
  NANDN U1079 ( .A(n965), .B(n964), .Z(n969) );
  NANDN U1080 ( .A(n967), .B(n966), .Z(n968) );
  AND U1081 ( .A(n969), .B(n968), .Z(n987) );
  XNOR U1082 ( .A(n988), .B(n987), .Z(n989) );
  NANDN U1083 ( .A(n971), .B(n970), .Z(n975) );
  NAND U1084 ( .A(n973), .B(n972), .Z(n974) );
  NAND U1085 ( .A(n975), .B(n974), .Z(n990) );
  XNOR U1086 ( .A(n989), .B(n990), .Z(n981) );
  XNOR U1087 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1088 ( .A(n984), .B(n983), .Z(n1017) );
  XNOR U1089 ( .A(sreg[147]), .B(n1017), .Z(n1019) );
  NANDN U1090 ( .A(sreg[146]), .B(n976), .Z(n980) );
  NAND U1091 ( .A(n978), .B(n977), .Z(n979) );
  NAND U1092 ( .A(n980), .B(n979), .Z(n1018) );
  XNOR U1093 ( .A(n1019), .B(n1018), .Z(c[147]) );
  NANDN U1094 ( .A(n982), .B(n981), .Z(n986) );
  NANDN U1095 ( .A(n984), .B(n983), .Z(n985) );
  AND U1096 ( .A(n986), .B(n985), .Z(n1025) );
  NANDN U1097 ( .A(n988), .B(n987), .Z(n992) );
  NANDN U1098 ( .A(n990), .B(n989), .Z(n991) );
  AND U1099 ( .A(n992), .B(n991), .Z(n1023) );
  NANDN U1100 ( .A(n5274), .B(n993), .Z(n995) );
  XOR U1101 ( .A(b[7]), .B(a[22]), .Z(n1034) );
  NANDN U1102 ( .A(n5275), .B(n1034), .Z(n994) );
  AND U1103 ( .A(n995), .B(n994), .Z(n1053) );
  NANDN U1104 ( .A(n5176), .B(n996), .Z(n998) );
  XOR U1105 ( .A(b[3]), .B(a[26]), .Z(n1037) );
  NANDN U1106 ( .A(n5177), .B(n1037), .Z(n997) );
  NAND U1107 ( .A(n998), .B(n997), .Z(n1052) );
  XNOR U1108 ( .A(n1053), .B(n1052), .Z(n1055) );
  NAND U1109 ( .A(b[0]), .B(a[28]), .Z(n999) );
  XNOR U1110 ( .A(b[1]), .B(n999), .Z(n1001) );
  NANDN U1111 ( .A(b[0]), .B(a[27]), .Z(n1000) );
  NAND U1112 ( .A(n1001), .B(n1000), .Z(n1049) );
  NANDN U1113 ( .A(n5249), .B(n1002), .Z(n1004) );
  XOR U1114 ( .A(b[5]), .B(a[24]), .Z(n1043) );
  NANDN U1115 ( .A(n5184), .B(n1043), .Z(n1003) );
  AND U1116 ( .A(n1004), .B(n1003), .Z(n1047) );
  AND U1117 ( .A(b[7]), .B(a[20]), .Z(n1046) );
  XNOR U1118 ( .A(n1047), .B(n1046), .Z(n1048) );
  XNOR U1119 ( .A(n1049), .B(n1048), .Z(n1054) );
  XOR U1120 ( .A(n1055), .B(n1054), .Z(n1029) );
  NANDN U1121 ( .A(n1006), .B(n1005), .Z(n1010) );
  NANDN U1122 ( .A(n1008), .B(n1007), .Z(n1009) );
  AND U1123 ( .A(n1010), .B(n1009), .Z(n1028) );
  XNOR U1124 ( .A(n1029), .B(n1028), .Z(n1030) );
  NANDN U1125 ( .A(n1012), .B(n1011), .Z(n1016) );
  NAND U1126 ( .A(n1014), .B(n1013), .Z(n1015) );
  NAND U1127 ( .A(n1016), .B(n1015), .Z(n1031) );
  XNOR U1128 ( .A(n1030), .B(n1031), .Z(n1022) );
  XNOR U1129 ( .A(n1023), .B(n1022), .Z(n1024) );
  XNOR U1130 ( .A(n1025), .B(n1024), .Z(n1058) );
  XNOR U1131 ( .A(sreg[148]), .B(n1058), .Z(n1060) );
  NANDN U1132 ( .A(sreg[147]), .B(n1017), .Z(n1021) );
  NAND U1133 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U1134 ( .A(n1021), .B(n1020), .Z(n1059) );
  XNOR U1135 ( .A(n1060), .B(n1059), .Z(c[148]) );
  NANDN U1136 ( .A(n1023), .B(n1022), .Z(n1027) );
  NANDN U1137 ( .A(n1025), .B(n1024), .Z(n1026) );
  AND U1138 ( .A(n1027), .B(n1026), .Z(n1066) );
  NANDN U1139 ( .A(n1029), .B(n1028), .Z(n1033) );
  NANDN U1140 ( .A(n1031), .B(n1030), .Z(n1032) );
  AND U1141 ( .A(n1033), .B(n1032), .Z(n1064) );
  NANDN U1142 ( .A(n5274), .B(n1034), .Z(n1036) );
  XOR U1143 ( .A(b[7]), .B(a[23]), .Z(n1075) );
  NANDN U1144 ( .A(n5275), .B(n1075), .Z(n1035) );
  AND U1145 ( .A(n1036), .B(n1035), .Z(n1094) );
  NANDN U1146 ( .A(n5176), .B(n1037), .Z(n1039) );
  XOR U1147 ( .A(b[3]), .B(a[27]), .Z(n1078) );
  NANDN U1148 ( .A(n5177), .B(n1078), .Z(n1038) );
  NAND U1149 ( .A(n1039), .B(n1038), .Z(n1093) );
  XNOR U1150 ( .A(n1094), .B(n1093), .Z(n1096) );
  NAND U1151 ( .A(b[0]), .B(a[29]), .Z(n1040) );
  XNOR U1152 ( .A(b[1]), .B(n1040), .Z(n1042) );
  NANDN U1153 ( .A(b[0]), .B(a[28]), .Z(n1041) );
  NAND U1154 ( .A(n1042), .B(n1041), .Z(n1090) );
  NANDN U1155 ( .A(n5249), .B(n1043), .Z(n1045) );
  XOR U1156 ( .A(b[5]), .B(a[25]), .Z(n1084) );
  NANDN U1157 ( .A(n5184), .B(n1084), .Z(n1044) );
  AND U1158 ( .A(n1045), .B(n1044), .Z(n1088) );
  AND U1159 ( .A(b[7]), .B(a[21]), .Z(n1087) );
  XNOR U1160 ( .A(n1088), .B(n1087), .Z(n1089) );
  XNOR U1161 ( .A(n1090), .B(n1089), .Z(n1095) );
  XOR U1162 ( .A(n1096), .B(n1095), .Z(n1070) );
  NANDN U1163 ( .A(n1047), .B(n1046), .Z(n1051) );
  NANDN U1164 ( .A(n1049), .B(n1048), .Z(n1050) );
  AND U1165 ( .A(n1051), .B(n1050), .Z(n1069) );
  XNOR U1166 ( .A(n1070), .B(n1069), .Z(n1071) );
  NANDN U1167 ( .A(n1053), .B(n1052), .Z(n1057) );
  NAND U1168 ( .A(n1055), .B(n1054), .Z(n1056) );
  NAND U1169 ( .A(n1057), .B(n1056), .Z(n1072) );
  XNOR U1170 ( .A(n1071), .B(n1072), .Z(n1063) );
  XNOR U1171 ( .A(n1064), .B(n1063), .Z(n1065) );
  XNOR U1172 ( .A(n1066), .B(n1065), .Z(n1099) );
  XNOR U1173 ( .A(sreg[149]), .B(n1099), .Z(n1101) );
  NANDN U1174 ( .A(sreg[148]), .B(n1058), .Z(n1062) );
  NAND U1175 ( .A(n1060), .B(n1059), .Z(n1061) );
  NAND U1176 ( .A(n1062), .B(n1061), .Z(n1100) );
  XNOR U1177 ( .A(n1101), .B(n1100), .Z(c[149]) );
  NANDN U1178 ( .A(n1064), .B(n1063), .Z(n1068) );
  NANDN U1179 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U1180 ( .A(n1068), .B(n1067), .Z(n1107) );
  NANDN U1181 ( .A(n1070), .B(n1069), .Z(n1074) );
  NANDN U1182 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1183 ( .A(n1074), .B(n1073), .Z(n1105) );
  NANDN U1184 ( .A(n5274), .B(n1075), .Z(n1077) );
  XOR U1185 ( .A(b[7]), .B(a[24]), .Z(n1116) );
  NANDN U1186 ( .A(n5275), .B(n1116), .Z(n1076) );
  AND U1187 ( .A(n1077), .B(n1076), .Z(n1135) );
  NANDN U1188 ( .A(n5176), .B(n1078), .Z(n1080) );
  XOR U1189 ( .A(b[3]), .B(a[28]), .Z(n1119) );
  NANDN U1190 ( .A(n5177), .B(n1119), .Z(n1079) );
  NAND U1191 ( .A(n1080), .B(n1079), .Z(n1134) );
  XNOR U1192 ( .A(n1135), .B(n1134), .Z(n1137) );
  NAND U1193 ( .A(b[0]), .B(a[30]), .Z(n1081) );
  XNOR U1194 ( .A(b[1]), .B(n1081), .Z(n1083) );
  NANDN U1195 ( .A(b[0]), .B(a[29]), .Z(n1082) );
  NAND U1196 ( .A(n1083), .B(n1082), .Z(n1131) );
  NANDN U1197 ( .A(n5249), .B(n1084), .Z(n1086) );
  XOR U1198 ( .A(b[5]), .B(a[26]), .Z(n1125) );
  NANDN U1199 ( .A(n5184), .B(n1125), .Z(n1085) );
  AND U1200 ( .A(n1086), .B(n1085), .Z(n1129) );
  AND U1201 ( .A(b[7]), .B(a[22]), .Z(n1128) );
  XNOR U1202 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1203 ( .A(n1131), .B(n1130), .Z(n1136) );
  XOR U1204 ( .A(n1137), .B(n1136), .Z(n1111) );
  NANDN U1205 ( .A(n1088), .B(n1087), .Z(n1092) );
  NANDN U1206 ( .A(n1090), .B(n1089), .Z(n1091) );
  AND U1207 ( .A(n1092), .B(n1091), .Z(n1110) );
  XNOR U1208 ( .A(n1111), .B(n1110), .Z(n1112) );
  NANDN U1209 ( .A(n1094), .B(n1093), .Z(n1098) );
  NAND U1210 ( .A(n1096), .B(n1095), .Z(n1097) );
  NAND U1211 ( .A(n1098), .B(n1097), .Z(n1113) );
  XNOR U1212 ( .A(n1112), .B(n1113), .Z(n1104) );
  XNOR U1213 ( .A(n1105), .B(n1104), .Z(n1106) );
  XNOR U1214 ( .A(n1107), .B(n1106), .Z(n1140) );
  XNOR U1215 ( .A(sreg[150]), .B(n1140), .Z(n1142) );
  NANDN U1216 ( .A(sreg[149]), .B(n1099), .Z(n1103) );
  NAND U1217 ( .A(n1101), .B(n1100), .Z(n1102) );
  NAND U1218 ( .A(n1103), .B(n1102), .Z(n1141) );
  XNOR U1219 ( .A(n1142), .B(n1141), .Z(c[150]) );
  NANDN U1220 ( .A(n1105), .B(n1104), .Z(n1109) );
  NANDN U1221 ( .A(n1107), .B(n1106), .Z(n1108) );
  AND U1222 ( .A(n1109), .B(n1108), .Z(n1148) );
  NANDN U1223 ( .A(n1111), .B(n1110), .Z(n1115) );
  NANDN U1224 ( .A(n1113), .B(n1112), .Z(n1114) );
  AND U1225 ( .A(n1115), .B(n1114), .Z(n1146) );
  NANDN U1226 ( .A(n5274), .B(n1116), .Z(n1118) );
  XOR U1227 ( .A(b[7]), .B(a[25]), .Z(n1157) );
  NANDN U1228 ( .A(n5275), .B(n1157), .Z(n1117) );
  AND U1229 ( .A(n1118), .B(n1117), .Z(n1176) );
  NANDN U1230 ( .A(n5176), .B(n1119), .Z(n1121) );
  XOR U1231 ( .A(b[3]), .B(a[29]), .Z(n1160) );
  NANDN U1232 ( .A(n5177), .B(n1160), .Z(n1120) );
  NAND U1233 ( .A(n1121), .B(n1120), .Z(n1175) );
  XNOR U1234 ( .A(n1176), .B(n1175), .Z(n1178) );
  NAND U1235 ( .A(b[0]), .B(a[31]), .Z(n1122) );
  XNOR U1236 ( .A(b[1]), .B(n1122), .Z(n1124) );
  NANDN U1237 ( .A(b[0]), .B(a[30]), .Z(n1123) );
  NAND U1238 ( .A(n1124), .B(n1123), .Z(n1172) );
  NANDN U1239 ( .A(n5249), .B(n1125), .Z(n1127) );
  XOR U1240 ( .A(b[5]), .B(a[27]), .Z(n1163) );
  NANDN U1241 ( .A(n5184), .B(n1163), .Z(n1126) );
  AND U1242 ( .A(n1127), .B(n1126), .Z(n1170) );
  AND U1243 ( .A(b[7]), .B(a[23]), .Z(n1169) );
  XNOR U1244 ( .A(n1170), .B(n1169), .Z(n1171) );
  XNOR U1245 ( .A(n1172), .B(n1171), .Z(n1177) );
  XOR U1246 ( .A(n1178), .B(n1177), .Z(n1152) );
  NANDN U1247 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U1248 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1249 ( .A(n1133), .B(n1132), .Z(n1151) );
  XNOR U1250 ( .A(n1152), .B(n1151), .Z(n1153) );
  NANDN U1251 ( .A(n1135), .B(n1134), .Z(n1139) );
  NAND U1252 ( .A(n1137), .B(n1136), .Z(n1138) );
  NAND U1253 ( .A(n1139), .B(n1138), .Z(n1154) );
  XNOR U1254 ( .A(n1153), .B(n1154), .Z(n1145) );
  XNOR U1255 ( .A(n1146), .B(n1145), .Z(n1147) );
  XNOR U1256 ( .A(n1148), .B(n1147), .Z(n1181) );
  XNOR U1257 ( .A(sreg[151]), .B(n1181), .Z(n1183) );
  NANDN U1258 ( .A(sreg[150]), .B(n1140), .Z(n1144) );
  NAND U1259 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1260 ( .A(n1144), .B(n1143), .Z(n1182) );
  XNOR U1261 ( .A(n1183), .B(n1182), .Z(c[151]) );
  NANDN U1262 ( .A(n1146), .B(n1145), .Z(n1150) );
  NANDN U1263 ( .A(n1148), .B(n1147), .Z(n1149) );
  AND U1264 ( .A(n1150), .B(n1149), .Z(n1189) );
  NANDN U1265 ( .A(n1152), .B(n1151), .Z(n1156) );
  NANDN U1266 ( .A(n1154), .B(n1153), .Z(n1155) );
  AND U1267 ( .A(n1156), .B(n1155), .Z(n1187) );
  NANDN U1268 ( .A(n5274), .B(n1157), .Z(n1159) );
  XOR U1269 ( .A(b[7]), .B(a[26]), .Z(n1198) );
  NANDN U1270 ( .A(n5275), .B(n1198), .Z(n1158) );
  AND U1271 ( .A(n1159), .B(n1158), .Z(n1217) );
  NANDN U1272 ( .A(n5176), .B(n1160), .Z(n1162) );
  XOR U1273 ( .A(b[3]), .B(a[30]), .Z(n1201) );
  NANDN U1274 ( .A(n5177), .B(n1201), .Z(n1161) );
  NAND U1275 ( .A(n1162), .B(n1161), .Z(n1216) );
  XNOR U1276 ( .A(n1217), .B(n1216), .Z(n1219) );
  NANDN U1277 ( .A(n5249), .B(n1163), .Z(n1165) );
  XOR U1278 ( .A(b[5]), .B(a[28]), .Z(n1207) );
  NANDN U1279 ( .A(n5184), .B(n1207), .Z(n1164) );
  AND U1280 ( .A(n1165), .B(n1164), .Z(n1211) );
  AND U1281 ( .A(b[7]), .B(a[24]), .Z(n1210) );
  XNOR U1282 ( .A(n1211), .B(n1210), .Z(n1212) );
  NAND U1283 ( .A(b[0]), .B(a[32]), .Z(n1166) );
  XNOR U1284 ( .A(b[1]), .B(n1166), .Z(n1168) );
  NANDN U1285 ( .A(b[0]), .B(a[31]), .Z(n1167) );
  NAND U1286 ( .A(n1168), .B(n1167), .Z(n1213) );
  XNOR U1287 ( .A(n1212), .B(n1213), .Z(n1218) );
  XOR U1288 ( .A(n1219), .B(n1218), .Z(n1193) );
  NANDN U1289 ( .A(n1170), .B(n1169), .Z(n1174) );
  NANDN U1290 ( .A(n1172), .B(n1171), .Z(n1173) );
  AND U1291 ( .A(n1174), .B(n1173), .Z(n1192) );
  XNOR U1292 ( .A(n1193), .B(n1192), .Z(n1194) );
  NANDN U1293 ( .A(n1176), .B(n1175), .Z(n1180) );
  NAND U1294 ( .A(n1178), .B(n1177), .Z(n1179) );
  NAND U1295 ( .A(n1180), .B(n1179), .Z(n1195) );
  XNOR U1296 ( .A(n1194), .B(n1195), .Z(n1186) );
  XNOR U1297 ( .A(n1187), .B(n1186), .Z(n1188) );
  XNOR U1298 ( .A(n1189), .B(n1188), .Z(n1222) );
  XNOR U1299 ( .A(sreg[152]), .B(n1222), .Z(n1224) );
  NANDN U1300 ( .A(sreg[151]), .B(n1181), .Z(n1185) );
  NAND U1301 ( .A(n1183), .B(n1182), .Z(n1184) );
  NAND U1302 ( .A(n1185), .B(n1184), .Z(n1223) );
  XNOR U1303 ( .A(n1224), .B(n1223), .Z(c[152]) );
  NANDN U1304 ( .A(n1187), .B(n1186), .Z(n1191) );
  NANDN U1305 ( .A(n1189), .B(n1188), .Z(n1190) );
  AND U1306 ( .A(n1191), .B(n1190), .Z(n1230) );
  NANDN U1307 ( .A(n1193), .B(n1192), .Z(n1197) );
  NANDN U1308 ( .A(n1195), .B(n1194), .Z(n1196) );
  AND U1309 ( .A(n1197), .B(n1196), .Z(n1228) );
  NANDN U1310 ( .A(n5274), .B(n1198), .Z(n1200) );
  XOR U1311 ( .A(b[7]), .B(a[27]), .Z(n1239) );
  NANDN U1312 ( .A(n5275), .B(n1239), .Z(n1199) );
  AND U1313 ( .A(n1200), .B(n1199), .Z(n1258) );
  NANDN U1314 ( .A(n5176), .B(n1201), .Z(n1203) );
  XOR U1315 ( .A(b[3]), .B(a[31]), .Z(n1242) );
  NANDN U1316 ( .A(n5177), .B(n1242), .Z(n1202) );
  NAND U1317 ( .A(n1203), .B(n1202), .Z(n1257) );
  XNOR U1318 ( .A(n1258), .B(n1257), .Z(n1260) );
  NAND U1319 ( .A(b[0]), .B(a[33]), .Z(n1204) );
  XNOR U1320 ( .A(b[1]), .B(n1204), .Z(n1206) );
  NANDN U1321 ( .A(b[0]), .B(a[32]), .Z(n1205) );
  NAND U1322 ( .A(n1206), .B(n1205), .Z(n1254) );
  NANDN U1323 ( .A(n5249), .B(n1207), .Z(n1209) );
  XOR U1324 ( .A(b[5]), .B(a[29]), .Z(n1248) );
  NANDN U1325 ( .A(n5184), .B(n1248), .Z(n1208) );
  AND U1326 ( .A(n1209), .B(n1208), .Z(n1252) );
  AND U1327 ( .A(b[7]), .B(a[25]), .Z(n1251) );
  XNOR U1328 ( .A(n1252), .B(n1251), .Z(n1253) );
  XNOR U1329 ( .A(n1254), .B(n1253), .Z(n1259) );
  XOR U1330 ( .A(n1260), .B(n1259), .Z(n1234) );
  NANDN U1331 ( .A(n1211), .B(n1210), .Z(n1215) );
  NANDN U1332 ( .A(n1213), .B(n1212), .Z(n1214) );
  AND U1333 ( .A(n1215), .B(n1214), .Z(n1233) );
  XNOR U1334 ( .A(n1234), .B(n1233), .Z(n1235) );
  NANDN U1335 ( .A(n1217), .B(n1216), .Z(n1221) );
  NAND U1336 ( .A(n1219), .B(n1218), .Z(n1220) );
  NAND U1337 ( .A(n1221), .B(n1220), .Z(n1236) );
  XNOR U1338 ( .A(n1235), .B(n1236), .Z(n1227) );
  XNOR U1339 ( .A(n1228), .B(n1227), .Z(n1229) );
  XNOR U1340 ( .A(n1230), .B(n1229), .Z(n1263) );
  XNOR U1341 ( .A(sreg[153]), .B(n1263), .Z(n1265) );
  NANDN U1342 ( .A(sreg[152]), .B(n1222), .Z(n1226) );
  NAND U1343 ( .A(n1224), .B(n1223), .Z(n1225) );
  NAND U1344 ( .A(n1226), .B(n1225), .Z(n1264) );
  XNOR U1345 ( .A(n1265), .B(n1264), .Z(c[153]) );
  NANDN U1346 ( .A(n1228), .B(n1227), .Z(n1232) );
  NANDN U1347 ( .A(n1230), .B(n1229), .Z(n1231) );
  AND U1348 ( .A(n1232), .B(n1231), .Z(n1271) );
  NANDN U1349 ( .A(n1234), .B(n1233), .Z(n1238) );
  NANDN U1350 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1351 ( .A(n1238), .B(n1237), .Z(n1269) );
  NANDN U1352 ( .A(n5274), .B(n1239), .Z(n1241) );
  XOR U1353 ( .A(b[7]), .B(a[28]), .Z(n1280) );
  NANDN U1354 ( .A(n5275), .B(n1280), .Z(n1240) );
  AND U1355 ( .A(n1241), .B(n1240), .Z(n1299) );
  NANDN U1356 ( .A(n5176), .B(n1242), .Z(n1244) );
  XOR U1357 ( .A(b[3]), .B(a[32]), .Z(n1283) );
  NANDN U1358 ( .A(n5177), .B(n1283), .Z(n1243) );
  NAND U1359 ( .A(n1244), .B(n1243), .Z(n1298) );
  XNOR U1360 ( .A(n1299), .B(n1298), .Z(n1301) );
  NAND U1361 ( .A(b[0]), .B(a[34]), .Z(n1245) );
  XNOR U1362 ( .A(b[1]), .B(n1245), .Z(n1247) );
  NANDN U1363 ( .A(b[0]), .B(a[33]), .Z(n1246) );
  NAND U1364 ( .A(n1247), .B(n1246), .Z(n1295) );
  NANDN U1365 ( .A(n5249), .B(n1248), .Z(n1250) );
  XOR U1366 ( .A(b[5]), .B(a[30]), .Z(n1289) );
  NANDN U1367 ( .A(n5184), .B(n1289), .Z(n1249) );
  AND U1368 ( .A(n1250), .B(n1249), .Z(n1293) );
  AND U1369 ( .A(b[7]), .B(a[26]), .Z(n1292) );
  XNOR U1370 ( .A(n1293), .B(n1292), .Z(n1294) );
  XNOR U1371 ( .A(n1295), .B(n1294), .Z(n1300) );
  XOR U1372 ( .A(n1301), .B(n1300), .Z(n1275) );
  NANDN U1373 ( .A(n1252), .B(n1251), .Z(n1256) );
  NANDN U1374 ( .A(n1254), .B(n1253), .Z(n1255) );
  AND U1375 ( .A(n1256), .B(n1255), .Z(n1274) );
  XNOR U1376 ( .A(n1275), .B(n1274), .Z(n1276) );
  NANDN U1377 ( .A(n1258), .B(n1257), .Z(n1262) );
  NAND U1378 ( .A(n1260), .B(n1259), .Z(n1261) );
  NAND U1379 ( .A(n1262), .B(n1261), .Z(n1277) );
  XNOR U1380 ( .A(n1276), .B(n1277), .Z(n1268) );
  XNOR U1381 ( .A(n1269), .B(n1268), .Z(n1270) );
  XNOR U1382 ( .A(n1271), .B(n1270), .Z(n1304) );
  XNOR U1383 ( .A(sreg[154]), .B(n1304), .Z(n1306) );
  NANDN U1384 ( .A(sreg[153]), .B(n1263), .Z(n1267) );
  NAND U1385 ( .A(n1265), .B(n1264), .Z(n1266) );
  NAND U1386 ( .A(n1267), .B(n1266), .Z(n1305) );
  XNOR U1387 ( .A(n1306), .B(n1305), .Z(c[154]) );
  NANDN U1388 ( .A(n1269), .B(n1268), .Z(n1273) );
  NANDN U1389 ( .A(n1271), .B(n1270), .Z(n1272) );
  AND U1390 ( .A(n1273), .B(n1272), .Z(n1312) );
  NANDN U1391 ( .A(n1275), .B(n1274), .Z(n1279) );
  NANDN U1392 ( .A(n1277), .B(n1276), .Z(n1278) );
  AND U1393 ( .A(n1279), .B(n1278), .Z(n1310) );
  NANDN U1394 ( .A(n5274), .B(n1280), .Z(n1282) );
  XOR U1395 ( .A(b[7]), .B(a[29]), .Z(n1321) );
  NANDN U1396 ( .A(n5275), .B(n1321), .Z(n1281) );
  AND U1397 ( .A(n1282), .B(n1281), .Z(n1340) );
  NANDN U1398 ( .A(n5176), .B(n1283), .Z(n1285) );
  XOR U1399 ( .A(b[3]), .B(a[33]), .Z(n1324) );
  NANDN U1400 ( .A(n5177), .B(n1324), .Z(n1284) );
  NAND U1401 ( .A(n1285), .B(n1284), .Z(n1339) );
  XNOR U1402 ( .A(n1340), .B(n1339), .Z(n1342) );
  NAND U1403 ( .A(b[0]), .B(a[35]), .Z(n1286) );
  XNOR U1404 ( .A(b[1]), .B(n1286), .Z(n1288) );
  NANDN U1405 ( .A(b[0]), .B(a[34]), .Z(n1287) );
  NAND U1406 ( .A(n1288), .B(n1287), .Z(n1336) );
  NANDN U1407 ( .A(n5249), .B(n1289), .Z(n1291) );
  XOR U1408 ( .A(b[5]), .B(a[31]), .Z(n1330) );
  NANDN U1409 ( .A(n5184), .B(n1330), .Z(n1290) );
  AND U1410 ( .A(n1291), .B(n1290), .Z(n1334) );
  AND U1411 ( .A(b[7]), .B(a[27]), .Z(n1333) );
  XNOR U1412 ( .A(n1334), .B(n1333), .Z(n1335) );
  XNOR U1413 ( .A(n1336), .B(n1335), .Z(n1341) );
  XOR U1414 ( .A(n1342), .B(n1341), .Z(n1316) );
  NANDN U1415 ( .A(n1293), .B(n1292), .Z(n1297) );
  NANDN U1416 ( .A(n1295), .B(n1294), .Z(n1296) );
  AND U1417 ( .A(n1297), .B(n1296), .Z(n1315) );
  XNOR U1418 ( .A(n1316), .B(n1315), .Z(n1317) );
  NANDN U1419 ( .A(n1299), .B(n1298), .Z(n1303) );
  NAND U1420 ( .A(n1301), .B(n1300), .Z(n1302) );
  NAND U1421 ( .A(n1303), .B(n1302), .Z(n1318) );
  XNOR U1422 ( .A(n1317), .B(n1318), .Z(n1309) );
  XNOR U1423 ( .A(n1310), .B(n1309), .Z(n1311) );
  XNOR U1424 ( .A(n1312), .B(n1311), .Z(n1345) );
  XNOR U1425 ( .A(sreg[155]), .B(n1345), .Z(n1347) );
  NANDN U1426 ( .A(sreg[154]), .B(n1304), .Z(n1308) );
  NAND U1427 ( .A(n1306), .B(n1305), .Z(n1307) );
  NAND U1428 ( .A(n1308), .B(n1307), .Z(n1346) );
  XNOR U1429 ( .A(n1347), .B(n1346), .Z(c[155]) );
  NANDN U1430 ( .A(n1310), .B(n1309), .Z(n1314) );
  NANDN U1431 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U1432 ( .A(n1314), .B(n1313), .Z(n1353) );
  NANDN U1433 ( .A(n1316), .B(n1315), .Z(n1320) );
  NANDN U1434 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U1435 ( .A(n1320), .B(n1319), .Z(n1351) );
  NANDN U1436 ( .A(n5274), .B(n1321), .Z(n1323) );
  XOR U1437 ( .A(b[7]), .B(a[30]), .Z(n1362) );
  NANDN U1438 ( .A(n5275), .B(n1362), .Z(n1322) );
  AND U1439 ( .A(n1323), .B(n1322), .Z(n1381) );
  NANDN U1440 ( .A(n5176), .B(n1324), .Z(n1326) );
  XOR U1441 ( .A(b[3]), .B(a[34]), .Z(n1365) );
  NANDN U1442 ( .A(n5177), .B(n1365), .Z(n1325) );
  NAND U1443 ( .A(n1326), .B(n1325), .Z(n1380) );
  XNOR U1444 ( .A(n1381), .B(n1380), .Z(n1383) );
  NAND U1445 ( .A(b[0]), .B(a[36]), .Z(n1327) );
  XNOR U1446 ( .A(b[1]), .B(n1327), .Z(n1329) );
  NANDN U1447 ( .A(b[0]), .B(a[35]), .Z(n1328) );
  NAND U1448 ( .A(n1329), .B(n1328), .Z(n1377) );
  NANDN U1449 ( .A(n5249), .B(n1330), .Z(n1332) );
  XOR U1450 ( .A(b[5]), .B(a[32]), .Z(n1371) );
  NANDN U1451 ( .A(n5184), .B(n1371), .Z(n1331) );
  AND U1452 ( .A(n1332), .B(n1331), .Z(n1375) );
  AND U1453 ( .A(b[7]), .B(a[28]), .Z(n1374) );
  XNOR U1454 ( .A(n1375), .B(n1374), .Z(n1376) );
  XNOR U1455 ( .A(n1377), .B(n1376), .Z(n1382) );
  XOR U1456 ( .A(n1383), .B(n1382), .Z(n1357) );
  NANDN U1457 ( .A(n1334), .B(n1333), .Z(n1338) );
  NANDN U1458 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U1459 ( .A(n1338), .B(n1337), .Z(n1356) );
  XNOR U1460 ( .A(n1357), .B(n1356), .Z(n1358) );
  NANDN U1461 ( .A(n1340), .B(n1339), .Z(n1344) );
  NAND U1462 ( .A(n1342), .B(n1341), .Z(n1343) );
  NAND U1463 ( .A(n1344), .B(n1343), .Z(n1359) );
  XNOR U1464 ( .A(n1358), .B(n1359), .Z(n1350) );
  XNOR U1465 ( .A(n1351), .B(n1350), .Z(n1352) );
  XNOR U1466 ( .A(n1353), .B(n1352), .Z(n1386) );
  XNOR U1467 ( .A(sreg[156]), .B(n1386), .Z(n1388) );
  NANDN U1468 ( .A(sreg[155]), .B(n1345), .Z(n1349) );
  NAND U1469 ( .A(n1347), .B(n1346), .Z(n1348) );
  NAND U1470 ( .A(n1349), .B(n1348), .Z(n1387) );
  XNOR U1471 ( .A(n1388), .B(n1387), .Z(c[156]) );
  NANDN U1472 ( .A(n1351), .B(n1350), .Z(n1355) );
  NANDN U1473 ( .A(n1353), .B(n1352), .Z(n1354) );
  AND U1474 ( .A(n1355), .B(n1354), .Z(n1394) );
  NANDN U1475 ( .A(n1357), .B(n1356), .Z(n1361) );
  NANDN U1476 ( .A(n1359), .B(n1358), .Z(n1360) );
  AND U1477 ( .A(n1361), .B(n1360), .Z(n1392) );
  NANDN U1478 ( .A(n5274), .B(n1362), .Z(n1364) );
  XOR U1479 ( .A(b[7]), .B(a[31]), .Z(n1403) );
  NANDN U1480 ( .A(n5275), .B(n1403), .Z(n1363) );
  AND U1481 ( .A(n1364), .B(n1363), .Z(n1422) );
  NANDN U1482 ( .A(n5176), .B(n1365), .Z(n1367) );
  XOR U1483 ( .A(b[3]), .B(a[35]), .Z(n1406) );
  NANDN U1484 ( .A(n5177), .B(n1406), .Z(n1366) );
  NAND U1485 ( .A(n1367), .B(n1366), .Z(n1421) );
  XNOR U1486 ( .A(n1422), .B(n1421), .Z(n1424) );
  NAND U1487 ( .A(b[0]), .B(a[37]), .Z(n1368) );
  XNOR U1488 ( .A(b[1]), .B(n1368), .Z(n1370) );
  NANDN U1489 ( .A(b[0]), .B(a[36]), .Z(n1369) );
  NAND U1490 ( .A(n1370), .B(n1369), .Z(n1418) );
  NANDN U1491 ( .A(n5249), .B(n1371), .Z(n1373) );
  XOR U1492 ( .A(b[5]), .B(a[33]), .Z(n1409) );
  NANDN U1493 ( .A(n5184), .B(n1409), .Z(n1372) );
  AND U1494 ( .A(n1373), .B(n1372), .Z(n1416) );
  AND U1495 ( .A(b[7]), .B(a[29]), .Z(n1415) );
  XNOR U1496 ( .A(n1416), .B(n1415), .Z(n1417) );
  XNOR U1497 ( .A(n1418), .B(n1417), .Z(n1423) );
  XOR U1498 ( .A(n1424), .B(n1423), .Z(n1398) );
  NANDN U1499 ( .A(n1375), .B(n1374), .Z(n1379) );
  NANDN U1500 ( .A(n1377), .B(n1376), .Z(n1378) );
  AND U1501 ( .A(n1379), .B(n1378), .Z(n1397) );
  XNOR U1502 ( .A(n1398), .B(n1397), .Z(n1399) );
  NANDN U1503 ( .A(n1381), .B(n1380), .Z(n1385) );
  NAND U1504 ( .A(n1383), .B(n1382), .Z(n1384) );
  NAND U1505 ( .A(n1385), .B(n1384), .Z(n1400) );
  XNOR U1506 ( .A(n1399), .B(n1400), .Z(n1391) );
  XNOR U1507 ( .A(n1392), .B(n1391), .Z(n1393) );
  XNOR U1508 ( .A(n1394), .B(n1393), .Z(n1427) );
  XNOR U1509 ( .A(sreg[157]), .B(n1427), .Z(n1429) );
  NANDN U1510 ( .A(sreg[156]), .B(n1386), .Z(n1390) );
  NAND U1511 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1512 ( .A(n1390), .B(n1389), .Z(n1428) );
  XNOR U1513 ( .A(n1429), .B(n1428), .Z(c[157]) );
  NANDN U1514 ( .A(n1392), .B(n1391), .Z(n1396) );
  NANDN U1515 ( .A(n1394), .B(n1393), .Z(n1395) );
  AND U1516 ( .A(n1396), .B(n1395), .Z(n1435) );
  NANDN U1517 ( .A(n1398), .B(n1397), .Z(n1402) );
  NANDN U1518 ( .A(n1400), .B(n1399), .Z(n1401) );
  AND U1519 ( .A(n1402), .B(n1401), .Z(n1433) );
  NANDN U1520 ( .A(n5274), .B(n1403), .Z(n1405) );
  XOR U1521 ( .A(b[7]), .B(a[32]), .Z(n1444) );
  NANDN U1522 ( .A(n5275), .B(n1444), .Z(n1404) );
  AND U1523 ( .A(n1405), .B(n1404), .Z(n1463) );
  NANDN U1524 ( .A(n5176), .B(n1406), .Z(n1408) );
  XOR U1525 ( .A(b[3]), .B(a[36]), .Z(n1447) );
  NANDN U1526 ( .A(n5177), .B(n1447), .Z(n1407) );
  NAND U1527 ( .A(n1408), .B(n1407), .Z(n1462) );
  XNOR U1528 ( .A(n1463), .B(n1462), .Z(n1465) );
  NANDN U1529 ( .A(n5249), .B(n1409), .Z(n1411) );
  XOR U1530 ( .A(b[5]), .B(a[34]), .Z(n1453) );
  NANDN U1531 ( .A(n5184), .B(n1453), .Z(n1410) );
  AND U1532 ( .A(n1411), .B(n1410), .Z(n1457) );
  AND U1533 ( .A(b[7]), .B(a[30]), .Z(n1456) );
  XNOR U1534 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U1535 ( .A(b[0]), .B(a[38]), .Z(n1412) );
  XNOR U1536 ( .A(b[1]), .B(n1412), .Z(n1414) );
  NANDN U1537 ( .A(b[0]), .B(a[37]), .Z(n1413) );
  NAND U1538 ( .A(n1414), .B(n1413), .Z(n1459) );
  XNOR U1539 ( .A(n1458), .B(n1459), .Z(n1464) );
  XOR U1540 ( .A(n1465), .B(n1464), .Z(n1439) );
  NANDN U1541 ( .A(n1416), .B(n1415), .Z(n1420) );
  NANDN U1542 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U1543 ( .A(n1420), .B(n1419), .Z(n1438) );
  XNOR U1544 ( .A(n1439), .B(n1438), .Z(n1440) );
  NANDN U1545 ( .A(n1422), .B(n1421), .Z(n1426) );
  NAND U1546 ( .A(n1424), .B(n1423), .Z(n1425) );
  NAND U1547 ( .A(n1426), .B(n1425), .Z(n1441) );
  XNOR U1548 ( .A(n1440), .B(n1441), .Z(n1432) );
  XNOR U1549 ( .A(n1433), .B(n1432), .Z(n1434) );
  XNOR U1550 ( .A(n1435), .B(n1434), .Z(n1468) );
  XNOR U1551 ( .A(sreg[158]), .B(n1468), .Z(n1470) );
  NANDN U1552 ( .A(sreg[157]), .B(n1427), .Z(n1431) );
  NAND U1553 ( .A(n1429), .B(n1428), .Z(n1430) );
  NAND U1554 ( .A(n1431), .B(n1430), .Z(n1469) );
  XNOR U1555 ( .A(n1470), .B(n1469), .Z(c[158]) );
  NANDN U1556 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1557 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1558 ( .A(n1437), .B(n1436), .Z(n1476) );
  NANDN U1559 ( .A(n1439), .B(n1438), .Z(n1443) );
  NANDN U1560 ( .A(n1441), .B(n1440), .Z(n1442) );
  AND U1561 ( .A(n1443), .B(n1442), .Z(n1474) );
  NANDN U1562 ( .A(n5274), .B(n1444), .Z(n1446) );
  XOR U1563 ( .A(b[7]), .B(a[33]), .Z(n1485) );
  NANDN U1564 ( .A(n5275), .B(n1485), .Z(n1445) );
  AND U1565 ( .A(n1446), .B(n1445), .Z(n1504) );
  NANDN U1566 ( .A(n5176), .B(n1447), .Z(n1449) );
  XOR U1567 ( .A(b[3]), .B(a[37]), .Z(n1488) );
  NANDN U1568 ( .A(n5177), .B(n1488), .Z(n1448) );
  NAND U1569 ( .A(n1449), .B(n1448), .Z(n1503) );
  XNOR U1570 ( .A(n1504), .B(n1503), .Z(n1506) );
  NAND U1571 ( .A(b[0]), .B(a[39]), .Z(n1450) );
  XNOR U1572 ( .A(b[1]), .B(n1450), .Z(n1452) );
  NANDN U1573 ( .A(b[0]), .B(a[38]), .Z(n1451) );
  NAND U1574 ( .A(n1452), .B(n1451), .Z(n1500) );
  NANDN U1575 ( .A(n5249), .B(n1453), .Z(n1455) );
  XOR U1576 ( .A(b[5]), .B(a[35]), .Z(n1491) );
  NANDN U1577 ( .A(n5184), .B(n1491), .Z(n1454) );
  AND U1578 ( .A(n1455), .B(n1454), .Z(n1498) );
  AND U1579 ( .A(b[7]), .B(a[31]), .Z(n1497) );
  XNOR U1580 ( .A(n1498), .B(n1497), .Z(n1499) );
  XNOR U1581 ( .A(n1500), .B(n1499), .Z(n1505) );
  XOR U1582 ( .A(n1506), .B(n1505), .Z(n1480) );
  NANDN U1583 ( .A(n1457), .B(n1456), .Z(n1461) );
  NANDN U1584 ( .A(n1459), .B(n1458), .Z(n1460) );
  AND U1585 ( .A(n1461), .B(n1460), .Z(n1479) );
  XNOR U1586 ( .A(n1480), .B(n1479), .Z(n1481) );
  NANDN U1587 ( .A(n1463), .B(n1462), .Z(n1467) );
  NAND U1588 ( .A(n1465), .B(n1464), .Z(n1466) );
  NAND U1589 ( .A(n1467), .B(n1466), .Z(n1482) );
  XNOR U1590 ( .A(n1481), .B(n1482), .Z(n1473) );
  XNOR U1591 ( .A(n1474), .B(n1473), .Z(n1475) );
  XNOR U1592 ( .A(n1476), .B(n1475), .Z(n1509) );
  XNOR U1593 ( .A(sreg[159]), .B(n1509), .Z(n1511) );
  NANDN U1594 ( .A(sreg[158]), .B(n1468), .Z(n1472) );
  NAND U1595 ( .A(n1470), .B(n1469), .Z(n1471) );
  NAND U1596 ( .A(n1472), .B(n1471), .Z(n1510) );
  XNOR U1597 ( .A(n1511), .B(n1510), .Z(c[159]) );
  NANDN U1598 ( .A(n1474), .B(n1473), .Z(n1478) );
  NANDN U1599 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U1600 ( .A(n1478), .B(n1477), .Z(n1517) );
  NANDN U1601 ( .A(n1480), .B(n1479), .Z(n1484) );
  NANDN U1602 ( .A(n1482), .B(n1481), .Z(n1483) );
  AND U1603 ( .A(n1484), .B(n1483), .Z(n1515) );
  NANDN U1604 ( .A(n5274), .B(n1485), .Z(n1487) );
  XOR U1605 ( .A(b[7]), .B(a[34]), .Z(n1526) );
  NANDN U1606 ( .A(n5275), .B(n1526), .Z(n1486) );
  AND U1607 ( .A(n1487), .B(n1486), .Z(n1545) );
  NANDN U1608 ( .A(n5176), .B(n1488), .Z(n1490) );
  XOR U1609 ( .A(b[3]), .B(a[38]), .Z(n1529) );
  NANDN U1610 ( .A(n5177), .B(n1529), .Z(n1489) );
  NAND U1611 ( .A(n1490), .B(n1489), .Z(n1544) );
  XNOR U1612 ( .A(n1545), .B(n1544), .Z(n1547) );
  NANDN U1613 ( .A(n5249), .B(n1491), .Z(n1493) );
  XOR U1614 ( .A(b[5]), .B(a[36]), .Z(n1535) );
  NANDN U1615 ( .A(n5184), .B(n1535), .Z(n1492) );
  AND U1616 ( .A(n1493), .B(n1492), .Z(n1539) );
  AND U1617 ( .A(b[7]), .B(a[32]), .Z(n1538) );
  XNOR U1618 ( .A(n1539), .B(n1538), .Z(n1540) );
  NAND U1619 ( .A(b[0]), .B(a[40]), .Z(n1494) );
  XNOR U1620 ( .A(b[1]), .B(n1494), .Z(n1496) );
  NANDN U1621 ( .A(b[0]), .B(a[39]), .Z(n1495) );
  NAND U1622 ( .A(n1496), .B(n1495), .Z(n1541) );
  XNOR U1623 ( .A(n1540), .B(n1541), .Z(n1546) );
  XOR U1624 ( .A(n1547), .B(n1546), .Z(n1521) );
  NANDN U1625 ( .A(n1498), .B(n1497), .Z(n1502) );
  NANDN U1626 ( .A(n1500), .B(n1499), .Z(n1501) );
  AND U1627 ( .A(n1502), .B(n1501), .Z(n1520) );
  XNOR U1628 ( .A(n1521), .B(n1520), .Z(n1522) );
  NANDN U1629 ( .A(n1504), .B(n1503), .Z(n1508) );
  NAND U1630 ( .A(n1506), .B(n1505), .Z(n1507) );
  NAND U1631 ( .A(n1508), .B(n1507), .Z(n1523) );
  XNOR U1632 ( .A(n1522), .B(n1523), .Z(n1514) );
  XNOR U1633 ( .A(n1515), .B(n1514), .Z(n1516) );
  XNOR U1634 ( .A(n1517), .B(n1516), .Z(n1550) );
  XNOR U1635 ( .A(sreg[160]), .B(n1550), .Z(n1552) );
  NANDN U1636 ( .A(sreg[159]), .B(n1509), .Z(n1513) );
  NAND U1637 ( .A(n1511), .B(n1510), .Z(n1512) );
  NAND U1638 ( .A(n1513), .B(n1512), .Z(n1551) );
  XNOR U1639 ( .A(n1552), .B(n1551), .Z(c[160]) );
  NANDN U1640 ( .A(n1515), .B(n1514), .Z(n1519) );
  NANDN U1641 ( .A(n1517), .B(n1516), .Z(n1518) );
  AND U1642 ( .A(n1519), .B(n1518), .Z(n1558) );
  NANDN U1643 ( .A(n1521), .B(n1520), .Z(n1525) );
  NANDN U1644 ( .A(n1523), .B(n1522), .Z(n1524) );
  AND U1645 ( .A(n1525), .B(n1524), .Z(n1556) );
  NANDN U1646 ( .A(n5274), .B(n1526), .Z(n1528) );
  XOR U1647 ( .A(b[7]), .B(a[35]), .Z(n1567) );
  NANDN U1648 ( .A(n5275), .B(n1567), .Z(n1527) );
  AND U1649 ( .A(n1528), .B(n1527), .Z(n1586) );
  NANDN U1650 ( .A(n5176), .B(n1529), .Z(n1531) );
  XOR U1651 ( .A(b[3]), .B(a[39]), .Z(n1570) );
  NANDN U1652 ( .A(n5177), .B(n1570), .Z(n1530) );
  NAND U1653 ( .A(n1531), .B(n1530), .Z(n1585) );
  XNOR U1654 ( .A(n1586), .B(n1585), .Z(n1588) );
  NAND U1655 ( .A(b[0]), .B(a[41]), .Z(n1532) );
  XNOR U1656 ( .A(b[1]), .B(n1532), .Z(n1534) );
  NANDN U1657 ( .A(b[0]), .B(a[40]), .Z(n1533) );
  NAND U1658 ( .A(n1534), .B(n1533), .Z(n1582) );
  NANDN U1659 ( .A(n5249), .B(n1535), .Z(n1537) );
  XOR U1660 ( .A(b[5]), .B(a[37]), .Z(n1576) );
  NANDN U1661 ( .A(n5184), .B(n1576), .Z(n1536) );
  AND U1662 ( .A(n1537), .B(n1536), .Z(n1580) );
  AND U1663 ( .A(b[7]), .B(a[33]), .Z(n1579) );
  XNOR U1664 ( .A(n1580), .B(n1579), .Z(n1581) );
  XNOR U1665 ( .A(n1582), .B(n1581), .Z(n1587) );
  XOR U1666 ( .A(n1588), .B(n1587), .Z(n1562) );
  NANDN U1667 ( .A(n1539), .B(n1538), .Z(n1543) );
  NANDN U1668 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1669 ( .A(n1543), .B(n1542), .Z(n1561) );
  XNOR U1670 ( .A(n1562), .B(n1561), .Z(n1563) );
  NANDN U1671 ( .A(n1545), .B(n1544), .Z(n1549) );
  NAND U1672 ( .A(n1547), .B(n1546), .Z(n1548) );
  NAND U1673 ( .A(n1549), .B(n1548), .Z(n1564) );
  XNOR U1674 ( .A(n1563), .B(n1564), .Z(n1555) );
  XNOR U1675 ( .A(n1556), .B(n1555), .Z(n1557) );
  XNOR U1676 ( .A(n1558), .B(n1557), .Z(n1591) );
  XNOR U1677 ( .A(sreg[161]), .B(n1591), .Z(n1593) );
  NANDN U1678 ( .A(sreg[160]), .B(n1550), .Z(n1554) );
  NAND U1679 ( .A(n1552), .B(n1551), .Z(n1553) );
  NAND U1680 ( .A(n1554), .B(n1553), .Z(n1592) );
  XNOR U1681 ( .A(n1593), .B(n1592), .Z(c[161]) );
  NANDN U1682 ( .A(n1556), .B(n1555), .Z(n1560) );
  NANDN U1683 ( .A(n1558), .B(n1557), .Z(n1559) );
  AND U1684 ( .A(n1560), .B(n1559), .Z(n1599) );
  NANDN U1685 ( .A(n1562), .B(n1561), .Z(n1566) );
  NANDN U1686 ( .A(n1564), .B(n1563), .Z(n1565) );
  AND U1687 ( .A(n1566), .B(n1565), .Z(n1597) );
  NANDN U1688 ( .A(n5274), .B(n1567), .Z(n1569) );
  XOR U1689 ( .A(b[7]), .B(a[36]), .Z(n1608) );
  NANDN U1690 ( .A(n5275), .B(n1608), .Z(n1568) );
  AND U1691 ( .A(n1569), .B(n1568), .Z(n1627) );
  NANDN U1692 ( .A(n5176), .B(n1570), .Z(n1572) );
  XOR U1693 ( .A(b[3]), .B(a[40]), .Z(n1611) );
  NANDN U1694 ( .A(n5177), .B(n1611), .Z(n1571) );
  NAND U1695 ( .A(n1572), .B(n1571), .Z(n1626) );
  XNOR U1696 ( .A(n1627), .B(n1626), .Z(n1629) );
  NAND U1697 ( .A(b[0]), .B(a[42]), .Z(n1573) );
  XNOR U1698 ( .A(b[1]), .B(n1573), .Z(n1575) );
  NANDN U1699 ( .A(b[0]), .B(a[41]), .Z(n1574) );
  NAND U1700 ( .A(n1575), .B(n1574), .Z(n1623) );
  NANDN U1701 ( .A(n5249), .B(n1576), .Z(n1578) );
  XOR U1702 ( .A(b[5]), .B(a[38]), .Z(n1617) );
  NANDN U1703 ( .A(n5184), .B(n1617), .Z(n1577) );
  AND U1704 ( .A(n1578), .B(n1577), .Z(n1621) );
  AND U1705 ( .A(b[7]), .B(a[34]), .Z(n1620) );
  XNOR U1706 ( .A(n1621), .B(n1620), .Z(n1622) );
  XNOR U1707 ( .A(n1623), .B(n1622), .Z(n1628) );
  XOR U1708 ( .A(n1629), .B(n1628), .Z(n1603) );
  NANDN U1709 ( .A(n1580), .B(n1579), .Z(n1584) );
  NANDN U1710 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U1711 ( .A(n1584), .B(n1583), .Z(n1602) );
  XNOR U1712 ( .A(n1603), .B(n1602), .Z(n1604) );
  NANDN U1713 ( .A(n1586), .B(n1585), .Z(n1590) );
  NAND U1714 ( .A(n1588), .B(n1587), .Z(n1589) );
  NAND U1715 ( .A(n1590), .B(n1589), .Z(n1605) );
  XNOR U1716 ( .A(n1604), .B(n1605), .Z(n1596) );
  XNOR U1717 ( .A(n1597), .B(n1596), .Z(n1598) );
  XNOR U1718 ( .A(n1599), .B(n1598), .Z(n1632) );
  XNOR U1719 ( .A(sreg[162]), .B(n1632), .Z(n1634) );
  NANDN U1720 ( .A(sreg[161]), .B(n1591), .Z(n1595) );
  NAND U1721 ( .A(n1593), .B(n1592), .Z(n1594) );
  NAND U1722 ( .A(n1595), .B(n1594), .Z(n1633) );
  XNOR U1723 ( .A(n1634), .B(n1633), .Z(c[162]) );
  NANDN U1724 ( .A(n1597), .B(n1596), .Z(n1601) );
  NANDN U1725 ( .A(n1599), .B(n1598), .Z(n1600) );
  AND U1726 ( .A(n1601), .B(n1600), .Z(n1640) );
  NANDN U1727 ( .A(n1603), .B(n1602), .Z(n1607) );
  NANDN U1728 ( .A(n1605), .B(n1604), .Z(n1606) );
  AND U1729 ( .A(n1607), .B(n1606), .Z(n1638) );
  NANDN U1730 ( .A(n5274), .B(n1608), .Z(n1610) );
  XOR U1731 ( .A(b[7]), .B(a[37]), .Z(n1649) );
  NANDN U1732 ( .A(n5275), .B(n1649), .Z(n1609) );
  AND U1733 ( .A(n1610), .B(n1609), .Z(n1668) );
  NANDN U1734 ( .A(n5176), .B(n1611), .Z(n1613) );
  XOR U1735 ( .A(b[3]), .B(a[41]), .Z(n1652) );
  NANDN U1736 ( .A(n5177), .B(n1652), .Z(n1612) );
  NAND U1737 ( .A(n1613), .B(n1612), .Z(n1667) );
  XNOR U1738 ( .A(n1668), .B(n1667), .Z(n1670) );
  NAND U1739 ( .A(b[0]), .B(a[43]), .Z(n1614) );
  XNOR U1740 ( .A(b[1]), .B(n1614), .Z(n1616) );
  NANDN U1741 ( .A(b[0]), .B(a[42]), .Z(n1615) );
  NAND U1742 ( .A(n1616), .B(n1615), .Z(n1664) );
  NANDN U1743 ( .A(n5249), .B(n1617), .Z(n1619) );
  XOR U1744 ( .A(b[5]), .B(a[39]), .Z(n1658) );
  NANDN U1745 ( .A(n5184), .B(n1658), .Z(n1618) );
  AND U1746 ( .A(n1619), .B(n1618), .Z(n1662) );
  AND U1747 ( .A(b[7]), .B(a[35]), .Z(n1661) );
  XNOR U1748 ( .A(n1662), .B(n1661), .Z(n1663) );
  XNOR U1749 ( .A(n1664), .B(n1663), .Z(n1669) );
  XOR U1750 ( .A(n1670), .B(n1669), .Z(n1644) );
  NANDN U1751 ( .A(n1621), .B(n1620), .Z(n1625) );
  NANDN U1752 ( .A(n1623), .B(n1622), .Z(n1624) );
  AND U1753 ( .A(n1625), .B(n1624), .Z(n1643) );
  XNOR U1754 ( .A(n1644), .B(n1643), .Z(n1645) );
  NANDN U1755 ( .A(n1627), .B(n1626), .Z(n1631) );
  NAND U1756 ( .A(n1629), .B(n1628), .Z(n1630) );
  NAND U1757 ( .A(n1631), .B(n1630), .Z(n1646) );
  XNOR U1758 ( .A(n1645), .B(n1646), .Z(n1637) );
  XNOR U1759 ( .A(n1638), .B(n1637), .Z(n1639) );
  XNOR U1760 ( .A(n1640), .B(n1639), .Z(n1673) );
  XNOR U1761 ( .A(sreg[163]), .B(n1673), .Z(n1675) );
  NANDN U1762 ( .A(sreg[162]), .B(n1632), .Z(n1636) );
  NAND U1763 ( .A(n1634), .B(n1633), .Z(n1635) );
  NAND U1764 ( .A(n1636), .B(n1635), .Z(n1674) );
  XNOR U1765 ( .A(n1675), .B(n1674), .Z(c[163]) );
  NANDN U1766 ( .A(n1638), .B(n1637), .Z(n1642) );
  NANDN U1767 ( .A(n1640), .B(n1639), .Z(n1641) );
  AND U1768 ( .A(n1642), .B(n1641), .Z(n1681) );
  NANDN U1769 ( .A(n1644), .B(n1643), .Z(n1648) );
  NANDN U1770 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U1771 ( .A(n1648), .B(n1647), .Z(n1679) );
  NANDN U1772 ( .A(n5274), .B(n1649), .Z(n1651) );
  XOR U1773 ( .A(b[7]), .B(a[38]), .Z(n1690) );
  NANDN U1774 ( .A(n5275), .B(n1690), .Z(n1650) );
  AND U1775 ( .A(n1651), .B(n1650), .Z(n1709) );
  NANDN U1776 ( .A(n5176), .B(n1652), .Z(n1654) );
  XOR U1777 ( .A(b[3]), .B(a[42]), .Z(n1693) );
  NANDN U1778 ( .A(n5177), .B(n1693), .Z(n1653) );
  NAND U1779 ( .A(n1654), .B(n1653), .Z(n1708) );
  XNOR U1780 ( .A(n1709), .B(n1708), .Z(n1711) );
  NAND U1781 ( .A(b[0]), .B(a[44]), .Z(n1655) );
  XNOR U1782 ( .A(b[1]), .B(n1655), .Z(n1657) );
  NANDN U1783 ( .A(b[0]), .B(a[43]), .Z(n1656) );
  NAND U1784 ( .A(n1657), .B(n1656), .Z(n1705) );
  NANDN U1785 ( .A(n5249), .B(n1658), .Z(n1660) );
  XOR U1786 ( .A(b[5]), .B(a[40]), .Z(n1696) );
  NANDN U1787 ( .A(n5184), .B(n1696), .Z(n1659) );
  AND U1788 ( .A(n1660), .B(n1659), .Z(n1703) );
  AND U1789 ( .A(b[7]), .B(a[36]), .Z(n1702) );
  XNOR U1790 ( .A(n1703), .B(n1702), .Z(n1704) );
  XNOR U1791 ( .A(n1705), .B(n1704), .Z(n1710) );
  XOR U1792 ( .A(n1711), .B(n1710), .Z(n1685) );
  NANDN U1793 ( .A(n1662), .B(n1661), .Z(n1666) );
  NANDN U1794 ( .A(n1664), .B(n1663), .Z(n1665) );
  AND U1795 ( .A(n1666), .B(n1665), .Z(n1684) );
  XNOR U1796 ( .A(n1685), .B(n1684), .Z(n1686) );
  NANDN U1797 ( .A(n1668), .B(n1667), .Z(n1672) );
  NAND U1798 ( .A(n1670), .B(n1669), .Z(n1671) );
  NAND U1799 ( .A(n1672), .B(n1671), .Z(n1687) );
  XNOR U1800 ( .A(n1686), .B(n1687), .Z(n1678) );
  XNOR U1801 ( .A(n1679), .B(n1678), .Z(n1680) );
  XNOR U1802 ( .A(n1681), .B(n1680), .Z(n1714) );
  XNOR U1803 ( .A(sreg[164]), .B(n1714), .Z(n1716) );
  NANDN U1804 ( .A(sreg[163]), .B(n1673), .Z(n1677) );
  NAND U1805 ( .A(n1675), .B(n1674), .Z(n1676) );
  NAND U1806 ( .A(n1677), .B(n1676), .Z(n1715) );
  XNOR U1807 ( .A(n1716), .B(n1715), .Z(c[164]) );
  NANDN U1808 ( .A(n1679), .B(n1678), .Z(n1683) );
  NANDN U1809 ( .A(n1681), .B(n1680), .Z(n1682) );
  AND U1810 ( .A(n1683), .B(n1682), .Z(n1722) );
  NANDN U1811 ( .A(n1685), .B(n1684), .Z(n1689) );
  NANDN U1812 ( .A(n1687), .B(n1686), .Z(n1688) );
  AND U1813 ( .A(n1689), .B(n1688), .Z(n1720) );
  NANDN U1814 ( .A(n5274), .B(n1690), .Z(n1692) );
  XOR U1815 ( .A(b[7]), .B(a[39]), .Z(n1731) );
  NANDN U1816 ( .A(n5275), .B(n1731), .Z(n1691) );
  AND U1817 ( .A(n1692), .B(n1691), .Z(n1750) );
  NANDN U1818 ( .A(n5176), .B(n1693), .Z(n1695) );
  XOR U1819 ( .A(b[3]), .B(a[43]), .Z(n1734) );
  NANDN U1820 ( .A(n5177), .B(n1734), .Z(n1694) );
  NAND U1821 ( .A(n1695), .B(n1694), .Z(n1749) );
  XNOR U1822 ( .A(n1750), .B(n1749), .Z(n1752) );
  NANDN U1823 ( .A(n5249), .B(n1696), .Z(n1698) );
  XOR U1824 ( .A(b[5]), .B(a[41]), .Z(n1740) );
  NANDN U1825 ( .A(n5184), .B(n1740), .Z(n1697) );
  AND U1826 ( .A(n1698), .B(n1697), .Z(n1744) );
  AND U1827 ( .A(b[7]), .B(a[37]), .Z(n1743) );
  XNOR U1828 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U1829 ( .A(b[0]), .B(a[45]), .Z(n1699) );
  XNOR U1830 ( .A(b[1]), .B(n1699), .Z(n1701) );
  NANDN U1831 ( .A(b[0]), .B(a[44]), .Z(n1700) );
  NAND U1832 ( .A(n1701), .B(n1700), .Z(n1746) );
  XNOR U1833 ( .A(n1745), .B(n1746), .Z(n1751) );
  XOR U1834 ( .A(n1752), .B(n1751), .Z(n1726) );
  NANDN U1835 ( .A(n1703), .B(n1702), .Z(n1707) );
  NANDN U1836 ( .A(n1705), .B(n1704), .Z(n1706) );
  AND U1837 ( .A(n1707), .B(n1706), .Z(n1725) );
  XNOR U1838 ( .A(n1726), .B(n1725), .Z(n1727) );
  NANDN U1839 ( .A(n1709), .B(n1708), .Z(n1713) );
  NAND U1840 ( .A(n1711), .B(n1710), .Z(n1712) );
  NAND U1841 ( .A(n1713), .B(n1712), .Z(n1728) );
  XNOR U1842 ( .A(n1727), .B(n1728), .Z(n1719) );
  XNOR U1843 ( .A(n1720), .B(n1719), .Z(n1721) );
  XNOR U1844 ( .A(n1722), .B(n1721), .Z(n1755) );
  XNOR U1845 ( .A(sreg[165]), .B(n1755), .Z(n1757) );
  NANDN U1846 ( .A(sreg[164]), .B(n1714), .Z(n1718) );
  NAND U1847 ( .A(n1716), .B(n1715), .Z(n1717) );
  NAND U1848 ( .A(n1718), .B(n1717), .Z(n1756) );
  XNOR U1849 ( .A(n1757), .B(n1756), .Z(c[165]) );
  NANDN U1850 ( .A(n1720), .B(n1719), .Z(n1724) );
  NANDN U1851 ( .A(n1722), .B(n1721), .Z(n1723) );
  AND U1852 ( .A(n1724), .B(n1723), .Z(n1763) );
  NANDN U1853 ( .A(n1726), .B(n1725), .Z(n1730) );
  NANDN U1854 ( .A(n1728), .B(n1727), .Z(n1729) );
  AND U1855 ( .A(n1730), .B(n1729), .Z(n1761) );
  NANDN U1856 ( .A(n5274), .B(n1731), .Z(n1733) );
  XOR U1857 ( .A(b[7]), .B(a[40]), .Z(n1772) );
  NANDN U1858 ( .A(n5275), .B(n1772), .Z(n1732) );
  AND U1859 ( .A(n1733), .B(n1732), .Z(n1791) );
  NANDN U1860 ( .A(n5176), .B(n1734), .Z(n1736) );
  XOR U1861 ( .A(b[3]), .B(a[44]), .Z(n1775) );
  NANDN U1862 ( .A(n5177), .B(n1775), .Z(n1735) );
  NAND U1863 ( .A(n1736), .B(n1735), .Z(n1790) );
  XNOR U1864 ( .A(n1791), .B(n1790), .Z(n1793) );
  NAND U1865 ( .A(b[0]), .B(a[46]), .Z(n1737) );
  XNOR U1866 ( .A(b[1]), .B(n1737), .Z(n1739) );
  NANDN U1867 ( .A(b[0]), .B(a[45]), .Z(n1738) );
  NAND U1868 ( .A(n1739), .B(n1738), .Z(n1787) );
  NANDN U1869 ( .A(n5249), .B(n1740), .Z(n1742) );
  XOR U1870 ( .A(b[5]), .B(a[42]), .Z(n1781) );
  NANDN U1871 ( .A(n5184), .B(n1781), .Z(n1741) );
  AND U1872 ( .A(n1742), .B(n1741), .Z(n1785) );
  AND U1873 ( .A(b[7]), .B(a[38]), .Z(n1784) );
  XNOR U1874 ( .A(n1785), .B(n1784), .Z(n1786) );
  XNOR U1875 ( .A(n1787), .B(n1786), .Z(n1792) );
  XOR U1876 ( .A(n1793), .B(n1792), .Z(n1767) );
  NANDN U1877 ( .A(n1744), .B(n1743), .Z(n1748) );
  NANDN U1878 ( .A(n1746), .B(n1745), .Z(n1747) );
  AND U1879 ( .A(n1748), .B(n1747), .Z(n1766) );
  XNOR U1880 ( .A(n1767), .B(n1766), .Z(n1768) );
  NANDN U1881 ( .A(n1750), .B(n1749), .Z(n1754) );
  NAND U1882 ( .A(n1752), .B(n1751), .Z(n1753) );
  NAND U1883 ( .A(n1754), .B(n1753), .Z(n1769) );
  XNOR U1884 ( .A(n1768), .B(n1769), .Z(n1760) );
  XNOR U1885 ( .A(n1761), .B(n1760), .Z(n1762) );
  XNOR U1886 ( .A(n1763), .B(n1762), .Z(n1796) );
  XNOR U1887 ( .A(sreg[166]), .B(n1796), .Z(n1798) );
  NANDN U1888 ( .A(sreg[165]), .B(n1755), .Z(n1759) );
  NAND U1889 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U1890 ( .A(n1759), .B(n1758), .Z(n1797) );
  XNOR U1891 ( .A(n1798), .B(n1797), .Z(c[166]) );
  NANDN U1892 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U1893 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U1894 ( .A(n1765), .B(n1764), .Z(n1804) );
  NANDN U1895 ( .A(n1767), .B(n1766), .Z(n1771) );
  NANDN U1896 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U1897 ( .A(n1771), .B(n1770), .Z(n1802) );
  NANDN U1898 ( .A(n5274), .B(n1772), .Z(n1774) );
  XOR U1899 ( .A(b[7]), .B(a[41]), .Z(n1813) );
  NANDN U1900 ( .A(n5275), .B(n1813), .Z(n1773) );
  AND U1901 ( .A(n1774), .B(n1773), .Z(n1832) );
  NANDN U1902 ( .A(n5176), .B(n1775), .Z(n1777) );
  XOR U1903 ( .A(b[3]), .B(a[45]), .Z(n1816) );
  NANDN U1904 ( .A(n5177), .B(n1816), .Z(n1776) );
  NAND U1905 ( .A(n1777), .B(n1776), .Z(n1831) );
  XNOR U1906 ( .A(n1832), .B(n1831), .Z(n1834) );
  NAND U1907 ( .A(b[0]), .B(a[47]), .Z(n1778) );
  XNOR U1908 ( .A(b[1]), .B(n1778), .Z(n1780) );
  NANDN U1909 ( .A(b[0]), .B(a[46]), .Z(n1779) );
  NAND U1910 ( .A(n1780), .B(n1779), .Z(n1828) );
  NANDN U1911 ( .A(n5249), .B(n1781), .Z(n1783) );
  XOR U1912 ( .A(b[5]), .B(a[43]), .Z(n1822) );
  NANDN U1913 ( .A(n5184), .B(n1822), .Z(n1782) );
  AND U1914 ( .A(n1783), .B(n1782), .Z(n1826) );
  AND U1915 ( .A(b[7]), .B(a[39]), .Z(n1825) );
  XNOR U1916 ( .A(n1826), .B(n1825), .Z(n1827) );
  XNOR U1917 ( .A(n1828), .B(n1827), .Z(n1833) );
  XOR U1918 ( .A(n1834), .B(n1833), .Z(n1808) );
  NANDN U1919 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U1920 ( .A(n1787), .B(n1786), .Z(n1788) );
  AND U1921 ( .A(n1789), .B(n1788), .Z(n1807) );
  XNOR U1922 ( .A(n1808), .B(n1807), .Z(n1809) );
  NANDN U1923 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U1924 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U1925 ( .A(n1795), .B(n1794), .Z(n1810) );
  XNOR U1926 ( .A(n1809), .B(n1810), .Z(n1801) );
  XNOR U1927 ( .A(n1802), .B(n1801), .Z(n1803) );
  XNOR U1928 ( .A(n1804), .B(n1803), .Z(n1837) );
  XNOR U1929 ( .A(sreg[167]), .B(n1837), .Z(n1839) );
  NANDN U1930 ( .A(sreg[166]), .B(n1796), .Z(n1800) );
  NAND U1931 ( .A(n1798), .B(n1797), .Z(n1799) );
  NAND U1932 ( .A(n1800), .B(n1799), .Z(n1838) );
  XNOR U1933 ( .A(n1839), .B(n1838), .Z(c[167]) );
  NANDN U1934 ( .A(n1802), .B(n1801), .Z(n1806) );
  NANDN U1935 ( .A(n1804), .B(n1803), .Z(n1805) );
  AND U1936 ( .A(n1806), .B(n1805), .Z(n1845) );
  NANDN U1937 ( .A(n1808), .B(n1807), .Z(n1812) );
  NANDN U1938 ( .A(n1810), .B(n1809), .Z(n1811) );
  AND U1939 ( .A(n1812), .B(n1811), .Z(n1843) );
  NANDN U1940 ( .A(n5274), .B(n1813), .Z(n1815) );
  XOR U1941 ( .A(b[7]), .B(a[42]), .Z(n1854) );
  NANDN U1942 ( .A(n5275), .B(n1854), .Z(n1814) );
  AND U1943 ( .A(n1815), .B(n1814), .Z(n1873) );
  NANDN U1944 ( .A(n5176), .B(n1816), .Z(n1818) );
  XOR U1945 ( .A(b[3]), .B(a[46]), .Z(n1857) );
  NANDN U1946 ( .A(n5177), .B(n1857), .Z(n1817) );
  NAND U1947 ( .A(n1818), .B(n1817), .Z(n1872) );
  XNOR U1948 ( .A(n1873), .B(n1872), .Z(n1875) );
  NAND U1949 ( .A(b[0]), .B(a[48]), .Z(n1819) );
  XNOR U1950 ( .A(b[1]), .B(n1819), .Z(n1821) );
  NANDN U1951 ( .A(b[0]), .B(a[47]), .Z(n1820) );
  NAND U1952 ( .A(n1821), .B(n1820), .Z(n1869) );
  NANDN U1953 ( .A(n5249), .B(n1822), .Z(n1824) );
  XOR U1954 ( .A(b[5]), .B(a[44]), .Z(n1860) );
  NANDN U1955 ( .A(n5184), .B(n1860), .Z(n1823) );
  AND U1956 ( .A(n1824), .B(n1823), .Z(n1867) );
  AND U1957 ( .A(b[7]), .B(a[40]), .Z(n1866) );
  XNOR U1958 ( .A(n1867), .B(n1866), .Z(n1868) );
  XNOR U1959 ( .A(n1869), .B(n1868), .Z(n1874) );
  XOR U1960 ( .A(n1875), .B(n1874), .Z(n1849) );
  NANDN U1961 ( .A(n1826), .B(n1825), .Z(n1830) );
  NANDN U1962 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U1963 ( .A(n1830), .B(n1829), .Z(n1848) );
  XNOR U1964 ( .A(n1849), .B(n1848), .Z(n1850) );
  NANDN U1965 ( .A(n1832), .B(n1831), .Z(n1836) );
  NAND U1966 ( .A(n1834), .B(n1833), .Z(n1835) );
  NAND U1967 ( .A(n1836), .B(n1835), .Z(n1851) );
  XNOR U1968 ( .A(n1850), .B(n1851), .Z(n1842) );
  XNOR U1969 ( .A(n1843), .B(n1842), .Z(n1844) );
  XNOR U1970 ( .A(n1845), .B(n1844), .Z(n1878) );
  XNOR U1971 ( .A(sreg[168]), .B(n1878), .Z(n1880) );
  NANDN U1972 ( .A(sreg[167]), .B(n1837), .Z(n1841) );
  NAND U1973 ( .A(n1839), .B(n1838), .Z(n1840) );
  NAND U1974 ( .A(n1841), .B(n1840), .Z(n1879) );
  XNOR U1975 ( .A(n1880), .B(n1879), .Z(c[168]) );
  NANDN U1976 ( .A(n1843), .B(n1842), .Z(n1847) );
  NANDN U1977 ( .A(n1845), .B(n1844), .Z(n1846) );
  AND U1978 ( .A(n1847), .B(n1846), .Z(n1886) );
  NANDN U1979 ( .A(n1849), .B(n1848), .Z(n1853) );
  NANDN U1980 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U1981 ( .A(n1853), .B(n1852), .Z(n1884) );
  NANDN U1982 ( .A(n5274), .B(n1854), .Z(n1856) );
  XOR U1983 ( .A(b[7]), .B(a[43]), .Z(n1895) );
  NANDN U1984 ( .A(n5275), .B(n1895), .Z(n1855) );
  AND U1985 ( .A(n1856), .B(n1855), .Z(n1914) );
  NANDN U1986 ( .A(n5176), .B(n1857), .Z(n1859) );
  XOR U1987 ( .A(b[3]), .B(a[47]), .Z(n1898) );
  NANDN U1988 ( .A(n5177), .B(n1898), .Z(n1858) );
  NAND U1989 ( .A(n1859), .B(n1858), .Z(n1913) );
  XNOR U1990 ( .A(n1914), .B(n1913), .Z(n1916) );
  NANDN U1991 ( .A(n5249), .B(n1860), .Z(n1862) );
  XOR U1992 ( .A(b[5]), .B(a[45]), .Z(n1904) );
  NANDN U1993 ( .A(n5184), .B(n1904), .Z(n1861) );
  AND U1994 ( .A(n1862), .B(n1861), .Z(n1908) );
  AND U1995 ( .A(b[7]), .B(a[41]), .Z(n1907) );
  XNOR U1996 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U1997 ( .A(b[0]), .B(a[49]), .Z(n1863) );
  XNOR U1998 ( .A(b[1]), .B(n1863), .Z(n1865) );
  NANDN U1999 ( .A(b[0]), .B(a[48]), .Z(n1864) );
  NAND U2000 ( .A(n1865), .B(n1864), .Z(n1910) );
  XNOR U2001 ( .A(n1909), .B(n1910), .Z(n1915) );
  XOR U2002 ( .A(n1916), .B(n1915), .Z(n1890) );
  NANDN U2003 ( .A(n1867), .B(n1866), .Z(n1871) );
  NANDN U2004 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2005 ( .A(n1871), .B(n1870), .Z(n1889) );
  XNOR U2006 ( .A(n1890), .B(n1889), .Z(n1891) );
  NANDN U2007 ( .A(n1873), .B(n1872), .Z(n1877) );
  NAND U2008 ( .A(n1875), .B(n1874), .Z(n1876) );
  NAND U2009 ( .A(n1877), .B(n1876), .Z(n1892) );
  XNOR U2010 ( .A(n1891), .B(n1892), .Z(n1883) );
  XNOR U2011 ( .A(n1884), .B(n1883), .Z(n1885) );
  XNOR U2012 ( .A(n1886), .B(n1885), .Z(n1919) );
  XNOR U2013 ( .A(sreg[169]), .B(n1919), .Z(n1921) );
  NANDN U2014 ( .A(sreg[168]), .B(n1878), .Z(n1882) );
  NAND U2015 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2016 ( .A(n1882), .B(n1881), .Z(n1920) );
  XNOR U2017 ( .A(n1921), .B(n1920), .Z(c[169]) );
  NANDN U2018 ( .A(n1884), .B(n1883), .Z(n1888) );
  NANDN U2019 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2020 ( .A(n1888), .B(n1887), .Z(n1927) );
  NANDN U2021 ( .A(n1890), .B(n1889), .Z(n1894) );
  NANDN U2022 ( .A(n1892), .B(n1891), .Z(n1893) );
  AND U2023 ( .A(n1894), .B(n1893), .Z(n1925) );
  NANDN U2024 ( .A(n5274), .B(n1895), .Z(n1897) );
  XOR U2025 ( .A(b[7]), .B(a[44]), .Z(n1936) );
  NANDN U2026 ( .A(n5275), .B(n1936), .Z(n1896) );
  AND U2027 ( .A(n1897), .B(n1896), .Z(n1955) );
  NANDN U2028 ( .A(n5176), .B(n1898), .Z(n1900) );
  XOR U2029 ( .A(b[3]), .B(a[48]), .Z(n1939) );
  NANDN U2030 ( .A(n5177), .B(n1939), .Z(n1899) );
  NAND U2031 ( .A(n1900), .B(n1899), .Z(n1954) );
  XNOR U2032 ( .A(n1955), .B(n1954), .Z(n1957) );
  NAND U2033 ( .A(b[0]), .B(a[50]), .Z(n1901) );
  XNOR U2034 ( .A(b[1]), .B(n1901), .Z(n1903) );
  NANDN U2035 ( .A(b[0]), .B(a[49]), .Z(n1902) );
  NAND U2036 ( .A(n1903), .B(n1902), .Z(n1951) );
  NANDN U2037 ( .A(n5249), .B(n1904), .Z(n1906) );
  XOR U2038 ( .A(b[5]), .B(a[46]), .Z(n1945) );
  NANDN U2039 ( .A(n5184), .B(n1945), .Z(n1905) );
  AND U2040 ( .A(n1906), .B(n1905), .Z(n1949) );
  AND U2041 ( .A(b[7]), .B(a[42]), .Z(n1948) );
  XNOR U2042 ( .A(n1949), .B(n1948), .Z(n1950) );
  XNOR U2043 ( .A(n1951), .B(n1950), .Z(n1956) );
  XOR U2044 ( .A(n1957), .B(n1956), .Z(n1931) );
  NANDN U2045 ( .A(n1908), .B(n1907), .Z(n1912) );
  NANDN U2046 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2047 ( .A(n1912), .B(n1911), .Z(n1930) );
  XNOR U2048 ( .A(n1931), .B(n1930), .Z(n1932) );
  NANDN U2049 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2050 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2051 ( .A(n1918), .B(n1917), .Z(n1933) );
  XNOR U2052 ( .A(n1932), .B(n1933), .Z(n1924) );
  XNOR U2053 ( .A(n1925), .B(n1924), .Z(n1926) );
  XNOR U2054 ( .A(n1927), .B(n1926), .Z(n1960) );
  XNOR U2055 ( .A(sreg[170]), .B(n1960), .Z(n1962) );
  NANDN U2056 ( .A(sreg[169]), .B(n1919), .Z(n1923) );
  NAND U2057 ( .A(n1921), .B(n1920), .Z(n1922) );
  NAND U2058 ( .A(n1923), .B(n1922), .Z(n1961) );
  XNOR U2059 ( .A(n1962), .B(n1961), .Z(c[170]) );
  NANDN U2060 ( .A(n1925), .B(n1924), .Z(n1929) );
  NANDN U2061 ( .A(n1927), .B(n1926), .Z(n1928) );
  AND U2062 ( .A(n1929), .B(n1928), .Z(n1968) );
  NANDN U2063 ( .A(n1931), .B(n1930), .Z(n1935) );
  NANDN U2064 ( .A(n1933), .B(n1932), .Z(n1934) );
  AND U2065 ( .A(n1935), .B(n1934), .Z(n1966) );
  NANDN U2066 ( .A(n5274), .B(n1936), .Z(n1938) );
  XOR U2067 ( .A(b[7]), .B(a[45]), .Z(n1977) );
  NANDN U2068 ( .A(n5275), .B(n1977), .Z(n1937) );
  AND U2069 ( .A(n1938), .B(n1937), .Z(n1996) );
  NANDN U2070 ( .A(n5176), .B(n1939), .Z(n1941) );
  XOR U2071 ( .A(b[3]), .B(a[49]), .Z(n1980) );
  NANDN U2072 ( .A(n5177), .B(n1980), .Z(n1940) );
  NAND U2073 ( .A(n1941), .B(n1940), .Z(n1995) );
  XNOR U2074 ( .A(n1996), .B(n1995), .Z(n1998) );
  NAND U2075 ( .A(b[0]), .B(a[51]), .Z(n1942) );
  XNOR U2076 ( .A(b[1]), .B(n1942), .Z(n1944) );
  NANDN U2077 ( .A(b[0]), .B(a[50]), .Z(n1943) );
  NAND U2078 ( .A(n1944), .B(n1943), .Z(n1992) );
  NANDN U2079 ( .A(n5249), .B(n1945), .Z(n1947) );
  XOR U2080 ( .A(b[5]), .B(a[47]), .Z(n1986) );
  NANDN U2081 ( .A(n5184), .B(n1986), .Z(n1946) );
  AND U2082 ( .A(n1947), .B(n1946), .Z(n1990) );
  AND U2083 ( .A(b[7]), .B(a[43]), .Z(n1989) );
  XNOR U2084 ( .A(n1990), .B(n1989), .Z(n1991) );
  XNOR U2085 ( .A(n1992), .B(n1991), .Z(n1997) );
  XOR U2086 ( .A(n1998), .B(n1997), .Z(n1972) );
  NANDN U2087 ( .A(n1949), .B(n1948), .Z(n1953) );
  NANDN U2088 ( .A(n1951), .B(n1950), .Z(n1952) );
  AND U2089 ( .A(n1953), .B(n1952), .Z(n1971) );
  XNOR U2090 ( .A(n1972), .B(n1971), .Z(n1973) );
  NANDN U2091 ( .A(n1955), .B(n1954), .Z(n1959) );
  NAND U2092 ( .A(n1957), .B(n1956), .Z(n1958) );
  NAND U2093 ( .A(n1959), .B(n1958), .Z(n1974) );
  XNOR U2094 ( .A(n1973), .B(n1974), .Z(n1965) );
  XNOR U2095 ( .A(n1966), .B(n1965), .Z(n1967) );
  XNOR U2096 ( .A(n1968), .B(n1967), .Z(n2001) );
  XNOR U2097 ( .A(sreg[171]), .B(n2001), .Z(n2003) );
  NANDN U2098 ( .A(sreg[170]), .B(n1960), .Z(n1964) );
  NAND U2099 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2100 ( .A(n1964), .B(n1963), .Z(n2002) );
  XNOR U2101 ( .A(n2003), .B(n2002), .Z(c[171]) );
  NANDN U2102 ( .A(n1966), .B(n1965), .Z(n1970) );
  NANDN U2103 ( .A(n1968), .B(n1967), .Z(n1969) );
  AND U2104 ( .A(n1970), .B(n1969), .Z(n2009) );
  NANDN U2105 ( .A(n1972), .B(n1971), .Z(n1976) );
  NANDN U2106 ( .A(n1974), .B(n1973), .Z(n1975) );
  AND U2107 ( .A(n1976), .B(n1975), .Z(n2007) );
  NANDN U2108 ( .A(n5274), .B(n1977), .Z(n1979) );
  XOR U2109 ( .A(b[7]), .B(a[46]), .Z(n2018) );
  NANDN U2110 ( .A(n5275), .B(n2018), .Z(n1978) );
  AND U2111 ( .A(n1979), .B(n1978), .Z(n2037) );
  NANDN U2112 ( .A(n5176), .B(n1980), .Z(n1982) );
  XOR U2113 ( .A(b[3]), .B(a[50]), .Z(n2021) );
  NANDN U2114 ( .A(n5177), .B(n2021), .Z(n1981) );
  NAND U2115 ( .A(n1982), .B(n1981), .Z(n2036) );
  XNOR U2116 ( .A(n2037), .B(n2036), .Z(n2039) );
  NAND U2117 ( .A(b[0]), .B(a[52]), .Z(n1983) );
  XNOR U2118 ( .A(b[1]), .B(n1983), .Z(n1985) );
  NANDN U2119 ( .A(b[0]), .B(a[51]), .Z(n1984) );
  NAND U2120 ( .A(n1985), .B(n1984), .Z(n2033) );
  NANDN U2121 ( .A(n5249), .B(n1986), .Z(n1988) );
  XOR U2122 ( .A(b[5]), .B(a[48]), .Z(n2024) );
  NANDN U2123 ( .A(n5184), .B(n2024), .Z(n1987) );
  AND U2124 ( .A(n1988), .B(n1987), .Z(n2031) );
  AND U2125 ( .A(b[7]), .B(a[44]), .Z(n2030) );
  XNOR U2126 ( .A(n2031), .B(n2030), .Z(n2032) );
  XNOR U2127 ( .A(n2033), .B(n2032), .Z(n2038) );
  XOR U2128 ( .A(n2039), .B(n2038), .Z(n2013) );
  NANDN U2129 ( .A(n1990), .B(n1989), .Z(n1994) );
  NANDN U2130 ( .A(n1992), .B(n1991), .Z(n1993) );
  AND U2131 ( .A(n1994), .B(n1993), .Z(n2012) );
  XNOR U2132 ( .A(n2013), .B(n2012), .Z(n2014) );
  NANDN U2133 ( .A(n1996), .B(n1995), .Z(n2000) );
  NAND U2134 ( .A(n1998), .B(n1997), .Z(n1999) );
  NAND U2135 ( .A(n2000), .B(n1999), .Z(n2015) );
  XNOR U2136 ( .A(n2014), .B(n2015), .Z(n2006) );
  XNOR U2137 ( .A(n2007), .B(n2006), .Z(n2008) );
  XNOR U2138 ( .A(n2009), .B(n2008), .Z(n2042) );
  XNOR U2139 ( .A(sreg[172]), .B(n2042), .Z(n2044) );
  NANDN U2140 ( .A(sreg[171]), .B(n2001), .Z(n2005) );
  NAND U2141 ( .A(n2003), .B(n2002), .Z(n2004) );
  NAND U2142 ( .A(n2005), .B(n2004), .Z(n2043) );
  XNOR U2143 ( .A(n2044), .B(n2043), .Z(c[172]) );
  NANDN U2144 ( .A(n2007), .B(n2006), .Z(n2011) );
  NANDN U2145 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U2146 ( .A(n2011), .B(n2010), .Z(n2050) );
  NANDN U2147 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2148 ( .A(n2015), .B(n2014), .Z(n2016) );
  AND U2149 ( .A(n2017), .B(n2016), .Z(n2048) );
  NANDN U2150 ( .A(n5274), .B(n2018), .Z(n2020) );
  XOR U2151 ( .A(b[7]), .B(a[47]), .Z(n2059) );
  NANDN U2152 ( .A(n5275), .B(n2059), .Z(n2019) );
  AND U2153 ( .A(n2020), .B(n2019), .Z(n2078) );
  NANDN U2154 ( .A(n5176), .B(n2021), .Z(n2023) );
  XOR U2155 ( .A(b[3]), .B(a[51]), .Z(n2062) );
  NANDN U2156 ( .A(n5177), .B(n2062), .Z(n2022) );
  NAND U2157 ( .A(n2023), .B(n2022), .Z(n2077) );
  XNOR U2158 ( .A(n2078), .B(n2077), .Z(n2080) );
  NANDN U2159 ( .A(n5249), .B(n2024), .Z(n2026) );
  XOR U2160 ( .A(b[5]), .B(a[49]), .Z(n2068) );
  NANDN U2161 ( .A(n5184), .B(n2068), .Z(n2025) );
  AND U2162 ( .A(n2026), .B(n2025), .Z(n2072) );
  AND U2163 ( .A(b[7]), .B(a[45]), .Z(n2071) );
  XNOR U2164 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U2165 ( .A(b[0]), .B(a[53]), .Z(n2027) );
  XNOR U2166 ( .A(b[1]), .B(n2027), .Z(n2029) );
  NANDN U2167 ( .A(b[0]), .B(a[52]), .Z(n2028) );
  NAND U2168 ( .A(n2029), .B(n2028), .Z(n2074) );
  XNOR U2169 ( .A(n2073), .B(n2074), .Z(n2079) );
  XOR U2170 ( .A(n2080), .B(n2079), .Z(n2054) );
  NANDN U2171 ( .A(n2031), .B(n2030), .Z(n2035) );
  NANDN U2172 ( .A(n2033), .B(n2032), .Z(n2034) );
  AND U2173 ( .A(n2035), .B(n2034), .Z(n2053) );
  XNOR U2174 ( .A(n2054), .B(n2053), .Z(n2055) );
  NANDN U2175 ( .A(n2037), .B(n2036), .Z(n2041) );
  NAND U2176 ( .A(n2039), .B(n2038), .Z(n2040) );
  NAND U2177 ( .A(n2041), .B(n2040), .Z(n2056) );
  XNOR U2178 ( .A(n2055), .B(n2056), .Z(n2047) );
  XNOR U2179 ( .A(n2048), .B(n2047), .Z(n2049) );
  XNOR U2180 ( .A(n2050), .B(n2049), .Z(n2083) );
  XNOR U2181 ( .A(sreg[173]), .B(n2083), .Z(n2085) );
  NANDN U2182 ( .A(sreg[172]), .B(n2042), .Z(n2046) );
  NAND U2183 ( .A(n2044), .B(n2043), .Z(n2045) );
  NAND U2184 ( .A(n2046), .B(n2045), .Z(n2084) );
  XNOR U2185 ( .A(n2085), .B(n2084), .Z(c[173]) );
  NANDN U2186 ( .A(n2048), .B(n2047), .Z(n2052) );
  NANDN U2187 ( .A(n2050), .B(n2049), .Z(n2051) );
  AND U2188 ( .A(n2052), .B(n2051), .Z(n2091) );
  NANDN U2189 ( .A(n2054), .B(n2053), .Z(n2058) );
  NANDN U2190 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U2191 ( .A(n2058), .B(n2057), .Z(n2089) );
  NANDN U2192 ( .A(n5274), .B(n2059), .Z(n2061) );
  XOR U2193 ( .A(b[7]), .B(a[48]), .Z(n2100) );
  NANDN U2194 ( .A(n5275), .B(n2100), .Z(n2060) );
  AND U2195 ( .A(n2061), .B(n2060), .Z(n2119) );
  NANDN U2196 ( .A(n5176), .B(n2062), .Z(n2064) );
  XOR U2197 ( .A(b[3]), .B(a[52]), .Z(n2103) );
  NANDN U2198 ( .A(n5177), .B(n2103), .Z(n2063) );
  NAND U2199 ( .A(n2064), .B(n2063), .Z(n2118) );
  XNOR U2200 ( .A(n2119), .B(n2118), .Z(n2121) );
  NAND U2201 ( .A(b[0]), .B(a[54]), .Z(n2065) );
  XNOR U2202 ( .A(b[1]), .B(n2065), .Z(n2067) );
  NANDN U2203 ( .A(b[0]), .B(a[53]), .Z(n2066) );
  NAND U2204 ( .A(n2067), .B(n2066), .Z(n2115) );
  NANDN U2205 ( .A(n5249), .B(n2068), .Z(n2070) );
  XOR U2206 ( .A(b[5]), .B(a[50]), .Z(n2106) );
  NANDN U2207 ( .A(n5184), .B(n2106), .Z(n2069) );
  AND U2208 ( .A(n2070), .B(n2069), .Z(n2113) );
  AND U2209 ( .A(b[7]), .B(a[46]), .Z(n2112) );
  XNOR U2210 ( .A(n2113), .B(n2112), .Z(n2114) );
  XNOR U2211 ( .A(n2115), .B(n2114), .Z(n2120) );
  XOR U2212 ( .A(n2121), .B(n2120), .Z(n2095) );
  NANDN U2213 ( .A(n2072), .B(n2071), .Z(n2076) );
  NANDN U2214 ( .A(n2074), .B(n2073), .Z(n2075) );
  AND U2215 ( .A(n2076), .B(n2075), .Z(n2094) );
  XNOR U2216 ( .A(n2095), .B(n2094), .Z(n2096) );
  NANDN U2217 ( .A(n2078), .B(n2077), .Z(n2082) );
  NAND U2218 ( .A(n2080), .B(n2079), .Z(n2081) );
  NAND U2219 ( .A(n2082), .B(n2081), .Z(n2097) );
  XNOR U2220 ( .A(n2096), .B(n2097), .Z(n2088) );
  XNOR U2221 ( .A(n2089), .B(n2088), .Z(n2090) );
  XNOR U2222 ( .A(n2091), .B(n2090), .Z(n2124) );
  XNOR U2223 ( .A(sreg[174]), .B(n2124), .Z(n2126) );
  NANDN U2224 ( .A(sreg[173]), .B(n2083), .Z(n2087) );
  NAND U2225 ( .A(n2085), .B(n2084), .Z(n2086) );
  NAND U2226 ( .A(n2087), .B(n2086), .Z(n2125) );
  XNOR U2227 ( .A(n2126), .B(n2125), .Z(c[174]) );
  NANDN U2228 ( .A(n2089), .B(n2088), .Z(n2093) );
  NANDN U2229 ( .A(n2091), .B(n2090), .Z(n2092) );
  AND U2230 ( .A(n2093), .B(n2092), .Z(n2132) );
  NANDN U2231 ( .A(n2095), .B(n2094), .Z(n2099) );
  NANDN U2232 ( .A(n2097), .B(n2096), .Z(n2098) );
  AND U2233 ( .A(n2099), .B(n2098), .Z(n2130) );
  NANDN U2234 ( .A(n5274), .B(n2100), .Z(n2102) );
  XOR U2235 ( .A(b[7]), .B(a[49]), .Z(n2141) );
  NANDN U2236 ( .A(n5275), .B(n2141), .Z(n2101) );
  AND U2237 ( .A(n2102), .B(n2101), .Z(n2160) );
  NANDN U2238 ( .A(n5176), .B(n2103), .Z(n2105) );
  XOR U2239 ( .A(b[3]), .B(a[53]), .Z(n2144) );
  NANDN U2240 ( .A(n5177), .B(n2144), .Z(n2104) );
  NAND U2241 ( .A(n2105), .B(n2104), .Z(n2159) );
  XNOR U2242 ( .A(n2160), .B(n2159), .Z(n2162) );
  NANDN U2243 ( .A(n5249), .B(n2106), .Z(n2108) );
  XOR U2244 ( .A(b[5]), .B(a[51]), .Z(n2150) );
  NANDN U2245 ( .A(n5184), .B(n2150), .Z(n2107) );
  AND U2246 ( .A(n2108), .B(n2107), .Z(n2154) );
  AND U2247 ( .A(b[7]), .B(a[47]), .Z(n2153) );
  XNOR U2248 ( .A(n2154), .B(n2153), .Z(n2155) );
  NAND U2249 ( .A(b[0]), .B(a[55]), .Z(n2109) );
  XNOR U2250 ( .A(b[1]), .B(n2109), .Z(n2111) );
  NANDN U2251 ( .A(b[0]), .B(a[54]), .Z(n2110) );
  NAND U2252 ( .A(n2111), .B(n2110), .Z(n2156) );
  XNOR U2253 ( .A(n2155), .B(n2156), .Z(n2161) );
  XOR U2254 ( .A(n2162), .B(n2161), .Z(n2136) );
  NANDN U2255 ( .A(n2113), .B(n2112), .Z(n2117) );
  NANDN U2256 ( .A(n2115), .B(n2114), .Z(n2116) );
  AND U2257 ( .A(n2117), .B(n2116), .Z(n2135) );
  XNOR U2258 ( .A(n2136), .B(n2135), .Z(n2137) );
  NANDN U2259 ( .A(n2119), .B(n2118), .Z(n2123) );
  NAND U2260 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U2261 ( .A(n2123), .B(n2122), .Z(n2138) );
  XNOR U2262 ( .A(n2137), .B(n2138), .Z(n2129) );
  XNOR U2263 ( .A(n2130), .B(n2129), .Z(n2131) );
  XNOR U2264 ( .A(n2132), .B(n2131), .Z(n2165) );
  XNOR U2265 ( .A(sreg[175]), .B(n2165), .Z(n2167) );
  NANDN U2266 ( .A(sreg[174]), .B(n2124), .Z(n2128) );
  NAND U2267 ( .A(n2126), .B(n2125), .Z(n2127) );
  NAND U2268 ( .A(n2128), .B(n2127), .Z(n2166) );
  XNOR U2269 ( .A(n2167), .B(n2166), .Z(c[175]) );
  NANDN U2270 ( .A(n2130), .B(n2129), .Z(n2134) );
  NANDN U2271 ( .A(n2132), .B(n2131), .Z(n2133) );
  AND U2272 ( .A(n2134), .B(n2133), .Z(n2173) );
  NANDN U2273 ( .A(n2136), .B(n2135), .Z(n2140) );
  NANDN U2274 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U2275 ( .A(n2140), .B(n2139), .Z(n2171) );
  NANDN U2276 ( .A(n5274), .B(n2141), .Z(n2143) );
  XOR U2277 ( .A(b[7]), .B(a[50]), .Z(n2182) );
  NANDN U2278 ( .A(n5275), .B(n2182), .Z(n2142) );
  AND U2279 ( .A(n2143), .B(n2142), .Z(n2201) );
  NANDN U2280 ( .A(n5176), .B(n2144), .Z(n2146) );
  XOR U2281 ( .A(b[3]), .B(a[54]), .Z(n2185) );
  NANDN U2282 ( .A(n5177), .B(n2185), .Z(n2145) );
  NAND U2283 ( .A(n2146), .B(n2145), .Z(n2200) );
  XNOR U2284 ( .A(n2201), .B(n2200), .Z(n2203) );
  NAND U2285 ( .A(b[0]), .B(a[56]), .Z(n2147) );
  XNOR U2286 ( .A(b[1]), .B(n2147), .Z(n2149) );
  NANDN U2287 ( .A(b[0]), .B(a[55]), .Z(n2148) );
  NAND U2288 ( .A(n2149), .B(n2148), .Z(n2197) );
  NANDN U2289 ( .A(n5249), .B(n2150), .Z(n2152) );
  XOR U2290 ( .A(b[5]), .B(a[52]), .Z(n2188) );
  NANDN U2291 ( .A(n5184), .B(n2188), .Z(n2151) );
  AND U2292 ( .A(n2152), .B(n2151), .Z(n2195) );
  AND U2293 ( .A(b[7]), .B(a[48]), .Z(n2194) );
  XNOR U2294 ( .A(n2195), .B(n2194), .Z(n2196) );
  XNOR U2295 ( .A(n2197), .B(n2196), .Z(n2202) );
  XOR U2296 ( .A(n2203), .B(n2202), .Z(n2177) );
  NANDN U2297 ( .A(n2154), .B(n2153), .Z(n2158) );
  NANDN U2298 ( .A(n2156), .B(n2155), .Z(n2157) );
  AND U2299 ( .A(n2158), .B(n2157), .Z(n2176) );
  XNOR U2300 ( .A(n2177), .B(n2176), .Z(n2178) );
  NANDN U2301 ( .A(n2160), .B(n2159), .Z(n2164) );
  NAND U2302 ( .A(n2162), .B(n2161), .Z(n2163) );
  NAND U2303 ( .A(n2164), .B(n2163), .Z(n2179) );
  XNOR U2304 ( .A(n2178), .B(n2179), .Z(n2170) );
  XNOR U2305 ( .A(n2171), .B(n2170), .Z(n2172) );
  XNOR U2306 ( .A(n2173), .B(n2172), .Z(n2206) );
  XNOR U2307 ( .A(sreg[176]), .B(n2206), .Z(n2208) );
  NANDN U2308 ( .A(sreg[175]), .B(n2165), .Z(n2169) );
  NAND U2309 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2310 ( .A(n2169), .B(n2168), .Z(n2207) );
  XNOR U2311 ( .A(n2208), .B(n2207), .Z(c[176]) );
  NANDN U2312 ( .A(n2171), .B(n2170), .Z(n2175) );
  NANDN U2313 ( .A(n2173), .B(n2172), .Z(n2174) );
  AND U2314 ( .A(n2175), .B(n2174), .Z(n2214) );
  NANDN U2315 ( .A(n2177), .B(n2176), .Z(n2181) );
  NANDN U2316 ( .A(n2179), .B(n2178), .Z(n2180) );
  AND U2317 ( .A(n2181), .B(n2180), .Z(n2212) );
  NANDN U2318 ( .A(n5274), .B(n2182), .Z(n2184) );
  XOR U2319 ( .A(b[7]), .B(a[51]), .Z(n2223) );
  NANDN U2320 ( .A(n5275), .B(n2223), .Z(n2183) );
  AND U2321 ( .A(n2184), .B(n2183), .Z(n2242) );
  NANDN U2322 ( .A(n5176), .B(n2185), .Z(n2187) );
  XOR U2323 ( .A(b[3]), .B(a[55]), .Z(n2226) );
  NANDN U2324 ( .A(n5177), .B(n2226), .Z(n2186) );
  NAND U2325 ( .A(n2187), .B(n2186), .Z(n2241) );
  XNOR U2326 ( .A(n2242), .B(n2241), .Z(n2244) );
  NANDN U2327 ( .A(n5249), .B(n2188), .Z(n2190) );
  XOR U2328 ( .A(b[5]), .B(a[53]), .Z(n2232) );
  NANDN U2329 ( .A(n5184), .B(n2232), .Z(n2189) );
  AND U2330 ( .A(n2190), .B(n2189), .Z(n2236) );
  AND U2331 ( .A(b[7]), .B(a[49]), .Z(n2235) );
  XNOR U2332 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2333 ( .A(b[0]), .B(a[57]), .Z(n2191) );
  XNOR U2334 ( .A(b[1]), .B(n2191), .Z(n2193) );
  NANDN U2335 ( .A(b[0]), .B(a[56]), .Z(n2192) );
  NAND U2336 ( .A(n2193), .B(n2192), .Z(n2238) );
  XNOR U2337 ( .A(n2237), .B(n2238), .Z(n2243) );
  XOR U2338 ( .A(n2244), .B(n2243), .Z(n2218) );
  NANDN U2339 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U2340 ( .A(n2197), .B(n2196), .Z(n2198) );
  AND U2341 ( .A(n2199), .B(n2198), .Z(n2217) );
  XNOR U2342 ( .A(n2218), .B(n2217), .Z(n2219) );
  NANDN U2343 ( .A(n2201), .B(n2200), .Z(n2205) );
  NAND U2344 ( .A(n2203), .B(n2202), .Z(n2204) );
  NAND U2345 ( .A(n2205), .B(n2204), .Z(n2220) );
  XNOR U2346 ( .A(n2219), .B(n2220), .Z(n2211) );
  XNOR U2347 ( .A(n2212), .B(n2211), .Z(n2213) );
  XNOR U2348 ( .A(n2214), .B(n2213), .Z(n2247) );
  XNOR U2349 ( .A(sreg[177]), .B(n2247), .Z(n2249) );
  NANDN U2350 ( .A(sreg[176]), .B(n2206), .Z(n2210) );
  NAND U2351 ( .A(n2208), .B(n2207), .Z(n2209) );
  NAND U2352 ( .A(n2210), .B(n2209), .Z(n2248) );
  XNOR U2353 ( .A(n2249), .B(n2248), .Z(c[177]) );
  NANDN U2354 ( .A(n2212), .B(n2211), .Z(n2216) );
  NANDN U2355 ( .A(n2214), .B(n2213), .Z(n2215) );
  AND U2356 ( .A(n2216), .B(n2215), .Z(n2255) );
  NANDN U2357 ( .A(n2218), .B(n2217), .Z(n2222) );
  NANDN U2358 ( .A(n2220), .B(n2219), .Z(n2221) );
  AND U2359 ( .A(n2222), .B(n2221), .Z(n2253) );
  NANDN U2360 ( .A(n5274), .B(n2223), .Z(n2225) );
  XOR U2361 ( .A(b[7]), .B(a[52]), .Z(n2264) );
  NANDN U2362 ( .A(n5275), .B(n2264), .Z(n2224) );
  AND U2363 ( .A(n2225), .B(n2224), .Z(n2283) );
  NANDN U2364 ( .A(n5176), .B(n2226), .Z(n2228) );
  XOR U2365 ( .A(b[3]), .B(a[56]), .Z(n2267) );
  NANDN U2366 ( .A(n5177), .B(n2267), .Z(n2227) );
  NAND U2367 ( .A(n2228), .B(n2227), .Z(n2282) );
  XNOR U2368 ( .A(n2283), .B(n2282), .Z(n2285) );
  NAND U2369 ( .A(b[0]), .B(a[58]), .Z(n2229) );
  XNOR U2370 ( .A(b[1]), .B(n2229), .Z(n2231) );
  NANDN U2371 ( .A(b[0]), .B(a[57]), .Z(n2230) );
  NAND U2372 ( .A(n2231), .B(n2230), .Z(n2279) );
  NANDN U2373 ( .A(n5249), .B(n2232), .Z(n2234) );
  XOR U2374 ( .A(b[5]), .B(a[54]), .Z(n2270) );
  NANDN U2375 ( .A(n5184), .B(n2270), .Z(n2233) );
  AND U2376 ( .A(n2234), .B(n2233), .Z(n2277) );
  AND U2377 ( .A(b[7]), .B(a[50]), .Z(n2276) );
  XNOR U2378 ( .A(n2277), .B(n2276), .Z(n2278) );
  XNOR U2379 ( .A(n2279), .B(n2278), .Z(n2284) );
  XOR U2380 ( .A(n2285), .B(n2284), .Z(n2259) );
  NANDN U2381 ( .A(n2236), .B(n2235), .Z(n2240) );
  NANDN U2382 ( .A(n2238), .B(n2237), .Z(n2239) );
  AND U2383 ( .A(n2240), .B(n2239), .Z(n2258) );
  XNOR U2384 ( .A(n2259), .B(n2258), .Z(n2260) );
  NANDN U2385 ( .A(n2242), .B(n2241), .Z(n2246) );
  NAND U2386 ( .A(n2244), .B(n2243), .Z(n2245) );
  NAND U2387 ( .A(n2246), .B(n2245), .Z(n2261) );
  XNOR U2388 ( .A(n2260), .B(n2261), .Z(n2252) );
  XNOR U2389 ( .A(n2253), .B(n2252), .Z(n2254) );
  XNOR U2390 ( .A(n2255), .B(n2254), .Z(n2288) );
  XNOR U2391 ( .A(sreg[178]), .B(n2288), .Z(n2290) );
  NANDN U2392 ( .A(sreg[177]), .B(n2247), .Z(n2251) );
  NAND U2393 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2394 ( .A(n2251), .B(n2250), .Z(n2289) );
  XNOR U2395 ( .A(n2290), .B(n2289), .Z(c[178]) );
  NANDN U2396 ( .A(n2253), .B(n2252), .Z(n2257) );
  NANDN U2397 ( .A(n2255), .B(n2254), .Z(n2256) );
  AND U2398 ( .A(n2257), .B(n2256), .Z(n2296) );
  NANDN U2399 ( .A(n2259), .B(n2258), .Z(n2263) );
  NANDN U2400 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U2401 ( .A(n2263), .B(n2262), .Z(n2294) );
  NANDN U2402 ( .A(n5274), .B(n2264), .Z(n2266) );
  XOR U2403 ( .A(b[7]), .B(a[53]), .Z(n2305) );
  NANDN U2404 ( .A(n5275), .B(n2305), .Z(n2265) );
  AND U2405 ( .A(n2266), .B(n2265), .Z(n2324) );
  NANDN U2406 ( .A(n5176), .B(n2267), .Z(n2269) );
  XOR U2407 ( .A(b[3]), .B(a[57]), .Z(n2308) );
  NANDN U2408 ( .A(n5177), .B(n2308), .Z(n2268) );
  NAND U2409 ( .A(n2269), .B(n2268), .Z(n2323) );
  XNOR U2410 ( .A(n2324), .B(n2323), .Z(n2326) );
  NANDN U2411 ( .A(n5249), .B(n2270), .Z(n2272) );
  XOR U2412 ( .A(b[5]), .B(a[55]), .Z(n2311) );
  NANDN U2413 ( .A(n5184), .B(n2311), .Z(n2271) );
  AND U2414 ( .A(n2272), .B(n2271), .Z(n2318) );
  AND U2415 ( .A(b[7]), .B(a[51]), .Z(n2317) );
  XNOR U2416 ( .A(n2318), .B(n2317), .Z(n2319) );
  NAND U2417 ( .A(b[0]), .B(a[59]), .Z(n2273) );
  XNOR U2418 ( .A(b[1]), .B(n2273), .Z(n2275) );
  NANDN U2419 ( .A(b[0]), .B(a[58]), .Z(n2274) );
  NAND U2420 ( .A(n2275), .B(n2274), .Z(n2320) );
  XNOR U2421 ( .A(n2319), .B(n2320), .Z(n2325) );
  XOR U2422 ( .A(n2326), .B(n2325), .Z(n2300) );
  NANDN U2423 ( .A(n2277), .B(n2276), .Z(n2281) );
  NANDN U2424 ( .A(n2279), .B(n2278), .Z(n2280) );
  AND U2425 ( .A(n2281), .B(n2280), .Z(n2299) );
  XNOR U2426 ( .A(n2300), .B(n2299), .Z(n2301) );
  NANDN U2427 ( .A(n2283), .B(n2282), .Z(n2287) );
  NAND U2428 ( .A(n2285), .B(n2284), .Z(n2286) );
  NAND U2429 ( .A(n2287), .B(n2286), .Z(n2302) );
  XNOR U2430 ( .A(n2301), .B(n2302), .Z(n2293) );
  XNOR U2431 ( .A(n2294), .B(n2293), .Z(n2295) );
  XNOR U2432 ( .A(n2296), .B(n2295), .Z(n2329) );
  XNOR U2433 ( .A(sreg[179]), .B(n2329), .Z(n2331) );
  NANDN U2434 ( .A(sreg[178]), .B(n2288), .Z(n2292) );
  NAND U2435 ( .A(n2290), .B(n2289), .Z(n2291) );
  NAND U2436 ( .A(n2292), .B(n2291), .Z(n2330) );
  XNOR U2437 ( .A(n2331), .B(n2330), .Z(c[179]) );
  NANDN U2438 ( .A(n2294), .B(n2293), .Z(n2298) );
  NANDN U2439 ( .A(n2296), .B(n2295), .Z(n2297) );
  AND U2440 ( .A(n2298), .B(n2297), .Z(n2337) );
  NANDN U2441 ( .A(n2300), .B(n2299), .Z(n2304) );
  NANDN U2442 ( .A(n2302), .B(n2301), .Z(n2303) );
  AND U2443 ( .A(n2304), .B(n2303), .Z(n2335) );
  NANDN U2444 ( .A(n5274), .B(n2305), .Z(n2307) );
  XOR U2445 ( .A(b[7]), .B(a[54]), .Z(n2346) );
  NANDN U2446 ( .A(n5275), .B(n2346), .Z(n2306) );
  AND U2447 ( .A(n2307), .B(n2306), .Z(n2365) );
  NANDN U2448 ( .A(n5176), .B(n2308), .Z(n2310) );
  XOR U2449 ( .A(b[3]), .B(a[58]), .Z(n2349) );
  NANDN U2450 ( .A(n5177), .B(n2349), .Z(n2309) );
  NAND U2451 ( .A(n2310), .B(n2309), .Z(n2364) );
  XNOR U2452 ( .A(n2365), .B(n2364), .Z(n2367) );
  NANDN U2453 ( .A(n5249), .B(n2311), .Z(n2313) );
  XOR U2454 ( .A(b[5]), .B(a[56]), .Z(n2355) );
  NANDN U2455 ( .A(n5184), .B(n2355), .Z(n2312) );
  AND U2456 ( .A(n2313), .B(n2312), .Z(n2359) );
  AND U2457 ( .A(b[7]), .B(a[52]), .Z(n2358) );
  XNOR U2458 ( .A(n2359), .B(n2358), .Z(n2360) );
  NAND U2459 ( .A(b[0]), .B(a[60]), .Z(n2314) );
  XNOR U2460 ( .A(b[1]), .B(n2314), .Z(n2316) );
  NANDN U2461 ( .A(b[0]), .B(a[59]), .Z(n2315) );
  NAND U2462 ( .A(n2316), .B(n2315), .Z(n2361) );
  XNOR U2463 ( .A(n2360), .B(n2361), .Z(n2366) );
  XOR U2464 ( .A(n2367), .B(n2366), .Z(n2341) );
  NANDN U2465 ( .A(n2318), .B(n2317), .Z(n2322) );
  NANDN U2466 ( .A(n2320), .B(n2319), .Z(n2321) );
  AND U2467 ( .A(n2322), .B(n2321), .Z(n2340) );
  XNOR U2468 ( .A(n2341), .B(n2340), .Z(n2342) );
  NANDN U2469 ( .A(n2324), .B(n2323), .Z(n2328) );
  NAND U2470 ( .A(n2326), .B(n2325), .Z(n2327) );
  NAND U2471 ( .A(n2328), .B(n2327), .Z(n2343) );
  XNOR U2472 ( .A(n2342), .B(n2343), .Z(n2334) );
  XNOR U2473 ( .A(n2335), .B(n2334), .Z(n2336) );
  XNOR U2474 ( .A(n2337), .B(n2336), .Z(n2370) );
  XNOR U2475 ( .A(sreg[180]), .B(n2370), .Z(n2372) );
  NANDN U2476 ( .A(sreg[179]), .B(n2329), .Z(n2333) );
  NAND U2477 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U2478 ( .A(n2333), .B(n2332), .Z(n2371) );
  XNOR U2479 ( .A(n2372), .B(n2371), .Z(c[180]) );
  NANDN U2480 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U2481 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U2482 ( .A(n2339), .B(n2338), .Z(n2382) );
  NANDN U2483 ( .A(n2341), .B(n2340), .Z(n2345) );
  NANDN U2484 ( .A(n2343), .B(n2342), .Z(n2344) );
  AND U2485 ( .A(n2345), .B(n2344), .Z(n2381) );
  NANDN U2486 ( .A(n5274), .B(n2346), .Z(n2348) );
  XOR U2487 ( .A(b[7]), .B(a[55]), .Z(n2392) );
  NANDN U2488 ( .A(n5275), .B(n2392), .Z(n2347) );
  AND U2489 ( .A(n2348), .B(n2347), .Z(n2411) );
  NANDN U2490 ( .A(n5176), .B(n2349), .Z(n2351) );
  XOR U2491 ( .A(b[3]), .B(a[59]), .Z(n2395) );
  NANDN U2492 ( .A(n5177), .B(n2395), .Z(n2350) );
  NAND U2493 ( .A(n2351), .B(n2350), .Z(n2410) );
  XNOR U2494 ( .A(n2411), .B(n2410), .Z(n2413) );
  NAND U2495 ( .A(b[0]), .B(a[61]), .Z(n2352) );
  XNOR U2496 ( .A(b[1]), .B(n2352), .Z(n2354) );
  NANDN U2497 ( .A(b[0]), .B(a[60]), .Z(n2353) );
  NAND U2498 ( .A(n2354), .B(n2353), .Z(n2407) );
  NANDN U2499 ( .A(n5249), .B(n2355), .Z(n2357) );
  XOR U2500 ( .A(b[5]), .B(a[57]), .Z(n2401) );
  NANDN U2501 ( .A(n5184), .B(n2401), .Z(n2356) );
  AND U2502 ( .A(n2357), .B(n2356), .Z(n2405) );
  AND U2503 ( .A(b[7]), .B(a[53]), .Z(n2404) );
  XNOR U2504 ( .A(n2405), .B(n2404), .Z(n2406) );
  XNOR U2505 ( .A(n2407), .B(n2406), .Z(n2412) );
  XOR U2506 ( .A(n2413), .B(n2412), .Z(n2387) );
  NANDN U2507 ( .A(n2359), .B(n2358), .Z(n2363) );
  NANDN U2508 ( .A(n2361), .B(n2360), .Z(n2362) );
  AND U2509 ( .A(n2363), .B(n2362), .Z(n2386) );
  XNOR U2510 ( .A(n2387), .B(n2386), .Z(n2388) );
  NANDN U2511 ( .A(n2365), .B(n2364), .Z(n2369) );
  NAND U2512 ( .A(n2367), .B(n2366), .Z(n2368) );
  NAND U2513 ( .A(n2369), .B(n2368), .Z(n2389) );
  XNOR U2514 ( .A(n2388), .B(n2389), .Z(n2380) );
  XOR U2515 ( .A(n2381), .B(n2380), .Z(n2383) );
  XOR U2516 ( .A(n2382), .B(n2383), .Z(n2375) );
  XNOR U2517 ( .A(n2375), .B(sreg[181]), .Z(n2377) );
  NANDN U2518 ( .A(sreg[180]), .B(n2370), .Z(n2374) );
  NAND U2519 ( .A(n2372), .B(n2371), .Z(n2373) );
  AND U2520 ( .A(n2374), .B(n2373), .Z(n2376) );
  XOR U2521 ( .A(n2377), .B(n2376), .Z(c[181]) );
  NANDN U2522 ( .A(n2375), .B(sreg[181]), .Z(n2379) );
  NAND U2523 ( .A(n2377), .B(n2376), .Z(n2378) );
  AND U2524 ( .A(n2379), .B(n2378), .Z(n2454) );
  NANDN U2525 ( .A(n2381), .B(n2380), .Z(n2385) );
  OR U2526 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U2527 ( .A(n2385), .B(n2384), .Z(n2419) );
  NANDN U2528 ( .A(n2387), .B(n2386), .Z(n2391) );
  NANDN U2529 ( .A(n2389), .B(n2388), .Z(n2390) );
  AND U2530 ( .A(n2391), .B(n2390), .Z(n2417) );
  NANDN U2531 ( .A(n5274), .B(n2392), .Z(n2394) );
  XOR U2532 ( .A(b[7]), .B(a[56]), .Z(n2428) );
  NANDN U2533 ( .A(n5275), .B(n2428), .Z(n2393) );
  AND U2534 ( .A(n2394), .B(n2393), .Z(n2447) );
  NANDN U2535 ( .A(n5176), .B(n2395), .Z(n2397) );
  XOR U2536 ( .A(b[3]), .B(a[60]), .Z(n2431) );
  NANDN U2537 ( .A(n5177), .B(n2431), .Z(n2396) );
  NAND U2538 ( .A(n2397), .B(n2396), .Z(n2446) );
  XNOR U2539 ( .A(n2447), .B(n2446), .Z(n2449) );
  NAND U2540 ( .A(b[0]), .B(a[62]), .Z(n2398) );
  XNOR U2541 ( .A(b[1]), .B(n2398), .Z(n2400) );
  NANDN U2542 ( .A(b[0]), .B(a[61]), .Z(n2399) );
  NAND U2543 ( .A(n2400), .B(n2399), .Z(n2443) );
  NANDN U2544 ( .A(n5249), .B(n2401), .Z(n2403) );
  XOR U2545 ( .A(b[5]), .B(a[58]), .Z(n2437) );
  NANDN U2546 ( .A(n5184), .B(n2437), .Z(n2402) );
  AND U2547 ( .A(n2403), .B(n2402), .Z(n2441) );
  AND U2548 ( .A(b[7]), .B(a[54]), .Z(n2440) );
  XNOR U2549 ( .A(n2441), .B(n2440), .Z(n2442) );
  XNOR U2550 ( .A(n2443), .B(n2442), .Z(n2448) );
  XOR U2551 ( .A(n2449), .B(n2448), .Z(n2423) );
  NANDN U2552 ( .A(n2405), .B(n2404), .Z(n2409) );
  NANDN U2553 ( .A(n2407), .B(n2406), .Z(n2408) );
  AND U2554 ( .A(n2409), .B(n2408), .Z(n2422) );
  XNOR U2555 ( .A(n2423), .B(n2422), .Z(n2424) );
  NANDN U2556 ( .A(n2411), .B(n2410), .Z(n2415) );
  NAND U2557 ( .A(n2413), .B(n2412), .Z(n2414) );
  NAND U2558 ( .A(n2415), .B(n2414), .Z(n2425) );
  XNOR U2559 ( .A(n2424), .B(n2425), .Z(n2416) );
  XNOR U2560 ( .A(n2417), .B(n2416), .Z(n2418) );
  XNOR U2561 ( .A(n2419), .B(n2418), .Z(n2452) );
  XNOR U2562 ( .A(sreg[182]), .B(n2452), .Z(n2453) );
  XNOR U2563 ( .A(n2454), .B(n2453), .Z(c[182]) );
  NANDN U2564 ( .A(n2417), .B(n2416), .Z(n2421) );
  NANDN U2565 ( .A(n2419), .B(n2418), .Z(n2420) );
  AND U2566 ( .A(n2421), .B(n2420), .Z(n2460) );
  NANDN U2567 ( .A(n2423), .B(n2422), .Z(n2427) );
  NANDN U2568 ( .A(n2425), .B(n2424), .Z(n2426) );
  AND U2569 ( .A(n2427), .B(n2426), .Z(n2458) );
  NANDN U2570 ( .A(n5274), .B(n2428), .Z(n2430) );
  XOR U2571 ( .A(b[7]), .B(a[57]), .Z(n2469) );
  NANDN U2572 ( .A(n5275), .B(n2469), .Z(n2429) );
  AND U2573 ( .A(n2430), .B(n2429), .Z(n2488) );
  NANDN U2574 ( .A(n5176), .B(n2431), .Z(n2433) );
  XOR U2575 ( .A(b[3]), .B(a[61]), .Z(n2472) );
  NANDN U2576 ( .A(n5177), .B(n2472), .Z(n2432) );
  NAND U2577 ( .A(n2433), .B(n2432), .Z(n2487) );
  XNOR U2578 ( .A(n2488), .B(n2487), .Z(n2490) );
  NAND U2579 ( .A(b[0]), .B(a[63]), .Z(n2434) );
  XNOR U2580 ( .A(b[1]), .B(n2434), .Z(n2436) );
  NANDN U2581 ( .A(b[0]), .B(a[62]), .Z(n2435) );
  NAND U2582 ( .A(n2436), .B(n2435), .Z(n2484) );
  NANDN U2583 ( .A(n5249), .B(n2437), .Z(n2439) );
  XOR U2584 ( .A(b[5]), .B(a[59]), .Z(n2475) );
  NANDN U2585 ( .A(n5184), .B(n2475), .Z(n2438) );
  AND U2586 ( .A(n2439), .B(n2438), .Z(n2482) );
  AND U2587 ( .A(b[7]), .B(a[55]), .Z(n2481) );
  XNOR U2588 ( .A(n2482), .B(n2481), .Z(n2483) );
  XNOR U2589 ( .A(n2484), .B(n2483), .Z(n2489) );
  XOR U2590 ( .A(n2490), .B(n2489), .Z(n2464) );
  NANDN U2591 ( .A(n2441), .B(n2440), .Z(n2445) );
  NANDN U2592 ( .A(n2443), .B(n2442), .Z(n2444) );
  AND U2593 ( .A(n2445), .B(n2444), .Z(n2463) );
  XNOR U2594 ( .A(n2464), .B(n2463), .Z(n2465) );
  NANDN U2595 ( .A(n2447), .B(n2446), .Z(n2451) );
  NAND U2596 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U2597 ( .A(n2451), .B(n2450), .Z(n2466) );
  XNOR U2598 ( .A(n2465), .B(n2466), .Z(n2457) );
  XNOR U2599 ( .A(n2458), .B(n2457), .Z(n2459) );
  XNOR U2600 ( .A(n2460), .B(n2459), .Z(n2493) );
  XNOR U2601 ( .A(sreg[183]), .B(n2493), .Z(n2495) );
  NANDN U2602 ( .A(sreg[182]), .B(n2452), .Z(n2456) );
  NAND U2603 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U2604 ( .A(n2456), .B(n2455), .Z(n2494) );
  XNOR U2605 ( .A(n2495), .B(n2494), .Z(c[183]) );
  NANDN U2606 ( .A(n2458), .B(n2457), .Z(n2462) );
  NANDN U2607 ( .A(n2460), .B(n2459), .Z(n2461) );
  AND U2608 ( .A(n2462), .B(n2461), .Z(n2501) );
  NANDN U2609 ( .A(n2464), .B(n2463), .Z(n2468) );
  NANDN U2610 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2611 ( .A(n2468), .B(n2467), .Z(n2499) );
  NANDN U2612 ( .A(n5274), .B(n2469), .Z(n2471) );
  XOR U2613 ( .A(b[7]), .B(a[58]), .Z(n2510) );
  NANDN U2614 ( .A(n5275), .B(n2510), .Z(n2470) );
  AND U2615 ( .A(n2471), .B(n2470), .Z(n2529) );
  NANDN U2616 ( .A(n5176), .B(n2472), .Z(n2474) );
  XOR U2617 ( .A(b[3]), .B(a[62]), .Z(n2513) );
  NANDN U2618 ( .A(n5177), .B(n2513), .Z(n2473) );
  NAND U2619 ( .A(n2474), .B(n2473), .Z(n2528) );
  XNOR U2620 ( .A(n2529), .B(n2528), .Z(n2531) );
  NANDN U2621 ( .A(n5249), .B(n2475), .Z(n2477) );
  XOR U2622 ( .A(b[5]), .B(a[60]), .Z(n2516) );
  NANDN U2623 ( .A(n5184), .B(n2516), .Z(n2476) );
  AND U2624 ( .A(n2477), .B(n2476), .Z(n2523) );
  AND U2625 ( .A(b[7]), .B(a[56]), .Z(n2522) );
  XNOR U2626 ( .A(n2523), .B(n2522), .Z(n2524) );
  NAND U2627 ( .A(b[0]), .B(a[64]), .Z(n2478) );
  XNOR U2628 ( .A(b[1]), .B(n2478), .Z(n2480) );
  NANDN U2629 ( .A(b[0]), .B(a[63]), .Z(n2479) );
  NAND U2630 ( .A(n2480), .B(n2479), .Z(n2525) );
  XNOR U2631 ( .A(n2524), .B(n2525), .Z(n2530) );
  XOR U2632 ( .A(n2531), .B(n2530), .Z(n2505) );
  NANDN U2633 ( .A(n2482), .B(n2481), .Z(n2486) );
  NANDN U2634 ( .A(n2484), .B(n2483), .Z(n2485) );
  AND U2635 ( .A(n2486), .B(n2485), .Z(n2504) );
  XNOR U2636 ( .A(n2505), .B(n2504), .Z(n2506) );
  NANDN U2637 ( .A(n2488), .B(n2487), .Z(n2492) );
  NAND U2638 ( .A(n2490), .B(n2489), .Z(n2491) );
  NAND U2639 ( .A(n2492), .B(n2491), .Z(n2507) );
  XNOR U2640 ( .A(n2506), .B(n2507), .Z(n2498) );
  XNOR U2641 ( .A(n2499), .B(n2498), .Z(n2500) );
  XNOR U2642 ( .A(n2501), .B(n2500), .Z(n2534) );
  XNOR U2643 ( .A(sreg[184]), .B(n2534), .Z(n2536) );
  NANDN U2644 ( .A(sreg[183]), .B(n2493), .Z(n2497) );
  NAND U2645 ( .A(n2495), .B(n2494), .Z(n2496) );
  NAND U2646 ( .A(n2497), .B(n2496), .Z(n2535) );
  XNOR U2647 ( .A(n2536), .B(n2535), .Z(c[184]) );
  NANDN U2648 ( .A(n2499), .B(n2498), .Z(n2503) );
  NANDN U2649 ( .A(n2501), .B(n2500), .Z(n2502) );
  AND U2650 ( .A(n2503), .B(n2502), .Z(n2542) );
  NANDN U2651 ( .A(n2505), .B(n2504), .Z(n2509) );
  NANDN U2652 ( .A(n2507), .B(n2506), .Z(n2508) );
  AND U2653 ( .A(n2509), .B(n2508), .Z(n2540) );
  NANDN U2654 ( .A(n5274), .B(n2510), .Z(n2512) );
  XOR U2655 ( .A(b[7]), .B(a[59]), .Z(n2551) );
  NANDN U2656 ( .A(n5275), .B(n2551), .Z(n2511) );
  AND U2657 ( .A(n2512), .B(n2511), .Z(n2570) );
  NANDN U2658 ( .A(n5176), .B(n2513), .Z(n2515) );
  XOR U2659 ( .A(b[3]), .B(a[63]), .Z(n2554) );
  NANDN U2660 ( .A(n5177), .B(n2554), .Z(n2514) );
  NAND U2661 ( .A(n2515), .B(n2514), .Z(n2569) );
  XNOR U2662 ( .A(n2570), .B(n2569), .Z(n2572) );
  NANDN U2663 ( .A(n5249), .B(n2516), .Z(n2518) );
  XOR U2664 ( .A(b[5]), .B(a[61]), .Z(n2560) );
  NANDN U2665 ( .A(n5184), .B(n2560), .Z(n2517) );
  AND U2666 ( .A(n2518), .B(n2517), .Z(n2564) );
  AND U2667 ( .A(b[7]), .B(a[57]), .Z(n2563) );
  XNOR U2668 ( .A(n2564), .B(n2563), .Z(n2565) );
  NAND U2669 ( .A(b[0]), .B(a[65]), .Z(n2519) );
  XNOR U2670 ( .A(b[1]), .B(n2519), .Z(n2521) );
  NANDN U2671 ( .A(b[0]), .B(a[64]), .Z(n2520) );
  NAND U2672 ( .A(n2521), .B(n2520), .Z(n2566) );
  XNOR U2673 ( .A(n2565), .B(n2566), .Z(n2571) );
  XOR U2674 ( .A(n2572), .B(n2571), .Z(n2546) );
  NANDN U2675 ( .A(n2523), .B(n2522), .Z(n2527) );
  NANDN U2676 ( .A(n2525), .B(n2524), .Z(n2526) );
  AND U2677 ( .A(n2527), .B(n2526), .Z(n2545) );
  XNOR U2678 ( .A(n2546), .B(n2545), .Z(n2547) );
  NANDN U2679 ( .A(n2529), .B(n2528), .Z(n2533) );
  NAND U2680 ( .A(n2531), .B(n2530), .Z(n2532) );
  NAND U2681 ( .A(n2533), .B(n2532), .Z(n2548) );
  XNOR U2682 ( .A(n2547), .B(n2548), .Z(n2539) );
  XNOR U2683 ( .A(n2540), .B(n2539), .Z(n2541) );
  XNOR U2684 ( .A(n2542), .B(n2541), .Z(n2575) );
  XNOR U2685 ( .A(sreg[185]), .B(n2575), .Z(n2577) );
  NANDN U2686 ( .A(sreg[184]), .B(n2534), .Z(n2538) );
  NAND U2687 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U2688 ( .A(n2538), .B(n2537), .Z(n2576) );
  XNOR U2689 ( .A(n2577), .B(n2576), .Z(c[185]) );
  NANDN U2690 ( .A(n2540), .B(n2539), .Z(n2544) );
  NANDN U2691 ( .A(n2542), .B(n2541), .Z(n2543) );
  AND U2692 ( .A(n2544), .B(n2543), .Z(n2583) );
  NANDN U2693 ( .A(n2546), .B(n2545), .Z(n2550) );
  NANDN U2694 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U2695 ( .A(n2550), .B(n2549), .Z(n2581) );
  NANDN U2696 ( .A(n5274), .B(n2551), .Z(n2553) );
  XOR U2697 ( .A(b[7]), .B(a[60]), .Z(n2592) );
  NANDN U2698 ( .A(n5275), .B(n2592), .Z(n2552) );
  AND U2699 ( .A(n2553), .B(n2552), .Z(n2611) );
  NANDN U2700 ( .A(n5176), .B(n2554), .Z(n2556) );
  XOR U2701 ( .A(b[3]), .B(a[64]), .Z(n2595) );
  NANDN U2702 ( .A(n5177), .B(n2595), .Z(n2555) );
  NAND U2703 ( .A(n2556), .B(n2555), .Z(n2610) );
  XNOR U2704 ( .A(n2611), .B(n2610), .Z(n2613) );
  NAND U2705 ( .A(b[0]), .B(a[66]), .Z(n2557) );
  XNOR U2706 ( .A(b[1]), .B(n2557), .Z(n2559) );
  NANDN U2707 ( .A(b[0]), .B(a[65]), .Z(n2558) );
  NAND U2708 ( .A(n2559), .B(n2558), .Z(n2607) );
  NANDN U2709 ( .A(n5249), .B(n2560), .Z(n2562) );
  XOR U2710 ( .A(b[5]), .B(a[62]), .Z(n2601) );
  NANDN U2711 ( .A(n5184), .B(n2601), .Z(n2561) );
  AND U2712 ( .A(n2562), .B(n2561), .Z(n2605) );
  AND U2713 ( .A(b[7]), .B(a[58]), .Z(n2604) );
  XNOR U2714 ( .A(n2605), .B(n2604), .Z(n2606) );
  XNOR U2715 ( .A(n2607), .B(n2606), .Z(n2612) );
  XOR U2716 ( .A(n2613), .B(n2612), .Z(n2587) );
  NANDN U2717 ( .A(n2564), .B(n2563), .Z(n2568) );
  NANDN U2718 ( .A(n2566), .B(n2565), .Z(n2567) );
  AND U2719 ( .A(n2568), .B(n2567), .Z(n2586) );
  XNOR U2720 ( .A(n2587), .B(n2586), .Z(n2588) );
  NANDN U2721 ( .A(n2570), .B(n2569), .Z(n2574) );
  NAND U2722 ( .A(n2572), .B(n2571), .Z(n2573) );
  NAND U2723 ( .A(n2574), .B(n2573), .Z(n2589) );
  XNOR U2724 ( .A(n2588), .B(n2589), .Z(n2580) );
  XNOR U2725 ( .A(n2581), .B(n2580), .Z(n2582) );
  XNOR U2726 ( .A(n2583), .B(n2582), .Z(n2616) );
  XNOR U2727 ( .A(sreg[186]), .B(n2616), .Z(n2618) );
  NANDN U2728 ( .A(sreg[185]), .B(n2575), .Z(n2579) );
  NAND U2729 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U2730 ( .A(n2579), .B(n2578), .Z(n2617) );
  XNOR U2731 ( .A(n2618), .B(n2617), .Z(c[186]) );
  NANDN U2732 ( .A(n2581), .B(n2580), .Z(n2585) );
  NANDN U2733 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U2734 ( .A(n2585), .B(n2584), .Z(n2624) );
  NANDN U2735 ( .A(n2587), .B(n2586), .Z(n2591) );
  NANDN U2736 ( .A(n2589), .B(n2588), .Z(n2590) );
  AND U2737 ( .A(n2591), .B(n2590), .Z(n2622) );
  NANDN U2738 ( .A(n5274), .B(n2592), .Z(n2594) );
  XOR U2739 ( .A(b[7]), .B(a[61]), .Z(n2633) );
  NANDN U2740 ( .A(n5275), .B(n2633), .Z(n2593) );
  AND U2741 ( .A(n2594), .B(n2593), .Z(n2652) );
  NANDN U2742 ( .A(n5176), .B(n2595), .Z(n2597) );
  XOR U2743 ( .A(b[3]), .B(a[65]), .Z(n2636) );
  NANDN U2744 ( .A(n5177), .B(n2636), .Z(n2596) );
  NAND U2745 ( .A(n2597), .B(n2596), .Z(n2651) );
  XNOR U2746 ( .A(n2652), .B(n2651), .Z(n2654) );
  NAND U2747 ( .A(b[0]), .B(a[67]), .Z(n2598) );
  XNOR U2748 ( .A(b[1]), .B(n2598), .Z(n2600) );
  NANDN U2749 ( .A(b[0]), .B(a[66]), .Z(n2599) );
  NAND U2750 ( .A(n2600), .B(n2599), .Z(n2648) );
  NANDN U2751 ( .A(n5249), .B(n2601), .Z(n2603) );
  XOR U2752 ( .A(b[5]), .B(a[63]), .Z(n2639) );
  NANDN U2753 ( .A(n5184), .B(n2639), .Z(n2602) );
  AND U2754 ( .A(n2603), .B(n2602), .Z(n2646) );
  AND U2755 ( .A(b[7]), .B(a[59]), .Z(n2645) );
  XNOR U2756 ( .A(n2646), .B(n2645), .Z(n2647) );
  XNOR U2757 ( .A(n2648), .B(n2647), .Z(n2653) );
  XOR U2758 ( .A(n2654), .B(n2653), .Z(n2628) );
  NANDN U2759 ( .A(n2605), .B(n2604), .Z(n2609) );
  NANDN U2760 ( .A(n2607), .B(n2606), .Z(n2608) );
  AND U2761 ( .A(n2609), .B(n2608), .Z(n2627) );
  XNOR U2762 ( .A(n2628), .B(n2627), .Z(n2629) );
  NANDN U2763 ( .A(n2611), .B(n2610), .Z(n2615) );
  NAND U2764 ( .A(n2613), .B(n2612), .Z(n2614) );
  NAND U2765 ( .A(n2615), .B(n2614), .Z(n2630) );
  XNOR U2766 ( .A(n2629), .B(n2630), .Z(n2621) );
  XNOR U2767 ( .A(n2622), .B(n2621), .Z(n2623) );
  XNOR U2768 ( .A(n2624), .B(n2623), .Z(n2657) );
  XNOR U2769 ( .A(sreg[187]), .B(n2657), .Z(n2659) );
  NANDN U2770 ( .A(sreg[186]), .B(n2616), .Z(n2620) );
  NAND U2771 ( .A(n2618), .B(n2617), .Z(n2619) );
  NAND U2772 ( .A(n2620), .B(n2619), .Z(n2658) );
  XNOR U2773 ( .A(n2659), .B(n2658), .Z(c[187]) );
  NANDN U2774 ( .A(n2622), .B(n2621), .Z(n2626) );
  NANDN U2775 ( .A(n2624), .B(n2623), .Z(n2625) );
  AND U2776 ( .A(n2626), .B(n2625), .Z(n2665) );
  NANDN U2777 ( .A(n2628), .B(n2627), .Z(n2632) );
  NANDN U2778 ( .A(n2630), .B(n2629), .Z(n2631) );
  AND U2779 ( .A(n2632), .B(n2631), .Z(n2663) );
  NANDN U2780 ( .A(n5274), .B(n2633), .Z(n2635) );
  XOR U2781 ( .A(b[7]), .B(a[62]), .Z(n2674) );
  NANDN U2782 ( .A(n5275), .B(n2674), .Z(n2634) );
  AND U2783 ( .A(n2635), .B(n2634), .Z(n2693) );
  NANDN U2784 ( .A(n5176), .B(n2636), .Z(n2638) );
  XOR U2785 ( .A(b[3]), .B(a[66]), .Z(n2677) );
  NANDN U2786 ( .A(n5177), .B(n2677), .Z(n2637) );
  NAND U2787 ( .A(n2638), .B(n2637), .Z(n2692) );
  XNOR U2788 ( .A(n2693), .B(n2692), .Z(n2695) );
  NANDN U2789 ( .A(n5249), .B(n2639), .Z(n2641) );
  XOR U2790 ( .A(b[5]), .B(a[64]), .Z(n2683) );
  NANDN U2791 ( .A(n5184), .B(n2683), .Z(n2640) );
  AND U2792 ( .A(n2641), .B(n2640), .Z(n2687) );
  AND U2793 ( .A(b[7]), .B(a[60]), .Z(n2686) );
  XNOR U2794 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U2795 ( .A(b[0]), .B(a[68]), .Z(n2642) );
  XNOR U2796 ( .A(b[1]), .B(n2642), .Z(n2644) );
  NANDN U2797 ( .A(b[0]), .B(a[67]), .Z(n2643) );
  NAND U2798 ( .A(n2644), .B(n2643), .Z(n2689) );
  XNOR U2799 ( .A(n2688), .B(n2689), .Z(n2694) );
  XOR U2800 ( .A(n2695), .B(n2694), .Z(n2669) );
  NANDN U2801 ( .A(n2646), .B(n2645), .Z(n2650) );
  NANDN U2802 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U2803 ( .A(n2650), .B(n2649), .Z(n2668) );
  XNOR U2804 ( .A(n2669), .B(n2668), .Z(n2670) );
  NANDN U2805 ( .A(n2652), .B(n2651), .Z(n2656) );
  NAND U2806 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U2807 ( .A(n2656), .B(n2655), .Z(n2671) );
  XNOR U2808 ( .A(n2670), .B(n2671), .Z(n2662) );
  XNOR U2809 ( .A(n2663), .B(n2662), .Z(n2664) );
  XNOR U2810 ( .A(n2665), .B(n2664), .Z(n2698) );
  XNOR U2811 ( .A(sreg[188]), .B(n2698), .Z(n2700) );
  NANDN U2812 ( .A(sreg[187]), .B(n2657), .Z(n2661) );
  NAND U2813 ( .A(n2659), .B(n2658), .Z(n2660) );
  NAND U2814 ( .A(n2661), .B(n2660), .Z(n2699) );
  XNOR U2815 ( .A(n2700), .B(n2699), .Z(c[188]) );
  NANDN U2816 ( .A(n2663), .B(n2662), .Z(n2667) );
  NANDN U2817 ( .A(n2665), .B(n2664), .Z(n2666) );
  AND U2818 ( .A(n2667), .B(n2666), .Z(n2706) );
  NANDN U2819 ( .A(n2669), .B(n2668), .Z(n2673) );
  NANDN U2820 ( .A(n2671), .B(n2670), .Z(n2672) );
  AND U2821 ( .A(n2673), .B(n2672), .Z(n2704) );
  NANDN U2822 ( .A(n5274), .B(n2674), .Z(n2676) );
  XOR U2823 ( .A(b[7]), .B(a[63]), .Z(n2715) );
  NANDN U2824 ( .A(n5275), .B(n2715), .Z(n2675) );
  AND U2825 ( .A(n2676), .B(n2675), .Z(n2734) );
  NANDN U2826 ( .A(n5176), .B(n2677), .Z(n2679) );
  XOR U2827 ( .A(b[3]), .B(a[67]), .Z(n2718) );
  NANDN U2828 ( .A(n5177), .B(n2718), .Z(n2678) );
  NAND U2829 ( .A(n2679), .B(n2678), .Z(n2733) );
  XNOR U2830 ( .A(n2734), .B(n2733), .Z(n2736) );
  NAND U2831 ( .A(b[0]), .B(a[69]), .Z(n2680) );
  XNOR U2832 ( .A(b[1]), .B(n2680), .Z(n2682) );
  NANDN U2833 ( .A(b[0]), .B(a[68]), .Z(n2681) );
  NAND U2834 ( .A(n2682), .B(n2681), .Z(n2730) );
  NANDN U2835 ( .A(n5249), .B(n2683), .Z(n2685) );
  XOR U2836 ( .A(b[5]), .B(a[65]), .Z(n2721) );
  NANDN U2837 ( .A(n5184), .B(n2721), .Z(n2684) );
  AND U2838 ( .A(n2685), .B(n2684), .Z(n2728) );
  AND U2839 ( .A(b[7]), .B(a[61]), .Z(n2727) );
  XNOR U2840 ( .A(n2728), .B(n2727), .Z(n2729) );
  XNOR U2841 ( .A(n2730), .B(n2729), .Z(n2735) );
  XOR U2842 ( .A(n2736), .B(n2735), .Z(n2710) );
  NANDN U2843 ( .A(n2687), .B(n2686), .Z(n2691) );
  NANDN U2844 ( .A(n2689), .B(n2688), .Z(n2690) );
  AND U2845 ( .A(n2691), .B(n2690), .Z(n2709) );
  XNOR U2846 ( .A(n2710), .B(n2709), .Z(n2711) );
  NANDN U2847 ( .A(n2693), .B(n2692), .Z(n2697) );
  NAND U2848 ( .A(n2695), .B(n2694), .Z(n2696) );
  NAND U2849 ( .A(n2697), .B(n2696), .Z(n2712) );
  XNOR U2850 ( .A(n2711), .B(n2712), .Z(n2703) );
  XNOR U2851 ( .A(n2704), .B(n2703), .Z(n2705) );
  XNOR U2852 ( .A(n2706), .B(n2705), .Z(n2739) );
  XNOR U2853 ( .A(sreg[189]), .B(n2739), .Z(n2741) );
  NANDN U2854 ( .A(sreg[188]), .B(n2698), .Z(n2702) );
  NAND U2855 ( .A(n2700), .B(n2699), .Z(n2701) );
  NAND U2856 ( .A(n2702), .B(n2701), .Z(n2740) );
  XNOR U2857 ( .A(n2741), .B(n2740), .Z(c[189]) );
  NANDN U2858 ( .A(n2704), .B(n2703), .Z(n2708) );
  NANDN U2859 ( .A(n2706), .B(n2705), .Z(n2707) );
  AND U2860 ( .A(n2708), .B(n2707), .Z(n2747) );
  NANDN U2861 ( .A(n2710), .B(n2709), .Z(n2714) );
  NANDN U2862 ( .A(n2712), .B(n2711), .Z(n2713) );
  AND U2863 ( .A(n2714), .B(n2713), .Z(n2745) );
  NANDN U2864 ( .A(n5274), .B(n2715), .Z(n2717) );
  XOR U2865 ( .A(b[7]), .B(a[64]), .Z(n2756) );
  NANDN U2866 ( .A(n5275), .B(n2756), .Z(n2716) );
  AND U2867 ( .A(n2717), .B(n2716), .Z(n2775) );
  NANDN U2868 ( .A(n5176), .B(n2718), .Z(n2720) );
  XOR U2869 ( .A(b[3]), .B(a[68]), .Z(n2759) );
  NANDN U2870 ( .A(n5177), .B(n2759), .Z(n2719) );
  NAND U2871 ( .A(n2720), .B(n2719), .Z(n2774) );
  XNOR U2872 ( .A(n2775), .B(n2774), .Z(n2777) );
  NANDN U2873 ( .A(n5249), .B(n2721), .Z(n2723) );
  XOR U2874 ( .A(b[5]), .B(a[66]), .Z(n2762) );
  NANDN U2875 ( .A(n5184), .B(n2762), .Z(n2722) );
  AND U2876 ( .A(n2723), .B(n2722), .Z(n2769) );
  AND U2877 ( .A(b[7]), .B(a[62]), .Z(n2768) );
  XNOR U2878 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U2879 ( .A(b[0]), .B(a[70]), .Z(n2724) );
  XNOR U2880 ( .A(b[1]), .B(n2724), .Z(n2726) );
  NANDN U2881 ( .A(b[0]), .B(a[69]), .Z(n2725) );
  NAND U2882 ( .A(n2726), .B(n2725), .Z(n2771) );
  XNOR U2883 ( .A(n2770), .B(n2771), .Z(n2776) );
  XOR U2884 ( .A(n2777), .B(n2776), .Z(n2751) );
  NANDN U2885 ( .A(n2728), .B(n2727), .Z(n2732) );
  NANDN U2886 ( .A(n2730), .B(n2729), .Z(n2731) );
  AND U2887 ( .A(n2732), .B(n2731), .Z(n2750) );
  XNOR U2888 ( .A(n2751), .B(n2750), .Z(n2752) );
  NANDN U2889 ( .A(n2734), .B(n2733), .Z(n2738) );
  NAND U2890 ( .A(n2736), .B(n2735), .Z(n2737) );
  NAND U2891 ( .A(n2738), .B(n2737), .Z(n2753) );
  XNOR U2892 ( .A(n2752), .B(n2753), .Z(n2744) );
  XNOR U2893 ( .A(n2745), .B(n2744), .Z(n2746) );
  XNOR U2894 ( .A(n2747), .B(n2746), .Z(n2780) );
  XNOR U2895 ( .A(sreg[190]), .B(n2780), .Z(n2782) );
  NANDN U2896 ( .A(sreg[189]), .B(n2739), .Z(n2743) );
  NAND U2897 ( .A(n2741), .B(n2740), .Z(n2742) );
  NAND U2898 ( .A(n2743), .B(n2742), .Z(n2781) );
  XNOR U2899 ( .A(n2782), .B(n2781), .Z(c[190]) );
  NANDN U2900 ( .A(n2745), .B(n2744), .Z(n2749) );
  NANDN U2901 ( .A(n2747), .B(n2746), .Z(n2748) );
  AND U2902 ( .A(n2749), .B(n2748), .Z(n2788) );
  NANDN U2903 ( .A(n2751), .B(n2750), .Z(n2755) );
  NANDN U2904 ( .A(n2753), .B(n2752), .Z(n2754) );
  AND U2905 ( .A(n2755), .B(n2754), .Z(n2786) );
  NANDN U2906 ( .A(n5274), .B(n2756), .Z(n2758) );
  XOR U2907 ( .A(b[7]), .B(a[65]), .Z(n2797) );
  NANDN U2908 ( .A(n5275), .B(n2797), .Z(n2757) );
  AND U2909 ( .A(n2758), .B(n2757), .Z(n2816) );
  NANDN U2910 ( .A(n5176), .B(n2759), .Z(n2761) );
  XOR U2911 ( .A(b[3]), .B(a[69]), .Z(n2800) );
  NANDN U2912 ( .A(n5177), .B(n2800), .Z(n2760) );
  NAND U2913 ( .A(n2761), .B(n2760), .Z(n2815) );
  XNOR U2914 ( .A(n2816), .B(n2815), .Z(n2818) );
  NANDN U2915 ( .A(n5249), .B(n2762), .Z(n2764) );
  XOR U2916 ( .A(b[5]), .B(a[67]), .Z(n2806) );
  NANDN U2917 ( .A(n5184), .B(n2806), .Z(n2763) );
  AND U2918 ( .A(n2764), .B(n2763), .Z(n2810) );
  AND U2919 ( .A(b[7]), .B(a[63]), .Z(n2809) );
  XNOR U2920 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U2921 ( .A(b[0]), .B(a[71]), .Z(n2765) );
  XNOR U2922 ( .A(b[1]), .B(n2765), .Z(n2767) );
  NANDN U2923 ( .A(b[0]), .B(a[70]), .Z(n2766) );
  NAND U2924 ( .A(n2767), .B(n2766), .Z(n2812) );
  XNOR U2925 ( .A(n2811), .B(n2812), .Z(n2817) );
  XOR U2926 ( .A(n2818), .B(n2817), .Z(n2792) );
  NANDN U2927 ( .A(n2769), .B(n2768), .Z(n2773) );
  NANDN U2928 ( .A(n2771), .B(n2770), .Z(n2772) );
  AND U2929 ( .A(n2773), .B(n2772), .Z(n2791) );
  XNOR U2930 ( .A(n2792), .B(n2791), .Z(n2793) );
  NANDN U2931 ( .A(n2775), .B(n2774), .Z(n2779) );
  NAND U2932 ( .A(n2777), .B(n2776), .Z(n2778) );
  NAND U2933 ( .A(n2779), .B(n2778), .Z(n2794) );
  XNOR U2934 ( .A(n2793), .B(n2794), .Z(n2785) );
  XNOR U2935 ( .A(n2786), .B(n2785), .Z(n2787) );
  XNOR U2936 ( .A(n2788), .B(n2787), .Z(n2821) );
  XNOR U2937 ( .A(sreg[191]), .B(n2821), .Z(n2823) );
  NANDN U2938 ( .A(sreg[190]), .B(n2780), .Z(n2784) );
  NAND U2939 ( .A(n2782), .B(n2781), .Z(n2783) );
  NAND U2940 ( .A(n2784), .B(n2783), .Z(n2822) );
  XNOR U2941 ( .A(n2823), .B(n2822), .Z(c[191]) );
  NANDN U2942 ( .A(n2786), .B(n2785), .Z(n2790) );
  NANDN U2943 ( .A(n2788), .B(n2787), .Z(n2789) );
  AND U2944 ( .A(n2790), .B(n2789), .Z(n2829) );
  NANDN U2945 ( .A(n2792), .B(n2791), .Z(n2796) );
  NANDN U2946 ( .A(n2794), .B(n2793), .Z(n2795) );
  AND U2947 ( .A(n2796), .B(n2795), .Z(n2827) );
  NANDN U2948 ( .A(n5274), .B(n2797), .Z(n2799) );
  XOR U2949 ( .A(b[7]), .B(a[66]), .Z(n2838) );
  NANDN U2950 ( .A(n5275), .B(n2838), .Z(n2798) );
  AND U2951 ( .A(n2799), .B(n2798), .Z(n2857) );
  NANDN U2952 ( .A(n5176), .B(n2800), .Z(n2802) );
  XOR U2953 ( .A(b[3]), .B(a[70]), .Z(n2841) );
  NANDN U2954 ( .A(n5177), .B(n2841), .Z(n2801) );
  NAND U2955 ( .A(n2802), .B(n2801), .Z(n2856) );
  XNOR U2956 ( .A(n2857), .B(n2856), .Z(n2859) );
  NAND U2957 ( .A(b[0]), .B(a[72]), .Z(n2803) );
  XNOR U2958 ( .A(b[1]), .B(n2803), .Z(n2805) );
  NANDN U2959 ( .A(b[0]), .B(a[71]), .Z(n2804) );
  NAND U2960 ( .A(n2805), .B(n2804), .Z(n2853) );
  NANDN U2961 ( .A(n5249), .B(n2806), .Z(n2808) );
  XOR U2962 ( .A(b[5]), .B(a[68]), .Z(n2847) );
  NANDN U2963 ( .A(n5184), .B(n2847), .Z(n2807) );
  AND U2964 ( .A(n2808), .B(n2807), .Z(n2851) );
  AND U2965 ( .A(b[7]), .B(a[64]), .Z(n2850) );
  XNOR U2966 ( .A(n2851), .B(n2850), .Z(n2852) );
  XNOR U2967 ( .A(n2853), .B(n2852), .Z(n2858) );
  XOR U2968 ( .A(n2859), .B(n2858), .Z(n2833) );
  NANDN U2969 ( .A(n2810), .B(n2809), .Z(n2814) );
  NANDN U2970 ( .A(n2812), .B(n2811), .Z(n2813) );
  AND U2971 ( .A(n2814), .B(n2813), .Z(n2832) );
  XNOR U2972 ( .A(n2833), .B(n2832), .Z(n2834) );
  NANDN U2973 ( .A(n2816), .B(n2815), .Z(n2820) );
  NAND U2974 ( .A(n2818), .B(n2817), .Z(n2819) );
  NAND U2975 ( .A(n2820), .B(n2819), .Z(n2835) );
  XNOR U2976 ( .A(n2834), .B(n2835), .Z(n2826) );
  XNOR U2977 ( .A(n2827), .B(n2826), .Z(n2828) );
  XNOR U2978 ( .A(n2829), .B(n2828), .Z(n2862) );
  XNOR U2979 ( .A(sreg[192]), .B(n2862), .Z(n2864) );
  NANDN U2980 ( .A(sreg[191]), .B(n2821), .Z(n2825) );
  NAND U2981 ( .A(n2823), .B(n2822), .Z(n2824) );
  NAND U2982 ( .A(n2825), .B(n2824), .Z(n2863) );
  XNOR U2983 ( .A(n2864), .B(n2863), .Z(c[192]) );
  NANDN U2984 ( .A(n2827), .B(n2826), .Z(n2831) );
  NANDN U2985 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U2986 ( .A(n2831), .B(n2830), .Z(n2870) );
  NANDN U2987 ( .A(n2833), .B(n2832), .Z(n2837) );
  NANDN U2988 ( .A(n2835), .B(n2834), .Z(n2836) );
  AND U2989 ( .A(n2837), .B(n2836), .Z(n2868) );
  NANDN U2990 ( .A(n5274), .B(n2838), .Z(n2840) );
  XOR U2991 ( .A(b[7]), .B(a[67]), .Z(n2879) );
  NANDN U2992 ( .A(n5275), .B(n2879), .Z(n2839) );
  AND U2993 ( .A(n2840), .B(n2839), .Z(n2898) );
  NANDN U2994 ( .A(n5176), .B(n2841), .Z(n2843) );
  XOR U2995 ( .A(b[3]), .B(a[71]), .Z(n2882) );
  NANDN U2996 ( .A(n5177), .B(n2882), .Z(n2842) );
  NAND U2997 ( .A(n2843), .B(n2842), .Z(n2897) );
  XNOR U2998 ( .A(n2898), .B(n2897), .Z(n2900) );
  AND U2999 ( .A(b[0]), .B(a[73]), .Z(n2844) );
  XOR U3000 ( .A(b[1]), .B(n2844), .Z(n2846) );
  NANDN U3001 ( .A(b[0]), .B(a[72]), .Z(n2845) );
  AND U3002 ( .A(n2846), .B(n2845), .Z(n2893) );
  NANDN U3003 ( .A(n5249), .B(n2847), .Z(n2849) );
  XOR U3004 ( .A(b[5]), .B(a[69]), .Z(n2888) );
  NANDN U3005 ( .A(n5184), .B(n2888), .Z(n2848) );
  AND U3006 ( .A(n2849), .B(n2848), .Z(n2892) );
  AND U3007 ( .A(b[7]), .B(a[65]), .Z(n2891) );
  XOR U3008 ( .A(n2892), .B(n2891), .Z(n2894) );
  XNOR U3009 ( .A(n2893), .B(n2894), .Z(n2899) );
  XOR U3010 ( .A(n2900), .B(n2899), .Z(n2874) );
  NANDN U3011 ( .A(n2851), .B(n2850), .Z(n2855) );
  NANDN U3012 ( .A(n2853), .B(n2852), .Z(n2854) );
  AND U3013 ( .A(n2855), .B(n2854), .Z(n2873) );
  XNOR U3014 ( .A(n2874), .B(n2873), .Z(n2875) );
  NANDN U3015 ( .A(n2857), .B(n2856), .Z(n2861) );
  NAND U3016 ( .A(n2859), .B(n2858), .Z(n2860) );
  NAND U3017 ( .A(n2861), .B(n2860), .Z(n2876) );
  XNOR U3018 ( .A(n2875), .B(n2876), .Z(n2867) );
  XNOR U3019 ( .A(n2868), .B(n2867), .Z(n2869) );
  XNOR U3020 ( .A(n2870), .B(n2869), .Z(n2903) );
  XNOR U3021 ( .A(sreg[193]), .B(n2903), .Z(n2905) );
  NANDN U3022 ( .A(sreg[192]), .B(n2862), .Z(n2866) );
  NAND U3023 ( .A(n2864), .B(n2863), .Z(n2865) );
  NAND U3024 ( .A(n2866), .B(n2865), .Z(n2904) );
  XNOR U3025 ( .A(n2905), .B(n2904), .Z(c[193]) );
  NANDN U3026 ( .A(n2868), .B(n2867), .Z(n2872) );
  NANDN U3027 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3028 ( .A(n2872), .B(n2871), .Z(n2911) );
  NANDN U3029 ( .A(n2874), .B(n2873), .Z(n2878) );
  NANDN U3030 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U3031 ( .A(n2878), .B(n2877), .Z(n2909) );
  NANDN U3032 ( .A(n5274), .B(n2879), .Z(n2881) );
  XOR U3033 ( .A(b[7]), .B(a[68]), .Z(n2920) );
  NANDN U3034 ( .A(n5275), .B(n2920), .Z(n2880) );
  AND U3035 ( .A(n2881), .B(n2880), .Z(n2939) );
  NANDN U3036 ( .A(n5176), .B(n2882), .Z(n2884) );
  XOR U3037 ( .A(b[3]), .B(a[72]), .Z(n2923) );
  NANDN U3038 ( .A(n5177), .B(n2923), .Z(n2883) );
  NAND U3039 ( .A(n2884), .B(n2883), .Z(n2938) );
  XNOR U3040 ( .A(n2939), .B(n2938), .Z(n2941) );
  NAND U3041 ( .A(b[0]), .B(a[74]), .Z(n2885) );
  XNOR U3042 ( .A(b[1]), .B(n2885), .Z(n2887) );
  NANDN U3043 ( .A(b[0]), .B(a[73]), .Z(n2886) );
  NAND U3044 ( .A(n2887), .B(n2886), .Z(n2935) );
  NANDN U3045 ( .A(n5249), .B(n2888), .Z(n2890) );
  XOR U3046 ( .A(b[5]), .B(a[70]), .Z(n2929) );
  NANDN U3047 ( .A(n5184), .B(n2929), .Z(n2889) );
  AND U3048 ( .A(n2890), .B(n2889), .Z(n2933) );
  AND U3049 ( .A(b[7]), .B(a[66]), .Z(n2932) );
  XNOR U3050 ( .A(n2933), .B(n2932), .Z(n2934) );
  XNOR U3051 ( .A(n2935), .B(n2934), .Z(n2940) );
  XOR U3052 ( .A(n2941), .B(n2940), .Z(n2915) );
  NANDN U3053 ( .A(n2892), .B(n2891), .Z(n2896) );
  NANDN U3054 ( .A(n2894), .B(n2893), .Z(n2895) );
  AND U3055 ( .A(n2896), .B(n2895), .Z(n2914) );
  XNOR U3056 ( .A(n2915), .B(n2914), .Z(n2916) );
  NANDN U3057 ( .A(n2898), .B(n2897), .Z(n2902) );
  NAND U3058 ( .A(n2900), .B(n2899), .Z(n2901) );
  NAND U3059 ( .A(n2902), .B(n2901), .Z(n2917) );
  XNOR U3060 ( .A(n2916), .B(n2917), .Z(n2908) );
  XNOR U3061 ( .A(n2909), .B(n2908), .Z(n2910) );
  XNOR U3062 ( .A(n2911), .B(n2910), .Z(n2944) );
  XNOR U3063 ( .A(sreg[194]), .B(n2944), .Z(n2946) );
  NANDN U3064 ( .A(sreg[193]), .B(n2903), .Z(n2907) );
  NAND U3065 ( .A(n2905), .B(n2904), .Z(n2906) );
  NAND U3066 ( .A(n2907), .B(n2906), .Z(n2945) );
  XNOR U3067 ( .A(n2946), .B(n2945), .Z(c[194]) );
  NANDN U3068 ( .A(n2909), .B(n2908), .Z(n2913) );
  NANDN U3069 ( .A(n2911), .B(n2910), .Z(n2912) );
  AND U3070 ( .A(n2913), .B(n2912), .Z(n2952) );
  NANDN U3071 ( .A(n2915), .B(n2914), .Z(n2919) );
  NANDN U3072 ( .A(n2917), .B(n2916), .Z(n2918) );
  AND U3073 ( .A(n2919), .B(n2918), .Z(n2950) );
  NANDN U3074 ( .A(n5274), .B(n2920), .Z(n2922) );
  XOR U3075 ( .A(b[7]), .B(a[69]), .Z(n2961) );
  NANDN U3076 ( .A(n5275), .B(n2961), .Z(n2921) );
  AND U3077 ( .A(n2922), .B(n2921), .Z(n2980) );
  NANDN U3078 ( .A(n5176), .B(n2923), .Z(n2925) );
  XOR U3079 ( .A(b[3]), .B(a[73]), .Z(n2964) );
  NANDN U3080 ( .A(n5177), .B(n2964), .Z(n2924) );
  NAND U3081 ( .A(n2925), .B(n2924), .Z(n2979) );
  XNOR U3082 ( .A(n2980), .B(n2979), .Z(n2982) );
  NAND U3083 ( .A(b[0]), .B(a[75]), .Z(n2926) );
  XNOR U3084 ( .A(b[1]), .B(n2926), .Z(n2928) );
  NANDN U3085 ( .A(b[0]), .B(a[74]), .Z(n2927) );
  NAND U3086 ( .A(n2928), .B(n2927), .Z(n2976) );
  NANDN U3087 ( .A(n5249), .B(n2929), .Z(n2931) );
  XOR U3088 ( .A(b[5]), .B(a[71]), .Z(n2970) );
  NANDN U3089 ( .A(n5184), .B(n2970), .Z(n2930) );
  AND U3090 ( .A(n2931), .B(n2930), .Z(n2974) );
  AND U3091 ( .A(b[7]), .B(a[67]), .Z(n2973) );
  XNOR U3092 ( .A(n2974), .B(n2973), .Z(n2975) );
  XNOR U3093 ( .A(n2976), .B(n2975), .Z(n2981) );
  XOR U3094 ( .A(n2982), .B(n2981), .Z(n2956) );
  NANDN U3095 ( .A(n2933), .B(n2932), .Z(n2937) );
  NANDN U3096 ( .A(n2935), .B(n2934), .Z(n2936) );
  AND U3097 ( .A(n2937), .B(n2936), .Z(n2955) );
  XNOR U3098 ( .A(n2956), .B(n2955), .Z(n2957) );
  NANDN U3099 ( .A(n2939), .B(n2938), .Z(n2943) );
  NAND U3100 ( .A(n2941), .B(n2940), .Z(n2942) );
  NAND U3101 ( .A(n2943), .B(n2942), .Z(n2958) );
  XNOR U3102 ( .A(n2957), .B(n2958), .Z(n2949) );
  XNOR U3103 ( .A(n2950), .B(n2949), .Z(n2951) );
  XNOR U3104 ( .A(n2952), .B(n2951), .Z(n2985) );
  XNOR U3105 ( .A(sreg[195]), .B(n2985), .Z(n2987) );
  NANDN U3106 ( .A(sreg[194]), .B(n2944), .Z(n2948) );
  NAND U3107 ( .A(n2946), .B(n2945), .Z(n2947) );
  NAND U3108 ( .A(n2948), .B(n2947), .Z(n2986) );
  XNOR U3109 ( .A(n2987), .B(n2986), .Z(c[195]) );
  NANDN U3110 ( .A(n2950), .B(n2949), .Z(n2954) );
  NANDN U3111 ( .A(n2952), .B(n2951), .Z(n2953) );
  AND U3112 ( .A(n2954), .B(n2953), .Z(n2993) );
  NANDN U3113 ( .A(n2956), .B(n2955), .Z(n2960) );
  NANDN U3114 ( .A(n2958), .B(n2957), .Z(n2959) );
  AND U3115 ( .A(n2960), .B(n2959), .Z(n2991) );
  NANDN U3116 ( .A(n5274), .B(n2961), .Z(n2963) );
  XOR U3117 ( .A(b[7]), .B(a[70]), .Z(n3002) );
  NANDN U3118 ( .A(n5275), .B(n3002), .Z(n2962) );
  AND U3119 ( .A(n2963), .B(n2962), .Z(n3021) );
  NANDN U3120 ( .A(n5176), .B(n2964), .Z(n2966) );
  XOR U3121 ( .A(b[3]), .B(a[74]), .Z(n3005) );
  NANDN U3122 ( .A(n5177), .B(n3005), .Z(n2965) );
  NAND U3123 ( .A(n2966), .B(n2965), .Z(n3020) );
  XNOR U3124 ( .A(n3021), .B(n3020), .Z(n3023) );
  NAND U3125 ( .A(b[0]), .B(a[76]), .Z(n2967) );
  XNOR U3126 ( .A(b[1]), .B(n2967), .Z(n2969) );
  NANDN U3127 ( .A(b[0]), .B(a[75]), .Z(n2968) );
  NAND U3128 ( .A(n2969), .B(n2968), .Z(n3017) );
  NANDN U3129 ( .A(n5249), .B(n2970), .Z(n2972) );
  XOR U3130 ( .A(b[5]), .B(a[72]), .Z(n3011) );
  NANDN U3131 ( .A(n5184), .B(n3011), .Z(n2971) );
  AND U3132 ( .A(n2972), .B(n2971), .Z(n3015) );
  AND U3133 ( .A(b[7]), .B(a[68]), .Z(n3014) );
  XNOR U3134 ( .A(n3015), .B(n3014), .Z(n3016) );
  XNOR U3135 ( .A(n3017), .B(n3016), .Z(n3022) );
  XOR U3136 ( .A(n3023), .B(n3022), .Z(n2997) );
  NANDN U3137 ( .A(n2974), .B(n2973), .Z(n2978) );
  NANDN U3138 ( .A(n2976), .B(n2975), .Z(n2977) );
  AND U3139 ( .A(n2978), .B(n2977), .Z(n2996) );
  XNOR U3140 ( .A(n2997), .B(n2996), .Z(n2998) );
  NANDN U3141 ( .A(n2980), .B(n2979), .Z(n2984) );
  NAND U3142 ( .A(n2982), .B(n2981), .Z(n2983) );
  NAND U3143 ( .A(n2984), .B(n2983), .Z(n2999) );
  XNOR U3144 ( .A(n2998), .B(n2999), .Z(n2990) );
  XNOR U3145 ( .A(n2991), .B(n2990), .Z(n2992) );
  XNOR U3146 ( .A(n2993), .B(n2992), .Z(n3026) );
  XNOR U3147 ( .A(sreg[196]), .B(n3026), .Z(n3028) );
  NANDN U3148 ( .A(sreg[195]), .B(n2985), .Z(n2989) );
  NAND U3149 ( .A(n2987), .B(n2986), .Z(n2988) );
  NAND U3150 ( .A(n2989), .B(n2988), .Z(n3027) );
  XNOR U3151 ( .A(n3028), .B(n3027), .Z(c[196]) );
  NANDN U3152 ( .A(n2991), .B(n2990), .Z(n2995) );
  NANDN U3153 ( .A(n2993), .B(n2992), .Z(n2994) );
  AND U3154 ( .A(n2995), .B(n2994), .Z(n3034) );
  NANDN U3155 ( .A(n2997), .B(n2996), .Z(n3001) );
  NANDN U3156 ( .A(n2999), .B(n2998), .Z(n3000) );
  AND U3157 ( .A(n3001), .B(n3000), .Z(n3032) );
  NANDN U3158 ( .A(n5274), .B(n3002), .Z(n3004) );
  XOR U3159 ( .A(b[7]), .B(a[71]), .Z(n3043) );
  NANDN U3160 ( .A(n5275), .B(n3043), .Z(n3003) );
  AND U3161 ( .A(n3004), .B(n3003), .Z(n3062) );
  NANDN U3162 ( .A(n5176), .B(n3005), .Z(n3007) );
  XOR U3163 ( .A(b[3]), .B(a[75]), .Z(n3046) );
  NANDN U3164 ( .A(n5177), .B(n3046), .Z(n3006) );
  NAND U3165 ( .A(n3007), .B(n3006), .Z(n3061) );
  XNOR U3166 ( .A(n3062), .B(n3061), .Z(n3064) );
  NAND U3167 ( .A(b[0]), .B(a[77]), .Z(n3008) );
  XNOR U3168 ( .A(b[1]), .B(n3008), .Z(n3010) );
  NANDN U3169 ( .A(b[0]), .B(a[76]), .Z(n3009) );
  NAND U3170 ( .A(n3010), .B(n3009), .Z(n3058) );
  NANDN U3171 ( .A(n5249), .B(n3011), .Z(n3013) );
  XOR U3172 ( .A(b[5]), .B(a[73]), .Z(n3049) );
  NANDN U3173 ( .A(n5184), .B(n3049), .Z(n3012) );
  AND U3174 ( .A(n3013), .B(n3012), .Z(n3056) );
  AND U3175 ( .A(b[7]), .B(a[69]), .Z(n3055) );
  XNOR U3176 ( .A(n3056), .B(n3055), .Z(n3057) );
  XNOR U3177 ( .A(n3058), .B(n3057), .Z(n3063) );
  XOR U3178 ( .A(n3064), .B(n3063), .Z(n3038) );
  NANDN U3179 ( .A(n3015), .B(n3014), .Z(n3019) );
  NANDN U3180 ( .A(n3017), .B(n3016), .Z(n3018) );
  AND U3181 ( .A(n3019), .B(n3018), .Z(n3037) );
  XNOR U3182 ( .A(n3038), .B(n3037), .Z(n3039) );
  NANDN U3183 ( .A(n3021), .B(n3020), .Z(n3025) );
  NAND U3184 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U3185 ( .A(n3025), .B(n3024), .Z(n3040) );
  XNOR U3186 ( .A(n3039), .B(n3040), .Z(n3031) );
  XNOR U3187 ( .A(n3032), .B(n3031), .Z(n3033) );
  XNOR U3188 ( .A(n3034), .B(n3033), .Z(n3067) );
  XNOR U3189 ( .A(sreg[197]), .B(n3067), .Z(n3069) );
  NANDN U3190 ( .A(sreg[196]), .B(n3026), .Z(n3030) );
  NAND U3191 ( .A(n3028), .B(n3027), .Z(n3029) );
  NAND U3192 ( .A(n3030), .B(n3029), .Z(n3068) );
  XNOR U3193 ( .A(n3069), .B(n3068), .Z(c[197]) );
  NANDN U3194 ( .A(n3032), .B(n3031), .Z(n3036) );
  NANDN U3195 ( .A(n3034), .B(n3033), .Z(n3035) );
  AND U3196 ( .A(n3036), .B(n3035), .Z(n3075) );
  NANDN U3197 ( .A(n3038), .B(n3037), .Z(n3042) );
  NANDN U3198 ( .A(n3040), .B(n3039), .Z(n3041) );
  AND U3199 ( .A(n3042), .B(n3041), .Z(n3073) );
  NANDN U3200 ( .A(n5274), .B(n3043), .Z(n3045) );
  XOR U3201 ( .A(b[7]), .B(a[72]), .Z(n3084) );
  NANDN U3202 ( .A(n5275), .B(n3084), .Z(n3044) );
  AND U3203 ( .A(n3045), .B(n3044), .Z(n3103) );
  NANDN U3204 ( .A(n5176), .B(n3046), .Z(n3048) );
  XOR U3205 ( .A(b[3]), .B(a[76]), .Z(n3087) );
  NANDN U3206 ( .A(n5177), .B(n3087), .Z(n3047) );
  NAND U3207 ( .A(n3048), .B(n3047), .Z(n3102) );
  XNOR U3208 ( .A(n3103), .B(n3102), .Z(n3105) );
  NANDN U3209 ( .A(n5249), .B(n3049), .Z(n3051) );
  XOR U3210 ( .A(b[5]), .B(a[74]), .Z(n3093) );
  NANDN U3211 ( .A(n5184), .B(n3093), .Z(n3050) );
  AND U3212 ( .A(n3051), .B(n3050), .Z(n3097) );
  AND U3213 ( .A(b[7]), .B(a[70]), .Z(n3096) );
  XNOR U3214 ( .A(n3097), .B(n3096), .Z(n3098) );
  NAND U3215 ( .A(b[0]), .B(a[78]), .Z(n3052) );
  XNOR U3216 ( .A(b[1]), .B(n3052), .Z(n3054) );
  NANDN U3217 ( .A(b[0]), .B(a[77]), .Z(n3053) );
  NAND U3218 ( .A(n3054), .B(n3053), .Z(n3099) );
  XNOR U3219 ( .A(n3098), .B(n3099), .Z(n3104) );
  XOR U3220 ( .A(n3105), .B(n3104), .Z(n3079) );
  NANDN U3221 ( .A(n3056), .B(n3055), .Z(n3060) );
  NANDN U3222 ( .A(n3058), .B(n3057), .Z(n3059) );
  AND U3223 ( .A(n3060), .B(n3059), .Z(n3078) );
  XNOR U3224 ( .A(n3079), .B(n3078), .Z(n3080) );
  NANDN U3225 ( .A(n3062), .B(n3061), .Z(n3066) );
  NAND U3226 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U3227 ( .A(n3066), .B(n3065), .Z(n3081) );
  XNOR U3228 ( .A(n3080), .B(n3081), .Z(n3072) );
  XNOR U3229 ( .A(n3073), .B(n3072), .Z(n3074) );
  XNOR U3230 ( .A(n3075), .B(n3074), .Z(n3108) );
  XNOR U3231 ( .A(sreg[198]), .B(n3108), .Z(n3110) );
  NANDN U3232 ( .A(sreg[197]), .B(n3067), .Z(n3071) );
  NAND U3233 ( .A(n3069), .B(n3068), .Z(n3070) );
  NAND U3234 ( .A(n3071), .B(n3070), .Z(n3109) );
  XNOR U3235 ( .A(n3110), .B(n3109), .Z(c[198]) );
  NANDN U3236 ( .A(n3073), .B(n3072), .Z(n3077) );
  NANDN U3237 ( .A(n3075), .B(n3074), .Z(n3076) );
  AND U3238 ( .A(n3077), .B(n3076), .Z(n3116) );
  NANDN U3239 ( .A(n3079), .B(n3078), .Z(n3083) );
  NANDN U3240 ( .A(n3081), .B(n3080), .Z(n3082) );
  AND U3241 ( .A(n3083), .B(n3082), .Z(n3114) );
  NANDN U3242 ( .A(n5274), .B(n3084), .Z(n3086) );
  XOR U3243 ( .A(b[7]), .B(a[73]), .Z(n3125) );
  NANDN U3244 ( .A(n5275), .B(n3125), .Z(n3085) );
  AND U3245 ( .A(n3086), .B(n3085), .Z(n3144) );
  NANDN U3246 ( .A(n5176), .B(n3087), .Z(n3089) );
  XOR U3247 ( .A(b[3]), .B(a[77]), .Z(n3128) );
  NANDN U3248 ( .A(n5177), .B(n3128), .Z(n3088) );
  NAND U3249 ( .A(n3089), .B(n3088), .Z(n3143) );
  XNOR U3250 ( .A(n3144), .B(n3143), .Z(n3146) );
  NAND U3251 ( .A(b[0]), .B(a[79]), .Z(n3090) );
  XNOR U3252 ( .A(b[1]), .B(n3090), .Z(n3092) );
  NANDN U3253 ( .A(b[0]), .B(a[78]), .Z(n3091) );
  NAND U3254 ( .A(n3092), .B(n3091), .Z(n3140) );
  NANDN U3255 ( .A(n5249), .B(n3093), .Z(n3095) );
  XOR U3256 ( .A(b[5]), .B(a[75]), .Z(n3134) );
  NANDN U3257 ( .A(n5184), .B(n3134), .Z(n3094) );
  AND U3258 ( .A(n3095), .B(n3094), .Z(n3138) );
  AND U3259 ( .A(b[7]), .B(a[71]), .Z(n3137) );
  XNOR U3260 ( .A(n3138), .B(n3137), .Z(n3139) );
  XNOR U3261 ( .A(n3140), .B(n3139), .Z(n3145) );
  XOR U3262 ( .A(n3146), .B(n3145), .Z(n3120) );
  NANDN U3263 ( .A(n3097), .B(n3096), .Z(n3101) );
  NANDN U3264 ( .A(n3099), .B(n3098), .Z(n3100) );
  AND U3265 ( .A(n3101), .B(n3100), .Z(n3119) );
  XNOR U3266 ( .A(n3120), .B(n3119), .Z(n3121) );
  NANDN U3267 ( .A(n3103), .B(n3102), .Z(n3107) );
  NAND U3268 ( .A(n3105), .B(n3104), .Z(n3106) );
  NAND U3269 ( .A(n3107), .B(n3106), .Z(n3122) );
  XNOR U3270 ( .A(n3121), .B(n3122), .Z(n3113) );
  XNOR U3271 ( .A(n3114), .B(n3113), .Z(n3115) );
  XNOR U3272 ( .A(n3116), .B(n3115), .Z(n3149) );
  XNOR U3273 ( .A(sreg[199]), .B(n3149), .Z(n3151) );
  NANDN U3274 ( .A(sreg[198]), .B(n3108), .Z(n3112) );
  NAND U3275 ( .A(n3110), .B(n3109), .Z(n3111) );
  NAND U3276 ( .A(n3112), .B(n3111), .Z(n3150) );
  XNOR U3277 ( .A(n3151), .B(n3150), .Z(c[199]) );
  NANDN U3278 ( .A(n3114), .B(n3113), .Z(n3118) );
  NANDN U3279 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U3280 ( .A(n3118), .B(n3117), .Z(n3157) );
  NANDN U3281 ( .A(n3120), .B(n3119), .Z(n3124) );
  NANDN U3282 ( .A(n3122), .B(n3121), .Z(n3123) );
  AND U3283 ( .A(n3124), .B(n3123), .Z(n3155) );
  NANDN U3284 ( .A(n5274), .B(n3125), .Z(n3127) );
  XOR U3285 ( .A(b[7]), .B(a[74]), .Z(n3166) );
  NANDN U3286 ( .A(n5275), .B(n3166), .Z(n3126) );
  AND U3287 ( .A(n3127), .B(n3126), .Z(n3185) );
  NANDN U3288 ( .A(n5176), .B(n3128), .Z(n3130) );
  XOR U3289 ( .A(b[3]), .B(a[78]), .Z(n3169) );
  NANDN U3290 ( .A(n5177), .B(n3169), .Z(n3129) );
  NAND U3291 ( .A(n3130), .B(n3129), .Z(n3184) );
  XNOR U3292 ( .A(n3185), .B(n3184), .Z(n3187) );
  NAND U3293 ( .A(b[0]), .B(a[80]), .Z(n3131) );
  XNOR U3294 ( .A(b[1]), .B(n3131), .Z(n3133) );
  NANDN U3295 ( .A(b[0]), .B(a[79]), .Z(n3132) );
  NAND U3296 ( .A(n3133), .B(n3132), .Z(n3181) );
  NANDN U3297 ( .A(n5249), .B(n3134), .Z(n3136) );
  XOR U3298 ( .A(b[5]), .B(a[76]), .Z(n3175) );
  NANDN U3299 ( .A(n5184), .B(n3175), .Z(n3135) );
  AND U3300 ( .A(n3136), .B(n3135), .Z(n3179) );
  AND U3301 ( .A(b[7]), .B(a[72]), .Z(n3178) );
  XNOR U3302 ( .A(n3179), .B(n3178), .Z(n3180) );
  XNOR U3303 ( .A(n3181), .B(n3180), .Z(n3186) );
  XOR U3304 ( .A(n3187), .B(n3186), .Z(n3161) );
  NANDN U3305 ( .A(n3138), .B(n3137), .Z(n3142) );
  NANDN U3306 ( .A(n3140), .B(n3139), .Z(n3141) );
  AND U3307 ( .A(n3142), .B(n3141), .Z(n3160) );
  XNOR U3308 ( .A(n3161), .B(n3160), .Z(n3162) );
  NANDN U3309 ( .A(n3144), .B(n3143), .Z(n3148) );
  NAND U3310 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3311 ( .A(n3148), .B(n3147), .Z(n3163) );
  XNOR U3312 ( .A(n3162), .B(n3163), .Z(n3154) );
  XNOR U3313 ( .A(n3155), .B(n3154), .Z(n3156) );
  XNOR U3314 ( .A(n3157), .B(n3156), .Z(n3190) );
  XNOR U3315 ( .A(sreg[200]), .B(n3190), .Z(n3192) );
  NANDN U3316 ( .A(sreg[199]), .B(n3149), .Z(n3153) );
  NAND U3317 ( .A(n3151), .B(n3150), .Z(n3152) );
  NAND U3318 ( .A(n3153), .B(n3152), .Z(n3191) );
  XNOR U3319 ( .A(n3192), .B(n3191), .Z(c[200]) );
  NANDN U3320 ( .A(n3155), .B(n3154), .Z(n3159) );
  NANDN U3321 ( .A(n3157), .B(n3156), .Z(n3158) );
  AND U3322 ( .A(n3159), .B(n3158), .Z(n3198) );
  NANDN U3323 ( .A(n3161), .B(n3160), .Z(n3165) );
  NANDN U3324 ( .A(n3163), .B(n3162), .Z(n3164) );
  AND U3325 ( .A(n3165), .B(n3164), .Z(n3196) );
  NANDN U3326 ( .A(n5274), .B(n3166), .Z(n3168) );
  XOR U3327 ( .A(b[7]), .B(a[75]), .Z(n3207) );
  NANDN U3328 ( .A(n5275), .B(n3207), .Z(n3167) );
  AND U3329 ( .A(n3168), .B(n3167), .Z(n3226) );
  NANDN U3330 ( .A(n5176), .B(n3169), .Z(n3171) );
  XOR U3331 ( .A(b[3]), .B(a[79]), .Z(n3210) );
  NANDN U3332 ( .A(n5177), .B(n3210), .Z(n3170) );
  NAND U3333 ( .A(n3171), .B(n3170), .Z(n3225) );
  XNOR U3334 ( .A(n3226), .B(n3225), .Z(n3228) );
  NAND U3335 ( .A(b[0]), .B(a[81]), .Z(n3172) );
  XNOR U3336 ( .A(b[1]), .B(n3172), .Z(n3174) );
  NANDN U3337 ( .A(b[0]), .B(a[80]), .Z(n3173) );
  NAND U3338 ( .A(n3174), .B(n3173), .Z(n3222) );
  NANDN U3339 ( .A(n5249), .B(n3175), .Z(n3177) );
  XOR U3340 ( .A(b[5]), .B(a[77]), .Z(n3216) );
  NANDN U3341 ( .A(n5184), .B(n3216), .Z(n3176) );
  AND U3342 ( .A(n3177), .B(n3176), .Z(n3220) );
  AND U3343 ( .A(b[7]), .B(a[73]), .Z(n3219) );
  XNOR U3344 ( .A(n3220), .B(n3219), .Z(n3221) );
  XNOR U3345 ( .A(n3222), .B(n3221), .Z(n3227) );
  XOR U3346 ( .A(n3228), .B(n3227), .Z(n3202) );
  NANDN U3347 ( .A(n3179), .B(n3178), .Z(n3183) );
  NANDN U3348 ( .A(n3181), .B(n3180), .Z(n3182) );
  AND U3349 ( .A(n3183), .B(n3182), .Z(n3201) );
  XNOR U3350 ( .A(n3202), .B(n3201), .Z(n3203) );
  NANDN U3351 ( .A(n3185), .B(n3184), .Z(n3189) );
  NAND U3352 ( .A(n3187), .B(n3186), .Z(n3188) );
  NAND U3353 ( .A(n3189), .B(n3188), .Z(n3204) );
  XNOR U3354 ( .A(n3203), .B(n3204), .Z(n3195) );
  XNOR U3355 ( .A(n3196), .B(n3195), .Z(n3197) );
  XNOR U3356 ( .A(n3198), .B(n3197), .Z(n3231) );
  XNOR U3357 ( .A(sreg[201]), .B(n3231), .Z(n3233) );
  NANDN U3358 ( .A(sreg[200]), .B(n3190), .Z(n3194) );
  NAND U3359 ( .A(n3192), .B(n3191), .Z(n3193) );
  NAND U3360 ( .A(n3194), .B(n3193), .Z(n3232) );
  XNOR U3361 ( .A(n3233), .B(n3232), .Z(c[201]) );
  NANDN U3362 ( .A(n3196), .B(n3195), .Z(n3200) );
  NANDN U3363 ( .A(n3198), .B(n3197), .Z(n3199) );
  AND U3364 ( .A(n3200), .B(n3199), .Z(n3239) );
  NANDN U3365 ( .A(n3202), .B(n3201), .Z(n3206) );
  NANDN U3366 ( .A(n3204), .B(n3203), .Z(n3205) );
  AND U3367 ( .A(n3206), .B(n3205), .Z(n3237) );
  NANDN U3368 ( .A(n5274), .B(n3207), .Z(n3209) );
  XOR U3369 ( .A(b[7]), .B(a[76]), .Z(n3248) );
  NANDN U3370 ( .A(n5275), .B(n3248), .Z(n3208) );
  AND U3371 ( .A(n3209), .B(n3208), .Z(n3267) );
  NANDN U3372 ( .A(n5176), .B(n3210), .Z(n3212) );
  XOR U3373 ( .A(b[3]), .B(a[80]), .Z(n3251) );
  NANDN U3374 ( .A(n5177), .B(n3251), .Z(n3211) );
  NAND U3375 ( .A(n3212), .B(n3211), .Z(n3266) );
  XNOR U3376 ( .A(n3267), .B(n3266), .Z(n3269) );
  NAND U3377 ( .A(b[0]), .B(a[82]), .Z(n3213) );
  XNOR U3378 ( .A(b[1]), .B(n3213), .Z(n3215) );
  NANDN U3379 ( .A(b[0]), .B(a[81]), .Z(n3214) );
  NAND U3380 ( .A(n3215), .B(n3214), .Z(n3263) );
  NANDN U3381 ( .A(n5249), .B(n3216), .Z(n3218) );
  XOR U3382 ( .A(b[5]), .B(a[78]), .Z(n3257) );
  NANDN U3383 ( .A(n5184), .B(n3257), .Z(n3217) );
  AND U3384 ( .A(n3218), .B(n3217), .Z(n3261) );
  AND U3385 ( .A(b[7]), .B(a[74]), .Z(n3260) );
  XNOR U3386 ( .A(n3261), .B(n3260), .Z(n3262) );
  XNOR U3387 ( .A(n3263), .B(n3262), .Z(n3268) );
  XOR U3388 ( .A(n3269), .B(n3268), .Z(n3243) );
  NANDN U3389 ( .A(n3220), .B(n3219), .Z(n3224) );
  NANDN U3390 ( .A(n3222), .B(n3221), .Z(n3223) );
  AND U3391 ( .A(n3224), .B(n3223), .Z(n3242) );
  XNOR U3392 ( .A(n3243), .B(n3242), .Z(n3244) );
  NANDN U3393 ( .A(n3226), .B(n3225), .Z(n3230) );
  NAND U3394 ( .A(n3228), .B(n3227), .Z(n3229) );
  NAND U3395 ( .A(n3230), .B(n3229), .Z(n3245) );
  XNOR U3396 ( .A(n3244), .B(n3245), .Z(n3236) );
  XNOR U3397 ( .A(n3237), .B(n3236), .Z(n3238) );
  XNOR U3398 ( .A(n3239), .B(n3238), .Z(n3272) );
  XNOR U3399 ( .A(sreg[202]), .B(n3272), .Z(n3274) );
  NANDN U3400 ( .A(sreg[201]), .B(n3231), .Z(n3235) );
  NAND U3401 ( .A(n3233), .B(n3232), .Z(n3234) );
  NAND U3402 ( .A(n3235), .B(n3234), .Z(n3273) );
  XNOR U3403 ( .A(n3274), .B(n3273), .Z(c[202]) );
  NANDN U3404 ( .A(n3237), .B(n3236), .Z(n3241) );
  NANDN U3405 ( .A(n3239), .B(n3238), .Z(n3240) );
  AND U3406 ( .A(n3241), .B(n3240), .Z(n3280) );
  NANDN U3407 ( .A(n3243), .B(n3242), .Z(n3247) );
  NANDN U3408 ( .A(n3245), .B(n3244), .Z(n3246) );
  AND U3409 ( .A(n3247), .B(n3246), .Z(n3278) );
  NANDN U3410 ( .A(n5274), .B(n3248), .Z(n3250) );
  XOR U3411 ( .A(b[7]), .B(a[77]), .Z(n3289) );
  NANDN U3412 ( .A(n5275), .B(n3289), .Z(n3249) );
  AND U3413 ( .A(n3250), .B(n3249), .Z(n3308) );
  NANDN U3414 ( .A(n5176), .B(n3251), .Z(n3253) );
  XOR U3415 ( .A(b[3]), .B(a[81]), .Z(n3292) );
  NANDN U3416 ( .A(n5177), .B(n3292), .Z(n3252) );
  NAND U3417 ( .A(n3253), .B(n3252), .Z(n3307) );
  XNOR U3418 ( .A(n3308), .B(n3307), .Z(n3310) );
  NAND U3419 ( .A(b[0]), .B(a[83]), .Z(n3254) );
  XNOR U3420 ( .A(b[1]), .B(n3254), .Z(n3256) );
  NANDN U3421 ( .A(b[0]), .B(a[82]), .Z(n3255) );
  NAND U3422 ( .A(n3256), .B(n3255), .Z(n3304) );
  NANDN U3423 ( .A(n5249), .B(n3257), .Z(n3259) );
  XOR U3424 ( .A(b[5]), .B(a[79]), .Z(n3298) );
  NANDN U3425 ( .A(n5184), .B(n3298), .Z(n3258) );
  AND U3426 ( .A(n3259), .B(n3258), .Z(n3302) );
  AND U3427 ( .A(b[7]), .B(a[75]), .Z(n3301) );
  XNOR U3428 ( .A(n3302), .B(n3301), .Z(n3303) );
  XNOR U3429 ( .A(n3304), .B(n3303), .Z(n3309) );
  XOR U3430 ( .A(n3310), .B(n3309), .Z(n3284) );
  NANDN U3431 ( .A(n3261), .B(n3260), .Z(n3265) );
  NANDN U3432 ( .A(n3263), .B(n3262), .Z(n3264) );
  AND U3433 ( .A(n3265), .B(n3264), .Z(n3283) );
  XNOR U3434 ( .A(n3284), .B(n3283), .Z(n3285) );
  NANDN U3435 ( .A(n3267), .B(n3266), .Z(n3271) );
  NAND U3436 ( .A(n3269), .B(n3268), .Z(n3270) );
  NAND U3437 ( .A(n3271), .B(n3270), .Z(n3286) );
  XNOR U3438 ( .A(n3285), .B(n3286), .Z(n3277) );
  XNOR U3439 ( .A(n3278), .B(n3277), .Z(n3279) );
  XNOR U3440 ( .A(n3280), .B(n3279), .Z(n3313) );
  XNOR U3441 ( .A(sreg[203]), .B(n3313), .Z(n3315) );
  NANDN U3442 ( .A(sreg[202]), .B(n3272), .Z(n3276) );
  NAND U3443 ( .A(n3274), .B(n3273), .Z(n3275) );
  NAND U3444 ( .A(n3276), .B(n3275), .Z(n3314) );
  XNOR U3445 ( .A(n3315), .B(n3314), .Z(c[203]) );
  NANDN U3446 ( .A(n3278), .B(n3277), .Z(n3282) );
  NANDN U3447 ( .A(n3280), .B(n3279), .Z(n3281) );
  AND U3448 ( .A(n3282), .B(n3281), .Z(n3321) );
  NANDN U3449 ( .A(n3284), .B(n3283), .Z(n3288) );
  NANDN U3450 ( .A(n3286), .B(n3285), .Z(n3287) );
  AND U3451 ( .A(n3288), .B(n3287), .Z(n3319) );
  NANDN U3452 ( .A(n5274), .B(n3289), .Z(n3291) );
  XOR U3453 ( .A(b[7]), .B(a[78]), .Z(n3330) );
  NANDN U3454 ( .A(n5275), .B(n3330), .Z(n3290) );
  AND U3455 ( .A(n3291), .B(n3290), .Z(n3349) );
  NANDN U3456 ( .A(n5176), .B(n3292), .Z(n3294) );
  XOR U3457 ( .A(b[3]), .B(a[82]), .Z(n3333) );
  NANDN U3458 ( .A(n5177), .B(n3333), .Z(n3293) );
  NAND U3459 ( .A(n3294), .B(n3293), .Z(n3348) );
  XNOR U3460 ( .A(n3349), .B(n3348), .Z(n3351) );
  NAND U3461 ( .A(b[0]), .B(a[84]), .Z(n3295) );
  XNOR U3462 ( .A(b[1]), .B(n3295), .Z(n3297) );
  NANDN U3463 ( .A(b[0]), .B(a[83]), .Z(n3296) );
  NAND U3464 ( .A(n3297), .B(n3296), .Z(n3345) );
  NANDN U3465 ( .A(n5249), .B(n3298), .Z(n3300) );
  XOR U3466 ( .A(b[5]), .B(a[80]), .Z(n3336) );
  NANDN U3467 ( .A(n5184), .B(n3336), .Z(n3299) );
  AND U3468 ( .A(n3300), .B(n3299), .Z(n3343) );
  AND U3469 ( .A(b[7]), .B(a[76]), .Z(n3342) );
  XNOR U3470 ( .A(n3343), .B(n3342), .Z(n3344) );
  XNOR U3471 ( .A(n3345), .B(n3344), .Z(n3350) );
  XOR U3472 ( .A(n3351), .B(n3350), .Z(n3325) );
  NANDN U3473 ( .A(n3302), .B(n3301), .Z(n3306) );
  NANDN U3474 ( .A(n3304), .B(n3303), .Z(n3305) );
  AND U3475 ( .A(n3306), .B(n3305), .Z(n3324) );
  XNOR U3476 ( .A(n3325), .B(n3324), .Z(n3326) );
  NANDN U3477 ( .A(n3308), .B(n3307), .Z(n3312) );
  NAND U3478 ( .A(n3310), .B(n3309), .Z(n3311) );
  NAND U3479 ( .A(n3312), .B(n3311), .Z(n3327) );
  XNOR U3480 ( .A(n3326), .B(n3327), .Z(n3318) );
  XNOR U3481 ( .A(n3319), .B(n3318), .Z(n3320) );
  XNOR U3482 ( .A(n3321), .B(n3320), .Z(n3354) );
  XNOR U3483 ( .A(sreg[204]), .B(n3354), .Z(n3356) );
  NANDN U3484 ( .A(sreg[203]), .B(n3313), .Z(n3317) );
  NAND U3485 ( .A(n3315), .B(n3314), .Z(n3316) );
  NAND U3486 ( .A(n3317), .B(n3316), .Z(n3355) );
  XNOR U3487 ( .A(n3356), .B(n3355), .Z(c[204]) );
  NANDN U3488 ( .A(n3319), .B(n3318), .Z(n3323) );
  NANDN U3489 ( .A(n3321), .B(n3320), .Z(n3322) );
  AND U3490 ( .A(n3323), .B(n3322), .Z(n3362) );
  NANDN U3491 ( .A(n3325), .B(n3324), .Z(n3329) );
  NANDN U3492 ( .A(n3327), .B(n3326), .Z(n3328) );
  AND U3493 ( .A(n3329), .B(n3328), .Z(n3360) );
  NANDN U3494 ( .A(n5274), .B(n3330), .Z(n3332) );
  XOR U3495 ( .A(b[7]), .B(a[79]), .Z(n3371) );
  NANDN U3496 ( .A(n5275), .B(n3371), .Z(n3331) );
  AND U3497 ( .A(n3332), .B(n3331), .Z(n3390) );
  NANDN U3498 ( .A(n5176), .B(n3333), .Z(n3335) );
  XOR U3499 ( .A(b[3]), .B(a[83]), .Z(n3374) );
  NANDN U3500 ( .A(n5177), .B(n3374), .Z(n3334) );
  NAND U3501 ( .A(n3335), .B(n3334), .Z(n3389) );
  XNOR U3502 ( .A(n3390), .B(n3389), .Z(n3392) );
  NANDN U3503 ( .A(n5249), .B(n3336), .Z(n3338) );
  XOR U3504 ( .A(b[5]), .B(a[81]), .Z(n3380) );
  NANDN U3505 ( .A(n5184), .B(n3380), .Z(n3337) );
  AND U3506 ( .A(n3338), .B(n3337), .Z(n3384) );
  AND U3507 ( .A(b[7]), .B(a[77]), .Z(n3383) );
  XNOR U3508 ( .A(n3384), .B(n3383), .Z(n3385) );
  NAND U3509 ( .A(b[0]), .B(a[85]), .Z(n3339) );
  XNOR U3510 ( .A(b[1]), .B(n3339), .Z(n3341) );
  NANDN U3511 ( .A(b[0]), .B(a[84]), .Z(n3340) );
  NAND U3512 ( .A(n3341), .B(n3340), .Z(n3386) );
  XNOR U3513 ( .A(n3385), .B(n3386), .Z(n3391) );
  XOR U3514 ( .A(n3392), .B(n3391), .Z(n3366) );
  NANDN U3515 ( .A(n3343), .B(n3342), .Z(n3347) );
  NANDN U3516 ( .A(n3345), .B(n3344), .Z(n3346) );
  AND U3517 ( .A(n3347), .B(n3346), .Z(n3365) );
  XNOR U3518 ( .A(n3366), .B(n3365), .Z(n3367) );
  NANDN U3519 ( .A(n3349), .B(n3348), .Z(n3353) );
  NAND U3520 ( .A(n3351), .B(n3350), .Z(n3352) );
  NAND U3521 ( .A(n3353), .B(n3352), .Z(n3368) );
  XNOR U3522 ( .A(n3367), .B(n3368), .Z(n3359) );
  XNOR U3523 ( .A(n3360), .B(n3359), .Z(n3361) );
  XNOR U3524 ( .A(n3362), .B(n3361), .Z(n3395) );
  XNOR U3525 ( .A(sreg[205]), .B(n3395), .Z(n3397) );
  NANDN U3526 ( .A(sreg[204]), .B(n3354), .Z(n3358) );
  NAND U3527 ( .A(n3356), .B(n3355), .Z(n3357) );
  NAND U3528 ( .A(n3358), .B(n3357), .Z(n3396) );
  XNOR U3529 ( .A(n3397), .B(n3396), .Z(c[205]) );
  NANDN U3530 ( .A(n3360), .B(n3359), .Z(n3364) );
  NANDN U3531 ( .A(n3362), .B(n3361), .Z(n3363) );
  AND U3532 ( .A(n3364), .B(n3363), .Z(n3403) );
  NANDN U3533 ( .A(n3366), .B(n3365), .Z(n3370) );
  NANDN U3534 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3535 ( .A(n3370), .B(n3369), .Z(n3401) );
  NANDN U3536 ( .A(n5274), .B(n3371), .Z(n3373) );
  XOR U3537 ( .A(b[7]), .B(a[80]), .Z(n3412) );
  NANDN U3538 ( .A(n5275), .B(n3412), .Z(n3372) );
  AND U3539 ( .A(n3373), .B(n3372), .Z(n3431) );
  NANDN U3540 ( .A(n5176), .B(n3374), .Z(n3376) );
  XOR U3541 ( .A(b[3]), .B(a[84]), .Z(n3415) );
  NANDN U3542 ( .A(n5177), .B(n3415), .Z(n3375) );
  NAND U3543 ( .A(n3376), .B(n3375), .Z(n3430) );
  XNOR U3544 ( .A(n3431), .B(n3430), .Z(n3433) );
  NAND U3545 ( .A(b[0]), .B(a[86]), .Z(n3377) );
  XNOR U3546 ( .A(b[1]), .B(n3377), .Z(n3379) );
  NANDN U3547 ( .A(b[0]), .B(a[85]), .Z(n3378) );
  NAND U3548 ( .A(n3379), .B(n3378), .Z(n3427) );
  NANDN U3549 ( .A(n5249), .B(n3380), .Z(n3382) );
  XOR U3550 ( .A(b[5]), .B(a[82]), .Z(n3418) );
  NANDN U3551 ( .A(n5184), .B(n3418), .Z(n3381) );
  AND U3552 ( .A(n3382), .B(n3381), .Z(n3425) );
  AND U3553 ( .A(b[7]), .B(a[78]), .Z(n3424) );
  XNOR U3554 ( .A(n3425), .B(n3424), .Z(n3426) );
  XNOR U3555 ( .A(n3427), .B(n3426), .Z(n3432) );
  XOR U3556 ( .A(n3433), .B(n3432), .Z(n3407) );
  NANDN U3557 ( .A(n3384), .B(n3383), .Z(n3388) );
  NANDN U3558 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U3559 ( .A(n3388), .B(n3387), .Z(n3406) );
  XNOR U3560 ( .A(n3407), .B(n3406), .Z(n3408) );
  NANDN U3561 ( .A(n3390), .B(n3389), .Z(n3394) );
  NAND U3562 ( .A(n3392), .B(n3391), .Z(n3393) );
  NAND U3563 ( .A(n3394), .B(n3393), .Z(n3409) );
  XNOR U3564 ( .A(n3408), .B(n3409), .Z(n3400) );
  XNOR U3565 ( .A(n3401), .B(n3400), .Z(n3402) );
  XNOR U3566 ( .A(n3403), .B(n3402), .Z(n3436) );
  XNOR U3567 ( .A(sreg[206]), .B(n3436), .Z(n3438) );
  NANDN U3568 ( .A(sreg[205]), .B(n3395), .Z(n3399) );
  NAND U3569 ( .A(n3397), .B(n3396), .Z(n3398) );
  NAND U3570 ( .A(n3399), .B(n3398), .Z(n3437) );
  XNOR U3571 ( .A(n3438), .B(n3437), .Z(c[206]) );
  NANDN U3572 ( .A(n3401), .B(n3400), .Z(n3405) );
  NANDN U3573 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U3574 ( .A(n3405), .B(n3404), .Z(n3444) );
  NANDN U3575 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U3576 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U3577 ( .A(n3411), .B(n3410), .Z(n3442) );
  NANDN U3578 ( .A(n5274), .B(n3412), .Z(n3414) );
  XOR U3579 ( .A(b[7]), .B(a[81]), .Z(n3453) );
  NANDN U3580 ( .A(n5275), .B(n3453), .Z(n3413) );
  AND U3581 ( .A(n3414), .B(n3413), .Z(n3472) );
  NANDN U3582 ( .A(n5176), .B(n3415), .Z(n3417) );
  XOR U3583 ( .A(b[3]), .B(a[85]), .Z(n3456) );
  NANDN U3584 ( .A(n5177), .B(n3456), .Z(n3416) );
  NAND U3585 ( .A(n3417), .B(n3416), .Z(n3471) );
  XNOR U3586 ( .A(n3472), .B(n3471), .Z(n3474) );
  NANDN U3587 ( .A(n5249), .B(n3418), .Z(n3420) );
  XOR U3588 ( .A(b[5]), .B(a[83]), .Z(n3459) );
  NANDN U3589 ( .A(n5184), .B(n3459), .Z(n3419) );
  AND U3590 ( .A(n3420), .B(n3419), .Z(n3466) );
  AND U3591 ( .A(b[7]), .B(a[79]), .Z(n3465) );
  XNOR U3592 ( .A(n3466), .B(n3465), .Z(n3467) );
  NAND U3593 ( .A(b[0]), .B(a[87]), .Z(n3421) );
  XNOR U3594 ( .A(b[1]), .B(n3421), .Z(n3423) );
  NANDN U3595 ( .A(b[0]), .B(a[86]), .Z(n3422) );
  NAND U3596 ( .A(n3423), .B(n3422), .Z(n3468) );
  XNOR U3597 ( .A(n3467), .B(n3468), .Z(n3473) );
  XOR U3598 ( .A(n3474), .B(n3473), .Z(n3448) );
  NANDN U3599 ( .A(n3425), .B(n3424), .Z(n3429) );
  NANDN U3600 ( .A(n3427), .B(n3426), .Z(n3428) );
  AND U3601 ( .A(n3429), .B(n3428), .Z(n3447) );
  XNOR U3602 ( .A(n3448), .B(n3447), .Z(n3449) );
  NANDN U3603 ( .A(n3431), .B(n3430), .Z(n3435) );
  NAND U3604 ( .A(n3433), .B(n3432), .Z(n3434) );
  NAND U3605 ( .A(n3435), .B(n3434), .Z(n3450) );
  XNOR U3606 ( .A(n3449), .B(n3450), .Z(n3441) );
  XNOR U3607 ( .A(n3442), .B(n3441), .Z(n3443) );
  XNOR U3608 ( .A(n3444), .B(n3443), .Z(n3477) );
  XNOR U3609 ( .A(sreg[207]), .B(n3477), .Z(n3479) );
  NANDN U3610 ( .A(sreg[206]), .B(n3436), .Z(n3440) );
  NAND U3611 ( .A(n3438), .B(n3437), .Z(n3439) );
  NAND U3612 ( .A(n3440), .B(n3439), .Z(n3478) );
  XNOR U3613 ( .A(n3479), .B(n3478), .Z(c[207]) );
  NANDN U3614 ( .A(n3442), .B(n3441), .Z(n3446) );
  NANDN U3615 ( .A(n3444), .B(n3443), .Z(n3445) );
  AND U3616 ( .A(n3446), .B(n3445), .Z(n3485) );
  NANDN U3617 ( .A(n3448), .B(n3447), .Z(n3452) );
  NANDN U3618 ( .A(n3450), .B(n3449), .Z(n3451) );
  AND U3619 ( .A(n3452), .B(n3451), .Z(n3483) );
  NANDN U3620 ( .A(n5274), .B(n3453), .Z(n3455) );
  XOR U3621 ( .A(b[7]), .B(a[82]), .Z(n3494) );
  NANDN U3622 ( .A(n5275), .B(n3494), .Z(n3454) );
  AND U3623 ( .A(n3455), .B(n3454), .Z(n3513) );
  NANDN U3624 ( .A(n5176), .B(n3456), .Z(n3458) );
  XOR U3625 ( .A(b[3]), .B(a[86]), .Z(n3497) );
  NANDN U3626 ( .A(n5177), .B(n3497), .Z(n3457) );
  NAND U3627 ( .A(n3458), .B(n3457), .Z(n3512) );
  XNOR U3628 ( .A(n3513), .B(n3512), .Z(n3515) );
  NANDN U3629 ( .A(n5249), .B(n3459), .Z(n3461) );
  XOR U3630 ( .A(b[5]), .B(a[84]), .Z(n3503) );
  NANDN U3631 ( .A(n5184), .B(n3503), .Z(n3460) );
  AND U3632 ( .A(n3461), .B(n3460), .Z(n3507) );
  AND U3633 ( .A(b[7]), .B(a[80]), .Z(n3506) );
  XNOR U3634 ( .A(n3507), .B(n3506), .Z(n3508) );
  NAND U3635 ( .A(b[0]), .B(a[88]), .Z(n3462) );
  XNOR U3636 ( .A(b[1]), .B(n3462), .Z(n3464) );
  NANDN U3637 ( .A(b[0]), .B(a[87]), .Z(n3463) );
  NAND U3638 ( .A(n3464), .B(n3463), .Z(n3509) );
  XNOR U3639 ( .A(n3508), .B(n3509), .Z(n3514) );
  XOR U3640 ( .A(n3515), .B(n3514), .Z(n3489) );
  NANDN U3641 ( .A(n3466), .B(n3465), .Z(n3470) );
  NANDN U3642 ( .A(n3468), .B(n3467), .Z(n3469) );
  AND U3643 ( .A(n3470), .B(n3469), .Z(n3488) );
  XNOR U3644 ( .A(n3489), .B(n3488), .Z(n3490) );
  NANDN U3645 ( .A(n3472), .B(n3471), .Z(n3476) );
  NAND U3646 ( .A(n3474), .B(n3473), .Z(n3475) );
  NAND U3647 ( .A(n3476), .B(n3475), .Z(n3491) );
  XNOR U3648 ( .A(n3490), .B(n3491), .Z(n3482) );
  XNOR U3649 ( .A(n3483), .B(n3482), .Z(n3484) );
  XNOR U3650 ( .A(n3485), .B(n3484), .Z(n3518) );
  XNOR U3651 ( .A(sreg[208]), .B(n3518), .Z(n3520) );
  NANDN U3652 ( .A(sreg[207]), .B(n3477), .Z(n3481) );
  NAND U3653 ( .A(n3479), .B(n3478), .Z(n3480) );
  NAND U3654 ( .A(n3481), .B(n3480), .Z(n3519) );
  XNOR U3655 ( .A(n3520), .B(n3519), .Z(c[208]) );
  NANDN U3656 ( .A(n3483), .B(n3482), .Z(n3487) );
  NANDN U3657 ( .A(n3485), .B(n3484), .Z(n3486) );
  AND U3658 ( .A(n3487), .B(n3486), .Z(n3526) );
  NANDN U3659 ( .A(n3489), .B(n3488), .Z(n3493) );
  NANDN U3660 ( .A(n3491), .B(n3490), .Z(n3492) );
  AND U3661 ( .A(n3493), .B(n3492), .Z(n3524) );
  NANDN U3662 ( .A(n5274), .B(n3494), .Z(n3496) );
  XOR U3663 ( .A(b[7]), .B(a[83]), .Z(n3535) );
  NANDN U3664 ( .A(n5275), .B(n3535), .Z(n3495) );
  AND U3665 ( .A(n3496), .B(n3495), .Z(n3554) );
  NANDN U3666 ( .A(n5176), .B(n3497), .Z(n3499) );
  XOR U3667 ( .A(b[3]), .B(a[87]), .Z(n3538) );
  NANDN U3668 ( .A(n5177), .B(n3538), .Z(n3498) );
  NAND U3669 ( .A(n3499), .B(n3498), .Z(n3553) );
  XNOR U3670 ( .A(n3554), .B(n3553), .Z(n3556) );
  NAND U3671 ( .A(b[0]), .B(a[89]), .Z(n3500) );
  XNOR U3672 ( .A(b[1]), .B(n3500), .Z(n3502) );
  NANDN U3673 ( .A(b[0]), .B(a[88]), .Z(n3501) );
  NAND U3674 ( .A(n3502), .B(n3501), .Z(n3550) );
  NANDN U3675 ( .A(n5249), .B(n3503), .Z(n3505) );
  XOR U3676 ( .A(b[5]), .B(a[85]), .Z(n3544) );
  NANDN U3677 ( .A(n5184), .B(n3544), .Z(n3504) );
  AND U3678 ( .A(n3505), .B(n3504), .Z(n3548) );
  AND U3679 ( .A(b[7]), .B(a[81]), .Z(n3547) );
  XNOR U3680 ( .A(n3548), .B(n3547), .Z(n3549) );
  XNOR U3681 ( .A(n3550), .B(n3549), .Z(n3555) );
  XOR U3682 ( .A(n3556), .B(n3555), .Z(n3530) );
  NANDN U3683 ( .A(n3507), .B(n3506), .Z(n3511) );
  NANDN U3684 ( .A(n3509), .B(n3508), .Z(n3510) );
  AND U3685 ( .A(n3511), .B(n3510), .Z(n3529) );
  XNOR U3686 ( .A(n3530), .B(n3529), .Z(n3531) );
  NANDN U3687 ( .A(n3513), .B(n3512), .Z(n3517) );
  NAND U3688 ( .A(n3515), .B(n3514), .Z(n3516) );
  NAND U3689 ( .A(n3517), .B(n3516), .Z(n3532) );
  XNOR U3690 ( .A(n3531), .B(n3532), .Z(n3523) );
  XNOR U3691 ( .A(n3524), .B(n3523), .Z(n3525) );
  XNOR U3692 ( .A(n3526), .B(n3525), .Z(n3559) );
  XNOR U3693 ( .A(sreg[209]), .B(n3559), .Z(n3561) );
  NANDN U3694 ( .A(sreg[208]), .B(n3518), .Z(n3522) );
  NAND U3695 ( .A(n3520), .B(n3519), .Z(n3521) );
  NAND U3696 ( .A(n3522), .B(n3521), .Z(n3560) );
  XNOR U3697 ( .A(n3561), .B(n3560), .Z(c[209]) );
  NANDN U3698 ( .A(n3524), .B(n3523), .Z(n3528) );
  NANDN U3699 ( .A(n3526), .B(n3525), .Z(n3527) );
  AND U3700 ( .A(n3528), .B(n3527), .Z(n3567) );
  NANDN U3701 ( .A(n3530), .B(n3529), .Z(n3534) );
  NANDN U3702 ( .A(n3532), .B(n3531), .Z(n3533) );
  AND U3703 ( .A(n3534), .B(n3533), .Z(n3565) );
  NANDN U3704 ( .A(n5274), .B(n3535), .Z(n3537) );
  XOR U3705 ( .A(b[7]), .B(a[84]), .Z(n3576) );
  NANDN U3706 ( .A(n5275), .B(n3576), .Z(n3536) );
  AND U3707 ( .A(n3537), .B(n3536), .Z(n3595) );
  NANDN U3708 ( .A(n5176), .B(n3538), .Z(n3540) );
  XOR U3709 ( .A(b[3]), .B(a[88]), .Z(n3579) );
  NANDN U3710 ( .A(n5177), .B(n3579), .Z(n3539) );
  NAND U3711 ( .A(n3540), .B(n3539), .Z(n3594) );
  XNOR U3712 ( .A(n3595), .B(n3594), .Z(n3597) );
  NAND U3713 ( .A(b[0]), .B(a[90]), .Z(n3541) );
  XNOR U3714 ( .A(b[1]), .B(n3541), .Z(n3543) );
  NANDN U3715 ( .A(b[0]), .B(a[89]), .Z(n3542) );
  NAND U3716 ( .A(n3543), .B(n3542), .Z(n3591) );
  NANDN U3717 ( .A(n5249), .B(n3544), .Z(n3546) );
  XOR U3718 ( .A(b[5]), .B(a[86]), .Z(n3585) );
  NANDN U3719 ( .A(n5184), .B(n3585), .Z(n3545) );
  AND U3720 ( .A(n3546), .B(n3545), .Z(n3589) );
  AND U3721 ( .A(b[7]), .B(a[82]), .Z(n3588) );
  XNOR U3722 ( .A(n3589), .B(n3588), .Z(n3590) );
  XNOR U3723 ( .A(n3591), .B(n3590), .Z(n3596) );
  XOR U3724 ( .A(n3597), .B(n3596), .Z(n3571) );
  NANDN U3725 ( .A(n3548), .B(n3547), .Z(n3552) );
  NANDN U3726 ( .A(n3550), .B(n3549), .Z(n3551) );
  AND U3727 ( .A(n3552), .B(n3551), .Z(n3570) );
  XNOR U3728 ( .A(n3571), .B(n3570), .Z(n3572) );
  NANDN U3729 ( .A(n3554), .B(n3553), .Z(n3558) );
  NAND U3730 ( .A(n3556), .B(n3555), .Z(n3557) );
  NAND U3731 ( .A(n3558), .B(n3557), .Z(n3573) );
  XNOR U3732 ( .A(n3572), .B(n3573), .Z(n3564) );
  XNOR U3733 ( .A(n3565), .B(n3564), .Z(n3566) );
  XNOR U3734 ( .A(n3567), .B(n3566), .Z(n3600) );
  XNOR U3735 ( .A(sreg[210]), .B(n3600), .Z(n3602) );
  NANDN U3736 ( .A(sreg[209]), .B(n3559), .Z(n3563) );
  NAND U3737 ( .A(n3561), .B(n3560), .Z(n3562) );
  NAND U3738 ( .A(n3563), .B(n3562), .Z(n3601) );
  XNOR U3739 ( .A(n3602), .B(n3601), .Z(c[210]) );
  NANDN U3740 ( .A(n3565), .B(n3564), .Z(n3569) );
  NANDN U3741 ( .A(n3567), .B(n3566), .Z(n3568) );
  AND U3742 ( .A(n3569), .B(n3568), .Z(n3608) );
  NANDN U3743 ( .A(n3571), .B(n3570), .Z(n3575) );
  NANDN U3744 ( .A(n3573), .B(n3572), .Z(n3574) );
  AND U3745 ( .A(n3575), .B(n3574), .Z(n3606) );
  NANDN U3746 ( .A(n5274), .B(n3576), .Z(n3578) );
  XOR U3747 ( .A(b[7]), .B(a[85]), .Z(n3617) );
  NANDN U3748 ( .A(n5275), .B(n3617), .Z(n3577) );
  AND U3749 ( .A(n3578), .B(n3577), .Z(n3636) );
  NANDN U3750 ( .A(n5176), .B(n3579), .Z(n3581) );
  XOR U3751 ( .A(b[3]), .B(a[89]), .Z(n3620) );
  NANDN U3752 ( .A(n5177), .B(n3620), .Z(n3580) );
  NAND U3753 ( .A(n3581), .B(n3580), .Z(n3635) );
  XNOR U3754 ( .A(n3636), .B(n3635), .Z(n3638) );
  NAND U3755 ( .A(b[0]), .B(a[91]), .Z(n3582) );
  XNOR U3756 ( .A(b[1]), .B(n3582), .Z(n3584) );
  NANDN U3757 ( .A(b[0]), .B(a[90]), .Z(n3583) );
  NAND U3758 ( .A(n3584), .B(n3583), .Z(n3632) );
  NANDN U3759 ( .A(n5249), .B(n3585), .Z(n3587) );
  XOR U3760 ( .A(b[5]), .B(a[87]), .Z(n3626) );
  NANDN U3761 ( .A(n5184), .B(n3626), .Z(n3586) );
  AND U3762 ( .A(n3587), .B(n3586), .Z(n3630) );
  AND U3763 ( .A(b[7]), .B(a[83]), .Z(n3629) );
  XNOR U3764 ( .A(n3630), .B(n3629), .Z(n3631) );
  XNOR U3765 ( .A(n3632), .B(n3631), .Z(n3637) );
  XOR U3766 ( .A(n3638), .B(n3637), .Z(n3612) );
  NANDN U3767 ( .A(n3589), .B(n3588), .Z(n3593) );
  NANDN U3768 ( .A(n3591), .B(n3590), .Z(n3592) );
  AND U3769 ( .A(n3593), .B(n3592), .Z(n3611) );
  XNOR U3770 ( .A(n3612), .B(n3611), .Z(n3613) );
  NANDN U3771 ( .A(n3595), .B(n3594), .Z(n3599) );
  NAND U3772 ( .A(n3597), .B(n3596), .Z(n3598) );
  NAND U3773 ( .A(n3599), .B(n3598), .Z(n3614) );
  XNOR U3774 ( .A(n3613), .B(n3614), .Z(n3605) );
  XNOR U3775 ( .A(n3606), .B(n3605), .Z(n3607) );
  XNOR U3776 ( .A(n3608), .B(n3607), .Z(n3641) );
  XNOR U3777 ( .A(sreg[211]), .B(n3641), .Z(n3643) );
  NANDN U3778 ( .A(sreg[210]), .B(n3600), .Z(n3604) );
  NAND U3779 ( .A(n3602), .B(n3601), .Z(n3603) );
  NAND U3780 ( .A(n3604), .B(n3603), .Z(n3642) );
  XNOR U3781 ( .A(n3643), .B(n3642), .Z(c[211]) );
  NANDN U3782 ( .A(n3606), .B(n3605), .Z(n3610) );
  NANDN U3783 ( .A(n3608), .B(n3607), .Z(n3609) );
  AND U3784 ( .A(n3610), .B(n3609), .Z(n3649) );
  NANDN U3785 ( .A(n3612), .B(n3611), .Z(n3616) );
  NANDN U3786 ( .A(n3614), .B(n3613), .Z(n3615) );
  AND U3787 ( .A(n3616), .B(n3615), .Z(n3647) );
  NANDN U3788 ( .A(n5274), .B(n3617), .Z(n3619) );
  XOR U3789 ( .A(b[7]), .B(a[86]), .Z(n3658) );
  NANDN U3790 ( .A(n5275), .B(n3658), .Z(n3618) );
  AND U3791 ( .A(n3619), .B(n3618), .Z(n3677) );
  NANDN U3792 ( .A(n5176), .B(n3620), .Z(n3622) );
  XOR U3793 ( .A(b[3]), .B(a[90]), .Z(n3661) );
  NANDN U3794 ( .A(n5177), .B(n3661), .Z(n3621) );
  NAND U3795 ( .A(n3622), .B(n3621), .Z(n3676) );
  XNOR U3796 ( .A(n3677), .B(n3676), .Z(n3679) );
  NAND U3797 ( .A(b[0]), .B(a[92]), .Z(n3623) );
  XNOR U3798 ( .A(b[1]), .B(n3623), .Z(n3625) );
  NANDN U3799 ( .A(b[0]), .B(a[91]), .Z(n3624) );
  NAND U3800 ( .A(n3625), .B(n3624), .Z(n3673) );
  NANDN U3801 ( .A(n5249), .B(n3626), .Z(n3628) );
  XOR U3802 ( .A(b[5]), .B(a[88]), .Z(n3667) );
  NANDN U3803 ( .A(n5184), .B(n3667), .Z(n3627) );
  AND U3804 ( .A(n3628), .B(n3627), .Z(n3671) );
  AND U3805 ( .A(b[7]), .B(a[84]), .Z(n3670) );
  XNOR U3806 ( .A(n3671), .B(n3670), .Z(n3672) );
  XNOR U3807 ( .A(n3673), .B(n3672), .Z(n3678) );
  XOR U3808 ( .A(n3679), .B(n3678), .Z(n3653) );
  NANDN U3809 ( .A(n3630), .B(n3629), .Z(n3634) );
  NANDN U3810 ( .A(n3632), .B(n3631), .Z(n3633) );
  AND U3811 ( .A(n3634), .B(n3633), .Z(n3652) );
  XNOR U3812 ( .A(n3653), .B(n3652), .Z(n3654) );
  NANDN U3813 ( .A(n3636), .B(n3635), .Z(n3640) );
  NAND U3814 ( .A(n3638), .B(n3637), .Z(n3639) );
  NAND U3815 ( .A(n3640), .B(n3639), .Z(n3655) );
  XNOR U3816 ( .A(n3654), .B(n3655), .Z(n3646) );
  XNOR U3817 ( .A(n3647), .B(n3646), .Z(n3648) );
  XNOR U3818 ( .A(n3649), .B(n3648), .Z(n3682) );
  XNOR U3819 ( .A(sreg[212]), .B(n3682), .Z(n3684) );
  NANDN U3820 ( .A(sreg[211]), .B(n3641), .Z(n3645) );
  NAND U3821 ( .A(n3643), .B(n3642), .Z(n3644) );
  NAND U3822 ( .A(n3645), .B(n3644), .Z(n3683) );
  XNOR U3823 ( .A(n3684), .B(n3683), .Z(c[212]) );
  NANDN U3824 ( .A(n3647), .B(n3646), .Z(n3651) );
  NANDN U3825 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U3826 ( .A(n3651), .B(n3650), .Z(n3690) );
  NANDN U3827 ( .A(n3653), .B(n3652), .Z(n3657) );
  NANDN U3828 ( .A(n3655), .B(n3654), .Z(n3656) );
  AND U3829 ( .A(n3657), .B(n3656), .Z(n3688) );
  NANDN U3830 ( .A(n5274), .B(n3658), .Z(n3660) );
  XOR U3831 ( .A(b[7]), .B(a[87]), .Z(n3699) );
  NANDN U3832 ( .A(n5275), .B(n3699), .Z(n3659) );
  AND U3833 ( .A(n3660), .B(n3659), .Z(n3718) );
  NANDN U3834 ( .A(n5176), .B(n3661), .Z(n3663) );
  XOR U3835 ( .A(b[3]), .B(a[91]), .Z(n3702) );
  NANDN U3836 ( .A(n5177), .B(n3702), .Z(n3662) );
  NAND U3837 ( .A(n3663), .B(n3662), .Z(n3717) );
  XNOR U3838 ( .A(n3718), .B(n3717), .Z(n3720) );
  NAND U3839 ( .A(b[0]), .B(a[93]), .Z(n3664) );
  XNOR U3840 ( .A(b[1]), .B(n3664), .Z(n3666) );
  NANDN U3841 ( .A(b[0]), .B(a[92]), .Z(n3665) );
  NAND U3842 ( .A(n3666), .B(n3665), .Z(n3714) );
  NANDN U3843 ( .A(n5249), .B(n3667), .Z(n3669) );
  XOR U3844 ( .A(b[5]), .B(a[89]), .Z(n3708) );
  NANDN U3845 ( .A(n5184), .B(n3708), .Z(n3668) );
  AND U3846 ( .A(n3669), .B(n3668), .Z(n3712) );
  AND U3847 ( .A(b[7]), .B(a[85]), .Z(n3711) );
  XNOR U3848 ( .A(n3712), .B(n3711), .Z(n3713) );
  XNOR U3849 ( .A(n3714), .B(n3713), .Z(n3719) );
  XOR U3850 ( .A(n3720), .B(n3719), .Z(n3694) );
  NANDN U3851 ( .A(n3671), .B(n3670), .Z(n3675) );
  NANDN U3852 ( .A(n3673), .B(n3672), .Z(n3674) );
  AND U3853 ( .A(n3675), .B(n3674), .Z(n3693) );
  XNOR U3854 ( .A(n3694), .B(n3693), .Z(n3695) );
  NANDN U3855 ( .A(n3677), .B(n3676), .Z(n3681) );
  NAND U3856 ( .A(n3679), .B(n3678), .Z(n3680) );
  NAND U3857 ( .A(n3681), .B(n3680), .Z(n3696) );
  XNOR U3858 ( .A(n3695), .B(n3696), .Z(n3687) );
  XNOR U3859 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U3860 ( .A(n3690), .B(n3689), .Z(n3723) );
  XNOR U3861 ( .A(sreg[213]), .B(n3723), .Z(n3725) );
  NANDN U3862 ( .A(sreg[212]), .B(n3682), .Z(n3686) );
  NAND U3863 ( .A(n3684), .B(n3683), .Z(n3685) );
  NAND U3864 ( .A(n3686), .B(n3685), .Z(n3724) );
  XNOR U3865 ( .A(n3725), .B(n3724), .Z(c[213]) );
  NANDN U3866 ( .A(n3688), .B(n3687), .Z(n3692) );
  NANDN U3867 ( .A(n3690), .B(n3689), .Z(n3691) );
  AND U3868 ( .A(n3692), .B(n3691), .Z(n3731) );
  NANDN U3869 ( .A(n3694), .B(n3693), .Z(n3698) );
  NANDN U3870 ( .A(n3696), .B(n3695), .Z(n3697) );
  AND U3871 ( .A(n3698), .B(n3697), .Z(n3729) );
  NANDN U3872 ( .A(n5274), .B(n3699), .Z(n3701) );
  XOR U3873 ( .A(b[7]), .B(a[88]), .Z(n3740) );
  NANDN U3874 ( .A(n5275), .B(n3740), .Z(n3700) );
  AND U3875 ( .A(n3701), .B(n3700), .Z(n3759) );
  NANDN U3876 ( .A(n5176), .B(n3702), .Z(n3704) );
  XOR U3877 ( .A(b[3]), .B(a[92]), .Z(n3743) );
  NANDN U3878 ( .A(n5177), .B(n3743), .Z(n3703) );
  NAND U3879 ( .A(n3704), .B(n3703), .Z(n3758) );
  XNOR U3880 ( .A(n3759), .B(n3758), .Z(n3761) );
  NAND U3881 ( .A(b[0]), .B(a[94]), .Z(n3705) );
  XNOR U3882 ( .A(b[1]), .B(n3705), .Z(n3707) );
  NANDN U3883 ( .A(b[0]), .B(a[93]), .Z(n3706) );
  NAND U3884 ( .A(n3707), .B(n3706), .Z(n3755) );
  NANDN U3885 ( .A(n5249), .B(n3708), .Z(n3710) );
  XOR U3886 ( .A(b[5]), .B(a[90]), .Z(n3749) );
  NANDN U3887 ( .A(n5184), .B(n3749), .Z(n3709) );
  AND U3888 ( .A(n3710), .B(n3709), .Z(n3753) );
  AND U3889 ( .A(b[7]), .B(a[86]), .Z(n3752) );
  XNOR U3890 ( .A(n3753), .B(n3752), .Z(n3754) );
  XNOR U3891 ( .A(n3755), .B(n3754), .Z(n3760) );
  XOR U3892 ( .A(n3761), .B(n3760), .Z(n3735) );
  NANDN U3893 ( .A(n3712), .B(n3711), .Z(n3716) );
  NANDN U3894 ( .A(n3714), .B(n3713), .Z(n3715) );
  AND U3895 ( .A(n3716), .B(n3715), .Z(n3734) );
  XNOR U3896 ( .A(n3735), .B(n3734), .Z(n3736) );
  NANDN U3897 ( .A(n3718), .B(n3717), .Z(n3722) );
  NAND U3898 ( .A(n3720), .B(n3719), .Z(n3721) );
  NAND U3899 ( .A(n3722), .B(n3721), .Z(n3737) );
  XNOR U3900 ( .A(n3736), .B(n3737), .Z(n3728) );
  XNOR U3901 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U3902 ( .A(n3731), .B(n3730), .Z(n3764) );
  XNOR U3903 ( .A(sreg[214]), .B(n3764), .Z(n3766) );
  NANDN U3904 ( .A(sreg[213]), .B(n3723), .Z(n3727) );
  NAND U3905 ( .A(n3725), .B(n3724), .Z(n3726) );
  NAND U3906 ( .A(n3727), .B(n3726), .Z(n3765) );
  XNOR U3907 ( .A(n3766), .B(n3765), .Z(c[214]) );
  NANDN U3908 ( .A(n3729), .B(n3728), .Z(n3733) );
  NANDN U3909 ( .A(n3731), .B(n3730), .Z(n3732) );
  AND U3910 ( .A(n3733), .B(n3732), .Z(n3772) );
  NANDN U3911 ( .A(n3735), .B(n3734), .Z(n3739) );
  NANDN U3912 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U3913 ( .A(n3739), .B(n3738), .Z(n3770) );
  NANDN U3914 ( .A(n5274), .B(n3740), .Z(n3742) );
  XOR U3915 ( .A(b[7]), .B(a[89]), .Z(n3781) );
  NANDN U3916 ( .A(n5275), .B(n3781), .Z(n3741) );
  AND U3917 ( .A(n3742), .B(n3741), .Z(n3800) );
  NANDN U3918 ( .A(n5176), .B(n3743), .Z(n3745) );
  XOR U3919 ( .A(b[3]), .B(a[93]), .Z(n3784) );
  NANDN U3920 ( .A(n5177), .B(n3784), .Z(n3744) );
  NAND U3921 ( .A(n3745), .B(n3744), .Z(n3799) );
  XNOR U3922 ( .A(n3800), .B(n3799), .Z(n3802) );
  NAND U3923 ( .A(b[0]), .B(a[95]), .Z(n3746) );
  XNOR U3924 ( .A(b[1]), .B(n3746), .Z(n3748) );
  NANDN U3925 ( .A(b[0]), .B(a[94]), .Z(n3747) );
  NAND U3926 ( .A(n3748), .B(n3747), .Z(n3796) );
  NANDN U3927 ( .A(n5249), .B(n3749), .Z(n3751) );
  XOR U3928 ( .A(b[5]), .B(a[91]), .Z(n3787) );
  NANDN U3929 ( .A(n5184), .B(n3787), .Z(n3750) );
  AND U3930 ( .A(n3751), .B(n3750), .Z(n3794) );
  AND U3931 ( .A(b[7]), .B(a[87]), .Z(n3793) );
  XNOR U3932 ( .A(n3794), .B(n3793), .Z(n3795) );
  XNOR U3933 ( .A(n3796), .B(n3795), .Z(n3801) );
  XOR U3934 ( .A(n3802), .B(n3801), .Z(n3776) );
  NANDN U3935 ( .A(n3753), .B(n3752), .Z(n3757) );
  NANDN U3936 ( .A(n3755), .B(n3754), .Z(n3756) );
  AND U3937 ( .A(n3757), .B(n3756), .Z(n3775) );
  XNOR U3938 ( .A(n3776), .B(n3775), .Z(n3777) );
  NANDN U3939 ( .A(n3759), .B(n3758), .Z(n3763) );
  NAND U3940 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U3941 ( .A(n3763), .B(n3762), .Z(n3778) );
  XNOR U3942 ( .A(n3777), .B(n3778), .Z(n3769) );
  XNOR U3943 ( .A(n3770), .B(n3769), .Z(n3771) );
  XNOR U3944 ( .A(n3772), .B(n3771), .Z(n3805) );
  XNOR U3945 ( .A(sreg[215]), .B(n3805), .Z(n3807) );
  NANDN U3946 ( .A(sreg[214]), .B(n3764), .Z(n3768) );
  NAND U3947 ( .A(n3766), .B(n3765), .Z(n3767) );
  NAND U3948 ( .A(n3768), .B(n3767), .Z(n3806) );
  XNOR U3949 ( .A(n3807), .B(n3806), .Z(c[215]) );
  NANDN U3950 ( .A(n3770), .B(n3769), .Z(n3774) );
  NANDN U3951 ( .A(n3772), .B(n3771), .Z(n3773) );
  AND U3952 ( .A(n3774), .B(n3773), .Z(n3813) );
  NANDN U3953 ( .A(n3776), .B(n3775), .Z(n3780) );
  NANDN U3954 ( .A(n3778), .B(n3777), .Z(n3779) );
  AND U3955 ( .A(n3780), .B(n3779), .Z(n3811) );
  NANDN U3956 ( .A(n5274), .B(n3781), .Z(n3783) );
  XOR U3957 ( .A(b[7]), .B(a[90]), .Z(n3822) );
  NANDN U3958 ( .A(n5275), .B(n3822), .Z(n3782) );
  AND U3959 ( .A(n3783), .B(n3782), .Z(n3841) );
  NANDN U3960 ( .A(n5176), .B(n3784), .Z(n3786) );
  XOR U3961 ( .A(b[3]), .B(a[94]), .Z(n3825) );
  NANDN U3962 ( .A(n5177), .B(n3825), .Z(n3785) );
  NAND U3963 ( .A(n3786), .B(n3785), .Z(n3840) );
  XNOR U3964 ( .A(n3841), .B(n3840), .Z(n3843) );
  NANDN U3965 ( .A(n5249), .B(n3787), .Z(n3789) );
  XOR U3966 ( .A(b[5]), .B(a[92]), .Z(n3831) );
  NANDN U3967 ( .A(n5184), .B(n3831), .Z(n3788) );
  AND U3968 ( .A(n3789), .B(n3788), .Z(n3835) );
  AND U3969 ( .A(b[7]), .B(a[88]), .Z(n3834) );
  XNOR U3970 ( .A(n3835), .B(n3834), .Z(n3836) );
  NAND U3971 ( .A(b[0]), .B(a[96]), .Z(n3790) );
  XNOR U3972 ( .A(b[1]), .B(n3790), .Z(n3792) );
  NANDN U3973 ( .A(b[0]), .B(a[95]), .Z(n3791) );
  NAND U3974 ( .A(n3792), .B(n3791), .Z(n3837) );
  XNOR U3975 ( .A(n3836), .B(n3837), .Z(n3842) );
  XOR U3976 ( .A(n3843), .B(n3842), .Z(n3817) );
  NANDN U3977 ( .A(n3794), .B(n3793), .Z(n3798) );
  NANDN U3978 ( .A(n3796), .B(n3795), .Z(n3797) );
  AND U3979 ( .A(n3798), .B(n3797), .Z(n3816) );
  XNOR U3980 ( .A(n3817), .B(n3816), .Z(n3818) );
  NANDN U3981 ( .A(n3800), .B(n3799), .Z(n3804) );
  NAND U3982 ( .A(n3802), .B(n3801), .Z(n3803) );
  NAND U3983 ( .A(n3804), .B(n3803), .Z(n3819) );
  XNOR U3984 ( .A(n3818), .B(n3819), .Z(n3810) );
  XNOR U3985 ( .A(n3811), .B(n3810), .Z(n3812) );
  XNOR U3986 ( .A(n3813), .B(n3812), .Z(n3846) );
  XNOR U3987 ( .A(sreg[216]), .B(n3846), .Z(n3848) );
  NANDN U3988 ( .A(sreg[215]), .B(n3805), .Z(n3809) );
  NAND U3989 ( .A(n3807), .B(n3806), .Z(n3808) );
  NAND U3990 ( .A(n3809), .B(n3808), .Z(n3847) );
  XNOR U3991 ( .A(n3848), .B(n3847), .Z(c[216]) );
  NANDN U3992 ( .A(n3811), .B(n3810), .Z(n3815) );
  NANDN U3993 ( .A(n3813), .B(n3812), .Z(n3814) );
  AND U3994 ( .A(n3815), .B(n3814), .Z(n3854) );
  NANDN U3995 ( .A(n3817), .B(n3816), .Z(n3821) );
  NANDN U3996 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U3997 ( .A(n3821), .B(n3820), .Z(n3852) );
  NANDN U3998 ( .A(n5274), .B(n3822), .Z(n3824) );
  XOR U3999 ( .A(b[7]), .B(a[91]), .Z(n3863) );
  NANDN U4000 ( .A(n5275), .B(n3863), .Z(n3823) );
  AND U4001 ( .A(n3824), .B(n3823), .Z(n3882) );
  NANDN U4002 ( .A(n5176), .B(n3825), .Z(n3827) );
  XOR U4003 ( .A(b[3]), .B(a[95]), .Z(n3866) );
  NANDN U4004 ( .A(n5177), .B(n3866), .Z(n3826) );
  NAND U4005 ( .A(n3827), .B(n3826), .Z(n3881) );
  XNOR U4006 ( .A(n3882), .B(n3881), .Z(n3884) );
  AND U4007 ( .A(b[0]), .B(a[97]), .Z(n3828) );
  XOR U4008 ( .A(b[1]), .B(n3828), .Z(n3830) );
  NANDN U4009 ( .A(b[0]), .B(a[96]), .Z(n3829) );
  AND U4010 ( .A(n3830), .B(n3829), .Z(n3877) );
  NANDN U4011 ( .A(n5249), .B(n3831), .Z(n3833) );
  XOR U4012 ( .A(b[5]), .B(a[93]), .Z(n3872) );
  NANDN U4013 ( .A(n5184), .B(n3872), .Z(n3832) );
  AND U4014 ( .A(n3833), .B(n3832), .Z(n3876) );
  AND U4015 ( .A(b[7]), .B(a[89]), .Z(n3875) );
  XOR U4016 ( .A(n3876), .B(n3875), .Z(n3878) );
  XNOR U4017 ( .A(n3877), .B(n3878), .Z(n3883) );
  XOR U4018 ( .A(n3884), .B(n3883), .Z(n3858) );
  NANDN U4019 ( .A(n3835), .B(n3834), .Z(n3839) );
  NANDN U4020 ( .A(n3837), .B(n3836), .Z(n3838) );
  AND U4021 ( .A(n3839), .B(n3838), .Z(n3857) );
  XNOR U4022 ( .A(n3858), .B(n3857), .Z(n3859) );
  NANDN U4023 ( .A(n3841), .B(n3840), .Z(n3845) );
  NAND U4024 ( .A(n3843), .B(n3842), .Z(n3844) );
  NAND U4025 ( .A(n3845), .B(n3844), .Z(n3860) );
  XNOR U4026 ( .A(n3859), .B(n3860), .Z(n3851) );
  XNOR U4027 ( .A(n3852), .B(n3851), .Z(n3853) );
  XNOR U4028 ( .A(n3854), .B(n3853), .Z(n3887) );
  XNOR U4029 ( .A(sreg[217]), .B(n3887), .Z(n3889) );
  NANDN U4030 ( .A(sreg[216]), .B(n3846), .Z(n3850) );
  NAND U4031 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U4032 ( .A(n3850), .B(n3849), .Z(n3888) );
  XNOR U4033 ( .A(n3889), .B(n3888), .Z(c[217]) );
  NANDN U4034 ( .A(n3852), .B(n3851), .Z(n3856) );
  NANDN U4035 ( .A(n3854), .B(n3853), .Z(n3855) );
  AND U4036 ( .A(n3856), .B(n3855), .Z(n3895) );
  NANDN U4037 ( .A(n3858), .B(n3857), .Z(n3862) );
  NANDN U4038 ( .A(n3860), .B(n3859), .Z(n3861) );
  AND U4039 ( .A(n3862), .B(n3861), .Z(n3893) );
  NANDN U4040 ( .A(n5274), .B(n3863), .Z(n3865) );
  XOR U4041 ( .A(b[7]), .B(a[92]), .Z(n3904) );
  NANDN U4042 ( .A(n5275), .B(n3904), .Z(n3864) );
  AND U4043 ( .A(n3865), .B(n3864), .Z(n3923) );
  NANDN U4044 ( .A(n5176), .B(n3866), .Z(n3868) );
  XOR U4045 ( .A(b[3]), .B(a[96]), .Z(n3907) );
  NANDN U4046 ( .A(n5177), .B(n3907), .Z(n3867) );
  NAND U4047 ( .A(n3868), .B(n3867), .Z(n3922) );
  XNOR U4048 ( .A(n3923), .B(n3922), .Z(n3925) );
  NAND U4049 ( .A(b[0]), .B(a[98]), .Z(n3869) );
  XNOR U4050 ( .A(b[1]), .B(n3869), .Z(n3871) );
  NANDN U4051 ( .A(b[0]), .B(a[97]), .Z(n3870) );
  NAND U4052 ( .A(n3871), .B(n3870), .Z(n3919) );
  NANDN U4053 ( .A(n5249), .B(n3872), .Z(n3874) );
  XOR U4054 ( .A(b[5]), .B(a[94]), .Z(n3913) );
  NANDN U4055 ( .A(n5184), .B(n3913), .Z(n3873) );
  AND U4056 ( .A(n3874), .B(n3873), .Z(n3917) );
  AND U4057 ( .A(b[7]), .B(a[90]), .Z(n3916) );
  XNOR U4058 ( .A(n3917), .B(n3916), .Z(n3918) );
  XNOR U4059 ( .A(n3919), .B(n3918), .Z(n3924) );
  XOR U4060 ( .A(n3925), .B(n3924), .Z(n3899) );
  NANDN U4061 ( .A(n3876), .B(n3875), .Z(n3880) );
  NANDN U4062 ( .A(n3878), .B(n3877), .Z(n3879) );
  AND U4063 ( .A(n3880), .B(n3879), .Z(n3898) );
  XNOR U4064 ( .A(n3899), .B(n3898), .Z(n3900) );
  NANDN U4065 ( .A(n3882), .B(n3881), .Z(n3886) );
  NAND U4066 ( .A(n3884), .B(n3883), .Z(n3885) );
  NAND U4067 ( .A(n3886), .B(n3885), .Z(n3901) );
  XNOR U4068 ( .A(n3900), .B(n3901), .Z(n3892) );
  XNOR U4069 ( .A(n3893), .B(n3892), .Z(n3894) );
  XNOR U4070 ( .A(n3895), .B(n3894), .Z(n3928) );
  XNOR U4071 ( .A(sreg[218]), .B(n3928), .Z(n3930) );
  NANDN U4072 ( .A(sreg[217]), .B(n3887), .Z(n3891) );
  NAND U4073 ( .A(n3889), .B(n3888), .Z(n3890) );
  NAND U4074 ( .A(n3891), .B(n3890), .Z(n3929) );
  XNOR U4075 ( .A(n3930), .B(n3929), .Z(c[218]) );
  NANDN U4076 ( .A(n3893), .B(n3892), .Z(n3897) );
  NANDN U4077 ( .A(n3895), .B(n3894), .Z(n3896) );
  AND U4078 ( .A(n3897), .B(n3896), .Z(n3936) );
  NANDN U4079 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4080 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4081 ( .A(n3903), .B(n3902), .Z(n3934) );
  NANDN U4082 ( .A(n5274), .B(n3904), .Z(n3906) );
  XOR U4083 ( .A(b[7]), .B(a[93]), .Z(n3945) );
  NANDN U4084 ( .A(n5275), .B(n3945), .Z(n3905) );
  AND U4085 ( .A(n3906), .B(n3905), .Z(n3964) );
  NANDN U4086 ( .A(n5176), .B(n3907), .Z(n3909) );
  XOR U4087 ( .A(b[3]), .B(a[97]), .Z(n3948) );
  NANDN U4088 ( .A(n5177), .B(n3948), .Z(n3908) );
  NAND U4089 ( .A(n3909), .B(n3908), .Z(n3963) );
  XNOR U4090 ( .A(n3964), .B(n3963), .Z(n3966) );
  NAND U4091 ( .A(b[0]), .B(a[99]), .Z(n3910) );
  XNOR U4092 ( .A(b[1]), .B(n3910), .Z(n3912) );
  NANDN U4093 ( .A(b[0]), .B(a[98]), .Z(n3911) );
  NAND U4094 ( .A(n3912), .B(n3911), .Z(n3960) );
  NANDN U4095 ( .A(n5249), .B(n3913), .Z(n3915) );
  XOR U4096 ( .A(b[5]), .B(a[95]), .Z(n3951) );
  NANDN U4097 ( .A(n5184), .B(n3951), .Z(n3914) );
  AND U4098 ( .A(n3915), .B(n3914), .Z(n3958) );
  AND U4099 ( .A(b[7]), .B(a[91]), .Z(n3957) );
  XNOR U4100 ( .A(n3958), .B(n3957), .Z(n3959) );
  XNOR U4101 ( .A(n3960), .B(n3959), .Z(n3965) );
  XOR U4102 ( .A(n3966), .B(n3965), .Z(n3940) );
  NANDN U4103 ( .A(n3917), .B(n3916), .Z(n3921) );
  NANDN U4104 ( .A(n3919), .B(n3918), .Z(n3920) );
  AND U4105 ( .A(n3921), .B(n3920), .Z(n3939) );
  XNOR U4106 ( .A(n3940), .B(n3939), .Z(n3941) );
  NANDN U4107 ( .A(n3923), .B(n3922), .Z(n3927) );
  NAND U4108 ( .A(n3925), .B(n3924), .Z(n3926) );
  NAND U4109 ( .A(n3927), .B(n3926), .Z(n3942) );
  XNOR U4110 ( .A(n3941), .B(n3942), .Z(n3933) );
  XNOR U4111 ( .A(n3934), .B(n3933), .Z(n3935) );
  XNOR U4112 ( .A(n3936), .B(n3935), .Z(n3969) );
  XNOR U4113 ( .A(sreg[219]), .B(n3969), .Z(n3971) );
  NANDN U4114 ( .A(sreg[218]), .B(n3928), .Z(n3932) );
  NAND U4115 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND U4116 ( .A(n3932), .B(n3931), .Z(n3970) );
  XNOR U4117 ( .A(n3971), .B(n3970), .Z(c[219]) );
  NANDN U4118 ( .A(n3934), .B(n3933), .Z(n3938) );
  NANDN U4119 ( .A(n3936), .B(n3935), .Z(n3937) );
  AND U4120 ( .A(n3938), .B(n3937), .Z(n3977) );
  NANDN U4121 ( .A(n3940), .B(n3939), .Z(n3944) );
  NANDN U4122 ( .A(n3942), .B(n3941), .Z(n3943) );
  AND U4123 ( .A(n3944), .B(n3943), .Z(n3975) );
  NANDN U4124 ( .A(n5274), .B(n3945), .Z(n3947) );
  XOR U4125 ( .A(b[7]), .B(a[94]), .Z(n3986) );
  NANDN U4126 ( .A(n5275), .B(n3986), .Z(n3946) );
  AND U4127 ( .A(n3947), .B(n3946), .Z(n4005) );
  NANDN U4128 ( .A(n5176), .B(n3948), .Z(n3950) );
  XOR U4129 ( .A(b[3]), .B(a[98]), .Z(n3989) );
  NANDN U4130 ( .A(n5177), .B(n3989), .Z(n3949) );
  NAND U4131 ( .A(n3950), .B(n3949), .Z(n4004) );
  XNOR U4132 ( .A(n4005), .B(n4004), .Z(n4007) );
  NANDN U4133 ( .A(n5249), .B(n3951), .Z(n3953) );
  XOR U4134 ( .A(b[5]), .B(a[96]), .Z(n3992) );
  NANDN U4135 ( .A(n5184), .B(n3992), .Z(n3952) );
  AND U4136 ( .A(n3953), .B(n3952), .Z(n3999) );
  AND U4137 ( .A(b[7]), .B(a[92]), .Z(n3998) );
  XNOR U4138 ( .A(n3999), .B(n3998), .Z(n4000) );
  NAND U4139 ( .A(b[0]), .B(a[100]), .Z(n3954) );
  XNOR U4140 ( .A(b[1]), .B(n3954), .Z(n3956) );
  NANDN U4141 ( .A(b[0]), .B(a[99]), .Z(n3955) );
  NAND U4142 ( .A(n3956), .B(n3955), .Z(n4001) );
  XNOR U4143 ( .A(n4000), .B(n4001), .Z(n4006) );
  XOR U4144 ( .A(n4007), .B(n4006), .Z(n3981) );
  NANDN U4145 ( .A(n3958), .B(n3957), .Z(n3962) );
  NANDN U4146 ( .A(n3960), .B(n3959), .Z(n3961) );
  AND U4147 ( .A(n3962), .B(n3961), .Z(n3980) );
  XNOR U4148 ( .A(n3981), .B(n3980), .Z(n3982) );
  NANDN U4149 ( .A(n3964), .B(n3963), .Z(n3968) );
  NAND U4150 ( .A(n3966), .B(n3965), .Z(n3967) );
  NAND U4151 ( .A(n3968), .B(n3967), .Z(n3983) );
  XNOR U4152 ( .A(n3982), .B(n3983), .Z(n3974) );
  XNOR U4153 ( .A(n3975), .B(n3974), .Z(n3976) );
  XNOR U4154 ( .A(n3977), .B(n3976), .Z(n4010) );
  XNOR U4155 ( .A(sreg[220]), .B(n4010), .Z(n4012) );
  NANDN U4156 ( .A(sreg[219]), .B(n3969), .Z(n3973) );
  NAND U4157 ( .A(n3971), .B(n3970), .Z(n3972) );
  NAND U4158 ( .A(n3973), .B(n3972), .Z(n4011) );
  XNOR U4159 ( .A(n4012), .B(n4011), .Z(c[220]) );
  NANDN U4160 ( .A(n3975), .B(n3974), .Z(n3979) );
  NANDN U4161 ( .A(n3977), .B(n3976), .Z(n3978) );
  AND U4162 ( .A(n3979), .B(n3978), .Z(n4018) );
  NANDN U4163 ( .A(n3981), .B(n3980), .Z(n3985) );
  NANDN U4164 ( .A(n3983), .B(n3982), .Z(n3984) );
  AND U4165 ( .A(n3985), .B(n3984), .Z(n4016) );
  NANDN U4166 ( .A(n5274), .B(n3986), .Z(n3988) );
  XOR U4167 ( .A(b[7]), .B(a[95]), .Z(n4027) );
  NANDN U4168 ( .A(n5275), .B(n4027), .Z(n3987) );
  AND U4169 ( .A(n3988), .B(n3987), .Z(n4046) );
  NANDN U4170 ( .A(n5176), .B(n3989), .Z(n3991) );
  XOR U4171 ( .A(b[3]), .B(a[99]), .Z(n4030) );
  NANDN U4172 ( .A(n5177), .B(n4030), .Z(n3990) );
  NAND U4173 ( .A(n3991), .B(n3990), .Z(n4045) );
  XNOR U4174 ( .A(n4046), .B(n4045), .Z(n4048) );
  NANDN U4175 ( .A(n5249), .B(n3992), .Z(n3994) );
  XOR U4176 ( .A(b[5]), .B(a[97]), .Z(n4036) );
  NANDN U4177 ( .A(n5184), .B(n4036), .Z(n3993) );
  AND U4178 ( .A(n3994), .B(n3993), .Z(n4040) );
  AND U4179 ( .A(b[7]), .B(a[93]), .Z(n4039) );
  XNOR U4180 ( .A(n4040), .B(n4039), .Z(n4041) );
  NAND U4181 ( .A(b[0]), .B(a[101]), .Z(n3995) );
  XNOR U4182 ( .A(b[1]), .B(n3995), .Z(n3997) );
  NANDN U4183 ( .A(b[0]), .B(a[100]), .Z(n3996) );
  NAND U4184 ( .A(n3997), .B(n3996), .Z(n4042) );
  XNOR U4185 ( .A(n4041), .B(n4042), .Z(n4047) );
  XOR U4186 ( .A(n4048), .B(n4047), .Z(n4022) );
  NANDN U4187 ( .A(n3999), .B(n3998), .Z(n4003) );
  NANDN U4188 ( .A(n4001), .B(n4000), .Z(n4002) );
  AND U4189 ( .A(n4003), .B(n4002), .Z(n4021) );
  XNOR U4190 ( .A(n4022), .B(n4021), .Z(n4023) );
  NANDN U4191 ( .A(n4005), .B(n4004), .Z(n4009) );
  NAND U4192 ( .A(n4007), .B(n4006), .Z(n4008) );
  NAND U4193 ( .A(n4009), .B(n4008), .Z(n4024) );
  XNOR U4194 ( .A(n4023), .B(n4024), .Z(n4015) );
  XNOR U4195 ( .A(n4016), .B(n4015), .Z(n4017) );
  XNOR U4196 ( .A(n4018), .B(n4017), .Z(n4051) );
  XNOR U4197 ( .A(sreg[221]), .B(n4051), .Z(n4053) );
  NANDN U4198 ( .A(sreg[220]), .B(n4010), .Z(n4014) );
  NAND U4199 ( .A(n4012), .B(n4011), .Z(n4013) );
  NAND U4200 ( .A(n4014), .B(n4013), .Z(n4052) );
  XNOR U4201 ( .A(n4053), .B(n4052), .Z(c[221]) );
  NANDN U4202 ( .A(n4016), .B(n4015), .Z(n4020) );
  NANDN U4203 ( .A(n4018), .B(n4017), .Z(n4019) );
  AND U4204 ( .A(n4020), .B(n4019), .Z(n4059) );
  NANDN U4205 ( .A(n4022), .B(n4021), .Z(n4026) );
  NANDN U4206 ( .A(n4024), .B(n4023), .Z(n4025) );
  AND U4207 ( .A(n4026), .B(n4025), .Z(n4057) );
  NANDN U4208 ( .A(n5274), .B(n4027), .Z(n4029) );
  XOR U4209 ( .A(b[7]), .B(a[96]), .Z(n4068) );
  NANDN U4210 ( .A(n5275), .B(n4068), .Z(n4028) );
  AND U4211 ( .A(n4029), .B(n4028), .Z(n4087) );
  NANDN U4212 ( .A(n5176), .B(n4030), .Z(n4032) );
  XOR U4213 ( .A(b[3]), .B(a[100]), .Z(n4071) );
  NANDN U4214 ( .A(n5177), .B(n4071), .Z(n4031) );
  NAND U4215 ( .A(n4032), .B(n4031), .Z(n4086) );
  XNOR U4216 ( .A(n4087), .B(n4086), .Z(n4089) );
  NAND U4217 ( .A(b[0]), .B(a[102]), .Z(n4033) );
  XNOR U4218 ( .A(b[1]), .B(n4033), .Z(n4035) );
  NANDN U4219 ( .A(b[0]), .B(a[101]), .Z(n4034) );
  NAND U4220 ( .A(n4035), .B(n4034), .Z(n4083) );
  NANDN U4221 ( .A(n5249), .B(n4036), .Z(n4038) );
  XOR U4222 ( .A(b[5]), .B(a[98]), .Z(n4077) );
  NANDN U4223 ( .A(n5184), .B(n4077), .Z(n4037) );
  AND U4224 ( .A(n4038), .B(n4037), .Z(n4081) );
  AND U4225 ( .A(b[7]), .B(a[94]), .Z(n4080) );
  XNOR U4226 ( .A(n4081), .B(n4080), .Z(n4082) );
  XNOR U4227 ( .A(n4083), .B(n4082), .Z(n4088) );
  XOR U4228 ( .A(n4089), .B(n4088), .Z(n4063) );
  NANDN U4229 ( .A(n4040), .B(n4039), .Z(n4044) );
  NANDN U4230 ( .A(n4042), .B(n4041), .Z(n4043) );
  AND U4231 ( .A(n4044), .B(n4043), .Z(n4062) );
  XNOR U4232 ( .A(n4063), .B(n4062), .Z(n4064) );
  NANDN U4233 ( .A(n4046), .B(n4045), .Z(n4050) );
  NAND U4234 ( .A(n4048), .B(n4047), .Z(n4049) );
  NAND U4235 ( .A(n4050), .B(n4049), .Z(n4065) );
  XNOR U4236 ( .A(n4064), .B(n4065), .Z(n4056) );
  XNOR U4237 ( .A(n4057), .B(n4056), .Z(n4058) );
  XNOR U4238 ( .A(n4059), .B(n4058), .Z(n4092) );
  XNOR U4239 ( .A(sreg[222]), .B(n4092), .Z(n4094) );
  NANDN U4240 ( .A(sreg[221]), .B(n4051), .Z(n4055) );
  NAND U4241 ( .A(n4053), .B(n4052), .Z(n4054) );
  NAND U4242 ( .A(n4055), .B(n4054), .Z(n4093) );
  XNOR U4243 ( .A(n4094), .B(n4093), .Z(c[222]) );
  NANDN U4244 ( .A(n4057), .B(n4056), .Z(n4061) );
  NANDN U4245 ( .A(n4059), .B(n4058), .Z(n4060) );
  AND U4246 ( .A(n4061), .B(n4060), .Z(n4100) );
  NANDN U4247 ( .A(n4063), .B(n4062), .Z(n4067) );
  NANDN U4248 ( .A(n4065), .B(n4064), .Z(n4066) );
  AND U4249 ( .A(n4067), .B(n4066), .Z(n4098) );
  NANDN U4250 ( .A(n5274), .B(n4068), .Z(n4070) );
  XOR U4251 ( .A(b[7]), .B(a[97]), .Z(n4109) );
  NANDN U4252 ( .A(n5275), .B(n4109), .Z(n4069) );
  AND U4253 ( .A(n4070), .B(n4069), .Z(n4128) );
  NANDN U4254 ( .A(n5176), .B(n4071), .Z(n4073) );
  XOR U4255 ( .A(b[3]), .B(a[101]), .Z(n4112) );
  NANDN U4256 ( .A(n5177), .B(n4112), .Z(n4072) );
  NAND U4257 ( .A(n4073), .B(n4072), .Z(n4127) );
  XNOR U4258 ( .A(n4128), .B(n4127), .Z(n4130) );
  NAND U4259 ( .A(b[0]), .B(a[103]), .Z(n4074) );
  XNOR U4260 ( .A(b[1]), .B(n4074), .Z(n4076) );
  NANDN U4261 ( .A(b[0]), .B(a[102]), .Z(n4075) );
  NAND U4262 ( .A(n4076), .B(n4075), .Z(n4124) );
  NANDN U4263 ( .A(n5249), .B(n4077), .Z(n4079) );
  XOR U4264 ( .A(b[5]), .B(a[99]), .Z(n4118) );
  NANDN U4265 ( .A(n5184), .B(n4118), .Z(n4078) );
  AND U4266 ( .A(n4079), .B(n4078), .Z(n4122) );
  AND U4267 ( .A(b[7]), .B(a[95]), .Z(n4121) );
  XNOR U4268 ( .A(n4122), .B(n4121), .Z(n4123) );
  XNOR U4269 ( .A(n4124), .B(n4123), .Z(n4129) );
  XOR U4270 ( .A(n4130), .B(n4129), .Z(n4104) );
  NANDN U4271 ( .A(n4081), .B(n4080), .Z(n4085) );
  NANDN U4272 ( .A(n4083), .B(n4082), .Z(n4084) );
  AND U4273 ( .A(n4085), .B(n4084), .Z(n4103) );
  XNOR U4274 ( .A(n4104), .B(n4103), .Z(n4105) );
  NANDN U4275 ( .A(n4087), .B(n4086), .Z(n4091) );
  NAND U4276 ( .A(n4089), .B(n4088), .Z(n4090) );
  NAND U4277 ( .A(n4091), .B(n4090), .Z(n4106) );
  XNOR U4278 ( .A(n4105), .B(n4106), .Z(n4097) );
  XNOR U4279 ( .A(n4098), .B(n4097), .Z(n4099) );
  XNOR U4280 ( .A(n4100), .B(n4099), .Z(n4133) );
  XNOR U4281 ( .A(sreg[223]), .B(n4133), .Z(n4135) );
  NANDN U4282 ( .A(sreg[222]), .B(n4092), .Z(n4096) );
  NAND U4283 ( .A(n4094), .B(n4093), .Z(n4095) );
  NAND U4284 ( .A(n4096), .B(n4095), .Z(n4134) );
  XNOR U4285 ( .A(n4135), .B(n4134), .Z(c[223]) );
  NANDN U4286 ( .A(n4098), .B(n4097), .Z(n4102) );
  NANDN U4287 ( .A(n4100), .B(n4099), .Z(n4101) );
  AND U4288 ( .A(n4102), .B(n4101), .Z(n4141) );
  NANDN U4289 ( .A(n4104), .B(n4103), .Z(n4108) );
  NANDN U4290 ( .A(n4106), .B(n4105), .Z(n4107) );
  AND U4291 ( .A(n4108), .B(n4107), .Z(n4139) );
  NANDN U4292 ( .A(n5274), .B(n4109), .Z(n4111) );
  XOR U4293 ( .A(b[7]), .B(a[98]), .Z(n4150) );
  NANDN U4294 ( .A(n5275), .B(n4150), .Z(n4110) );
  AND U4295 ( .A(n4111), .B(n4110), .Z(n4169) );
  NANDN U4296 ( .A(n5176), .B(n4112), .Z(n4114) );
  XOR U4297 ( .A(b[3]), .B(a[102]), .Z(n4153) );
  NANDN U4298 ( .A(n5177), .B(n4153), .Z(n4113) );
  NAND U4299 ( .A(n4114), .B(n4113), .Z(n4168) );
  XNOR U4300 ( .A(n4169), .B(n4168), .Z(n4171) );
  NAND U4301 ( .A(b[0]), .B(a[104]), .Z(n4115) );
  XNOR U4302 ( .A(b[1]), .B(n4115), .Z(n4117) );
  NANDN U4303 ( .A(b[0]), .B(a[103]), .Z(n4116) );
  NAND U4304 ( .A(n4117), .B(n4116), .Z(n4165) );
  NANDN U4305 ( .A(n5249), .B(n4118), .Z(n4120) );
  XOR U4306 ( .A(b[5]), .B(a[100]), .Z(n4159) );
  NANDN U4307 ( .A(n5184), .B(n4159), .Z(n4119) );
  AND U4308 ( .A(n4120), .B(n4119), .Z(n4163) );
  AND U4309 ( .A(b[7]), .B(a[96]), .Z(n4162) );
  XNOR U4310 ( .A(n4163), .B(n4162), .Z(n4164) );
  XNOR U4311 ( .A(n4165), .B(n4164), .Z(n4170) );
  XOR U4312 ( .A(n4171), .B(n4170), .Z(n4145) );
  NANDN U4313 ( .A(n4122), .B(n4121), .Z(n4126) );
  NANDN U4314 ( .A(n4124), .B(n4123), .Z(n4125) );
  AND U4315 ( .A(n4126), .B(n4125), .Z(n4144) );
  XNOR U4316 ( .A(n4145), .B(n4144), .Z(n4146) );
  NANDN U4317 ( .A(n4128), .B(n4127), .Z(n4132) );
  NAND U4318 ( .A(n4130), .B(n4129), .Z(n4131) );
  NAND U4319 ( .A(n4132), .B(n4131), .Z(n4147) );
  XNOR U4320 ( .A(n4146), .B(n4147), .Z(n4138) );
  XNOR U4321 ( .A(n4139), .B(n4138), .Z(n4140) );
  XNOR U4322 ( .A(n4141), .B(n4140), .Z(n4174) );
  XNOR U4323 ( .A(sreg[224]), .B(n4174), .Z(n4176) );
  NANDN U4324 ( .A(sreg[223]), .B(n4133), .Z(n4137) );
  NAND U4325 ( .A(n4135), .B(n4134), .Z(n4136) );
  NAND U4326 ( .A(n4137), .B(n4136), .Z(n4175) );
  XNOR U4327 ( .A(n4176), .B(n4175), .Z(c[224]) );
  NANDN U4328 ( .A(n4139), .B(n4138), .Z(n4143) );
  NANDN U4329 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U4330 ( .A(n4143), .B(n4142), .Z(n4182) );
  NANDN U4331 ( .A(n4145), .B(n4144), .Z(n4149) );
  NANDN U4332 ( .A(n4147), .B(n4146), .Z(n4148) );
  AND U4333 ( .A(n4149), .B(n4148), .Z(n4180) );
  NANDN U4334 ( .A(n5274), .B(n4150), .Z(n4152) );
  XOR U4335 ( .A(b[7]), .B(a[99]), .Z(n4191) );
  NANDN U4336 ( .A(n5275), .B(n4191), .Z(n4151) );
  AND U4337 ( .A(n4152), .B(n4151), .Z(n4210) );
  NANDN U4338 ( .A(n5176), .B(n4153), .Z(n4155) );
  XOR U4339 ( .A(b[3]), .B(a[103]), .Z(n4194) );
  NANDN U4340 ( .A(n5177), .B(n4194), .Z(n4154) );
  NAND U4341 ( .A(n4155), .B(n4154), .Z(n4209) );
  XNOR U4342 ( .A(n4210), .B(n4209), .Z(n4212) );
  NAND U4343 ( .A(b[0]), .B(a[105]), .Z(n4156) );
  XNOR U4344 ( .A(b[1]), .B(n4156), .Z(n4158) );
  NANDN U4345 ( .A(b[0]), .B(a[104]), .Z(n4157) );
  NAND U4346 ( .A(n4158), .B(n4157), .Z(n4206) );
  NANDN U4347 ( .A(n5249), .B(n4159), .Z(n4161) );
  XOR U4348 ( .A(b[5]), .B(a[101]), .Z(n4200) );
  NANDN U4349 ( .A(n5184), .B(n4200), .Z(n4160) );
  AND U4350 ( .A(n4161), .B(n4160), .Z(n4204) );
  AND U4351 ( .A(b[7]), .B(a[97]), .Z(n4203) );
  XNOR U4352 ( .A(n4204), .B(n4203), .Z(n4205) );
  XNOR U4353 ( .A(n4206), .B(n4205), .Z(n4211) );
  XOR U4354 ( .A(n4212), .B(n4211), .Z(n4186) );
  NANDN U4355 ( .A(n4163), .B(n4162), .Z(n4167) );
  NANDN U4356 ( .A(n4165), .B(n4164), .Z(n4166) );
  AND U4357 ( .A(n4167), .B(n4166), .Z(n4185) );
  XNOR U4358 ( .A(n4186), .B(n4185), .Z(n4187) );
  NANDN U4359 ( .A(n4169), .B(n4168), .Z(n4173) );
  NAND U4360 ( .A(n4171), .B(n4170), .Z(n4172) );
  NAND U4361 ( .A(n4173), .B(n4172), .Z(n4188) );
  XNOR U4362 ( .A(n4187), .B(n4188), .Z(n4179) );
  XNOR U4363 ( .A(n4180), .B(n4179), .Z(n4181) );
  XNOR U4364 ( .A(n4182), .B(n4181), .Z(n4215) );
  XNOR U4365 ( .A(sreg[225]), .B(n4215), .Z(n4217) );
  NANDN U4366 ( .A(sreg[224]), .B(n4174), .Z(n4178) );
  NAND U4367 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U4368 ( .A(n4178), .B(n4177), .Z(n4216) );
  XNOR U4369 ( .A(n4217), .B(n4216), .Z(c[225]) );
  NANDN U4370 ( .A(n4180), .B(n4179), .Z(n4184) );
  NANDN U4371 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U4372 ( .A(n4184), .B(n4183), .Z(n4223) );
  NANDN U4373 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4374 ( .A(n4188), .B(n4187), .Z(n4189) );
  AND U4375 ( .A(n4190), .B(n4189), .Z(n4221) );
  NANDN U4376 ( .A(n5274), .B(n4191), .Z(n4193) );
  XOR U4377 ( .A(b[7]), .B(a[100]), .Z(n4232) );
  NANDN U4378 ( .A(n5275), .B(n4232), .Z(n4192) );
  AND U4379 ( .A(n4193), .B(n4192), .Z(n4251) );
  NANDN U4380 ( .A(n5176), .B(n4194), .Z(n4196) );
  XOR U4381 ( .A(b[3]), .B(a[104]), .Z(n4235) );
  NANDN U4382 ( .A(n5177), .B(n4235), .Z(n4195) );
  NAND U4383 ( .A(n4196), .B(n4195), .Z(n4250) );
  XNOR U4384 ( .A(n4251), .B(n4250), .Z(n4253) );
  NAND U4385 ( .A(b[0]), .B(a[106]), .Z(n4197) );
  XNOR U4386 ( .A(b[1]), .B(n4197), .Z(n4199) );
  NANDN U4387 ( .A(b[0]), .B(a[105]), .Z(n4198) );
  NAND U4388 ( .A(n4199), .B(n4198), .Z(n4247) );
  NANDN U4389 ( .A(n5249), .B(n4200), .Z(n4202) );
  XOR U4390 ( .A(b[5]), .B(a[102]), .Z(n4241) );
  NANDN U4391 ( .A(n5184), .B(n4241), .Z(n4201) );
  AND U4392 ( .A(n4202), .B(n4201), .Z(n4245) );
  AND U4393 ( .A(b[7]), .B(a[98]), .Z(n4244) );
  XNOR U4394 ( .A(n4245), .B(n4244), .Z(n4246) );
  XNOR U4395 ( .A(n4247), .B(n4246), .Z(n4252) );
  XOR U4396 ( .A(n4253), .B(n4252), .Z(n4227) );
  NANDN U4397 ( .A(n4204), .B(n4203), .Z(n4208) );
  NANDN U4398 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U4399 ( .A(n4208), .B(n4207), .Z(n4226) );
  XNOR U4400 ( .A(n4227), .B(n4226), .Z(n4228) );
  NANDN U4401 ( .A(n4210), .B(n4209), .Z(n4214) );
  NAND U4402 ( .A(n4212), .B(n4211), .Z(n4213) );
  NAND U4403 ( .A(n4214), .B(n4213), .Z(n4229) );
  XNOR U4404 ( .A(n4228), .B(n4229), .Z(n4220) );
  XNOR U4405 ( .A(n4221), .B(n4220), .Z(n4222) );
  XNOR U4406 ( .A(n4223), .B(n4222), .Z(n4256) );
  XNOR U4407 ( .A(sreg[226]), .B(n4256), .Z(n4258) );
  NANDN U4408 ( .A(sreg[225]), .B(n4215), .Z(n4219) );
  NAND U4409 ( .A(n4217), .B(n4216), .Z(n4218) );
  NAND U4410 ( .A(n4219), .B(n4218), .Z(n4257) );
  XNOR U4411 ( .A(n4258), .B(n4257), .Z(c[226]) );
  NANDN U4412 ( .A(n4221), .B(n4220), .Z(n4225) );
  NANDN U4413 ( .A(n4223), .B(n4222), .Z(n4224) );
  AND U4414 ( .A(n4225), .B(n4224), .Z(n4264) );
  NANDN U4415 ( .A(n4227), .B(n4226), .Z(n4231) );
  NANDN U4416 ( .A(n4229), .B(n4228), .Z(n4230) );
  AND U4417 ( .A(n4231), .B(n4230), .Z(n4262) );
  NANDN U4418 ( .A(n5274), .B(n4232), .Z(n4234) );
  XOR U4419 ( .A(b[7]), .B(a[101]), .Z(n4273) );
  NANDN U4420 ( .A(n5275), .B(n4273), .Z(n4233) );
  AND U4421 ( .A(n4234), .B(n4233), .Z(n4292) );
  NANDN U4422 ( .A(n5176), .B(n4235), .Z(n4237) );
  XOR U4423 ( .A(b[3]), .B(a[105]), .Z(n4276) );
  NANDN U4424 ( .A(n5177), .B(n4276), .Z(n4236) );
  NAND U4425 ( .A(n4237), .B(n4236), .Z(n4291) );
  XNOR U4426 ( .A(n4292), .B(n4291), .Z(n4294) );
  NAND U4427 ( .A(b[0]), .B(a[107]), .Z(n4238) );
  XNOR U4428 ( .A(b[1]), .B(n4238), .Z(n4240) );
  NANDN U4429 ( .A(b[0]), .B(a[106]), .Z(n4239) );
  NAND U4430 ( .A(n4240), .B(n4239), .Z(n4288) );
  NANDN U4431 ( .A(n5249), .B(n4241), .Z(n4243) );
  XOR U4432 ( .A(b[5]), .B(a[103]), .Z(n4282) );
  NANDN U4433 ( .A(n5184), .B(n4282), .Z(n4242) );
  AND U4434 ( .A(n4243), .B(n4242), .Z(n4286) );
  AND U4435 ( .A(b[7]), .B(a[99]), .Z(n4285) );
  XNOR U4436 ( .A(n4286), .B(n4285), .Z(n4287) );
  XNOR U4437 ( .A(n4288), .B(n4287), .Z(n4293) );
  XOR U4438 ( .A(n4294), .B(n4293), .Z(n4268) );
  NANDN U4439 ( .A(n4245), .B(n4244), .Z(n4249) );
  NANDN U4440 ( .A(n4247), .B(n4246), .Z(n4248) );
  AND U4441 ( .A(n4249), .B(n4248), .Z(n4267) );
  XNOR U4442 ( .A(n4268), .B(n4267), .Z(n4269) );
  NANDN U4443 ( .A(n4251), .B(n4250), .Z(n4255) );
  NAND U4444 ( .A(n4253), .B(n4252), .Z(n4254) );
  NAND U4445 ( .A(n4255), .B(n4254), .Z(n4270) );
  XNOR U4446 ( .A(n4269), .B(n4270), .Z(n4261) );
  XNOR U4447 ( .A(n4262), .B(n4261), .Z(n4263) );
  XNOR U4448 ( .A(n4264), .B(n4263), .Z(n4297) );
  XNOR U4449 ( .A(sreg[227]), .B(n4297), .Z(n4299) );
  NANDN U4450 ( .A(sreg[226]), .B(n4256), .Z(n4260) );
  NAND U4451 ( .A(n4258), .B(n4257), .Z(n4259) );
  NAND U4452 ( .A(n4260), .B(n4259), .Z(n4298) );
  XNOR U4453 ( .A(n4299), .B(n4298), .Z(c[227]) );
  NANDN U4454 ( .A(n4262), .B(n4261), .Z(n4266) );
  NANDN U4455 ( .A(n4264), .B(n4263), .Z(n4265) );
  AND U4456 ( .A(n4266), .B(n4265), .Z(n4305) );
  NANDN U4457 ( .A(n4268), .B(n4267), .Z(n4272) );
  NANDN U4458 ( .A(n4270), .B(n4269), .Z(n4271) );
  AND U4459 ( .A(n4272), .B(n4271), .Z(n4303) );
  NANDN U4460 ( .A(n5274), .B(n4273), .Z(n4275) );
  XOR U4461 ( .A(b[7]), .B(a[102]), .Z(n4314) );
  NANDN U4462 ( .A(n5275), .B(n4314), .Z(n4274) );
  AND U4463 ( .A(n4275), .B(n4274), .Z(n4333) );
  NANDN U4464 ( .A(n5176), .B(n4276), .Z(n4278) );
  XOR U4465 ( .A(b[3]), .B(a[106]), .Z(n4317) );
  NANDN U4466 ( .A(n5177), .B(n4317), .Z(n4277) );
  NAND U4467 ( .A(n4278), .B(n4277), .Z(n4332) );
  XNOR U4468 ( .A(n4333), .B(n4332), .Z(n4335) );
  NAND U4469 ( .A(b[0]), .B(a[108]), .Z(n4279) );
  XNOR U4470 ( .A(b[1]), .B(n4279), .Z(n4281) );
  NANDN U4471 ( .A(b[0]), .B(a[107]), .Z(n4280) );
  NAND U4472 ( .A(n4281), .B(n4280), .Z(n4329) );
  NANDN U4473 ( .A(n5249), .B(n4282), .Z(n4284) );
  XOR U4474 ( .A(b[5]), .B(a[104]), .Z(n4323) );
  NANDN U4475 ( .A(n5184), .B(n4323), .Z(n4283) );
  AND U4476 ( .A(n4284), .B(n4283), .Z(n4327) );
  AND U4477 ( .A(b[7]), .B(a[100]), .Z(n4326) );
  XNOR U4478 ( .A(n4327), .B(n4326), .Z(n4328) );
  XNOR U4479 ( .A(n4329), .B(n4328), .Z(n4334) );
  XOR U4480 ( .A(n4335), .B(n4334), .Z(n4309) );
  NANDN U4481 ( .A(n4286), .B(n4285), .Z(n4290) );
  NANDN U4482 ( .A(n4288), .B(n4287), .Z(n4289) );
  AND U4483 ( .A(n4290), .B(n4289), .Z(n4308) );
  XNOR U4484 ( .A(n4309), .B(n4308), .Z(n4310) );
  NANDN U4485 ( .A(n4292), .B(n4291), .Z(n4296) );
  NAND U4486 ( .A(n4294), .B(n4293), .Z(n4295) );
  NAND U4487 ( .A(n4296), .B(n4295), .Z(n4311) );
  XNOR U4488 ( .A(n4310), .B(n4311), .Z(n4302) );
  XNOR U4489 ( .A(n4303), .B(n4302), .Z(n4304) );
  XNOR U4490 ( .A(n4305), .B(n4304), .Z(n4338) );
  XNOR U4491 ( .A(sreg[228]), .B(n4338), .Z(n4340) );
  NANDN U4492 ( .A(sreg[227]), .B(n4297), .Z(n4301) );
  NAND U4493 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U4494 ( .A(n4301), .B(n4300), .Z(n4339) );
  XNOR U4495 ( .A(n4340), .B(n4339), .Z(c[228]) );
  NANDN U4496 ( .A(n4303), .B(n4302), .Z(n4307) );
  NANDN U4497 ( .A(n4305), .B(n4304), .Z(n4306) );
  AND U4498 ( .A(n4307), .B(n4306), .Z(n4346) );
  NANDN U4499 ( .A(n4309), .B(n4308), .Z(n4313) );
  NANDN U4500 ( .A(n4311), .B(n4310), .Z(n4312) );
  AND U4501 ( .A(n4313), .B(n4312), .Z(n4344) );
  NANDN U4502 ( .A(n5274), .B(n4314), .Z(n4316) );
  XOR U4503 ( .A(b[7]), .B(a[103]), .Z(n4355) );
  NANDN U4504 ( .A(n5275), .B(n4355), .Z(n4315) );
  AND U4505 ( .A(n4316), .B(n4315), .Z(n4374) );
  NANDN U4506 ( .A(n5176), .B(n4317), .Z(n4319) );
  XOR U4507 ( .A(b[3]), .B(a[107]), .Z(n4358) );
  NANDN U4508 ( .A(n5177), .B(n4358), .Z(n4318) );
  NAND U4509 ( .A(n4319), .B(n4318), .Z(n4373) );
  XNOR U4510 ( .A(n4374), .B(n4373), .Z(n4376) );
  NAND U4511 ( .A(b[0]), .B(a[109]), .Z(n4320) );
  XNOR U4512 ( .A(b[1]), .B(n4320), .Z(n4322) );
  NANDN U4513 ( .A(b[0]), .B(a[108]), .Z(n4321) );
  NAND U4514 ( .A(n4322), .B(n4321), .Z(n4370) );
  NANDN U4515 ( .A(n5249), .B(n4323), .Z(n4325) );
  XOR U4516 ( .A(b[5]), .B(a[105]), .Z(n4361) );
  NANDN U4517 ( .A(n5184), .B(n4361), .Z(n4324) );
  AND U4518 ( .A(n4325), .B(n4324), .Z(n4368) );
  AND U4519 ( .A(b[7]), .B(a[101]), .Z(n4367) );
  XNOR U4520 ( .A(n4368), .B(n4367), .Z(n4369) );
  XNOR U4521 ( .A(n4370), .B(n4369), .Z(n4375) );
  XOR U4522 ( .A(n4376), .B(n4375), .Z(n4350) );
  NANDN U4523 ( .A(n4327), .B(n4326), .Z(n4331) );
  NANDN U4524 ( .A(n4329), .B(n4328), .Z(n4330) );
  AND U4525 ( .A(n4331), .B(n4330), .Z(n4349) );
  XNOR U4526 ( .A(n4350), .B(n4349), .Z(n4351) );
  NANDN U4527 ( .A(n4333), .B(n4332), .Z(n4337) );
  NAND U4528 ( .A(n4335), .B(n4334), .Z(n4336) );
  NAND U4529 ( .A(n4337), .B(n4336), .Z(n4352) );
  XNOR U4530 ( .A(n4351), .B(n4352), .Z(n4343) );
  XNOR U4531 ( .A(n4344), .B(n4343), .Z(n4345) );
  XNOR U4532 ( .A(n4346), .B(n4345), .Z(n4379) );
  XNOR U4533 ( .A(sreg[229]), .B(n4379), .Z(n4381) );
  NANDN U4534 ( .A(sreg[228]), .B(n4338), .Z(n4342) );
  NAND U4535 ( .A(n4340), .B(n4339), .Z(n4341) );
  NAND U4536 ( .A(n4342), .B(n4341), .Z(n4380) );
  XNOR U4537 ( .A(n4381), .B(n4380), .Z(c[229]) );
  NANDN U4538 ( .A(n4344), .B(n4343), .Z(n4348) );
  NANDN U4539 ( .A(n4346), .B(n4345), .Z(n4347) );
  AND U4540 ( .A(n4348), .B(n4347), .Z(n4387) );
  NANDN U4541 ( .A(n4350), .B(n4349), .Z(n4354) );
  NANDN U4542 ( .A(n4352), .B(n4351), .Z(n4353) );
  AND U4543 ( .A(n4354), .B(n4353), .Z(n4385) );
  NANDN U4544 ( .A(n5274), .B(n4355), .Z(n4357) );
  XOR U4545 ( .A(b[7]), .B(a[104]), .Z(n4396) );
  NANDN U4546 ( .A(n5275), .B(n4396), .Z(n4356) );
  AND U4547 ( .A(n4357), .B(n4356), .Z(n4415) );
  NANDN U4548 ( .A(n5176), .B(n4358), .Z(n4360) );
  XOR U4549 ( .A(b[3]), .B(a[108]), .Z(n4399) );
  NANDN U4550 ( .A(n5177), .B(n4399), .Z(n4359) );
  NAND U4551 ( .A(n4360), .B(n4359), .Z(n4414) );
  XNOR U4552 ( .A(n4415), .B(n4414), .Z(n4417) );
  NANDN U4553 ( .A(n5249), .B(n4361), .Z(n4363) );
  XOR U4554 ( .A(b[5]), .B(a[106]), .Z(n4405) );
  NANDN U4555 ( .A(n5184), .B(n4405), .Z(n4362) );
  AND U4556 ( .A(n4363), .B(n4362), .Z(n4409) );
  AND U4557 ( .A(b[7]), .B(a[102]), .Z(n4408) );
  XNOR U4558 ( .A(n4409), .B(n4408), .Z(n4410) );
  NAND U4559 ( .A(b[0]), .B(a[110]), .Z(n4364) );
  XNOR U4560 ( .A(b[1]), .B(n4364), .Z(n4366) );
  NANDN U4561 ( .A(b[0]), .B(a[109]), .Z(n4365) );
  NAND U4562 ( .A(n4366), .B(n4365), .Z(n4411) );
  XNOR U4563 ( .A(n4410), .B(n4411), .Z(n4416) );
  XOR U4564 ( .A(n4417), .B(n4416), .Z(n4391) );
  NANDN U4565 ( .A(n4368), .B(n4367), .Z(n4372) );
  NANDN U4566 ( .A(n4370), .B(n4369), .Z(n4371) );
  AND U4567 ( .A(n4372), .B(n4371), .Z(n4390) );
  XNOR U4568 ( .A(n4391), .B(n4390), .Z(n4392) );
  NANDN U4569 ( .A(n4374), .B(n4373), .Z(n4378) );
  NAND U4570 ( .A(n4376), .B(n4375), .Z(n4377) );
  NAND U4571 ( .A(n4378), .B(n4377), .Z(n4393) );
  XNOR U4572 ( .A(n4392), .B(n4393), .Z(n4384) );
  XNOR U4573 ( .A(n4385), .B(n4384), .Z(n4386) );
  XNOR U4574 ( .A(n4387), .B(n4386), .Z(n4420) );
  XNOR U4575 ( .A(sreg[230]), .B(n4420), .Z(n4422) );
  NANDN U4576 ( .A(sreg[229]), .B(n4379), .Z(n4383) );
  NAND U4577 ( .A(n4381), .B(n4380), .Z(n4382) );
  NAND U4578 ( .A(n4383), .B(n4382), .Z(n4421) );
  XNOR U4579 ( .A(n4422), .B(n4421), .Z(c[230]) );
  NANDN U4580 ( .A(n4385), .B(n4384), .Z(n4389) );
  NANDN U4581 ( .A(n4387), .B(n4386), .Z(n4388) );
  AND U4582 ( .A(n4389), .B(n4388), .Z(n4428) );
  NANDN U4583 ( .A(n4391), .B(n4390), .Z(n4395) );
  NANDN U4584 ( .A(n4393), .B(n4392), .Z(n4394) );
  AND U4585 ( .A(n4395), .B(n4394), .Z(n4426) );
  NANDN U4586 ( .A(n5274), .B(n4396), .Z(n4398) );
  XOR U4587 ( .A(b[7]), .B(a[105]), .Z(n4437) );
  NANDN U4588 ( .A(n5275), .B(n4437), .Z(n4397) );
  AND U4589 ( .A(n4398), .B(n4397), .Z(n4456) );
  NANDN U4590 ( .A(n5176), .B(n4399), .Z(n4401) );
  XOR U4591 ( .A(b[3]), .B(a[109]), .Z(n4440) );
  NANDN U4592 ( .A(n5177), .B(n4440), .Z(n4400) );
  NAND U4593 ( .A(n4401), .B(n4400), .Z(n4455) );
  XNOR U4594 ( .A(n4456), .B(n4455), .Z(n4458) );
  NAND U4595 ( .A(b[0]), .B(a[111]), .Z(n4402) );
  XNOR U4596 ( .A(b[1]), .B(n4402), .Z(n4404) );
  NANDN U4597 ( .A(b[0]), .B(a[110]), .Z(n4403) );
  NAND U4598 ( .A(n4404), .B(n4403), .Z(n4452) );
  NANDN U4599 ( .A(n5249), .B(n4405), .Z(n4407) );
  XOR U4600 ( .A(b[5]), .B(a[107]), .Z(n4446) );
  NANDN U4601 ( .A(n5184), .B(n4446), .Z(n4406) );
  AND U4602 ( .A(n4407), .B(n4406), .Z(n4450) );
  AND U4603 ( .A(b[7]), .B(a[103]), .Z(n4449) );
  XNOR U4604 ( .A(n4450), .B(n4449), .Z(n4451) );
  XNOR U4605 ( .A(n4452), .B(n4451), .Z(n4457) );
  XOR U4606 ( .A(n4458), .B(n4457), .Z(n4432) );
  NANDN U4607 ( .A(n4409), .B(n4408), .Z(n4413) );
  NANDN U4608 ( .A(n4411), .B(n4410), .Z(n4412) );
  AND U4609 ( .A(n4413), .B(n4412), .Z(n4431) );
  XNOR U4610 ( .A(n4432), .B(n4431), .Z(n4433) );
  NANDN U4611 ( .A(n4415), .B(n4414), .Z(n4419) );
  NAND U4612 ( .A(n4417), .B(n4416), .Z(n4418) );
  NAND U4613 ( .A(n4419), .B(n4418), .Z(n4434) );
  XNOR U4614 ( .A(n4433), .B(n4434), .Z(n4425) );
  XNOR U4615 ( .A(n4426), .B(n4425), .Z(n4427) );
  XNOR U4616 ( .A(n4428), .B(n4427), .Z(n4461) );
  XNOR U4617 ( .A(sreg[231]), .B(n4461), .Z(n4463) );
  NANDN U4618 ( .A(sreg[230]), .B(n4420), .Z(n4424) );
  NAND U4619 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U4620 ( .A(n4424), .B(n4423), .Z(n4462) );
  XNOR U4621 ( .A(n4463), .B(n4462), .Z(c[231]) );
  NANDN U4622 ( .A(n4426), .B(n4425), .Z(n4430) );
  NANDN U4623 ( .A(n4428), .B(n4427), .Z(n4429) );
  AND U4624 ( .A(n4430), .B(n4429), .Z(n4469) );
  NANDN U4625 ( .A(n4432), .B(n4431), .Z(n4436) );
  NANDN U4626 ( .A(n4434), .B(n4433), .Z(n4435) );
  AND U4627 ( .A(n4436), .B(n4435), .Z(n4467) );
  NANDN U4628 ( .A(n5274), .B(n4437), .Z(n4439) );
  XOR U4629 ( .A(b[7]), .B(a[106]), .Z(n4478) );
  NANDN U4630 ( .A(n5275), .B(n4478), .Z(n4438) );
  AND U4631 ( .A(n4439), .B(n4438), .Z(n4497) );
  NANDN U4632 ( .A(n5176), .B(n4440), .Z(n4442) );
  XOR U4633 ( .A(b[3]), .B(a[110]), .Z(n4481) );
  NANDN U4634 ( .A(n5177), .B(n4481), .Z(n4441) );
  NAND U4635 ( .A(n4442), .B(n4441), .Z(n4496) );
  XNOR U4636 ( .A(n4497), .B(n4496), .Z(n4499) );
  NAND U4637 ( .A(b[0]), .B(a[112]), .Z(n4443) );
  XNOR U4638 ( .A(b[1]), .B(n4443), .Z(n4445) );
  NANDN U4639 ( .A(b[0]), .B(a[111]), .Z(n4444) );
  NAND U4640 ( .A(n4445), .B(n4444), .Z(n4493) );
  NANDN U4641 ( .A(n5249), .B(n4446), .Z(n4448) );
  XOR U4642 ( .A(b[5]), .B(a[108]), .Z(n4484) );
  NANDN U4643 ( .A(n5184), .B(n4484), .Z(n4447) );
  AND U4644 ( .A(n4448), .B(n4447), .Z(n4491) );
  AND U4645 ( .A(b[7]), .B(a[104]), .Z(n4490) );
  XNOR U4646 ( .A(n4491), .B(n4490), .Z(n4492) );
  XNOR U4647 ( .A(n4493), .B(n4492), .Z(n4498) );
  XOR U4648 ( .A(n4499), .B(n4498), .Z(n4473) );
  NANDN U4649 ( .A(n4450), .B(n4449), .Z(n4454) );
  NANDN U4650 ( .A(n4452), .B(n4451), .Z(n4453) );
  AND U4651 ( .A(n4454), .B(n4453), .Z(n4472) );
  XNOR U4652 ( .A(n4473), .B(n4472), .Z(n4474) );
  NANDN U4653 ( .A(n4456), .B(n4455), .Z(n4460) );
  NAND U4654 ( .A(n4458), .B(n4457), .Z(n4459) );
  NAND U4655 ( .A(n4460), .B(n4459), .Z(n4475) );
  XNOR U4656 ( .A(n4474), .B(n4475), .Z(n4466) );
  XNOR U4657 ( .A(n4467), .B(n4466), .Z(n4468) );
  XNOR U4658 ( .A(n4469), .B(n4468), .Z(n4502) );
  XNOR U4659 ( .A(sreg[232]), .B(n4502), .Z(n4504) );
  NANDN U4660 ( .A(sreg[231]), .B(n4461), .Z(n4465) );
  NAND U4661 ( .A(n4463), .B(n4462), .Z(n4464) );
  NAND U4662 ( .A(n4465), .B(n4464), .Z(n4503) );
  XNOR U4663 ( .A(n4504), .B(n4503), .Z(c[232]) );
  NANDN U4664 ( .A(n4467), .B(n4466), .Z(n4471) );
  NANDN U4665 ( .A(n4469), .B(n4468), .Z(n4470) );
  AND U4666 ( .A(n4471), .B(n4470), .Z(n4510) );
  NANDN U4667 ( .A(n4473), .B(n4472), .Z(n4477) );
  NANDN U4668 ( .A(n4475), .B(n4474), .Z(n4476) );
  AND U4669 ( .A(n4477), .B(n4476), .Z(n4508) );
  NANDN U4670 ( .A(n5274), .B(n4478), .Z(n4480) );
  XOR U4671 ( .A(b[7]), .B(a[107]), .Z(n4519) );
  NANDN U4672 ( .A(n5275), .B(n4519), .Z(n4479) );
  AND U4673 ( .A(n4480), .B(n4479), .Z(n4538) );
  NANDN U4674 ( .A(n5176), .B(n4481), .Z(n4483) );
  XOR U4675 ( .A(b[3]), .B(a[111]), .Z(n4522) );
  NANDN U4676 ( .A(n5177), .B(n4522), .Z(n4482) );
  NAND U4677 ( .A(n4483), .B(n4482), .Z(n4537) );
  XNOR U4678 ( .A(n4538), .B(n4537), .Z(n4540) );
  NANDN U4679 ( .A(n5249), .B(n4484), .Z(n4486) );
  XOR U4680 ( .A(b[5]), .B(a[109]), .Z(n4528) );
  NANDN U4681 ( .A(n5184), .B(n4528), .Z(n4485) );
  AND U4682 ( .A(n4486), .B(n4485), .Z(n4532) );
  AND U4683 ( .A(b[7]), .B(a[105]), .Z(n4531) );
  XNOR U4684 ( .A(n4532), .B(n4531), .Z(n4533) );
  NAND U4685 ( .A(b[0]), .B(a[113]), .Z(n4487) );
  XNOR U4686 ( .A(b[1]), .B(n4487), .Z(n4489) );
  NANDN U4687 ( .A(b[0]), .B(a[112]), .Z(n4488) );
  NAND U4688 ( .A(n4489), .B(n4488), .Z(n4534) );
  XNOR U4689 ( .A(n4533), .B(n4534), .Z(n4539) );
  XOR U4690 ( .A(n4540), .B(n4539), .Z(n4514) );
  NANDN U4691 ( .A(n4491), .B(n4490), .Z(n4495) );
  NANDN U4692 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U4693 ( .A(n4495), .B(n4494), .Z(n4513) );
  XNOR U4694 ( .A(n4514), .B(n4513), .Z(n4515) );
  NANDN U4695 ( .A(n4497), .B(n4496), .Z(n4501) );
  NAND U4696 ( .A(n4499), .B(n4498), .Z(n4500) );
  NAND U4697 ( .A(n4501), .B(n4500), .Z(n4516) );
  XNOR U4698 ( .A(n4515), .B(n4516), .Z(n4507) );
  XNOR U4699 ( .A(n4508), .B(n4507), .Z(n4509) );
  XNOR U4700 ( .A(n4510), .B(n4509), .Z(n4543) );
  XNOR U4701 ( .A(sreg[233]), .B(n4543), .Z(n4545) );
  NANDN U4702 ( .A(sreg[232]), .B(n4502), .Z(n4506) );
  NAND U4703 ( .A(n4504), .B(n4503), .Z(n4505) );
  NAND U4704 ( .A(n4506), .B(n4505), .Z(n4544) );
  XNOR U4705 ( .A(n4545), .B(n4544), .Z(c[233]) );
  NANDN U4706 ( .A(n4508), .B(n4507), .Z(n4512) );
  NANDN U4707 ( .A(n4510), .B(n4509), .Z(n4511) );
  AND U4708 ( .A(n4512), .B(n4511), .Z(n4551) );
  NANDN U4709 ( .A(n4514), .B(n4513), .Z(n4518) );
  NANDN U4710 ( .A(n4516), .B(n4515), .Z(n4517) );
  AND U4711 ( .A(n4518), .B(n4517), .Z(n4549) );
  NANDN U4712 ( .A(n5274), .B(n4519), .Z(n4521) );
  XOR U4713 ( .A(b[7]), .B(a[108]), .Z(n4560) );
  NANDN U4714 ( .A(n5275), .B(n4560), .Z(n4520) );
  AND U4715 ( .A(n4521), .B(n4520), .Z(n4579) );
  NANDN U4716 ( .A(n5176), .B(n4522), .Z(n4524) );
  XOR U4717 ( .A(b[3]), .B(a[112]), .Z(n4563) );
  NANDN U4718 ( .A(n5177), .B(n4563), .Z(n4523) );
  NAND U4719 ( .A(n4524), .B(n4523), .Z(n4578) );
  XNOR U4720 ( .A(n4579), .B(n4578), .Z(n4581) );
  NAND U4721 ( .A(b[0]), .B(a[114]), .Z(n4525) );
  XNOR U4722 ( .A(b[1]), .B(n4525), .Z(n4527) );
  NANDN U4723 ( .A(b[0]), .B(a[113]), .Z(n4526) );
  NAND U4724 ( .A(n4527), .B(n4526), .Z(n4575) );
  NANDN U4725 ( .A(n5249), .B(n4528), .Z(n4530) );
  XOR U4726 ( .A(b[5]), .B(a[110]), .Z(n4569) );
  NANDN U4727 ( .A(n5184), .B(n4569), .Z(n4529) );
  AND U4728 ( .A(n4530), .B(n4529), .Z(n4573) );
  AND U4729 ( .A(b[7]), .B(a[106]), .Z(n4572) );
  XNOR U4730 ( .A(n4573), .B(n4572), .Z(n4574) );
  XNOR U4731 ( .A(n4575), .B(n4574), .Z(n4580) );
  XOR U4732 ( .A(n4581), .B(n4580), .Z(n4555) );
  NANDN U4733 ( .A(n4532), .B(n4531), .Z(n4536) );
  NANDN U4734 ( .A(n4534), .B(n4533), .Z(n4535) );
  AND U4735 ( .A(n4536), .B(n4535), .Z(n4554) );
  XNOR U4736 ( .A(n4555), .B(n4554), .Z(n4556) );
  NANDN U4737 ( .A(n4538), .B(n4537), .Z(n4542) );
  NAND U4738 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U4739 ( .A(n4542), .B(n4541), .Z(n4557) );
  XNOR U4740 ( .A(n4556), .B(n4557), .Z(n4548) );
  XNOR U4741 ( .A(n4549), .B(n4548), .Z(n4550) );
  XNOR U4742 ( .A(n4551), .B(n4550), .Z(n4584) );
  XNOR U4743 ( .A(sreg[234]), .B(n4584), .Z(n4586) );
  NANDN U4744 ( .A(sreg[233]), .B(n4543), .Z(n4547) );
  NAND U4745 ( .A(n4545), .B(n4544), .Z(n4546) );
  NAND U4746 ( .A(n4547), .B(n4546), .Z(n4585) );
  XNOR U4747 ( .A(n4586), .B(n4585), .Z(c[234]) );
  NANDN U4748 ( .A(n4549), .B(n4548), .Z(n4553) );
  NANDN U4749 ( .A(n4551), .B(n4550), .Z(n4552) );
  AND U4750 ( .A(n4553), .B(n4552), .Z(n4592) );
  NANDN U4751 ( .A(n4555), .B(n4554), .Z(n4559) );
  NANDN U4752 ( .A(n4557), .B(n4556), .Z(n4558) );
  AND U4753 ( .A(n4559), .B(n4558), .Z(n4590) );
  NANDN U4754 ( .A(n5274), .B(n4560), .Z(n4562) );
  XOR U4755 ( .A(b[7]), .B(a[109]), .Z(n4601) );
  NANDN U4756 ( .A(n5275), .B(n4601), .Z(n4561) );
  AND U4757 ( .A(n4562), .B(n4561), .Z(n4620) );
  NANDN U4758 ( .A(n5176), .B(n4563), .Z(n4565) );
  XOR U4759 ( .A(b[3]), .B(a[113]), .Z(n4604) );
  NANDN U4760 ( .A(n5177), .B(n4604), .Z(n4564) );
  NAND U4761 ( .A(n4565), .B(n4564), .Z(n4619) );
  XNOR U4762 ( .A(n4620), .B(n4619), .Z(n4622) );
  NAND U4763 ( .A(b[0]), .B(a[115]), .Z(n4566) );
  XNOR U4764 ( .A(b[1]), .B(n4566), .Z(n4568) );
  NANDN U4765 ( .A(b[0]), .B(a[114]), .Z(n4567) );
  NAND U4766 ( .A(n4568), .B(n4567), .Z(n4616) );
  NANDN U4767 ( .A(n5249), .B(n4569), .Z(n4571) );
  XOR U4768 ( .A(b[5]), .B(a[111]), .Z(n4607) );
  NANDN U4769 ( .A(n5184), .B(n4607), .Z(n4570) );
  AND U4770 ( .A(n4571), .B(n4570), .Z(n4614) );
  AND U4771 ( .A(b[7]), .B(a[107]), .Z(n4613) );
  XNOR U4772 ( .A(n4614), .B(n4613), .Z(n4615) );
  XNOR U4773 ( .A(n4616), .B(n4615), .Z(n4621) );
  XOR U4774 ( .A(n4622), .B(n4621), .Z(n4596) );
  NANDN U4775 ( .A(n4573), .B(n4572), .Z(n4577) );
  NANDN U4776 ( .A(n4575), .B(n4574), .Z(n4576) );
  AND U4777 ( .A(n4577), .B(n4576), .Z(n4595) );
  XNOR U4778 ( .A(n4596), .B(n4595), .Z(n4597) );
  NANDN U4779 ( .A(n4579), .B(n4578), .Z(n4583) );
  NAND U4780 ( .A(n4581), .B(n4580), .Z(n4582) );
  NAND U4781 ( .A(n4583), .B(n4582), .Z(n4598) );
  XNOR U4782 ( .A(n4597), .B(n4598), .Z(n4589) );
  XNOR U4783 ( .A(n4590), .B(n4589), .Z(n4591) );
  XNOR U4784 ( .A(n4592), .B(n4591), .Z(n4625) );
  XNOR U4785 ( .A(sreg[235]), .B(n4625), .Z(n4627) );
  NANDN U4786 ( .A(sreg[234]), .B(n4584), .Z(n4588) );
  NAND U4787 ( .A(n4586), .B(n4585), .Z(n4587) );
  NAND U4788 ( .A(n4588), .B(n4587), .Z(n4626) );
  XNOR U4789 ( .A(n4627), .B(n4626), .Z(c[235]) );
  NANDN U4790 ( .A(n4590), .B(n4589), .Z(n4594) );
  NANDN U4791 ( .A(n4592), .B(n4591), .Z(n4593) );
  AND U4792 ( .A(n4594), .B(n4593), .Z(n4633) );
  NANDN U4793 ( .A(n4596), .B(n4595), .Z(n4600) );
  NANDN U4794 ( .A(n4598), .B(n4597), .Z(n4599) );
  AND U4795 ( .A(n4600), .B(n4599), .Z(n4631) );
  NANDN U4796 ( .A(n5274), .B(n4601), .Z(n4603) );
  XOR U4797 ( .A(b[7]), .B(a[110]), .Z(n4642) );
  NANDN U4798 ( .A(n5275), .B(n4642), .Z(n4602) );
  AND U4799 ( .A(n4603), .B(n4602), .Z(n4661) );
  NANDN U4800 ( .A(n5176), .B(n4604), .Z(n4606) );
  XOR U4801 ( .A(b[3]), .B(a[114]), .Z(n4645) );
  NANDN U4802 ( .A(n5177), .B(n4645), .Z(n4605) );
  NAND U4803 ( .A(n4606), .B(n4605), .Z(n4660) );
  XNOR U4804 ( .A(n4661), .B(n4660), .Z(n4663) );
  NANDN U4805 ( .A(n5249), .B(n4607), .Z(n4609) );
  XOR U4806 ( .A(b[5]), .B(a[112]), .Z(n4651) );
  NANDN U4807 ( .A(n5184), .B(n4651), .Z(n4608) );
  AND U4808 ( .A(n4609), .B(n4608), .Z(n4655) );
  AND U4809 ( .A(b[7]), .B(a[108]), .Z(n4654) );
  XNOR U4810 ( .A(n4655), .B(n4654), .Z(n4656) );
  NAND U4811 ( .A(b[0]), .B(a[116]), .Z(n4610) );
  XNOR U4812 ( .A(b[1]), .B(n4610), .Z(n4612) );
  NANDN U4813 ( .A(b[0]), .B(a[115]), .Z(n4611) );
  NAND U4814 ( .A(n4612), .B(n4611), .Z(n4657) );
  XNOR U4815 ( .A(n4656), .B(n4657), .Z(n4662) );
  XOR U4816 ( .A(n4663), .B(n4662), .Z(n4637) );
  NANDN U4817 ( .A(n4614), .B(n4613), .Z(n4618) );
  NANDN U4818 ( .A(n4616), .B(n4615), .Z(n4617) );
  AND U4819 ( .A(n4618), .B(n4617), .Z(n4636) );
  XNOR U4820 ( .A(n4637), .B(n4636), .Z(n4638) );
  NANDN U4821 ( .A(n4620), .B(n4619), .Z(n4624) );
  NAND U4822 ( .A(n4622), .B(n4621), .Z(n4623) );
  NAND U4823 ( .A(n4624), .B(n4623), .Z(n4639) );
  XNOR U4824 ( .A(n4638), .B(n4639), .Z(n4630) );
  XNOR U4825 ( .A(n4631), .B(n4630), .Z(n4632) );
  XNOR U4826 ( .A(n4633), .B(n4632), .Z(n4666) );
  XNOR U4827 ( .A(sreg[236]), .B(n4666), .Z(n4668) );
  NANDN U4828 ( .A(sreg[235]), .B(n4625), .Z(n4629) );
  NAND U4829 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U4830 ( .A(n4629), .B(n4628), .Z(n4667) );
  XNOR U4831 ( .A(n4668), .B(n4667), .Z(c[236]) );
  NANDN U4832 ( .A(n4631), .B(n4630), .Z(n4635) );
  NANDN U4833 ( .A(n4633), .B(n4632), .Z(n4634) );
  AND U4834 ( .A(n4635), .B(n4634), .Z(n4674) );
  NANDN U4835 ( .A(n4637), .B(n4636), .Z(n4641) );
  NANDN U4836 ( .A(n4639), .B(n4638), .Z(n4640) );
  AND U4837 ( .A(n4641), .B(n4640), .Z(n4672) );
  NANDN U4838 ( .A(n5274), .B(n4642), .Z(n4644) );
  XOR U4839 ( .A(b[7]), .B(a[111]), .Z(n4683) );
  NANDN U4840 ( .A(n5275), .B(n4683), .Z(n4643) );
  AND U4841 ( .A(n4644), .B(n4643), .Z(n4702) );
  NANDN U4842 ( .A(n5176), .B(n4645), .Z(n4647) );
  XOR U4843 ( .A(b[3]), .B(a[115]), .Z(n4686) );
  NANDN U4844 ( .A(n5177), .B(n4686), .Z(n4646) );
  NAND U4845 ( .A(n4647), .B(n4646), .Z(n4701) );
  XNOR U4846 ( .A(n4702), .B(n4701), .Z(n4704) );
  NAND U4847 ( .A(b[0]), .B(a[117]), .Z(n4648) );
  XNOR U4848 ( .A(b[1]), .B(n4648), .Z(n4650) );
  NANDN U4849 ( .A(b[0]), .B(a[116]), .Z(n4649) );
  NAND U4850 ( .A(n4650), .B(n4649), .Z(n4698) );
  NANDN U4851 ( .A(n5249), .B(n4651), .Z(n4653) );
  XOR U4852 ( .A(b[5]), .B(a[113]), .Z(n4692) );
  NANDN U4853 ( .A(n5184), .B(n4692), .Z(n4652) );
  AND U4854 ( .A(n4653), .B(n4652), .Z(n4696) );
  AND U4855 ( .A(b[7]), .B(a[109]), .Z(n4695) );
  XNOR U4856 ( .A(n4696), .B(n4695), .Z(n4697) );
  XNOR U4857 ( .A(n4698), .B(n4697), .Z(n4703) );
  XOR U4858 ( .A(n4704), .B(n4703), .Z(n4678) );
  NANDN U4859 ( .A(n4655), .B(n4654), .Z(n4659) );
  NANDN U4860 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U4861 ( .A(n4659), .B(n4658), .Z(n4677) );
  XNOR U4862 ( .A(n4678), .B(n4677), .Z(n4679) );
  NANDN U4863 ( .A(n4661), .B(n4660), .Z(n4665) );
  NAND U4864 ( .A(n4663), .B(n4662), .Z(n4664) );
  NAND U4865 ( .A(n4665), .B(n4664), .Z(n4680) );
  XNOR U4866 ( .A(n4679), .B(n4680), .Z(n4671) );
  XNOR U4867 ( .A(n4672), .B(n4671), .Z(n4673) );
  XNOR U4868 ( .A(n4674), .B(n4673), .Z(n4707) );
  XNOR U4869 ( .A(sreg[237]), .B(n4707), .Z(n4709) );
  NANDN U4870 ( .A(sreg[236]), .B(n4666), .Z(n4670) );
  NAND U4871 ( .A(n4668), .B(n4667), .Z(n4669) );
  NAND U4872 ( .A(n4670), .B(n4669), .Z(n4708) );
  XNOR U4873 ( .A(n4709), .B(n4708), .Z(c[237]) );
  NANDN U4874 ( .A(n4672), .B(n4671), .Z(n4676) );
  NANDN U4875 ( .A(n4674), .B(n4673), .Z(n4675) );
  AND U4876 ( .A(n4676), .B(n4675), .Z(n4715) );
  NANDN U4877 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U4878 ( .A(n4680), .B(n4679), .Z(n4681) );
  AND U4879 ( .A(n4682), .B(n4681), .Z(n4713) );
  NANDN U4880 ( .A(n5274), .B(n4683), .Z(n4685) );
  XOR U4881 ( .A(b[7]), .B(a[112]), .Z(n4724) );
  NANDN U4882 ( .A(n5275), .B(n4724), .Z(n4684) );
  AND U4883 ( .A(n4685), .B(n4684), .Z(n4743) );
  NANDN U4884 ( .A(n5176), .B(n4686), .Z(n4688) );
  XOR U4885 ( .A(b[3]), .B(a[116]), .Z(n4727) );
  NANDN U4886 ( .A(n5177), .B(n4727), .Z(n4687) );
  NAND U4887 ( .A(n4688), .B(n4687), .Z(n4742) );
  XNOR U4888 ( .A(n4743), .B(n4742), .Z(n4745) );
  NAND U4889 ( .A(b[0]), .B(a[118]), .Z(n4689) );
  XNOR U4890 ( .A(b[1]), .B(n4689), .Z(n4691) );
  NANDN U4891 ( .A(b[0]), .B(a[117]), .Z(n4690) );
  NAND U4892 ( .A(n4691), .B(n4690), .Z(n4739) );
  NANDN U4893 ( .A(n5249), .B(n4692), .Z(n4694) );
  XOR U4894 ( .A(b[5]), .B(a[114]), .Z(n4733) );
  NANDN U4895 ( .A(n5184), .B(n4733), .Z(n4693) );
  AND U4896 ( .A(n4694), .B(n4693), .Z(n4737) );
  AND U4897 ( .A(b[7]), .B(a[110]), .Z(n4736) );
  XNOR U4898 ( .A(n4737), .B(n4736), .Z(n4738) );
  XNOR U4899 ( .A(n4739), .B(n4738), .Z(n4744) );
  XOR U4900 ( .A(n4745), .B(n4744), .Z(n4719) );
  NANDN U4901 ( .A(n4696), .B(n4695), .Z(n4700) );
  NANDN U4902 ( .A(n4698), .B(n4697), .Z(n4699) );
  AND U4903 ( .A(n4700), .B(n4699), .Z(n4718) );
  XNOR U4904 ( .A(n4719), .B(n4718), .Z(n4720) );
  NANDN U4905 ( .A(n4702), .B(n4701), .Z(n4706) );
  NAND U4906 ( .A(n4704), .B(n4703), .Z(n4705) );
  NAND U4907 ( .A(n4706), .B(n4705), .Z(n4721) );
  XNOR U4908 ( .A(n4720), .B(n4721), .Z(n4712) );
  XNOR U4909 ( .A(n4713), .B(n4712), .Z(n4714) );
  XNOR U4910 ( .A(n4715), .B(n4714), .Z(n4748) );
  XNOR U4911 ( .A(sreg[238]), .B(n4748), .Z(n4750) );
  NANDN U4912 ( .A(sreg[237]), .B(n4707), .Z(n4711) );
  NAND U4913 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U4914 ( .A(n4711), .B(n4710), .Z(n4749) );
  XNOR U4915 ( .A(n4750), .B(n4749), .Z(c[238]) );
  NANDN U4916 ( .A(n4713), .B(n4712), .Z(n4717) );
  NANDN U4917 ( .A(n4715), .B(n4714), .Z(n4716) );
  AND U4918 ( .A(n4717), .B(n4716), .Z(n4756) );
  NANDN U4919 ( .A(n4719), .B(n4718), .Z(n4723) );
  NANDN U4920 ( .A(n4721), .B(n4720), .Z(n4722) );
  AND U4921 ( .A(n4723), .B(n4722), .Z(n4754) );
  NANDN U4922 ( .A(n5274), .B(n4724), .Z(n4726) );
  XOR U4923 ( .A(b[7]), .B(a[113]), .Z(n4765) );
  NANDN U4924 ( .A(n5275), .B(n4765), .Z(n4725) );
  AND U4925 ( .A(n4726), .B(n4725), .Z(n4784) );
  NANDN U4926 ( .A(n5176), .B(n4727), .Z(n4729) );
  XOR U4927 ( .A(b[3]), .B(a[117]), .Z(n4768) );
  NANDN U4928 ( .A(n5177), .B(n4768), .Z(n4728) );
  NAND U4929 ( .A(n4729), .B(n4728), .Z(n4783) );
  XNOR U4930 ( .A(n4784), .B(n4783), .Z(n4786) );
  NAND U4931 ( .A(b[0]), .B(a[119]), .Z(n4730) );
  XNOR U4932 ( .A(b[1]), .B(n4730), .Z(n4732) );
  NANDN U4933 ( .A(b[0]), .B(a[118]), .Z(n4731) );
  NAND U4934 ( .A(n4732), .B(n4731), .Z(n4780) );
  NANDN U4935 ( .A(n5249), .B(n4733), .Z(n4735) );
  XOR U4936 ( .A(b[5]), .B(a[115]), .Z(n4774) );
  NANDN U4937 ( .A(n5184), .B(n4774), .Z(n4734) );
  AND U4938 ( .A(n4735), .B(n4734), .Z(n4778) );
  AND U4939 ( .A(b[7]), .B(a[111]), .Z(n4777) );
  XNOR U4940 ( .A(n4778), .B(n4777), .Z(n4779) );
  XNOR U4941 ( .A(n4780), .B(n4779), .Z(n4785) );
  XOR U4942 ( .A(n4786), .B(n4785), .Z(n4760) );
  NANDN U4943 ( .A(n4737), .B(n4736), .Z(n4741) );
  NANDN U4944 ( .A(n4739), .B(n4738), .Z(n4740) );
  AND U4945 ( .A(n4741), .B(n4740), .Z(n4759) );
  XNOR U4946 ( .A(n4760), .B(n4759), .Z(n4761) );
  NANDN U4947 ( .A(n4743), .B(n4742), .Z(n4747) );
  NAND U4948 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U4949 ( .A(n4747), .B(n4746), .Z(n4762) );
  XNOR U4950 ( .A(n4761), .B(n4762), .Z(n4753) );
  XNOR U4951 ( .A(n4754), .B(n4753), .Z(n4755) );
  XNOR U4952 ( .A(n4756), .B(n4755), .Z(n4789) );
  XNOR U4953 ( .A(sreg[239]), .B(n4789), .Z(n4791) );
  NANDN U4954 ( .A(sreg[238]), .B(n4748), .Z(n4752) );
  NAND U4955 ( .A(n4750), .B(n4749), .Z(n4751) );
  NAND U4956 ( .A(n4752), .B(n4751), .Z(n4790) );
  XNOR U4957 ( .A(n4791), .B(n4790), .Z(c[239]) );
  NANDN U4958 ( .A(n4754), .B(n4753), .Z(n4758) );
  NANDN U4959 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U4960 ( .A(n4758), .B(n4757), .Z(n4797) );
  NANDN U4961 ( .A(n4760), .B(n4759), .Z(n4764) );
  NANDN U4962 ( .A(n4762), .B(n4761), .Z(n4763) );
  AND U4963 ( .A(n4764), .B(n4763), .Z(n4795) );
  NANDN U4964 ( .A(n5274), .B(n4765), .Z(n4767) );
  XOR U4965 ( .A(b[7]), .B(a[114]), .Z(n4806) );
  NANDN U4966 ( .A(n5275), .B(n4806), .Z(n4766) );
  AND U4967 ( .A(n4767), .B(n4766), .Z(n4825) );
  NANDN U4968 ( .A(n5176), .B(n4768), .Z(n4770) );
  XOR U4969 ( .A(b[3]), .B(a[118]), .Z(n4809) );
  NANDN U4970 ( .A(n5177), .B(n4809), .Z(n4769) );
  NAND U4971 ( .A(n4770), .B(n4769), .Z(n4824) );
  XNOR U4972 ( .A(n4825), .B(n4824), .Z(n4827) );
  NAND U4973 ( .A(b[0]), .B(a[120]), .Z(n4771) );
  XNOR U4974 ( .A(b[1]), .B(n4771), .Z(n4773) );
  NANDN U4975 ( .A(b[0]), .B(a[119]), .Z(n4772) );
  NAND U4976 ( .A(n4773), .B(n4772), .Z(n4821) );
  NANDN U4977 ( .A(n5249), .B(n4774), .Z(n4776) );
  XOR U4978 ( .A(b[5]), .B(a[116]), .Z(n4815) );
  NANDN U4979 ( .A(n5184), .B(n4815), .Z(n4775) );
  AND U4980 ( .A(n4776), .B(n4775), .Z(n4819) );
  AND U4981 ( .A(b[7]), .B(a[112]), .Z(n4818) );
  XNOR U4982 ( .A(n4819), .B(n4818), .Z(n4820) );
  XNOR U4983 ( .A(n4821), .B(n4820), .Z(n4826) );
  XOR U4984 ( .A(n4827), .B(n4826), .Z(n4801) );
  NANDN U4985 ( .A(n4778), .B(n4777), .Z(n4782) );
  NANDN U4986 ( .A(n4780), .B(n4779), .Z(n4781) );
  AND U4987 ( .A(n4782), .B(n4781), .Z(n4800) );
  XNOR U4988 ( .A(n4801), .B(n4800), .Z(n4802) );
  NANDN U4989 ( .A(n4784), .B(n4783), .Z(n4788) );
  NAND U4990 ( .A(n4786), .B(n4785), .Z(n4787) );
  NAND U4991 ( .A(n4788), .B(n4787), .Z(n4803) );
  XNOR U4992 ( .A(n4802), .B(n4803), .Z(n4794) );
  XNOR U4993 ( .A(n4795), .B(n4794), .Z(n4796) );
  XNOR U4994 ( .A(n4797), .B(n4796), .Z(n4830) );
  XNOR U4995 ( .A(sreg[240]), .B(n4830), .Z(n4832) );
  NANDN U4996 ( .A(sreg[239]), .B(n4789), .Z(n4793) );
  NAND U4997 ( .A(n4791), .B(n4790), .Z(n4792) );
  NAND U4998 ( .A(n4793), .B(n4792), .Z(n4831) );
  XNOR U4999 ( .A(n4832), .B(n4831), .Z(c[240]) );
  NANDN U5000 ( .A(n4795), .B(n4794), .Z(n4799) );
  NANDN U5001 ( .A(n4797), .B(n4796), .Z(n4798) );
  AND U5002 ( .A(n4799), .B(n4798), .Z(n4838) );
  NANDN U5003 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U5004 ( .A(n4803), .B(n4802), .Z(n4804) );
  AND U5005 ( .A(n4805), .B(n4804), .Z(n4836) );
  NANDN U5006 ( .A(n5274), .B(n4806), .Z(n4808) );
  XOR U5007 ( .A(b[7]), .B(a[115]), .Z(n4847) );
  NANDN U5008 ( .A(n5275), .B(n4847), .Z(n4807) );
  AND U5009 ( .A(n4808), .B(n4807), .Z(n4866) );
  NANDN U5010 ( .A(n5176), .B(n4809), .Z(n4811) );
  XOR U5011 ( .A(b[3]), .B(a[119]), .Z(n4850) );
  NANDN U5012 ( .A(n5177), .B(n4850), .Z(n4810) );
  NAND U5013 ( .A(n4811), .B(n4810), .Z(n4865) );
  XNOR U5014 ( .A(n4866), .B(n4865), .Z(n4868) );
  NAND U5015 ( .A(b[0]), .B(a[121]), .Z(n4812) );
  XNOR U5016 ( .A(b[1]), .B(n4812), .Z(n4814) );
  NANDN U5017 ( .A(b[0]), .B(a[120]), .Z(n4813) );
  NAND U5018 ( .A(n4814), .B(n4813), .Z(n4862) );
  NANDN U5019 ( .A(n5249), .B(n4815), .Z(n4817) );
  XOR U5020 ( .A(b[5]), .B(a[117]), .Z(n4856) );
  NANDN U5021 ( .A(n5184), .B(n4856), .Z(n4816) );
  AND U5022 ( .A(n4817), .B(n4816), .Z(n4860) );
  AND U5023 ( .A(b[7]), .B(a[113]), .Z(n4859) );
  XNOR U5024 ( .A(n4860), .B(n4859), .Z(n4861) );
  XNOR U5025 ( .A(n4862), .B(n4861), .Z(n4867) );
  XOR U5026 ( .A(n4868), .B(n4867), .Z(n4842) );
  NANDN U5027 ( .A(n4819), .B(n4818), .Z(n4823) );
  NANDN U5028 ( .A(n4821), .B(n4820), .Z(n4822) );
  AND U5029 ( .A(n4823), .B(n4822), .Z(n4841) );
  XNOR U5030 ( .A(n4842), .B(n4841), .Z(n4843) );
  NANDN U5031 ( .A(n4825), .B(n4824), .Z(n4829) );
  NAND U5032 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5033 ( .A(n4829), .B(n4828), .Z(n4844) );
  XNOR U5034 ( .A(n4843), .B(n4844), .Z(n4835) );
  XNOR U5035 ( .A(n4836), .B(n4835), .Z(n4837) );
  XNOR U5036 ( .A(n4838), .B(n4837), .Z(n4871) );
  XNOR U5037 ( .A(sreg[241]), .B(n4871), .Z(n4873) );
  NANDN U5038 ( .A(sreg[240]), .B(n4830), .Z(n4834) );
  NAND U5039 ( .A(n4832), .B(n4831), .Z(n4833) );
  NAND U5040 ( .A(n4834), .B(n4833), .Z(n4872) );
  XNOR U5041 ( .A(n4873), .B(n4872), .Z(c[241]) );
  NANDN U5042 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U5043 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U5044 ( .A(n4840), .B(n4839), .Z(n4879) );
  NANDN U5045 ( .A(n4842), .B(n4841), .Z(n4846) );
  NANDN U5046 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U5047 ( .A(n4846), .B(n4845), .Z(n4877) );
  NANDN U5048 ( .A(n5274), .B(n4847), .Z(n4849) );
  XOR U5049 ( .A(b[7]), .B(a[116]), .Z(n4888) );
  NANDN U5050 ( .A(n5275), .B(n4888), .Z(n4848) );
  AND U5051 ( .A(n4849), .B(n4848), .Z(n4907) );
  NANDN U5052 ( .A(n5176), .B(n4850), .Z(n4852) );
  XOR U5053 ( .A(b[3]), .B(a[120]), .Z(n4891) );
  NANDN U5054 ( .A(n5177), .B(n4891), .Z(n4851) );
  NAND U5055 ( .A(n4852), .B(n4851), .Z(n4906) );
  XNOR U5056 ( .A(n4907), .B(n4906), .Z(n4909) );
  NAND U5057 ( .A(b[0]), .B(a[122]), .Z(n4853) );
  XNOR U5058 ( .A(b[1]), .B(n4853), .Z(n4855) );
  NANDN U5059 ( .A(b[0]), .B(a[121]), .Z(n4854) );
  NAND U5060 ( .A(n4855), .B(n4854), .Z(n4903) );
  NANDN U5061 ( .A(n5249), .B(n4856), .Z(n4858) );
  XOR U5062 ( .A(b[5]), .B(a[118]), .Z(n4897) );
  NANDN U5063 ( .A(n5184), .B(n4897), .Z(n4857) );
  AND U5064 ( .A(n4858), .B(n4857), .Z(n4901) );
  AND U5065 ( .A(b[7]), .B(a[114]), .Z(n4900) );
  XNOR U5066 ( .A(n4901), .B(n4900), .Z(n4902) );
  XNOR U5067 ( .A(n4903), .B(n4902), .Z(n4908) );
  XOR U5068 ( .A(n4909), .B(n4908), .Z(n4883) );
  NANDN U5069 ( .A(n4860), .B(n4859), .Z(n4864) );
  NANDN U5070 ( .A(n4862), .B(n4861), .Z(n4863) );
  AND U5071 ( .A(n4864), .B(n4863), .Z(n4882) );
  XNOR U5072 ( .A(n4883), .B(n4882), .Z(n4884) );
  NANDN U5073 ( .A(n4866), .B(n4865), .Z(n4870) );
  NAND U5074 ( .A(n4868), .B(n4867), .Z(n4869) );
  NAND U5075 ( .A(n4870), .B(n4869), .Z(n4885) );
  XNOR U5076 ( .A(n4884), .B(n4885), .Z(n4876) );
  XNOR U5077 ( .A(n4877), .B(n4876), .Z(n4878) );
  XNOR U5078 ( .A(n4879), .B(n4878), .Z(n4912) );
  XNOR U5079 ( .A(sreg[242]), .B(n4912), .Z(n4914) );
  NANDN U5080 ( .A(sreg[241]), .B(n4871), .Z(n4875) );
  NAND U5081 ( .A(n4873), .B(n4872), .Z(n4874) );
  NAND U5082 ( .A(n4875), .B(n4874), .Z(n4913) );
  XNOR U5083 ( .A(n4914), .B(n4913), .Z(c[242]) );
  NANDN U5084 ( .A(n4877), .B(n4876), .Z(n4881) );
  NANDN U5085 ( .A(n4879), .B(n4878), .Z(n4880) );
  AND U5086 ( .A(n4881), .B(n4880), .Z(n4920) );
  NANDN U5087 ( .A(n4883), .B(n4882), .Z(n4887) );
  NANDN U5088 ( .A(n4885), .B(n4884), .Z(n4886) );
  AND U5089 ( .A(n4887), .B(n4886), .Z(n4918) );
  NANDN U5090 ( .A(n5274), .B(n4888), .Z(n4890) );
  XOR U5091 ( .A(b[7]), .B(a[117]), .Z(n4929) );
  NANDN U5092 ( .A(n5275), .B(n4929), .Z(n4889) );
  AND U5093 ( .A(n4890), .B(n4889), .Z(n4948) );
  NANDN U5094 ( .A(n5176), .B(n4891), .Z(n4893) );
  XOR U5095 ( .A(b[3]), .B(a[121]), .Z(n4932) );
  NANDN U5096 ( .A(n5177), .B(n4932), .Z(n4892) );
  NAND U5097 ( .A(n4893), .B(n4892), .Z(n4947) );
  XNOR U5098 ( .A(n4948), .B(n4947), .Z(n4950) );
  NAND U5099 ( .A(b[0]), .B(a[123]), .Z(n4894) );
  XNOR U5100 ( .A(b[1]), .B(n4894), .Z(n4896) );
  NANDN U5101 ( .A(b[0]), .B(a[122]), .Z(n4895) );
  NAND U5102 ( .A(n4896), .B(n4895), .Z(n4944) );
  NANDN U5103 ( .A(n5249), .B(n4897), .Z(n4899) );
  XOR U5104 ( .A(b[5]), .B(a[119]), .Z(n4938) );
  NANDN U5105 ( .A(n5184), .B(n4938), .Z(n4898) );
  AND U5106 ( .A(n4899), .B(n4898), .Z(n4942) );
  AND U5107 ( .A(b[7]), .B(a[115]), .Z(n4941) );
  XNOR U5108 ( .A(n4942), .B(n4941), .Z(n4943) );
  XNOR U5109 ( .A(n4944), .B(n4943), .Z(n4949) );
  XOR U5110 ( .A(n4950), .B(n4949), .Z(n4924) );
  NANDN U5111 ( .A(n4901), .B(n4900), .Z(n4905) );
  NANDN U5112 ( .A(n4903), .B(n4902), .Z(n4904) );
  AND U5113 ( .A(n4905), .B(n4904), .Z(n4923) );
  XNOR U5114 ( .A(n4924), .B(n4923), .Z(n4925) );
  NANDN U5115 ( .A(n4907), .B(n4906), .Z(n4911) );
  NAND U5116 ( .A(n4909), .B(n4908), .Z(n4910) );
  NAND U5117 ( .A(n4911), .B(n4910), .Z(n4926) );
  XNOR U5118 ( .A(n4925), .B(n4926), .Z(n4917) );
  XNOR U5119 ( .A(n4918), .B(n4917), .Z(n4919) );
  XNOR U5120 ( .A(n4920), .B(n4919), .Z(n4953) );
  XNOR U5121 ( .A(sreg[243]), .B(n4953), .Z(n4955) );
  NANDN U5122 ( .A(sreg[242]), .B(n4912), .Z(n4916) );
  NAND U5123 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U5124 ( .A(n4916), .B(n4915), .Z(n4954) );
  XNOR U5125 ( .A(n4955), .B(n4954), .Z(c[243]) );
  NANDN U5126 ( .A(n4918), .B(n4917), .Z(n4922) );
  NANDN U5127 ( .A(n4920), .B(n4919), .Z(n4921) );
  AND U5128 ( .A(n4922), .B(n4921), .Z(n4961) );
  NANDN U5129 ( .A(n4924), .B(n4923), .Z(n4928) );
  NANDN U5130 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U5131 ( .A(n4928), .B(n4927), .Z(n4959) );
  NANDN U5132 ( .A(n5274), .B(n4929), .Z(n4931) );
  XOR U5133 ( .A(b[7]), .B(a[118]), .Z(n4970) );
  NANDN U5134 ( .A(n5275), .B(n4970), .Z(n4930) );
  AND U5135 ( .A(n4931), .B(n4930), .Z(n4989) );
  NANDN U5136 ( .A(n5176), .B(n4932), .Z(n4934) );
  XOR U5137 ( .A(b[3]), .B(a[122]), .Z(n4973) );
  NANDN U5138 ( .A(n5177), .B(n4973), .Z(n4933) );
  NAND U5139 ( .A(n4934), .B(n4933), .Z(n4988) );
  XNOR U5140 ( .A(n4989), .B(n4988), .Z(n4991) );
  NAND U5141 ( .A(b[0]), .B(a[124]), .Z(n4935) );
  XNOR U5142 ( .A(b[1]), .B(n4935), .Z(n4937) );
  NANDN U5143 ( .A(b[0]), .B(a[123]), .Z(n4936) );
  NAND U5144 ( .A(n4937), .B(n4936), .Z(n4985) );
  NANDN U5145 ( .A(n5249), .B(n4938), .Z(n4940) );
  XOR U5146 ( .A(b[5]), .B(a[120]), .Z(n4979) );
  NANDN U5147 ( .A(n5184), .B(n4979), .Z(n4939) );
  AND U5148 ( .A(n4940), .B(n4939), .Z(n4983) );
  AND U5149 ( .A(b[7]), .B(a[116]), .Z(n4982) );
  XNOR U5150 ( .A(n4983), .B(n4982), .Z(n4984) );
  XNOR U5151 ( .A(n4985), .B(n4984), .Z(n4990) );
  XOR U5152 ( .A(n4991), .B(n4990), .Z(n4965) );
  NANDN U5153 ( .A(n4942), .B(n4941), .Z(n4946) );
  NANDN U5154 ( .A(n4944), .B(n4943), .Z(n4945) );
  AND U5155 ( .A(n4946), .B(n4945), .Z(n4964) );
  XNOR U5156 ( .A(n4965), .B(n4964), .Z(n4966) );
  NANDN U5157 ( .A(n4948), .B(n4947), .Z(n4952) );
  NAND U5158 ( .A(n4950), .B(n4949), .Z(n4951) );
  NAND U5159 ( .A(n4952), .B(n4951), .Z(n4967) );
  XNOR U5160 ( .A(n4966), .B(n4967), .Z(n4958) );
  XNOR U5161 ( .A(n4959), .B(n4958), .Z(n4960) );
  XNOR U5162 ( .A(n4961), .B(n4960), .Z(n4994) );
  XNOR U5163 ( .A(sreg[244]), .B(n4994), .Z(n4996) );
  NANDN U5164 ( .A(sreg[243]), .B(n4953), .Z(n4957) );
  NAND U5165 ( .A(n4955), .B(n4954), .Z(n4956) );
  NAND U5166 ( .A(n4957), .B(n4956), .Z(n4995) );
  XNOR U5167 ( .A(n4996), .B(n4995), .Z(c[244]) );
  NANDN U5168 ( .A(n4959), .B(n4958), .Z(n4963) );
  NANDN U5169 ( .A(n4961), .B(n4960), .Z(n4962) );
  AND U5170 ( .A(n4963), .B(n4962), .Z(n5002) );
  NANDN U5171 ( .A(n4965), .B(n4964), .Z(n4969) );
  NANDN U5172 ( .A(n4967), .B(n4966), .Z(n4968) );
  AND U5173 ( .A(n4969), .B(n4968), .Z(n5000) );
  NANDN U5174 ( .A(n5274), .B(n4970), .Z(n4972) );
  XOR U5175 ( .A(b[7]), .B(a[119]), .Z(n5011) );
  NANDN U5176 ( .A(n5275), .B(n5011), .Z(n4971) );
  AND U5177 ( .A(n4972), .B(n4971), .Z(n5030) );
  NANDN U5178 ( .A(n5176), .B(n4973), .Z(n4975) );
  XOR U5179 ( .A(b[3]), .B(a[123]), .Z(n5014) );
  NANDN U5180 ( .A(n5177), .B(n5014), .Z(n4974) );
  NAND U5181 ( .A(n4975), .B(n4974), .Z(n5029) );
  XNOR U5182 ( .A(n5030), .B(n5029), .Z(n5032) );
  NAND U5183 ( .A(b[0]), .B(a[125]), .Z(n4976) );
  XNOR U5184 ( .A(b[1]), .B(n4976), .Z(n4978) );
  NANDN U5185 ( .A(b[0]), .B(a[124]), .Z(n4977) );
  NAND U5186 ( .A(n4978), .B(n4977), .Z(n5026) );
  NANDN U5187 ( .A(n5249), .B(n4979), .Z(n4981) );
  XOR U5188 ( .A(b[5]), .B(a[121]), .Z(n5020) );
  NANDN U5189 ( .A(n5184), .B(n5020), .Z(n4980) );
  AND U5190 ( .A(n4981), .B(n4980), .Z(n5024) );
  AND U5191 ( .A(b[7]), .B(a[117]), .Z(n5023) );
  XNOR U5192 ( .A(n5024), .B(n5023), .Z(n5025) );
  XNOR U5193 ( .A(n5026), .B(n5025), .Z(n5031) );
  XOR U5194 ( .A(n5032), .B(n5031), .Z(n5006) );
  NANDN U5195 ( .A(n4983), .B(n4982), .Z(n4987) );
  NANDN U5196 ( .A(n4985), .B(n4984), .Z(n4986) );
  AND U5197 ( .A(n4987), .B(n4986), .Z(n5005) );
  XNOR U5198 ( .A(n5006), .B(n5005), .Z(n5007) );
  NANDN U5199 ( .A(n4989), .B(n4988), .Z(n4993) );
  NAND U5200 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U5201 ( .A(n4993), .B(n4992), .Z(n5008) );
  XNOR U5202 ( .A(n5007), .B(n5008), .Z(n4999) );
  XNOR U5203 ( .A(n5000), .B(n4999), .Z(n5001) );
  XNOR U5204 ( .A(n5002), .B(n5001), .Z(n5035) );
  XNOR U5205 ( .A(sreg[245]), .B(n5035), .Z(n5037) );
  NANDN U5206 ( .A(sreg[244]), .B(n4994), .Z(n4998) );
  NAND U5207 ( .A(n4996), .B(n4995), .Z(n4997) );
  NAND U5208 ( .A(n4998), .B(n4997), .Z(n5036) );
  XNOR U5209 ( .A(n5037), .B(n5036), .Z(c[245]) );
  NANDN U5210 ( .A(n5000), .B(n4999), .Z(n5004) );
  NANDN U5211 ( .A(n5002), .B(n5001), .Z(n5003) );
  AND U5212 ( .A(n5004), .B(n5003), .Z(n5043) );
  NANDN U5213 ( .A(n5006), .B(n5005), .Z(n5010) );
  NANDN U5214 ( .A(n5008), .B(n5007), .Z(n5009) );
  AND U5215 ( .A(n5010), .B(n5009), .Z(n5041) );
  NANDN U5216 ( .A(n5274), .B(n5011), .Z(n5013) );
  XOR U5217 ( .A(b[7]), .B(a[120]), .Z(n5064) );
  NANDN U5218 ( .A(n5275), .B(n5064), .Z(n5012) );
  AND U5219 ( .A(n5013), .B(n5012), .Z(n5053) );
  NANDN U5220 ( .A(n5176), .B(n5014), .Z(n5016) );
  XOR U5221 ( .A(b[3]), .B(a[124]), .Z(n5067) );
  NANDN U5222 ( .A(n5177), .B(n5067), .Z(n5015) );
  NAND U5223 ( .A(n5016), .B(n5015), .Z(n5052) );
  NAND U5224 ( .A(b[0]), .B(a[126]), .Z(n5017) );
  XNOR U5225 ( .A(b[1]), .B(n5017), .Z(n5019) );
  NANDN U5226 ( .A(b[0]), .B(a[125]), .Z(n5018) );
  NAND U5227 ( .A(n5019), .B(n5018), .Z(n5061) );
  NANDN U5228 ( .A(n5249), .B(n5020), .Z(n5022) );
  XOR U5229 ( .A(b[5]), .B(a[122]), .Z(n5070) );
  NANDN U5230 ( .A(n5184), .B(n5070), .Z(n5021) );
  AND U5231 ( .A(n5022), .B(n5021), .Z(n5059) );
  AND U5232 ( .A(b[7]), .B(a[118]), .Z(n5058) );
  XNOR U5233 ( .A(n5061), .B(n5060), .Z(n5054) );
  XOR U5234 ( .A(n5055), .B(n5054), .Z(n5047) );
  NANDN U5235 ( .A(n5024), .B(n5023), .Z(n5028) );
  NANDN U5236 ( .A(n5026), .B(n5025), .Z(n5027) );
  AND U5237 ( .A(n5028), .B(n5027), .Z(n5046) );
  NANDN U5238 ( .A(n5030), .B(n5029), .Z(n5034) );
  NAND U5239 ( .A(n5032), .B(n5031), .Z(n5033) );
  NAND U5240 ( .A(n5034), .B(n5033), .Z(n5049) );
  XNOR U5241 ( .A(n5041), .B(n5040), .Z(n5042) );
  XNOR U5242 ( .A(n5043), .B(n5042), .Z(n5076) );
  XNOR U5243 ( .A(sreg[246]), .B(n5076), .Z(n5078) );
  NANDN U5244 ( .A(sreg[245]), .B(n5035), .Z(n5039) );
  NAND U5245 ( .A(n5037), .B(n5036), .Z(n5038) );
  NAND U5246 ( .A(n5039), .B(n5038), .Z(n5077) );
  XNOR U5247 ( .A(n5078), .B(n5077), .Z(c[246]) );
  NANDN U5248 ( .A(n5041), .B(n5040), .Z(n5045) );
  NANDN U5249 ( .A(n5043), .B(n5042), .Z(n5044) );
  AND U5250 ( .A(n5045), .B(n5044), .Z(n5089) );
  NANDN U5251 ( .A(n5047), .B(n5046), .Z(n5051) );
  NANDN U5252 ( .A(n5049), .B(n5048), .Z(n5050) );
  AND U5253 ( .A(n5051), .B(n5050), .Z(n5087) );
  NANDN U5254 ( .A(n5053), .B(n5052), .Z(n5057) );
  NAND U5255 ( .A(n5055), .B(n5054), .Z(n5056) );
  AND U5256 ( .A(n5057), .B(n5056), .Z(n5116) );
  NANDN U5257 ( .A(n5059), .B(n5058), .Z(n5063) );
  NANDN U5258 ( .A(n5061), .B(n5060), .Z(n5062) );
  AND U5259 ( .A(n5063), .B(n5062), .Z(n5114) );
  NANDN U5260 ( .A(n5274), .B(n5064), .Z(n5066) );
  XOR U5261 ( .A(b[7]), .B(a[121]), .Z(n5104) );
  NANDN U5262 ( .A(n5275), .B(n5104), .Z(n5065) );
  AND U5263 ( .A(n5066), .B(n5065), .Z(n5095) );
  NANDN U5264 ( .A(n5176), .B(n5067), .Z(n5069) );
  XOR U5265 ( .A(b[3]), .B(a[125]), .Z(n5107) );
  NANDN U5266 ( .A(n5177), .B(n5107), .Z(n5068) );
  AND U5267 ( .A(n5069), .B(n5068), .Z(n5093) );
  NANDN U5268 ( .A(n5249), .B(n5070), .Z(n5072) );
  XOR U5269 ( .A(b[5]), .B(a[123]), .Z(n5110) );
  NANDN U5270 ( .A(n5184), .B(n5110), .Z(n5071) );
  AND U5271 ( .A(n5072), .B(n5071), .Z(n5099) );
  AND U5272 ( .A(b[7]), .B(a[119]), .Z(n5098) );
  NAND U5273 ( .A(b[0]), .B(a[127]), .Z(n5073) );
  XNOR U5274 ( .A(b[1]), .B(n5073), .Z(n5075) );
  NANDN U5275 ( .A(b[0]), .B(a[126]), .Z(n5074) );
  NAND U5276 ( .A(n5075), .B(n5074), .Z(n5101) );
  XNOR U5277 ( .A(n5100), .B(n5101), .Z(n5092) );
  XOR U5278 ( .A(n5116), .B(n5115), .Z(n5086) );
  XNOR U5279 ( .A(sreg[247]), .B(n5081), .Z(n5083) );
  NANDN U5280 ( .A(sreg[246]), .B(n5076), .Z(n5080) );
  NAND U5281 ( .A(n5078), .B(n5077), .Z(n5079) );
  NAND U5282 ( .A(n5080), .B(n5079), .Z(n5082) );
  XNOR U5283 ( .A(n5083), .B(n5082), .Z(c[247]) );
  NANDN U5284 ( .A(sreg[247]), .B(n5081), .Z(n5085) );
  NAND U5285 ( .A(n5083), .B(n5082), .Z(n5084) );
  AND U5286 ( .A(n5085), .B(n5084), .Z(n5120) );
  NANDN U5287 ( .A(n5087), .B(n5086), .Z(n5091) );
  NANDN U5288 ( .A(n5089), .B(n5088), .Z(n5090) );
  AND U5289 ( .A(n5091), .B(n5090), .Z(n5124) );
  NANDN U5290 ( .A(n5093), .B(n5092), .Z(n5097) );
  NANDN U5291 ( .A(n5095), .B(n5094), .Z(n5096) );
  AND U5292 ( .A(n5097), .B(n5096), .Z(n5153) );
  NANDN U5293 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U5294 ( .A(n5101), .B(n5100), .Z(n5102) );
  AND U5295 ( .A(n5103), .B(n5102), .Z(n5151) );
  NANDN U5296 ( .A(n5274), .B(n5104), .Z(n5106) );
  XOR U5297 ( .A(b[7]), .B(a[122]), .Z(n5127) );
  NANDN U5298 ( .A(n5275), .B(n5127), .Z(n5105) );
  AND U5299 ( .A(n5106), .B(n5105), .Z(n5147) );
  NANDN U5300 ( .A(n5176), .B(n5107), .Z(n5109) );
  XOR U5301 ( .A(a[126]), .B(b[3]), .Z(n5133) );
  NANDN U5302 ( .A(n5177), .B(n5133), .Z(n5108) );
  AND U5303 ( .A(n5109), .B(n5108), .Z(n5145) );
  NANDN U5304 ( .A(n5249), .B(n5110), .Z(n5112) );
  XOR U5305 ( .A(b[5]), .B(a[124]), .Z(n5130) );
  NANDN U5306 ( .A(n5184), .B(n5130), .Z(n5111) );
  AND U5307 ( .A(n5112), .B(n5111), .Z(n5139) );
  AND U5308 ( .A(b[7]), .B(a[120]), .Z(n5138) );
  NANDN U5309 ( .A(n5114), .B(n5113), .Z(n5118) );
  NANDN U5310 ( .A(n5116), .B(n5115), .Z(n5117) );
  AND U5311 ( .A(n5118), .B(n5117), .Z(n5122) );
  XOR U5312 ( .A(n5121), .B(n5122), .Z(n5123) );
  XOR U5313 ( .A(n5124), .B(n5123), .Z(n5119) );
  XOR U5314 ( .A(n5120), .B(n5119), .Z(c[248]) );
  AND U5315 ( .A(n5120), .B(n5119), .Z(n5157) );
  NAND U5316 ( .A(n5122), .B(n5121), .Z(n5126) );
  NANDN U5317 ( .A(n5124), .B(n5123), .Z(n5125) );
  AND U5318 ( .A(n5126), .B(n5125), .Z(n5161) );
  NANDN U5319 ( .A(n5274), .B(n5127), .Z(n5129) );
  XOR U5320 ( .A(b[7]), .B(a[123]), .Z(n5180) );
  NANDN U5321 ( .A(n5275), .B(n5180), .Z(n5128) );
  AND U5322 ( .A(n5129), .B(n5128), .Z(n5189) );
  NAND U5323 ( .A(b[7]), .B(a[121]), .Z(n5243) );
  NANDN U5324 ( .A(n5249), .B(n5130), .Z(n5132) );
  XOR U5325 ( .A(b[5]), .B(a[125]), .Z(n5183) );
  NANDN U5326 ( .A(n5184), .B(n5183), .Z(n5131) );
  NAND U5327 ( .A(n5132), .B(n5131), .Z(n5187) );
  XOR U5328 ( .A(n5243), .B(n5187), .Z(n5188) );
  NAND U5329 ( .A(n5134), .B(n5133), .Z(n5137) );
  XOR U5330 ( .A(a[127]), .B(b[3]), .Z(n5175) );
  NAND U5331 ( .A(n5135), .B(n5175), .Z(n5136) );
  NAND U5332 ( .A(n5137), .B(n5136), .Z(n5170) );
  XOR U5333 ( .A(n5171), .B(n5172), .Z(n5164) );
  NANDN U5334 ( .A(n5139), .B(n5138), .Z(n5143) );
  NANDN U5335 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5336 ( .A(n5143), .B(n5142), .Z(n5165) );
  NANDN U5337 ( .A(n5145), .B(n5144), .Z(n5149) );
  NANDN U5338 ( .A(n5147), .B(n5146), .Z(n5148) );
  NAND U5339 ( .A(n5149), .B(n5148), .Z(n5167) );
  NANDN U5340 ( .A(n5151), .B(n5150), .Z(n5155) );
  NANDN U5341 ( .A(n5153), .B(n5152), .Z(n5154) );
  NAND U5342 ( .A(n5155), .B(n5154), .Z(n5159) );
  XOR U5343 ( .A(n5161), .B(n5160), .Z(n5156) );
  XOR U5344 ( .A(n5157), .B(n5156), .Z(c[249]) );
  AND U5345 ( .A(n5157), .B(n5156), .Z(n5193) );
  NANDN U5346 ( .A(n5159), .B(n5158), .Z(n5163) );
  NANDN U5347 ( .A(n5161), .B(n5160), .Z(n5162) );
  AND U5348 ( .A(n5163), .B(n5162), .Z(n5197) );
  NANDN U5349 ( .A(n5165), .B(n5164), .Z(n5169) );
  NANDN U5350 ( .A(n5167), .B(n5166), .Z(n5168) );
  AND U5351 ( .A(n5169), .B(n5168), .Z(n5195) );
  NANDN U5352 ( .A(n5170), .B(b[1]), .Z(n5174) );
  NAND U5353 ( .A(n5172), .B(n5171), .Z(n5173) );
  AND U5354 ( .A(n5174), .B(n5173), .Z(n5203) );
  NANDN U5355 ( .A(n5176), .B(n5175), .Z(n5179) );
  NANDN U5356 ( .A(n5177), .B(b[3]), .Z(n5178) );
  AND U5357 ( .A(n5179), .B(n5178), .Z(n5221) );
  AND U5358 ( .A(b[7]), .B(a[122]), .Z(n5220) );
  XOR U5359 ( .A(n5243), .B(n5222), .Z(n5209) );
  NANDN U5360 ( .A(n5274), .B(n5180), .Z(n5182) );
  XOR U5361 ( .A(b[7]), .B(a[124]), .Z(n5212) );
  NANDN U5362 ( .A(n5275), .B(n5212), .Z(n5181) );
  AND U5363 ( .A(n5182), .B(n5181), .Z(n5207) );
  NANDN U5364 ( .A(n5249), .B(n5183), .Z(n5186) );
  XOR U5365 ( .A(b[5]), .B(a[126]), .Z(n5215) );
  NANDN U5366 ( .A(n5184), .B(n5215), .Z(n5185) );
  NAND U5367 ( .A(n5186), .B(n5185), .Z(n5206) );
  XOR U5368 ( .A(n5209), .B(n5208), .Z(n5201) );
  IV U5369 ( .A(n5243), .Z(n5223) );
  NANDN U5370 ( .A(n5223), .B(n5187), .Z(n5191) );
  NANDN U5371 ( .A(n5189), .B(n5188), .Z(n5190) );
  AND U5372 ( .A(n5191), .B(n5190), .Z(n5200) );
  XOR U5373 ( .A(n5197), .B(n5196), .Z(n5192) );
  XOR U5374 ( .A(n5193), .B(n5192), .Z(c[250]) );
  AND U5375 ( .A(n5193), .B(n5192), .Z(n5227) );
  NANDN U5376 ( .A(n5195), .B(n5194), .Z(n5199) );
  NANDN U5377 ( .A(n5197), .B(n5196), .Z(n5198) );
  AND U5378 ( .A(n5199), .B(n5198), .Z(n5231) );
  NANDN U5379 ( .A(n5201), .B(n5200), .Z(n5205) );
  NANDN U5380 ( .A(n5203), .B(n5202), .Z(n5204) );
  AND U5381 ( .A(n5205), .B(n5204), .Z(n5229) );
  NANDN U5382 ( .A(n5207), .B(n5206), .Z(n5211) );
  NAND U5383 ( .A(n5209), .B(n5208), .Z(n5210) );
  AND U5384 ( .A(n5211), .B(n5210), .Z(n5257) );
  NANDN U5385 ( .A(n5274), .B(n5212), .Z(n5214) );
  XOR U5386 ( .A(b[7]), .B(a[125]), .Z(n5246) );
  NANDN U5387 ( .A(n5275), .B(n5246), .Z(n5213) );
  AND U5388 ( .A(n5214), .B(n5213), .Z(n5235) );
  XOR U5389 ( .A(a[127]), .B(b[5]), .Z(n5250) );
  NAND U5390 ( .A(n5251), .B(n5250), .Z(n5218) );
  NAND U5391 ( .A(n5216), .B(n5215), .Z(n5217) );
  NAND U5392 ( .A(n5218), .B(n5217), .Z(n5234) );
  AND U5393 ( .A(b[7]), .B(a[123]), .Z(n5240) );
  XOR U5394 ( .A(n5219), .B(n5240), .Z(n5242) );
  XOR U5395 ( .A(n5223), .B(n5242), .Z(n5236) );
  XOR U5396 ( .A(n5237), .B(n5236), .Z(n5255) );
  NANDN U5397 ( .A(n5221), .B(n5220), .Z(n5225) );
  NANDN U5398 ( .A(n5223), .B(n5222), .Z(n5224) );
  AND U5399 ( .A(n5225), .B(n5224), .Z(n5254) );
  XOR U5400 ( .A(n5257), .B(n5256), .Z(n5228) );
  XOR U5401 ( .A(n5231), .B(n5230), .Z(n5226) );
  XOR U5402 ( .A(n5227), .B(n5226), .Z(c[251]) );
  AND U5403 ( .A(n5227), .B(n5226), .Z(n5261) );
  NANDN U5404 ( .A(n5229), .B(n5228), .Z(n5233) );
  NANDN U5405 ( .A(n5231), .B(n5230), .Z(n5232) );
  AND U5406 ( .A(n5233), .B(n5232), .Z(n5265) );
  NANDN U5407 ( .A(n5235), .B(n5234), .Z(n5239) );
  NAND U5408 ( .A(n5237), .B(n5236), .Z(n5238) );
  AND U5409 ( .A(n5239), .B(n5238), .Z(n5282) );
  NANDN U5410 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U5411 ( .A(n5243), .B(n5242), .Z(n5244) );
  AND U5412 ( .A(n5245), .B(n5244), .Z(n5280) );
  NANDN U5413 ( .A(n5274), .B(n5246), .Z(n5248) );
  XOR U5414 ( .A(b[7]), .B(a[126]), .Z(n5273) );
  NANDN U5415 ( .A(n5275), .B(n5273), .Z(n5247) );
  AND U5416 ( .A(n5248), .B(n5247), .Z(n5270) );
  AND U5417 ( .A(b[7]), .B(a[124]), .Z(n5278) );
  IV U5418 ( .A(n5278), .Z(n5288) );
  ANDN U5419 ( .B(n5250), .A(n5249), .Z(n5253) );
  NAND U5420 ( .A(b[5]), .B(n5251), .Z(n5252) );
  NANDN U5421 ( .A(n5253), .B(n5252), .Z(n5268) );
  XOR U5422 ( .A(n5288), .B(n5268), .Z(n5269) );
  NANDN U5423 ( .A(n5255), .B(n5254), .Z(n5259) );
  NAND U5424 ( .A(n5257), .B(n5256), .Z(n5258) );
  NAND U5425 ( .A(n5259), .B(n5258), .Z(n5262) );
  XOR U5426 ( .A(n5263), .B(n5262), .Z(n5264) );
  XOR U5427 ( .A(n5265), .B(n5264), .Z(n5260) );
  XOR U5428 ( .A(n5261), .B(n5260), .Z(c[252]) );
  AND U5429 ( .A(n5261), .B(n5260), .Z(n5297) );
  NAND U5430 ( .A(n5263), .B(n5262), .Z(n5267) );
  NANDN U5431 ( .A(n5265), .B(n5264), .Z(n5266) );
  AND U5432 ( .A(n5267), .B(n5266), .Z(n5307) );
  NANDN U5433 ( .A(n5278), .B(n5268), .Z(n5272) );
  NANDN U5434 ( .A(n5270), .B(n5269), .Z(n5271) );
  AND U5435 ( .A(n5272), .B(n5271), .Z(n5301) );
  NANDN U5436 ( .A(n5274), .B(n5273), .Z(n5277) );
  XOR U5437 ( .A(a[127]), .B(b[7]), .Z(n5292) );
  NANDN U5438 ( .A(n5275), .B(n5292), .Z(n5276) );
  AND U5439 ( .A(n5277), .B(n5276), .Z(n5299) );
  AND U5440 ( .A(b[7]), .B(a[125]), .Z(n5286) );
  XNOR U5441 ( .A(n5285), .B(n5286), .Z(n5287) );
  XOR U5442 ( .A(n5287), .B(n5278), .Z(n5298) );
  NANDN U5443 ( .A(n5280), .B(n5279), .Z(n5284) );
  NANDN U5444 ( .A(n5282), .B(n5281), .Z(n5283) );
  AND U5445 ( .A(n5284), .B(n5283), .Z(n5305) );
  XOR U5446 ( .A(n5304), .B(n5305), .Z(n5306) );
  XOR U5447 ( .A(n5307), .B(n5306), .Z(n5296) );
  XOR U5448 ( .A(n5297), .B(n5296), .Z(c[253]) );
  ANDN U5449 ( .B(n5286), .A(n5285), .Z(n5290) );
  NANDN U5450 ( .A(n5288), .B(n5287), .Z(n5289) );
  NANDN U5451 ( .A(n5290), .B(n5289), .Z(n5319) );
  NAND U5452 ( .A(b[7]), .B(a[126]), .Z(n5317) );
  NAND U5453 ( .A(b[7]), .B(n5291), .Z(n5295) );
  NAND U5454 ( .A(n5293), .B(n5292), .Z(n5294) );
  NAND U5455 ( .A(n5295), .B(n5294), .Z(n5316) );
  XNOR U5456 ( .A(n5317), .B(n5316), .Z(n5318) );
  AND U5457 ( .A(n5297), .B(n5296), .Z(n5315) );
  XNOR U5458 ( .A(n5314), .B(n5315), .Z(n5311) );
  NANDN U5459 ( .A(n5299), .B(n5298), .Z(n5303) );
  NANDN U5460 ( .A(n5301), .B(n5300), .Z(n5302) );
  AND U5461 ( .A(n5303), .B(n5302), .Z(n5312) );
  NAND U5462 ( .A(n5305), .B(n5304), .Z(n5309) );
  NANDN U5463 ( .A(n5307), .B(n5306), .Z(n5308) );
  AND U5464 ( .A(n5309), .B(n5308), .Z(n5313) );
  XOR U5465 ( .A(n5312), .B(n5313), .Z(n5310) );
  XNOR U5466 ( .A(n5311), .B(n5310), .Z(c[254]) );
endmodule

