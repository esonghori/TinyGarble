
module FA_0 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_1023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_1000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_99 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_98 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_97 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_95 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_94 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_93 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_92 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_91 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_90 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_89 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_88 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_87 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_86 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_85 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_84 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_83 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_82 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_81 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_80 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_79 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_78 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_77 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_76 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_75 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_74 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_73 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_72 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_71 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_70 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_69 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_68 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_67 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_66 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_65 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_63 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_62 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_61 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_60 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_59 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_58 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_57 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_56 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_55 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_54 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_53 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_52 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_51 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_50 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_49 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_48 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_47 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_46 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_45 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_44 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_43 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_42 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_41 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_40 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_39 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_38 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_37 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_36 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_35 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_34 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_33 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_31 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_30 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_29 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_28 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_27 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_26 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_25 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_24 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_23 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_22 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_21 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_20 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_19 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_18 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_17 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_16 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_15 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_14 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_13 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_12 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_11 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_10 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_9 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_8 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_7 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_6 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_5 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(CI), .B(A), .Z(n1) );
endmodule


module FA_4 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(B), .Z(S) );
  AND U2 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_3 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(B), .Z(S) );
  AND U2 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_2 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(B), .Z(S) );
  AND U2 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_1 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(B), .Z(S) );
endmodule


module ADD_N1024 ( A, B, CI, S, CO );
  input [1023:0] A;
  input [1023:0] B;
  output [1023:0] S;
  input CI;
  output CO;

  wire   [1023:1] C;

  FA_0 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(
        S[0]), .CO(C[1]) );
  FA_1023 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_1022 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_1021 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_1020 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_1019 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_1018 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_1017 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_1016 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_1015 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_1014 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_1013 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_1012 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_1011 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_1010 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_1009 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_1008 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_1007 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_1006 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_1005 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_1004 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_1003 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_1002 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_1001 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_1000 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_999 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_998 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_997 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_996 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_995 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_994 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_993 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_992 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_991 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_990 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_989 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_988 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_987 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_986 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_985 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_984 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_983 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_982 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_981 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_980 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_979 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_978 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_977 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_976 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_975 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_974 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_973 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_972 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_971 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_970 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_969 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_968 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_967 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_966 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_965 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_964 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_963 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_962 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_961 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_960 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_959 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_958 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_957 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_956 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_955 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_954 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_953 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_952 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_951 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_950 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_949 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_948 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_947 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_946 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_945 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_944 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_943 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_942 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_941 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_940 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_939 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_938 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_937 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_936 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_935 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_934 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_933 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_932 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_931 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_930 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_929 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_928 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_927 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_926 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_925 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_924 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_923 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_922 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_921 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_920 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_919 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_918 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_917 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_916 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_915 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_914 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_913 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_912 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_911 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_910 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_909 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_908 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_907 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_906 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_905 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_904 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_903 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_902 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_901 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_900 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_899 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_898 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_897 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_896 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_895 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_894 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_893 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_892 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_891 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_890 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_889 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_888 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_887 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_886 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_885 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_884 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_883 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_882 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_881 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_880 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_879 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_878 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_877 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_876 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_875 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_874 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_873 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_872 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_871 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_870 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_869 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_868 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_867 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_866 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_865 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_864 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_863 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_862 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_861 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_860 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_859 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_858 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_857 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_856 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_855 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_854 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_853 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_852 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_851 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_850 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_849 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_848 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_847 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_846 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_845 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_844 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_843 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_842 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_841 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_840 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_839 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_838 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_837 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_836 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_835 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_834 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_833 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_832 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_831 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_830 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_829 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_828 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_827 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_826 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_825 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_824 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_823 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_822 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_821 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_820 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_819 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_818 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_817 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_816 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_815 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_814 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_813 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_812 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_811 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_810 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_809 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_808 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_807 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_806 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_805 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_804 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_803 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_802 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_801 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_800 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_799 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_798 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_797 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_796 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_795 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_794 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_793 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_792 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_791 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_790 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_789 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_788 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_787 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_786 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_785 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_784 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_783 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_782 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_781 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_780 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_779 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_778 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_777 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_776 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_775 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_774 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_773 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_772 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_771 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_770 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_769 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_768 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_767 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_766 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_765 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_764 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_763 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_762 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_761 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_760 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_759 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_758 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_757 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_756 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_755 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_754 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_753 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_752 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_751 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_750 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_749 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_748 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_747 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_746 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_745 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_744 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_743 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_742 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_741 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_740 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_739 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_738 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_737 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_736 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_735 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_734 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_733 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_732 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_731 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_730 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_729 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_728 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_727 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_726 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_725 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_724 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_723 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_722 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_721 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_720 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_719 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_718 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_717 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_716 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_715 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_714 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_713 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_712 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_711 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_710 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_709 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_708 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_707 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_706 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_705 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_704 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_703 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_702 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_701 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_700 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_699 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_698 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_697 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_696 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_695 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_694 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_693 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_692 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_691 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_690 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_689 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_688 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_687 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_686 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_685 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_684 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_683 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_682 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_681 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_680 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_679 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_678 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_677 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_676 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_675 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_674 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_673 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_672 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_671 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_670 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_669 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_668 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_667 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_666 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_665 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_664 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_663 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_662 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_661 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_660 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_659 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_658 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_657 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_656 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_655 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_654 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_653 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_652 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_651 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_650 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_649 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_648 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_647 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_646 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_645 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_644 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_643 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_642 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_641 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_640 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_639 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_638 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_637 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_636 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_635 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_634 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_633 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_632 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_631 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_630 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_629 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_628 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_627 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_626 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_625 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_624 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_623 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_622 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_621 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_620 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_619 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_618 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_617 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_616 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_615 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_614 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_613 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_612 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_611 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_610 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_609 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_608 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_607 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_606 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_605 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_604 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_603 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_602 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_601 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_600 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_599 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_598 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_597 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_596 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_595 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_594 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_593 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_592 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_591 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_590 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_589 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_588 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_587 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_586 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_585 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_584 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_583 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_582 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_581 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_580 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_579 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_578 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_577 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_576 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_575 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_574 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_573 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_572 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_571 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_570 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_569 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_568 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_567 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_566 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_565 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_564 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_563 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_562 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_561 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_560 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_559 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_558 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_557 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_556 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_555 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_554 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_553 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_552 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_551 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_550 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_549 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_548 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_547 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_546 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_545 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_544 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_543 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_542 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_541 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_540 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_539 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_538 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_537 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_536 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_535 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_534 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_533 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_532 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_531 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_530 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_529 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_528 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_527 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_526 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_525 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_524 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_523 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_522 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_521 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_520 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_519 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_518 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_517 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_516 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_515 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_514 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_513 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_512 \FA_INST_0[1].FA_INST_1[0].FA_  ( .A(A[512]), .B(B[512]), .CI(C[512]), 
        .S(S[512]), .CO(C[513]) );
  FA_511 \FA_INST_0[1].FA_INST_1[1].FA_  ( .A(A[513]), .B(B[513]), .CI(C[513]), 
        .S(S[513]), .CO(C[514]) );
  FA_510 \FA_INST_0[1].FA_INST_1[2].FA_  ( .A(A[514]), .B(B[514]), .CI(C[514]), 
        .S(S[514]), .CO(C[515]) );
  FA_509 \FA_INST_0[1].FA_INST_1[3].FA_  ( .A(A[515]), .B(B[515]), .CI(C[515]), 
        .S(S[515]), .CO(C[516]) );
  FA_508 \FA_INST_0[1].FA_INST_1[4].FA_  ( .A(A[516]), .B(B[516]), .CI(C[516]), 
        .S(S[516]), .CO(C[517]) );
  FA_507 \FA_INST_0[1].FA_INST_1[5].FA_  ( .A(A[517]), .B(B[517]), .CI(C[517]), 
        .S(S[517]), .CO(C[518]) );
  FA_506 \FA_INST_0[1].FA_INST_1[6].FA_  ( .A(A[518]), .B(B[518]), .CI(C[518]), 
        .S(S[518]), .CO(C[519]) );
  FA_505 \FA_INST_0[1].FA_INST_1[7].FA_  ( .A(A[519]), .B(B[519]), .CI(C[519]), 
        .S(S[519]), .CO(C[520]) );
  FA_504 \FA_INST_0[1].FA_INST_1[8].FA_  ( .A(A[520]), .B(B[520]), .CI(C[520]), 
        .S(S[520]), .CO(C[521]) );
  FA_503 \FA_INST_0[1].FA_INST_1[9].FA_  ( .A(A[521]), .B(B[521]), .CI(C[521]), 
        .S(S[521]), .CO(C[522]) );
  FA_502 \FA_INST_0[1].FA_INST_1[10].FA_  ( .A(A[522]), .B(B[522]), .CI(C[522]), .S(S[522]), .CO(C[523]) );
  FA_501 \FA_INST_0[1].FA_INST_1[11].FA_  ( .A(A[523]), .B(B[523]), .CI(C[523]), .S(S[523]), .CO(C[524]) );
  FA_500 \FA_INST_0[1].FA_INST_1[12].FA_  ( .A(A[524]), .B(B[524]), .CI(C[524]), .S(S[524]), .CO(C[525]) );
  FA_499 \FA_INST_0[1].FA_INST_1[13].FA_  ( .A(A[525]), .B(B[525]), .CI(C[525]), .S(S[525]), .CO(C[526]) );
  FA_498 \FA_INST_0[1].FA_INST_1[14].FA_  ( .A(A[526]), .B(B[526]), .CI(C[526]), .S(S[526]), .CO(C[527]) );
  FA_497 \FA_INST_0[1].FA_INST_1[15].FA_  ( .A(A[527]), .B(B[527]), .CI(C[527]), .S(S[527]), .CO(C[528]) );
  FA_496 \FA_INST_0[1].FA_INST_1[16].FA_  ( .A(A[528]), .B(B[528]), .CI(C[528]), .S(S[528]), .CO(C[529]) );
  FA_495 \FA_INST_0[1].FA_INST_1[17].FA_  ( .A(A[529]), .B(B[529]), .CI(C[529]), .S(S[529]), .CO(C[530]) );
  FA_494 \FA_INST_0[1].FA_INST_1[18].FA_  ( .A(A[530]), .B(B[530]), .CI(C[530]), .S(S[530]), .CO(C[531]) );
  FA_493 \FA_INST_0[1].FA_INST_1[19].FA_  ( .A(A[531]), .B(B[531]), .CI(C[531]), .S(S[531]), .CO(C[532]) );
  FA_492 \FA_INST_0[1].FA_INST_1[20].FA_  ( .A(A[532]), .B(B[532]), .CI(C[532]), .S(S[532]), .CO(C[533]) );
  FA_491 \FA_INST_0[1].FA_INST_1[21].FA_  ( .A(A[533]), .B(B[533]), .CI(C[533]), .S(S[533]), .CO(C[534]) );
  FA_490 \FA_INST_0[1].FA_INST_1[22].FA_  ( .A(A[534]), .B(B[534]), .CI(C[534]), .S(S[534]), .CO(C[535]) );
  FA_489 \FA_INST_0[1].FA_INST_1[23].FA_  ( .A(A[535]), .B(B[535]), .CI(C[535]), .S(S[535]), .CO(C[536]) );
  FA_488 \FA_INST_0[1].FA_INST_1[24].FA_  ( .A(A[536]), .B(B[536]), .CI(C[536]), .S(S[536]), .CO(C[537]) );
  FA_487 \FA_INST_0[1].FA_INST_1[25].FA_  ( .A(A[537]), .B(B[537]), .CI(C[537]), .S(S[537]), .CO(C[538]) );
  FA_486 \FA_INST_0[1].FA_INST_1[26].FA_  ( .A(A[538]), .B(B[538]), .CI(C[538]), .S(S[538]), .CO(C[539]) );
  FA_485 \FA_INST_0[1].FA_INST_1[27].FA_  ( .A(A[539]), .B(B[539]), .CI(C[539]), .S(S[539]), .CO(C[540]) );
  FA_484 \FA_INST_0[1].FA_INST_1[28].FA_  ( .A(A[540]), .B(B[540]), .CI(C[540]), .S(S[540]), .CO(C[541]) );
  FA_483 \FA_INST_0[1].FA_INST_1[29].FA_  ( .A(A[541]), .B(B[541]), .CI(C[541]), .S(S[541]), .CO(C[542]) );
  FA_482 \FA_INST_0[1].FA_INST_1[30].FA_  ( .A(A[542]), .B(B[542]), .CI(C[542]), .S(S[542]), .CO(C[543]) );
  FA_481 \FA_INST_0[1].FA_INST_1[31].FA_  ( .A(A[543]), .B(B[543]), .CI(C[543]), .S(S[543]), .CO(C[544]) );
  FA_480 \FA_INST_0[1].FA_INST_1[32].FA_  ( .A(A[544]), .B(B[544]), .CI(C[544]), .S(S[544]), .CO(C[545]) );
  FA_479 \FA_INST_0[1].FA_INST_1[33].FA_  ( .A(A[545]), .B(B[545]), .CI(C[545]), .S(S[545]), .CO(C[546]) );
  FA_478 \FA_INST_0[1].FA_INST_1[34].FA_  ( .A(A[546]), .B(B[546]), .CI(C[546]), .S(S[546]), .CO(C[547]) );
  FA_477 \FA_INST_0[1].FA_INST_1[35].FA_  ( .A(A[547]), .B(B[547]), .CI(C[547]), .S(S[547]), .CO(C[548]) );
  FA_476 \FA_INST_0[1].FA_INST_1[36].FA_  ( .A(A[548]), .B(B[548]), .CI(C[548]), .S(S[548]), .CO(C[549]) );
  FA_475 \FA_INST_0[1].FA_INST_1[37].FA_  ( .A(A[549]), .B(B[549]), .CI(C[549]), .S(S[549]), .CO(C[550]) );
  FA_474 \FA_INST_0[1].FA_INST_1[38].FA_  ( .A(A[550]), .B(B[550]), .CI(C[550]), .S(S[550]), .CO(C[551]) );
  FA_473 \FA_INST_0[1].FA_INST_1[39].FA_  ( .A(A[551]), .B(B[551]), .CI(C[551]), .S(S[551]), .CO(C[552]) );
  FA_472 \FA_INST_0[1].FA_INST_1[40].FA_  ( .A(A[552]), .B(B[552]), .CI(C[552]), .S(S[552]), .CO(C[553]) );
  FA_471 \FA_INST_0[1].FA_INST_1[41].FA_  ( .A(A[553]), .B(B[553]), .CI(C[553]), .S(S[553]), .CO(C[554]) );
  FA_470 \FA_INST_0[1].FA_INST_1[42].FA_  ( .A(A[554]), .B(B[554]), .CI(C[554]), .S(S[554]), .CO(C[555]) );
  FA_469 \FA_INST_0[1].FA_INST_1[43].FA_  ( .A(A[555]), .B(B[555]), .CI(C[555]), .S(S[555]), .CO(C[556]) );
  FA_468 \FA_INST_0[1].FA_INST_1[44].FA_  ( .A(A[556]), .B(B[556]), .CI(C[556]), .S(S[556]), .CO(C[557]) );
  FA_467 \FA_INST_0[1].FA_INST_1[45].FA_  ( .A(A[557]), .B(B[557]), .CI(C[557]), .S(S[557]), .CO(C[558]) );
  FA_466 \FA_INST_0[1].FA_INST_1[46].FA_  ( .A(A[558]), .B(B[558]), .CI(C[558]), .S(S[558]), .CO(C[559]) );
  FA_465 \FA_INST_0[1].FA_INST_1[47].FA_  ( .A(A[559]), .B(B[559]), .CI(C[559]), .S(S[559]), .CO(C[560]) );
  FA_464 \FA_INST_0[1].FA_INST_1[48].FA_  ( .A(A[560]), .B(B[560]), .CI(C[560]), .S(S[560]), .CO(C[561]) );
  FA_463 \FA_INST_0[1].FA_INST_1[49].FA_  ( .A(A[561]), .B(B[561]), .CI(C[561]), .S(S[561]), .CO(C[562]) );
  FA_462 \FA_INST_0[1].FA_INST_1[50].FA_  ( .A(A[562]), .B(B[562]), .CI(C[562]), .S(S[562]), .CO(C[563]) );
  FA_461 \FA_INST_0[1].FA_INST_1[51].FA_  ( .A(A[563]), .B(B[563]), .CI(C[563]), .S(S[563]), .CO(C[564]) );
  FA_460 \FA_INST_0[1].FA_INST_1[52].FA_  ( .A(A[564]), .B(B[564]), .CI(C[564]), .S(S[564]), .CO(C[565]) );
  FA_459 \FA_INST_0[1].FA_INST_1[53].FA_  ( .A(A[565]), .B(B[565]), .CI(C[565]), .S(S[565]), .CO(C[566]) );
  FA_458 \FA_INST_0[1].FA_INST_1[54].FA_  ( .A(A[566]), .B(B[566]), .CI(C[566]), .S(S[566]), .CO(C[567]) );
  FA_457 \FA_INST_0[1].FA_INST_1[55].FA_  ( .A(A[567]), .B(B[567]), .CI(C[567]), .S(S[567]), .CO(C[568]) );
  FA_456 \FA_INST_0[1].FA_INST_1[56].FA_  ( .A(A[568]), .B(B[568]), .CI(C[568]), .S(S[568]), .CO(C[569]) );
  FA_455 \FA_INST_0[1].FA_INST_1[57].FA_  ( .A(A[569]), .B(B[569]), .CI(C[569]), .S(S[569]), .CO(C[570]) );
  FA_454 \FA_INST_0[1].FA_INST_1[58].FA_  ( .A(A[570]), .B(B[570]), .CI(C[570]), .S(S[570]), .CO(C[571]) );
  FA_453 \FA_INST_0[1].FA_INST_1[59].FA_  ( .A(A[571]), .B(B[571]), .CI(C[571]), .S(S[571]), .CO(C[572]) );
  FA_452 \FA_INST_0[1].FA_INST_1[60].FA_  ( .A(A[572]), .B(B[572]), .CI(C[572]), .S(S[572]), .CO(C[573]) );
  FA_451 \FA_INST_0[1].FA_INST_1[61].FA_  ( .A(A[573]), .B(B[573]), .CI(C[573]), .S(S[573]), .CO(C[574]) );
  FA_450 \FA_INST_0[1].FA_INST_1[62].FA_  ( .A(A[574]), .B(B[574]), .CI(C[574]), .S(S[574]), .CO(C[575]) );
  FA_449 \FA_INST_0[1].FA_INST_1[63].FA_  ( .A(A[575]), .B(B[575]), .CI(C[575]), .S(S[575]), .CO(C[576]) );
  FA_448 \FA_INST_0[1].FA_INST_1[64].FA_  ( .A(A[576]), .B(B[576]), .CI(C[576]), .S(S[576]), .CO(C[577]) );
  FA_447 \FA_INST_0[1].FA_INST_1[65].FA_  ( .A(A[577]), .B(B[577]), .CI(C[577]), .S(S[577]), .CO(C[578]) );
  FA_446 \FA_INST_0[1].FA_INST_1[66].FA_  ( .A(A[578]), .B(B[578]), .CI(C[578]), .S(S[578]), .CO(C[579]) );
  FA_445 \FA_INST_0[1].FA_INST_1[67].FA_  ( .A(A[579]), .B(B[579]), .CI(C[579]), .S(S[579]), .CO(C[580]) );
  FA_444 \FA_INST_0[1].FA_INST_1[68].FA_  ( .A(A[580]), .B(B[580]), .CI(C[580]), .S(S[580]), .CO(C[581]) );
  FA_443 \FA_INST_0[1].FA_INST_1[69].FA_  ( .A(A[581]), .B(B[581]), .CI(C[581]), .S(S[581]), .CO(C[582]) );
  FA_442 \FA_INST_0[1].FA_INST_1[70].FA_  ( .A(A[582]), .B(B[582]), .CI(C[582]), .S(S[582]), .CO(C[583]) );
  FA_441 \FA_INST_0[1].FA_INST_1[71].FA_  ( .A(A[583]), .B(B[583]), .CI(C[583]), .S(S[583]), .CO(C[584]) );
  FA_440 \FA_INST_0[1].FA_INST_1[72].FA_  ( .A(A[584]), .B(B[584]), .CI(C[584]), .S(S[584]), .CO(C[585]) );
  FA_439 \FA_INST_0[1].FA_INST_1[73].FA_  ( .A(A[585]), .B(B[585]), .CI(C[585]), .S(S[585]), .CO(C[586]) );
  FA_438 \FA_INST_0[1].FA_INST_1[74].FA_  ( .A(A[586]), .B(B[586]), .CI(C[586]), .S(S[586]), .CO(C[587]) );
  FA_437 \FA_INST_0[1].FA_INST_1[75].FA_  ( .A(A[587]), .B(B[587]), .CI(C[587]), .S(S[587]), .CO(C[588]) );
  FA_436 \FA_INST_0[1].FA_INST_1[76].FA_  ( .A(A[588]), .B(B[588]), .CI(C[588]), .S(S[588]), .CO(C[589]) );
  FA_435 \FA_INST_0[1].FA_INST_1[77].FA_  ( .A(A[589]), .B(B[589]), .CI(C[589]), .S(S[589]), .CO(C[590]) );
  FA_434 \FA_INST_0[1].FA_INST_1[78].FA_  ( .A(A[590]), .B(B[590]), .CI(C[590]), .S(S[590]), .CO(C[591]) );
  FA_433 \FA_INST_0[1].FA_INST_1[79].FA_  ( .A(A[591]), .B(B[591]), .CI(C[591]), .S(S[591]), .CO(C[592]) );
  FA_432 \FA_INST_0[1].FA_INST_1[80].FA_  ( .A(A[592]), .B(B[592]), .CI(C[592]), .S(S[592]), .CO(C[593]) );
  FA_431 \FA_INST_0[1].FA_INST_1[81].FA_  ( .A(A[593]), .B(B[593]), .CI(C[593]), .S(S[593]), .CO(C[594]) );
  FA_430 \FA_INST_0[1].FA_INST_1[82].FA_  ( .A(A[594]), .B(B[594]), .CI(C[594]), .S(S[594]), .CO(C[595]) );
  FA_429 \FA_INST_0[1].FA_INST_1[83].FA_  ( .A(A[595]), .B(B[595]), .CI(C[595]), .S(S[595]), .CO(C[596]) );
  FA_428 \FA_INST_0[1].FA_INST_1[84].FA_  ( .A(A[596]), .B(B[596]), .CI(C[596]), .S(S[596]), .CO(C[597]) );
  FA_427 \FA_INST_0[1].FA_INST_1[85].FA_  ( .A(A[597]), .B(B[597]), .CI(C[597]), .S(S[597]), .CO(C[598]) );
  FA_426 \FA_INST_0[1].FA_INST_1[86].FA_  ( .A(A[598]), .B(B[598]), .CI(C[598]), .S(S[598]), .CO(C[599]) );
  FA_425 \FA_INST_0[1].FA_INST_1[87].FA_  ( .A(A[599]), .B(B[599]), .CI(C[599]), .S(S[599]), .CO(C[600]) );
  FA_424 \FA_INST_0[1].FA_INST_1[88].FA_  ( .A(A[600]), .B(B[600]), .CI(C[600]), .S(S[600]), .CO(C[601]) );
  FA_423 \FA_INST_0[1].FA_INST_1[89].FA_  ( .A(A[601]), .B(B[601]), .CI(C[601]), .S(S[601]), .CO(C[602]) );
  FA_422 \FA_INST_0[1].FA_INST_1[90].FA_  ( .A(A[602]), .B(B[602]), .CI(C[602]), .S(S[602]), .CO(C[603]) );
  FA_421 \FA_INST_0[1].FA_INST_1[91].FA_  ( .A(A[603]), .B(B[603]), .CI(C[603]), .S(S[603]), .CO(C[604]) );
  FA_420 \FA_INST_0[1].FA_INST_1[92].FA_  ( .A(A[604]), .B(B[604]), .CI(C[604]), .S(S[604]), .CO(C[605]) );
  FA_419 \FA_INST_0[1].FA_INST_1[93].FA_  ( .A(A[605]), .B(B[605]), .CI(C[605]), .S(S[605]), .CO(C[606]) );
  FA_418 \FA_INST_0[1].FA_INST_1[94].FA_  ( .A(A[606]), .B(B[606]), .CI(C[606]), .S(S[606]), .CO(C[607]) );
  FA_417 \FA_INST_0[1].FA_INST_1[95].FA_  ( .A(A[607]), .B(B[607]), .CI(C[607]), .S(S[607]), .CO(C[608]) );
  FA_416 \FA_INST_0[1].FA_INST_1[96].FA_  ( .A(A[608]), .B(B[608]), .CI(C[608]), .S(S[608]), .CO(C[609]) );
  FA_415 \FA_INST_0[1].FA_INST_1[97].FA_  ( .A(A[609]), .B(B[609]), .CI(C[609]), .S(S[609]), .CO(C[610]) );
  FA_414 \FA_INST_0[1].FA_INST_1[98].FA_  ( .A(A[610]), .B(B[610]), .CI(C[610]), .S(S[610]), .CO(C[611]) );
  FA_413 \FA_INST_0[1].FA_INST_1[99].FA_  ( .A(A[611]), .B(B[611]), .CI(C[611]), .S(S[611]), .CO(C[612]) );
  FA_412 \FA_INST_0[1].FA_INST_1[100].FA_  ( .A(A[612]), .B(B[612]), .CI(
        C[612]), .S(S[612]), .CO(C[613]) );
  FA_411 \FA_INST_0[1].FA_INST_1[101].FA_  ( .A(A[613]), .B(B[613]), .CI(
        C[613]), .S(S[613]), .CO(C[614]) );
  FA_410 \FA_INST_0[1].FA_INST_1[102].FA_  ( .A(A[614]), .B(B[614]), .CI(
        C[614]), .S(S[614]), .CO(C[615]) );
  FA_409 \FA_INST_0[1].FA_INST_1[103].FA_  ( .A(A[615]), .B(B[615]), .CI(
        C[615]), .S(S[615]), .CO(C[616]) );
  FA_408 \FA_INST_0[1].FA_INST_1[104].FA_  ( .A(A[616]), .B(B[616]), .CI(
        C[616]), .S(S[616]), .CO(C[617]) );
  FA_407 \FA_INST_0[1].FA_INST_1[105].FA_  ( .A(A[617]), .B(B[617]), .CI(
        C[617]), .S(S[617]), .CO(C[618]) );
  FA_406 \FA_INST_0[1].FA_INST_1[106].FA_  ( .A(A[618]), .B(B[618]), .CI(
        C[618]), .S(S[618]), .CO(C[619]) );
  FA_405 \FA_INST_0[1].FA_INST_1[107].FA_  ( .A(A[619]), .B(B[619]), .CI(
        C[619]), .S(S[619]), .CO(C[620]) );
  FA_404 \FA_INST_0[1].FA_INST_1[108].FA_  ( .A(A[620]), .B(B[620]), .CI(
        C[620]), .S(S[620]), .CO(C[621]) );
  FA_403 \FA_INST_0[1].FA_INST_1[109].FA_  ( .A(A[621]), .B(B[621]), .CI(
        C[621]), .S(S[621]), .CO(C[622]) );
  FA_402 \FA_INST_0[1].FA_INST_1[110].FA_  ( .A(A[622]), .B(B[622]), .CI(
        C[622]), .S(S[622]), .CO(C[623]) );
  FA_401 \FA_INST_0[1].FA_INST_1[111].FA_  ( .A(A[623]), .B(B[623]), .CI(
        C[623]), .S(S[623]), .CO(C[624]) );
  FA_400 \FA_INST_0[1].FA_INST_1[112].FA_  ( .A(A[624]), .B(B[624]), .CI(
        C[624]), .S(S[624]), .CO(C[625]) );
  FA_399 \FA_INST_0[1].FA_INST_1[113].FA_  ( .A(A[625]), .B(B[625]), .CI(
        C[625]), .S(S[625]), .CO(C[626]) );
  FA_398 \FA_INST_0[1].FA_INST_1[114].FA_  ( .A(A[626]), .B(B[626]), .CI(
        C[626]), .S(S[626]), .CO(C[627]) );
  FA_397 \FA_INST_0[1].FA_INST_1[115].FA_  ( .A(A[627]), .B(B[627]), .CI(
        C[627]), .S(S[627]), .CO(C[628]) );
  FA_396 \FA_INST_0[1].FA_INST_1[116].FA_  ( .A(A[628]), .B(B[628]), .CI(
        C[628]), .S(S[628]), .CO(C[629]) );
  FA_395 \FA_INST_0[1].FA_INST_1[117].FA_  ( .A(A[629]), .B(B[629]), .CI(
        C[629]), .S(S[629]), .CO(C[630]) );
  FA_394 \FA_INST_0[1].FA_INST_1[118].FA_  ( .A(A[630]), .B(B[630]), .CI(
        C[630]), .S(S[630]), .CO(C[631]) );
  FA_393 \FA_INST_0[1].FA_INST_1[119].FA_  ( .A(A[631]), .B(B[631]), .CI(
        C[631]), .S(S[631]), .CO(C[632]) );
  FA_392 \FA_INST_0[1].FA_INST_1[120].FA_  ( .A(A[632]), .B(B[632]), .CI(
        C[632]), .S(S[632]), .CO(C[633]) );
  FA_391 \FA_INST_0[1].FA_INST_1[121].FA_  ( .A(A[633]), .B(B[633]), .CI(
        C[633]), .S(S[633]), .CO(C[634]) );
  FA_390 \FA_INST_0[1].FA_INST_1[122].FA_  ( .A(A[634]), .B(B[634]), .CI(
        C[634]), .S(S[634]), .CO(C[635]) );
  FA_389 \FA_INST_0[1].FA_INST_1[123].FA_  ( .A(A[635]), .B(B[635]), .CI(
        C[635]), .S(S[635]), .CO(C[636]) );
  FA_388 \FA_INST_0[1].FA_INST_1[124].FA_  ( .A(A[636]), .B(B[636]), .CI(
        C[636]), .S(S[636]), .CO(C[637]) );
  FA_387 \FA_INST_0[1].FA_INST_1[125].FA_  ( .A(A[637]), .B(B[637]), .CI(
        C[637]), .S(S[637]), .CO(C[638]) );
  FA_386 \FA_INST_0[1].FA_INST_1[126].FA_  ( .A(A[638]), .B(B[638]), .CI(
        C[638]), .S(S[638]), .CO(C[639]) );
  FA_385 \FA_INST_0[1].FA_INST_1[127].FA_  ( .A(A[639]), .B(B[639]), .CI(
        C[639]), .S(S[639]), .CO(C[640]) );
  FA_384 \FA_INST_0[1].FA_INST_1[128].FA_  ( .A(A[640]), .B(B[640]), .CI(
        C[640]), .S(S[640]), .CO(C[641]) );
  FA_383 \FA_INST_0[1].FA_INST_1[129].FA_  ( .A(A[641]), .B(B[641]), .CI(
        C[641]), .S(S[641]), .CO(C[642]) );
  FA_382 \FA_INST_0[1].FA_INST_1[130].FA_  ( .A(A[642]), .B(B[642]), .CI(
        C[642]), .S(S[642]), .CO(C[643]) );
  FA_381 \FA_INST_0[1].FA_INST_1[131].FA_  ( .A(A[643]), .B(B[643]), .CI(
        C[643]), .S(S[643]), .CO(C[644]) );
  FA_380 \FA_INST_0[1].FA_INST_1[132].FA_  ( .A(A[644]), .B(B[644]), .CI(
        C[644]), .S(S[644]), .CO(C[645]) );
  FA_379 \FA_INST_0[1].FA_INST_1[133].FA_  ( .A(A[645]), .B(B[645]), .CI(
        C[645]), .S(S[645]), .CO(C[646]) );
  FA_378 \FA_INST_0[1].FA_INST_1[134].FA_  ( .A(A[646]), .B(B[646]), .CI(
        C[646]), .S(S[646]), .CO(C[647]) );
  FA_377 \FA_INST_0[1].FA_INST_1[135].FA_  ( .A(A[647]), .B(B[647]), .CI(
        C[647]), .S(S[647]), .CO(C[648]) );
  FA_376 \FA_INST_0[1].FA_INST_1[136].FA_  ( .A(A[648]), .B(B[648]), .CI(
        C[648]), .S(S[648]), .CO(C[649]) );
  FA_375 \FA_INST_0[1].FA_INST_1[137].FA_  ( .A(A[649]), .B(B[649]), .CI(
        C[649]), .S(S[649]), .CO(C[650]) );
  FA_374 \FA_INST_0[1].FA_INST_1[138].FA_  ( .A(A[650]), .B(B[650]), .CI(
        C[650]), .S(S[650]), .CO(C[651]) );
  FA_373 \FA_INST_0[1].FA_INST_1[139].FA_  ( .A(A[651]), .B(B[651]), .CI(
        C[651]), .S(S[651]), .CO(C[652]) );
  FA_372 \FA_INST_0[1].FA_INST_1[140].FA_  ( .A(A[652]), .B(B[652]), .CI(
        C[652]), .S(S[652]), .CO(C[653]) );
  FA_371 \FA_INST_0[1].FA_INST_1[141].FA_  ( .A(A[653]), .B(B[653]), .CI(
        C[653]), .S(S[653]), .CO(C[654]) );
  FA_370 \FA_INST_0[1].FA_INST_1[142].FA_  ( .A(A[654]), .B(B[654]), .CI(
        C[654]), .S(S[654]), .CO(C[655]) );
  FA_369 \FA_INST_0[1].FA_INST_1[143].FA_  ( .A(A[655]), .B(B[655]), .CI(
        C[655]), .S(S[655]), .CO(C[656]) );
  FA_368 \FA_INST_0[1].FA_INST_1[144].FA_  ( .A(A[656]), .B(B[656]), .CI(
        C[656]), .S(S[656]), .CO(C[657]) );
  FA_367 \FA_INST_0[1].FA_INST_1[145].FA_  ( .A(A[657]), .B(B[657]), .CI(
        C[657]), .S(S[657]), .CO(C[658]) );
  FA_366 \FA_INST_0[1].FA_INST_1[146].FA_  ( .A(A[658]), .B(B[658]), .CI(
        C[658]), .S(S[658]), .CO(C[659]) );
  FA_365 \FA_INST_0[1].FA_INST_1[147].FA_  ( .A(A[659]), .B(B[659]), .CI(
        C[659]), .S(S[659]), .CO(C[660]) );
  FA_364 \FA_INST_0[1].FA_INST_1[148].FA_  ( .A(A[660]), .B(B[660]), .CI(
        C[660]), .S(S[660]), .CO(C[661]) );
  FA_363 \FA_INST_0[1].FA_INST_1[149].FA_  ( .A(A[661]), .B(B[661]), .CI(
        C[661]), .S(S[661]), .CO(C[662]) );
  FA_362 \FA_INST_0[1].FA_INST_1[150].FA_  ( .A(A[662]), .B(B[662]), .CI(
        C[662]), .S(S[662]), .CO(C[663]) );
  FA_361 \FA_INST_0[1].FA_INST_1[151].FA_  ( .A(A[663]), .B(B[663]), .CI(
        C[663]), .S(S[663]), .CO(C[664]) );
  FA_360 \FA_INST_0[1].FA_INST_1[152].FA_  ( .A(A[664]), .B(B[664]), .CI(
        C[664]), .S(S[664]), .CO(C[665]) );
  FA_359 \FA_INST_0[1].FA_INST_1[153].FA_  ( .A(A[665]), .B(B[665]), .CI(
        C[665]), .S(S[665]), .CO(C[666]) );
  FA_358 \FA_INST_0[1].FA_INST_1[154].FA_  ( .A(A[666]), .B(B[666]), .CI(
        C[666]), .S(S[666]), .CO(C[667]) );
  FA_357 \FA_INST_0[1].FA_INST_1[155].FA_  ( .A(A[667]), .B(B[667]), .CI(
        C[667]), .S(S[667]), .CO(C[668]) );
  FA_356 \FA_INST_0[1].FA_INST_1[156].FA_  ( .A(A[668]), .B(B[668]), .CI(
        C[668]), .S(S[668]), .CO(C[669]) );
  FA_355 \FA_INST_0[1].FA_INST_1[157].FA_  ( .A(A[669]), .B(B[669]), .CI(
        C[669]), .S(S[669]), .CO(C[670]) );
  FA_354 \FA_INST_0[1].FA_INST_1[158].FA_  ( .A(A[670]), .B(B[670]), .CI(
        C[670]), .S(S[670]), .CO(C[671]) );
  FA_353 \FA_INST_0[1].FA_INST_1[159].FA_  ( .A(A[671]), .B(B[671]), .CI(
        C[671]), .S(S[671]), .CO(C[672]) );
  FA_352 \FA_INST_0[1].FA_INST_1[160].FA_  ( .A(A[672]), .B(B[672]), .CI(
        C[672]), .S(S[672]), .CO(C[673]) );
  FA_351 \FA_INST_0[1].FA_INST_1[161].FA_  ( .A(A[673]), .B(B[673]), .CI(
        C[673]), .S(S[673]), .CO(C[674]) );
  FA_350 \FA_INST_0[1].FA_INST_1[162].FA_  ( .A(A[674]), .B(B[674]), .CI(
        C[674]), .S(S[674]), .CO(C[675]) );
  FA_349 \FA_INST_0[1].FA_INST_1[163].FA_  ( .A(A[675]), .B(B[675]), .CI(
        C[675]), .S(S[675]), .CO(C[676]) );
  FA_348 \FA_INST_0[1].FA_INST_1[164].FA_  ( .A(A[676]), .B(B[676]), .CI(
        C[676]), .S(S[676]), .CO(C[677]) );
  FA_347 \FA_INST_0[1].FA_INST_1[165].FA_  ( .A(A[677]), .B(B[677]), .CI(
        C[677]), .S(S[677]), .CO(C[678]) );
  FA_346 \FA_INST_0[1].FA_INST_1[166].FA_  ( .A(A[678]), .B(B[678]), .CI(
        C[678]), .S(S[678]), .CO(C[679]) );
  FA_345 \FA_INST_0[1].FA_INST_1[167].FA_  ( .A(A[679]), .B(B[679]), .CI(
        C[679]), .S(S[679]), .CO(C[680]) );
  FA_344 \FA_INST_0[1].FA_INST_1[168].FA_  ( .A(A[680]), .B(B[680]), .CI(
        C[680]), .S(S[680]), .CO(C[681]) );
  FA_343 \FA_INST_0[1].FA_INST_1[169].FA_  ( .A(A[681]), .B(B[681]), .CI(
        C[681]), .S(S[681]), .CO(C[682]) );
  FA_342 \FA_INST_0[1].FA_INST_1[170].FA_  ( .A(A[682]), .B(B[682]), .CI(
        C[682]), .S(S[682]), .CO(C[683]) );
  FA_341 \FA_INST_0[1].FA_INST_1[171].FA_  ( .A(A[683]), .B(B[683]), .CI(
        C[683]), .S(S[683]), .CO(C[684]) );
  FA_340 \FA_INST_0[1].FA_INST_1[172].FA_  ( .A(A[684]), .B(B[684]), .CI(
        C[684]), .S(S[684]), .CO(C[685]) );
  FA_339 \FA_INST_0[1].FA_INST_1[173].FA_  ( .A(A[685]), .B(B[685]), .CI(
        C[685]), .S(S[685]), .CO(C[686]) );
  FA_338 \FA_INST_0[1].FA_INST_1[174].FA_  ( .A(A[686]), .B(B[686]), .CI(
        C[686]), .S(S[686]), .CO(C[687]) );
  FA_337 \FA_INST_0[1].FA_INST_1[175].FA_  ( .A(A[687]), .B(B[687]), .CI(
        C[687]), .S(S[687]), .CO(C[688]) );
  FA_336 \FA_INST_0[1].FA_INST_1[176].FA_  ( .A(A[688]), .B(B[688]), .CI(
        C[688]), .S(S[688]), .CO(C[689]) );
  FA_335 \FA_INST_0[1].FA_INST_1[177].FA_  ( .A(A[689]), .B(B[689]), .CI(
        C[689]), .S(S[689]), .CO(C[690]) );
  FA_334 \FA_INST_0[1].FA_INST_1[178].FA_  ( .A(A[690]), .B(B[690]), .CI(
        C[690]), .S(S[690]), .CO(C[691]) );
  FA_333 \FA_INST_0[1].FA_INST_1[179].FA_  ( .A(A[691]), .B(B[691]), .CI(
        C[691]), .S(S[691]), .CO(C[692]) );
  FA_332 \FA_INST_0[1].FA_INST_1[180].FA_  ( .A(A[692]), .B(B[692]), .CI(
        C[692]), .S(S[692]), .CO(C[693]) );
  FA_331 \FA_INST_0[1].FA_INST_1[181].FA_  ( .A(A[693]), .B(B[693]), .CI(
        C[693]), .S(S[693]), .CO(C[694]) );
  FA_330 \FA_INST_0[1].FA_INST_1[182].FA_  ( .A(A[694]), .B(B[694]), .CI(
        C[694]), .S(S[694]), .CO(C[695]) );
  FA_329 \FA_INST_0[1].FA_INST_1[183].FA_  ( .A(A[695]), .B(B[695]), .CI(
        C[695]), .S(S[695]), .CO(C[696]) );
  FA_328 \FA_INST_0[1].FA_INST_1[184].FA_  ( .A(A[696]), .B(B[696]), .CI(
        C[696]), .S(S[696]), .CO(C[697]) );
  FA_327 \FA_INST_0[1].FA_INST_1[185].FA_  ( .A(A[697]), .B(B[697]), .CI(
        C[697]), .S(S[697]), .CO(C[698]) );
  FA_326 \FA_INST_0[1].FA_INST_1[186].FA_  ( .A(A[698]), .B(B[698]), .CI(
        C[698]), .S(S[698]), .CO(C[699]) );
  FA_325 \FA_INST_0[1].FA_INST_1[187].FA_  ( .A(A[699]), .B(B[699]), .CI(
        C[699]), .S(S[699]), .CO(C[700]) );
  FA_324 \FA_INST_0[1].FA_INST_1[188].FA_  ( .A(A[700]), .B(B[700]), .CI(
        C[700]), .S(S[700]), .CO(C[701]) );
  FA_323 \FA_INST_0[1].FA_INST_1[189].FA_  ( .A(A[701]), .B(B[701]), .CI(
        C[701]), .S(S[701]), .CO(C[702]) );
  FA_322 \FA_INST_0[1].FA_INST_1[190].FA_  ( .A(A[702]), .B(B[702]), .CI(
        C[702]), .S(S[702]), .CO(C[703]) );
  FA_321 \FA_INST_0[1].FA_INST_1[191].FA_  ( .A(A[703]), .B(B[703]), .CI(
        C[703]), .S(S[703]), .CO(C[704]) );
  FA_320 \FA_INST_0[1].FA_INST_1[192].FA_  ( .A(A[704]), .B(B[704]), .CI(
        C[704]), .S(S[704]), .CO(C[705]) );
  FA_319 \FA_INST_0[1].FA_INST_1[193].FA_  ( .A(A[705]), .B(B[705]), .CI(
        C[705]), .S(S[705]), .CO(C[706]) );
  FA_318 \FA_INST_0[1].FA_INST_1[194].FA_  ( .A(A[706]), .B(B[706]), .CI(
        C[706]), .S(S[706]), .CO(C[707]) );
  FA_317 \FA_INST_0[1].FA_INST_1[195].FA_  ( .A(A[707]), .B(B[707]), .CI(
        C[707]), .S(S[707]), .CO(C[708]) );
  FA_316 \FA_INST_0[1].FA_INST_1[196].FA_  ( .A(A[708]), .B(B[708]), .CI(
        C[708]), .S(S[708]), .CO(C[709]) );
  FA_315 \FA_INST_0[1].FA_INST_1[197].FA_  ( .A(A[709]), .B(B[709]), .CI(
        C[709]), .S(S[709]), .CO(C[710]) );
  FA_314 \FA_INST_0[1].FA_INST_1[198].FA_  ( .A(A[710]), .B(B[710]), .CI(
        C[710]), .S(S[710]), .CO(C[711]) );
  FA_313 \FA_INST_0[1].FA_INST_1[199].FA_  ( .A(A[711]), .B(B[711]), .CI(
        C[711]), .S(S[711]), .CO(C[712]) );
  FA_312 \FA_INST_0[1].FA_INST_1[200].FA_  ( .A(A[712]), .B(B[712]), .CI(
        C[712]), .S(S[712]), .CO(C[713]) );
  FA_311 \FA_INST_0[1].FA_INST_1[201].FA_  ( .A(A[713]), .B(B[713]), .CI(
        C[713]), .S(S[713]), .CO(C[714]) );
  FA_310 \FA_INST_0[1].FA_INST_1[202].FA_  ( .A(A[714]), .B(B[714]), .CI(
        C[714]), .S(S[714]), .CO(C[715]) );
  FA_309 \FA_INST_0[1].FA_INST_1[203].FA_  ( .A(A[715]), .B(B[715]), .CI(
        C[715]), .S(S[715]), .CO(C[716]) );
  FA_308 \FA_INST_0[1].FA_INST_1[204].FA_  ( .A(A[716]), .B(B[716]), .CI(
        C[716]), .S(S[716]), .CO(C[717]) );
  FA_307 \FA_INST_0[1].FA_INST_1[205].FA_  ( .A(A[717]), .B(B[717]), .CI(
        C[717]), .S(S[717]), .CO(C[718]) );
  FA_306 \FA_INST_0[1].FA_INST_1[206].FA_  ( .A(A[718]), .B(B[718]), .CI(
        C[718]), .S(S[718]), .CO(C[719]) );
  FA_305 \FA_INST_0[1].FA_INST_1[207].FA_  ( .A(A[719]), .B(B[719]), .CI(
        C[719]), .S(S[719]), .CO(C[720]) );
  FA_304 \FA_INST_0[1].FA_INST_1[208].FA_  ( .A(A[720]), .B(B[720]), .CI(
        C[720]), .S(S[720]), .CO(C[721]) );
  FA_303 \FA_INST_0[1].FA_INST_1[209].FA_  ( .A(A[721]), .B(B[721]), .CI(
        C[721]), .S(S[721]), .CO(C[722]) );
  FA_302 \FA_INST_0[1].FA_INST_1[210].FA_  ( .A(A[722]), .B(B[722]), .CI(
        C[722]), .S(S[722]), .CO(C[723]) );
  FA_301 \FA_INST_0[1].FA_INST_1[211].FA_  ( .A(A[723]), .B(B[723]), .CI(
        C[723]), .S(S[723]), .CO(C[724]) );
  FA_300 \FA_INST_0[1].FA_INST_1[212].FA_  ( .A(A[724]), .B(B[724]), .CI(
        C[724]), .S(S[724]), .CO(C[725]) );
  FA_299 \FA_INST_0[1].FA_INST_1[213].FA_  ( .A(A[725]), .B(B[725]), .CI(
        C[725]), .S(S[725]), .CO(C[726]) );
  FA_298 \FA_INST_0[1].FA_INST_1[214].FA_  ( .A(A[726]), .B(B[726]), .CI(
        C[726]), .S(S[726]), .CO(C[727]) );
  FA_297 \FA_INST_0[1].FA_INST_1[215].FA_  ( .A(A[727]), .B(B[727]), .CI(
        C[727]), .S(S[727]), .CO(C[728]) );
  FA_296 \FA_INST_0[1].FA_INST_1[216].FA_  ( .A(A[728]), .B(B[728]), .CI(
        C[728]), .S(S[728]), .CO(C[729]) );
  FA_295 \FA_INST_0[1].FA_INST_1[217].FA_  ( .A(A[729]), .B(B[729]), .CI(
        C[729]), .S(S[729]), .CO(C[730]) );
  FA_294 \FA_INST_0[1].FA_INST_1[218].FA_  ( .A(A[730]), .B(B[730]), .CI(
        C[730]), .S(S[730]), .CO(C[731]) );
  FA_293 \FA_INST_0[1].FA_INST_1[219].FA_  ( .A(A[731]), .B(B[731]), .CI(
        C[731]), .S(S[731]), .CO(C[732]) );
  FA_292 \FA_INST_0[1].FA_INST_1[220].FA_  ( .A(A[732]), .B(B[732]), .CI(
        C[732]), .S(S[732]), .CO(C[733]) );
  FA_291 \FA_INST_0[1].FA_INST_1[221].FA_  ( .A(A[733]), .B(B[733]), .CI(
        C[733]), .S(S[733]), .CO(C[734]) );
  FA_290 \FA_INST_0[1].FA_INST_1[222].FA_  ( .A(A[734]), .B(B[734]), .CI(
        C[734]), .S(S[734]), .CO(C[735]) );
  FA_289 \FA_INST_0[1].FA_INST_1[223].FA_  ( .A(A[735]), .B(B[735]), .CI(
        C[735]), .S(S[735]), .CO(C[736]) );
  FA_288 \FA_INST_0[1].FA_INST_1[224].FA_  ( .A(A[736]), .B(B[736]), .CI(
        C[736]), .S(S[736]), .CO(C[737]) );
  FA_287 \FA_INST_0[1].FA_INST_1[225].FA_  ( .A(A[737]), .B(B[737]), .CI(
        C[737]), .S(S[737]), .CO(C[738]) );
  FA_286 \FA_INST_0[1].FA_INST_1[226].FA_  ( .A(A[738]), .B(B[738]), .CI(
        C[738]), .S(S[738]), .CO(C[739]) );
  FA_285 \FA_INST_0[1].FA_INST_1[227].FA_  ( .A(A[739]), .B(B[739]), .CI(
        C[739]), .S(S[739]), .CO(C[740]) );
  FA_284 \FA_INST_0[1].FA_INST_1[228].FA_  ( .A(A[740]), .B(B[740]), .CI(
        C[740]), .S(S[740]), .CO(C[741]) );
  FA_283 \FA_INST_0[1].FA_INST_1[229].FA_  ( .A(A[741]), .B(B[741]), .CI(
        C[741]), .S(S[741]), .CO(C[742]) );
  FA_282 \FA_INST_0[1].FA_INST_1[230].FA_  ( .A(A[742]), .B(B[742]), .CI(
        C[742]), .S(S[742]), .CO(C[743]) );
  FA_281 \FA_INST_0[1].FA_INST_1[231].FA_  ( .A(A[743]), .B(B[743]), .CI(
        C[743]), .S(S[743]), .CO(C[744]) );
  FA_280 \FA_INST_0[1].FA_INST_1[232].FA_  ( .A(A[744]), .B(B[744]), .CI(
        C[744]), .S(S[744]), .CO(C[745]) );
  FA_279 \FA_INST_0[1].FA_INST_1[233].FA_  ( .A(A[745]), .B(B[745]), .CI(
        C[745]), .S(S[745]), .CO(C[746]) );
  FA_278 \FA_INST_0[1].FA_INST_1[234].FA_  ( .A(A[746]), .B(B[746]), .CI(
        C[746]), .S(S[746]), .CO(C[747]) );
  FA_277 \FA_INST_0[1].FA_INST_1[235].FA_  ( .A(A[747]), .B(B[747]), .CI(
        C[747]), .S(S[747]), .CO(C[748]) );
  FA_276 \FA_INST_0[1].FA_INST_1[236].FA_  ( .A(A[748]), .B(B[748]), .CI(
        C[748]), .S(S[748]), .CO(C[749]) );
  FA_275 \FA_INST_0[1].FA_INST_1[237].FA_  ( .A(A[749]), .B(B[749]), .CI(
        C[749]), .S(S[749]), .CO(C[750]) );
  FA_274 \FA_INST_0[1].FA_INST_1[238].FA_  ( .A(A[750]), .B(B[750]), .CI(
        C[750]), .S(S[750]), .CO(C[751]) );
  FA_273 \FA_INST_0[1].FA_INST_1[239].FA_  ( .A(A[751]), .B(B[751]), .CI(
        C[751]), .S(S[751]), .CO(C[752]) );
  FA_272 \FA_INST_0[1].FA_INST_1[240].FA_  ( .A(A[752]), .B(B[752]), .CI(
        C[752]), .S(S[752]), .CO(C[753]) );
  FA_271 \FA_INST_0[1].FA_INST_1[241].FA_  ( .A(A[753]), .B(B[753]), .CI(
        C[753]), .S(S[753]), .CO(C[754]) );
  FA_270 \FA_INST_0[1].FA_INST_1[242].FA_  ( .A(A[754]), .B(B[754]), .CI(
        C[754]), .S(S[754]), .CO(C[755]) );
  FA_269 \FA_INST_0[1].FA_INST_1[243].FA_  ( .A(A[755]), .B(B[755]), .CI(
        C[755]), .S(S[755]), .CO(C[756]) );
  FA_268 \FA_INST_0[1].FA_INST_1[244].FA_  ( .A(A[756]), .B(B[756]), .CI(
        C[756]), .S(S[756]), .CO(C[757]) );
  FA_267 \FA_INST_0[1].FA_INST_1[245].FA_  ( .A(A[757]), .B(B[757]), .CI(
        C[757]), .S(S[757]), .CO(C[758]) );
  FA_266 \FA_INST_0[1].FA_INST_1[246].FA_  ( .A(A[758]), .B(B[758]), .CI(
        C[758]), .S(S[758]), .CO(C[759]) );
  FA_265 \FA_INST_0[1].FA_INST_1[247].FA_  ( .A(A[759]), .B(B[759]), .CI(
        C[759]), .S(S[759]), .CO(C[760]) );
  FA_264 \FA_INST_0[1].FA_INST_1[248].FA_  ( .A(A[760]), .B(B[760]), .CI(
        C[760]), .S(S[760]), .CO(C[761]) );
  FA_263 \FA_INST_0[1].FA_INST_1[249].FA_  ( .A(A[761]), .B(B[761]), .CI(
        C[761]), .S(S[761]), .CO(C[762]) );
  FA_262 \FA_INST_0[1].FA_INST_1[250].FA_  ( .A(A[762]), .B(B[762]), .CI(
        C[762]), .S(S[762]), .CO(C[763]) );
  FA_261 \FA_INST_0[1].FA_INST_1[251].FA_  ( .A(A[763]), .B(B[763]), .CI(
        C[763]), .S(S[763]), .CO(C[764]) );
  FA_260 \FA_INST_0[1].FA_INST_1[252].FA_  ( .A(A[764]), .B(B[764]), .CI(
        C[764]), .S(S[764]), .CO(C[765]) );
  FA_259 \FA_INST_0[1].FA_INST_1[253].FA_  ( .A(A[765]), .B(B[765]), .CI(
        C[765]), .S(S[765]), .CO(C[766]) );
  FA_258 \FA_INST_0[1].FA_INST_1[254].FA_  ( .A(A[766]), .B(B[766]), .CI(
        C[766]), .S(S[766]), .CO(C[767]) );
  FA_257 \FA_INST_0[1].FA_INST_1[255].FA_  ( .A(A[767]), .B(B[767]), .CI(
        C[767]), .S(S[767]), .CO(C[768]) );
  FA_256 \FA_INST_0[1].FA_INST_1[256].FA_  ( .A(A[768]), .B(B[768]), .CI(
        C[768]), .S(S[768]), .CO(C[769]) );
  FA_255 \FA_INST_0[1].FA_INST_1[257].FA_  ( .A(A[769]), .B(B[769]), .CI(
        C[769]), .S(S[769]), .CO(C[770]) );
  FA_254 \FA_INST_0[1].FA_INST_1[258].FA_  ( .A(A[770]), .B(B[770]), .CI(
        C[770]), .S(S[770]), .CO(C[771]) );
  FA_253 \FA_INST_0[1].FA_INST_1[259].FA_  ( .A(A[771]), .B(B[771]), .CI(
        C[771]), .S(S[771]), .CO(C[772]) );
  FA_252 \FA_INST_0[1].FA_INST_1[260].FA_  ( .A(A[772]), .B(B[772]), .CI(
        C[772]), .S(S[772]), .CO(C[773]) );
  FA_251 \FA_INST_0[1].FA_INST_1[261].FA_  ( .A(A[773]), .B(B[773]), .CI(
        C[773]), .S(S[773]), .CO(C[774]) );
  FA_250 \FA_INST_0[1].FA_INST_1[262].FA_  ( .A(A[774]), .B(B[774]), .CI(
        C[774]), .S(S[774]), .CO(C[775]) );
  FA_249 \FA_INST_0[1].FA_INST_1[263].FA_  ( .A(A[775]), .B(B[775]), .CI(
        C[775]), .S(S[775]), .CO(C[776]) );
  FA_248 \FA_INST_0[1].FA_INST_1[264].FA_  ( .A(A[776]), .B(B[776]), .CI(
        C[776]), .S(S[776]), .CO(C[777]) );
  FA_247 \FA_INST_0[1].FA_INST_1[265].FA_  ( .A(A[777]), .B(B[777]), .CI(
        C[777]), .S(S[777]), .CO(C[778]) );
  FA_246 \FA_INST_0[1].FA_INST_1[266].FA_  ( .A(A[778]), .B(B[778]), .CI(
        C[778]), .S(S[778]), .CO(C[779]) );
  FA_245 \FA_INST_0[1].FA_INST_1[267].FA_  ( .A(A[779]), .B(B[779]), .CI(
        C[779]), .S(S[779]), .CO(C[780]) );
  FA_244 \FA_INST_0[1].FA_INST_1[268].FA_  ( .A(A[780]), .B(B[780]), .CI(
        C[780]), .S(S[780]), .CO(C[781]) );
  FA_243 \FA_INST_0[1].FA_INST_1[269].FA_  ( .A(A[781]), .B(B[781]), .CI(
        C[781]), .S(S[781]), .CO(C[782]) );
  FA_242 \FA_INST_0[1].FA_INST_1[270].FA_  ( .A(A[782]), .B(B[782]), .CI(
        C[782]), .S(S[782]), .CO(C[783]) );
  FA_241 \FA_INST_0[1].FA_INST_1[271].FA_  ( .A(A[783]), .B(B[783]), .CI(
        C[783]), .S(S[783]), .CO(C[784]) );
  FA_240 \FA_INST_0[1].FA_INST_1[272].FA_  ( .A(A[784]), .B(B[784]), .CI(
        C[784]), .S(S[784]), .CO(C[785]) );
  FA_239 \FA_INST_0[1].FA_INST_1[273].FA_  ( .A(A[785]), .B(B[785]), .CI(
        C[785]), .S(S[785]), .CO(C[786]) );
  FA_238 \FA_INST_0[1].FA_INST_1[274].FA_  ( .A(A[786]), .B(B[786]), .CI(
        C[786]), .S(S[786]), .CO(C[787]) );
  FA_237 \FA_INST_0[1].FA_INST_1[275].FA_  ( .A(A[787]), .B(B[787]), .CI(
        C[787]), .S(S[787]), .CO(C[788]) );
  FA_236 \FA_INST_0[1].FA_INST_1[276].FA_  ( .A(A[788]), .B(B[788]), .CI(
        C[788]), .S(S[788]), .CO(C[789]) );
  FA_235 \FA_INST_0[1].FA_INST_1[277].FA_  ( .A(A[789]), .B(B[789]), .CI(
        C[789]), .S(S[789]), .CO(C[790]) );
  FA_234 \FA_INST_0[1].FA_INST_1[278].FA_  ( .A(A[790]), .B(B[790]), .CI(
        C[790]), .S(S[790]), .CO(C[791]) );
  FA_233 \FA_INST_0[1].FA_INST_1[279].FA_  ( .A(A[791]), .B(B[791]), .CI(
        C[791]), .S(S[791]), .CO(C[792]) );
  FA_232 \FA_INST_0[1].FA_INST_1[280].FA_  ( .A(A[792]), .B(B[792]), .CI(
        C[792]), .S(S[792]), .CO(C[793]) );
  FA_231 \FA_INST_0[1].FA_INST_1[281].FA_  ( .A(A[793]), .B(B[793]), .CI(
        C[793]), .S(S[793]), .CO(C[794]) );
  FA_230 \FA_INST_0[1].FA_INST_1[282].FA_  ( .A(A[794]), .B(B[794]), .CI(
        C[794]), .S(S[794]), .CO(C[795]) );
  FA_229 \FA_INST_0[1].FA_INST_1[283].FA_  ( .A(A[795]), .B(B[795]), .CI(
        C[795]), .S(S[795]), .CO(C[796]) );
  FA_228 \FA_INST_0[1].FA_INST_1[284].FA_  ( .A(A[796]), .B(B[796]), .CI(
        C[796]), .S(S[796]), .CO(C[797]) );
  FA_227 \FA_INST_0[1].FA_INST_1[285].FA_  ( .A(A[797]), .B(B[797]), .CI(
        C[797]), .S(S[797]), .CO(C[798]) );
  FA_226 \FA_INST_0[1].FA_INST_1[286].FA_  ( .A(A[798]), .B(B[798]), .CI(
        C[798]), .S(S[798]), .CO(C[799]) );
  FA_225 \FA_INST_0[1].FA_INST_1[287].FA_  ( .A(A[799]), .B(B[799]), .CI(
        C[799]), .S(S[799]), .CO(C[800]) );
  FA_224 \FA_INST_0[1].FA_INST_1[288].FA_  ( .A(A[800]), .B(B[800]), .CI(
        C[800]), .S(S[800]), .CO(C[801]) );
  FA_223 \FA_INST_0[1].FA_INST_1[289].FA_  ( .A(A[801]), .B(B[801]), .CI(
        C[801]), .S(S[801]), .CO(C[802]) );
  FA_222 \FA_INST_0[1].FA_INST_1[290].FA_  ( .A(A[802]), .B(B[802]), .CI(
        C[802]), .S(S[802]), .CO(C[803]) );
  FA_221 \FA_INST_0[1].FA_INST_1[291].FA_  ( .A(A[803]), .B(B[803]), .CI(
        C[803]), .S(S[803]), .CO(C[804]) );
  FA_220 \FA_INST_0[1].FA_INST_1[292].FA_  ( .A(A[804]), .B(B[804]), .CI(
        C[804]), .S(S[804]), .CO(C[805]) );
  FA_219 \FA_INST_0[1].FA_INST_1[293].FA_  ( .A(A[805]), .B(B[805]), .CI(
        C[805]), .S(S[805]), .CO(C[806]) );
  FA_218 \FA_INST_0[1].FA_INST_1[294].FA_  ( .A(A[806]), .B(B[806]), .CI(
        C[806]), .S(S[806]), .CO(C[807]) );
  FA_217 \FA_INST_0[1].FA_INST_1[295].FA_  ( .A(A[807]), .B(B[807]), .CI(
        C[807]), .S(S[807]), .CO(C[808]) );
  FA_216 \FA_INST_0[1].FA_INST_1[296].FA_  ( .A(A[808]), .B(B[808]), .CI(
        C[808]), .S(S[808]), .CO(C[809]) );
  FA_215 \FA_INST_0[1].FA_INST_1[297].FA_  ( .A(A[809]), .B(B[809]), .CI(
        C[809]), .S(S[809]), .CO(C[810]) );
  FA_214 \FA_INST_0[1].FA_INST_1[298].FA_  ( .A(A[810]), .B(B[810]), .CI(
        C[810]), .S(S[810]), .CO(C[811]) );
  FA_213 \FA_INST_0[1].FA_INST_1[299].FA_  ( .A(A[811]), .B(B[811]), .CI(
        C[811]), .S(S[811]), .CO(C[812]) );
  FA_212 \FA_INST_0[1].FA_INST_1[300].FA_  ( .A(A[812]), .B(B[812]), .CI(
        C[812]), .S(S[812]), .CO(C[813]) );
  FA_211 \FA_INST_0[1].FA_INST_1[301].FA_  ( .A(A[813]), .B(B[813]), .CI(
        C[813]), .S(S[813]), .CO(C[814]) );
  FA_210 \FA_INST_0[1].FA_INST_1[302].FA_  ( .A(A[814]), .B(B[814]), .CI(
        C[814]), .S(S[814]), .CO(C[815]) );
  FA_209 \FA_INST_0[1].FA_INST_1[303].FA_  ( .A(A[815]), .B(B[815]), .CI(
        C[815]), .S(S[815]), .CO(C[816]) );
  FA_208 \FA_INST_0[1].FA_INST_1[304].FA_  ( .A(A[816]), .B(B[816]), .CI(
        C[816]), .S(S[816]), .CO(C[817]) );
  FA_207 \FA_INST_0[1].FA_INST_1[305].FA_  ( .A(A[817]), .B(B[817]), .CI(
        C[817]), .S(S[817]), .CO(C[818]) );
  FA_206 \FA_INST_0[1].FA_INST_1[306].FA_  ( .A(A[818]), .B(B[818]), .CI(
        C[818]), .S(S[818]), .CO(C[819]) );
  FA_205 \FA_INST_0[1].FA_INST_1[307].FA_  ( .A(A[819]), .B(B[819]), .CI(
        C[819]), .S(S[819]), .CO(C[820]) );
  FA_204 \FA_INST_0[1].FA_INST_1[308].FA_  ( .A(A[820]), .B(B[820]), .CI(
        C[820]), .S(S[820]), .CO(C[821]) );
  FA_203 \FA_INST_0[1].FA_INST_1[309].FA_  ( .A(A[821]), .B(B[821]), .CI(
        C[821]), .S(S[821]), .CO(C[822]) );
  FA_202 \FA_INST_0[1].FA_INST_1[310].FA_  ( .A(A[822]), .B(B[822]), .CI(
        C[822]), .S(S[822]), .CO(C[823]) );
  FA_201 \FA_INST_0[1].FA_INST_1[311].FA_  ( .A(A[823]), .B(B[823]), .CI(
        C[823]), .S(S[823]), .CO(C[824]) );
  FA_200 \FA_INST_0[1].FA_INST_1[312].FA_  ( .A(A[824]), .B(B[824]), .CI(
        C[824]), .S(S[824]), .CO(C[825]) );
  FA_199 \FA_INST_0[1].FA_INST_1[313].FA_  ( .A(A[825]), .B(B[825]), .CI(
        C[825]), .S(S[825]), .CO(C[826]) );
  FA_198 \FA_INST_0[1].FA_INST_1[314].FA_  ( .A(A[826]), .B(B[826]), .CI(
        C[826]), .S(S[826]), .CO(C[827]) );
  FA_197 \FA_INST_0[1].FA_INST_1[315].FA_  ( .A(A[827]), .B(B[827]), .CI(
        C[827]), .S(S[827]), .CO(C[828]) );
  FA_196 \FA_INST_0[1].FA_INST_1[316].FA_  ( .A(A[828]), .B(B[828]), .CI(
        C[828]), .S(S[828]), .CO(C[829]) );
  FA_195 \FA_INST_0[1].FA_INST_1[317].FA_  ( .A(A[829]), .B(B[829]), .CI(
        C[829]), .S(S[829]), .CO(C[830]) );
  FA_194 \FA_INST_0[1].FA_INST_1[318].FA_  ( .A(A[830]), .B(B[830]), .CI(
        C[830]), .S(S[830]), .CO(C[831]) );
  FA_193 \FA_INST_0[1].FA_INST_1[319].FA_  ( .A(A[831]), .B(B[831]), .CI(
        C[831]), .S(S[831]), .CO(C[832]) );
  FA_192 \FA_INST_0[1].FA_INST_1[320].FA_  ( .A(A[832]), .B(B[832]), .CI(
        C[832]), .S(S[832]), .CO(C[833]) );
  FA_191 \FA_INST_0[1].FA_INST_1[321].FA_  ( .A(A[833]), .B(B[833]), .CI(
        C[833]), .S(S[833]), .CO(C[834]) );
  FA_190 \FA_INST_0[1].FA_INST_1[322].FA_  ( .A(A[834]), .B(B[834]), .CI(
        C[834]), .S(S[834]), .CO(C[835]) );
  FA_189 \FA_INST_0[1].FA_INST_1[323].FA_  ( .A(A[835]), .B(B[835]), .CI(
        C[835]), .S(S[835]), .CO(C[836]) );
  FA_188 \FA_INST_0[1].FA_INST_1[324].FA_  ( .A(A[836]), .B(B[836]), .CI(
        C[836]), .S(S[836]), .CO(C[837]) );
  FA_187 \FA_INST_0[1].FA_INST_1[325].FA_  ( .A(A[837]), .B(B[837]), .CI(
        C[837]), .S(S[837]), .CO(C[838]) );
  FA_186 \FA_INST_0[1].FA_INST_1[326].FA_  ( .A(A[838]), .B(B[838]), .CI(
        C[838]), .S(S[838]), .CO(C[839]) );
  FA_185 \FA_INST_0[1].FA_INST_1[327].FA_  ( .A(A[839]), .B(B[839]), .CI(
        C[839]), .S(S[839]), .CO(C[840]) );
  FA_184 \FA_INST_0[1].FA_INST_1[328].FA_  ( .A(A[840]), .B(B[840]), .CI(
        C[840]), .S(S[840]), .CO(C[841]) );
  FA_183 \FA_INST_0[1].FA_INST_1[329].FA_  ( .A(A[841]), .B(B[841]), .CI(
        C[841]), .S(S[841]), .CO(C[842]) );
  FA_182 \FA_INST_0[1].FA_INST_1[330].FA_  ( .A(A[842]), .B(B[842]), .CI(
        C[842]), .S(S[842]), .CO(C[843]) );
  FA_181 \FA_INST_0[1].FA_INST_1[331].FA_  ( .A(A[843]), .B(B[843]), .CI(
        C[843]), .S(S[843]), .CO(C[844]) );
  FA_180 \FA_INST_0[1].FA_INST_1[332].FA_  ( .A(A[844]), .B(B[844]), .CI(
        C[844]), .S(S[844]), .CO(C[845]) );
  FA_179 \FA_INST_0[1].FA_INST_1[333].FA_  ( .A(A[845]), .B(B[845]), .CI(
        C[845]), .S(S[845]), .CO(C[846]) );
  FA_178 \FA_INST_0[1].FA_INST_1[334].FA_  ( .A(A[846]), .B(B[846]), .CI(
        C[846]), .S(S[846]), .CO(C[847]) );
  FA_177 \FA_INST_0[1].FA_INST_1[335].FA_  ( .A(A[847]), .B(B[847]), .CI(
        C[847]), .S(S[847]), .CO(C[848]) );
  FA_176 \FA_INST_0[1].FA_INST_1[336].FA_  ( .A(A[848]), .B(B[848]), .CI(
        C[848]), .S(S[848]), .CO(C[849]) );
  FA_175 \FA_INST_0[1].FA_INST_1[337].FA_  ( .A(A[849]), .B(B[849]), .CI(
        C[849]), .S(S[849]), .CO(C[850]) );
  FA_174 \FA_INST_0[1].FA_INST_1[338].FA_  ( .A(A[850]), .B(B[850]), .CI(
        C[850]), .S(S[850]), .CO(C[851]) );
  FA_173 \FA_INST_0[1].FA_INST_1[339].FA_  ( .A(A[851]), .B(B[851]), .CI(
        C[851]), .S(S[851]), .CO(C[852]) );
  FA_172 \FA_INST_0[1].FA_INST_1[340].FA_  ( .A(A[852]), .B(B[852]), .CI(
        C[852]), .S(S[852]), .CO(C[853]) );
  FA_171 \FA_INST_0[1].FA_INST_1[341].FA_  ( .A(A[853]), .B(B[853]), .CI(
        C[853]), .S(S[853]), .CO(C[854]) );
  FA_170 \FA_INST_0[1].FA_INST_1[342].FA_  ( .A(A[854]), .B(B[854]), .CI(
        C[854]), .S(S[854]), .CO(C[855]) );
  FA_169 \FA_INST_0[1].FA_INST_1[343].FA_  ( .A(A[855]), .B(B[855]), .CI(
        C[855]), .S(S[855]), .CO(C[856]) );
  FA_168 \FA_INST_0[1].FA_INST_1[344].FA_  ( .A(A[856]), .B(B[856]), .CI(
        C[856]), .S(S[856]), .CO(C[857]) );
  FA_167 \FA_INST_0[1].FA_INST_1[345].FA_  ( .A(A[857]), .B(B[857]), .CI(
        C[857]), .S(S[857]), .CO(C[858]) );
  FA_166 \FA_INST_0[1].FA_INST_1[346].FA_  ( .A(A[858]), .B(B[858]), .CI(
        C[858]), .S(S[858]), .CO(C[859]) );
  FA_165 \FA_INST_0[1].FA_INST_1[347].FA_  ( .A(A[859]), .B(B[859]), .CI(
        C[859]), .S(S[859]), .CO(C[860]) );
  FA_164 \FA_INST_0[1].FA_INST_1[348].FA_  ( .A(A[860]), .B(B[860]), .CI(
        C[860]), .S(S[860]), .CO(C[861]) );
  FA_163 \FA_INST_0[1].FA_INST_1[349].FA_  ( .A(A[861]), .B(B[861]), .CI(
        C[861]), .S(S[861]), .CO(C[862]) );
  FA_162 \FA_INST_0[1].FA_INST_1[350].FA_  ( .A(A[862]), .B(B[862]), .CI(
        C[862]), .S(S[862]), .CO(C[863]) );
  FA_161 \FA_INST_0[1].FA_INST_1[351].FA_  ( .A(A[863]), .B(B[863]), .CI(
        C[863]), .S(S[863]), .CO(C[864]) );
  FA_160 \FA_INST_0[1].FA_INST_1[352].FA_  ( .A(A[864]), .B(B[864]), .CI(
        C[864]), .S(S[864]), .CO(C[865]) );
  FA_159 \FA_INST_0[1].FA_INST_1[353].FA_  ( .A(A[865]), .B(B[865]), .CI(
        C[865]), .S(S[865]), .CO(C[866]) );
  FA_158 \FA_INST_0[1].FA_INST_1[354].FA_  ( .A(A[866]), .B(B[866]), .CI(
        C[866]), .S(S[866]), .CO(C[867]) );
  FA_157 \FA_INST_0[1].FA_INST_1[355].FA_  ( .A(A[867]), .B(B[867]), .CI(
        C[867]), .S(S[867]), .CO(C[868]) );
  FA_156 \FA_INST_0[1].FA_INST_1[356].FA_  ( .A(A[868]), .B(B[868]), .CI(
        C[868]), .S(S[868]), .CO(C[869]) );
  FA_155 \FA_INST_0[1].FA_INST_1[357].FA_  ( .A(A[869]), .B(B[869]), .CI(
        C[869]), .S(S[869]), .CO(C[870]) );
  FA_154 \FA_INST_0[1].FA_INST_1[358].FA_  ( .A(A[870]), .B(B[870]), .CI(
        C[870]), .S(S[870]), .CO(C[871]) );
  FA_153 \FA_INST_0[1].FA_INST_1[359].FA_  ( .A(A[871]), .B(B[871]), .CI(
        C[871]), .S(S[871]), .CO(C[872]) );
  FA_152 \FA_INST_0[1].FA_INST_1[360].FA_  ( .A(A[872]), .B(B[872]), .CI(
        C[872]), .S(S[872]), .CO(C[873]) );
  FA_151 \FA_INST_0[1].FA_INST_1[361].FA_  ( .A(A[873]), .B(B[873]), .CI(
        C[873]), .S(S[873]), .CO(C[874]) );
  FA_150 \FA_INST_0[1].FA_INST_1[362].FA_  ( .A(A[874]), .B(B[874]), .CI(
        C[874]), .S(S[874]), .CO(C[875]) );
  FA_149 \FA_INST_0[1].FA_INST_1[363].FA_  ( .A(A[875]), .B(B[875]), .CI(
        C[875]), .S(S[875]), .CO(C[876]) );
  FA_148 \FA_INST_0[1].FA_INST_1[364].FA_  ( .A(A[876]), .B(B[876]), .CI(
        C[876]), .S(S[876]), .CO(C[877]) );
  FA_147 \FA_INST_0[1].FA_INST_1[365].FA_  ( .A(A[877]), .B(B[877]), .CI(
        C[877]), .S(S[877]), .CO(C[878]) );
  FA_146 \FA_INST_0[1].FA_INST_1[366].FA_  ( .A(A[878]), .B(B[878]), .CI(
        C[878]), .S(S[878]), .CO(C[879]) );
  FA_145 \FA_INST_0[1].FA_INST_1[367].FA_  ( .A(A[879]), .B(B[879]), .CI(
        C[879]), .S(S[879]), .CO(C[880]) );
  FA_144 \FA_INST_0[1].FA_INST_1[368].FA_  ( .A(A[880]), .B(B[880]), .CI(
        C[880]), .S(S[880]), .CO(C[881]) );
  FA_143 \FA_INST_0[1].FA_INST_1[369].FA_  ( .A(A[881]), .B(B[881]), .CI(
        C[881]), .S(S[881]), .CO(C[882]) );
  FA_142 \FA_INST_0[1].FA_INST_1[370].FA_  ( .A(A[882]), .B(B[882]), .CI(
        C[882]), .S(S[882]), .CO(C[883]) );
  FA_141 \FA_INST_0[1].FA_INST_1[371].FA_  ( .A(A[883]), .B(B[883]), .CI(
        C[883]), .S(S[883]), .CO(C[884]) );
  FA_140 \FA_INST_0[1].FA_INST_1[372].FA_  ( .A(A[884]), .B(B[884]), .CI(
        C[884]), .S(S[884]), .CO(C[885]) );
  FA_139 \FA_INST_0[1].FA_INST_1[373].FA_  ( .A(A[885]), .B(B[885]), .CI(
        C[885]), .S(S[885]), .CO(C[886]) );
  FA_138 \FA_INST_0[1].FA_INST_1[374].FA_  ( .A(A[886]), .B(B[886]), .CI(
        C[886]), .S(S[886]), .CO(C[887]) );
  FA_137 \FA_INST_0[1].FA_INST_1[375].FA_  ( .A(A[887]), .B(B[887]), .CI(
        C[887]), .S(S[887]), .CO(C[888]) );
  FA_136 \FA_INST_0[1].FA_INST_1[376].FA_  ( .A(A[888]), .B(B[888]), .CI(
        C[888]), .S(S[888]), .CO(C[889]) );
  FA_135 \FA_INST_0[1].FA_INST_1[377].FA_  ( .A(A[889]), .B(B[889]), .CI(
        C[889]), .S(S[889]), .CO(C[890]) );
  FA_134 \FA_INST_0[1].FA_INST_1[378].FA_  ( .A(A[890]), .B(B[890]), .CI(
        C[890]), .S(S[890]), .CO(C[891]) );
  FA_133 \FA_INST_0[1].FA_INST_1[379].FA_  ( .A(A[891]), .B(B[891]), .CI(
        C[891]), .S(S[891]), .CO(C[892]) );
  FA_132 \FA_INST_0[1].FA_INST_1[380].FA_  ( .A(A[892]), .B(B[892]), .CI(
        C[892]), .S(S[892]), .CO(C[893]) );
  FA_131 \FA_INST_0[1].FA_INST_1[381].FA_  ( .A(A[893]), .B(B[893]), .CI(
        C[893]), .S(S[893]), .CO(C[894]) );
  FA_130 \FA_INST_0[1].FA_INST_1[382].FA_  ( .A(A[894]), .B(B[894]), .CI(
        C[894]), .S(S[894]), .CO(C[895]) );
  FA_129 \FA_INST_0[1].FA_INST_1[383].FA_  ( .A(A[895]), .B(B[895]), .CI(
        C[895]), .S(S[895]), .CO(C[896]) );
  FA_128 \FA_INST_0[1].FA_INST_1[384].FA_  ( .A(A[896]), .B(B[896]), .CI(
        C[896]), .S(S[896]), .CO(C[897]) );
  FA_127 \FA_INST_0[1].FA_INST_1[385].FA_  ( .A(A[897]), .B(B[897]), .CI(
        C[897]), .S(S[897]), .CO(C[898]) );
  FA_126 \FA_INST_0[1].FA_INST_1[386].FA_  ( .A(A[898]), .B(B[898]), .CI(
        C[898]), .S(S[898]), .CO(C[899]) );
  FA_125 \FA_INST_0[1].FA_INST_1[387].FA_  ( .A(A[899]), .B(B[899]), .CI(
        C[899]), .S(S[899]), .CO(C[900]) );
  FA_124 \FA_INST_0[1].FA_INST_1[388].FA_  ( .A(A[900]), .B(B[900]), .CI(
        C[900]), .S(S[900]), .CO(C[901]) );
  FA_123 \FA_INST_0[1].FA_INST_1[389].FA_  ( .A(A[901]), .B(B[901]), .CI(
        C[901]), .S(S[901]), .CO(C[902]) );
  FA_122 \FA_INST_0[1].FA_INST_1[390].FA_  ( .A(A[902]), .B(B[902]), .CI(
        C[902]), .S(S[902]), .CO(C[903]) );
  FA_121 \FA_INST_0[1].FA_INST_1[391].FA_  ( .A(A[903]), .B(B[903]), .CI(
        C[903]), .S(S[903]), .CO(C[904]) );
  FA_120 \FA_INST_0[1].FA_INST_1[392].FA_  ( .A(A[904]), .B(B[904]), .CI(
        C[904]), .S(S[904]), .CO(C[905]) );
  FA_119 \FA_INST_0[1].FA_INST_1[393].FA_  ( .A(A[905]), .B(B[905]), .CI(
        C[905]), .S(S[905]), .CO(C[906]) );
  FA_118 \FA_INST_0[1].FA_INST_1[394].FA_  ( .A(A[906]), .B(B[906]), .CI(
        C[906]), .S(S[906]), .CO(C[907]) );
  FA_117 \FA_INST_0[1].FA_INST_1[395].FA_  ( .A(A[907]), .B(B[907]), .CI(
        C[907]), .S(S[907]), .CO(C[908]) );
  FA_116 \FA_INST_0[1].FA_INST_1[396].FA_  ( .A(A[908]), .B(B[908]), .CI(
        C[908]), .S(S[908]), .CO(C[909]) );
  FA_115 \FA_INST_0[1].FA_INST_1[397].FA_  ( .A(A[909]), .B(B[909]), .CI(
        C[909]), .S(S[909]), .CO(C[910]) );
  FA_114 \FA_INST_0[1].FA_INST_1[398].FA_  ( .A(A[910]), .B(B[910]), .CI(
        C[910]), .S(S[910]), .CO(C[911]) );
  FA_113 \FA_INST_0[1].FA_INST_1[399].FA_  ( .A(A[911]), .B(B[911]), .CI(
        C[911]), .S(S[911]), .CO(C[912]) );
  FA_112 \FA_INST_0[1].FA_INST_1[400].FA_  ( .A(A[912]), .B(B[912]), .CI(
        C[912]), .S(S[912]), .CO(C[913]) );
  FA_111 \FA_INST_0[1].FA_INST_1[401].FA_  ( .A(A[913]), .B(B[913]), .CI(
        C[913]), .S(S[913]), .CO(C[914]) );
  FA_110 \FA_INST_0[1].FA_INST_1[402].FA_  ( .A(A[914]), .B(B[914]), .CI(
        C[914]), .S(S[914]), .CO(C[915]) );
  FA_109 \FA_INST_0[1].FA_INST_1[403].FA_  ( .A(A[915]), .B(B[915]), .CI(
        C[915]), .S(S[915]), .CO(C[916]) );
  FA_108 \FA_INST_0[1].FA_INST_1[404].FA_  ( .A(A[916]), .B(B[916]), .CI(
        C[916]), .S(S[916]), .CO(C[917]) );
  FA_107 \FA_INST_0[1].FA_INST_1[405].FA_  ( .A(A[917]), .B(B[917]), .CI(
        C[917]), .S(S[917]), .CO(C[918]) );
  FA_106 \FA_INST_0[1].FA_INST_1[406].FA_  ( .A(A[918]), .B(B[918]), .CI(
        C[918]), .S(S[918]), .CO(C[919]) );
  FA_105 \FA_INST_0[1].FA_INST_1[407].FA_  ( .A(A[919]), .B(B[919]), .CI(
        C[919]), .S(S[919]), .CO(C[920]) );
  FA_104 \FA_INST_0[1].FA_INST_1[408].FA_  ( .A(A[920]), .B(B[920]), .CI(
        C[920]), .S(S[920]), .CO(C[921]) );
  FA_103 \FA_INST_0[1].FA_INST_1[409].FA_  ( .A(A[921]), .B(B[921]), .CI(
        C[921]), .S(S[921]), .CO(C[922]) );
  FA_102 \FA_INST_0[1].FA_INST_1[410].FA_  ( .A(A[922]), .B(B[922]), .CI(
        C[922]), .S(S[922]), .CO(C[923]) );
  FA_101 \FA_INST_0[1].FA_INST_1[411].FA_  ( .A(A[923]), .B(B[923]), .CI(
        C[923]), .S(S[923]), .CO(C[924]) );
  FA_100 \FA_INST_0[1].FA_INST_1[412].FA_  ( .A(A[924]), .B(B[924]), .CI(
        C[924]), .S(S[924]), .CO(C[925]) );
  FA_99 \FA_INST_0[1].FA_INST_1[413].FA_  ( .A(A[925]), .B(B[925]), .CI(C[925]), .S(S[925]), .CO(C[926]) );
  FA_98 \FA_INST_0[1].FA_INST_1[414].FA_  ( .A(A[926]), .B(B[926]), .CI(C[926]), .S(S[926]), .CO(C[927]) );
  FA_97 \FA_INST_0[1].FA_INST_1[415].FA_  ( .A(A[927]), .B(B[927]), .CI(C[927]), .S(S[927]), .CO(C[928]) );
  FA_96 \FA_INST_0[1].FA_INST_1[416].FA_  ( .A(A[928]), .B(B[928]), .CI(C[928]), .S(S[928]), .CO(C[929]) );
  FA_95 \FA_INST_0[1].FA_INST_1[417].FA_  ( .A(A[929]), .B(B[929]), .CI(C[929]), .S(S[929]), .CO(C[930]) );
  FA_94 \FA_INST_0[1].FA_INST_1[418].FA_  ( .A(A[930]), .B(B[930]), .CI(C[930]), .S(S[930]), .CO(C[931]) );
  FA_93 \FA_INST_0[1].FA_INST_1[419].FA_  ( .A(A[931]), .B(B[931]), .CI(C[931]), .S(S[931]), .CO(C[932]) );
  FA_92 \FA_INST_0[1].FA_INST_1[420].FA_  ( .A(A[932]), .B(B[932]), .CI(C[932]), .S(S[932]), .CO(C[933]) );
  FA_91 \FA_INST_0[1].FA_INST_1[421].FA_  ( .A(A[933]), .B(B[933]), .CI(C[933]), .S(S[933]), .CO(C[934]) );
  FA_90 \FA_INST_0[1].FA_INST_1[422].FA_  ( .A(A[934]), .B(B[934]), .CI(C[934]), .S(S[934]), .CO(C[935]) );
  FA_89 \FA_INST_0[1].FA_INST_1[423].FA_  ( .A(A[935]), .B(B[935]), .CI(C[935]), .S(S[935]), .CO(C[936]) );
  FA_88 \FA_INST_0[1].FA_INST_1[424].FA_  ( .A(A[936]), .B(B[936]), .CI(C[936]), .S(S[936]), .CO(C[937]) );
  FA_87 \FA_INST_0[1].FA_INST_1[425].FA_  ( .A(A[937]), .B(B[937]), .CI(C[937]), .S(S[937]), .CO(C[938]) );
  FA_86 \FA_INST_0[1].FA_INST_1[426].FA_  ( .A(A[938]), .B(B[938]), .CI(C[938]), .S(S[938]), .CO(C[939]) );
  FA_85 \FA_INST_0[1].FA_INST_1[427].FA_  ( .A(A[939]), .B(B[939]), .CI(C[939]), .S(S[939]), .CO(C[940]) );
  FA_84 \FA_INST_0[1].FA_INST_1[428].FA_  ( .A(A[940]), .B(B[940]), .CI(C[940]), .S(S[940]), .CO(C[941]) );
  FA_83 \FA_INST_0[1].FA_INST_1[429].FA_  ( .A(A[941]), .B(B[941]), .CI(C[941]), .S(S[941]), .CO(C[942]) );
  FA_82 \FA_INST_0[1].FA_INST_1[430].FA_  ( .A(A[942]), .B(B[942]), .CI(C[942]), .S(S[942]), .CO(C[943]) );
  FA_81 \FA_INST_0[1].FA_INST_1[431].FA_  ( .A(A[943]), .B(B[943]), .CI(C[943]), .S(S[943]), .CO(C[944]) );
  FA_80 \FA_INST_0[1].FA_INST_1[432].FA_  ( .A(A[944]), .B(B[944]), .CI(C[944]), .S(S[944]), .CO(C[945]) );
  FA_79 \FA_INST_0[1].FA_INST_1[433].FA_  ( .A(A[945]), .B(B[945]), .CI(C[945]), .S(S[945]), .CO(C[946]) );
  FA_78 \FA_INST_0[1].FA_INST_1[434].FA_  ( .A(A[946]), .B(B[946]), .CI(C[946]), .S(S[946]), .CO(C[947]) );
  FA_77 \FA_INST_0[1].FA_INST_1[435].FA_  ( .A(A[947]), .B(B[947]), .CI(C[947]), .S(S[947]), .CO(C[948]) );
  FA_76 \FA_INST_0[1].FA_INST_1[436].FA_  ( .A(A[948]), .B(B[948]), .CI(C[948]), .S(S[948]), .CO(C[949]) );
  FA_75 \FA_INST_0[1].FA_INST_1[437].FA_  ( .A(A[949]), .B(B[949]), .CI(C[949]), .S(S[949]), .CO(C[950]) );
  FA_74 \FA_INST_0[1].FA_INST_1[438].FA_  ( .A(A[950]), .B(B[950]), .CI(C[950]), .S(S[950]), .CO(C[951]) );
  FA_73 \FA_INST_0[1].FA_INST_1[439].FA_  ( .A(A[951]), .B(B[951]), .CI(C[951]), .S(S[951]), .CO(C[952]) );
  FA_72 \FA_INST_0[1].FA_INST_1[440].FA_  ( .A(A[952]), .B(B[952]), .CI(C[952]), .S(S[952]), .CO(C[953]) );
  FA_71 \FA_INST_0[1].FA_INST_1[441].FA_  ( .A(A[953]), .B(B[953]), .CI(C[953]), .S(S[953]), .CO(C[954]) );
  FA_70 \FA_INST_0[1].FA_INST_1[442].FA_  ( .A(A[954]), .B(B[954]), .CI(C[954]), .S(S[954]), .CO(C[955]) );
  FA_69 \FA_INST_0[1].FA_INST_1[443].FA_  ( .A(A[955]), .B(B[955]), .CI(C[955]), .S(S[955]), .CO(C[956]) );
  FA_68 \FA_INST_0[1].FA_INST_1[444].FA_  ( .A(A[956]), .B(B[956]), .CI(C[956]), .S(S[956]), .CO(C[957]) );
  FA_67 \FA_INST_0[1].FA_INST_1[445].FA_  ( .A(A[957]), .B(B[957]), .CI(C[957]), .S(S[957]), .CO(C[958]) );
  FA_66 \FA_INST_0[1].FA_INST_1[446].FA_  ( .A(A[958]), .B(B[958]), .CI(C[958]), .S(S[958]), .CO(C[959]) );
  FA_65 \FA_INST_0[1].FA_INST_1[447].FA_  ( .A(A[959]), .B(B[959]), .CI(C[959]), .S(S[959]), .CO(C[960]) );
  FA_64 \FA_INST_0[1].FA_INST_1[448].FA_  ( .A(A[960]), .B(B[960]), .CI(C[960]), .S(S[960]), .CO(C[961]) );
  FA_63 \FA_INST_0[1].FA_INST_1[449].FA_  ( .A(A[961]), .B(B[961]), .CI(C[961]), .S(S[961]), .CO(C[962]) );
  FA_62 \FA_INST_0[1].FA_INST_1[450].FA_  ( .A(A[962]), .B(B[962]), .CI(C[962]), .S(S[962]), .CO(C[963]) );
  FA_61 \FA_INST_0[1].FA_INST_1[451].FA_  ( .A(A[963]), .B(B[963]), .CI(C[963]), .S(S[963]), .CO(C[964]) );
  FA_60 \FA_INST_0[1].FA_INST_1[452].FA_  ( .A(A[964]), .B(B[964]), .CI(C[964]), .S(S[964]), .CO(C[965]) );
  FA_59 \FA_INST_0[1].FA_INST_1[453].FA_  ( .A(A[965]), .B(B[965]), .CI(C[965]), .S(S[965]), .CO(C[966]) );
  FA_58 \FA_INST_0[1].FA_INST_1[454].FA_  ( .A(A[966]), .B(B[966]), .CI(C[966]), .S(S[966]), .CO(C[967]) );
  FA_57 \FA_INST_0[1].FA_INST_1[455].FA_  ( .A(A[967]), .B(B[967]), .CI(C[967]), .S(S[967]), .CO(C[968]) );
  FA_56 \FA_INST_0[1].FA_INST_1[456].FA_  ( .A(A[968]), .B(B[968]), .CI(C[968]), .S(S[968]), .CO(C[969]) );
  FA_55 \FA_INST_0[1].FA_INST_1[457].FA_  ( .A(A[969]), .B(B[969]), .CI(C[969]), .S(S[969]), .CO(C[970]) );
  FA_54 \FA_INST_0[1].FA_INST_1[458].FA_  ( .A(A[970]), .B(B[970]), .CI(C[970]), .S(S[970]), .CO(C[971]) );
  FA_53 \FA_INST_0[1].FA_INST_1[459].FA_  ( .A(A[971]), .B(B[971]), .CI(C[971]), .S(S[971]), .CO(C[972]) );
  FA_52 \FA_INST_0[1].FA_INST_1[460].FA_  ( .A(A[972]), .B(B[972]), .CI(C[972]), .S(S[972]), .CO(C[973]) );
  FA_51 \FA_INST_0[1].FA_INST_1[461].FA_  ( .A(A[973]), .B(B[973]), .CI(C[973]), .S(S[973]), .CO(C[974]) );
  FA_50 \FA_INST_0[1].FA_INST_1[462].FA_  ( .A(A[974]), .B(B[974]), .CI(C[974]), .S(S[974]), .CO(C[975]) );
  FA_49 \FA_INST_0[1].FA_INST_1[463].FA_  ( .A(A[975]), .B(B[975]), .CI(C[975]), .S(S[975]), .CO(C[976]) );
  FA_48 \FA_INST_0[1].FA_INST_1[464].FA_  ( .A(A[976]), .B(B[976]), .CI(C[976]), .S(S[976]), .CO(C[977]) );
  FA_47 \FA_INST_0[1].FA_INST_1[465].FA_  ( .A(A[977]), .B(B[977]), .CI(C[977]), .S(S[977]), .CO(C[978]) );
  FA_46 \FA_INST_0[1].FA_INST_1[466].FA_  ( .A(A[978]), .B(B[978]), .CI(C[978]), .S(S[978]), .CO(C[979]) );
  FA_45 \FA_INST_0[1].FA_INST_1[467].FA_  ( .A(A[979]), .B(B[979]), .CI(C[979]), .S(S[979]), .CO(C[980]) );
  FA_44 \FA_INST_0[1].FA_INST_1[468].FA_  ( .A(A[980]), .B(B[980]), .CI(C[980]), .S(S[980]), .CO(C[981]) );
  FA_43 \FA_INST_0[1].FA_INST_1[469].FA_  ( .A(A[981]), .B(B[981]), .CI(C[981]), .S(S[981]), .CO(C[982]) );
  FA_42 \FA_INST_0[1].FA_INST_1[470].FA_  ( .A(A[982]), .B(B[982]), .CI(C[982]), .S(S[982]), .CO(C[983]) );
  FA_41 \FA_INST_0[1].FA_INST_1[471].FA_  ( .A(A[983]), .B(B[983]), .CI(C[983]), .S(S[983]), .CO(C[984]) );
  FA_40 \FA_INST_0[1].FA_INST_1[472].FA_  ( .A(A[984]), .B(B[984]), .CI(C[984]), .S(S[984]), .CO(C[985]) );
  FA_39 \FA_INST_0[1].FA_INST_1[473].FA_  ( .A(A[985]), .B(B[985]), .CI(C[985]), .S(S[985]), .CO(C[986]) );
  FA_38 \FA_INST_0[1].FA_INST_1[474].FA_  ( .A(A[986]), .B(B[986]), .CI(C[986]), .S(S[986]), .CO(C[987]) );
  FA_37 \FA_INST_0[1].FA_INST_1[475].FA_  ( .A(A[987]), .B(B[987]), .CI(C[987]), .S(S[987]), .CO(C[988]) );
  FA_36 \FA_INST_0[1].FA_INST_1[476].FA_  ( .A(A[988]), .B(B[988]), .CI(C[988]), .S(S[988]), .CO(C[989]) );
  FA_35 \FA_INST_0[1].FA_INST_1[477].FA_  ( .A(A[989]), .B(B[989]), .CI(C[989]), .S(S[989]), .CO(C[990]) );
  FA_34 \FA_INST_0[1].FA_INST_1[478].FA_  ( .A(A[990]), .B(B[990]), .CI(C[990]), .S(S[990]), .CO(C[991]) );
  FA_33 \FA_INST_0[1].FA_INST_1[479].FA_  ( .A(A[991]), .B(B[991]), .CI(C[991]), .S(S[991]), .CO(C[992]) );
  FA_32 \FA_INST_0[1].FA_INST_1[480].FA_  ( .A(A[992]), .B(B[992]), .CI(C[992]), .S(S[992]), .CO(C[993]) );
  FA_31 \FA_INST_0[1].FA_INST_1[481].FA_  ( .A(A[993]), .B(B[993]), .CI(C[993]), .S(S[993]), .CO(C[994]) );
  FA_30 \FA_INST_0[1].FA_INST_1[482].FA_  ( .A(A[994]), .B(B[994]), .CI(C[994]), .S(S[994]), .CO(C[995]) );
  FA_29 \FA_INST_0[1].FA_INST_1[483].FA_  ( .A(A[995]), .B(B[995]), .CI(C[995]), .S(S[995]), .CO(C[996]) );
  FA_28 \FA_INST_0[1].FA_INST_1[484].FA_  ( .A(A[996]), .B(B[996]), .CI(C[996]), .S(S[996]), .CO(C[997]) );
  FA_27 \FA_INST_0[1].FA_INST_1[485].FA_  ( .A(A[997]), .B(B[997]), .CI(C[997]), .S(S[997]), .CO(C[998]) );
  FA_26 \FA_INST_0[1].FA_INST_1[486].FA_  ( .A(A[998]), .B(B[998]), .CI(C[998]), .S(S[998]), .CO(C[999]) );
  FA_25 \FA_INST_0[1].FA_INST_1[487].FA_  ( .A(A[999]), .B(B[999]), .CI(C[999]), .S(S[999]), .CO(C[1000]) );
  FA_24 \FA_INST_0[1].FA_INST_1[488].FA_  ( .A(A[1000]), .B(B[1000]), .CI(
        C[1000]), .S(S[1000]), .CO(C[1001]) );
  FA_23 \FA_INST_0[1].FA_INST_1[489].FA_  ( .A(A[1001]), .B(B[1001]), .CI(
        C[1001]), .S(S[1001]), .CO(C[1002]) );
  FA_22 \FA_INST_0[1].FA_INST_1[490].FA_  ( .A(A[1002]), .B(B[1002]), .CI(
        C[1002]), .S(S[1002]), .CO(C[1003]) );
  FA_21 \FA_INST_0[1].FA_INST_1[491].FA_  ( .A(A[1003]), .B(B[1003]), .CI(
        C[1003]), .S(S[1003]), .CO(C[1004]) );
  FA_20 \FA_INST_0[1].FA_INST_1[492].FA_  ( .A(A[1004]), .B(B[1004]), .CI(
        C[1004]), .S(S[1004]), .CO(C[1005]) );
  FA_19 \FA_INST_0[1].FA_INST_1[493].FA_  ( .A(A[1005]), .B(B[1005]), .CI(
        C[1005]), .S(S[1005]), .CO(C[1006]) );
  FA_18 \FA_INST_0[1].FA_INST_1[494].FA_  ( .A(A[1006]), .B(B[1006]), .CI(
        C[1006]), .S(S[1006]), .CO(C[1007]) );
  FA_17 \FA_INST_0[1].FA_INST_1[495].FA_  ( .A(A[1007]), .B(B[1007]), .CI(
        C[1007]), .S(S[1007]), .CO(C[1008]) );
  FA_16 \FA_INST_0[1].FA_INST_1[496].FA_  ( .A(A[1008]), .B(B[1008]), .CI(
        C[1008]), .S(S[1008]), .CO(C[1009]) );
  FA_15 \FA_INST_0[1].FA_INST_1[497].FA_  ( .A(A[1009]), .B(B[1009]), .CI(
        C[1009]), .S(S[1009]), .CO(C[1010]) );
  FA_14 \FA_INST_0[1].FA_INST_1[498].FA_  ( .A(A[1010]), .B(B[1010]), .CI(
        C[1010]), .S(S[1010]), .CO(C[1011]) );
  FA_13 \FA_INST_0[1].FA_INST_1[499].FA_  ( .A(A[1011]), .B(B[1011]), .CI(
        C[1011]), .S(S[1011]), .CO(C[1012]) );
  FA_12 \FA_INST_0[1].FA_INST_1[500].FA_  ( .A(A[1012]), .B(B[1012]), .CI(
        C[1012]), .S(S[1012]), .CO(C[1013]) );
  FA_11 \FA_INST_0[1].FA_INST_1[501].FA_  ( .A(A[1013]), .B(B[1013]), .CI(
        C[1013]), .S(S[1013]), .CO(C[1014]) );
  FA_10 \FA_INST_0[1].FA_INST_1[502].FA_  ( .A(A[1014]), .B(B[1014]), .CI(
        C[1014]), .S(S[1014]), .CO(C[1015]) );
  FA_9 \FA_INST_0[1].FA_INST_1[503].FA_  ( .A(A[1015]), .B(B[1015]), .CI(
        C[1015]), .S(S[1015]), .CO(C[1016]) );
  FA_8 \FA_INST_0[1].FA_INST_1[504].FA_  ( .A(A[1016]), .B(B[1016]), .CI(
        C[1016]), .S(S[1016]), .CO(C[1017]) );
  FA_7 \FA_INST_0[1].FA_INST_1[505].FA_  ( .A(A[1017]), .B(B[1017]), .CI(
        C[1017]), .S(S[1017]), .CO(C[1018]) );
  FA_6 \FA_INST_0[1].FA_INST_1[506].FA_  ( .A(A[1018]), .B(B[1018]), .CI(
        C[1018]), .S(S[1018]), .CO(C[1019]) );
  FA_5 \FA_INST_0[1].FA_INST_1[507].FA_  ( .A(A[1019]), .B(B[1019]), .CI(
        C[1019]), .S(S[1019]), .CO(C[1020]) );
  FA_4 \FA_INST_0[1].FA_INST_1[508].FA_  ( .A(1'b0), .B(B[1020]), .CI(C[1020]), 
        .S(S[1020]), .CO(C[1021]) );
  FA_3 \FA_INST_0[1].FA_INST_1[509].FA_  ( .A(1'b0), .B(B[1021]), .CI(C[1021]), 
        .S(S[1021]), .CO(C[1022]) );
  FA_2 \FA_INST_0[1].FA_INST_1[510].FA_  ( .A(1'b0), .B(B[1022]), .CI(C[1022]), 
        .S(S[1022]), .CO(C[1023]) );
  FA_1 \FA_INST_0[1].FA_INST_1[511].FA_  ( .A(1'b0), .B(B[1023]), .CI(C[1023]), 
        .S(S[1023]) );
endmodule


module mult_N1024_CC256_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [1023:0] A;
  input [3:0] B;
  output [1027:0] PRODUCT;
  input TC;
  wire   \ab[1023][0] , \ab[1022][1] , \ab[1022][0] , \ab[1021][2] ,
         \ab[1021][1] , \ab[1021][0] , \ab[1020][3] , \ab[1020][2] ,
         \ab[1020][1] , \ab[1020][0] , \ab[1019][3] , \ab[1019][2] ,
         \ab[1019][1] , \ab[1019][0] , \ab[1018][3] , \ab[1018][2] ,
         \ab[1018][1] , \ab[1018][0] , \ab[1017][3] , \ab[1017][2] ,
         \ab[1017][1] , \ab[1017][0] , \ab[1016][3] , \ab[1016][2] ,
         \ab[1016][1] , \ab[1016][0] , \ab[1015][3] , \ab[1015][2] ,
         \ab[1015][1] , \ab[1015][0] , \ab[1014][3] , \ab[1014][2] ,
         \ab[1014][1] , \ab[1014][0] , \ab[1013][3] , \ab[1013][2] ,
         \ab[1013][1] , \ab[1013][0] , \ab[1012][3] , \ab[1012][2] ,
         \ab[1012][1] , \ab[1012][0] , \ab[1011][3] , \ab[1011][2] ,
         \ab[1011][1] , \ab[1011][0] , \ab[1010][3] , \ab[1010][2] ,
         \ab[1010][1] , \ab[1010][0] , \ab[1009][3] , \ab[1009][2] ,
         \ab[1009][1] , \ab[1009][0] , \ab[1008][3] , \ab[1008][2] ,
         \ab[1008][1] , \ab[1008][0] , \ab[1007][3] , \ab[1007][2] ,
         \ab[1007][1] , \ab[1007][0] , \ab[1006][3] , \ab[1006][2] ,
         \ab[1006][1] , \ab[1006][0] , \ab[1005][3] , \ab[1005][2] ,
         \ab[1005][1] , \ab[1005][0] , \ab[1004][3] , \ab[1004][2] ,
         \ab[1004][1] , \ab[1004][0] , \ab[1003][3] , \ab[1003][2] ,
         \ab[1003][1] , \ab[1003][0] , \ab[1002][3] , \ab[1002][2] ,
         \ab[1002][1] , \ab[1002][0] , \ab[1001][3] , \ab[1001][2] ,
         \ab[1001][1] , \ab[1001][0] , \ab[1000][3] , \ab[1000][2] ,
         \ab[1000][1] , \ab[1000][0] , \ab[999][3] , \ab[999][2] ,
         \ab[999][1] , \ab[999][0] , \ab[998][3] , \ab[998][2] , \ab[998][1] ,
         \ab[998][0] , \ab[997][3] , \ab[997][2] , \ab[997][1] , \ab[997][0] ,
         \ab[996][3] , \ab[996][2] , \ab[996][1] , \ab[996][0] , \ab[995][3] ,
         \ab[995][2] , \ab[995][1] , \ab[995][0] , \ab[994][3] , \ab[994][2] ,
         \ab[994][1] , \ab[994][0] , \ab[993][3] , \ab[993][2] , \ab[993][1] ,
         \ab[993][0] , \ab[992][3] , \ab[992][2] , \ab[992][1] , \ab[992][0] ,
         \ab[991][3] , \ab[991][2] , \ab[991][1] , \ab[991][0] , \ab[990][3] ,
         \ab[990][2] , \ab[990][1] , \ab[990][0] , \ab[989][3] , \ab[989][2] ,
         \ab[989][1] , \ab[989][0] , \ab[988][3] , \ab[988][2] , \ab[988][1] ,
         \ab[988][0] , \ab[987][3] , \ab[987][2] , \ab[987][1] , \ab[987][0] ,
         \ab[986][3] , \ab[986][2] , \ab[986][1] , \ab[986][0] , \ab[985][3] ,
         \ab[985][2] , \ab[985][1] , \ab[985][0] , \ab[984][3] , \ab[984][2] ,
         \ab[984][1] , \ab[984][0] , \ab[983][3] , \ab[983][2] , \ab[983][1] ,
         \ab[983][0] , \ab[982][3] , \ab[982][2] , \ab[982][1] , \ab[982][0] ,
         \ab[981][3] , \ab[981][2] , \ab[981][1] , \ab[981][0] , \ab[980][3] ,
         \ab[980][2] , \ab[980][1] , \ab[980][0] , \ab[979][3] , \ab[979][2] ,
         \ab[979][1] , \ab[979][0] , \ab[978][3] , \ab[978][2] , \ab[978][1] ,
         \ab[978][0] , \ab[977][3] , \ab[977][2] , \ab[977][1] , \ab[977][0] ,
         \ab[976][3] , \ab[976][2] , \ab[976][1] , \ab[976][0] , \ab[975][3] ,
         \ab[975][2] , \ab[975][1] , \ab[975][0] , \ab[974][3] , \ab[974][2] ,
         \ab[974][1] , \ab[974][0] , \ab[973][3] , \ab[973][2] , \ab[973][1] ,
         \ab[973][0] , \ab[972][3] , \ab[972][2] , \ab[972][1] , \ab[972][0] ,
         \ab[971][3] , \ab[971][2] , \ab[971][1] , \ab[971][0] , \ab[970][3] ,
         \ab[970][2] , \ab[970][1] , \ab[970][0] , \ab[969][3] , \ab[969][2] ,
         \ab[969][1] , \ab[969][0] , \ab[968][3] , \ab[968][2] , \ab[968][1] ,
         \ab[968][0] , \ab[967][3] , \ab[967][2] , \ab[967][1] , \ab[967][0] ,
         \ab[966][3] , \ab[966][2] , \ab[966][1] , \ab[966][0] , \ab[965][3] ,
         \ab[965][2] , \ab[965][1] , \ab[965][0] , \ab[964][3] , \ab[964][2] ,
         \ab[964][1] , \ab[964][0] , \ab[963][3] , \ab[963][2] , \ab[963][1] ,
         \ab[963][0] , \ab[962][3] , \ab[962][2] , \ab[962][1] , \ab[962][0] ,
         \ab[961][3] , \ab[961][2] , \ab[961][1] , \ab[961][0] , \ab[960][3] ,
         \ab[960][2] , \ab[960][1] , \ab[960][0] , \ab[959][3] , \ab[959][2] ,
         \ab[959][1] , \ab[959][0] , \ab[958][3] , \ab[958][2] , \ab[958][1] ,
         \ab[958][0] , \ab[957][3] , \ab[957][2] , \ab[957][1] , \ab[957][0] ,
         \ab[956][3] , \ab[956][2] , \ab[956][1] , \ab[956][0] , \ab[955][3] ,
         \ab[955][2] , \ab[955][1] , \ab[955][0] , \ab[954][3] , \ab[954][2] ,
         \ab[954][1] , \ab[954][0] , \ab[953][3] , \ab[953][2] , \ab[953][1] ,
         \ab[953][0] , \ab[952][3] , \ab[952][2] , \ab[952][1] , \ab[952][0] ,
         \ab[951][3] , \ab[951][2] , \ab[951][1] , \ab[951][0] , \ab[950][3] ,
         \ab[950][2] , \ab[950][1] , \ab[950][0] , \ab[949][3] , \ab[949][2] ,
         \ab[949][1] , \ab[949][0] , \ab[948][3] , \ab[948][2] , \ab[948][1] ,
         \ab[948][0] , \ab[947][3] , \ab[947][2] , \ab[947][1] , \ab[947][0] ,
         \ab[946][3] , \ab[946][2] , \ab[946][1] , \ab[946][0] , \ab[945][3] ,
         \ab[945][2] , \ab[945][1] , \ab[945][0] , \ab[944][3] , \ab[944][2] ,
         \ab[944][1] , \ab[944][0] , \ab[943][3] , \ab[943][2] , \ab[943][1] ,
         \ab[943][0] , \ab[942][3] , \ab[942][2] , \ab[942][1] , \ab[942][0] ,
         \ab[941][3] , \ab[941][2] , \ab[941][1] , \ab[941][0] , \ab[940][3] ,
         \ab[940][2] , \ab[940][1] , \ab[940][0] , \ab[939][3] , \ab[939][2] ,
         \ab[939][1] , \ab[939][0] , \ab[938][3] , \ab[938][2] , \ab[938][1] ,
         \ab[938][0] , \ab[937][3] , \ab[937][2] , \ab[937][1] , \ab[937][0] ,
         \ab[936][3] , \ab[936][2] , \ab[936][1] , \ab[936][0] , \ab[935][3] ,
         \ab[935][2] , \ab[935][1] , \ab[935][0] , \ab[934][3] , \ab[934][2] ,
         \ab[934][1] , \ab[934][0] , \ab[933][3] , \ab[933][2] , \ab[933][1] ,
         \ab[933][0] , \ab[932][3] , \ab[932][2] , \ab[932][1] , \ab[932][0] ,
         \ab[931][3] , \ab[931][2] , \ab[931][1] , \ab[931][0] , \ab[930][3] ,
         \ab[930][2] , \ab[930][1] , \ab[930][0] , \ab[929][3] , \ab[929][2] ,
         \ab[929][1] , \ab[929][0] , \ab[928][3] , \ab[928][2] , \ab[928][1] ,
         \ab[928][0] , \ab[927][3] , \ab[927][2] , \ab[927][1] , \ab[927][0] ,
         \ab[926][3] , \ab[926][2] , \ab[926][1] , \ab[926][0] , \ab[925][3] ,
         \ab[925][2] , \ab[925][1] , \ab[925][0] , \ab[924][3] , \ab[924][2] ,
         \ab[924][1] , \ab[924][0] , \ab[923][3] , \ab[923][2] , \ab[923][1] ,
         \ab[923][0] , \ab[922][3] , \ab[922][2] , \ab[922][1] , \ab[922][0] ,
         \ab[921][3] , \ab[921][2] , \ab[921][1] , \ab[921][0] , \ab[920][3] ,
         \ab[920][2] , \ab[920][1] , \ab[920][0] , \ab[919][3] , \ab[919][2] ,
         \ab[919][1] , \ab[919][0] , \ab[918][3] , \ab[918][2] , \ab[918][1] ,
         \ab[918][0] , \ab[917][3] , \ab[917][2] , \ab[917][1] , \ab[917][0] ,
         \ab[916][3] , \ab[916][2] , \ab[916][1] , \ab[916][0] , \ab[915][3] ,
         \ab[915][2] , \ab[915][1] , \ab[915][0] , \ab[914][3] , \ab[914][2] ,
         \ab[914][1] , \ab[914][0] , \ab[913][3] , \ab[913][2] , \ab[913][1] ,
         \ab[913][0] , \ab[912][3] , \ab[912][2] , \ab[912][1] , \ab[912][0] ,
         \ab[911][3] , \ab[911][2] , \ab[911][1] , \ab[911][0] , \ab[910][3] ,
         \ab[910][2] , \ab[910][1] , \ab[910][0] , \ab[909][3] , \ab[909][2] ,
         \ab[909][1] , \ab[909][0] , \ab[908][3] , \ab[908][2] , \ab[908][1] ,
         \ab[908][0] , \ab[907][3] , \ab[907][2] , \ab[907][1] , \ab[907][0] ,
         \ab[906][3] , \ab[906][2] , \ab[906][1] , \ab[906][0] , \ab[905][3] ,
         \ab[905][2] , \ab[905][1] , \ab[905][0] , \ab[904][3] , \ab[904][2] ,
         \ab[904][1] , \ab[904][0] , \ab[903][3] , \ab[903][2] , \ab[903][1] ,
         \ab[903][0] , \ab[902][3] , \ab[902][2] , \ab[902][1] , \ab[902][0] ,
         \ab[901][3] , \ab[901][2] , \ab[901][1] , \ab[901][0] , \ab[900][3] ,
         \ab[900][2] , \ab[900][1] , \ab[900][0] , \ab[899][3] , \ab[899][2] ,
         \ab[899][1] , \ab[899][0] , \ab[898][3] , \ab[898][2] , \ab[898][1] ,
         \ab[898][0] , \ab[897][3] , \ab[897][2] , \ab[897][1] , \ab[897][0] ,
         \ab[896][3] , \ab[896][2] , \ab[896][1] , \ab[896][0] , \ab[895][3] ,
         \ab[895][2] , \ab[895][1] , \ab[895][0] , \ab[894][3] , \ab[894][2] ,
         \ab[894][1] , \ab[894][0] , \ab[893][3] , \ab[893][2] , \ab[893][1] ,
         \ab[893][0] , \ab[892][3] , \ab[892][2] , \ab[892][1] , \ab[892][0] ,
         \ab[891][3] , \ab[891][2] , \ab[891][1] , \ab[891][0] , \ab[890][3] ,
         \ab[890][2] , \ab[890][1] , \ab[890][0] , \ab[889][3] , \ab[889][2] ,
         \ab[889][1] , \ab[889][0] , \ab[888][3] , \ab[888][2] , \ab[888][1] ,
         \ab[888][0] , \ab[887][3] , \ab[887][2] , \ab[887][1] , \ab[887][0] ,
         \ab[886][3] , \ab[886][2] , \ab[886][1] , \ab[886][0] , \ab[885][3] ,
         \ab[885][2] , \ab[885][1] , \ab[885][0] , \ab[884][3] , \ab[884][2] ,
         \ab[884][1] , \ab[884][0] , \ab[883][3] , \ab[883][2] , \ab[883][1] ,
         \ab[883][0] , \ab[882][3] , \ab[882][2] , \ab[882][1] , \ab[882][0] ,
         \ab[881][3] , \ab[881][2] , \ab[881][1] , \ab[881][0] , \ab[880][3] ,
         \ab[880][2] , \ab[880][1] , \ab[880][0] , \ab[879][3] , \ab[879][2] ,
         \ab[879][1] , \ab[879][0] , \ab[878][3] , \ab[878][2] , \ab[878][1] ,
         \ab[878][0] , \ab[877][3] , \ab[877][2] , \ab[877][1] , \ab[877][0] ,
         \ab[876][3] , \ab[876][2] , \ab[876][1] , \ab[876][0] , \ab[875][3] ,
         \ab[875][2] , \ab[875][1] , \ab[875][0] , \ab[874][3] , \ab[874][2] ,
         \ab[874][1] , \ab[874][0] , \ab[873][3] , \ab[873][2] , \ab[873][1] ,
         \ab[873][0] , \ab[872][3] , \ab[872][2] , \ab[872][1] , \ab[872][0] ,
         \ab[871][3] , \ab[871][2] , \ab[871][1] , \ab[871][0] , \ab[870][3] ,
         \ab[870][2] , \ab[870][1] , \ab[870][0] , \ab[869][3] , \ab[869][2] ,
         \ab[869][1] , \ab[869][0] , \ab[868][3] , \ab[868][2] , \ab[868][1] ,
         \ab[868][0] , \ab[867][3] , \ab[867][2] , \ab[867][1] , \ab[867][0] ,
         \ab[866][3] , \ab[866][2] , \ab[866][1] , \ab[866][0] , \ab[865][3] ,
         \ab[865][2] , \ab[865][1] , \ab[865][0] , \ab[864][3] , \ab[864][2] ,
         \ab[864][1] , \ab[864][0] , \ab[863][3] , \ab[863][2] , \ab[863][1] ,
         \ab[863][0] , \ab[862][3] , \ab[862][2] , \ab[862][1] , \ab[862][0] ,
         \ab[861][3] , \ab[861][2] , \ab[861][1] , \ab[861][0] , \ab[860][3] ,
         \ab[860][2] , \ab[860][1] , \ab[860][0] , \ab[859][3] , \ab[859][2] ,
         \ab[859][1] , \ab[859][0] , \ab[858][3] , \ab[858][2] , \ab[858][1] ,
         \ab[858][0] , \ab[857][3] , \ab[857][2] , \ab[857][1] , \ab[857][0] ,
         \ab[856][3] , \ab[856][2] , \ab[856][1] , \ab[856][0] , \ab[855][3] ,
         \ab[855][2] , \ab[855][1] , \ab[855][0] , \ab[854][3] , \ab[854][2] ,
         \ab[854][1] , \ab[854][0] , \ab[853][3] , \ab[853][2] , \ab[853][1] ,
         \ab[853][0] , \ab[852][3] , \ab[852][2] , \ab[852][1] , \ab[852][0] ,
         \ab[851][3] , \ab[851][2] , \ab[851][1] , \ab[851][0] , \ab[850][3] ,
         \ab[850][2] , \ab[850][1] , \ab[850][0] , \ab[849][3] , \ab[849][2] ,
         \ab[849][1] , \ab[849][0] , \ab[848][3] , \ab[848][2] , \ab[848][1] ,
         \ab[848][0] , \ab[847][3] , \ab[847][2] , \ab[847][1] , \ab[847][0] ,
         \ab[846][3] , \ab[846][2] , \ab[846][1] , \ab[846][0] , \ab[845][3] ,
         \ab[845][2] , \ab[845][1] , \ab[845][0] , \ab[844][3] , \ab[844][2] ,
         \ab[844][1] , \ab[844][0] , \ab[843][3] , \ab[843][2] , \ab[843][1] ,
         \ab[843][0] , \ab[842][3] , \ab[842][2] , \ab[842][1] , \ab[842][0] ,
         \ab[841][3] , \ab[841][2] , \ab[841][1] , \ab[841][0] , \ab[840][3] ,
         \ab[840][2] , \ab[840][1] , \ab[840][0] , \ab[839][3] , \ab[839][2] ,
         \ab[839][1] , \ab[839][0] , \ab[838][3] , \ab[838][2] , \ab[838][1] ,
         \ab[838][0] , \ab[837][3] , \ab[837][2] , \ab[837][1] , \ab[837][0] ,
         \ab[836][3] , \ab[836][2] , \ab[836][1] , \ab[836][0] , \ab[835][3] ,
         \ab[835][2] , \ab[835][1] , \ab[835][0] , \ab[834][3] , \ab[834][2] ,
         \ab[834][1] , \ab[834][0] , \ab[833][3] , \ab[833][2] , \ab[833][1] ,
         \ab[833][0] , \ab[832][3] , \ab[832][2] , \ab[832][1] , \ab[832][0] ,
         \ab[831][3] , \ab[831][2] , \ab[831][1] , \ab[831][0] , \ab[830][3] ,
         \ab[830][2] , \ab[830][1] , \ab[830][0] , \ab[829][3] , \ab[829][2] ,
         \ab[829][1] , \ab[829][0] , \ab[828][3] , \ab[828][2] , \ab[828][1] ,
         \ab[828][0] , \ab[827][3] , \ab[827][2] , \ab[827][1] , \ab[827][0] ,
         \ab[826][3] , \ab[826][2] , \ab[826][1] , \ab[826][0] , \ab[825][3] ,
         \ab[825][2] , \ab[825][1] , \ab[825][0] , \ab[824][3] , \ab[824][2] ,
         \ab[824][1] , \ab[824][0] , \ab[823][3] , \ab[823][2] , \ab[823][1] ,
         \ab[823][0] , \ab[822][3] , \ab[822][2] , \ab[822][1] , \ab[822][0] ,
         \ab[821][3] , \ab[821][2] , \ab[821][1] , \ab[821][0] , \ab[820][3] ,
         \ab[820][2] , \ab[820][1] , \ab[820][0] , \ab[819][3] , \ab[819][2] ,
         \ab[819][1] , \ab[819][0] , \ab[818][3] , \ab[818][2] , \ab[818][1] ,
         \ab[818][0] , \ab[817][3] , \ab[817][2] , \ab[817][1] , \ab[817][0] ,
         \ab[816][3] , \ab[816][2] , \ab[816][1] , \ab[816][0] , \ab[815][3] ,
         \ab[815][2] , \ab[815][1] , \ab[815][0] , \ab[814][3] , \ab[814][2] ,
         \ab[814][1] , \ab[814][0] , \ab[813][3] , \ab[813][2] , \ab[813][1] ,
         \ab[813][0] , \ab[812][3] , \ab[812][2] , \ab[812][1] , \ab[812][0] ,
         \ab[811][3] , \ab[811][2] , \ab[811][1] , \ab[811][0] , \ab[810][3] ,
         \ab[810][2] , \ab[810][1] , \ab[810][0] , \ab[809][3] , \ab[809][2] ,
         \ab[809][1] , \ab[809][0] , \ab[808][3] , \ab[808][2] , \ab[808][1] ,
         \ab[808][0] , \ab[807][3] , \ab[807][2] , \ab[807][1] , \ab[807][0] ,
         \ab[806][3] , \ab[806][2] , \ab[806][1] , \ab[806][0] , \ab[805][3] ,
         \ab[805][2] , \ab[805][1] , \ab[805][0] , \ab[804][3] , \ab[804][2] ,
         \ab[804][1] , \ab[804][0] , \ab[803][3] , \ab[803][2] , \ab[803][1] ,
         \ab[803][0] , \ab[802][3] , \ab[802][2] , \ab[802][1] , \ab[802][0] ,
         \ab[801][3] , \ab[801][2] , \ab[801][1] , \ab[801][0] , \ab[800][3] ,
         \ab[800][2] , \ab[800][1] , \ab[800][0] , \ab[799][3] , \ab[799][2] ,
         \ab[799][1] , \ab[799][0] , \ab[798][3] , \ab[798][2] , \ab[798][1] ,
         \ab[798][0] , \ab[797][3] , \ab[797][2] , \ab[797][1] , \ab[797][0] ,
         \ab[796][3] , \ab[796][2] , \ab[796][1] , \ab[796][0] , \ab[795][3] ,
         \ab[795][2] , \ab[795][1] , \ab[795][0] , \ab[794][3] , \ab[794][2] ,
         \ab[794][1] , \ab[794][0] , \ab[793][3] , \ab[793][2] , \ab[793][1] ,
         \ab[793][0] , \ab[792][3] , \ab[792][2] , \ab[792][1] , \ab[792][0] ,
         \ab[791][3] , \ab[791][2] , \ab[791][1] , \ab[791][0] , \ab[790][3] ,
         \ab[790][2] , \ab[790][1] , \ab[790][0] , \ab[789][3] , \ab[789][2] ,
         \ab[789][1] , \ab[789][0] , \ab[788][3] , \ab[788][2] , \ab[788][1] ,
         \ab[788][0] , \ab[787][3] , \ab[787][2] , \ab[787][1] , \ab[787][0] ,
         \ab[786][3] , \ab[786][2] , \ab[786][1] , \ab[786][0] , \ab[785][3] ,
         \ab[785][2] , \ab[785][1] , \ab[785][0] , \ab[784][3] , \ab[784][2] ,
         \ab[784][1] , \ab[784][0] , \ab[783][3] , \ab[783][2] , \ab[783][1] ,
         \ab[783][0] , \ab[782][3] , \ab[782][2] , \ab[782][1] , \ab[782][0] ,
         \ab[781][3] , \ab[781][2] , \ab[781][1] , \ab[781][0] , \ab[780][3] ,
         \ab[780][2] , \ab[780][1] , \ab[780][0] , \ab[779][3] , \ab[779][2] ,
         \ab[779][1] , \ab[779][0] , \ab[778][3] , \ab[778][2] , \ab[778][1] ,
         \ab[778][0] , \ab[777][3] , \ab[777][2] , \ab[777][1] , \ab[777][0] ,
         \ab[776][3] , \ab[776][2] , \ab[776][1] , \ab[776][0] , \ab[775][3] ,
         \ab[775][2] , \ab[775][1] , \ab[775][0] , \ab[774][3] , \ab[774][2] ,
         \ab[774][1] , \ab[774][0] , \ab[773][3] , \ab[773][2] , \ab[773][1] ,
         \ab[773][0] , \ab[772][3] , \ab[772][2] , \ab[772][1] , \ab[772][0] ,
         \ab[771][3] , \ab[771][2] , \ab[771][1] , \ab[771][0] , \ab[770][3] ,
         \ab[770][2] , \ab[770][1] , \ab[770][0] , \ab[769][3] , \ab[769][2] ,
         \ab[769][1] , \ab[769][0] , \ab[768][3] , \ab[768][2] , \ab[768][1] ,
         \ab[768][0] , \ab[767][3] , \ab[767][2] , \ab[767][1] , \ab[767][0] ,
         \ab[766][3] , \ab[766][2] , \ab[766][1] , \ab[766][0] , \ab[765][3] ,
         \ab[765][2] , \ab[765][1] , \ab[765][0] , \ab[764][3] , \ab[764][2] ,
         \ab[764][1] , \ab[764][0] , \ab[763][3] , \ab[763][2] , \ab[763][1] ,
         \ab[763][0] , \ab[762][3] , \ab[762][2] , \ab[762][1] , \ab[762][0] ,
         \ab[761][3] , \ab[761][2] , \ab[761][1] , \ab[761][0] , \ab[760][3] ,
         \ab[760][2] , \ab[760][1] , \ab[760][0] , \ab[759][3] , \ab[759][2] ,
         \ab[759][1] , \ab[759][0] , \ab[758][3] , \ab[758][2] , \ab[758][1] ,
         \ab[758][0] , \ab[757][3] , \ab[757][2] , \ab[757][1] , \ab[757][0] ,
         \ab[756][3] , \ab[756][2] , \ab[756][1] , \ab[756][0] , \ab[755][3] ,
         \ab[755][2] , \ab[755][1] , \ab[755][0] , \ab[754][3] , \ab[754][2] ,
         \ab[754][1] , \ab[754][0] , \ab[753][3] , \ab[753][2] , \ab[753][1] ,
         \ab[753][0] , \ab[752][3] , \ab[752][2] , \ab[752][1] , \ab[752][0] ,
         \ab[751][3] , \ab[751][2] , \ab[751][1] , \ab[751][0] , \ab[750][3] ,
         \ab[750][2] , \ab[750][1] , \ab[750][0] , \ab[749][3] , \ab[749][2] ,
         \ab[749][1] , \ab[749][0] , \ab[748][3] , \ab[748][2] , \ab[748][1] ,
         \ab[748][0] , \ab[747][3] , \ab[747][2] , \ab[747][1] , \ab[747][0] ,
         \ab[746][3] , \ab[746][2] , \ab[746][1] , \ab[746][0] , \ab[745][3] ,
         \ab[745][2] , \ab[745][1] , \ab[745][0] , \ab[744][3] , \ab[744][2] ,
         \ab[744][1] , \ab[744][0] , \ab[743][3] , \ab[743][2] , \ab[743][1] ,
         \ab[743][0] , \ab[742][3] , \ab[742][2] , \ab[742][1] , \ab[742][0] ,
         \ab[741][3] , \ab[741][2] , \ab[741][1] , \ab[741][0] , \ab[740][3] ,
         \ab[740][2] , \ab[740][1] , \ab[740][0] , \ab[739][3] , \ab[739][2] ,
         \ab[739][1] , \ab[739][0] , \ab[738][3] , \ab[738][2] , \ab[738][1] ,
         \ab[738][0] , \ab[737][3] , \ab[737][2] , \ab[737][1] , \ab[737][0] ,
         \ab[736][3] , \ab[736][2] , \ab[736][1] , \ab[736][0] , \ab[735][3] ,
         \ab[735][2] , \ab[735][1] , \ab[735][0] , \ab[734][3] , \ab[734][2] ,
         \ab[734][1] , \ab[734][0] , \ab[733][3] , \ab[733][2] , \ab[733][1] ,
         \ab[733][0] , \ab[732][3] , \ab[732][2] , \ab[732][1] , \ab[732][0] ,
         \ab[731][3] , \ab[731][2] , \ab[731][1] , \ab[731][0] , \ab[730][3] ,
         \ab[730][2] , \ab[730][1] , \ab[730][0] , \ab[729][3] , \ab[729][2] ,
         \ab[729][1] , \ab[729][0] , \ab[728][3] , \ab[728][2] , \ab[728][1] ,
         \ab[728][0] , \ab[727][3] , \ab[727][2] , \ab[727][1] , \ab[727][0] ,
         \ab[726][3] , \ab[726][2] , \ab[726][1] , \ab[726][0] , \ab[725][3] ,
         \ab[725][2] , \ab[725][1] , \ab[725][0] , \ab[724][3] , \ab[724][2] ,
         \ab[724][1] , \ab[724][0] , \ab[723][3] , \ab[723][2] , \ab[723][1] ,
         \ab[723][0] , \ab[722][3] , \ab[722][2] , \ab[722][1] , \ab[722][0] ,
         \ab[721][3] , \ab[721][2] , \ab[721][1] , \ab[721][0] , \ab[720][3] ,
         \ab[720][2] , \ab[720][1] , \ab[720][0] , \ab[719][3] , \ab[719][2] ,
         \ab[719][1] , \ab[719][0] , \ab[718][3] , \ab[718][2] , \ab[718][1] ,
         \ab[718][0] , \ab[717][3] , \ab[717][2] , \ab[717][1] , \ab[717][0] ,
         \ab[716][3] , \ab[716][2] , \ab[716][1] , \ab[716][0] , \ab[715][3] ,
         \ab[715][2] , \ab[715][1] , \ab[715][0] , \ab[714][3] , \ab[714][2] ,
         \ab[714][1] , \ab[714][0] , \ab[713][3] , \ab[713][2] , \ab[713][1] ,
         \ab[713][0] , \ab[712][3] , \ab[712][2] , \ab[712][1] , \ab[712][0] ,
         \ab[711][3] , \ab[711][2] , \ab[711][1] , \ab[711][0] , \ab[710][3] ,
         \ab[710][2] , \ab[710][1] , \ab[710][0] , \ab[709][3] , \ab[709][2] ,
         \ab[709][1] , \ab[709][0] , \ab[708][3] , \ab[708][2] , \ab[708][1] ,
         \ab[708][0] , \ab[707][3] , \ab[707][2] , \ab[707][1] , \ab[707][0] ,
         \ab[706][3] , \ab[706][2] , \ab[706][1] , \ab[706][0] , \ab[705][3] ,
         \ab[705][2] , \ab[705][1] , \ab[705][0] , \ab[704][3] , \ab[704][2] ,
         \ab[704][1] , \ab[704][0] , \ab[703][3] , \ab[703][2] , \ab[703][1] ,
         \ab[703][0] , \ab[702][3] , \ab[702][2] , \ab[702][1] , \ab[702][0] ,
         \ab[701][3] , \ab[701][2] , \ab[701][1] , \ab[701][0] , \ab[700][3] ,
         \ab[700][2] , \ab[700][1] , \ab[700][0] , \ab[699][3] , \ab[699][2] ,
         \ab[699][1] , \ab[699][0] , \ab[698][3] , \ab[698][2] , \ab[698][1] ,
         \ab[698][0] , \ab[697][3] , \ab[697][2] , \ab[697][1] , \ab[697][0] ,
         \ab[696][3] , \ab[696][2] , \ab[696][1] , \ab[696][0] , \ab[695][3] ,
         \ab[695][2] , \ab[695][1] , \ab[695][0] , \ab[694][3] , \ab[694][2] ,
         \ab[694][1] , \ab[694][0] , \ab[693][3] , \ab[693][2] , \ab[693][1] ,
         \ab[693][0] , \ab[692][3] , \ab[692][2] , \ab[692][1] , \ab[692][0] ,
         \ab[691][3] , \ab[691][2] , \ab[691][1] , \ab[691][0] , \ab[690][3] ,
         \ab[690][2] , \ab[690][1] , \ab[690][0] , \ab[689][3] , \ab[689][2] ,
         \ab[689][1] , \ab[689][0] , \ab[688][3] , \ab[688][2] , \ab[688][1] ,
         \ab[688][0] , \ab[687][3] , \ab[687][2] , \ab[687][1] , \ab[687][0] ,
         \ab[686][3] , \ab[686][2] , \ab[686][1] , \ab[686][0] , \ab[685][3] ,
         \ab[685][2] , \ab[685][1] , \ab[685][0] , \ab[684][3] , \ab[684][2] ,
         \ab[684][1] , \ab[684][0] , \ab[683][3] , \ab[683][2] , \ab[683][1] ,
         \ab[683][0] , \ab[682][3] , \ab[682][2] , \ab[682][1] , \ab[682][0] ,
         \ab[681][3] , \ab[681][2] , \ab[681][1] , \ab[681][0] , \ab[680][3] ,
         \ab[680][2] , \ab[680][1] , \ab[680][0] , \ab[679][3] , \ab[679][2] ,
         \ab[679][1] , \ab[679][0] , \ab[678][3] , \ab[678][2] , \ab[678][1] ,
         \ab[678][0] , \ab[677][3] , \ab[677][2] , \ab[677][1] , \ab[677][0] ,
         \ab[676][3] , \ab[676][2] , \ab[676][1] , \ab[676][0] , \ab[675][3] ,
         \ab[675][2] , \ab[675][1] , \ab[675][0] , \ab[674][3] , \ab[674][2] ,
         \ab[674][1] , \ab[674][0] , \ab[673][3] , \ab[673][2] , \ab[673][1] ,
         \ab[673][0] , \ab[672][3] , \ab[672][2] , \ab[672][1] , \ab[672][0] ,
         \ab[671][3] , \ab[671][2] , \ab[671][1] , \ab[671][0] , \ab[670][3] ,
         \ab[670][2] , \ab[670][1] , \ab[670][0] , \ab[669][3] , \ab[669][2] ,
         \ab[669][1] , \ab[669][0] , \ab[668][3] , \ab[668][2] , \ab[668][1] ,
         \ab[668][0] , \ab[667][3] , \ab[667][2] , \ab[667][1] , \ab[667][0] ,
         \ab[666][3] , \ab[666][2] , \ab[666][1] , \ab[666][0] , \ab[665][3] ,
         \ab[665][2] , \ab[665][1] , \ab[665][0] , \ab[664][3] , \ab[664][2] ,
         \ab[664][1] , \ab[664][0] , \ab[663][3] , \ab[663][2] , \ab[663][1] ,
         \ab[663][0] , \ab[662][3] , \ab[662][2] , \ab[662][1] , \ab[662][0] ,
         \ab[661][3] , \ab[661][2] , \ab[661][1] , \ab[661][0] , \ab[660][3] ,
         \ab[660][2] , \ab[660][1] , \ab[660][0] , \ab[659][3] , \ab[659][2] ,
         \ab[659][1] , \ab[659][0] , \ab[658][3] , \ab[658][2] , \ab[658][1] ,
         \ab[658][0] , \ab[657][3] , \ab[657][2] , \ab[657][1] , \ab[657][0] ,
         \ab[656][3] , \ab[656][2] , \ab[656][1] , \ab[656][0] , \ab[655][3] ,
         \ab[655][2] , \ab[655][1] , \ab[655][0] , \ab[654][3] , \ab[654][2] ,
         \ab[654][1] , \ab[654][0] , \ab[653][3] , \ab[653][2] , \ab[653][1] ,
         \ab[653][0] , \ab[652][3] , \ab[652][2] , \ab[652][1] , \ab[652][0] ,
         \ab[651][3] , \ab[651][2] , \ab[651][1] , \ab[651][0] , \ab[650][3] ,
         \ab[650][2] , \ab[650][1] , \ab[650][0] , \ab[649][3] , \ab[649][2] ,
         \ab[649][1] , \ab[649][0] , \ab[648][3] , \ab[648][2] , \ab[648][1] ,
         \ab[648][0] , \ab[647][3] , \ab[647][2] , \ab[647][1] , \ab[647][0] ,
         \ab[646][3] , \ab[646][2] , \ab[646][1] , \ab[646][0] , \ab[645][3] ,
         \ab[645][2] , \ab[645][1] , \ab[645][0] , \ab[644][3] , \ab[644][2] ,
         \ab[644][1] , \ab[644][0] , \ab[643][3] , \ab[643][2] , \ab[643][1] ,
         \ab[643][0] , \ab[642][3] , \ab[642][2] , \ab[642][1] , \ab[642][0] ,
         \ab[641][3] , \ab[641][2] , \ab[641][1] , \ab[641][0] , \ab[640][3] ,
         \ab[640][2] , \ab[640][1] , \ab[640][0] , \ab[639][3] , \ab[639][2] ,
         \ab[639][1] , \ab[639][0] , \ab[638][3] , \ab[638][2] , \ab[638][1] ,
         \ab[638][0] , \ab[637][3] , \ab[637][2] , \ab[637][1] , \ab[637][0] ,
         \ab[636][3] , \ab[636][2] , \ab[636][1] , \ab[636][0] , \ab[635][3] ,
         \ab[635][2] , \ab[635][1] , \ab[635][0] , \ab[634][3] , \ab[634][2] ,
         \ab[634][1] , \ab[634][0] , \ab[633][3] , \ab[633][2] , \ab[633][1] ,
         \ab[633][0] , \ab[632][3] , \ab[632][2] , \ab[632][1] , \ab[632][0] ,
         \ab[631][3] , \ab[631][2] , \ab[631][1] , \ab[631][0] , \ab[630][3] ,
         \ab[630][2] , \ab[630][1] , \ab[630][0] , \ab[629][3] , \ab[629][2] ,
         \ab[629][1] , \ab[629][0] , \ab[628][3] , \ab[628][2] , \ab[628][1] ,
         \ab[628][0] , \ab[627][3] , \ab[627][2] , \ab[627][1] , \ab[627][0] ,
         \ab[626][3] , \ab[626][2] , \ab[626][1] , \ab[626][0] , \ab[625][3] ,
         \ab[625][2] , \ab[625][1] , \ab[625][0] , \ab[624][3] , \ab[624][2] ,
         \ab[624][1] , \ab[624][0] , \ab[623][3] , \ab[623][2] , \ab[623][1] ,
         \ab[623][0] , \ab[622][3] , \ab[622][2] , \ab[622][1] , \ab[622][0] ,
         \ab[621][3] , \ab[621][2] , \ab[621][1] , \ab[621][0] , \ab[620][3] ,
         \ab[620][2] , \ab[620][1] , \ab[620][0] , \ab[619][3] , \ab[619][2] ,
         \ab[619][1] , \ab[619][0] , \ab[618][3] , \ab[618][2] , \ab[618][1] ,
         \ab[618][0] , \ab[617][3] , \ab[617][2] , \ab[617][1] , \ab[617][0] ,
         \ab[616][3] , \ab[616][2] , \ab[616][1] , \ab[616][0] , \ab[615][3] ,
         \ab[615][2] , \ab[615][1] , \ab[615][0] , \ab[614][3] , \ab[614][2] ,
         \ab[614][1] , \ab[614][0] , \ab[613][3] , \ab[613][2] , \ab[613][1] ,
         \ab[613][0] , \ab[612][3] , \ab[612][2] , \ab[612][1] , \ab[612][0] ,
         \ab[611][3] , \ab[611][2] , \ab[611][1] , \ab[611][0] , \ab[610][3] ,
         \ab[610][2] , \ab[610][1] , \ab[610][0] , \ab[609][3] , \ab[609][2] ,
         \ab[609][1] , \ab[609][0] , \ab[608][3] , \ab[608][2] , \ab[608][1] ,
         \ab[608][0] , \ab[607][3] , \ab[607][2] , \ab[607][1] , \ab[607][0] ,
         \ab[606][3] , \ab[606][2] , \ab[606][1] , \ab[606][0] , \ab[605][3] ,
         \ab[605][2] , \ab[605][1] , \ab[605][0] , \ab[604][3] , \ab[604][2] ,
         \ab[604][1] , \ab[604][0] , \ab[603][3] , \ab[603][2] , \ab[603][1] ,
         \ab[603][0] , \ab[602][3] , \ab[602][2] , \ab[602][1] , \ab[602][0] ,
         \ab[601][3] , \ab[601][2] , \ab[601][1] , \ab[601][0] , \ab[600][3] ,
         \ab[600][2] , \ab[600][1] , \ab[600][0] , \ab[599][3] , \ab[599][2] ,
         \ab[599][1] , \ab[599][0] , \ab[598][3] , \ab[598][2] , \ab[598][1] ,
         \ab[598][0] , \ab[597][3] , \ab[597][2] , \ab[597][1] , \ab[597][0] ,
         \ab[596][3] , \ab[596][2] , \ab[596][1] , \ab[596][0] , \ab[595][3] ,
         \ab[595][2] , \ab[595][1] , \ab[595][0] , \ab[594][3] , \ab[594][2] ,
         \ab[594][1] , \ab[594][0] , \ab[593][3] , \ab[593][2] , \ab[593][1] ,
         \ab[593][0] , \ab[592][3] , \ab[592][2] , \ab[592][1] , \ab[592][0] ,
         \ab[591][3] , \ab[591][2] , \ab[591][1] , \ab[591][0] , \ab[590][3] ,
         \ab[590][2] , \ab[590][1] , \ab[590][0] , \ab[589][3] , \ab[589][2] ,
         \ab[589][1] , \ab[589][0] , \ab[588][3] , \ab[588][2] , \ab[588][1] ,
         \ab[588][0] , \ab[587][3] , \ab[587][2] , \ab[587][1] , \ab[587][0] ,
         \ab[586][3] , \ab[586][2] , \ab[586][1] , \ab[586][0] , \ab[585][3] ,
         \ab[585][2] , \ab[585][1] , \ab[585][0] , \ab[584][3] , \ab[584][2] ,
         \ab[584][1] , \ab[584][0] , \ab[583][3] , \ab[583][2] , \ab[583][1] ,
         \ab[583][0] , \ab[582][3] , \ab[582][2] , \ab[582][1] , \ab[582][0] ,
         \ab[581][3] , \ab[581][2] , \ab[581][1] , \ab[581][0] , \ab[580][3] ,
         \ab[580][2] , \ab[580][1] , \ab[580][0] , \ab[579][3] , \ab[579][2] ,
         \ab[579][1] , \ab[579][0] , \ab[578][3] , \ab[578][2] , \ab[578][1] ,
         \ab[578][0] , \ab[577][3] , \ab[577][2] , \ab[577][1] , \ab[577][0] ,
         \ab[576][3] , \ab[576][2] , \ab[576][1] , \ab[576][0] , \ab[575][3] ,
         \ab[575][2] , \ab[575][1] , \ab[575][0] , \ab[574][3] , \ab[574][2] ,
         \ab[574][1] , \ab[574][0] , \ab[573][3] , \ab[573][2] , \ab[573][1] ,
         \ab[573][0] , \ab[572][3] , \ab[572][2] , \ab[572][1] , \ab[572][0] ,
         \ab[571][3] , \ab[571][2] , \ab[571][1] , \ab[571][0] , \ab[570][3] ,
         \ab[570][2] , \ab[570][1] , \ab[570][0] , \ab[569][3] , \ab[569][2] ,
         \ab[569][1] , \ab[569][0] , \ab[568][3] , \ab[568][2] , \ab[568][1] ,
         \ab[568][0] , \ab[567][3] , \ab[567][2] , \ab[567][1] , \ab[567][0] ,
         \ab[566][3] , \ab[566][2] , \ab[566][1] , \ab[566][0] , \ab[565][3] ,
         \ab[565][2] , \ab[565][1] , \ab[565][0] , \ab[564][3] , \ab[564][2] ,
         \ab[564][1] , \ab[564][0] , \ab[563][3] , \ab[563][2] , \ab[563][1] ,
         \ab[563][0] , \ab[562][3] , \ab[562][2] , \ab[562][1] , \ab[562][0] ,
         \ab[561][3] , \ab[561][2] , \ab[561][1] , \ab[561][0] , \ab[560][3] ,
         \ab[560][2] , \ab[560][1] , \ab[560][0] , \ab[559][3] , \ab[559][2] ,
         \ab[559][1] , \ab[559][0] , \ab[558][3] , \ab[558][2] , \ab[558][1] ,
         \ab[558][0] , \ab[557][3] , \ab[557][2] , \ab[557][1] , \ab[557][0] ,
         \ab[556][3] , \ab[556][2] , \ab[556][1] , \ab[556][0] , \ab[555][3] ,
         \ab[555][2] , \ab[555][1] , \ab[555][0] , \ab[554][3] , \ab[554][2] ,
         \ab[554][1] , \ab[554][0] , \ab[553][3] , \ab[553][2] , \ab[553][1] ,
         \ab[553][0] , \ab[552][3] , \ab[552][2] , \ab[552][1] , \ab[552][0] ,
         \ab[551][3] , \ab[551][2] , \ab[551][1] , \ab[551][0] , \ab[550][3] ,
         \ab[550][2] , \ab[550][1] , \ab[550][0] , \ab[549][3] , \ab[549][2] ,
         \ab[549][1] , \ab[549][0] , \ab[548][3] , \ab[548][2] , \ab[548][1] ,
         \ab[548][0] , \ab[547][3] , \ab[547][2] , \ab[547][1] , \ab[547][0] ,
         \ab[546][3] , \ab[546][2] , \ab[546][1] , \ab[546][0] , \ab[545][3] ,
         \ab[545][2] , \ab[545][1] , \ab[545][0] , \ab[544][3] , \ab[544][2] ,
         \ab[544][1] , \ab[544][0] , \ab[543][3] , \ab[543][2] , \ab[543][1] ,
         \ab[543][0] , \ab[542][3] , \ab[542][2] , \ab[542][1] , \ab[542][0] ,
         \ab[541][3] , \ab[541][2] , \ab[541][1] , \ab[541][0] , \ab[540][3] ,
         \ab[540][2] , \ab[540][1] , \ab[540][0] , \ab[539][3] , \ab[539][2] ,
         \ab[539][1] , \ab[539][0] , \ab[538][3] , \ab[538][2] , \ab[538][1] ,
         \ab[538][0] , \ab[537][3] , \ab[537][2] , \ab[537][1] , \ab[537][0] ,
         \ab[536][3] , \ab[536][2] , \ab[536][1] , \ab[536][0] , \ab[535][3] ,
         \ab[535][2] , \ab[535][1] , \ab[535][0] , \ab[534][3] , \ab[534][2] ,
         \ab[534][1] , \ab[534][0] , \ab[533][3] , \ab[533][2] , \ab[533][1] ,
         \ab[533][0] , \ab[532][3] , \ab[532][2] , \ab[532][1] , \ab[532][0] ,
         \ab[531][3] , \ab[531][2] , \ab[531][1] , \ab[531][0] , \ab[530][3] ,
         \ab[530][2] , \ab[530][1] , \ab[530][0] , \ab[529][3] , \ab[529][2] ,
         \ab[529][1] , \ab[529][0] , \ab[528][3] , \ab[528][2] , \ab[528][1] ,
         \ab[528][0] , \ab[527][3] , \ab[527][2] , \ab[527][1] , \ab[527][0] ,
         \ab[526][3] , \ab[526][2] , \ab[526][1] , \ab[526][0] , \ab[525][3] ,
         \ab[525][2] , \ab[525][1] , \ab[525][0] , \ab[524][3] , \ab[524][2] ,
         \ab[524][1] , \ab[524][0] , \ab[523][3] , \ab[523][2] , \ab[523][1] ,
         \ab[523][0] , \ab[522][3] , \ab[522][2] , \ab[522][1] , \ab[522][0] ,
         \ab[521][3] , \ab[521][2] , \ab[521][1] , \ab[521][0] , \ab[520][3] ,
         \ab[520][2] , \ab[520][1] , \ab[520][0] , \ab[519][3] , \ab[519][2] ,
         \ab[519][1] , \ab[519][0] , \ab[518][3] , \ab[518][2] , \ab[518][1] ,
         \ab[518][0] , \ab[517][3] , \ab[517][2] , \ab[517][1] , \ab[517][0] ,
         \ab[516][3] , \ab[516][2] , \ab[516][1] , \ab[516][0] , \ab[515][3] ,
         \ab[515][2] , \ab[515][1] , \ab[515][0] , \ab[514][3] , \ab[514][2] ,
         \ab[514][1] , \ab[514][0] , \ab[513][3] , \ab[513][2] , \ab[513][1] ,
         \ab[513][0] , \ab[512][3] , \ab[512][2] , \ab[512][1] , \ab[512][0] ,
         \ab[511][3] , \ab[511][2] , \ab[511][1] , \ab[511][0] , \ab[510][3] ,
         \ab[510][2] , \ab[510][1] , \ab[510][0] , \ab[509][3] , \ab[509][2] ,
         \ab[509][1] , \ab[509][0] , \ab[508][3] , \ab[508][2] , \ab[508][1] ,
         \ab[508][0] , \ab[507][3] , \ab[507][2] , \ab[507][1] , \ab[507][0] ,
         \ab[506][3] , \ab[506][2] , \ab[506][1] , \ab[506][0] , \ab[505][3] ,
         \ab[505][2] , \ab[505][1] , \ab[505][0] , \ab[504][3] , \ab[504][2] ,
         \ab[504][1] , \ab[504][0] , \ab[503][3] , \ab[503][2] , \ab[503][1] ,
         \ab[503][0] , \ab[502][3] , \ab[502][2] , \ab[502][1] , \ab[502][0] ,
         \ab[501][3] , \ab[501][2] , \ab[501][1] , \ab[501][0] , \ab[500][3] ,
         \ab[500][2] , \ab[500][1] , \ab[500][0] , \ab[499][3] , \ab[499][2] ,
         \ab[499][1] , \ab[499][0] , \ab[498][3] , \ab[498][2] , \ab[498][1] ,
         \ab[498][0] , \ab[497][3] , \ab[497][2] , \ab[497][1] , \ab[497][0] ,
         \ab[496][3] , \ab[496][2] , \ab[496][1] , \ab[496][0] , \ab[495][3] ,
         \ab[495][2] , \ab[495][1] , \ab[495][0] , \ab[494][3] , \ab[494][2] ,
         \ab[494][1] , \ab[494][0] , \ab[493][3] , \ab[493][2] , \ab[493][1] ,
         \ab[493][0] , \ab[492][3] , \ab[492][2] , \ab[492][1] , \ab[492][0] ,
         \ab[491][3] , \ab[491][2] , \ab[491][1] , \ab[491][0] , \ab[490][3] ,
         \ab[490][2] , \ab[490][1] , \ab[490][0] , \ab[489][3] , \ab[489][2] ,
         \ab[489][1] , \ab[489][0] , \ab[488][3] , \ab[488][2] , \ab[488][1] ,
         \ab[488][0] , \ab[487][3] , \ab[487][2] , \ab[487][1] , \ab[487][0] ,
         \ab[486][3] , \ab[486][2] , \ab[486][1] , \ab[486][0] , \ab[485][3] ,
         \ab[485][2] , \ab[485][1] , \ab[485][0] , \ab[484][3] , \ab[484][2] ,
         \ab[484][1] , \ab[484][0] , \ab[483][3] , \ab[483][2] , \ab[483][1] ,
         \ab[483][0] , \ab[482][3] , \ab[482][2] , \ab[482][1] , \ab[482][0] ,
         \ab[481][3] , \ab[481][2] , \ab[481][1] , \ab[481][0] , \ab[480][3] ,
         \ab[480][2] , \ab[480][1] , \ab[480][0] , \ab[479][3] , \ab[479][2] ,
         \ab[479][1] , \ab[479][0] , \ab[478][3] , \ab[478][2] , \ab[478][1] ,
         \ab[478][0] , \ab[477][3] , \ab[477][2] , \ab[477][1] , \ab[477][0] ,
         \ab[476][3] , \ab[476][2] , \ab[476][1] , \ab[476][0] , \ab[475][3] ,
         \ab[475][2] , \ab[475][1] , \ab[475][0] , \ab[474][3] , \ab[474][2] ,
         \ab[474][1] , \ab[474][0] , \ab[473][3] , \ab[473][2] , \ab[473][1] ,
         \ab[473][0] , \ab[472][3] , \ab[472][2] , \ab[472][1] , \ab[472][0] ,
         \ab[471][3] , \ab[471][2] , \ab[471][1] , \ab[471][0] , \ab[470][3] ,
         \ab[470][2] , \ab[470][1] , \ab[470][0] , \ab[469][3] , \ab[469][2] ,
         \ab[469][1] , \ab[469][0] , \ab[468][3] , \ab[468][2] , \ab[468][1] ,
         \ab[468][0] , \ab[467][3] , \ab[467][2] , \ab[467][1] , \ab[467][0] ,
         \ab[466][3] , \ab[466][2] , \ab[466][1] , \ab[466][0] , \ab[465][3] ,
         \ab[465][2] , \ab[465][1] , \ab[465][0] , \ab[464][3] , \ab[464][2] ,
         \ab[464][1] , \ab[464][0] , \ab[463][3] , \ab[463][2] , \ab[463][1] ,
         \ab[463][0] , \ab[462][3] , \ab[462][2] , \ab[462][1] , \ab[462][0] ,
         \ab[461][3] , \ab[461][2] , \ab[461][1] , \ab[461][0] , \ab[460][3] ,
         \ab[460][2] , \ab[460][1] , \ab[460][0] , \ab[459][3] , \ab[459][2] ,
         \ab[459][1] , \ab[459][0] , \ab[458][3] , \ab[458][2] , \ab[458][1] ,
         \ab[458][0] , \ab[457][3] , \ab[457][2] , \ab[457][1] , \ab[457][0] ,
         \ab[456][3] , \ab[456][2] , \ab[456][1] , \ab[456][0] , \ab[455][3] ,
         \ab[455][2] , \ab[455][1] , \ab[455][0] , \ab[454][3] , \ab[454][2] ,
         \ab[454][1] , \ab[454][0] , \ab[453][3] , \ab[453][2] , \ab[453][1] ,
         \ab[453][0] , \ab[452][3] , \ab[452][2] , \ab[452][1] , \ab[452][0] ,
         \ab[451][3] , \ab[451][2] , \ab[451][1] , \ab[451][0] , \ab[450][3] ,
         \ab[450][2] , \ab[450][1] , \ab[450][0] , \ab[449][3] , \ab[449][2] ,
         \ab[449][1] , \ab[449][0] , \ab[448][3] , \ab[448][2] , \ab[448][1] ,
         \ab[448][0] , \ab[447][3] , \ab[447][2] , \ab[447][1] , \ab[447][0] ,
         \ab[446][3] , \ab[446][2] , \ab[446][1] , \ab[446][0] , \ab[445][3] ,
         \ab[445][2] , \ab[445][1] , \ab[445][0] , \ab[444][3] , \ab[444][2] ,
         \ab[444][1] , \ab[444][0] , \ab[443][3] , \ab[443][2] , \ab[443][1] ,
         \ab[443][0] , \ab[442][3] , \ab[442][2] , \ab[442][1] , \ab[442][0] ,
         \ab[441][3] , \ab[441][2] , \ab[441][1] , \ab[441][0] , \ab[440][3] ,
         \ab[440][2] , \ab[440][1] , \ab[440][0] , \ab[439][3] , \ab[439][2] ,
         \ab[439][1] , \ab[439][0] , \ab[438][3] , \ab[438][2] , \ab[438][1] ,
         \ab[438][0] , \ab[437][3] , \ab[437][2] , \ab[437][1] , \ab[437][0] ,
         \ab[436][3] , \ab[436][2] , \ab[436][1] , \ab[436][0] , \ab[435][3] ,
         \ab[435][2] , \ab[435][1] , \ab[435][0] , \ab[434][3] , \ab[434][2] ,
         \ab[434][1] , \ab[434][0] , \ab[433][3] , \ab[433][2] , \ab[433][1] ,
         \ab[433][0] , \ab[432][3] , \ab[432][2] , \ab[432][1] , \ab[432][0] ,
         \ab[431][3] , \ab[431][2] , \ab[431][1] , \ab[431][0] , \ab[430][3] ,
         \ab[430][2] , \ab[430][1] , \ab[430][0] , \ab[429][3] , \ab[429][2] ,
         \ab[429][1] , \ab[429][0] , \ab[428][3] , \ab[428][2] , \ab[428][1] ,
         \ab[428][0] , \ab[427][3] , \ab[427][2] , \ab[427][1] , \ab[427][0] ,
         \ab[426][3] , \ab[426][2] , \ab[426][1] , \ab[426][0] , \ab[425][3] ,
         \ab[425][2] , \ab[425][1] , \ab[425][0] , \ab[424][3] , \ab[424][2] ,
         \ab[424][1] , \ab[424][0] , \ab[423][3] , \ab[423][2] , \ab[423][1] ,
         \ab[423][0] , \ab[422][3] , \ab[422][2] , \ab[422][1] , \ab[422][0] ,
         \ab[421][3] , \ab[421][2] , \ab[421][1] , \ab[421][0] , \ab[420][3] ,
         \ab[420][2] , \ab[420][1] , \ab[420][0] , \ab[419][3] , \ab[419][2] ,
         \ab[419][1] , \ab[419][0] , \ab[418][3] , \ab[418][2] , \ab[418][1] ,
         \ab[418][0] , \ab[417][3] , \ab[417][2] , \ab[417][1] , \ab[417][0] ,
         \ab[416][3] , \ab[416][2] , \ab[416][1] , \ab[416][0] , \ab[415][3] ,
         \ab[415][2] , \ab[415][1] , \ab[415][0] , \ab[414][3] , \ab[414][2] ,
         \ab[414][1] , \ab[414][0] , \ab[413][3] , \ab[413][2] , \ab[413][1] ,
         \ab[413][0] , \ab[412][3] , \ab[412][2] , \ab[412][1] , \ab[412][0] ,
         \ab[411][3] , \ab[411][2] , \ab[411][1] , \ab[411][0] , \ab[410][3] ,
         \ab[410][2] , \ab[410][1] , \ab[410][0] , \ab[409][3] , \ab[409][2] ,
         \ab[409][1] , \ab[409][0] , \ab[408][3] , \ab[408][2] , \ab[408][1] ,
         \ab[408][0] , \ab[407][3] , \ab[407][2] , \ab[407][1] , \ab[407][0] ,
         \ab[406][3] , \ab[406][2] , \ab[406][1] , \ab[406][0] , \ab[405][3] ,
         \ab[405][2] , \ab[405][1] , \ab[405][0] , \ab[404][3] , \ab[404][2] ,
         \ab[404][1] , \ab[404][0] , \ab[403][3] , \ab[403][2] , \ab[403][1] ,
         \ab[403][0] , \ab[402][3] , \ab[402][2] , \ab[402][1] , \ab[402][0] ,
         \ab[401][3] , \ab[401][2] , \ab[401][1] , \ab[401][0] , \ab[400][3] ,
         \ab[400][2] , \ab[400][1] , \ab[400][0] , \ab[399][3] , \ab[399][2] ,
         \ab[399][1] , \ab[399][0] , \ab[398][3] , \ab[398][2] , \ab[398][1] ,
         \ab[398][0] , \ab[397][3] , \ab[397][2] , \ab[397][1] , \ab[397][0] ,
         \ab[396][3] , \ab[396][2] , \ab[396][1] , \ab[396][0] , \ab[395][3] ,
         \ab[395][2] , \ab[395][1] , \ab[395][0] , \ab[394][3] , \ab[394][2] ,
         \ab[394][1] , \ab[394][0] , \ab[393][3] , \ab[393][2] , \ab[393][1] ,
         \ab[393][0] , \ab[392][3] , \ab[392][2] , \ab[392][1] , \ab[392][0] ,
         \ab[391][3] , \ab[391][2] , \ab[391][1] , \ab[391][0] , \ab[390][3] ,
         \ab[390][2] , \ab[390][1] , \ab[390][0] , \ab[389][3] , \ab[389][2] ,
         \ab[389][1] , \ab[389][0] , \ab[388][3] , \ab[388][2] , \ab[388][1] ,
         \ab[388][0] , \ab[387][3] , \ab[387][2] , \ab[387][1] , \ab[387][0] ,
         \ab[386][3] , \ab[386][2] , \ab[386][1] , \ab[386][0] , \ab[385][3] ,
         \ab[385][2] , \ab[385][1] , \ab[385][0] , \ab[384][3] , \ab[384][2] ,
         \ab[384][1] , \ab[384][0] , \ab[383][3] , \ab[383][2] , \ab[383][1] ,
         \ab[383][0] , \ab[382][3] , \ab[382][2] , \ab[382][1] , \ab[382][0] ,
         \ab[381][3] , \ab[381][2] , \ab[381][1] , \ab[381][0] , \ab[380][3] ,
         \ab[380][2] , \ab[380][1] , \ab[380][0] , \ab[379][3] , \ab[379][2] ,
         \ab[379][1] , \ab[379][0] , \ab[378][3] , \ab[378][2] , \ab[378][1] ,
         \ab[378][0] , \ab[377][3] , \ab[377][2] , \ab[377][1] , \ab[377][0] ,
         \ab[376][3] , \ab[376][2] , \ab[376][1] , \ab[376][0] , \ab[375][3] ,
         \ab[375][2] , \ab[375][1] , \ab[375][0] , \ab[374][3] , \ab[374][2] ,
         \ab[374][1] , \ab[374][0] , \ab[373][3] , \ab[373][2] , \ab[373][1] ,
         \ab[373][0] , \ab[372][3] , \ab[372][2] , \ab[372][1] , \ab[372][0] ,
         \ab[371][3] , \ab[371][2] , \ab[371][1] , \ab[371][0] , \ab[370][3] ,
         \ab[370][2] , \ab[370][1] , \ab[370][0] , \ab[369][3] , \ab[369][2] ,
         \ab[369][1] , \ab[369][0] , \ab[368][3] , \ab[368][2] , \ab[368][1] ,
         \ab[368][0] , \ab[367][3] , \ab[367][2] , \ab[367][1] , \ab[367][0] ,
         \ab[366][3] , \ab[366][2] , \ab[366][1] , \ab[366][0] , \ab[365][3] ,
         \ab[365][2] , \ab[365][1] , \ab[365][0] , \ab[364][3] , \ab[364][2] ,
         \ab[364][1] , \ab[364][0] , \ab[363][3] , \ab[363][2] , \ab[363][1] ,
         \ab[363][0] , \ab[362][3] , \ab[362][2] , \ab[362][1] , \ab[362][0] ,
         \ab[361][3] , \ab[361][2] , \ab[361][1] , \ab[361][0] , \ab[360][3] ,
         \ab[360][2] , \ab[360][1] , \ab[360][0] , \ab[359][3] , \ab[359][2] ,
         \ab[359][1] , \ab[359][0] , \ab[358][3] , \ab[358][2] , \ab[358][1] ,
         \ab[358][0] , \ab[357][3] , \ab[357][2] , \ab[357][1] , \ab[357][0] ,
         \ab[356][3] , \ab[356][2] , \ab[356][1] , \ab[356][0] , \ab[355][3] ,
         \ab[355][2] , \ab[355][1] , \ab[355][0] , \ab[354][3] , \ab[354][2] ,
         \ab[354][1] , \ab[354][0] , \ab[353][3] , \ab[353][2] , \ab[353][1] ,
         \ab[353][0] , \ab[352][3] , \ab[352][2] , \ab[352][1] , \ab[352][0] ,
         \ab[351][3] , \ab[351][2] , \ab[351][1] , \ab[351][0] , \ab[350][3] ,
         \ab[350][2] , \ab[350][1] , \ab[350][0] , \ab[349][3] , \ab[349][2] ,
         \ab[349][1] , \ab[349][0] , \ab[348][3] , \ab[348][2] , \ab[348][1] ,
         \ab[348][0] , \ab[347][3] , \ab[347][2] , \ab[347][1] , \ab[347][0] ,
         \ab[346][3] , \ab[346][2] , \ab[346][1] , \ab[346][0] , \ab[345][3] ,
         \ab[345][2] , \ab[345][1] , \ab[345][0] , \ab[344][3] , \ab[344][2] ,
         \ab[344][1] , \ab[344][0] , \ab[343][3] , \ab[343][2] , \ab[343][1] ,
         \ab[343][0] , \ab[342][3] , \ab[342][2] , \ab[342][1] , \ab[342][0] ,
         \ab[341][3] , \ab[341][2] , \ab[341][1] , \ab[341][0] , \ab[340][3] ,
         \ab[340][2] , \ab[340][1] , \ab[340][0] , \ab[339][3] , \ab[339][2] ,
         \ab[339][1] , \ab[339][0] , \ab[338][3] , \ab[338][2] , \ab[338][1] ,
         \ab[338][0] , \ab[337][3] , \ab[337][2] , \ab[337][1] , \ab[337][0] ,
         \ab[336][3] , \ab[336][2] , \ab[336][1] , \ab[336][0] , \ab[335][3] ,
         \ab[335][2] , \ab[335][1] , \ab[335][0] , \ab[334][3] , \ab[334][2] ,
         \ab[334][1] , \ab[334][0] , \ab[333][3] , \ab[333][2] , \ab[333][1] ,
         \ab[333][0] , \ab[332][3] , \ab[332][2] , \ab[332][1] , \ab[332][0] ,
         \ab[331][3] , \ab[331][2] , \ab[331][1] , \ab[331][0] , \ab[330][3] ,
         \ab[330][2] , \ab[330][1] , \ab[330][0] , \ab[329][3] , \ab[329][2] ,
         \ab[329][1] , \ab[329][0] , \ab[328][3] , \ab[328][2] , \ab[328][1] ,
         \ab[328][0] , \ab[327][3] , \ab[327][2] , \ab[327][1] , \ab[327][0] ,
         \ab[326][3] , \ab[326][2] , \ab[326][1] , \ab[326][0] , \ab[325][3] ,
         \ab[325][2] , \ab[325][1] , \ab[325][0] , \ab[324][3] , \ab[324][2] ,
         \ab[324][1] , \ab[324][0] , \ab[323][3] , \ab[323][2] , \ab[323][1] ,
         \ab[323][0] , \ab[322][3] , \ab[322][2] , \ab[322][1] , \ab[322][0] ,
         \ab[321][3] , \ab[321][2] , \ab[321][1] , \ab[321][0] , \ab[320][3] ,
         \ab[320][2] , \ab[320][1] , \ab[320][0] , \ab[319][3] , \ab[319][2] ,
         \ab[319][1] , \ab[319][0] , \ab[318][3] , \ab[318][2] , \ab[318][1] ,
         \ab[318][0] , \ab[317][3] , \ab[317][2] , \ab[317][1] , \ab[317][0] ,
         \ab[316][3] , \ab[316][2] , \ab[316][1] , \ab[316][0] , \ab[315][3] ,
         \ab[315][2] , \ab[315][1] , \ab[315][0] , \ab[314][3] , \ab[314][2] ,
         \ab[314][1] , \ab[314][0] , \ab[313][3] , \ab[313][2] , \ab[313][1] ,
         \ab[313][0] , \ab[312][3] , \ab[312][2] , \ab[312][1] , \ab[312][0] ,
         \ab[311][3] , \ab[311][2] , \ab[311][1] , \ab[311][0] , \ab[310][3] ,
         \ab[310][2] , \ab[310][1] , \ab[310][0] , \ab[309][3] , \ab[309][2] ,
         \ab[309][1] , \ab[309][0] , \ab[308][3] , \ab[308][2] , \ab[308][1] ,
         \ab[308][0] , \ab[307][3] , \ab[307][2] , \ab[307][1] , \ab[307][0] ,
         \ab[306][3] , \ab[306][2] , \ab[306][1] , \ab[306][0] , \ab[305][3] ,
         \ab[305][2] , \ab[305][1] , \ab[305][0] , \ab[304][3] , \ab[304][2] ,
         \ab[304][1] , \ab[304][0] , \ab[303][3] , \ab[303][2] , \ab[303][1] ,
         \ab[303][0] , \ab[302][3] , \ab[302][2] , \ab[302][1] , \ab[302][0] ,
         \ab[301][3] , \ab[301][2] , \ab[301][1] , \ab[301][0] , \ab[300][3] ,
         \ab[300][2] , \ab[300][1] , \ab[300][0] , \ab[299][3] , \ab[299][2] ,
         \ab[299][1] , \ab[299][0] , \ab[298][3] , \ab[298][2] , \ab[298][1] ,
         \ab[298][0] , \ab[297][3] , \ab[297][2] , \ab[297][1] , \ab[297][0] ,
         \ab[296][3] , \ab[296][2] , \ab[296][1] , \ab[296][0] , \ab[295][3] ,
         \ab[295][2] , \ab[295][1] , \ab[295][0] , \ab[294][3] , \ab[294][2] ,
         \ab[294][1] , \ab[294][0] , \ab[293][3] , \ab[293][2] , \ab[293][1] ,
         \ab[293][0] , \ab[292][3] , \ab[292][2] , \ab[292][1] , \ab[292][0] ,
         \ab[291][3] , \ab[291][2] , \ab[291][1] , \ab[291][0] , \ab[290][3] ,
         \ab[290][2] , \ab[290][1] , \ab[290][0] , \ab[289][3] , \ab[289][2] ,
         \ab[289][1] , \ab[289][0] , \ab[288][3] , \ab[288][2] , \ab[288][1] ,
         \ab[288][0] , \ab[287][3] , \ab[287][2] , \ab[287][1] , \ab[287][0] ,
         \ab[286][3] , \ab[286][2] , \ab[286][1] , \ab[286][0] , \ab[285][3] ,
         \ab[285][2] , \ab[285][1] , \ab[285][0] , \ab[284][3] , \ab[284][2] ,
         \ab[284][1] , \ab[284][0] , \ab[283][3] , \ab[283][2] , \ab[283][1] ,
         \ab[283][0] , \ab[282][3] , \ab[282][2] , \ab[282][1] , \ab[282][0] ,
         \ab[281][3] , \ab[281][2] , \ab[281][1] , \ab[281][0] , \ab[280][3] ,
         \ab[280][2] , \ab[280][1] , \ab[280][0] , \ab[279][3] , \ab[279][2] ,
         \ab[279][1] , \ab[279][0] , \ab[278][3] , \ab[278][2] , \ab[278][1] ,
         \ab[278][0] , \ab[277][3] , \ab[277][2] , \ab[277][1] , \ab[277][0] ,
         \ab[276][3] , \ab[276][2] , \ab[276][1] , \ab[276][0] , \ab[275][3] ,
         \ab[275][2] , \ab[275][1] , \ab[275][0] , \ab[274][3] , \ab[274][2] ,
         \ab[274][1] , \ab[274][0] , \ab[273][3] , \ab[273][2] , \ab[273][1] ,
         \ab[273][0] , \ab[272][3] , \ab[272][2] , \ab[272][1] , \ab[272][0] ,
         \ab[271][3] , \ab[271][2] , \ab[271][1] , \ab[271][0] , \ab[270][3] ,
         \ab[270][2] , \ab[270][1] , \ab[270][0] , \ab[269][3] , \ab[269][2] ,
         \ab[269][1] , \ab[269][0] , \ab[268][3] , \ab[268][2] , \ab[268][1] ,
         \ab[268][0] , \ab[267][3] , \ab[267][2] , \ab[267][1] , \ab[267][0] ,
         \ab[266][3] , \ab[266][2] , \ab[266][1] , \ab[266][0] , \ab[265][3] ,
         \ab[265][2] , \ab[265][1] , \ab[265][0] , \ab[264][3] , \ab[264][2] ,
         \ab[264][1] , \ab[264][0] , \ab[263][3] , \ab[263][2] , \ab[263][1] ,
         \ab[263][0] , \ab[262][3] , \ab[262][2] , \ab[262][1] , \ab[262][0] ,
         \ab[261][3] , \ab[261][2] , \ab[261][1] , \ab[261][0] , \ab[260][3] ,
         \ab[260][2] , \ab[260][1] , \ab[260][0] , \ab[259][3] , \ab[259][2] ,
         \ab[259][1] , \ab[259][0] , \ab[258][3] , \ab[258][2] , \ab[258][1] ,
         \ab[258][0] , \ab[257][3] , \ab[257][2] , \ab[257][1] , \ab[257][0] ,
         \ab[256][3] , \ab[256][2] , \ab[256][1] , \ab[256][0] , \ab[255][3] ,
         \ab[255][2] , \ab[255][1] , \ab[255][0] , \ab[254][3] , \ab[254][2] ,
         \ab[254][1] , \ab[254][0] , \ab[253][3] , \ab[253][2] , \ab[253][1] ,
         \ab[253][0] , \ab[252][3] , \ab[252][2] , \ab[252][1] , \ab[252][0] ,
         \ab[251][3] , \ab[251][2] , \ab[251][1] , \ab[251][0] , \ab[250][3] ,
         \ab[250][2] , \ab[250][1] , \ab[250][0] , \ab[249][3] , \ab[249][2] ,
         \ab[249][1] , \ab[249][0] , \ab[248][3] , \ab[248][2] , \ab[248][1] ,
         \ab[248][0] , \ab[247][3] , \ab[247][2] , \ab[247][1] , \ab[247][0] ,
         \ab[246][3] , \ab[246][2] , \ab[246][1] , \ab[246][0] , \ab[245][3] ,
         \ab[245][2] , \ab[245][1] , \ab[245][0] , \ab[244][3] , \ab[244][2] ,
         \ab[244][1] , \ab[244][0] , \ab[243][3] , \ab[243][2] , \ab[243][1] ,
         \ab[243][0] , \ab[242][3] , \ab[242][2] , \ab[242][1] , \ab[242][0] ,
         \ab[241][3] , \ab[241][2] , \ab[241][1] , \ab[241][0] , \ab[240][3] ,
         \ab[240][2] , \ab[240][1] , \ab[240][0] , \ab[239][3] , \ab[239][2] ,
         \ab[239][1] , \ab[239][0] , \ab[238][3] , \ab[238][2] , \ab[238][1] ,
         \ab[238][0] , \ab[237][3] , \ab[237][2] , \ab[237][1] , \ab[237][0] ,
         \ab[236][3] , \ab[236][2] , \ab[236][1] , \ab[236][0] , \ab[235][3] ,
         \ab[235][2] , \ab[235][1] , \ab[235][0] , \ab[234][3] , \ab[234][2] ,
         \ab[234][1] , \ab[234][0] , \ab[233][3] , \ab[233][2] , \ab[233][1] ,
         \ab[233][0] , \ab[232][3] , \ab[232][2] , \ab[232][1] , \ab[232][0] ,
         \ab[231][3] , \ab[231][2] , \ab[231][1] , \ab[231][0] , \ab[230][3] ,
         \ab[230][2] , \ab[230][1] , \ab[230][0] , \ab[229][3] , \ab[229][2] ,
         \ab[229][1] , \ab[229][0] , \ab[228][3] , \ab[228][2] , \ab[228][1] ,
         \ab[228][0] , \ab[227][3] , \ab[227][2] , \ab[227][1] , \ab[227][0] ,
         \ab[226][3] , \ab[226][2] , \ab[226][1] , \ab[226][0] , \ab[225][3] ,
         \ab[225][2] , \ab[225][1] , \ab[225][0] , \ab[224][3] , \ab[224][2] ,
         \ab[224][1] , \ab[224][0] , \ab[223][3] , \ab[223][2] , \ab[223][1] ,
         \ab[223][0] , \ab[222][3] , \ab[222][2] , \ab[222][1] , \ab[222][0] ,
         \ab[221][3] , \ab[221][2] , \ab[221][1] , \ab[221][0] , \ab[220][3] ,
         \ab[220][2] , \ab[220][1] , \ab[220][0] , \ab[219][3] , \ab[219][2] ,
         \ab[219][1] , \ab[219][0] , \ab[218][3] , \ab[218][2] , \ab[218][1] ,
         \ab[218][0] , \ab[217][3] , \ab[217][2] , \ab[217][1] , \ab[217][0] ,
         \ab[216][3] , \ab[216][2] , \ab[216][1] , \ab[216][0] , \ab[215][3] ,
         \ab[215][2] , \ab[215][1] , \ab[215][0] , \ab[214][3] , \ab[214][2] ,
         \ab[214][1] , \ab[214][0] , \ab[213][3] , \ab[213][2] , \ab[213][1] ,
         \ab[213][0] , \ab[212][3] , \ab[212][2] , \ab[212][1] , \ab[212][0] ,
         \ab[211][3] , \ab[211][2] , \ab[211][1] , \ab[211][0] , \ab[210][3] ,
         \ab[210][2] , \ab[210][1] , \ab[210][0] , \ab[209][3] , \ab[209][2] ,
         \ab[209][1] , \ab[209][0] , \ab[208][3] , \ab[208][2] , \ab[208][1] ,
         \ab[208][0] , \ab[207][3] , \ab[207][2] , \ab[207][1] , \ab[207][0] ,
         \ab[206][3] , \ab[206][2] , \ab[206][1] , \ab[206][0] , \ab[205][3] ,
         \ab[205][2] , \ab[205][1] , \ab[205][0] , \ab[204][3] , \ab[204][2] ,
         \ab[204][1] , \ab[204][0] , \ab[203][3] , \ab[203][2] , \ab[203][1] ,
         \ab[203][0] , \ab[202][3] , \ab[202][2] , \ab[202][1] , \ab[202][0] ,
         \ab[201][3] , \ab[201][2] , \ab[201][1] , \ab[201][0] , \ab[200][3] ,
         \ab[200][2] , \ab[200][1] , \ab[200][0] , \ab[199][3] , \ab[199][2] ,
         \ab[199][1] , \ab[199][0] , \ab[198][3] , \ab[198][2] , \ab[198][1] ,
         \ab[198][0] , \ab[197][3] , \ab[197][2] , \ab[197][1] , \ab[197][0] ,
         \ab[196][3] , \ab[196][2] , \ab[196][1] , \ab[196][0] , \ab[195][3] ,
         \ab[195][2] , \ab[195][1] , \ab[195][0] , \ab[194][3] , \ab[194][2] ,
         \ab[194][1] , \ab[194][0] , \ab[193][3] , \ab[193][2] , \ab[193][1] ,
         \ab[193][0] , \ab[192][3] , \ab[192][2] , \ab[192][1] , \ab[192][0] ,
         \ab[191][3] , \ab[191][2] , \ab[191][1] , \ab[191][0] , \ab[190][3] ,
         \ab[190][2] , \ab[190][1] , \ab[190][0] , \ab[189][3] , \ab[189][2] ,
         \ab[189][1] , \ab[189][0] , \ab[188][3] , \ab[188][2] , \ab[188][1] ,
         \ab[188][0] , \ab[187][3] , \ab[187][2] , \ab[187][1] , \ab[187][0] ,
         \ab[186][3] , \ab[186][2] , \ab[186][1] , \ab[186][0] , \ab[185][3] ,
         \ab[185][2] , \ab[185][1] , \ab[185][0] , \ab[184][3] , \ab[184][2] ,
         \ab[184][1] , \ab[184][0] , \ab[183][3] , \ab[183][2] , \ab[183][1] ,
         \ab[183][0] , \ab[182][3] , \ab[182][2] , \ab[182][1] , \ab[182][0] ,
         \ab[181][3] , \ab[181][2] , \ab[181][1] , \ab[181][0] , \ab[180][3] ,
         \ab[180][2] , \ab[180][1] , \ab[180][0] , \ab[179][3] , \ab[179][2] ,
         \ab[179][1] , \ab[179][0] , \ab[178][3] , \ab[178][2] , \ab[178][1] ,
         \ab[178][0] , \ab[177][3] , \ab[177][2] , \ab[177][1] , \ab[177][0] ,
         \ab[176][3] , \ab[176][2] , \ab[176][1] , \ab[176][0] , \ab[175][3] ,
         \ab[175][2] , \ab[175][1] , \ab[175][0] , \ab[174][3] , \ab[174][2] ,
         \ab[174][1] , \ab[174][0] , \ab[173][3] , \ab[173][2] , \ab[173][1] ,
         \ab[173][0] , \ab[172][3] , \ab[172][2] , \ab[172][1] , \ab[172][0] ,
         \ab[171][3] , \ab[171][2] , \ab[171][1] , \ab[171][0] , \ab[170][3] ,
         \ab[170][2] , \ab[170][1] , \ab[170][0] , \ab[169][3] , \ab[169][2] ,
         \ab[169][1] , \ab[169][0] , \ab[168][3] , \ab[168][2] , \ab[168][1] ,
         \ab[168][0] , \ab[167][3] , \ab[167][2] , \ab[167][1] , \ab[167][0] ,
         \ab[166][3] , \ab[166][2] , \ab[166][1] , \ab[166][0] , \ab[165][3] ,
         \ab[165][2] , \ab[165][1] , \ab[165][0] , \ab[164][3] , \ab[164][2] ,
         \ab[164][1] , \ab[164][0] , \ab[163][3] , \ab[163][2] , \ab[163][1] ,
         \ab[163][0] , \ab[162][3] , \ab[162][2] , \ab[162][1] , \ab[162][0] ,
         \ab[161][3] , \ab[161][2] , \ab[161][1] , \ab[161][0] , \ab[160][3] ,
         \ab[160][2] , \ab[160][1] , \ab[160][0] , \ab[159][3] , \ab[159][2] ,
         \ab[159][1] , \ab[159][0] , \ab[158][3] , \ab[158][2] , \ab[158][1] ,
         \ab[158][0] , \ab[157][3] , \ab[157][2] , \ab[157][1] , \ab[157][0] ,
         \ab[156][3] , \ab[156][2] , \ab[156][1] , \ab[156][0] , \ab[155][3] ,
         \ab[155][2] , \ab[155][1] , \ab[155][0] , \ab[154][3] , \ab[154][2] ,
         \ab[154][1] , \ab[154][0] , \ab[153][3] , \ab[153][2] , \ab[153][1] ,
         \ab[153][0] , \ab[152][3] , \ab[152][2] , \ab[152][1] , \ab[152][0] ,
         \ab[151][3] , \ab[151][2] , \ab[151][1] , \ab[151][0] , \ab[150][3] ,
         \ab[150][2] , \ab[150][1] , \ab[150][0] , \ab[149][3] , \ab[149][2] ,
         \ab[149][1] , \ab[149][0] , \ab[148][3] , \ab[148][2] , \ab[148][1] ,
         \ab[148][0] , \ab[147][3] , \ab[147][2] , \ab[147][1] , \ab[147][0] ,
         \ab[146][3] , \ab[146][2] , \ab[146][1] , \ab[146][0] , \ab[145][3] ,
         \ab[145][2] , \ab[145][1] , \ab[145][0] , \ab[144][3] , \ab[144][2] ,
         \ab[144][1] , \ab[144][0] , \ab[143][3] , \ab[143][2] , \ab[143][1] ,
         \ab[143][0] , \ab[142][3] , \ab[142][2] , \ab[142][1] , \ab[142][0] ,
         \ab[141][3] , \ab[141][2] , \ab[141][1] , \ab[141][0] , \ab[140][3] ,
         \ab[140][2] , \ab[140][1] , \ab[140][0] , \ab[139][3] , \ab[139][2] ,
         \ab[139][1] , \ab[139][0] , \ab[138][3] , \ab[138][2] , \ab[138][1] ,
         \ab[138][0] , \ab[137][3] , \ab[137][2] , \ab[137][1] , \ab[137][0] ,
         \ab[136][3] , \ab[136][2] , \ab[136][1] , \ab[136][0] , \ab[135][3] ,
         \ab[135][2] , \ab[135][1] , \ab[135][0] , \ab[134][3] , \ab[134][2] ,
         \ab[134][1] , \ab[134][0] , \ab[133][3] , \ab[133][2] , \ab[133][1] ,
         \ab[133][0] , \ab[132][3] , \ab[132][2] , \ab[132][1] , \ab[132][0] ,
         \ab[131][3] , \ab[131][2] , \ab[131][1] , \ab[131][0] , \ab[130][3] ,
         \ab[130][2] , \ab[130][1] , \ab[130][0] , \ab[129][3] , \ab[129][2] ,
         \ab[129][1] , \ab[129][0] , \ab[128][3] , \ab[128][2] , \ab[128][1] ,
         \ab[128][0] , \ab[127][3] , \ab[127][2] , \ab[127][1] , \ab[127][0] ,
         \ab[126][3] , \ab[126][2] , \ab[126][1] , \ab[126][0] , \ab[125][3] ,
         \ab[125][2] , \ab[125][1] , \ab[125][0] , \ab[124][3] , \ab[124][2] ,
         \ab[124][1] , \ab[124][0] , \ab[123][3] , \ab[123][2] , \ab[123][1] ,
         \ab[123][0] , \ab[122][3] , \ab[122][2] , \ab[122][1] , \ab[122][0] ,
         \ab[121][3] , \ab[121][2] , \ab[121][1] , \ab[121][0] , \ab[120][3] ,
         \ab[120][2] , \ab[120][1] , \ab[120][0] , \ab[119][3] , \ab[119][2] ,
         \ab[119][1] , \ab[119][0] , \ab[118][3] , \ab[118][2] , \ab[118][1] ,
         \ab[118][0] , \ab[117][3] , \ab[117][2] , \ab[117][1] , \ab[117][0] ,
         \ab[116][3] , \ab[116][2] , \ab[116][1] , \ab[116][0] , \ab[115][3] ,
         \ab[115][2] , \ab[115][1] , \ab[115][0] , \ab[114][3] , \ab[114][2] ,
         \ab[114][1] , \ab[114][0] , \ab[113][3] , \ab[113][2] , \ab[113][1] ,
         \ab[113][0] , \ab[112][3] , \ab[112][2] , \ab[112][1] , \ab[112][0] ,
         \ab[111][3] , \ab[111][2] , \ab[111][1] , \ab[111][0] , \ab[110][3] ,
         \ab[110][2] , \ab[110][1] , \ab[110][0] , \ab[109][3] , \ab[109][2] ,
         \ab[109][1] , \ab[109][0] , \ab[108][3] , \ab[108][2] , \ab[108][1] ,
         \ab[108][0] , \ab[107][3] , \ab[107][2] , \ab[107][1] , \ab[107][0] ,
         \ab[106][3] , \ab[106][2] , \ab[106][1] , \ab[106][0] , \ab[105][3] ,
         \ab[105][2] , \ab[105][1] , \ab[105][0] , \ab[104][3] , \ab[104][2] ,
         \ab[104][1] , \ab[104][0] , \ab[103][3] , \ab[103][2] , \ab[103][1] ,
         \ab[103][0] , \ab[102][3] , \ab[102][2] , \ab[102][1] , \ab[102][0] ,
         \ab[101][3] , \ab[101][2] , \ab[101][1] , \ab[101][0] , \ab[100][3] ,
         \ab[100][2] , \ab[100][1] , \ab[100][0] , \ab[99][3] , \ab[99][2] ,
         \ab[99][1] , \ab[99][0] , \ab[98][3] , \ab[98][2] , \ab[98][1] ,
         \ab[98][0] , \ab[97][3] , \ab[97][2] , \ab[97][1] , \ab[97][0] ,
         \ab[96][3] , \ab[96][2] , \ab[96][1] , \ab[96][0] , \ab[95][3] ,
         \ab[95][2] , \ab[95][1] , \ab[95][0] , \ab[94][3] , \ab[94][2] ,
         \ab[94][1] , \ab[94][0] , \ab[93][3] , \ab[93][2] , \ab[93][1] ,
         \ab[93][0] , \ab[92][3] , \ab[92][2] , \ab[92][1] , \ab[92][0] ,
         \ab[91][3] , \ab[91][2] , \ab[91][1] , \ab[91][0] , \ab[90][3] ,
         \ab[90][2] , \ab[90][1] , \ab[90][0] , \ab[89][3] , \ab[89][2] ,
         \ab[89][1] , \ab[89][0] , \ab[88][3] , \ab[88][2] , \ab[88][1] ,
         \ab[88][0] , \ab[87][3] , \ab[87][2] , \ab[87][1] , \ab[87][0] ,
         \ab[86][3] , \ab[86][2] , \ab[86][1] , \ab[86][0] , \ab[85][3] ,
         \ab[85][2] , \ab[85][1] , \ab[85][0] , \ab[84][3] , \ab[84][2] ,
         \ab[84][1] , \ab[84][0] , \ab[83][3] , \ab[83][2] , \ab[83][1] ,
         \ab[83][0] , \ab[82][3] , \ab[82][2] , \ab[82][1] , \ab[82][0] ,
         \ab[81][3] , \ab[81][2] , \ab[81][1] , \ab[81][0] , \ab[80][3] ,
         \ab[80][2] , \ab[80][1] , \ab[80][0] , \ab[79][3] , \ab[79][2] ,
         \ab[79][1] , \ab[79][0] , \ab[78][3] , \ab[78][2] , \ab[78][1] ,
         \ab[78][0] , \ab[77][3] , \ab[77][2] , \ab[77][1] , \ab[77][0] ,
         \ab[76][3] , \ab[76][2] , \ab[76][1] , \ab[76][0] , \ab[75][3] ,
         \ab[75][2] , \ab[75][1] , \ab[75][0] , \ab[74][3] , \ab[74][2] ,
         \ab[74][1] , \ab[74][0] , \ab[73][3] , \ab[73][2] , \ab[73][1] ,
         \ab[73][0] , \ab[72][3] , \ab[72][2] , \ab[72][1] , \ab[72][0] ,
         \ab[71][3] , \ab[71][2] , \ab[71][1] , \ab[71][0] , \ab[70][3] ,
         \ab[70][2] , \ab[70][1] , \ab[70][0] , \ab[69][3] , \ab[69][2] ,
         \ab[69][1] , \ab[69][0] , \ab[68][3] , \ab[68][2] , \ab[68][1] ,
         \ab[68][0] , \ab[67][3] , \ab[67][2] , \ab[67][1] , \ab[67][0] ,
         \ab[66][3] , \ab[66][2] , \ab[66][1] , \ab[66][0] , \ab[65][3] ,
         \ab[65][2] , \ab[65][1] , \ab[65][0] , \ab[64][3] , \ab[64][2] ,
         \ab[64][1] , \ab[64][0] , \ab[63][3] , \ab[63][2] , \ab[63][1] ,
         \ab[63][0] , \ab[62][3] , \ab[62][2] , \ab[62][1] , \ab[62][0] ,
         \ab[61][3] , \ab[61][2] , \ab[61][1] , \ab[61][0] , \ab[60][3] ,
         \ab[60][2] , \ab[60][1] , \ab[60][0] , \ab[59][3] , \ab[59][2] ,
         \ab[59][1] , \ab[59][0] , \ab[58][3] , \ab[58][2] , \ab[58][1] ,
         \ab[58][0] , \ab[57][3] , \ab[57][2] , \ab[57][1] , \ab[57][0] ,
         \ab[56][3] , \ab[56][2] , \ab[56][1] , \ab[56][0] , \ab[55][3] ,
         \ab[55][2] , \ab[55][1] , \ab[55][0] , \ab[54][3] , \ab[54][2] ,
         \ab[54][1] , \ab[54][0] , \ab[53][3] , \ab[53][2] , \ab[53][1] ,
         \ab[53][0] , \ab[52][3] , \ab[52][2] , \ab[52][1] , \ab[52][0] ,
         \ab[51][3] , \ab[51][2] , \ab[51][1] , \ab[51][0] , \ab[50][3] ,
         \ab[50][2] , \ab[50][1] , \ab[50][0] , \ab[49][3] , \ab[49][2] ,
         \ab[49][1] , \ab[49][0] , \ab[48][3] , \ab[48][2] , \ab[48][1] ,
         \ab[48][0] , \ab[47][3] , \ab[47][2] , \ab[47][1] , \ab[47][0] ,
         \ab[46][3] , \ab[46][2] , \ab[46][1] , \ab[46][0] , \ab[45][3] ,
         \ab[45][2] , \ab[45][1] , \ab[45][0] , \ab[44][3] , \ab[44][2] ,
         \ab[44][1] , \ab[44][0] , \ab[43][3] , \ab[43][2] , \ab[43][1] ,
         \ab[43][0] , \ab[42][3] , \ab[42][2] , \ab[42][1] , \ab[42][0] ,
         \ab[41][3] , \ab[41][2] , \ab[41][1] , \ab[41][0] , \ab[40][3] ,
         \ab[40][2] , \ab[40][1] , \ab[40][0] , \ab[39][3] , \ab[39][2] ,
         \ab[39][1] , \ab[39][0] , \ab[38][3] , \ab[38][2] , \ab[38][1] ,
         \ab[38][0] , \ab[37][3] , \ab[37][2] , \ab[37][1] , \ab[37][0] ,
         \ab[36][3] , \ab[36][2] , \ab[36][1] , \ab[36][0] , \ab[35][3] ,
         \ab[35][2] , \ab[35][1] , \ab[35][0] , \ab[34][3] , \ab[34][2] ,
         \ab[34][1] , \ab[34][0] , \ab[33][3] , \ab[33][2] , \ab[33][1] ,
         \ab[33][0] , \ab[32][3] , \ab[32][2] , \ab[32][1] , \ab[32][0] ,
         \ab[31][3] , \ab[31][2] , \ab[31][1] , \ab[31][0] , \ab[30][3] ,
         \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][3] , \ab[29][2] ,
         \ab[29][1] , \ab[29][0] , \ab[28][3] , \ab[28][2] , \ab[28][1] ,
         \ab[28][0] , \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] ,
         \ab[26][3] , \ab[26][2] , \ab[26][1] , \ab[26][0] , \ab[25][3] ,
         \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][3] , \ab[24][2] ,
         \ab[24][1] , \ab[24][0] , \ab[23][3] , \ab[23][2] , \ab[23][1] ,
         \ab[23][0] , \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] ,
         \ab[21][3] , \ab[21][2] , \ab[21][1] , \ab[21][0] , \ab[20][3] ,
         \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][3] , \ab[19][2] ,
         \ab[19][1] , \ab[19][0] , \ab[18][3] , \ab[18][2] , \ab[18][1] ,
         \ab[18][0] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][3] , \ab[16][2] , \ab[16][1] , \ab[16][0] , \ab[15][3] ,
         \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][3] , \ab[13][2] , \ab[13][1] ,
         \ab[13][0] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][3] , \ab[8][2] , \ab[8][1] ,
         \ab[8][0] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[127][2] , \CARRYB[127][1] ,
         \CARRYB[127][0] , \CARRYB[126][2] , \CARRYB[126][1] ,
         \CARRYB[126][0] , \CARRYB[125][2] , \CARRYB[125][1] ,
         \CARRYB[125][0] , \CARRYB[124][2] , \CARRYB[124][1] ,
         \CARRYB[124][0] , \CARRYB[123][2] , \CARRYB[123][1] ,
         \CARRYB[123][0] , \CARRYB[122][2] , \CARRYB[122][1] ,
         \CARRYB[122][0] , \CARRYB[121][2] , \CARRYB[121][1] ,
         \CARRYB[121][0] , \CARRYB[120][2] , \CARRYB[120][1] ,
         \CARRYB[120][0] , \CARRYB[119][2] , \CARRYB[119][1] ,
         \CARRYB[119][0] , \CARRYB[118][2] , \CARRYB[118][1] ,
         \CARRYB[118][0] , \CARRYB[117][2] , \CARRYB[117][1] ,
         \CARRYB[117][0] , \CARRYB[116][2] , \CARRYB[116][1] ,
         \CARRYB[116][0] , \CARRYB[115][2] , \CARRYB[115][1] ,
         \CARRYB[115][0] , \CARRYB[114][2] , \CARRYB[114][1] ,
         \CARRYB[114][0] , \CARRYB[113][2] , \CARRYB[113][1] ,
         \CARRYB[113][0] , \CARRYB[112][2] , \CARRYB[112][1] ,
         \CARRYB[112][0] , \CARRYB[111][2] , \CARRYB[111][1] ,
         \CARRYB[111][0] , \CARRYB[110][2] , \CARRYB[110][1] ,
         \CARRYB[110][0] , \CARRYB[109][2] , \CARRYB[109][1] ,
         \CARRYB[109][0] , \CARRYB[108][2] , \CARRYB[108][1] ,
         \CARRYB[108][0] , \CARRYB[107][2] , \CARRYB[107][1] ,
         \CARRYB[107][0] , \CARRYB[106][2] , \CARRYB[106][1] ,
         \CARRYB[106][0] , \CARRYB[105][2] , \CARRYB[105][1] ,
         \CARRYB[105][0] , \CARRYB[104][2] , \CARRYB[104][1] ,
         \CARRYB[104][0] , \CARRYB[103][2] , \CARRYB[103][1] ,
         \CARRYB[103][0] , \CARRYB[102][2] , \CARRYB[102][1] ,
         \CARRYB[102][0] , \CARRYB[101][2] , \CARRYB[101][1] ,
         \CARRYB[101][0] , \CARRYB[100][2] , \CARRYB[100][1] ,
         \CARRYB[100][0] , \CARRYB[99][2] , \CARRYB[99][1] , \CARRYB[99][0] ,
         \CARRYB[98][2] , \CARRYB[98][1] , \CARRYB[98][0] , \CARRYB[97][2] ,
         \CARRYB[97][1] , \CARRYB[97][0] , \CARRYB[96][2] , \CARRYB[96][1] ,
         \CARRYB[96][0] , \CARRYB[95][2] , \CARRYB[95][1] , \CARRYB[95][0] ,
         \CARRYB[94][2] , \CARRYB[94][1] , \CARRYB[94][0] , \CARRYB[93][2] ,
         \CARRYB[93][1] , \CARRYB[93][0] , \CARRYB[92][2] , \CARRYB[92][1] ,
         \CARRYB[92][0] , \CARRYB[91][2] , \CARRYB[91][1] , \CARRYB[91][0] ,
         \CARRYB[90][2] , \CARRYB[90][1] , \CARRYB[90][0] , \CARRYB[89][2] ,
         \CARRYB[89][1] , \CARRYB[89][0] , \CARRYB[88][2] , \CARRYB[88][1] ,
         \CARRYB[88][0] , \CARRYB[87][2] , \CARRYB[87][1] , \CARRYB[87][0] ,
         \CARRYB[86][2] , \CARRYB[86][1] , \CARRYB[86][0] , \CARRYB[85][2] ,
         \CARRYB[85][1] , \CARRYB[85][0] , \CARRYB[84][2] , \CARRYB[84][1] ,
         \CARRYB[84][0] , \CARRYB[83][2] , \CARRYB[83][1] , \CARRYB[83][0] ,
         \CARRYB[82][2] , \CARRYB[82][1] , \CARRYB[82][0] , \CARRYB[81][2] ,
         \CARRYB[81][1] , \CARRYB[81][0] , \CARRYB[80][2] , \CARRYB[80][1] ,
         \CARRYB[80][0] , \CARRYB[79][2] , \CARRYB[79][1] , \CARRYB[79][0] ,
         \CARRYB[78][2] , \CARRYB[78][1] , \CARRYB[78][0] , \CARRYB[77][2] ,
         \CARRYB[77][1] , \CARRYB[77][0] , \CARRYB[76][2] , \CARRYB[76][1] ,
         \CARRYB[76][0] , \CARRYB[75][2] , \CARRYB[75][1] , \CARRYB[75][0] ,
         \CARRYB[74][2] , \CARRYB[74][1] , \CARRYB[74][0] , \CARRYB[73][2] ,
         \CARRYB[73][1] , \CARRYB[73][0] , \CARRYB[72][2] , \CARRYB[72][1] ,
         \CARRYB[72][0] , \CARRYB[71][2] , \CARRYB[71][1] , \CARRYB[71][0] ,
         \CARRYB[70][2] , \CARRYB[70][1] , \CARRYB[70][0] , \CARRYB[69][2] ,
         \CARRYB[69][1] , \CARRYB[69][0] , \CARRYB[68][2] , \CARRYB[68][1] ,
         \CARRYB[68][0] , \CARRYB[67][2] , \CARRYB[67][1] , \CARRYB[67][0] ,
         \CARRYB[66][2] , \CARRYB[66][1] , \CARRYB[66][0] , \CARRYB[65][2] ,
         \CARRYB[65][1] , \CARRYB[65][0] , \CARRYB[64][2] , \CARRYB[64][1] ,
         \CARRYB[64][0] , \CARRYB[63][2] , \CARRYB[63][1] , \CARRYB[63][0] ,
         \CARRYB[62][2] , \CARRYB[62][1] , \CARRYB[62][0] , \CARRYB[61][2] ,
         \CARRYB[61][1] , \CARRYB[61][0] , \CARRYB[60][2] , \CARRYB[60][1] ,
         \CARRYB[60][0] , \CARRYB[59][2] , \CARRYB[59][1] , \CARRYB[59][0] ,
         \CARRYB[58][2] , \CARRYB[58][1] , \CARRYB[58][0] , \CARRYB[57][2] ,
         \CARRYB[57][1] , \CARRYB[57][0] , \CARRYB[56][2] , \CARRYB[56][1] ,
         \CARRYB[56][0] , \CARRYB[55][2] , \CARRYB[55][1] , \CARRYB[55][0] ,
         \CARRYB[54][2] , \CARRYB[54][1] , \CARRYB[54][0] , \CARRYB[53][2] ,
         \CARRYB[53][1] , \CARRYB[53][0] , \CARRYB[52][2] , \CARRYB[52][1] ,
         \CARRYB[52][0] , \CARRYB[51][2] , \CARRYB[51][1] , \CARRYB[51][0] ,
         \CARRYB[50][2] , \CARRYB[50][1] , \CARRYB[50][0] , \CARRYB[49][2] ,
         \CARRYB[49][1] , \CARRYB[49][0] , \CARRYB[48][2] , \CARRYB[48][1] ,
         \CARRYB[48][0] , \CARRYB[47][2] , \CARRYB[47][1] , \CARRYB[47][0] ,
         \CARRYB[46][2] , \CARRYB[46][1] , \CARRYB[46][0] , \CARRYB[45][2] ,
         \CARRYB[45][1] , \CARRYB[45][0] , \CARRYB[44][2] , \CARRYB[44][1] ,
         \CARRYB[44][0] , \CARRYB[43][2] , \CARRYB[43][1] , \CARRYB[43][0] ,
         \CARRYB[42][2] , \CARRYB[42][1] , \CARRYB[42][0] , \CARRYB[41][2] ,
         \CARRYB[41][1] , \CARRYB[41][0] , \CARRYB[40][2] , \CARRYB[40][1] ,
         \CARRYB[40][0] , \CARRYB[39][2] , \CARRYB[39][1] , \CARRYB[39][0] ,
         \CARRYB[38][2] , \CARRYB[38][1] , \CARRYB[38][0] , \CARRYB[37][2] ,
         \CARRYB[37][1] , \CARRYB[37][0] , \CARRYB[36][2] , \CARRYB[36][1] ,
         \CARRYB[36][0] , \CARRYB[35][2] , \CARRYB[35][1] , \CARRYB[35][0] ,
         \CARRYB[34][2] , \CARRYB[34][1] , \CARRYB[34][0] , \CARRYB[33][2] ,
         \CARRYB[33][1] , \CARRYB[33][0] , \CARRYB[32][2] , \CARRYB[32][1] ,
         \CARRYB[32][0] , \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] ,
         \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] , \CARRYB[29][2] ,
         \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] ,
         \CARRYB[26][2] , \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][2] ,
         \CARRYB[25][1] , \CARRYB[25][0] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][2] ,
         \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] ,
         \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][2] ,
         \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][2] ,
         \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[127][2] , \SUMB[127][1] ,
         \SUMB[126][2] , \SUMB[126][1] , \SUMB[125][2] , \SUMB[125][1] ,
         \SUMB[124][2] , \SUMB[124][1] , \SUMB[123][2] , \SUMB[123][1] ,
         \SUMB[122][2] , \SUMB[122][1] , \SUMB[121][2] , \SUMB[121][1] ,
         \SUMB[120][2] , \SUMB[120][1] , \SUMB[119][2] , \SUMB[119][1] ,
         \SUMB[118][2] , \SUMB[118][1] , \SUMB[117][2] , \SUMB[117][1] ,
         \SUMB[116][2] , \SUMB[116][1] , \SUMB[115][2] , \SUMB[115][1] ,
         \SUMB[114][2] , \SUMB[114][1] , \SUMB[113][2] , \SUMB[113][1] ,
         \SUMB[112][2] , \SUMB[112][1] , \SUMB[111][2] , \SUMB[111][1] ,
         \SUMB[110][2] , \SUMB[110][1] , \SUMB[109][2] , \SUMB[109][1] ,
         \SUMB[108][2] , \SUMB[108][1] , \SUMB[107][2] , \SUMB[107][1] ,
         \SUMB[106][2] , \SUMB[106][1] , \SUMB[105][2] , \SUMB[105][1] ,
         \SUMB[104][2] , \SUMB[104][1] , \SUMB[103][2] , \SUMB[103][1] ,
         \SUMB[102][2] , \SUMB[102][1] , \SUMB[101][2] , \SUMB[101][1] ,
         \SUMB[100][2] , \SUMB[100][1] , \SUMB[99][2] , \SUMB[99][1] ,
         \SUMB[98][2] , \SUMB[98][1] , \SUMB[97][2] , \SUMB[97][1] ,
         \SUMB[96][2] , \SUMB[96][1] , \SUMB[95][2] , \SUMB[95][1] ,
         \SUMB[94][2] , \SUMB[94][1] , \SUMB[93][2] , \SUMB[93][1] ,
         \SUMB[92][2] , \SUMB[92][1] , \SUMB[91][2] , \SUMB[91][1] ,
         \SUMB[90][2] , \SUMB[90][1] , \SUMB[89][2] , \SUMB[89][1] ,
         \SUMB[88][2] , \SUMB[88][1] , \SUMB[87][2] , \SUMB[87][1] ,
         \SUMB[86][2] , \SUMB[86][1] , \SUMB[85][2] , \SUMB[85][1] ,
         \SUMB[84][2] , \SUMB[84][1] , \SUMB[83][2] , \SUMB[83][1] ,
         \SUMB[82][2] , \SUMB[82][1] , \SUMB[81][2] , \SUMB[81][1] ,
         \SUMB[80][2] , \SUMB[80][1] , \SUMB[79][2] , \SUMB[79][1] ,
         \SUMB[78][2] , \SUMB[78][1] , \SUMB[77][2] , \SUMB[77][1] ,
         \SUMB[76][2] , \SUMB[76][1] , \SUMB[75][2] , \SUMB[75][1] ,
         \SUMB[74][2] , \SUMB[74][1] , \SUMB[73][2] , \SUMB[73][1] ,
         \SUMB[72][2] , \SUMB[72][1] , \SUMB[71][2] , \SUMB[71][1] ,
         \SUMB[70][2] , \SUMB[70][1] , \SUMB[69][2] , \SUMB[69][1] ,
         \SUMB[68][2] , \SUMB[68][1] , \SUMB[67][2] , \SUMB[67][1] ,
         \SUMB[66][2] , \SUMB[66][1] , \SUMB[65][2] , \SUMB[65][1] ,
         \SUMB[64][2] , \SUMB[64][1] , \SUMB[63][2] , \SUMB[63][1] ,
         \SUMB[62][2] , \SUMB[62][1] , \SUMB[61][2] , \SUMB[61][1] ,
         \SUMB[60][2] , \SUMB[60][1] , \SUMB[59][2] , \SUMB[59][1] ,
         \SUMB[58][2] , \SUMB[58][1] , \SUMB[57][2] , \SUMB[57][1] ,
         \SUMB[56][2] , \SUMB[56][1] , \SUMB[55][2] , \SUMB[55][1] ,
         \SUMB[54][2] , \SUMB[54][1] , \SUMB[53][2] , \SUMB[53][1] ,
         \SUMB[52][2] , \SUMB[52][1] , \SUMB[51][2] , \SUMB[51][1] ,
         \SUMB[50][2] , \SUMB[50][1] , \SUMB[49][2] , \SUMB[49][1] ,
         \SUMB[48][2] , \SUMB[48][1] , \SUMB[47][2] , \SUMB[47][1] ,
         \SUMB[46][2] , \SUMB[46][1] , \SUMB[45][2] , \SUMB[45][1] ,
         \SUMB[44][2] , \SUMB[44][1] , \SUMB[43][2] , \SUMB[43][1] ,
         \SUMB[42][2] , \SUMB[42][1] , \SUMB[41][2] , \SUMB[41][1] ,
         \SUMB[40][2] , \SUMB[40][1] , \SUMB[39][2] , \SUMB[39][1] ,
         \SUMB[38][2] , \SUMB[38][1] , \SUMB[37][2] , \SUMB[37][1] ,
         \SUMB[36][2] , \SUMB[36][1] , \SUMB[35][2] , \SUMB[35][1] ,
         \SUMB[34][2] , \SUMB[34][1] , \SUMB[33][2] , \SUMB[33][1] ,
         \SUMB[32][2] , \SUMB[32][1] , \SUMB[31][2] , \SUMB[31][1] ,
         \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][2] , \SUMB[29][1] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][2] , \SUMB[27][1] ,
         \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][2] , \SUMB[25][1] ,
         \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][2] , \SUMB[23][1] ,
         \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][2] , \SUMB[21][1] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][2] , \SUMB[19][1] ,
         \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][2] , \SUMB[17][1] ,
         \SUMB[16][2] , \SUMB[16][1] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][2] , \SUMB[11][1] ,
         \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][2] ,
         \SUMB[6][1] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][2] ,
         \SUMB[1][1] , \CARRYB[255][2] , \CARRYB[255][1] , \CARRYB[255][0] ,
         \CARRYB[254][2] , \CARRYB[254][1] , \CARRYB[254][0] ,
         \CARRYB[253][2] , \CARRYB[253][1] , \CARRYB[253][0] ,
         \CARRYB[252][2] , \CARRYB[252][1] , \CARRYB[252][0] ,
         \CARRYB[251][2] , \CARRYB[251][1] , \CARRYB[251][0] ,
         \CARRYB[250][2] , \CARRYB[250][1] , \CARRYB[250][0] ,
         \CARRYB[249][2] , \CARRYB[249][1] , \CARRYB[249][0] ,
         \CARRYB[248][2] , \CARRYB[248][1] , \CARRYB[248][0] ,
         \CARRYB[247][2] , \CARRYB[247][1] , \CARRYB[247][0] ,
         \CARRYB[246][2] , \CARRYB[246][1] , \CARRYB[246][0] ,
         \CARRYB[245][2] , \CARRYB[245][1] , \CARRYB[245][0] ,
         \CARRYB[244][2] , \CARRYB[244][1] , \CARRYB[244][0] ,
         \CARRYB[243][2] , \CARRYB[243][1] , \CARRYB[243][0] ,
         \CARRYB[242][2] , \CARRYB[242][1] , \CARRYB[242][0] ,
         \CARRYB[241][2] , \CARRYB[241][1] , \CARRYB[241][0] ,
         \CARRYB[240][2] , \CARRYB[240][1] , \CARRYB[240][0] ,
         \CARRYB[239][2] , \CARRYB[239][1] , \CARRYB[239][0] ,
         \CARRYB[238][2] , \CARRYB[238][1] , \CARRYB[238][0] ,
         \CARRYB[237][2] , \CARRYB[237][1] , \CARRYB[237][0] ,
         \CARRYB[236][2] , \CARRYB[236][1] , \CARRYB[236][0] ,
         \CARRYB[235][2] , \CARRYB[235][1] , \CARRYB[235][0] ,
         \CARRYB[234][2] , \CARRYB[234][1] , \CARRYB[234][0] ,
         \CARRYB[233][2] , \CARRYB[233][1] , \CARRYB[233][0] ,
         \CARRYB[232][2] , \CARRYB[232][1] , \CARRYB[232][0] ,
         \CARRYB[231][2] , \CARRYB[231][1] , \CARRYB[231][0] ,
         \CARRYB[230][2] , \CARRYB[230][1] , \CARRYB[230][0] ,
         \CARRYB[229][2] , \CARRYB[229][1] , \CARRYB[229][0] ,
         \CARRYB[228][2] , \CARRYB[228][1] , \CARRYB[228][0] ,
         \CARRYB[227][2] , \CARRYB[227][1] , \CARRYB[227][0] ,
         \CARRYB[226][2] , \CARRYB[226][1] , \CARRYB[226][0] ,
         \CARRYB[225][2] , \CARRYB[225][1] , \CARRYB[225][0] ,
         \CARRYB[224][2] , \CARRYB[224][1] , \CARRYB[224][0] ,
         \CARRYB[223][2] , \CARRYB[223][1] , \CARRYB[223][0] ,
         \CARRYB[222][2] , \CARRYB[222][1] , \CARRYB[222][0] ,
         \CARRYB[221][2] , \CARRYB[221][1] , \CARRYB[221][0] ,
         \CARRYB[220][2] , \CARRYB[220][1] , \CARRYB[220][0] ,
         \CARRYB[219][2] , \CARRYB[219][1] , \CARRYB[219][0] ,
         \CARRYB[218][2] , \CARRYB[218][1] , \CARRYB[218][0] ,
         \CARRYB[217][2] , \CARRYB[217][1] , \CARRYB[217][0] ,
         \CARRYB[216][2] , \CARRYB[216][1] , \CARRYB[216][0] ,
         \CARRYB[215][2] , \CARRYB[215][1] , \CARRYB[215][0] ,
         \CARRYB[214][2] , \CARRYB[214][1] , \CARRYB[214][0] ,
         \CARRYB[213][2] , \CARRYB[213][1] , \CARRYB[213][0] ,
         \CARRYB[212][2] , \CARRYB[212][1] , \CARRYB[212][0] ,
         \CARRYB[211][2] , \CARRYB[211][1] , \CARRYB[211][0] ,
         \CARRYB[210][2] , \CARRYB[210][1] , \CARRYB[210][0] ,
         \CARRYB[209][2] , \CARRYB[209][1] , \CARRYB[209][0] ,
         \CARRYB[208][2] , \CARRYB[208][1] , \CARRYB[208][0] ,
         \CARRYB[207][2] , \CARRYB[207][1] , \CARRYB[207][0] ,
         \CARRYB[206][2] , \CARRYB[206][1] , \CARRYB[206][0] ,
         \CARRYB[205][2] , \CARRYB[205][1] , \CARRYB[205][0] ,
         \CARRYB[204][2] , \CARRYB[204][1] , \CARRYB[204][0] ,
         \CARRYB[203][2] , \CARRYB[203][1] , \CARRYB[203][0] ,
         \CARRYB[202][2] , \CARRYB[202][1] , \CARRYB[202][0] ,
         \CARRYB[201][2] , \CARRYB[201][1] , \CARRYB[201][0] ,
         \CARRYB[200][2] , \CARRYB[200][1] , \CARRYB[200][0] ,
         \CARRYB[199][2] , \CARRYB[199][1] , \CARRYB[199][0] ,
         \CARRYB[198][2] , \CARRYB[198][1] , \CARRYB[198][0] ,
         \CARRYB[197][2] , \CARRYB[197][1] , \CARRYB[197][0] ,
         \CARRYB[196][2] , \CARRYB[196][1] , \CARRYB[196][0] ,
         \CARRYB[195][2] , \CARRYB[195][1] , \CARRYB[195][0] ,
         \CARRYB[194][2] , \CARRYB[194][1] , \CARRYB[194][0] ,
         \CARRYB[193][2] , \CARRYB[193][1] , \CARRYB[193][0] ,
         \CARRYB[192][2] , \CARRYB[192][1] , \CARRYB[192][0] ,
         \CARRYB[191][2] , \CARRYB[191][1] , \CARRYB[191][0] ,
         \CARRYB[190][2] , \CARRYB[190][1] , \CARRYB[190][0] ,
         \CARRYB[189][2] , \CARRYB[189][1] , \CARRYB[189][0] ,
         \CARRYB[188][2] , \CARRYB[188][1] , \CARRYB[188][0] ,
         \CARRYB[187][2] , \CARRYB[187][1] , \CARRYB[187][0] ,
         \CARRYB[186][2] , \CARRYB[186][1] , \CARRYB[186][0] ,
         \CARRYB[185][2] , \CARRYB[185][1] , \CARRYB[185][0] ,
         \CARRYB[184][2] , \CARRYB[184][1] , \CARRYB[184][0] ,
         \CARRYB[183][2] , \CARRYB[183][1] , \CARRYB[183][0] ,
         \CARRYB[182][2] , \CARRYB[182][1] , \CARRYB[182][0] ,
         \CARRYB[181][2] , \CARRYB[181][1] , \CARRYB[181][0] ,
         \CARRYB[180][2] , \CARRYB[180][1] , \CARRYB[180][0] ,
         \CARRYB[179][2] , \CARRYB[179][1] , \CARRYB[179][0] ,
         \CARRYB[178][2] , \CARRYB[178][1] , \CARRYB[178][0] ,
         \CARRYB[177][2] , \CARRYB[177][1] , \CARRYB[177][0] ,
         \CARRYB[176][2] , \CARRYB[176][1] , \CARRYB[176][0] ,
         \CARRYB[175][2] , \CARRYB[175][1] , \CARRYB[175][0] ,
         \CARRYB[174][2] , \CARRYB[174][1] , \CARRYB[174][0] ,
         \CARRYB[173][2] , \CARRYB[173][1] , \CARRYB[173][0] ,
         \CARRYB[172][2] , \CARRYB[172][1] , \CARRYB[172][0] ,
         \CARRYB[171][2] , \CARRYB[171][1] , \CARRYB[171][0] ,
         \CARRYB[170][2] , \CARRYB[170][1] , \CARRYB[170][0] ,
         \CARRYB[169][2] , \CARRYB[169][1] , \CARRYB[169][0] ,
         \CARRYB[168][2] , \CARRYB[168][1] , \CARRYB[168][0] ,
         \CARRYB[167][2] , \CARRYB[167][1] , \CARRYB[167][0] ,
         \CARRYB[166][2] , \CARRYB[166][1] , \CARRYB[166][0] ,
         \CARRYB[165][2] , \CARRYB[165][1] , \CARRYB[165][0] ,
         \CARRYB[164][2] , \CARRYB[164][1] , \CARRYB[164][0] ,
         \CARRYB[163][2] , \CARRYB[163][1] , \CARRYB[163][0] ,
         \CARRYB[162][2] , \CARRYB[162][1] , \CARRYB[162][0] ,
         \CARRYB[161][2] , \CARRYB[161][1] , \CARRYB[161][0] ,
         \CARRYB[160][2] , \CARRYB[160][1] , \CARRYB[160][0] ,
         \CARRYB[159][2] , \CARRYB[159][1] , \CARRYB[159][0] ,
         \CARRYB[158][2] , \CARRYB[158][1] , \CARRYB[158][0] ,
         \CARRYB[157][2] , \CARRYB[157][1] , \CARRYB[157][0] ,
         \CARRYB[156][2] , \CARRYB[156][1] , \CARRYB[156][0] ,
         \CARRYB[155][2] , \CARRYB[155][1] , \CARRYB[155][0] ,
         \CARRYB[154][2] , \CARRYB[154][1] , \CARRYB[154][0] ,
         \CARRYB[153][2] , \CARRYB[153][1] , \CARRYB[153][0] ,
         \CARRYB[152][2] , \CARRYB[152][1] , \CARRYB[152][0] ,
         \CARRYB[151][2] , \CARRYB[151][1] , \CARRYB[151][0] ,
         \CARRYB[150][2] , \CARRYB[150][1] , \CARRYB[150][0] ,
         \CARRYB[149][2] , \CARRYB[149][1] , \CARRYB[149][0] ,
         \CARRYB[148][2] , \CARRYB[148][1] , \CARRYB[148][0] ,
         \CARRYB[147][2] , \CARRYB[147][1] , \CARRYB[147][0] ,
         \CARRYB[146][2] , \CARRYB[146][1] , \CARRYB[146][0] ,
         \CARRYB[145][2] , \CARRYB[145][1] , \CARRYB[145][0] ,
         \CARRYB[144][2] , \CARRYB[144][1] , \CARRYB[144][0] ,
         \CARRYB[143][2] , \CARRYB[143][1] , \CARRYB[143][0] ,
         \CARRYB[142][2] , \CARRYB[142][1] , \CARRYB[142][0] ,
         \CARRYB[141][2] , \CARRYB[141][1] , \CARRYB[141][0] ,
         \CARRYB[140][2] , \CARRYB[140][1] , \CARRYB[140][0] ,
         \CARRYB[139][2] , \CARRYB[139][1] , \CARRYB[139][0] ,
         \CARRYB[138][2] , \CARRYB[138][1] , \CARRYB[138][0] ,
         \CARRYB[137][2] , \CARRYB[137][1] , \CARRYB[137][0] ,
         \CARRYB[136][2] , \CARRYB[136][1] , \CARRYB[136][0] ,
         \CARRYB[135][2] , \CARRYB[135][1] , \CARRYB[135][0] ,
         \CARRYB[134][2] , \CARRYB[134][1] , \CARRYB[134][0] ,
         \CARRYB[133][2] , \CARRYB[133][1] , \CARRYB[133][0] ,
         \CARRYB[132][2] , \CARRYB[132][1] , \CARRYB[132][0] ,
         \CARRYB[131][2] , \CARRYB[131][1] , \CARRYB[131][0] ,
         \CARRYB[130][2] , \CARRYB[130][1] , \CARRYB[130][0] ,
         \CARRYB[129][2] , \CARRYB[129][1] , \CARRYB[129][0] ,
         \CARRYB[128][2] , \CARRYB[128][1] , \CARRYB[128][0] , \SUMB[255][2] ,
         \SUMB[255][1] , \SUMB[254][2] , \SUMB[254][1] , \SUMB[253][2] ,
         \SUMB[253][1] , \SUMB[252][2] , \SUMB[252][1] , \SUMB[251][2] ,
         \SUMB[251][1] , \SUMB[250][2] , \SUMB[250][1] , \SUMB[249][2] ,
         \SUMB[249][1] , \SUMB[248][2] , \SUMB[248][1] , \SUMB[247][2] ,
         \SUMB[247][1] , \SUMB[246][2] , \SUMB[246][1] , \SUMB[245][2] ,
         \SUMB[245][1] , \SUMB[244][2] , \SUMB[244][1] , \SUMB[243][2] ,
         \SUMB[243][1] , \SUMB[242][2] , \SUMB[242][1] , \SUMB[241][2] ,
         \SUMB[241][1] , \SUMB[240][2] , \SUMB[240][1] , \SUMB[239][2] ,
         \SUMB[239][1] , \SUMB[238][2] , \SUMB[238][1] , \SUMB[237][2] ,
         \SUMB[237][1] , \SUMB[236][2] , \SUMB[236][1] , \SUMB[235][2] ,
         \SUMB[235][1] , \SUMB[234][2] , \SUMB[234][1] , \SUMB[233][2] ,
         \SUMB[233][1] , \SUMB[232][2] , \SUMB[232][1] , \SUMB[231][2] ,
         \SUMB[231][1] , \SUMB[230][2] , \SUMB[230][1] , \SUMB[229][2] ,
         \SUMB[229][1] , \SUMB[228][2] , \SUMB[228][1] , \SUMB[227][2] ,
         \SUMB[227][1] , \SUMB[226][2] , \SUMB[226][1] , \SUMB[225][2] ,
         \SUMB[225][1] , \SUMB[224][2] , \SUMB[224][1] , \SUMB[223][2] ,
         \SUMB[223][1] , \SUMB[222][2] , \SUMB[222][1] , \SUMB[221][2] ,
         \SUMB[221][1] , \SUMB[220][2] , \SUMB[220][1] , \SUMB[219][2] ,
         \SUMB[219][1] , \SUMB[218][2] , \SUMB[218][1] , \SUMB[217][2] ,
         \SUMB[217][1] , \SUMB[216][2] , \SUMB[216][1] , \SUMB[215][2] ,
         \SUMB[215][1] , \SUMB[214][2] , \SUMB[214][1] , \SUMB[213][2] ,
         \SUMB[213][1] , \SUMB[212][2] , \SUMB[212][1] , \SUMB[211][2] ,
         \SUMB[211][1] , \SUMB[210][2] , \SUMB[210][1] , \SUMB[209][2] ,
         \SUMB[209][1] , \SUMB[208][2] , \SUMB[208][1] , \SUMB[207][2] ,
         \SUMB[207][1] , \SUMB[206][2] , \SUMB[206][1] , \SUMB[205][2] ,
         \SUMB[205][1] , \SUMB[204][2] , \SUMB[204][1] , \SUMB[203][2] ,
         \SUMB[203][1] , \SUMB[202][2] , \SUMB[202][1] , \SUMB[201][2] ,
         \SUMB[201][1] , \SUMB[200][2] , \SUMB[200][1] , \SUMB[199][2] ,
         \SUMB[199][1] , \SUMB[198][2] , \SUMB[198][1] , \SUMB[197][2] ,
         \SUMB[197][1] , \SUMB[196][2] , \SUMB[196][1] , \SUMB[195][2] ,
         \SUMB[195][1] , \SUMB[194][2] , \SUMB[194][1] , \SUMB[193][2] ,
         \SUMB[193][1] , \SUMB[192][2] , \SUMB[192][1] , \SUMB[191][2] ,
         \SUMB[191][1] , \SUMB[190][2] , \SUMB[190][1] , \SUMB[189][2] ,
         \SUMB[189][1] , \SUMB[188][2] , \SUMB[188][1] , \SUMB[187][2] ,
         \SUMB[187][1] , \SUMB[186][2] , \SUMB[186][1] , \SUMB[185][2] ,
         \SUMB[185][1] , \SUMB[184][2] , \SUMB[184][1] , \SUMB[183][2] ,
         \SUMB[183][1] , \SUMB[182][2] , \SUMB[182][1] , \SUMB[181][2] ,
         \SUMB[181][1] , \SUMB[180][2] , \SUMB[180][1] , \SUMB[179][2] ,
         \SUMB[179][1] , \SUMB[178][2] , \SUMB[178][1] , \SUMB[177][2] ,
         \SUMB[177][1] , \SUMB[176][2] , \SUMB[176][1] , \SUMB[175][2] ,
         \SUMB[175][1] , \SUMB[174][2] , \SUMB[174][1] , \SUMB[173][2] ,
         \SUMB[173][1] , \SUMB[172][2] , \SUMB[172][1] , \SUMB[171][2] ,
         \SUMB[171][1] , \SUMB[170][2] , \SUMB[170][1] , \SUMB[169][2] ,
         \SUMB[169][1] , \SUMB[168][2] , \SUMB[168][1] , \SUMB[167][2] ,
         \SUMB[167][1] , \SUMB[166][2] , \SUMB[166][1] , \SUMB[165][2] ,
         \SUMB[165][1] , \SUMB[164][2] , \SUMB[164][1] , \SUMB[163][2] ,
         \SUMB[163][1] , \SUMB[162][2] , \SUMB[162][1] , \SUMB[161][2] ,
         \SUMB[161][1] , \SUMB[160][2] , \SUMB[160][1] , \SUMB[159][2] ,
         \SUMB[159][1] , \SUMB[158][2] , \SUMB[158][1] , \SUMB[157][2] ,
         \SUMB[157][1] , \SUMB[156][2] , \SUMB[156][1] , \SUMB[155][2] ,
         \SUMB[155][1] , \SUMB[154][2] , \SUMB[154][1] , \SUMB[153][2] ,
         \SUMB[153][1] , \SUMB[152][2] , \SUMB[152][1] , \SUMB[151][2] ,
         \SUMB[151][1] , \SUMB[150][2] , \SUMB[150][1] , \SUMB[149][2] ,
         \SUMB[149][1] , \SUMB[148][2] , \SUMB[148][1] , \SUMB[147][2] ,
         \SUMB[147][1] , \SUMB[146][2] , \SUMB[146][1] , \SUMB[145][2] ,
         \SUMB[145][1] , \SUMB[144][2] , \SUMB[144][1] , \SUMB[143][2] ,
         \SUMB[143][1] , \SUMB[142][2] , \SUMB[142][1] , \SUMB[141][2] ,
         \SUMB[141][1] , \SUMB[140][2] , \SUMB[140][1] , \SUMB[139][2] ,
         \SUMB[139][1] , \SUMB[138][2] , \SUMB[138][1] , \SUMB[137][2] ,
         \SUMB[137][1] , \SUMB[136][2] , \SUMB[136][1] , \SUMB[135][2] ,
         \SUMB[135][1] , \SUMB[134][2] , \SUMB[134][1] , \SUMB[133][2] ,
         \SUMB[133][1] , \SUMB[132][2] , \SUMB[132][1] , \SUMB[131][2] ,
         \SUMB[131][1] , \SUMB[130][2] , \SUMB[130][1] , \SUMB[129][2] ,
         \SUMB[129][1] , \SUMB[128][2] , \SUMB[128][1] , \CARRYB[383][2] ,
         \CARRYB[383][1] , \CARRYB[383][0] , \CARRYB[382][2] ,
         \CARRYB[382][1] , \CARRYB[382][0] , \CARRYB[381][2] ,
         \CARRYB[381][1] , \CARRYB[381][0] , \CARRYB[380][2] ,
         \CARRYB[380][1] , \CARRYB[380][0] , \CARRYB[379][2] ,
         \CARRYB[379][1] , \CARRYB[379][0] , \CARRYB[378][2] ,
         \CARRYB[378][1] , \CARRYB[378][0] , \CARRYB[377][2] ,
         \CARRYB[377][1] , \CARRYB[377][0] , \CARRYB[376][2] ,
         \CARRYB[376][1] , \CARRYB[376][0] , \CARRYB[375][2] ,
         \CARRYB[375][1] , \CARRYB[375][0] , \CARRYB[374][2] ,
         \CARRYB[374][1] , \CARRYB[374][0] , \CARRYB[373][2] ,
         \CARRYB[373][1] , \CARRYB[373][0] , \CARRYB[372][2] ,
         \CARRYB[372][1] , \CARRYB[372][0] , \CARRYB[371][2] ,
         \CARRYB[371][1] , \CARRYB[371][0] , \CARRYB[370][2] ,
         \CARRYB[370][1] , \CARRYB[370][0] , \CARRYB[369][2] ,
         \CARRYB[369][1] , \CARRYB[369][0] , \CARRYB[368][2] ,
         \CARRYB[368][1] , \CARRYB[368][0] , \CARRYB[367][2] ,
         \CARRYB[367][1] , \CARRYB[367][0] , \CARRYB[366][2] ,
         \CARRYB[366][1] , \CARRYB[366][0] , \CARRYB[365][2] ,
         \CARRYB[365][1] , \CARRYB[365][0] , \CARRYB[364][2] ,
         \CARRYB[364][1] , \CARRYB[364][0] , \CARRYB[363][2] ,
         \CARRYB[363][1] , \CARRYB[363][0] , \CARRYB[362][2] ,
         \CARRYB[362][1] , \CARRYB[362][0] , \CARRYB[361][2] ,
         \CARRYB[361][1] , \CARRYB[361][0] , \CARRYB[360][2] ,
         \CARRYB[360][1] , \CARRYB[360][0] , \CARRYB[359][2] ,
         \CARRYB[359][1] , \CARRYB[359][0] , \CARRYB[358][2] ,
         \CARRYB[358][1] , \CARRYB[358][0] , \CARRYB[357][2] ,
         \CARRYB[357][1] , \CARRYB[357][0] , \CARRYB[356][2] ,
         \CARRYB[356][1] , \CARRYB[356][0] , \CARRYB[355][2] ,
         \CARRYB[355][1] , \CARRYB[355][0] , \CARRYB[354][2] ,
         \CARRYB[354][1] , \CARRYB[354][0] , \CARRYB[353][2] ,
         \CARRYB[353][1] , \CARRYB[353][0] , \CARRYB[352][2] ,
         \CARRYB[352][1] , \CARRYB[352][0] , \CARRYB[351][2] ,
         \CARRYB[351][1] , \CARRYB[351][0] , \CARRYB[350][2] ,
         \CARRYB[350][1] , \CARRYB[350][0] , \CARRYB[349][2] ,
         \CARRYB[349][1] , \CARRYB[349][0] , \CARRYB[348][2] ,
         \CARRYB[348][1] , \CARRYB[348][0] , \CARRYB[347][2] ,
         \CARRYB[347][1] , \CARRYB[347][0] , \CARRYB[346][2] ,
         \CARRYB[346][1] , \CARRYB[346][0] , \CARRYB[345][2] ,
         \CARRYB[345][1] , \CARRYB[345][0] , \CARRYB[344][2] ,
         \CARRYB[344][1] , \CARRYB[344][0] , \CARRYB[343][2] ,
         \CARRYB[343][1] , \CARRYB[343][0] , \CARRYB[342][2] ,
         \CARRYB[342][1] , \CARRYB[342][0] , \CARRYB[341][2] ,
         \CARRYB[341][1] , \CARRYB[341][0] , \CARRYB[340][2] ,
         \CARRYB[340][1] , \CARRYB[340][0] , \CARRYB[339][2] ,
         \CARRYB[339][1] , \CARRYB[339][0] , \CARRYB[338][2] ,
         \CARRYB[338][1] , \CARRYB[338][0] , \CARRYB[337][2] ,
         \CARRYB[337][1] , \CARRYB[337][0] , \CARRYB[336][2] ,
         \CARRYB[336][1] , \CARRYB[336][0] , \CARRYB[335][2] ,
         \CARRYB[335][1] , \CARRYB[335][0] , \CARRYB[334][2] ,
         \CARRYB[334][1] , \CARRYB[334][0] , \CARRYB[333][2] ,
         \CARRYB[333][1] , \CARRYB[333][0] , \CARRYB[332][2] ,
         \CARRYB[332][1] , \CARRYB[332][0] , \CARRYB[331][2] ,
         \CARRYB[331][1] , \CARRYB[331][0] , \CARRYB[330][2] ,
         \CARRYB[330][1] , \CARRYB[330][0] , \CARRYB[329][2] ,
         \CARRYB[329][1] , \CARRYB[329][0] , \CARRYB[328][2] ,
         \CARRYB[328][1] , \CARRYB[328][0] , \CARRYB[327][2] ,
         \CARRYB[327][1] , \CARRYB[327][0] , \CARRYB[326][2] ,
         \CARRYB[326][1] , \CARRYB[326][0] , \CARRYB[325][2] ,
         \CARRYB[325][1] , \CARRYB[325][0] , \CARRYB[324][2] ,
         \CARRYB[324][1] , \CARRYB[324][0] , \CARRYB[323][2] ,
         \CARRYB[323][1] , \CARRYB[323][0] , \CARRYB[322][2] ,
         \CARRYB[322][1] , \CARRYB[322][0] , \CARRYB[321][2] ,
         \CARRYB[321][1] , \CARRYB[321][0] , \CARRYB[320][2] ,
         \CARRYB[320][1] , \CARRYB[320][0] , \CARRYB[319][2] ,
         \CARRYB[319][1] , \CARRYB[319][0] , \CARRYB[318][2] ,
         \CARRYB[318][1] , \CARRYB[318][0] , \CARRYB[317][2] ,
         \CARRYB[317][1] , \CARRYB[317][0] , \CARRYB[316][2] ,
         \CARRYB[316][1] , \CARRYB[316][0] , \CARRYB[315][2] ,
         \CARRYB[315][1] , \CARRYB[315][0] , \CARRYB[314][2] ,
         \CARRYB[314][1] , \CARRYB[314][0] , \CARRYB[313][2] ,
         \CARRYB[313][1] , \CARRYB[313][0] , \CARRYB[312][2] ,
         \CARRYB[312][1] , \CARRYB[312][0] , \CARRYB[311][2] ,
         \CARRYB[311][1] , \CARRYB[311][0] , \CARRYB[310][2] ,
         \CARRYB[310][1] , \CARRYB[310][0] , \CARRYB[309][2] ,
         \CARRYB[309][1] , \CARRYB[309][0] , \CARRYB[308][2] ,
         \CARRYB[308][1] , \CARRYB[308][0] , \CARRYB[307][2] ,
         \CARRYB[307][1] , \CARRYB[307][0] , \CARRYB[306][2] ,
         \CARRYB[306][1] , \CARRYB[306][0] , \CARRYB[305][2] ,
         \CARRYB[305][1] , \CARRYB[305][0] , \CARRYB[304][2] ,
         \CARRYB[304][1] , \CARRYB[304][0] , \CARRYB[303][2] ,
         \CARRYB[303][1] , \CARRYB[303][0] , \CARRYB[302][2] ,
         \CARRYB[302][1] , \CARRYB[302][0] , \CARRYB[301][2] ,
         \CARRYB[301][1] , \CARRYB[301][0] , \CARRYB[300][2] ,
         \CARRYB[300][1] , \CARRYB[300][0] , \CARRYB[299][2] ,
         \CARRYB[299][1] , \CARRYB[299][0] , \CARRYB[298][2] ,
         \CARRYB[298][1] , \CARRYB[298][0] , \CARRYB[297][2] ,
         \CARRYB[297][1] , \CARRYB[297][0] , \CARRYB[296][2] ,
         \CARRYB[296][1] , \CARRYB[296][0] , \CARRYB[295][2] ,
         \CARRYB[295][1] , \CARRYB[295][0] , \CARRYB[294][2] ,
         \CARRYB[294][1] , \CARRYB[294][0] , \CARRYB[293][2] ,
         \CARRYB[293][1] , \CARRYB[293][0] , \CARRYB[292][2] ,
         \CARRYB[292][1] , \CARRYB[292][0] , \CARRYB[291][2] ,
         \CARRYB[291][1] , \CARRYB[291][0] , \CARRYB[290][2] ,
         \CARRYB[290][1] , \CARRYB[290][0] , \CARRYB[289][2] ,
         \CARRYB[289][1] , \CARRYB[289][0] , \CARRYB[288][2] ,
         \CARRYB[288][1] , \CARRYB[288][0] , \CARRYB[287][2] ,
         \CARRYB[287][1] , \CARRYB[287][0] , \CARRYB[286][2] ,
         \CARRYB[286][1] , \CARRYB[286][0] , \CARRYB[285][2] ,
         \CARRYB[285][1] , \CARRYB[285][0] , \CARRYB[284][2] ,
         \CARRYB[284][1] , \CARRYB[284][0] , \CARRYB[283][2] ,
         \CARRYB[283][1] , \CARRYB[283][0] , \CARRYB[282][2] ,
         \CARRYB[282][1] , \CARRYB[282][0] , \CARRYB[281][2] ,
         \CARRYB[281][1] , \CARRYB[281][0] , \CARRYB[280][2] ,
         \CARRYB[280][1] , \CARRYB[280][0] , \CARRYB[279][2] ,
         \CARRYB[279][1] , \CARRYB[279][0] , \CARRYB[278][2] ,
         \CARRYB[278][1] , \CARRYB[278][0] , \CARRYB[277][2] ,
         \CARRYB[277][1] , \CARRYB[277][0] , \CARRYB[276][2] ,
         \CARRYB[276][1] , \CARRYB[276][0] , \CARRYB[275][2] ,
         \CARRYB[275][1] , \CARRYB[275][0] , \CARRYB[274][2] ,
         \CARRYB[274][1] , \CARRYB[274][0] , \CARRYB[273][2] ,
         \CARRYB[273][1] , \CARRYB[273][0] , \CARRYB[272][2] ,
         \CARRYB[272][1] , \CARRYB[272][0] , \CARRYB[271][2] ,
         \CARRYB[271][1] , \CARRYB[271][0] , \CARRYB[270][2] ,
         \CARRYB[270][1] , \CARRYB[270][0] , \CARRYB[269][2] ,
         \CARRYB[269][1] , \CARRYB[269][0] , \CARRYB[268][2] ,
         \CARRYB[268][1] , \CARRYB[268][0] , \CARRYB[267][2] ,
         \CARRYB[267][1] , \CARRYB[267][0] , \CARRYB[266][2] ,
         \CARRYB[266][1] , \CARRYB[266][0] , \CARRYB[265][2] ,
         \CARRYB[265][1] , \CARRYB[265][0] , \CARRYB[264][2] ,
         \CARRYB[264][1] , \CARRYB[264][0] , \CARRYB[263][2] ,
         \CARRYB[263][1] , \CARRYB[263][0] , \CARRYB[262][2] ,
         \CARRYB[262][1] , \CARRYB[262][0] , \CARRYB[261][2] ,
         \CARRYB[261][1] , \CARRYB[261][0] , \CARRYB[260][2] ,
         \CARRYB[260][1] , \CARRYB[260][0] , \CARRYB[259][2] ,
         \CARRYB[259][1] , \CARRYB[259][0] , \CARRYB[258][2] ,
         \CARRYB[258][1] , \CARRYB[258][0] , \CARRYB[257][2] ,
         \CARRYB[257][1] , \CARRYB[257][0] , \CARRYB[256][2] ,
         \CARRYB[256][1] , \CARRYB[256][0] , \SUMB[383][2] , \SUMB[383][1] ,
         \SUMB[382][2] , \SUMB[382][1] , \SUMB[381][2] , \SUMB[381][1] ,
         \SUMB[380][2] , \SUMB[380][1] , \SUMB[379][2] , \SUMB[379][1] ,
         \SUMB[378][2] , \SUMB[378][1] , \SUMB[377][2] , \SUMB[377][1] ,
         \SUMB[376][2] , \SUMB[376][1] , \SUMB[375][2] , \SUMB[375][1] ,
         \SUMB[374][2] , \SUMB[374][1] , \SUMB[373][2] , \SUMB[373][1] ,
         \SUMB[372][2] , \SUMB[372][1] , \SUMB[371][2] , \SUMB[371][1] ,
         \SUMB[370][2] , \SUMB[370][1] , \SUMB[369][2] , \SUMB[369][1] ,
         \SUMB[368][2] , \SUMB[368][1] , \SUMB[367][2] , \SUMB[367][1] ,
         \SUMB[366][2] , \SUMB[366][1] , \SUMB[365][2] , \SUMB[365][1] ,
         \SUMB[364][2] , \SUMB[364][1] , \SUMB[363][2] , \SUMB[363][1] ,
         \SUMB[362][2] , \SUMB[362][1] , \SUMB[361][2] , \SUMB[361][1] ,
         \SUMB[360][2] , \SUMB[360][1] , \SUMB[359][2] , \SUMB[359][1] ,
         \SUMB[358][2] , \SUMB[358][1] , \SUMB[357][2] , \SUMB[357][1] ,
         \SUMB[356][2] , \SUMB[356][1] , \SUMB[355][2] , \SUMB[355][1] ,
         \SUMB[354][2] , \SUMB[354][1] , \SUMB[353][2] , \SUMB[353][1] ,
         \SUMB[352][2] , \SUMB[352][1] , \SUMB[351][2] , \SUMB[351][1] ,
         \SUMB[350][2] , \SUMB[350][1] , \SUMB[349][2] , \SUMB[349][1] ,
         \SUMB[348][2] , \SUMB[348][1] , \SUMB[347][2] , \SUMB[347][1] ,
         \SUMB[346][2] , \SUMB[346][1] , \SUMB[345][2] , \SUMB[345][1] ,
         \SUMB[344][2] , \SUMB[344][1] , \SUMB[343][2] , \SUMB[343][1] ,
         \SUMB[342][2] , \SUMB[342][1] , \SUMB[341][2] , \SUMB[341][1] ,
         \SUMB[340][2] , \SUMB[340][1] , \SUMB[339][2] , \SUMB[339][1] ,
         \SUMB[338][2] , \SUMB[338][1] , \SUMB[337][2] , \SUMB[337][1] ,
         \SUMB[336][2] , \SUMB[336][1] , \SUMB[335][2] , \SUMB[335][1] ,
         \SUMB[334][2] , \SUMB[334][1] , \SUMB[333][2] , \SUMB[333][1] ,
         \SUMB[332][2] , \SUMB[332][1] , \SUMB[331][2] , \SUMB[331][1] ,
         \SUMB[330][2] , \SUMB[330][1] , \SUMB[329][2] , \SUMB[329][1] ,
         \SUMB[328][2] , \SUMB[328][1] , \SUMB[327][2] , \SUMB[327][1] ,
         \SUMB[326][2] , \SUMB[326][1] , \SUMB[325][2] , \SUMB[325][1] ,
         \SUMB[324][2] , \SUMB[324][1] , \SUMB[323][2] , \SUMB[323][1] ,
         \SUMB[322][2] , \SUMB[322][1] , \SUMB[321][2] , \SUMB[321][1] ,
         \SUMB[320][2] , \SUMB[320][1] , \SUMB[319][2] , \SUMB[319][1] ,
         \SUMB[318][2] , \SUMB[318][1] , \SUMB[317][2] , \SUMB[317][1] ,
         \SUMB[316][2] , \SUMB[316][1] , \SUMB[315][2] , \SUMB[315][1] ,
         \SUMB[314][2] , \SUMB[314][1] , \SUMB[313][2] , \SUMB[313][1] ,
         \SUMB[312][2] , \SUMB[312][1] , \SUMB[311][2] , \SUMB[311][1] ,
         \SUMB[310][2] , \SUMB[310][1] , \SUMB[309][2] , \SUMB[309][1] ,
         \SUMB[308][2] , \SUMB[308][1] , \SUMB[307][2] , \SUMB[307][1] ,
         \SUMB[306][2] , \SUMB[306][1] , \SUMB[305][2] , \SUMB[305][1] ,
         \SUMB[304][2] , \SUMB[304][1] , \SUMB[303][2] , \SUMB[303][1] ,
         \SUMB[302][2] , \SUMB[302][1] , \SUMB[301][2] , \SUMB[301][1] ,
         \SUMB[300][2] , \SUMB[300][1] , \SUMB[299][2] , \SUMB[299][1] ,
         \SUMB[298][2] , \SUMB[298][1] , \SUMB[297][2] , \SUMB[297][1] ,
         \SUMB[296][2] , \SUMB[296][1] , \SUMB[295][2] , \SUMB[295][1] ,
         \SUMB[294][2] , \SUMB[294][1] , \SUMB[293][2] , \SUMB[293][1] ,
         \SUMB[292][2] , \SUMB[292][1] , \SUMB[291][2] , \SUMB[291][1] ,
         \SUMB[290][2] , \SUMB[290][1] , \SUMB[289][2] , \SUMB[289][1] ,
         \SUMB[288][2] , \SUMB[288][1] , \SUMB[287][2] , \SUMB[287][1] ,
         \SUMB[286][2] , \SUMB[286][1] , \SUMB[285][2] , \SUMB[285][1] ,
         \SUMB[284][2] , \SUMB[284][1] , \SUMB[283][2] , \SUMB[283][1] ,
         \SUMB[282][2] , \SUMB[282][1] , \SUMB[281][2] , \SUMB[281][1] ,
         \SUMB[280][2] , \SUMB[280][1] , \SUMB[279][2] , \SUMB[279][1] ,
         \SUMB[278][2] , \SUMB[278][1] , \SUMB[277][2] , \SUMB[277][1] ,
         \SUMB[276][2] , \SUMB[276][1] , \SUMB[275][2] , \SUMB[275][1] ,
         \SUMB[274][2] , \SUMB[274][1] , \SUMB[273][2] , \SUMB[273][1] ,
         \SUMB[272][2] , \SUMB[272][1] , \SUMB[271][2] , \SUMB[271][1] ,
         \SUMB[270][2] , \SUMB[270][1] , \SUMB[269][2] , \SUMB[269][1] ,
         \SUMB[268][2] , \SUMB[268][1] , \SUMB[267][2] , \SUMB[267][1] ,
         \SUMB[266][2] , \SUMB[266][1] , \SUMB[265][2] , \SUMB[265][1] ,
         \SUMB[264][2] , \SUMB[264][1] , \SUMB[263][2] , \SUMB[263][1] ,
         \SUMB[262][2] , \SUMB[262][1] , \SUMB[261][2] , \SUMB[261][1] ,
         \SUMB[260][2] , \SUMB[260][1] , \SUMB[259][2] , \SUMB[259][1] ,
         \SUMB[258][2] , \SUMB[258][1] , \SUMB[257][2] , \SUMB[257][1] ,
         \SUMB[256][2] , \SUMB[256][1] , \CARRYB[511][2] , \CARRYB[511][1] ,
         \CARRYB[511][0] , \CARRYB[510][2] , \CARRYB[510][1] ,
         \CARRYB[510][0] , \CARRYB[509][2] , \CARRYB[509][1] ,
         \CARRYB[509][0] , \CARRYB[508][2] , \CARRYB[508][1] ,
         \CARRYB[508][0] , \CARRYB[507][2] , \CARRYB[507][1] ,
         \CARRYB[507][0] , \CARRYB[506][2] , \CARRYB[506][1] ,
         \CARRYB[506][0] , \CARRYB[505][2] , \CARRYB[505][1] ,
         \CARRYB[505][0] , \CARRYB[504][2] , \CARRYB[504][1] ,
         \CARRYB[504][0] , \CARRYB[503][2] , \CARRYB[503][1] ,
         \CARRYB[503][0] , \CARRYB[502][2] , \CARRYB[502][1] ,
         \CARRYB[502][0] , \CARRYB[501][2] , \CARRYB[501][1] ,
         \CARRYB[501][0] , \CARRYB[500][2] , \CARRYB[500][1] ,
         \CARRYB[500][0] , \CARRYB[499][2] , \CARRYB[499][1] ,
         \CARRYB[499][0] , \CARRYB[498][2] , \CARRYB[498][1] ,
         \CARRYB[498][0] , \CARRYB[497][2] , \CARRYB[497][1] ,
         \CARRYB[497][0] , \CARRYB[496][2] , \CARRYB[496][1] ,
         \CARRYB[496][0] , \CARRYB[495][2] , \CARRYB[495][1] ,
         \CARRYB[495][0] , \CARRYB[494][2] , \CARRYB[494][1] ,
         \CARRYB[494][0] , \CARRYB[493][2] , \CARRYB[493][1] ,
         \CARRYB[493][0] , \CARRYB[492][2] , \CARRYB[492][1] ,
         \CARRYB[492][0] , \CARRYB[491][2] , \CARRYB[491][1] ,
         \CARRYB[491][0] , \CARRYB[490][2] , \CARRYB[490][1] ,
         \CARRYB[490][0] , \CARRYB[489][2] , \CARRYB[489][1] ,
         \CARRYB[489][0] , \CARRYB[488][2] , \CARRYB[488][1] ,
         \CARRYB[488][0] , \CARRYB[487][2] , \CARRYB[487][1] ,
         \CARRYB[487][0] , \CARRYB[486][2] , \CARRYB[486][1] ,
         \CARRYB[486][0] , \CARRYB[485][2] , \CARRYB[485][1] ,
         \CARRYB[485][0] , \CARRYB[484][2] , \CARRYB[484][1] ,
         \CARRYB[484][0] , \CARRYB[483][2] , \CARRYB[483][1] ,
         \CARRYB[483][0] , \CARRYB[482][2] , \CARRYB[482][1] ,
         \CARRYB[482][0] , \CARRYB[481][2] , \CARRYB[481][1] ,
         \CARRYB[481][0] , \CARRYB[480][2] , \CARRYB[480][1] ,
         \CARRYB[480][0] , \CARRYB[479][2] , \CARRYB[479][1] ,
         \CARRYB[479][0] , \CARRYB[478][2] , \CARRYB[478][1] ,
         \CARRYB[478][0] , \CARRYB[477][2] , \CARRYB[477][1] ,
         \CARRYB[477][0] , \CARRYB[476][2] , \CARRYB[476][1] ,
         \CARRYB[476][0] , \CARRYB[475][2] , \CARRYB[475][1] ,
         \CARRYB[475][0] , \CARRYB[474][2] , \CARRYB[474][1] ,
         \CARRYB[474][0] , \CARRYB[473][2] , \CARRYB[473][1] ,
         \CARRYB[473][0] , \CARRYB[472][2] , \CARRYB[472][1] ,
         \CARRYB[472][0] , \CARRYB[471][2] , \CARRYB[471][1] ,
         \CARRYB[471][0] , \CARRYB[470][2] , \CARRYB[470][1] ,
         \CARRYB[470][0] , \CARRYB[469][2] , \CARRYB[469][1] ,
         \CARRYB[469][0] , \CARRYB[468][2] , \CARRYB[468][1] ,
         \CARRYB[468][0] , \CARRYB[467][2] , \CARRYB[467][1] ,
         \CARRYB[467][0] , \CARRYB[466][2] , \CARRYB[466][1] ,
         \CARRYB[466][0] , \CARRYB[465][2] , \CARRYB[465][1] ,
         \CARRYB[465][0] , \CARRYB[464][2] , \CARRYB[464][1] ,
         \CARRYB[464][0] , \CARRYB[463][2] , \CARRYB[463][1] ,
         \CARRYB[463][0] , \CARRYB[462][2] , \CARRYB[462][1] ,
         \CARRYB[462][0] , \CARRYB[461][2] , \CARRYB[461][1] ,
         \CARRYB[461][0] , \CARRYB[460][2] , \CARRYB[460][1] ,
         \CARRYB[460][0] , \CARRYB[459][2] , \CARRYB[459][1] ,
         \CARRYB[459][0] , \CARRYB[458][2] , \CARRYB[458][1] ,
         \CARRYB[458][0] , \CARRYB[457][2] , \CARRYB[457][1] ,
         \CARRYB[457][0] , \CARRYB[456][2] , \CARRYB[456][1] ,
         \CARRYB[456][0] , \CARRYB[455][2] , \CARRYB[455][1] ,
         \CARRYB[455][0] , \CARRYB[454][2] , \CARRYB[454][1] ,
         \CARRYB[454][0] , \CARRYB[453][2] , \CARRYB[453][1] ,
         \CARRYB[453][0] , \CARRYB[452][2] , \CARRYB[452][1] ,
         \CARRYB[452][0] , \CARRYB[451][2] , \CARRYB[451][1] ,
         \CARRYB[451][0] , \CARRYB[450][2] , \CARRYB[450][1] ,
         \CARRYB[450][0] , \CARRYB[449][2] , \CARRYB[449][1] ,
         \CARRYB[449][0] , \CARRYB[448][2] , \CARRYB[448][1] ,
         \CARRYB[448][0] , \CARRYB[447][2] , \CARRYB[447][1] ,
         \CARRYB[447][0] , \CARRYB[446][2] , \CARRYB[446][1] ,
         \CARRYB[446][0] , \CARRYB[445][2] , \CARRYB[445][1] ,
         \CARRYB[445][0] , \CARRYB[444][2] , \CARRYB[444][1] ,
         \CARRYB[444][0] , \CARRYB[443][2] , \CARRYB[443][1] ,
         \CARRYB[443][0] , \CARRYB[442][2] , \CARRYB[442][1] ,
         \CARRYB[442][0] , \CARRYB[441][2] , \CARRYB[441][1] ,
         \CARRYB[441][0] , \CARRYB[440][2] , \CARRYB[440][1] ,
         \CARRYB[440][0] , \CARRYB[439][2] , \CARRYB[439][1] ,
         \CARRYB[439][0] , \CARRYB[438][2] , \CARRYB[438][1] ,
         \CARRYB[438][0] , \CARRYB[437][2] , \CARRYB[437][1] ,
         \CARRYB[437][0] , \CARRYB[436][2] , \CARRYB[436][1] ,
         \CARRYB[436][0] , \CARRYB[435][2] , \CARRYB[435][1] ,
         \CARRYB[435][0] , \CARRYB[434][2] , \CARRYB[434][1] ,
         \CARRYB[434][0] , \CARRYB[433][2] , \CARRYB[433][1] ,
         \CARRYB[433][0] , \CARRYB[432][2] , \CARRYB[432][1] ,
         \CARRYB[432][0] , \CARRYB[431][2] , \CARRYB[431][1] ,
         \CARRYB[431][0] , \CARRYB[430][2] , \CARRYB[430][1] ,
         \CARRYB[430][0] , \CARRYB[429][2] , \CARRYB[429][1] ,
         \CARRYB[429][0] , \CARRYB[428][2] , \CARRYB[428][1] ,
         \CARRYB[428][0] , \CARRYB[427][2] , \CARRYB[427][1] ,
         \CARRYB[427][0] , \CARRYB[426][2] , \CARRYB[426][1] ,
         \CARRYB[426][0] , \CARRYB[425][2] , \CARRYB[425][1] ,
         \CARRYB[425][0] , \CARRYB[424][2] , \CARRYB[424][1] ,
         \CARRYB[424][0] , \CARRYB[423][2] , \CARRYB[423][1] ,
         \CARRYB[423][0] , \CARRYB[422][2] , \CARRYB[422][1] ,
         \CARRYB[422][0] , \CARRYB[421][2] , \CARRYB[421][1] ,
         \CARRYB[421][0] , \CARRYB[420][2] , \CARRYB[420][1] ,
         \CARRYB[420][0] , \CARRYB[419][2] , \CARRYB[419][1] ,
         \CARRYB[419][0] , \CARRYB[418][2] , \CARRYB[418][1] ,
         \CARRYB[418][0] , \CARRYB[417][2] , \CARRYB[417][1] ,
         \CARRYB[417][0] , \CARRYB[416][2] , \CARRYB[416][1] ,
         \CARRYB[416][0] , \CARRYB[415][2] , \CARRYB[415][1] ,
         \CARRYB[415][0] , \CARRYB[414][2] , \CARRYB[414][1] ,
         \CARRYB[414][0] , \CARRYB[413][2] , \CARRYB[413][1] ,
         \CARRYB[413][0] , \CARRYB[412][2] , \CARRYB[412][1] ,
         \CARRYB[412][0] , \CARRYB[411][2] , \CARRYB[411][1] ,
         \CARRYB[411][0] , \CARRYB[410][2] , \CARRYB[410][1] ,
         \CARRYB[410][0] , \CARRYB[409][2] , \CARRYB[409][1] ,
         \CARRYB[409][0] , \CARRYB[408][2] , \CARRYB[408][1] ,
         \CARRYB[408][0] , \CARRYB[407][2] , \CARRYB[407][1] ,
         \CARRYB[407][0] , \CARRYB[406][2] , \CARRYB[406][1] ,
         \CARRYB[406][0] , \CARRYB[405][2] , \CARRYB[405][1] ,
         \CARRYB[405][0] , \CARRYB[404][2] , \CARRYB[404][1] ,
         \CARRYB[404][0] , \CARRYB[403][2] , \CARRYB[403][1] ,
         \CARRYB[403][0] , \CARRYB[402][2] , \CARRYB[402][1] ,
         \CARRYB[402][0] , \CARRYB[401][2] , \CARRYB[401][1] ,
         \CARRYB[401][0] , \CARRYB[400][2] , \CARRYB[400][1] ,
         \CARRYB[400][0] , \CARRYB[399][2] , \CARRYB[399][1] ,
         \CARRYB[399][0] , \CARRYB[398][2] , \CARRYB[398][1] ,
         \CARRYB[398][0] , \CARRYB[397][2] , \CARRYB[397][1] ,
         \CARRYB[397][0] , \CARRYB[396][2] , \CARRYB[396][1] ,
         \CARRYB[396][0] , \CARRYB[395][2] , \CARRYB[395][1] ,
         \CARRYB[395][0] , \CARRYB[394][2] , \CARRYB[394][1] ,
         \CARRYB[394][0] , \CARRYB[393][2] , \CARRYB[393][1] ,
         \CARRYB[393][0] , \CARRYB[392][2] , \CARRYB[392][1] ,
         \CARRYB[392][0] , \CARRYB[391][2] , \CARRYB[391][1] ,
         \CARRYB[391][0] , \CARRYB[390][2] , \CARRYB[390][1] ,
         \CARRYB[390][0] , \CARRYB[389][2] , \CARRYB[389][1] ,
         \CARRYB[389][0] , \CARRYB[388][2] , \CARRYB[388][1] ,
         \CARRYB[388][0] , \CARRYB[387][2] , \CARRYB[387][1] ,
         \CARRYB[387][0] , \CARRYB[386][2] , \CARRYB[386][1] ,
         \CARRYB[386][0] , \CARRYB[385][2] , \CARRYB[385][1] ,
         \CARRYB[385][0] , \CARRYB[384][2] , \CARRYB[384][1] ,
         \CARRYB[384][0] , \SUMB[511][2] , \SUMB[511][1] , \SUMB[510][2] ,
         \SUMB[510][1] , \SUMB[509][2] , \SUMB[509][1] , \SUMB[508][2] ,
         \SUMB[508][1] , \SUMB[507][2] , \SUMB[507][1] , \SUMB[506][2] ,
         \SUMB[506][1] , \SUMB[505][2] , \SUMB[505][1] , \SUMB[504][2] ,
         \SUMB[504][1] , \SUMB[503][2] , \SUMB[503][1] , \SUMB[502][2] ,
         \SUMB[502][1] , \SUMB[501][2] , \SUMB[501][1] , \SUMB[500][2] ,
         \SUMB[500][1] , \SUMB[499][2] , \SUMB[499][1] , \SUMB[498][2] ,
         \SUMB[498][1] , \SUMB[497][2] , \SUMB[497][1] , \SUMB[496][2] ,
         \SUMB[496][1] , \SUMB[495][2] , \SUMB[495][1] , \SUMB[494][2] ,
         \SUMB[494][1] , \SUMB[493][2] , \SUMB[493][1] , \SUMB[492][2] ,
         \SUMB[492][1] , \SUMB[491][2] , \SUMB[491][1] , \SUMB[490][2] ,
         \SUMB[490][1] , \SUMB[489][2] , \SUMB[489][1] , \SUMB[488][2] ,
         \SUMB[488][1] , \SUMB[487][2] , \SUMB[487][1] , \SUMB[486][2] ,
         \SUMB[486][1] , \SUMB[485][2] , \SUMB[485][1] , \SUMB[484][2] ,
         \SUMB[484][1] , \SUMB[483][2] , \SUMB[483][1] , \SUMB[482][2] ,
         \SUMB[482][1] , \SUMB[481][2] , \SUMB[481][1] , \SUMB[480][2] ,
         \SUMB[480][1] , \SUMB[479][2] , \SUMB[479][1] , \SUMB[478][2] ,
         \SUMB[478][1] , \SUMB[477][2] , \SUMB[477][1] , \SUMB[476][2] ,
         \SUMB[476][1] , \SUMB[475][2] , \SUMB[475][1] , \SUMB[474][2] ,
         \SUMB[474][1] , \SUMB[473][2] , \SUMB[473][1] , \SUMB[472][2] ,
         \SUMB[472][1] , \SUMB[471][2] , \SUMB[471][1] , \SUMB[470][2] ,
         \SUMB[470][1] , \SUMB[469][2] , \SUMB[469][1] , \SUMB[468][2] ,
         \SUMB[468][1] , \SUMB[467][2] , \SUMB[467][1] , \SUMB[466][2] ,
         \SUMB[466][1] , \SUMB[465][2] , \SUMB[465][1] , \SUMB[464][2] ,
         \SUMB[464][1] , \SUMB[463][2] , \SUMB[463][1] , \SUMB[462][2] ,
         \SUMB[462][1] , \SUMB[461][2] , \SUMB[461][1] , \SUMB[460][2] ,
         \SUMB[460][1] , \SUMB[459][2] , \SUMB[459][1] , \SUMB[458][2] ,
         \SUMB[458][1] , \SUMB[457][2] , \SUMB[457][1] , \SUMB[456][2] ,
         \SUMB[456][1] , \SUMB[455][2] , \SUMB[455][1] , \SUMB[454][2] ,
         \SUMB[454][1] , \SUMB[453][2] , \SUMB[453][1] , \SUMB[452][2] ,
         \SUMB[452][1] , \SUMB[451][2] , \SUMB[451][1] , \SUMB[450][2] ,
         \SUMB[450][1] , \SUMB[449][2] , \SUMB[449][1] , \SUMB[448][2] ,
         \SUMB[448][1] , \SUMB[447][2] , \SUMB[447][1] , \SUMB[446][2] ,
         \SUMB[446][1] , \SUMB[445][2] , \SUMB[445][1] , \SUMB[444][2] ,
         \SUMB[444][1] , \SUMB[443][2] , \SUMB[443][1] , \SUMB[442][2] ,
         \SUMB[442][1] , \SUMB[441][2] , \SUMB[441][1] , \SUMB[440][2] ,
         \SUMB[440][1] , \SUMB[439][2] , \SUMB[439][1] , \SUMB[438][2] ,
         \SUMB[438][1] , \SUMB[437][2] , \SUMB[437][1] , \SUMB[436][2] ,
         \SUMB[436][1] , \SUMB[435][2] , \SUMB[435][1] , \SUMB[434][2] ,
         \SUMB[434][1] , \SUMB[433][2] , \SUMB[433][1] , \SUMB[432][2] ,
         \SUMB[432][1] , \SUMB[431][2] , \SUMB[431][1] , \SUMB[430][2] ,
         \SUMB[430][1] , \SUMB[429][2] , \SUMB[429][1] , \SUMB[428][2] ,
         \SUMB[428][1] , \SUMB[427][2] , \SUMB[427][1] , \SUMB[426][2] ,
         \SUMB[426][1] , \SUMB[425][2] , \SUMB[425][1] , \SUMB[424][2] ,
         \SUMB[424][1] , \SUMB[423][2] , \SUMB[423][1] , \SUMB[422][2] ,
         \SUMB[422][1] , \SUMB[421][2] , \SUMB[421][1] , \SUMB[420][2] ,
         \SUMB[420][1] , \SUMB[419][2] , \SUMB[419][1] , \SUMB[418][2] ,
         \SUMB[418][1] , \SUMB[417][2] , \SUMB[417][1] , \SUMB[416][2] ,
         \SUMB[416][1] , \SUMB[415][2] , \SUMB[415][1] , \SUMB[414][2] ,
         \SUMB[414][1] , \SUMB[413][2] , \SUMB[413][1] , \SUMB[412][2] ,
         \SUMB[412][1] , \SUMB[411][2] , \SUMB[411][1] , \SUMB[410][2] ,
         \SUMB[410][1] , \SUMB[409][2] , \SUMB[409][1] , \SUMB[408][2] ,
         \SUMB[408][1] , \SUMB[407][2] , \SUMB[407][1] , \SUMB[406][2] ,
         \SUMB[406][1] , \SUMB[405][2] , \SUMB[405][1] , \SUMB[404][2] ,
         \SUMB[404][1] , \SUMB[403][2] , \SUMB[403][1] , \SUMB[402][2] ,
         \SUMB[402][1] , \SUMB[401][2] , \SUMB[401][1] , \SUMB[400][2] ,
         \SUMB[400][1] , \SUMB[399][2] , \SUMB[399][1] , \SUMB[398][2] ,
         \SUMB[398][1] , \SUMB[397][2] , \SUMB[397][1] , \SUMB[396][2] ,
         \SUMB[396][1] , \SUMB[395][2] , \SUMB[395][1] , \SUMB[394][2] ,
         \SUMB[394][1] , \SUMB[393][2] , \SUMB[393][1] , \SUMB[392][2] ,
         \SUMB[392][1] , \SUMB[391][2] , \SUMB[391][1] , \SUMB[390][2] ,
         \SUMB[390][1] , \SUMB[389][2] , \SUMB[389][1] , \SUMB[388][2] ,
         \SUMB[388][1] , \SUMB[387][2] , \SUMB[387][1] , \SUMB[386][2] ,
         \SUMB[386][1] , \SUMB[385][2] , \SUMB[385][1] , \SUMB[384][2] ,
         \SUMB[384][1] , \CARRYB[639][2] , \CARRYB[639][1] , \CARRYB[639][0] ,
         \CARRYB[638][2] , \CARRYB[638][1] , \CARRYB[638][0] ,
         \CARRYB[637][2] , \CARRYB[637][1] , \CARRYB[637][0] ,
         \CARRYB[636][2] , \CARRYB[636][1] , \CARRYB[636][0] ,
         \CARRYB[635][2] , \CARRYB[635][1] , \CARRYB[635][0] ,
         \CARRYB[634][2] , \CARRYB[634][1] , \CARRYB[634][0] ,
         \CARRYB[633][2] , \CARRYB[633][1] , \CARRYB[633][0] ,
         \CARRYB[632][2] , \CARRYB[632][1] , \CARRYB[632][0] ,
         \CARRYB[631][2] , \CARRYB[631][1] , \CARRYB[631][0] ,
         \CARRYB[630][2] , \CARRYB[630][1] , \CARRYB[630][0] ,
         \CARRYB[629][2] , \CARRYB[629][1] , \CARRYB[629][0] ,
         \CARRYB[628][2] , \CARRYB[628][1] , \CARRYB[628][0] ,
         \CARRYB[627][2] , \CARRYB[627][1] , \CARRYB[627][0] ,
         \CARRYB[626][2] , \CARRYB[626][1] , \CARRYB[626][0] ,
         \CARRYB[625][2] , \CARRYB[625][1] , \CARRYB[625][0] ,
         \CARRYB[624][2] , \CARRYB[624][1] , \CARRYB[624][0] ,
         \CARRYB[623][2] , \CARRYB[623][1] , \CARRYB[623][0] ,
         \CARRYB[622][2] , \CARRYB[622][1] , \CARRYB[622][0] ,
         \CARRYB[621][2] , \CARRYB[621][1] , \CARRYB[621][0] ,
         \CARRYB[620][2] , \CARRYB[620][1] , \CARRYB[620][0] ,
         \CARRYB[619][2] , \CARRYB[619][1] , \CARRYB[619][0] ,
         \CARRYB[618][2] , \CARRYB[618][1] , \CARRYB[618][0] ,
         \CARRYB[617][2] , \CARRYB[617][1] , \CARRYB[617][0] ,
         \CARRYB[616][2] , \CARRYB[616][1] , \CARRYB[616][0] ,
         \CARRYB[615][2] , \CARRYB[615][1] , \CARRYB[615][0] ,
         \CARRYB[614][2] , \CARRYB[614][1] , \CARRYB[614][0] ,
         \CARRYB[613][2] , \CARRYB[613][1] , \CARRYB[613][0] ,
         \CARRYB[612][2] , \CARRYB[612][1] , \CARRYB[612][0] ,
         \CARRYB[611][2] , \CARRYB[611][1] , \CARRYB[611][0] ,
         \CARRYB[610][2] , \CARRYB[610][1] , \CARRYB[610][0] ,
         \CARRYB[609][2] , \CARRYB[609][1] , \CARRYB[609][0] ,
         \CARRYB[608][2] , \CARRYB[608][1] , \CARRYB[608][0] ,
         \CARRYB[607][2] , \CARRYB[607][1] , \CARRYB[607][0] ,
         \CARRYB[606][2] , \CARRYB[606][1] , \CARRYB[606][0] ,
         \CARRYB[605][2] , \CARRYB[605][1] , \CARRYB[605][0] ,
         \CARRYB[604][2] , \CARRYB[604][1] , \CARRYB[604][0] ,
         \CARRYB[603][2] , \CARRYB[603][1] , \CARRYB[603][0] ,
         \CARRYB[602][2] , \CARRYB[602][1] , \CARRYB[602][0] ,
         \CARRYB[601][2] , \CARRYB[601][1] , \CARRYB[601][0] ,
         \CARRYB[600][2] , \CARRYB[600][1] , \CARRYB[600][0] ,
         \CARRYB[599][2] , \CARRYB[599][1] , \CARRYB[599][0] ,
         \CARRYB[598][2] , \CARRYB[598][1] , \CARRYB[598][0] ,
         \CARRYB[597][2] , \CARRYB[597][1] , \CARRYB[597][0] ,
         \CARRYB[596][2] , \CARRYB[596][1] , \CARRYB[596][0] ,
         \CARRYB[595][2] , \CARRYB[595][1] , \CARRYB[595][0] ,
         \CARRYB[594][2] , \CARRYB[594][1] , \CARRYB[594][0] ,
         \CARRYB[593][2] , \CARRYB[593][1] , \CARRYB[593][0] ,
         \CARRYB[592][2] , \CARRYB[592][1] , \CARRYB[592][0] ,
         \CARRYB[591][2] , \CARRYB[591][1] , \CARRYB[591][0] ,
         \CARRYB[590][2] , \CARRYB[590][1] , \CARRYB[590][0] ,
         \CARRYB[589][2] , \CARRYB[589][1] , \CARRYB[589][0] ,
         \CARRYB[588][2] , \CARRYB[588][1] , \CARRYB[588][0] ,
         \CARRYB[587][2] , \CARRYB[587][1] , \CARRYB[587][0] ,
         \CARRYB[586][2] , \CARRYB[586][1] , \CARRYB[586][0] ,
         \CARRYB[585][2] , \CARRYB[585][1] , \CARRYB[585][0] ,
         \CARRYB[584][2] , \CARRYB[584][1] , \CARRYB[584][0] ,
         \CARRYB[583][2] , \CARRYB[583][1] , \CARRYB[583][0] ,
         \CARRYB[582][2] , \CARRYB[582][1] , \CARRYB[582][0] ,
         \CARRYB[581][2] , \CARRYB[581][1] , \CARRYB[581][0] ,
         \CARRYB[580][2] , \CARRYB[580][1] , \CARRYB[580][0] ,
         \CARRYB[579][2] , \CARRYB[579][1] , \CARRYB[579][0] ,
         \CARRYB[578][2] , \CARRYB[578][1] , \CARRYB[578][0] ,
         \CARRYB[577][2] , \CARRYB[577][1] , \CARRYB[577][0] ,
         \CARRYB[576][2] , \CARRYB[576][1] , \CARRYB[576][0] ,
         \CARRYB[575][2] , \CARRYB[575][1] , \CARRYB[575][0] ,
         \CARRYB[574][2] , \CARRYB[574][1] , \CARRYB[574][0] ,
         \CARRYB[573][2] , \CARRYB[573][1] , \CARRYB[573][0] ,
         \CARRYB[572][2] , \CARRYB[572][1] , \CARRYB[572][0] ,
         \CARRYB[571][2] , \CARRYB[571][1] , \CARRYB[571][0] ,
         \CARRYB[570][2] , \CARRYB[570][1] , \CARRYB[570][0] ,
         \CARRYB[569][2] , \CARRYB[569][1] , \CARRYB[569][0] ,
         \CARRYB[568][2] , \CARRYB[568][1] , \CARRYB[568][0] ,
         \CARRYB[567][2] , \CARRYB[567][1] , \CARRYB[567][0] ,
         \CARRYB[566][2] , \CARRYB[566][1] , \CARRYB[566][0] ,
         \CARRYB[565][2] , \CARRYB[565][1] , \CARRYB[565][0] ,
         \CARRYB[564][2] , \CARRYB[564][1] , \CARRYB[564][0] ,
         \CARRYB[563][2] , \CARRYB[563][1] , \CARRYB[563][0] ,
         \CARRYB[562][2] , \CARRYB[562][1] , \CARRYB[562][0] ,
         \CARRYB[561][2] , \CARRYB[561][1] , \CARRYB[561][0] ,
         \CARRYB[560][2] , \CARRYB[560][1] , \CARRYB[560][0] ,
         \CARRYB[559][2] , \CARRYB[559][1] , \CARRYB[559][0] ,
         \CARRYB[558][2] , \CARRYB[558][1] , \CARRYB[558][0] ,
         \CARRYB[557][2] , \CARRYB[557][1] , \CARRYB[557][0] ,
         \CARRYB[556][2] , \CARRYB[556][1] , \CARRYB[556][0] ,
         \CARRYB[555][2] , \CARRYB[555][1] , \CARRYB[555][0] ,
         \CARRYB[554][2] , \CARRYB[554][1] , \CARRYB[554][0] ,
         \CARRYB[553][2] , \CARRYB[553][1] , \CARRYB[553][0] ,
         \CARRYB[552][2] , \CARRYB[552][1] , \CARRYB[552][0] ,
         \CARRYB[551][2] , \CARRYB[551][1] , \CARRYB[551][0] ,
         \CARRYB[550][2] , \CARRYB[550][1] , \CARRYB[550][0] ,
         \CARRYB[549][2] , \CARRYB[549][1] , \CARRYB[549][0] ,
         \CARRYB[548][2] , \CARRYB[548][1] , \CARRYB[548][0] ,
         \CARRYB[547][2] , \CARRYB[547][1] , \CARRYB[547][0] ,
         \CARRYB[546][2] , \CARRYB[546][1] , \CARRYB[546][0] ,
         \CARRYB[545][2] , \CARRYB[545][1] , \CARRYB[545][0] ,
         \CARRYB[544][2] , \CARRYB[544][1] , \CARRYB[544][0] ,
         \CARRYB[543][2] , \CARRYB[543][1] , \CARRYB[543][0] ,
         \CARRYB[542][2] , \CARRYB[542][1] , \CARRYB[542][0] ,
         \CARRYB[541][2] , \CARRYB[541][1] , \CARRYB[541][0] ,
         \CARRYB[540][2] , \CARRYB[540][1] , \CARRYB[540][0] ,
         \CARRYB[539][2] , \CARRYB[539][1] , \CARRYB[539][0] ,
         \CARRYB[538][2] , \CARRYB[538][1] , \CARRYB[538][0] ,
         \CARRYB[537][2] , \CARRYB[537][1] , \CARRYB[537][0] ,
         \CARRYB[536][2] , \CARRYB[536][1] , \CARRYB[536][0] ,
         \CARRYB[535][2] , \CARRYB[535][1] , \CARRYB[535][0] ,
         \CARRYB[534][2] , \CARRYB[534][1] , \CARRYB[534][0] ,
         \CARRYB[533][2] , \CARRYB[533][1] , \CARRYB[533][0] ,
         \CARRYB[532][2] , \CARRYB[532][1] , \CARRYB[532][0] ,
         \CARRYB[531][2] , \CARRYB[531][1] , \CARRYB[531][0] ,
         \CARRYB[530][2] , \CARRYB[530][1] , \CARRYB[530][0] ,
         \CARRYB[529][2] , \CARRYB[529][1] , \CARRYB[529][0] ,
         \CARRYB[528][2] , \CARRYB[528][1] , \CARRYB[528][0] ,
         \CARRYB[527][2] , \CARRYB[527][1] , \CARRYB[527][0] ,
         \CARRYB[526][2] , \CARRYB[526][1] , \CARRYB[526][0] ,
         \CARRYB[525][2] , \CARRYB[525][1] , \CARRYB[525][0] ,
         \CARRYB[524][2] , \CARRYB[524][1] , \CARRYB[524][0] ,
         \CARRYB[523][2] , \CARRYB[523][1] , \CARRYB[523][0] ,
         \CARRYB[522][2] , \CARRYB[522][1] , \CARRYB[522][0] ,
         \CARRYB[521][2] , \CARRYB[521][1] , \CARRYB[521][0] ,
         \CARRYB[520][2] , \CARRYB[520][1] , \CARRYB[520][0] ,
         \CARRYB[519][2] , \CARRYB[519][1] , \CARRYB[519][0] ,
         \CARRYB[518][2] , \CARRYB[518][1] , \CARRYB[518][0] ,
         \CARRYB[517][2] , \CARRYB[517][1] , \CARRYB[517][0] ,
         \CARRYB[516][2] , \CARRYB[516][1] , \CARRYB[516][0] ,
         \CARRYB[515][2] , \CARRYB[515][1] , \CARRYB[515][0] ,
         \CARRYB[514][2] , \CARRYB[514][1] , \CARRYB[514][0] ,
         \CARRYB[513][2] , \CARRYB[513][1] , \CARRYB[513][0] ,
         \CARRYB[512][2] , \CARRYB[512][1] , \CARRYB[512][0] , \SUMB[639][2] ,
         \SUMB[639][1] , \SUMB[638][2] , \SUMB[638][1] , \SUMB[637][2] ,
         \SUMB[637][1] , \SUMB[636][2] , \SUMB[636][1] , \SUMB[635][2] ,
         \SUMB[635][1] , \SUMB[634][2] , \SUMB[634][1] , \SUMB[633][2] ,
         \SUMB[633][1] , \SUMB[632][2] , \SUMB[632][1] , \SUMB[631][2] ,
         \SUMB[631][1] , \SUMB[630][2] , \SUMB[630][1] , \SUMB[629][2] ,
         \SUMB[629][1] , \SUMB[628][2] , \SUMB[628][1] , \SUMB[627][2] ,
         \SUMB[627][1] , \SUMB[626][2] , \SUMB[626][1] , \SUMB[625][2] ,
         \SUMB[625][1] , \SUMB[624][2] , \SUMB[624][1] , \SUMB[623][2] ,
         \SUMB[623][1] , \SUMB[622][2] , \SUMB[622][1] , \SUMB[621][2] ,
         \SUMB[621][1] , \SUMB[620][2] , \SUMB[620][1] , \SUMB[619][2] ,
         \SUMB[619][1] , \SUMB[618][2] , \SUMB[618][1] , \SUMB[617][2] ,
         \SUMB[617][1] , \SUMB[616][2] , \SUMB[616][1] , \SUMB[615][2] ,
         \SUMB[615][1] , \SUMB[614][2] , \SUMB[614][1] , \SUMB[613][2] ,
         \SUMB[613][1] , \SUMB[612][2] , \SUMB[612][1] , \SUMB[611][2] ,
         \SUMB[611][1] , \SUMB[610][2] , \SUMB[610][1] , \SUMB[609][2] ,
         \SUMB[609][1] , \SUMB[608][2] , \SUMB[608][1] , \SUMB[607][2] ,
         \SUMB[607][1] , \SUMB[606][2] , \SUMB[606][1] , \SUMB[605][2] ,
         \SUMB[605][1] , \SUMB[604][2] , \SUMB[604][1] , \SUMB[603][2] ,
         \SUMB[603][1] , \SUMB[602][2] , \SUMB[602][1] , \SUMB[601][2] ,
         \SUMB[601][1] , \SUMB[600][2] , \SUMB[600][1] , \SUMB[599][2] ,
         \SUMB[599][1] , \SUMB[598][2] , \SUMB[598][1] , \SUMB[597][2] ,
         \SUMB[597][1] , \SUMB[596][2] , \SUMB[596][1] , \SUMB[595][2] ,
         \SUMB[595][1] , \SUMB[594][2] , \SUMB[594][1] , \SUMB[593][2] ,
         \SUMB[593][1] , \SUMB[592][2] , \SUMB[592][1] , \SUMB[591][2] ,
         \SUMB[591][1] , \SUMB[590][2] , \SUMB[590][1] , \SUMB[589][2] ,
         \SUMB[589][1] , \SUMB[588][2] , \SUMB[588][1] , \SUMB[587][2] ,
         \SUMB[587][1] , \SUMB[586][2] , \SUMB[586][1] , \SUMB[585][2] ,
         \SUMB[585][1] , \SUMB[584][2] , \SUMB[584][1] , \SUMB[583][2] ,
         \SUMB[583][1] , \SUMB[582][2] , \SUMB[582][1] , \SUMB[581][2] ,
         \SUMB[581][1] , \SUMB[580][2] , \SUMB[580][1] , \SUMB[579][2] ,
         \SUMB[579][1] , \SUMB[578][2] , \SUMB[578][1] , \SUMB[577][2] ,
         \SUMB[577][1] , \SUMB[576][2] , \SUMB[576][1] , \SUMB[575][2] ,
         \SUMB[575][1] , \SUMB[574][2] , \SUMB[574][1] , \SUMB[573][2] ,
         \SUMB[573][1] , \SUMB[572][2] , \SUMB[572][1] , \SUMB[571][2] ,
         \SUMB[571][1] , \SUMB[570][2] , \SUMB[570][1] , \SUMB[569][2] ,
         \SUMB[569][1] , \SUMB[568][2] , \SUMB[568][1] , \SUMB[567][2] ,
         \SUMB[567][1] , \SUMB[566][2] , \SUMB[566][1] , \SUMB[565][2] ,
         \SUMB[565][1] , \SUMB[564][2] , \SUMB[564][1] , \SUMB[563][2] ,
         \SUMB[563][1] , \SUMB[562][2] , \SUMB[562][1] , \SUMB[561][2] ,
         \SUMB[561][1] , \SUMB[560][2] , \SUMB[560][1] , \SUMB[559][2] ,
         \SUMB[559][1] , \SUMB[558][2] , \SUMB[558][1] , \SUMB[557][2] ,
         \SUMB[557][1] , \SUMB[556][2] , \SUMB[556][1] , \SUMB[555][2] ,
         \SUMB[555][1] , \SUMB[554][2] , \SUMB[554][1] , \SUMB[553][2] ,
         \SUMB[553][1] , \SUMB[552][2] , \SUMB[552][1] , \SUMB[551][2] ,
         \SUMB[551][1] , \SUMB[550][2] , \SUMB[550][1] , \SUMB[549][2] ,
         \SUMB[549][1] , \SUMB[548][2] , \SUMB[548][1] , \SUMB[547][2] ,
         \SUMB[547][1] , \SUMB[546][2] , \SUMB[546][1] , \SUMB[545][2] ,
         \SUMB[545][1] , \SUMB[544][2] , \SUMB[544][1] , \SUMB[543][2] ,
         \SUMB[543][1] , \SUMB[542][2] , \SUMB[542][1] , \SUMB[541][2] ,
         \SUMB[541][1] , \SUMB[540][2] , \SUMB[540][1] , \SUMB[539][2] ,
         \SUMB[539][1] , \SUMB[538][2] , \SUMB[538][1] , \SUMB[537][2] ,
         \SUMB[537][1] , \SUMB[536][2] , \SUMB[536][1] , \SUMB[535][2] ,
         \SUMB[535][1] , \SUMB[534][2] , \SUMB[534][1] , \SUMB[533][2] ,
         \SUMB[533][1] , \SUMB[532][2] , \SUMB[532][1] , \SUMB[531][2] ,
         \SUMB[531][1] , \SUMB[530][2] , \SUMB[530][1] , \SUMB[529][2] ,
         \SUMB[529][1] , \SUMB[528][2] , \SUMB[528][1] , \SUMB[527][2] ,
         \SUMB[527][1] , \SUMB[526][2] , \SUMB[526][1] , \SUMB[525][2] ,
         \SUMB[525][1] , \SUMB[524][2] , \SUMB[524][1] , \SUMB[523][2] ,
         \SUMB[523][1] , \SUMB[522][2] , \SUMB[522][1] , \SUMB[521][2] ,
         \SUMB[521][1] , \SUMB[520][2] , \SUMB[520][1] , \SUMB[519][2] ,
         \SUMB[519][1] , \SUMB[518][2] , \SUMB[518][1] , \SUMB[517][2] ,
         \SUMB[517][1] , \SUMB[516][2] , \SUMB[516][1] , \SUMB[515][2] ,
         \SUMB[515][1] , \SUMB[514][2] , \SUMB[514][1] , \SUMB[513][2] ,
         \SUMB[513][1] , \SUMB[512][2] , \SUMB[512][1] , \CARRYB[767][2] ,
         \CARRYB[767][1] , \CARRYB[767][0] , \CARRYB[766][2] ,
         \CARRYB[766][1] , \CARRYB[766][0] , \CARRYB[765][2] ,
         \CARRYB[765][1] , \CARRYB[765][0] , \CARRYB[764][2] ,
         \CARRYB[764][1] , \CARRYB[764][0] , \CARRYB[763][2] ,
         \CARRYB[763][1] , \CARRYB[763][0] , \CARRYB[762][2] ,
         \CARRYB[762][1] , \CARRYB[762][0] , \CARRYB[761][2] ,
         \CARRYB[761][1] , \CARRYB[761][0] , \CARRYB[760][2] ,
         \CARRYB[760][1] , \CARRYB[760][0] , \CARRYB[759][2] ,
         \CARRYB[759][1] , \CARRYB[759][0] , \CARRYB[758][2] ,
         \CARRYB[758][1] , \CARRYB[758][0] , \CARRYB[757][2] ,
         \CARRYB[757][1] , \CARRYB[757][0] , \CARRYB[756][2] ,
         \CARRYB[756][1] , \CARRYB[756][0] , \CARRYB[755][2] ,
         \CARRYB[755][1] , \CARRYB[755][0] , \CARRYB[754][2] ,
         \CARRYB[754][1] , \CARRYB[754][0] , \CARRYB[753][2] ,
         \CARRYB[753][1] , \CARRYB[753][0] , \CARRYB[752][2] ,
         \CARRYB[752][1] , \CARRYB[752][0] , \CARRYB[751][2] ,
         \CARRYB[751][1] , \CARRYB[751][0] , \CARRYB[750][2] ,
         \CARRYB[750][1] , \CARRYB[750][0] , \CARRYB[749][2] ,
         \CARRYB[749][1] , \CARRYB[749][0] , \CARRYB[748][2] ,
         \CARRYB[748][1] , \CARRYB[748][0] , \CARRYB[747][2] ,
         \CARRYB[747][1] , \CARRYB[747][0] , \CARRYB[746][2] ,
         \CARRYB[746][1] , \CARRYB[746][0] , \CARRYB[745][2] ,
         \CARRYB[745][1] , \CARRYB[745][0] , \CARRYB[744][2] ,
         \CARRYB[744][1] , \CARRYB[744][0] , \CARRYB[743][2] ,
         \CARRYB[743][1] , \CARRYB[743][0] , \CARRYB[742][2] ,
         \CARRYB[742][1] , \CARRYB[742][0] , \CARRYB[741][2] ,
         \CARRYB[741][1] , \CARRYB[741][0] , \CARRYB[740][2] ,
         \CARRYB[740][1] , \CARRYB[740][0] , \CARRYB[739][2] ,
         \CARRYB[739][1] , \CARRYB[739][0] , \CARRYB[738][2] ,
         \CARRYB[738][1] , \CARRYB[738][0] , \CARRYB[737][2] ,
         \CARRYB[737][1] , \CARRYB[737][0] , \CARRYB[736][2] ,
         \CARRYB[736][1] , \CARRYB[736][0] , \CARRYB[735][2] ,
         \CARRYB[735][1] , \CARRYB[735][0] , \CARRYB[734][2] ,
         \CARRYB[734][1] , \CARRYB[734][0] , \CARRYB[733][2] ,
         \CARRYB[733][1] , \CARRYB[733][0] , \CARRYB[732][2] ,
         \CARRYB[732][1] , \CARRYB[732][0] , \CARRYB[731][2] ,
         \CARRYB[731][1] , \CARRYB[731][0] , \CARRYB[730][2] ,
         \CARRYB[730][1] , \CARRYB[730][0] , \CARRYB[729][2] ,
         \CARRYB[729][1] , \CARRYB[729][0] , \CARRYB[728][2] ,
         \CARRYB[728][1] , \CARRYB[728][0] , \CARRYB[727][2] ,
         \CARRYB[727][1] , \CARRYB[727][0] , \CARRYB[726][2] ,
         \CARRYB[726][1] , \CARRYB[726][0] , \CARRYB[725][2] ,
         \CARRYB[725][1] , \CARRYB[725][0] , \CARRYB[724][2] ,
         \CARRYB[724][1] , \CARRYB[724][0] , \CARRYB[723][2] ,
         \CARRYB[723][1] , \CARRYB[723][0] , \CARRYB[722][2] ,
         \CARRYB[722][1] , \CARRYB[722][0] , \CARRYB[721][2] ,
         \CARRYB[721][1] , \CARRYB[721][0] , \CARRYB[720][2] ,
         \CARRYB[720][1] , \CARRYB[720][0] , \CARRYB[719][2] ,
         \CARRYB[719][1] , \CARRYB[719][0] , \CARRYB[718][2] ,
         \CARRYB[718][1] , \CARRYB[718][0] , \CARRYB[717][2] ,
         \CARRYB[717][1] , \CARRYB[717][0] , \CARRYB[716][2] ,
         \CARRYB[716][1] , \CARRYB[716][0] , \CARRYB[715][2] ,
         \CARRYB[715][1] , \CARRYB[715][0] , \CARRYB[714][2] ,
         \CARRYB[714][1] , \CARRYB[714][0] , \CARRYB[713][2] ,
         \CARRYB[713][1] , \CARRYB[713][0] , \CARRYB[712][2] ,
         \CARRYB[712][1] , \CARRYB[712][0] , \CARRYB[711][2] ,
         \CARRYB[711][1] , \CARRYB[711][0] , \CARRYB[710][2] ,
         \CARRYB[710][1] , \CARRYB[710][0] , \CARRYB[709][2] ,
         \CARRYB[709][1] , \CARRYB[709][0] , \CARRYB[708][2] ,
         \CARRYB[708][1] , \CARRYB[708][0] , \CARRYB[707][2] ,
         \CARRYB[707][1] , \CARRYB[707][0] , \CARRYB[706][2] ,
         \CARRYB[706][1] , \CARRYB[706][0] , \CARRYB[705][2] ,
         \CARRYB[705][1] , \CARRYB[705][0] , \CARRYB[704][2] ,
         \CARRYB[704][1] , \CARRYB[704][0] , \CARRYB[703][2] ,
         \CARRYB[703][1] , \CARRYB[703][0] , \CARRYB[702][2] ,
         \CARRYB[702][1] , \CARRYB[702][0] , \CARRYB[701][2] ,
         \CARRYB[701][1] , \CARRYB[701][0] , \CARRYB[700][2] ,
         \CARRYB[700][1] , \CARRYB[700][0] , \CARRYB[699][2] ,
         \CARRYB[699][1] , \CARRYB[699][0] , \CARRYB[698][2] ,
         \CARRYB[698][1] , \CARRYB[698][0] , \CARRYB[697][2] ,
         \CARRYB[697][1] , \CARRYB[697][0] , \CARRYB[696][2] ,
         \CARRYB[696][1] , \CARRYB[696][0] , \CARRYB[695][2] ,
         \CARRYB[695][1] , \CARRYB[695][0] , \CARRYB[694][2] ,
         \CARRYB[694][1] , \CARRYB[694][0] , \CARRYB[693][2] ,
         \CARRYB[693][1] , \CARRYB[693][0] , \CARRYB[692][2] ,
         \CARRYB[692][1] , \CARRYB[692][0] , \CARRYB[691][2] ,
         \CARRYB[691][1] , \CARRYB[691][0] , \CARRYB[690][2] ,
         \CARRYB[690][1] , \CARRYB[690][0] , \CARRYB[689][2] ,
         \CARRYB[689][1] , \CARRYB[689][0] , \CARRYB[688][2] ,
         \CARRYB[688][1] , \CARRYB[688][0] , \CARRYB[687][2] ,
         \CARRYB[687][1] , \CARRYB[687][0] , \CARRYB[686][2] ,
         \CARRYB[686][1] , \CARRYB[686][0] , \CARRYB[685][2] ,
         \CARRYB[685][1] , \CARRYB[685][0] , \CARRYB[684][2] ,
         \CARRYB[684][1] , \CARRYB[684][0] , \CARRYB[683][2] ,
         \CARRYB[683][1] , \CARRYB[683][0] , \CARRYB[682][2] ,
         \CARRYB[682][1] , \CARRYB[682][0] , \CARRYB[681][2] ,
         \CARRYB[681][1] , \CARRYB[681][0] , \CARRYB[680][2] ,
         \CARRYB[680][1] , \CARRYB[680][0] , \CARRYB[679][2] ,
         \CARRYB[679][1] , \CARRYB[679][0] , \CARRYB[678][2] ,
         \CARRYB[678][1] , \CARRYB[678][0] , \CARRYB[677][2] ,
         \CARRYB[677][1] , \CARRYB[677][0] , \CARRYB[676][2] ,
         \CARRYB[676][1] , \CARRYB[676][0] , \CARRYB[675][2] ,
         \CARRYB[675][1] , \CARRYB[675][0] , \CARRYB[674][2] ,
         \CARRYB[674][1] , \CARRYB[674][0] , \CARRYB[673][2] ,
         \CARRYB[673][1] , \CARRYB[673][0] , \CARRYB[672][2] ,
         \CARRYB[672][1] , \CARRYB[672][0] , \CARRYB[671][2] ,
         \CARRYB[671][1] , \CARRYB[671][0] , \CARRYB[670][2] ,
         \CARRYB[670][1] , \CARRYB[670][0] , \CARRYB[669][2] ,
         \CARRYB[669][1] , \CARRYB[669][0] , \CARRYB[668][2] ,
         \CARRYB[668][1] , \CARRYB[668][0] , \CARRYB[667][2] ,
         \CARRYB[667][1] , \CARRYB[667][0] , \CARRYB[666][2] ,
         \CARRYB[666][1] , \CARRYB[666][0] , \CARRYB[665][2] ,
         \CARRYB[665][1] , \CARRYB[665][0] , \CARRYB[664][2] ,
         \CARRYB[664][1] , \CARRYB[664][0] , \CARRYB[663][2] ,
         \CARRYB[663][1] , \CARRYB[663][0] , \CARRYB[662][2] ,
         \CARRYB[662][1] , \CARRYB[662][0] , \CARRYB[661][2] ,
         \CARRYB[661][1] , \CARRYB[661][0] , \CARRYB[660][2] ,
         \CARRYB[660][1] , \CARRYB[660][0] , \CARRYB[659][2] ,
         \CARRYB[659][1] , \CARRYB[659][0] , \CARRYB[658][2] ,
         \CARRYB[658][1] , \CARRYB[658][0] , \CARRYB[657][2] ,
         \CARRYB[657][1] , \CARRYB[657][0] , \CARRYB[656][2] ,
         \CARRYB[656][1] , \CARRYB[656][0] , \CARRYB[655][2] ,
         \CARRYB[655][1] , \CARRYB[655][0] , \CARRYB[654][2] ,
         \CARRYB[654][1] , \CARRYB[654][0] , \CARRYB[653][2] ,
         \CARRYB[653][1] , \CARRYB[653][0] , \CARRYB[652][2] ,
         \CARRYB[652][1] , \CARRYB[652][0] , \CARRYB[651][2] ,
         \CARRYB[651][1] , \CARRYB[651][0] , \CARRYB[650][2] ,
         \CARRYB[650][1] , \CARRYB[650][0] , \CARRYB[649][2] ,
         \CARRYB[649][1] , \CARRYB[649][0] , \CARRYB[648][2] ,
         \CARRYB[648][1] , \CARRYB[648][0] , \CARRYB[647][2] ,
         \CARRYB[647][1] , \CARRYB[647][0] , \CARRYB[646][2] ,
         \CARRYB[646][1] , \CARRYB[646][0] , \CARRYB[645][2] ,
         \CARRYB[645][1] , \CARRYB[645][0] , \CARRYB[644][2] ,
         \CARRYB[644][1] , \CARRYB[644][0] , \CARRYB[643][2] ,
         \CARRYB[643][1] , \CARRYB[643][0] , \CARRYB[642][2] ,
         \CARRYB[642][1] , \CARRYB[642][0] , \CARRYB[641][2] ,
         \CARRYB[641][1] , \CARRYB[641][0] , \CARRYB[640][2] ,
         \CARRYB[640][1] , \CARRYB[640][0] , \SUMB[767][2] , \SUMB[767][1] ,
         \SUMB[766][2] , \SUMB[766][1] , \SUMB[765][2] , \SUMB[765][1] ,
         \SUMB[764][2] , \SUMB[764][1] , \SUMB[763][2] , \SUMB[763][1] ,
         \SUMB[762][2] , \SUMB[762][1] , \SUMB[761][2] , \SUMB[761][1] ,
         \SUMB[760][2] , \SUMB[760][1] , \SUMB[759][2] , \SUMB[759][1] ,
         \SUMB[758][2] , \SUMB[758][1] , \SUMB[757][2] , \SUMB[757][1] ,
         \SUMB[756][2] , \SUMB[756][1] , \SUMB[755][2] , \SUMB[755][1] ,
         \SUMB[754][2] , \SUMB[754][1] , \SUMB[753][2] , \SUMB[753][1] ,
         \SUMB[752][2] , \SUMB[752][1] , \SUMB[751][2] , \SUMB[751][1] ,
         \SUMB[750][2] , \SUMB[750][1] , \SUMB[749][2] , \SUMB[749][1] ,
         \SUMB[748][2] , \SUMB[748][1] , \SUMB[747][2] , \SUMB[747][1] ,
         \SUMB[746][2] , \SUMB[746][1] , \SUMB[745][2] , \SUMB[745][1] ,
         \SUMB[744][2] , \SUMB[744][1] , \SUMB[743][2] , \SUMB[743][1] ,
         \SUMB[742][2] , \SUMB[742][1] , \SUMB[741][2] , \SUMB[741][1] ,
         \SUMB[740][2] , \SUMB[740][1] , \SUMB[739][2] , \SUMB[739][1] ,
         \SUMB[738][2] , \SUMB[738][1] , \SUMB[737][2] , \SUMB[737][1] ,
         \SUMB[736][2] , \SUMB[736][1] , \SUMB[735][2] , \SUMB[735][1] ,
         \SUMB[734][2] , \SUMB[734][1] , \SUMB[733][2] , \SUMB[733][1] ,
         \SUMB[732][2] , \SUMB[732][1] , \SUMB[731][2] , \SUMB[731][1] ,
         \SUMB[730][2] , \SUMB[730][1] , \SUMB[729][2] , \SUMB[729][1] ,
         \SUMB[728][2] , \SUMB[728][1] , \SUMB[727][2] , \SUMB[727][1] ,
         \SUMB[726][2] , \SUMB[726][1] , \SUMB[725][2] , \SUMB[725][1] ,
         \SUMB[724][2] , \SUMB[724][1] , \SUMB[723][2] , \SUMB[723][1] ,
         \SUMB[722][2] , \SUMB[722][1] , \SUMB[721][2] , \SUMB[721][1] ,
         \SUMB[720][2] , \SUMB[720][1] , \SUMB[719][2] , \SUMB[719][1] ,
         \SUMB[718][2] , \SUMB[718][1] , \SUMB[717][2] , \SUMB[717][1] ,
         \SUMB[716][2] , \SUMB[716][1] , \SUMB[715][2] , \SUMB[715][1] ,
         \SUMB[714][2] , \SUMB[714][1] , \SUMB[713][2] , \SUMB[713][1] ,
         \SUMB[712][2] , \SUMB[712][1] , \SUMB[711][2] , \SUMB[711][1] ,
         \SUMB[710][2] , \SUMB[710][1] , \SUMB[709][2] , \SUMB[709][1] ,
         \SUMB[708][2] , \SUMB[708][1] , \SUMB[707][2] , \SUMB[707][1] ,
         \SUMB[706][2] , \SUMB[706][1] , \SUMB[705][2] , \SUMB[705][1] ,
         \SUMB[704][2] , \SUMB[704][1] , \SUMB[703][2] , \SUMB[703][1] ,
         \SUMB[702][2] , \SUMB[702][1] , \SUMB[701][2] , \SUMB[701][1] ,
         \SUMB[700][2] , \SUMB[700][1] , \SUMB[699][2] , \SUMB[699][1] ,
         \SUMB[698][2] , \SUMB[698][1] , \SUMB[697][2] , \SUMB[697][1] ,
         \SUMB[696][2] , \SUMB[696][1] , \SUMB[695][2] , \SUMB[695][1] ,
         \SUMB[694][2] , \SUMB[694][1] , \SUMB[693][2] , \SUMB[693][1] ,
         \SUMB[692][2] , \SUMB[692][1] , \SUMB[691][2] , \SUMB[691][1] ,
         \SUMB[690][2] , \SUMB[690][1] , \SUMB[689][2] , \SUMB[689][1] ,
         \SUMB[688][2] , \SUMB[688][1] , \SUMB[687][2] , \SUMB[687][1] ,
         \SUMB[686][2] , \SUMB[686][1] , \SUMB[685][2] , \SUMB[685][1] ,
         \SUMB[684][2] , \SUMB[684][1] , \SUMB[683][2] , \SUMB[683][1] ,
         \SUMB[682][2] , \SUMB[682][1] , \SUMB[681][2] , \SUMB[681][1] ,
         \SUMB[680][2] , \SUMB[680][1] , \SUMB[679][2] , \SUMB[679][1] ,
         \SUMB[678][2] , \SUMB[678][1] , \SUMB[677][2] , \SUMB[677][1] ,
         \SUMB[676][2] , \SUMB[676][1] , \SUMB[675][2] , \SUMB[675][1] ,
         \SUMB[674][2] , \SUMB[674][1] , \SUMB[673][2] , \SUMB[673][1] ,
         \SUMB[672][2] , \SUMB[672][1] , \SUMB[671][2] , \SUMB[671][1] ,
         \SUMB[670][2] , \SUMB[670][1] , \SUMB[669][2] , \SUMB[669][1] ,
         \SUMB[668][2] , \SUMB[668][1] , \SUMB[667][2] , \SUMB[667][1] ,
         \SUMB[666][2] , \SUMB[666][1] , \SUMB[665][2] , \SUMB[665][1] ,
         \SUMB[664][2] , \SUMB[664][1] , \SUMB[663][2] , \SUMB[663][1] ,
         \SUMB[662][2] , \SUMB[662][1] , \SUMB[661][2] , \SUMB[661][1] ,
         \SUMB[660][2] , \SUMB[660][1] , \SUMB[659][2] , \SUMB[659][1] ,
         \SUMB[658][2] , \SUMB[658][1] , \SUMB[657][2] , \SUMB[657][1] ,
         \SUMB[656][2] , \SUMB[656][1] , \SUMB[655][2] , \SUMB[655][1] ,
         \SUMB[654][2] , \SUMB[654][1] , \SUMB[653][2] , \SUMB[653][1] ,
         \SUMB[652][2] , \SUMB[652][1] , \SUMB[651][2] , \SUMB[651][1] ,
         \SUMB[650][2] , \SUMB[650][1] , \SUMB[649][2] , \SUMB[649][1] ,
         \SUMB[648][2] , \SUMB[648][1] , \SUMB[647][2] , \SUMB[647][1] ,
         \SUMB[646][2] , \SUMB[646][1] , \SUMB[645][2] , \SUMB[645][1] ,
         \SUMB[644][2] , \SUMB[644][1] , \SUMB[643][2] , \SUMB[643][1] ,
         \SUMB[642][2] , \SUMB[642][1] , \SUMB[641][2] , \SUMB[641][1] ,
         \SUMB[640][2] , \SUMB[640][1] , \CARRYB[895][2] , \CARRYB[895][1] ,
         \CARRYB[895][0] , \CARRYB[894][2] , \CARRYB[894][1] ,
         \CARRYB[894][0] , \CARRYB[893][2] , \CARRYB[893][1] ,
         \CARRYB[893][0] , \CARRYB[892][2] , \CARRYB[892][1] ,
         \CARRYB[892][0] , \CARRYB[891][2] , \CARRYB[891][1] ,
         \CARRYB[891][0] , \CARRYB[890][2] , \CARRYB[890][1] ,
         \CARRYB[890][0] , \CARRYB[889][2] , \CARRYB[889][1] ,
         \CARRYB[889][0] , \CARRYB[888][2] , \CARRYB[888][1] ,
         \CARRYB[888][0] , \CARRYB[887][2] , \CARRYB[887][1] ,
         \CARRYB[887][0] , \CARRYB[886][2] , \CARRYB[886][1] ,
         \CARRYB[886][0] , \CARRYB[885][2] , \CARRYB[885][1] ,
         \CARRYB[885][0] , \CARRYB[884][2] , \CARRYB[884][1] ,
         \CARRYB[884][0] , \CARRYB[883][2] , \CARRYB[883][1] ,
         \CARRYB[883][0] , \CARRYB[882][2] , \CARRYB[882][1] ,
         \CARRYB[882][0] , \CARRYB[881][2] , \CARRYB[881][1] ,
         \CARRYB[881][0] , \CARRYB[880][2] , \CARRYB[880][1] ,
         \CARRYB[880][0] , \CARRYB[879][2] , \CARRYB[879][1] ,
         \CARRYB[879][0] , \CARRYB[878][2] , \CARRYB[878][1] ,
         \CARRYB[878][0] , \CARRYB[877][2] , \CARRYB[877][1] ,
         \CARRYB[877][0] , \CARRYB[876][2] , \CARRYB[876][1] ,
         \CARRYB[876][0] , \CARRYB[875][2] , \CARRYB[875][1] ,
         \CARRYB[875][0] , \CARRYB[874][2] , \CARRYB[874][1] ,
         \CARRYB[874][0] , \CARRYB[873][2] , \CARRYB[873][1] ,
         \CARRYB[873][0] , \CARRYB[872][2] , \CARRYB[872][1] ,
         \CARRYB[872][0] , \CARRYB[871][2] , \CARRYB[871][1] ,
         \CARRYB[871][0] , \CARRYB[870][2] , \CARRYB[870][1] ,
         \CARRYB[870][0] , \CARRYB[869][2] , \CARRYB[869][1] ,
         \CARRYB[869][0] , \CARRYB[868][2] , \CARRYB[868][1] ,
         \CARRYB[868][0] , \CARRYB[867][2] , \CARRYB[867][1] ,
         \CARRYB[867][0] , \CARRYB[866][2] , \CARRYB[866][1] ,
         \CARRYB[866][0] , \CARRYB[865][2] , \CARRYB[865][1] ,
         \CARRYB[865][0] , \CARRYB[864][2] , \CARRYB[864][1] ,
         \CARRYB[864][0] , \CARRYB[863][2] , \CARRYB[863][1] ,
         \CARRYB[863][0] , \CARRYB[862][2] , \CARRYB[862][1] ,
         \CARRYB[862][0] , \CARRYB[861][2] , \CARRYB[861][1] ,
         \CARRYB[861][0] , \CARRYB[860][2] , \CARRYB[860][1] ,
         \CARRYB[860][0] , \CARRYB[859][2] , \CARRYB[859][1] ,
         \CARRYB[859][0] , \CARRYB[858][2] , \CARRYB[858][1] ,
         \CARRYB[858][0] , \CARRYB[857][2] , \CARRYB[857][1] ,
         \CARRYB[857][0] , \CARRYB[856][2] , \CARRYB[856][1] ,
         \CARRYB[856][0] , \CARRYB[855][2] , \CARRYB[855][1] ,
         \CARRYB[855][0] , \CARRYB[854][2] , \CARRYB[854][1] ,
         \CARRYB[854][0] , \CARRYB[853][2] , \CARRYB[853][1] ,
         \CARRYB[853][0] , \CARRYB[852][2] , \CARRYB[852][1] ,
         \CARRYB[852][0] , \CARRYB[851][2] , \CARRYB[851][1] ,
         \CARRYB[851][0] , \CARRYB[850][2] , \CARRYB[850][1] ,
         \CARRYB[850][0] , \CARRYB[849][2] , \CARRYB[849][1] ,
         \CARRYB[849][0] , \CARRYB[848][2] , \CARRYB[848][1] ,
         \CARRYB[848][0] , \CARRYB[847][2] , \CARRYB[847][1] ,
         \CARRYB[847][0] , \CARRYB[846][2] , \CARRYB[846][1] ,
         \CARRYB[846][0] , \CARRYB[845][2] , \CARRYB[845][1] ,
         \CARRYB[845][0] , \CARRYB[844][2] , \CARRYB[844][1] ,
         \CARRYB[844][0] , \CARRYB[843][2] , \CARRYB[843][1] ,
         \CARRYB[843][0] , \CARRYB[842][2] , \CARRYB[842][1] ,
         \CARRYB[842][0] , \CARRYB[841][2] , \CARRYB[841][1] ,
         \CARRYB[841][0] , \CARRYB[840][2] , \CARRYB[840][1] ,
         \CARRYB[840][0] , \CARRYB[839][2] , \CARRYB[839][1] ,
         \CARRYB[839][0] , \CARRYB[838][2] , \CARRYB[838][1] ,
         \CARRYB[838][0] , \CARRYB[837][2] , \CARRYB[837][1] ,
         \CARRYB[837][0] , \CARRYB[836][2] , \CARRYB[836][1] ,
         \CARRYB[836][0] , \CARRYB[835][2] , \CARRYB[835][1] ,
         \CARRYB[835][0] , \CARRYB[834][2] , \CARRYB[834][1] ,
         \CARRYB[834][0] , \CARRYB[833][2] , \CARRYB[833][1] ,
         \CARRYB[833][0] , \CARRYB[832][2] , \CARRYB[832][1] ,
         \CARRYB[832][0] , \CARRYB[831][2] , \CARRYB[831][1] ,
         \CARRYB[831][0] , \CARRYB[830][2] , \CARRYB[830][1] ,
         \CARRYB[830][0] , \CARRYB[829][2] , \CARRYB[829][1] ,
         \CARRYB[829][0] , \CARRYB[828][2] , \CARRYB[828][1] ,
         \CARRYB[828][0] , \CARRYB[827][2] , \CARRYB[827][1] ,
         \CARRYB[827][0] , \CARRYB[826][2] , \CARRYB[826][1] ,
         \CARRYB[826][0] , \CARRYB[825][2] , \CARRYB[825][1] ,
         \CARRYB[825][0] , \CARRYB[824][2] , \CARRYB[824][1] ,
         \CARRYB[824][0] , \CARRYB[823][2] , \CARRYB[823][1] ,
         \CARRYB[823][0] , \CARRYB[822][2] , \CARRYB[822][1] ,
         \CARRYB[822][0] , \CARRYB[821][2] , \CARRYB[821][1] ,
         \CARRYB[821][0] , \CARRYB[820][2] , \CARRYB[820][1] ,
         \CARRYB[820][0] , \CARRYB[819][2] , \CARRYB[819][1] ,
         \CARRYB[819][0] , \CARRYB[818][2] , \CARRYB[818][1] ,
         \CARRYB[818][0] , \CARRYB[817][2] , \CARRYB[817][1] ,
         \CARRYB[817][0] , \CARRYB[816][2] , \CARRYB[816][1] ,
         \CARRYB[816][0] , \CARRYB[815][2] , \CARRYB[815][1] ,
         \CARRYB[815][0] , \CARRYB[814][2] , \CARRYB[814][1] ,
         \CARRYB[814][0] , \CARRYB[813][2] , \CARRYB[813][1] ,
         \CARRYB[813][0] , \CARRYB[812][2] , \CARRYB[812][1] ,
         \CARRYB[812][0] , \CARRYB[811][2] , \CARRYB[811][1] ,
         \CARRYB[811][0] , \CARRYB[810][2] , \CARRYB[810][1] ,
         \CARRYB[810][0] , \CARRYB[809][2] , \CARRYB[809][1] ,
         \CARRYB[809][0] , \CARRYB[808][2] , \CARRYB[808][1] ,
         \CARRYB[808][0] , \CARRYB[807][2] , \CARRYB[807][1] ,
         \CARRYB[807][0] , \CARRYB[806][2] , \CARRYB[806][1] ,
         \CARRYB[806][0] , \CARRYB[805][2] , \CARRYB[805][1] ,
         \CARRYB[805][0] , \CARRYB[804][2] , \CARRYB[804][1] ,
         \CARRYB[804][0] , \CARRYB[803][2] , \CARRYB[803][1] ,
         \CARRYB[803][0] , \CARRYB[802][2] , \CARRYB[802][1] ,
         \CARRYB[802][0] , \CARRYB[801][2] , \CARRYB[801][1] ,
         \CARRYB[801][0] , \CARRYB[800][2] , \CARRYB[800][1] ,
         \CARRYB[800][0] , \CARRYB[799][2] , \CARRYB[799][1] ,
         \CARRYB[799][0] , \CARRYB[798][2] , \CARRYB[798][1] ,
         \CARRYB[798][0] , \CARRYB[797][2] , \CARRYB[797][1] ,
         \CARRYB[797][0] , \CARRYB[796][2] , \CARRYB[796][1] ,
         \CARRYB[796][0] , \CARRYB[795][2] , \CARRYB[795][1] ,
         \CARRYB[795][0] , \CARRYB[794][2] , \CARRYB[794][1] ,
         \CARRYB[794][0] , \CARRYB[793][2] , \CARRYB[793][1] ,
         \CARRYB[793][0] , \CARRYB[792][2] , \CARRYB[792][1] ,
         \CARRYB[792][0] , \CARRYB[791][2] , \CARRYB[791][1] ,
         \CARRYB[791][0] , \CARRYB[790][2] , \CARRYB[790][1] ,
         \CARRYB[790][0] , \CARRYB[789][2] , \CARRYB[789][1] ,
         \CARRYB[789][0] , \CARRYB[788][2] , \CARRYB[788][1] ,
         \CARRYB[788][0] , \CARRYB[787][2] , \CARRYB[787][1] ,
         \CARRYB[787][0] , \CARRYB[786][2] , \CARRYB[786][1] ,
         \CARRYB[786][0] , \CARRYB[785][2] , \CARRYB[785][1] ,
         \CARRYB[785][0] , \CARRYB[784][2] , \CARRYB[784][1] ,
         \CARRYB[784][0] , \CARRYB[783][2] , \CARRYB[783][1] ,
         \CARRYB[783][0] , \CARRYB[782][2] , \CARRYB[782][1] ,
         \CARRYB[782][0] , \CARRYB[781][2] , \CARRYB[781][1] ,
         \CARRYB[781][0] , \CARRYB[780][2] , \CARRYB[780][1] ,
         \CARRYB[780][0] , \CARRYB[779][2] , \CARRYB[779][1] ,
         \CARRYB[779][0] , \CARRYB[778][2] , \CARRYB[778][1] ,
         \CARRYB[778][0] , \CARRYB[777][2] , \CARRYB[777][1] ,
         \CARRYB[777][0] , \CARRYB[776][2] , \CARRYB[776][1] ,
         \CARRYB[776][0] , \CARRYB[775][2] , \CARRYB[775][1] ,
         \CARRYB[775][0] , \CARRYB[774][2] , \CARRYB[774][1] ,
         \CARRYB[774][0] , \CARRYB[773][2] , \CARRYB[773][1] ,
         \CARRYB[773][0] , \CARRYB[772][2] , \CARRYB[772][1] ,
         \CARRYB[772][0] , \CARRYB[771][2] , \CARRYB[771][1] ,
         \CARRYB[771][0] , \CARRYB[770][2] , \CARRYB[770][1] ,
         \CARRYB[770][0] , \CARRYB[769][2] , \CARRYB[769][1] ,
         \CARRYB[769][0] , \CARRYB[768][2] , \CARRYB[768][1] ,
         \CARRYB[768][0] , \SUMB[895][2] , \SUMB[895][1] , \SUMB[894][2] ,
         \SUMB[894][1] , \SUMB[893][2] , \SUMB[893][1] , \SUMB[892][2] ,
         \SUMB[892][1] , \SUMB[891][2] , \SUMB[891][1] , \SUMB[890][2] ,
         \SUMB[890][1] , \SUMB[889][2] , \SUMB[889][1] , \SUMB[888][2] ,
         \SUMB[888][1] , \SUMB[887][2] , \SUMB[887][1] , \SUMB[886][2] ,
         \SUMB[886][1] , \SUMB[885][2] , \SUMB[885][1] , \SUMB[884][2] ,
         \SUMB[884][1] , \SUMB[883][2] , \SUMB[883][1] , \SUMB[882][2] ,
         \SUMB[882][1] , \SUMB[881][2] , \SUMB[881][1] , \SUMB[880][2] ,
         \SUMB[880][1] , \SUMB[879][2] , \SUMB[879][1] , \SUMB[878][2] ,
         \SUMB[878][1] , \SUMB[877][2] , \SUMB[877][1] , \SUMB[876][2] ,
         \SUMB[876][1] , \SUMB[875][2] , \SUMB[875][1] , \SUMB[874][2] ,
         \SUMB[874][1] , \SUMB[873][2] , \SUMB[873][1] , \SUMB[872][2] ,
         \SUMB[872][1] , \SUMB[871][2] , \SUMB[871][1] , \SUMB[870][2] ,
         \SUMB[870][1] , \SUMB[869][2] , \SUMB[869][1] , \SUMB[868][2] ,
         \SUMB[868][1] , \SUMB[867][2] , \SUMB[867][1] , \SUMB[866][2] ,
         \SUMB[866][1] , \SUMB[865][2] , \SUMB[865][1] , \SUMB[864][2] ,
         \SUMB[864][1] , \SUMB[863][2] , \SUMB[863][1] , \SUMB[862][2] ,
         \SUMB[862][1] , \SUMB[861][2] , \SUMB[861][1] , \SUMB[860][2] ,
         \SUMB[860][1] , \SUMB[859][2] , \SUMB[859][1] , \SUMB[858][2] ,
         \SUMB[858][1] , \SUMB[857][2] , \SUMB[857][1] , \SUMB[856][2] ,
         \SUMB[856][1] , \SUMB[855][2] , \SUMB[855][1] , \SUMB[854][2] ,
         \SUMB[854][1] , \SUMB[853][2] , \SUMB[853][1] , \SUMB[852][2] ,
         \SUMB[852][1] , \SUMB[851][2] , \SUMB[851][1] , \SUMB[850][2] ,
         \SUMB[850][1] , \SUMB[849][2] , \SUMB[849][1] , \SUMB[848][2] ,
         \SUMB[848][1] , \SUMB[847][2] , \SUMB[847][1] , \SUMB[846][2] ,
         \SUMB[846][1] , \SUMB[845][2] , \SUMB[845][1] , \SUMB[844][2] ,
         \SUMB[844][1] , \SUMB[843][2] , \SUMB[843][1] , \SUMB[842][2] ,
         \SUMB[842][1] , \SUMB[841][2] , \SUMB[841][1] , \SUMB[840][2] ,
         \SUMB[840][1] , \SUMB[839][2] , \SUMB[839][1] , \SUMB[838][2] ,
         \SUMB[838][1] , \SUMB[837][2] , \SUMB[837][1] , \SUMB[836][2] ,
         \SUMB[836][1] , \SUMB[835][2] , \SUMB[835][1] , \SUMB[834][2] ,
         \SUMB[834][1] , \SUMB[833][2] , \SUMB[833][1] , \SUMB[832][2] ,
         \SUMB[832][1] , \SUMB[831][2] , \SUMB[831][1] , \SUMB[830][2] ,
         \SUMB[830][1] , \SUMB[829][2] , \SUMB[829][1] , \SUMB[828][2] ,
         \SUMB[828][1] , \SUMB[827][2] , \SUMB[827][1] , \SUMB[826][2] ,
         \SUMB[826][1] , \SUMB[825][2] , \SUMB[825][1] , \SUMB[824][2] ,
         \SUMB[824][1] , \SUMB[823][2] , \SUMB[823][1] , \SUMB[822][2] ,
         \SUMB[822][1] , \SUMB[821][2] , \SUMB[821][1] , \SUMB[820][2] ,
         \SUMB[820][1] , \SUMB[819][2] , \SUMB[819][1] , \SUMB[818][2] ,
         \SUMB[818][1] , \SUMB[817][2] , \SUMB[817][1] , \SUMB[816][2] ,
         \SUMB[816][1] , \SUMB[815][2] , \SUMB[815][1] , \SUMB[814][2] ,
         \SUMB[814][1] , \SUMB[813][2] , \SUMB[813][1] , \SUMB[812][2] ,
         \SUMB[812][1] , \SUMB[811][2] , \SUMB[811][1] , \SUMB[810][2] ,
         \SUMB[810][1] , \SUMB[809][2] , \SUMB[809][1] , \SUMB[808][2] ,
         \SUMB[808][1] , \SUMB[807][2] , \SUMB[807][1] , \SUMB[806][2] ,
         \SUMB[806][1] , \SUMB[805][2] , \SUMB[805][1] , \SUMB[804][2] ,
         \SUMB[804][1] , \SUMB[803][2] , \SUMB[803][1] , \SUMB[802][2] ,
         \SUMB[802][1] , \SUMB[801][2] , \SUMB[801][1] , \SUMB[800][2] ,
         \SUMB[800][1] , \SUMB[799][2] , \SUMB[799][1] , \SUMB[798][2] ,
         \SUMB[798][1] , \SUMB[797][2] , \SUMB[797][1] , \SUMB[796][2] ,
         \SUMB[796][1] , \SUMB[795][2] , \SUMB[795][1] , \SUMB[794][2] ,
         \SUMB[794][1] , \SUMB[793][2] , \SUMB[793][1] , \SUMB[792][2] ,
         \SUMB[792][1] , \SUMB[791][2] , \SUMB[791][1] , \SUMB[790][2] ,
         \SUMB[790][1] , \SUMB[789][2] , \SUMB[789][1] , \SUMB[788][2] ,
         \SUMB[788][1] , \SUMB[787][2] , \SUMB[787][1] , \SUMB[786][2] ,
         \SUMB[786][1] , \SUMB[785][2] , \SUMB[785][1] , \SUMB[784][2] ,
         \SUMB[784][1] , \SUMB[783][2] , \SUMB[783][1] , \SUMB[782][2] ,
         \SUMB[782][1] , \SUMB[781][2] , \SUMB[781][1] , \SUMB[780][2] ,
         \SUMB[780][1] , \SUMB[779][2] , \SUMB[779][1] , \SUMB[778][2] ,
         \SUMB[778][1] , \SUMB[777][2] , \SUMB[777][1] , \SUMB[776][2] ,
         \SUMB[776][1] , \SUMB[775][2] , \SUMB[775][1] , \SUMB[774][2] ,
         \SUMB[774][1] , \SUMB[773][2] , \SUMB[773][1] , \SUMB[772][2] ,
         \SUMB[772][1] , \SUMB[771][2] , \SUMB[771][1] , \SUMB[770][2] ,
         \SUMB[770][1] , \SUMB[769][2] , \SUMB[769][1] , \SUMB[768][2] ,
         \SUMB[768][1] , \CARRYB[1022][0] , \CARRYB[1021][1] ,
         \CARRYB[1021][0] , \CARRYB[1020][2] , \CARRYB[1020][1] ,
         \CARRYB[1020][0] , \CARRYB[1019][2] , \CARRYB[1019][1] ,
         \CARRYB[1019][0] , \CARRYB[1018][2] , \CARRYB[1018][1] ,
         \CARRYB[1018][0] , \CARRYB[1017][2] , \CARRYB[1017][1] ,
         \CARRYB[1017][0] , \CARRYB[1016][2] , \CARRYB[1016][1] ,
         \CARRYB[1016][0] , \CARRYB[1015][2] , \CARRYB[1015][1] ,
         \CARRYB[1015][0] , \CARRYB[1014][2] , \CARRYB[1014][1] ,
         \CARRYB[1014][0] , \CARRYB[1013][2] , \CARRYB[1013][1] ,
         \CARRYB[1013][0] , \CARRYB[1012][2] , \CARRYB[1012][1] ,
         \CARRYB[1012][0] , \CARRYB[1011][2] , \CARRYB[1011][1] ,
         \CARRYB[1011][0] , \CARRYB[1010][2] , \CARRYB[1010][1] ,
         \CARRYB[1010][0] , \CARRYB[1009][2] , \CARRYB[1009][1] ,
         \CARRYB[1009][0] , \CARRYB[1008][2] , \CARRYB[1008][1] ,
         \CARRYB[1008][0] , \CARRYB[1007][2] , \CARRYB[1007][1] ,
         \CARRYB[1007][0] , \CARRYB[1006][2] , \CARRYB[1006][1] ,
         \CARRYB[1006][0] , \CARRYB[1005][2] , \CARRYB[1005][1] ,
         \CARRYB[1005][0] , \CARRYB[1004][2] , \CARRYB[1004][1] ,
         \CARRYB[1004][0] , \CARRYB[1003][2] , \CARRYB[1003][1] ,
         \CARRYB[1003][0] , \CARRYB[1002][2] , \CARRYB[1002][1] ,
         \CARRYB[1002][0] , \CARRYB[1001][2] , \CARRYB[1001][1] ,
         \CARRYB[1001][0] , \CARRYB[1000][2] , \CARRYB[1000][1] ,
         \CARRYB[1000][0] , \CARRYB[999][2] , \CARRYB[999][1] ,
         \CARRYB[999][0] , \CARRYB[998][2] , \CARRYB[998][1] ,
         \CARRYB[998][0] , \CARRYB[997][2] , \CARRYB[997][1] ,
         \CARRYB[997][0] , \CARRYB[996][2] , \CARRYB[996][1] ,
         \CARRYB[996][0] , \CARRYB[995][2] , \CARRYB[995][1] ,
         \CARRYB[995][0] , \CARRYB[994][2] , \CARRYB[994][1] ,
         \CARRYB[994][0] , \CARRYB[993][2] , \CARRYB[993][1] ,
         \CARRYB[993][0] , \CARRYB[992][2] , \CARRYB[992][1] ,
         \CARRYB[992][0] , \CARRYB[991][2] , \CARRYB[991][1] ,
         \CARRYB[991][0] , \CARRYB[990][2] , \CARRYB[990][1] ,
         \CARRYB[990][0] , \CARRYB[989][2] , \CARRYB[989][1] ,
         \CARRYB[989][0] , \CARRYB[988][2] , \CARRYB[988][1] ,
         \CARRYB[988][0] , \CARRYB[987][2] , \CARRYB[987][1] ,
         \CARRYB[987][0] , \CARRYB[986][2] , \CARRYB[986][1] ,
         \CARRYB[986][0] , \CARRYB[985][2] , \CARRYB[985][1] ,
         \CARRYB[985][0] , \CARRYB[984][2] , \CARRYB[984][1] ,
         \CARRYB[984][0] , \CARRYB[983][2] , \CARRYB[983][1] ,
         \CARRYB[983][0] , \CARRYB[982][2] , \CARRYB[982][1] ,
         \CARRYB[982][0] , \CARRYB[981][2] , \CARRYB[981][1] ,
         \CARRYB[981][0] , \CARRYB[980][2] , \CARRYB[980][1] ,
         \CARRYB[980][0] , \CARRYB[979][2] , \CARRYB[979][1] ,
         \CARRYB[979][0] , \CARRYB[978][2] , \CARRYB[978][1] ,
         \CARRYB[978][0] , \CARRYB[977][2] , \CARRYB[977][1] ,
         \CARRYB[977][0] , \CARRYB[976][2] , \CARRYB[976][1] ,
         \CARRYB[976][0] , \CARRYB[975][2] , \CARRYB[975][1] ,
         \CARRYB[975][0] , \CARRYB[974][2] , \CARRYB[974][1] ,
         \CARRYB[974][0] , \CARRYB[973][2] , \CARRYB[973][1] ,
         \CARRYB[973][0] , \CARRYB[972][2] , \CARRYB[972][1] ,
         \CARRYB[972][0] , \CARRYB[971][2] , \CARRYB[971][1] ,
         \CARRYB[971][0] , \CARRYB[970][2] , \CARRYB[970][1] ,
         \CARRYB[970][0] , \CARRYB[969][2] , \CARRYB[969][1] ,
         \CARRYB[969][0] , \CARRYB[968][2] , \CARRYB[968][1] ,
         \CARRYB[968][0] , \CARRYB[967][2] , \CARRYB[967][1] ,
         \CARRYB[967][0] , \CARRYB[966][2] , \CARRYB[966][1] ,
         \CARRYB[966][0] , \CARRYB[965][2] , \CARRYB[965][1] ,
         \CARRYB[965][0] , \CARRYB[964][2] , \CARRYB[964][1] ,
         \CARRYB[964][0] , \CARRYB[963][2] , \CARRYB[963][1] ,
         \CARRYB[963][0] , \CARRYB[962][2] , \CARRYB[962][1] ,
         \CARRYB[962][0] , \CARRYB[961][2] , \CARRYB[961][1] ,
         \CARRYB[961][0] , \CARRYB[960][2] , \CARRYB[960][1] ,
         \CARRYB[960][0] , \CARRYB[959][2] , \CARRYB[959][1] ,
         \CARRYB[959][0] , \CARRYB[958][2] , \CARRYB[958][1] ,
         \CARRYB[958][0] , \CARRYB[957][2] , \CARRYB[957][1] ,
         \CARRYB[957][0] , \CARRYB[956][2] , \CARRYB[956][1] ,
         \CARRYB[956][0] , \CARRYB[955][2] , \CARRYB[955][1] ,
         \CARRYB[955][0] , \CARRYB[954][2] , \CARRYB[954][1] ,
         \CARRYB[954][0] , \CARRYB[953][2] , \CARRYB[953][1] ,
         \CARRYB[953][0] , \CARRYB[952][2] , \CARRYB[952][1] ,
         \CARRYB[952][0] , \CARRYB[951][2] , \CARRYB[951][1] ,
         \CARRYB[951][0] , \CARRYB[950][2] , \CARRYB[950][1] ,
         \CARRYB[950][0] , \CARRYB[949][2] , \CARRYB[949][1] ,
         \CARRYB[949][0] , \CARRYB[948][2] , \CARRYB[948][1] ,
         \CARRYB[948][0] , \CARRYB[947][2] , \CARRYB[947][1] ,
         \CARRYB[947][0] , \CARRYB[946][2] , \CARRYB[946][1] ,
         \CARRYB[946][0] , \CARRYB[945][2] , \CARRYB[945][1] ,
         \CARRYB[945][0] , \CARRYB[944][2] , \CARRYB[944][1] ,
         \CARRYB[944][0] , \CARRYB[943][2] , \CARRYB[943][1] ,
         \CARRYB[943][0] , \CARRYB[942][2] , \CARRYB[942][1] ,
         \CARRYB[942][0] , \CARRYB[941][2] , \CARRYB[941][1] ,
         \CARRYB[941][0] , \CARRYB[940][2] , \CARRYB[940][1] ,
         \CARRYB[940][0] , \CARRYB[939][2] , \CARRYB[939][1] ,
         \CARRYB[939][0] , \CARRYB[938][2] , \CARRYB[938][1] ,
         \CARRYB[938][0] , \CARRYB[937][2] , \CARRYB[937][1] ,
         \CARRYB[937][0] , \CARRYB[936][2] , \CARRYB[936][1] ,
         \CARRYB[936][0] , \CARRYB[935][2] , \CARRYB[935][1] ,
         \CARRYB[935][0] , \CARRYB[934][2] , \CARRYB[934][1] ,
         \CARRYB[934][0] , \CARRYB[933][2] , \CARRYB[933][1] ,
         \CARRYB[933][0] , \CARRYB[932][2] , \CARRYB[932][1] ,
         \CARRYB[932][0] , \CARRYB[931][2] , \CARRYB[931][1] ,
         \CARRYB[931][0] , \CARRYB[930][2] , \CARRYB[930][1] ,
         \CARRYB[930][0] , \CARRYB[929][2] , \CARRYB[929][1] ,
         \CARRYB[929][0] , \CARRYB[928][2] , \CARRYB[928][1] ,
         \CARRYB[928][0] , \CARRYB[927][2] , \CARRYB[927][1] ,
         \CARRYB[927][0] , \CARRYB[926][2] , \CARRYB[926][1] ,
         \CARRYB[926][0] , \CARRYB[925][2] , \CARRYB[925][1] ,
         \CARRYB[925][0] , \CARRYB[924][2] , \CARRYB[924][1] ,
         \CARRYB[924][0] , \CARRYB[923][2] , \CARRYB[923][1] ,
         \CARRYB[923][0] , \CARRYB[922][2] , \CARRYB[922][1] ,
         \CARRYB[922][0] , \CARRYB[921][2] , \CARRYB[921][1] ,
         \CARRYB[921][0] , \CARRYB[920][2] , \CARRYB[920][1] ,
         \CARRYB[920][0] , \CARRYB[919][2] , \CARRYB[919][1] ,
         \CARRYB[919][0] , \CARRYB[918][2] , \CARRYB[918][1] ,
         \CARRYB[918][0] , \CARRYB[917][2] , \CARRYB[917][1] ,
         \CARRYB[917][0] , \CARRYB[916][2] , \CARRYB[916][1] ,
         \CARRYB[916][0] , \CARRYB[915][2] , \CARRYB[915][1] ,
         \CARRYB[915][0] , \CARRYB[914][2] , \CARRYB[914][1] ,
         \CARRYB[914][0] , \CARRYB[913][2] , \CARRYB[913][1] ,
         \CARRYB[913][0] , \CARRYB[912][2] , \CARRYB[912][1] ,
         \CARRYB[912][0] , \CARRYB[911][2] , \CARRYB[911][1] ,
         \CARRYB[911][0] , \CARRYB[910][2] , \CARRYB[910][1] ,
         \CARRYB[910][0] , \CARRYB[909][2] , \CARRYB[909][1] ,
         \CARRYB[909][0] , \CARRYB[908][2] , \CARRYB[908][1] ,
         \CARRYB[908][0] , \CARRYB[907][2] , \CARRYB[907][1] ,
         \CARRYB[907][0] , \CARRYB[906][2] , \CARRYB[906][1] ,
         \CARRYB[906][0] , \CARRYB[905][2] , \CARRYB[905][1] ,
         \CARRYB[905][0] , \CARRYB[904][2] , \CARRYB[904][1] ,
         \CARRYB[904][0] , \CARRYB[903][2] , \CARRYB[903][1] ,
         \CARRYB[903][0] , \CARRYB[902][2] , \CARRYB[902][1] ,
         \CARRYB[902][0] , \CARRYB[901][2] , \CARRYB[901][1] ,
         \CARRYB[901][0] , \CARRYB[900][2] , \CARRYB[900][1] ,
         \CARRYB[900][0] , \CARRYB[899][2] , \CARRYB[899][1] ,
         \CARRYB[899][0] , \CARRYB[898][2] , \CARRYB[898][1] ,
         \CARRYB[898][0] , \CARRYB[897][2] , \CARRYB[897][1] ,
         \CARRYB[897][0] , \CARRYB[896][2] , \CARRYB[896][1] ,
         \CARRYB[896][0] , \SUMB[1022][1] , \SUMB[1021][2] , \SUMB[1021][1] ,
         \SUMB[1020][2] , \SUMB[1020][1] , \SUMB[1019][2] , \SUMB[1019][1] ,
         \SUMB[1018][2] , \SUMB[1018][1] , \SUMB[1017][2] , \SUMB[1017][1] ,
         \SUMB[1016][2] , \SUMB[1016][1] , \SUMB[1015][2] , \SUMB[1015][1] ,
         \SUMB[1014][2] , \SUMB[1014][1] , \SUMB[1013][2] , \SUMB[1013][1] ,
         \SUMB[1012][2] , \SUMB[1012][1] , \SUMB[1011][2] , \SUMB[1011][1] ,
         \SUMB[1010][2] , \SUMB[1010][1] , \SUMB[1009][2] , \SUMB[1009][1] ,
         \SUMB[1008][2] , \SUMB[1008][1] , \SUMB[1007][2] , \SUMB[1007][1] ,
         \SUMB[1006][2] , \SUMB[1006][1] , \SUMB[1005][2] , \SUMB[1005][1] ,
         \SUMB[1004][2] , \SUMB[1004][1] , \SUMB[1003][2] , \SUMB[1003][1] ,
         \SUMB[1002][2] , \SUMB[1002][1] , \SUMB[1001][2] , \SUMB[1001][1] ,
         \SUMB[1000][2] , \SUMB[1000][1] , \SUMB[999][2] , \SUMB[999][1] ,
         \SUMB[998][2] , \SUMB[998][1] , \SUMB[997][2] , \SUMB[997][1] ,
         \SUMB[996][2] , \SUMB[996][1] , \SUMB[995][2] , \SUMB[995][1] ,
         \SUMB[994][2] , \SUMB[994][1] , \SUMB[993][2] , \SUMB[993][1] ,
         \SUMB[992][2] , \SUMB[992][1] , \SUMB[991][2] , \SUMB[991][1] ,
         \SUMB[990][2] , \SUMB[990][1] , \SUMB[989][2] , \SUMB[989][1] ,
         \SUMB[988][2] , \SUMB[988][1] , \SUMB[987][2] , \SUMB[987][1] ,
         \SUMB[986][2] , \SUMB[986][1] , \SUMB[985][2] , \SUMB[985][1] ,
         \SUMB[984][2] , \SUMB[984][1] , \SUMB[983][2] , \SUMB[983][1] ,
         \SUMB[982][2] , \SUMB[982][1] , \SUMB[981][2] , \SUMB[981][1] ,
         \SUMB[980][2] , \SUMB[980][1] , \SUMB[979][2] , \SUMB[979][1] ,
         \SUMB[978][2] , \SUMB[978][1] , \SUMB[977][2] , \SUMB[977][1] ,
         \SUMB[976][2] , \SUMB[976][1] , \SUMB[975][2] , \SUMB[975][1] ,
         \SUMB[974][2] , \SUMB[974][1] , \SUMB[973][2] , \SUMB[973][1] ,
         \SUMB[972][2] , \SUMB[972][1] , \SUMB[971][2] , \SUMB[971][1] ,
         \SUMB[970][2] , \SUMB[970][1] , \SUMB[969][2] , \SUMB[969][1] ,
         \SUMB[968][2] , \SUMB[968][1] , \SUMB[967][2] , \SUMB[967][1] ,
         \SUMB[966][2] , \SUMB[966][1] , \SUMB[965][2] , \SUMB[965][1] ,
         \SUMB[964][2] , \SUMB[964][1] , \SUMB[963][2] , \SUMB[963][1] ,
         \SUMB[962][2] , \SUMB[962][1] , \SUMB[961][2] , \SUMB[961][1] ,
         \SUMB[960][2] , \SUMB[960][1] , \SUMB[959][2] , \SUMB[959][1] ,
         \SUMB[958][2] , \SUMB[958][1] , \SUMB[957][2] , \SUMB[957][1] ,
         \SUMB[956][2] , \SUMB[956][1] , \SUMB[955][2] , \SUMB[955][1] ,
         \SUMB[954][2] , \SUMB[954][1] , \SUMB[953][2] , \SUMB[953][1] ,
         \SUMB[952][2] , \SUMB[952][1] , \SUMB[951][2] , \SUMB[951][1] ,
         \SUMB[950][2] , \SUMB[950][1] , \SUMB[949][2] , \SUMB[949][1] ,
         \SUMB[948][2] , \SUMB[948][1] , \SUMB[947][2] , \SUMB[947][1] ,
         \SUMB[946][2] , \SUMB[946][1] , \SUMB[945][2] , \SUMB[945][1] ,
         \SUMB[944][2] , \SUMB[944][1] , \SUMB[943][2] , \SUMB[943][1] ,
         \SUMB[942][2] , \SUMB[942][1] , \SUMB[941][2] , \SUMB[941][1] ,
         \SUMB[940][2] , \SUMB[940][1] , \SUMB[939][2] , \SUMB[939][1] ,
         \SUMB[938][2] , \SUMB[938][1] , \SUMB[937][2] , \SUMB[937][1] ,
         \SUMB[936][2] , \SUMB[936][1] , \SUMB[935][2] , \SUMB[935][1] ,
         \SUMB[934][2] , \SUMB[934][1] , \SUMB[933][2] , \SUMB[933][1] ,
         \SUMB[932][2] , \SUMB[932][1] , \SUMB[931][2] , \SUMB[931][1] ,
         \SUMB[930][2] , \SUMB[930][1] , \SUMB[929][2] , \SUMB[929][1] ,
         \SUMB[928][2] , \SUMB[928][1] , \SUMB[927][2] , \SUMB[927][1] ,
         \SUMB[926][2] , \SUMB[926][1] , \SUMB[925][2] , \SUMB[925][1] ,
         \SUMB[924][2] , \SUMB[924][1] , \SUMB[923][2] , \SUMB[923][1] ,
         \SUMB[922][2] , \SUMB[922][1] , \SUMB[921][2] , \SUMB[921][1] ,
         \SUMB[920][2] , \SUMB[920][1] , \SUMB[919][2] , \SUMB[919][1] ,
         \SUMB[918][2] , \SUMB[918][1] , \SUMB[917][2] , \SUMB[917][1] ,
         \SUMB[916][2] , \SUMB[916][1] , \SUMB[915][2] , \SUMB[915][1] ,
         \SUMB[914][2] , \SUMB[914][1] , \SUMB[913][2] , \SUMB[913][1] ,
         \SUMB[912][2] , \SUMB[912][1] , \SUMB[911][2] , \SUMB[911][1] ,
         \SUMB[910][2] , \SUMB[910][1] , \SUMB[909][2] , \SUMB[909][1] ,
         \SUMB[908][2] , \SUMB[908][1] , \SUMB[907][2] , \SUMB[907][1] ,
         \SUMB[906][2] , \SUMB[906][1] , \SUMB[905][2] , \SUMB[905][1] ,
         \SUMB[904][2] , \SUMB[904][1] , \SUMB[903][2] , \SUMB[903][1] ,
         \SUMB[902][2] , \SUMB[902][1] , \SUMB[901][2] , \SUMB[901][1] ,
         \SUMB[900][2] , \SUMB[900][1] , \SUMB[899][2] , \SUMB[899][1] ,
         \SUMB[898][2] , \SUMB[898][1] , \SUMB[897][2] , \SUMB[897][1] ,
         \SUMB[896][2] , \SUMB[896][1] ;

  FADDER S4_0 ( .CIN(\ab[1023][0] ), .IN0(\CARRYB[1022][0] ), .IN1(
        \SUMB[1022][1] ), .SUM(PRODUCT[1023]) );
  FADDER S1_1022_0 ( .CIN(\ab[1022][0] ), .IN0(\CARRYB[1021][0] ), .IN1(
        \SUMB[1021][1] ), .COUT(\CARRYB[1022][0] ), .SUM(PRODUCT[1022]) );
  FADDER S2_1022_1 ( .CIN(\ab[1022][1] ), .IN0(\CARRYB[1021][1] ), .IN1(
        \SUMB[1021][2] ), .SUM(\SUMB[1022][1] ) );
  FADDER S1_1021_0 ( .CIN(\ab[1021][0] ), .IN0(\CARRYB[1020][0] ), .IN1(
        \SUMB[1020][1] ), .COUT(\CARRYB[1021][0] ), .SUM(PRODUCT[1021]) );
  FADDER S2_1021_1 ( .CIN(\ab[1021][1] ), .IN0(\CARRYB[1020][1] ), .IN1(
        \SUMB[1020][2] ), .COUT(\CARRYB[1021][1] ), .SUM(\SUMB[1021][1] ) );
  FADDER S3_1021_2 ( .CIN(\ab[1021][2] ), .IN0(\CARRYB[1020][2] ), .IN1(
        \ab[1020][3] ), .SUM(\SUMB[1021][2] ) );
  FADDER S1_1020_0 ( .CIN(\ab[1020][0] ), .IN0(\CARRYB[1019][0] ), .IN1(
        \SUMB[1019][1] ), .COUT(\CARRYB[1020][0] ), .SUM(PRODUCT[1020]) );
  FADDER S2_1020_1 ( .CIN(\ab[1020][1] ), .IN0(\CARRYB[1019][1] ), .IN1(
        \SUMB[1019][2] ), .COUT(\CARRYB[1020][1] ), .SUM(\SUMB[1020][1] ) );
  FADDER S3_1020_2 ( .CIN(\ab[1020][2] ), .IN0(\CARRYB[1019][2] ), .IN1(
        \ab[1019][3] ), .COUT(\CARRYB[1020][2] ), .SUM(\SUMB[1020][2] ) );
  FADDER S1_1019_0 ( .CIN(\ab[1019][0] ), .IN0(\CARRYB[1018][0] ), .IN1(
        \SUMB[1018][1] ), .COUT(\CARRYB[1019][0] ), .SUM(PRODUCT[1019]) );
  FADDER S2_1019_1 ( .CIN(\ab[1019][1] ), .IN0(\CARRYB[1018][1] ), .IN1(
        \SUMB[1018][2] ), .COUT(\CARRYB[1019][1] ), .SUM(\SUMB[1019][1] ) );
  FADDER S3_1019_2 ( .CIN(\ab[1019][2] ), .IN0(\CARRYB[1018][2] ), .IN1(
        \ab[1018][3] ), .COUT(\CARRYB[1019][2] ), .SUM(\SUMB[1019][2] ) );
  FADDER S1_1018_0 ( .CIN(\ab[1018][0] ), .IN0(\CARRYB[1017][0] ), .IN1(
        \SUMB[1017][1] ), .COUT(\CARRYB[1018][0] ), .SUM(PRODUCT[1018]) );
  FADDER S2_1018_1 ( .CIN(\ab[1018][1] ), .IN0(\CARRYB[1017][1] ), .IN1(
        \SUMB[1017][2] ), .COUT(\CARRYB[1018][1] ), .SUM(\SUMB[1018][1] ) );
  FADDER S3_1018_2 ( .CIN(\ab[1018][2] ), .IN0(\CARRYB[1017][2] ), .IN1(
        \ab[1017][3] ), .COUT(\CARRYB[1018][2] ), .SUM(\SUMB[1018][2] ) );
  FADDER S1_1017_0 ( .CIN(\ab[1017][0] ), .IN0(\CARRYB[1016][0] ), .IN1(
        \SUMB[1016][1] ), .COUT(\CARRYB[1017][0] ), .SUM(PRODUCT[1017]) );
  FADDER S2_1017_1 ( .CIN(\ab[1017][1] ), .IN0(\CARRYB[1016][1] ), .IN1(
        \SUMB[1016][2] ), .COUT(\CARRYB[1017][1] ), .SUM(\SUMB[1017][1] ) );
  FADDER S3_1017_2 ( .CIN(\ab[1017][2] ), .IN0(\CARRYB[1016][2] ), .IN1(
        \ab[1016][3] ), .COUT(\CARRYB[1017][2] ), .SUM(\SUMB[1017][2] ) );
  FADDER S1_1016_0 ( .CIN(\ab[1016][0] ), .IN0(\CARRYB[1015][0] ), .IN1(
        \SUMB[1015][1] ), .COUT(\CARRYB[1016][0] ), .SUM(PRODUCT[1016]) );
  FADDER S2_1016_1 ( .CIN(\ab[1016][1] ), .IN0(\CARRYB[1015][1] ), .IN1(
        \SUMB[1015][2] ), .COUT(\CARRYB[1016][1] ), .SUM(\SUMB[1016][1] ) );
  FADDER S3_1016_2 ( .CIN(\ab[1016][2] ), .IN0(\CARRYB[1015][2] ), .IN1(
        \ab[1015][3] ), .COUT(\CARRYB[1016][2] ), .SUM(\SUMB[1016][2] ) );
  FADDER S1_1015_0 ( .CIN(\ab[1015][0] ), .IN0(\CARRYB[1014][0] ), .IN1(
        \SUMB[1014][1] ), .COUT(\CARRYB[1015][0] ), .SUM(PRODUCT[1015]) );
  FADDER S2_1015_1 ( .CIN(\ab[1015][1] ), .IN0(\CARRYB[1014][1] ), .IN1(
        \SUMB[1014][2] ), .COUT(\CARRYB[1015][1] ), .SUM(\SUMB[1015][1] ) );
  FADDER S3_1015_2 ( .CIN(\ab[1015][2] ), .IN0(\CARRYB[1014][2] ), .IN1(
        \ab[1014][3] ), .COUT(\CARRYB[1015][2] ), .SUM(\SUMB[1015][2] ) );
  FADDER S1_1014_0 ( .CIN(\ab[1014][0] ), .IN0(\CARRYB[1013][0] ), .IN1(
        \SUMB[1013][1] ), .COUT(\CARRYB[1014][0] ), .SUM(PRODUCT[1014]) );
  FADDER S2_1014_1 ( .CIN(\ab[1014][1] ), .IN0(\CARRYB[1013][1] ), .IN1(
        \SUMB[1013][2] ), .COUT(\CARRYB[1014][1] ), .SUM(\SUMB[1014][1] ) );
  FADDER S3_1014_2 ( .CIN(\ab[1014][2] ), .IN0(\CARRYB[1013][2] ), .IN1(
        \ab[1013][3] ), .COUT(\CARRYB[1014][2] ), .SUM(\SUMB[1014][2] ) );
  FADDER S1_1013_0 ( .CIN(\ab[1013][0] ), .IN0(\CARRYB[1012][0] ), .IN1(
        \SUMB[1012][1] ), .COUT(\CARRYB[1013][0] ), .SUM(PRODUCT[1013]) );
  FADDER S2_1013_1 ( .CIN(\ab[1013][1] ), .IN0(\CARRYB[1012][1] ), .IN1(
        \SUMB[1012][2] ), .COUT(\CARRYB[1013][1] ), .SUM(\SUMB[1013][1] ) );
  FADDER S3_1013_2 ( .CIN(\ab[1013][2] ), .IN0(\CARRYB[1012][2] ), .IN1(
        \ab[1012][3] ), .COUT(\CARRYB[1013][2] ), .SUM(\SUMB[1013][2] ) );
  FADDER S1_1012_0 ( .CIN(\ab[1012][0] ), .IN0(\CARRYB[1011][0] ), .IN1(
        \SUMB[1011][1] ), .COUT(\CARRYB[1012][0] ), .SUM(PRODUCT[1012]) );
  FADDER S2_1012_1 ( .CIN(\ab[1012][1] ), .IN0(\CARRYB[1011][1] ), .IN1(
        \SUMB[1011][2] ), .COUT(\CARRYB[1012][1] ), .SUM(\SUMB[1012][1] ) );
  FADDER S3_1012_2 ( .CIN(\ab[1012][2] ), .IN0(\CARRYB[1011][2] ), .IN1(
        \ab[1011][3] ), .COUT(\CARRYB[1012][2] ), .SUM(\SUMB[1012][2] ) );
  FADDER S1_1011_0 ( .CIN(\ab[1011][0] ), .IN0(\CARRYB[1010][0] ), .IN1(
        \SUMB[1010][1] ), .COUT(\CARRYB[1011][0] ), .SUM(PRODUCT[1011]) );
  FADDER S2_1011_1 ( .CIN(\ab[1011][1] ), .IN0(\CARRYB[1010][1] ), .IN1(
        \SUMB[1010][2] ), .COUT(\CARRYB[1011][1] ), .SUM(\SUMB[1011][1] ) );
  FADDER S3_1011_2 ( .CIN(\ab[1011][2] ), .IN0(\CARRYB[1010][2] ), .IN1(
        \ab[1010][3] ), .COUT(\CARRYB[1011][2] ), .SUM(\SUMB[1011][2] ) );
  FADDER S1_1010_0 ( .CIN(\ab[1010][0] ), .IN0(\CARRYB[1009][0] ), .IN1(
        \SUMB[1009][1] ), .COUT(\CARRYB[1010][0] ), .SUM(PRODUCT[1010]) );
  FADDER S2_1010_1 ( .CIN(\ab[1010][1] ), .IN0(\CARRYB[1009][1] ), .IN1(
        \SUMB[1009][2] ), .COUT(\CARRYB[1010][1] ), .SUM(\SUMB[1010][1] ) );
  FADDER S3_1010_2 ( .CIN(\ab[1010][2] ), .IN0(\CARRYB[1009][2] ), .IN1(
        \ab[1009][3] ), .COUT(\CARRYB[1010][2] ), .SUM(\SUMB[1010][2] ) );
  FADDER S1_1009_0 ( .CIN(\ab[1009][0] ), .IN0(\CARRYB[1008][0] ), .IN1(
        \SUMB[1008][1] ), .COUT(\CARRYB[1009][0] ), .SUM(PRODUCT[1009]) );
  FADDER S2_1009_1 ( .CIN(\ab[1009][1] ), .IN0(\CARRYB[1008][1] ), .IN1(
        \SUMB[1008][2] ), .COUT(\CARRYB[1009][1] ), .SUM(\SUMB[1009][1] ) );
  FADDER S3_1009_2 ( .CIN(\ab[1009][2] ), .IN0(\CARRYB[1008][2] ), .IN1(
        \ab[1008][3] ), .COUT(\CARRYB[1009][2] ), .SUM(\SUMB[1009][2] ) );
  FADDER S1_1008_0 ( .CIN(\ab[1008][0] ), .IN0(\CARRYB[1007][0] ), .IN1(
        \SUMB[1007][1] ), .COUT(\CARRYB[1008][0] ), .SUM(PRODUCT[1008]) );
  FADDER S2_1008_1 ( .CIN(\ab[1008][1] ), .IN0(\CARRYB[1007][1] ), .IN1(
        \SUMB[1007][2] ), .COUT(\CARRYB[1008][1] ), .SUM(\SUMB[1008][1] ) );
  FADDER S3_1008_2 ( .CIN(\ab[1008][2] ), .IN0(\CARRYB[1007][2] ), .IN1(
        \ab[1007][3] ), .COUT(\CARRYB[1008][2] ), .SUM(\SUMB[1008][2] ) );
  FADDER S1_1007_0 ( .CIN(\ab[1007][0] ), .IN0(\CARRYB[1006][0] ), .IN1(
        \SUMB[1006][1] ), .COUT(\CARRYB[1007][0] ), .SUM(PRODUCT[1007]) );
  FADDER S2_1007_1 ( .CIN(\ab[1007][1] ), .IN0(\CARRYB[1006][1] ), .IN1(
        \SUMB[1006][2] ), .COUT(\CARRYB[1007][1] ), .SUM(\SUMB[1007][1] ) );
  FADDER S3_1007_2 ( .CIN(\ab[1007][2] ), .IN0(\CARRYB[1006][2] ), .IN1(
        \ab[1006][3] ), .COUT(\CARRYB[1007][2] ), .SUM(\SUMB[1007][2] ) );
  FADDER S1_1006_0 ( .CIN(\ab[1006][0] ), .IN0(\CARRYB[1005][0] ), .IN1(
        \SUMB[1005][1] ), .COUT(\CARRYB[1006][0] ), .SUM(PRODUCT[1006]) );
  FADDER S2_1006_1 ( .CIN(\ab[1006][1] ), .IN0(\CARRYB[1005][1] ), .IN1(
        \SUMB[1005][2] ), .COUT(\CARRYB[1006][1] ), .SUM(\SUMB[1006][1] ) );
  FADDER S3_1006_2 ( .CIN(\ab[1006][2] ), .IN0(\CARRYB[1005][2] ), .IN1(
        \ab[1005][3] ), .COUT(\CARRYB[1006][2] ), .SUM(\SUMB[1006][2] ) );
  FADDER S1_1005_0 ( .CIN(\ab[1005][0] ), .IN0(\CARRYB[1004][0] ), .IN1(
        \SUMB[1004][1] ), .COUT(\CARRYB[1005][0] ), .SUM(PRODUCT[1005]) );
  FADDER S2_1005_1 ( .CIN(\ab[1005][1] ), .IN0(\CARRYB[1004][1] ), .IN1(
        \SUMB[1004][2] ), .COUT(\CARRYB[1005][1] ), .SUM(\SUMB[1005][1] ) );
  FADDER S3_1005_2 ( .CIN(\ab[1005][2] ), .IN0(\CARRYB[1004][2] ), .IN1(
        \ab[1004][3] ), .COUT(\CARRYB[1005][2] ), .SUM(\SUMB[1005][2] ) );
  FADDER S1_1004_0 ( .CIN(\ab[1004][0] ), .IN0(\CARRYB[1003][0] ), .IN1(
        \SUMB[1003][1] ), .COUT(\CARRYB[1004][0] ), .SUM(PRODUCT[1004]) );
  FADDER S2_1004_1 ( .CIN(\ab[1004][1] ), .IN0(\CARRYB[1003][1] ), .IN1(
        \SUMB[1003][2] ), .COUT(\CARRYB[1004][1] ), .SUM(\SUMB[1004][1] ) );
  FADDER S3_1004_2 ( .CIN(\ab[1004][2] ), .IN0(\CARRYB[1003][2] ), .IN1(
        \ab[1003][3] ), .COUT(\CARRYB[1004][2] ), .SUM(\SUMB[1004][2] ) );
  FADDER S1_1003_0 ( .CIN(\ab[1003][0] ), .IN0(\CARRYB[1002][0] ), .IN1(
        \SUMB[1002][1] ), .COUT(\CARRYB[1003][0] ), .SUM(PRODUCT[1003]) );
  FADDER S2_1003_1 ( .CIN(\ab[1003][1] ), .IN0(\CARRYB[1002][1] ), .IN1(
        \SUMB[1002][2] ), .COUT(\CARRYB[1003][1] ), .SUM(\SUMB[1003][1] ) );
  FADDER S3_1003_2 ( .CIN(\ab[1003][2] ), .IN0(\CARRYB[1002][2] ), .IN1(
        \ab[1002][3] ), .COUT(\CARRYB[1003][2] ), .SUM(\SUMB[1003][2] ) );
  FADDER S1_1002_0 ( .CIN(\ab[1002][0] ), .IN0(\CARRYB[1001][0] ), .IN1(
        \SUMB[1001][1] ), .COUT(\CARRYB[1002][0] ), .SUM(PRODUCT[1002]) );
  FADDER S2_1002_1 ( .CIN(\ab[1002][1] ), .IN0(\CARRYB[1001][1] ), .IN1(
        \SUMB[1001][2] ), .COUT(\CARRYB[1002][1] ), .SUM(\SUMB[1002][1] ) );
  FADDER S3_1002_2 ( .CIN(\ab[1002][2] ), .IN0(\CARRYB[1001][2] ), .IN1(
        \ab[1001][3] ), .COUT(\CARRYB[1002][2] ), .SUM(\SUMB[1002][2] ) );
  FADDER S1_1001_0 ( .CIN(\ab[1001][0] ), .IN0(\CARRYB[1000][0] ), .IN1(
        \SUMB[1000][1] ), .COUT(\CARRYB[1001][0] ), .SUM(PRODUCT[1001]) );
  FADDER S2_1001_1 ( .CIN(\ab[1001][1] ), .IN0(\CARRYB[1000][1] ), .IN1(
        \SUMB[1000][2] ), .COUT(\CARRYB[1001][1] ), .SUM(\SUMB[1001][1] ) );
  FADDER S3_1001_2 ( .CIN(\ab[1001][2] ), .IN0(\CARRYB[1000][2] ), .IN1(
        \ab[1000][3] ), .COUT(\CARRYB[1001][2] ), .SUM(\SUMB[1001][2] ) );
  FADDER S1_1000_0 ( .CIN(\ab[1000][0] ), .IN0(\CARRYB[999][0] ), .IN1(
        \SUMB[999][1] ), .COUT(\CARRYB[1000][0] ), .SUM(PRODUCT[1000]) );
  FADDER S2_1000_1 ( .CIN(\ab[1000][1] ), .IN0(\CARRYB[999][1] ), .IN1(
        \SUMB[999][2] ), .COUT(\CARRYB[1000][1] ), .SUM(\SUMB[1000][1] ) );
  FADDER S3_1000_2 ( .CIN(\ab[1000][2] ), .IN0(\CARRYB[999][2] ), .IN1(
        \ab[999][3] ), .COUT(\CARRYB[1000][2] ), .SUM(\SUMB[1000][2] ) );
  FADDER S1_999_0 ( .CIN(\ab[999][0] ), .IN0(\CARRYB[998][0] ), .IN1(
        \SUMB[998][1] ), .COUT(\CARRYB[999][0] ), .SUM(PRODUCT[999]) );
  FADDER S2_999_1 ( .CIN(\ab[999][1] ), .IN0(\CARRYB[998][1] ), .IN1(
        \SUMB[998][2] ), .COUT(\CARRYB[999][1] ), .SUM(\SUMB[999][1] ) );
  FADDER S3_999_2 ( .CIN(\ab[999][2] ), .IN0(\CARRYB[998][2] ), .IN1(
        \ab[998][3] ), .COUT(\CARRYB[999][2] ), .SUM(\SUMB[999][2] ) );
  FADDER S1_998_0 ( .CIN(\ab[998][0] ), .IN0(\CARRYB[997][0] ), .IN1(
        \SUMB[997][1] ), .COUT(\CARRYB[998][0] ), .SUM(PRODUCT[998]) );
  FADDER S2_998_1 ( .CIN(\ab[998][1] ), .IN0(\CARRYB[997][1] ), .IN1(
        \SUMB[997][2] ), .COUT(\CARRYB[998][1] ), .SUM(\SUMB[998][1] ) );
  FADDER S3_998_2 ( .CIN(\ab[998][2] ), .IN0(\CARRYB[997][2] ), .IN1(
        \ab[997][3] ), .COUT(\CARRYB[998][2] ), .SUM(\SUMB[998][2] ) );
  FADDER S1_997_0 ( .CIN(\ab[997][0] ), .IN0(\CARRYB[996][0] ), .IN1(
        \SUMB[996][1] ), .COUT(\CARRYB[997][0] ), .SUM(PRODUCT[997]) );
  FADDER S2_997_1 ( .CIN(\ab[997][1] ), .IN0(\CARRYB[996][1] ), .IN1(
        \SUMB[996][2] ), .COUT(\CARRYB[997][1] ), .SUM(\SUMB[997][1] ) );
  FADDER S3_997_2 ( .CIN(\ab[997][2] ), .IN0(\CARRYB[996][2] ), .IN1(
        \ab[996][3] ), .COUT(\CARRYB[997][2] ), .SUM(\SUMB[997][2] ) );
  FADDER S1_996_0 ( .CIN(\ab[996][0] ), .IN0(\CARRYB[995][0] ), .IN1(
        \SUMB[995][1] ), .COUT(\CARRYB[996][0] ), .SUM(PRODUCT[996]) );
  FADDER S2_996_1 ( .CIN(\ab[996][1] ), .IN0(\CARRYB[995][1] ), .IN1(
        \SUMB[995][2] ), .COUT(\CARRYB[996][1] ), .SUM(\SUMB[996][1] ) );
  FADDER S3_996_2 ( .CIN(\ab[996][2] ), .IN0(\CARRYB[995][2] ), .IN1(
        \ab[995][3] ), .COUT(\CARRYB[996][2] ), .SUM(\SUMB[996][2] ) );
  FADDER S1_995_0 ( .CIN(\ab[995][0] ), .IN0(\CARRYB[994][0] ), .IN1(
        \SUMB[994][1] ), .COUT(\CARRYB[995][0] ), .SUM(PRODUCT[995]) );
  FADDER S2_995_1 ( .CIN(\ab[995][1] ), .IN0(\CARRYB[994][1] ), .IN1(
        \SUMB[994][2] ), .COUT(\CARRYB[995][1] ), .SUM(\SUMB[995][1] ) );
  FADDER S3_995_2 ( .CIN(\ab[995][2] ), .IN0(\CARRYB[994][2] ), .IN1(
        \ab[994][3] ), .COUT(\CARRYB[995][2] ), .SUM(\SUMB[995][2] ) );
  FADDER S1_994_0 ( .CIN(\ab[994][0] ), .IN0(\CARRYB[993][0] ), .IN1(
        \SUMB[993][1] ), .COUT(\CARRYB[994][0] ), .SUM(PRODUCT[994]) );
  FADDER S2_994_1 ( .CIN(\ab[994][1] ), .IN0(\CARRYB[993][1] ), .IN1(
        \SUMB[993][2] ), .COUT(\CARRYB[994][1] ), .SUM(\SUMB[994][1] ) );
  FADDER S3_994_2 ( .CIN(\ab[994][2] ), .IN0(\CARRYB[993][2] ), .IN1(
        \ab[993][3] ), .COUT(\CARRYB[994][2] ), .SUM(\SUMB[994][2] ) );
  FADDER S1_993_0 ( .CIN(\ab[993][0] ), .IN0(\CARRYB[992][0] ), .IN1(
        \SUMB[992][1] ), .COUT(\CARRYB[993][0] ), .SUM(PRODUCT[993]) );
  FADDER S2_993_1 ( .CIN(\ab[993][1] ), .IN0(\CARRYB[992][1] ), .IN1(
        \SUMB[992][2] ), .COUT(\CARRYB[993][1] ), .SUM(\SUMB[993][1] ) );
  FADDER S3_993_2 ( .CIN(\ab[993][2] ), .IN0(\CARRYB[992][2] ), .IN1(
        \ab[992][3] ), .COUT(\CARRYB[993][2] ), .SUM(\SUMB[993][2] ) );
  FADDER S1_992_0 ( .CIN(\ab[992][0] ), .IN0(\CARRYB[991][0] ), .IN1(
        \SUMB[991][1] ), .COUT(\CARRYB[992][0] ), .SUM(PRODUCT[992]) );
  FADDER S2_992_1 ( .CIN(\ab[992][1] ), .IN0(\CARRYB[991][1] ), .IN1(
        \SUMB[991][2] ), .COUT(\CARRYB[992][1] ), .SUM(\SUMB[992][1] ) );
  FADDER S3_992_2 ( .CIN(\ab[992][2] ), .IN0(\CARRYB[991][2] ), .IN1(
        \ab[991][3] ), .COUT(\CARRYB[992][2] ), .SUM(\SUMB[992][2] ) );
  FADDER S1_991_0 ( .CIN(\ab[991][0] ), .IN0(\CARRYB[990][0] ), .IN1(
        \SUMB[990][1] ), .COUT(\CARRYB[991][0] ), .SUM(PRODUCT[991]) );
  FADDER S2_991_1 ( .CIN(\ab[991][1] ), .IN0(\CARRYB[990][1] ), .IN1(
        \SUMB[990][2] ), .COUT(\CARRYB[991][1] ), .SUM(\SUMB[991][1] ) );
  FADDER S3_991_2 ( .CIN(\ab[991][2] ), .IN0(\CARRYB[990][2] ), .IN1(
        \ab[990][3] ), .COUT(\CARRYB[991][2] ), .SUM(\SUMB[991][2] ) );
  FADDER S1_990_0 ( .CIN(\ab[990][0] ), .IN0(\CARRYB[989][0] ), .IN1(
        \SUMB[989][1] ), .COUT(\CARRYB[990][0] ), .SUM(PRODUCT[990]) );
  FADDER S2_990_1 ( .CIN(\ab[990][1] ), .IN0(\CARRYB[989][1] ), .IN1(
        \SUMB[989][2] ), .COUT(\CARRYB[990][1] ), .SUM(\SUMB[990][1] ) );
  FADDER S3_990_2 ( .CIN(\ab[990][2] ), .IN0(\CARRYB[989][2] ), .IN1(
        \ab[989][3] ), .COUT(\CARRYB[990][2] ), .SUM(\SUMB[990][2] ) );
  FADDER S1_989_0 ( .CIN(\ab[989][0] ), .IN0(\CARRYB[988][0] ), .IN1(
        \SUMB[988][1] ), .COUT(\CARRYB[989][0] ), .SUM(PRODUCT[989]) );
  FADDER S2_989_1 ( .CIN(\ab[989][1] ), .IN0(\CARRYB[988][1] ), .IN1(
        \SUMB[988][2] ), .COUT(\CARRYB[989][1] ), .SUM(\SUMB[989][1] ) );
  FADDER S3_989_2 ( .CIN(\ab[989][2] ), .IN0(\CARRYB[988][2] ), .IN1(
        \ab[988][3] ), .COUT(\CARRYB[989][2] ), .SUM(\SUMB[989][2] ) );
  FADDER S1_988_0 ( .CIN(\ab[988][0] ), .IN0(\CARRYB[987][0] ), .IN1(
        \SUMB[987][1] ), .COUT(\CARRYB[988][0] ), .SUM(PRODUCT[988]) );
  FADDER S2_988_1 ( .CIN(\ab[988][1] ), .IN0(\CARRYB[987][1] ), .IN1(
        \SUMB[987][2] ), .COUT(\CARRYB[988][1] ), .SUM(\SUMB[988][1] ) );
  FADDER S3_988_2 ( .CIN(\ab[988][2] ), .IN0(\CARRYB[987][2] ), .IN1(
        \ab[987][3] ), .COUT(\CARRYB[988][2] ), .SUM(\SUMB[988][2] ) );
  FADDER S1_987_0 ( .CIN(\ab[987][0] ), .IN0(\CARRYB[986][0] ), .IN1(
        \SUMB[986][1] ), .COUT(\CARRYB[987][0] ), .SUM(PRODUCT[987]) );
  FADDER S2_987_1 ( .CIN(\ab[987][1] ), .IN0(\CARRYB[986][1] ), .IN1(
        \SUMB[986][2] ), .COUT(\CARRYB[987][1] ), .SUM(\SUMB[987][1] ) );
  FADDER S3_987_2 ( .CIN(\ab[987][2] ), .IN0(\CARRYB[986][2] ), .IN1(
        \ab[986][3] ), .COUT(\CARRYB[987][2] ), .SUM(\SUMB[987][2] ) );
  FADDER S1_986_0 ( .CIN(\ab[986][0] ), .IN0(\CARRYB[985][0] ), .IN1(
        \SUMB[985][1] ), .COUT(\CARRYB[986][0] ), .SUM(PRODUCT[986]) );
  FADDER S2_986_1 ( .CIN(\ab[986][1] ), .IN0(\CARRYB[985][1] ), .IN1(
        \SUMB[985][2] ), .COUT(\CARRYB[986][1] ), .SUM(\SUMB[986][1] ) );
  FADDER S3_986_2 ( .CIN(\ab[986][2] ), .IN0(\CARRYB[985][2] ), .IN1(
        \ab[985][3] ), .COUT(\CARRYB[986][2] ), .SUM(\SUMB[986][2] ) );
  FADDER S1_985_0 ( .CIN(\ab[985][0] ), .IN0(\CARRYB[984][0] ), .IN1(
        \SUMB[984][1] ), .COUT(\CARRYB[985][0] ), .SUM(PRODUCT[985]) );
  FADDER S2_985_1 ( .CIN(\ab[985][1] ), .IN0(\CARRYB[984][1] ), .IN1(
        \SUMB[984][2] ), .COUT(\CARRYB[985][1] ), .SUM(\SUMB[985][1] ) );
  FADDER S3_985_2 ( .CIN(\ab[985][2] ), .IN0(\CARRYB[984][2] ), .IN1(
        \ab[984][3] ), .COUT(\CARRYB[985][2] ), .SUM(\SUMB[985][2] ) );
  FADDER S1_984_0 ( .CIN(\ab[984][0] ), .IN0(\CARRYB[983][0] ), .IN1(
        \SUMB[983][1] ), .COUT(\CARRYB[984][0] ), .SUM(PRODUCT[984]) );
  FADDER S2_984_1 ( .CIN(\ab[984][1] ), .IN0(\CARRYB[983][1] ), .IN1(
        \SUMB[983][2] ), .COUT(\CARRYB[984][1] ), .SUM(\SUMB[984][1] ) );
  FADDER S3_984_2 ( .CIN(\ab[984][2] ), .IN0(\CARRYB[983][2] ), .IN1(
        \ab[983][3] ), .COUT(\CARRYB[984][2] ), .SUM(\SUMB[984][2] ) );
  FADDER S1_983_0 ( .CIN(\ab[983][0] ), .IN0(\CARRYB[982][0] ), .IN1(
        \SUMB[982][1] ), .COUT(\CARRYB[983][0] ), .SUM(PRODUCT[983]) );
  FADDER S2_983_1 ( .CIN(\ab[983][1] ), .IN0(\CARRYB[982][1] ), .IN1(
        \SUMB[982][2] ), .COUT(\CARRYB[983][1] ), .SUM(\SUMB[983][1] ) );
  FADDER S3_983_2 ( .CIN(\ab[983][2] ), .IN0(\CARRYB[982][2] ), .IN1(
        \ab[982][3] ), .COUT(\CARRYB[983][2] ), .SUM(\SUMB[983][2] ) );
  FADDER S1_982_0 ( .CIN(\ab[982][0] ), .IN0(\CARRYB[981][0] ), .IN1(
        \SUMB[981][1] ), .COUT(\CARRYB[982][0] ), .SUM(PRODUCT[982]) );
  FADDER S2_982_1 ( .CIN(\ab[982][1] ), .IN0(\CARRYB[981][1] ), .IN1(
        \SUMB[981][2] ), .COUT(\CARRYB[982][1] ), .SUM(\SUMB[982][1] ) );
  FADDER S3_982_2 ( .CIN(\ab[982][2] ), .IN0(\CARRYB[981][2] ), .IN1(
        \ab[981][3] ), .COUT(\CARRYB[982][2] ), .SUM(\SUMB[982][2] ) );
  FADDER S1_981_0 ( .CIN(\ab[981][0] ), .IN0(\CARRYB[980][0] ), .IN1(
        \SUMB[980][1] ), .COUT(\CARRYB[981][0] ), .SUM(PRODUCT[981]) );
  FADDER S2_981_1 ( .CIN(\ab[981][1] ), .IN0(\CARRYB[980][1] ), .IN1(
        \SUMB[980][2] ), .COUT(\CARRYB[981][1] ), .SUM(\SUMB[981][1] ) );
  FADDER S3_981_2 ( .CIN(\ab[981][2] ), .IN0(\CARRYB[980][2] ), .IN1(
        \ab[980][3] ), .COUT(\CARRYB[981][2] ), .SUM(\SUMB[981][2] ) );
  FADDER S1_980_0 ( .CIN(\ab[980][0] ), .IN0(\CARRYB[979][0] ), .IN1(
        \SUMB[979][1] ), .COUT(\CARRYB[980][0] ), .SUM(PRODUCT[980]) );
  FADDER S2_980_1 ( .CIN(\ab[980][1] ), .IN0(\CARRYB[979][1] ), .IN1(
        \SUMB[979][2] ), .COUT(\CARRYB[980][1] ), .SUM(\SUMB[980][1] ) );
  FADDER S3_980_2 ( .CIN(\ab[980][2] ), .IN0(\CARRYB[979][2] ), .IN1(
        \ab[979][3] ), .COUT(\CARRYB[980][2] ), .SUM(\SUMB[980][2] ) );
  FADDER S1_979_0 ( .CIN(\ab[979][0] ), .IN0(\CARRYB[978][0] ), .IN1(
        \SUMB[978][1] ), .COUT(\CARRYB[979][0] ), .SUM(PRODUCT[979]) );
  FADDER S2_979_1 ( .CIN(\ab[979][1] ), .IN0(\CARRYB[978][1] ), .IN1(
        \SUMB[978][2] ), .COUT(\CARRYB[979][1] ), .SUM(\SUMB[979][1] ) );
  FADDER S3_979_2 ( .CIN(\ab[979][2] ), .IN0(\CARRYB[978][2] ), .IN1(
        \ab[978][3] ), .COUT(\CARRYB[979][2] ), .SUM(\SUMB[979][2] ) );
  FADDER S1_978_0 ( .CIN(\ab[978][0] ), .IN0(\CARRYB[977][0] ), .IN1(
        \SUMB[977][1] ), .COUT(\CARRYB[978][0] ), .SUM(PRODUCT[978]) );
  FADDER S2_978_1 ( .CIN(\ab[978][1] ), .IN0(\CARRYB[977][1] ), .IN1(
        \SUMB[977][2] ), .COUT(\CARRYB[978][1] ), .SUM(\SUMB[978][1] ) );
  FADDER S3_978_2 ( .CIN(\ab[978][2] ), .IN0(\CARRYB[977][2] ), .IN1(
        \ab[977][3] ), .COUT(\CARRYB[978][2] ), .SUM(\SUMB[978][2] ) );
  FADDER S1_977_0 ( .CIN(\ab[977][0] ), .IN0(\CARRYB[976][0] ), .IN1(
        \SUMB[976][1] ), .COUT(\CARRYB[977][0] ), .SUM(PRODUCT[977]) );
  FADDER S2_977_1 ( .CIN(\ab[977][1] ), .IN0(\CARRYB[976][1] ), .IN1(
        \SUMB[976][2] ), .COUT(\CARRYB[977][1] ), .SUM(\SUMB[977][1] ) );
  FADDER S3_977_2 ( .CIN(\ab[977][2] ), .IN0(\CARRYB[976][2] ), .IN1(
        \ab[976][3] ), .COUT(\CARRYB[977][2] ), .SUM(\SUMB[977][2] ) );
  FADDER S1_976_0 ( .CIN(\ab[976][0] ), .IN0(\CARRYB[975][0] ), .IN1(
        \SUMB[975][1] ), .COUT(\CARRYB[976][0] ), .SUM(PRODUCT[976]) );
  FADDER S2_976_1 ( .CIN(\ab[976][1] ), .IN0(\CARRYB[975][1] ), .IN1(
        \SUMB[975][2] ), .COUT(\CARRYB[976][1] ), .SUM(\SUMB[976][1] ) );
  FADDER S3_976_2 ( .CIN(\ab[976][2] ), .IN0(\CARRYB[975][2] ), .IN1(
        \ab[975][3] ), .COUT(\CARRYB[976][2] ), .SUM(\SUMB[976][2] ) );
  FADDER S1_975_0 ( .CIN(\ab[975][0] ), .IN0(\CARRYB[974][0] ), .IN1(
        \SUMB[974][1] ), .COUT(\CARRYB[975][0] ), .SUM(PRODUCT[975]) );
  FADDER S2_975_1 ( .CIN(\ab[975][1] ), .IN0(\CARRYB[974][1] ), .IN1(
        \SUMB[974][2] ), .COUT(\CARRYB[975][1] ), .SUM(\SUMB[975][1] ) );
  FADDER S3_975_2 ( .CIN(\ab[975][2] ), .IN0(\CARRYB[974][2] ), .IN1(
        \ab[974][3] ), .COUT(\CARRYB[975][2] ), .SUM(\SUMB[975][2] ) );
  FADDER S1_974_0 ( .CIN(\ab[974][0] ), .IN0(\CARRYB[973][0] ), .IN1(
        \SUMB[973][1] ), .COUT(\CARRYB[974][0] ), .SUM(PRODUCT[974]) );
  FADDER S2_974_1 ( .CIN(\ab[974][1] ), .IN0(\CARRYB[973][1] ), .IN1(
        \SUMB[973][2] ), .COUT(\CARRYB[974][1] ), .SUM(\SUMB[974][1] ) );
  FADDER S3_974_2 ( .CIN(\ab[974][2] ), .IN0(\CARRYB[973][2] ), .IN1(
        \ab[973][3] ), .COUT(\CARRYB[974][2] ), .SUM(\SUMB[974][2] ) );
  FADDER S1_973_0 ( .CIN(\ab[973][0] ), .IN0(\CARRYB[972][0] ), .IN1(
        \SUMB[972][1] ), .COUT(\CARRYB[973][0] ), .SUM(PRODUCT[973]) );
  FADDER S2_973_1 ( .CIN(\ab[973][1] ), .IN0(\CARRYB[972][1] ), .IN1(
        \SUMB[972][2] ), .COUT(\CARRYB[973][1] ), .SUM(\SUMB[973][1] ) );
  FADDER S3_973_2 ( .CIN(\ab[973][2] ), .IN0(\CARRYB[972][2] ), .IN1(
        \ab[972][3] ), .COUT(\CARRYB[973][2] ), .SUM(\SUMB[973][2] ) );
  FADDER S1_972_0 ( .CIN(\ab[972][0] ), .IN0(\CARRYB[971][0] ), .IN1(
        \SUMB[971][1] ), .COUT(\CARRYB[972][0] ), .SUM(PRODUCT[972]) );
  FADDER S2_972_1 ( .CIN(\ab[972][1] ), .IN0(\CARRYB[971][1] ), .IN1(
        \SUMB[971][2] ), .COUT(\CARRYB[972][1] ), .SUM(\SUMB[972][1] ) );
  FADDER S3_972_2 ( .CIN(\ab[972][2] ), .IN0(\CARRYB[971][2] ), .IN1(
        \ab[971][3] ), .COUT(\CARRYB[972][2] ), .SUM(\SUMB[972][2] ) );
  FADDER S1_971_0 ( .CIN(\ab[971][0] ), .IN0(\CARRYB[970][0] ), .IN1(
        \SUMB[970][1] ), .COUT(\CARRYB[971][0] ), .SUM(PRODUCT[971]) );
  FADDER S2_971_1 ( .CIN(\ab[971][1] ), .IN0(\CARRYB[970][1] ), .IN1(
        \SUMB[970][2] ), .COUT(\CARRYB[971][1] ), .SUM(\SUMB[971][1] ) );
  FADDER S3_971_2 ( .CIN(\ab[971][2] ), .IN0(\CARRYB[970][2] ), .IN1(
        \ab[970][3] ), .COUT(\CARRYB[971][2] ), .SUM(\SUMB[971][2] ) );
  FADDER S1_970_0 ( .CIN(\ab[970][0] ), .IN0(\CARRYB[969][0] ), .IN1(
        \SUMB[969][1] ), .COUT(\CARRYB[970][0] ), .SUM(PRODUCT[970]) );
  FADDER S2_970_1 ( .CIN(\ab[970][1] ), .IN0(\CARRYB[969][1] ), .IN1(
        \SUMB[969][2] ), .COUT(\CARRYB[970][1] ), .SUM(\SUMB[970][1] ) );
  FADDER S3_970_2 ( .CIN(\ab[970][2] ), .IN0(\CARRYB[969][2] ), .IN1(
        \ab[969][3] ), .COUT(\CARRYB[970][2] ), .SUM(\SUMB[970][2] ) );
  FADDER S1_969_0 ( .CIN(\ab[969][0] ), .IN0(\CARRYB[968][0] ), .IN1(
        \SUMB[968][1] ), .COUT(\CARRYB[969][0] ), .SUM(PRODUCT[969]) );
  FADDER S2_969_1 ( .CIN(\ab[969][1] ), .IN0(\CARRYB[968][1] ), .IN1(
        \SUMB[968][2] ), .COUT(\CARRYB[969][1] ), .SUM(\SUMB[969][1] ) );
  FADDER S3_969_2 ( .CIN(\ab[969][2] ), .IN0(\CARRYB[968][2] ), .IN1(
        \ab[968][3] ), .COUT(\CARRYB[969][2] ), .SUM(\SUMB[969][2] ) );
  FADDER S1_968_0 ( .CIN(\ab[968][0] ), .IN0(\CARRYB[967][0] ), .IN1(
        \SUMB[967][1] ), .COUT(\CARRYB[968][0] ), .SUM(PRODUCT[968]) );
  FADDER S2_968_1 ( .CIN(\ab[968][1] ), .IN0(\CARRYB[967][1] ), .IN1(
        \SUMB[967][2] ), .COUT(\CARRYB[968][1] ), .SUM(\SUMB[968][1] ) );
  FADDER S3_968_2 ( .CIN(\ab[968][2] ), .IN0(\CARRYB[967][2] ), .IN1(
        \ab[967][3] ), .COUT(\CARRYB[968][2] ), .SUM(\SUMB[968][2] ) );
  FADDER S1_967_0 ( .CIN(\ab[967][0] ), .IN0(\CARRYB[966][0] ), .IN1(
        \SUMB[966][1] ), .COUT(\CARRYB[967][0] ), .SUM(PRODUCT[967]) );
  FADDER S2_967_1 ( .CIN(\ab[967][1] ), .IN0(\CARRYB[966][1] ), .IN1(
        \SUMB[966][2] ), .COUT(\CARRYB[967][1] ), .SUM(\SUMB[967][1] ) );
  FADDER S3_967_2 ( .CIN(\ab[967][2] ), .IN0(\CARRYB[966][2] ), .IN1(
        \ab[966][3] ), .COUT(\CARRYB[967][2] ), .SUM(\SUMB[967][2] ) );
  FADDER S1_966_0 ( .CIN(\ab[966][0] ), .IN0(\CARRYB[965][0] ), .IN1(
        \SUMB[965][1] ), .COUT(\CARRYB[966][0] ), .SUM(PRODUCT[966]) );
  FADDER S2_966_1 ( .CIN(\ab[966][1] ), .IN0(\CARRYB[965][1] ), .IN1(
        \SUMB[965][2] ), .COUT(\CARRYB[966][1] ), .SUM(\SUMB[966][1] ) );
  FADDER S3_966_2 ( .CIN(\ab[966][2] ), .IN0(\CARRYB[965][2] ), .IN1(
        \ab[965][3] ), .COUT(\CARRYB[966][2] ), .SUM(\SUMB[966][2] ) );
  FADDER S1_965_0 ( .CIN(\ab[965][0] ), .IN0(\CARRYB[964][0] ), .IN1(
        \SUMB[964][1] ), .COUT(\CARRYB[965][0] ), .SUM(PRODUCT[965]) );
  FADDER S2_965_1 ( .CIN(\ab[965][1] ), .IN0(\CARRYB[964][1] ), .IN1(
        \SUMB[964][2] ), .COUT(\CARRYB[965][1] ), .SUM(\SUMB[965][1] ) );
  FADDER S3_965_2 ( .CIN(\ab[965][2] ), .IN0(\CARRYB[964][2] ), .IN1(
        \ab[964][3] ), .COUT(\CARRYB[965][2] ), .SUM(\SUMB[965][2] ) );
  FADDER S1_964_0 ( .CIN(\ab[964][0] ), .IN0(\CARRYB[963][0] ), .IN1(
        \SUMB[963][1] ), .COUT(\CARRYB[964][0] ), .SUM(PRODUCT[964]) );
  FADDER S2_964_1 ( .CIN(\ab[964][1] ), .IN0(\CARRYB[963][1] ), .IN1(
        \SUMB[963][2] ), .COUT(\CARRYB[964][1] ), .SUM(\SUMB[964][1] ) );
  FADDER S3_964_2 ( .CIN(\ab[964][2] ), .IN0(\CARRYB[963][2] ), .IN1(
        \ab[963][3] ), .COUT(\CARRYB[964][2] ), .SUM(\SUMB[964][2] ) );
  FADDER S1_963_0 ( .CIN(\ab[963][0] ), .IN0(\CARRYB[962][0] ), .IN1(
        \SUMB[962][1] ), .COUT(\CARRYB[963][0] ), .SUM(PRODUCT[963]) );
  FADDER S2_963_1 ( .CIN(\ab[963][1] ), .IN0(\CARRYB[962][1] ), .IN1(
        \SUMB[962][2] ), .COUT(\CARRYB[963][1] ), .SUM(\SUMB[963][1] ) );
  FADDER S3_963_2 ( .CIN(\ab[963][2] ), .IN0(\CARRYB[962][2] ), .IN1(
        \ab[962][3] ), .COUT(\CARRYB[963][2] ), .SUM(\SUMB[963][2] ) );
  FADDER S1_962_0 ( .CIN(\ab[962][0] ), .IN0(\CARRYB[961][0] ), .IN1(
        \SUMB[961][1] ), .COUT(\CARRYB[962][0] ), .SUM(PRODUCT[962]) );
  FADDER S2_962_1 ( .CIN(\ab[962][1] ), .IN0(\CARRYB[961][1] ), .IN1(
        \SUMB[961][2] ), .COUT(\CARRYB[962][1] ), .SUM(\SUMB[962][1] ) );
  FADDER S3_962_2 ( .CIN(\ab[962][2] ), .IN0(\CARRYB[961][2] ), .IN1(
        \ab[961][3] ), .COUT(\CARRYB[962][2] ), .SUM(\SUMB[962][2] ) );
  FADDER S1_961_0 ( .CIN(\ab[961][0] ), .IN0(\CARRYB[960][0] ), .IN1(
        \SUMB[960][1] ), .COUT(\CARRYB[961][0] ), .SUM(PRODUCT[961]) );
  FADDER S2_961_1 ( .CIN(\ab[961][1] ), .IN0(\CARRYB[960][1] ), .IN1(
        \SUMB[960][2] ), .COUT(\CARRYB[961][1] ), .SUM(\SUMB[961][1] ) );
  FADDER S3_961_2 ( .CIN(\ab[961][2] ), .IN0(\CARRYB[960][2] ), .IN1(
        \ab[960][3] ), .COUT(\CARRYB[961][2] ), .SUM(\SUMB[961][2] ) );
  FADDER S1_960_0 ( .CIN(\ab[960][0] ), .IN0(\CARRYB[959][0] ), .IN1(
        \SUMB[959][1] ), .COUT(\CARRYB[960][0] ), .SUM(PRODUCT[960]) );
  FADDER S2_960_1 ( .CIN(\ab[960][1] ), .IN0(\CARRYB[959][1] ), .IN1(
        \SUMB[959][2] ), .COUT(\CARRYB[960][1] ), .SUM(\SUMB[960][1] ) );
  FADDER S3_960_2 ( .CIN(\ab[960][2] ), .IN0(\CARRYB[959][2] ), .IN1(
        \ab[959][3] ), .COUT(\CARRYB[960][2] ), .SUM(\SUMB[960][2] ) );
  FADDER S1_959_0 ( .CIN(\ab[959][0] ), .IN0(\CARRYB[958][0] ), .IN1(
        \SUMB[958][1] ), .COUT(\CARRYB[959][0] ), .SUM(PRODUCT[959]) );
  FADDER S2_959_1 ( .CIN(\ab[959][1] ), .IN0(\CARRYB[958][1] ), .IN1(
        \SUMB[958][2] ), .COUT(\CARRYB[959][1] ), .SUM(\SUMB[959][1] ) );
  FADDER S3_959_2 ( .CIN(\ab[959][2] ), .IN0(\CARRYB[958][2] ), .IN1(
        \ab[958][3] ), .COUT(\CARRYB[959][2] ), .SUM(\SUMB[959][2] ) );
  FADDER S1_958_0 ( .CIN(\ab[958][0] ), .IN0(\CARRYB[957][0] ), .IN1(
        \SUMB[957][1] ), .COUT(\CARRYB[958][0] ), .SUM(PRODUCT[958]) );
  FADDER S2_958_1 ( .CIN(\ab[958][1] ), .IN0(\CARRYB[957][1] ), .IN1(
        \SUMB[957][2] ), .COUT(\CARRYB[958][1] ), .SUM(\SUMB[958][1] ) );
  FADDER S3_958_2 ( .CIN(\ab[958][2] ), .IN0(\CARRYB[957][2] ), .IN1(
        \ab[957][3] ), .COUT(\CARRYB[958][2] ), .SUM(\SUMB[958][2] ) );
  FADDER S1_957_0 ( .CIN(\ab[957][0] ), .IN0(\CARRYB[956][0] ), .IN1(
        \SUMB[956][1] ), .COUT(\CARRYB[957][0] ), .SUM(PRODUCT[957]) );
  FADDER S2_957_1 ( .CIN(\ab[957][1] ), .IN0(\CARRYB[956][1] ), .IN1(
        \SUMB[956][2] ), .COUT(\CARRYB[957][1] ), .SUM(\SUMB[957][1] ) );
  FADDER S3_957_2 ( .CIN(\ab[957][2] ), .IN0(\CARRYB[956][2] ), .IN1(
        \ab[956][3] ), .COUT(\CARRYB[957][2] ), .SUM(\SUMB[957][2] ) );
  FADDER S1_956_0 ( .CIN(\ab[956][0] ), .IN0(\CARRYB[955][0] ), .IN1(
        \SUMB[955][1] ), .COUT(\CARRYB[956][0] ), .SUM(PRODUCT[956]) );
  FADDER S2_956_1 ( .CIN(\ab[956][1] ), .IN0(\CARRYB[955][1] ), .IN1(
        \SUMB[955][2] ), .COUT(\CARRYB[956][1] ), .SUM(\SUMB[956][1] ) );
  FADDER S3_956_2 ( .CIN(\ab[956][2] ), .IN0(\CARRYB[955][2] ), .IN1(
        \ab[955][3] ), .COUT(\CARRYB[956][2] ), .SUM(\SUMB[956][2] ) );
  FADDER S1_955_0 ( .CIN(\ab[955][0] ), .IN0(\CARRYB[954][0] ), .IN1(
        \SUMB[954][1] ), .COUT(\CARRYB[955][0] ), .SUM(PRODUCT[955]) );
  FADDER S2_955_1 ( .CIN(\ab[955][1] ), .IN0(\CARRYB[954][1] ), .IN1(
        \SUMB[954][2] ), .COUT(\CARRYB[955][1] ), .SUM(\SUMB[955][1] ) );
  FADDER S3_955_2 ( .CIN(\ab[955][2] ), .IN0(\CARRYB[954][2] ), .IN1(
        \ab[954][3] ), .COUT(\CARRYB[955][2] ), .SUM(\SUMB[955][2] ) );
  FADDER S1_954_0 ( .CIN(\ab[954][0] ), .IN0(\CARRYB[953][0] ), .IN1(
        \SUMB[953][1] ), .COUT(\CARRYB[954][0] ), .SUM(PRODUCT[954]) );
  FADDER S2_954_1 ( .CIN(\ab[954][1] ), .IN0(\CARRYB[953][1] ), .IN1(
        \SUMB[953][2] ), .COUT(\CARRYB[954][1] ), .SUM(\SUMB[954][1] ) );
  FADDER S3_954_2 ( .CIN(\ab[954][2] ), .IN0(\CARRYB[953][2] ), .IN1(
        \ab[953][3] ), .COUT(\CARRYB[954][2] ), .SUM(\SUMB[954][2] ) );
  FADDER S1_953_0 ( .CIN(\ab[953][0] ), .IN0(\CARRYB[952][0] ), .IN1(
        \SUMB[952][1] ), .COUT(\CARRYB[953][0] ), .SUM(PRODUCT[953]) );
  FADDER S2_953_1 ( .CIN(\ab[953][1] ), .IN0(\CARRYB[952][1] ), .IN1(
        \SUMB[952][2] ), .COUT(\CARRYB[953][1] ), .SUM(\SUMB[953][1] ) );
  FADDER S3_953_2 ( .CIN(\ab[953][2] ), .IN0(\CARRYB[952][2] ), .IN1(
        \ab[952][3] ), .COUT(\CARRYB[953][2] ), .SUM(\SUMB[953][2] ) );
  FADDER S1_952_0 ( .CIN(\ab[952][0] ), .IN0(\CARRYB[951][0] ), .IN1(
        \SUMB[951][1] ), .COUT(\CARRYB[952][0] ), .SUM(PRODUCT[952]) );
  FADDER S2_952_1 ( .CIN(\ab[952][1] ), .IN0(\CARRYB[951][1] ), .IN1(
        \SUMB[951][2] ), .COUT(\CARRYB[952][1] ), .SUM(\SUMB[952][1] ) );
  FADDER S3_952_2 ( .CIN(\ab[952][2] ), .IN0(\CARRYB[951][2] ), .IN1(
        \ab[951][3] ), .COUT(\CARRYB[952][2] ), .SUM(\SUMB[952][2] ) );
  FADDER S1_951_0 ( .CIN(\ab[951][0] ), .IN0(\CARRYB[950][0] ), .IN1(
        \SUMB[950][1] ), .COUT(\CARRYB[951][0] ), .SUM(PRODUCT[951]) );
  FADDER S2_951_1 ( .CIN(\ab[951][1] ), .IN0(\CARRYB[950][1] ), .IN1(
        \SUMB[950][2] ), .COUT(\CARRYB[951][1] ), .SUM(\SUMB[951][1] ) );
  FADDER S3_951_2 ( .CIN(\ab[951][2] ), .IN0(\CARRYB[950][2] ), .IN1(
        \ab[950][3] ), .COUT(\CARRYB[951][2] ), .SUM(\SUMB[951][2] ) );
  FADDER S1_950_0 ( .CIN(\ab[950][0] ), .IN0(\CARRYB[949][0] ), .IN1(
        \SUMB[949][1] ), .COUT(\CARRYB[950][0] ), .SUM(PRODUCT[950]) );
  FADDER S2_950_1 ( .CIN(\ab[950][1] ), .IN0(\CARRYB[949][1] ), .IN1(
        \SUMB[949][2] ), .COUT(\CARRYB[950][1] ), .SUM(\SUMB[950][1] ) );
  FADDER S3_950_2 ( .CIN(\ab[950][2] ), .IN0(\CARRYB[949][2] ), .IN1(
        \ab[949][3] ), .COUT(\CARRYB[950][2] ), .SUM(\SUMB[950][2] ) );
  FADDER S1_949_0 ( .CIN(\ab[949][0] ), .IN0(\CARRYB[948][0] ), .IN1(
        \SUMB[948][1] ), .COUT(\CARRYB[949][0] ), .SUM(PRODUCT[949]) );
  FADDER S2_949_1 ( .CIN(\ab[949][1] ), .IN0(\CARRYB[948][1] ), .IN1(
        \SUMB[948][2] ), .COUT(\CARRYB[949][1] ), .SUM(\SUMB[949][1] ) );
  FADDER S3_949_2 ( .CIN(\ab[949][2] ), .IN0(\CARRYB[948][2] ), .IN1(
        \ab[948][3] ), .COUT(\CARRYB[949][2] ), .SUM(\SUMB[949][2] ) );
  FADDER S1_948_0 ( .CIN(\ab[948][0] ), .IN0(\CARRYB[947][0] ), .IN1(
        \SUMB[947][1] ), .COUT(\CARRYB[948][0] ), .SUM(PRODUCT[948]) );
  FADDER S2_948_1 ( .CIN(\ab[948][1] ), .IN0(\CARRYB[947][1] ), .IN1(
        \SUMB[947][2] ), .COUT(\CARRYB[948][1] ), .SUM(\SUMB[948][1] ) );
  FADDER S3_948_2 ( .CIN(\ab[948][2] ), .IN0(\CARRYB[947][2] ), .IN1(
        \ab[947][3] ), .COUT(\CARRYB[948][2] ), .SUM(\SUMB[948][2] ) );
  FADDER S1_947_0 ( .CIN(\ab[947][0] ), .IN0(\CARRYB[946][0] ), .IN1(
        \SUMB[946][1] ), .COUT(\CARRYB[947][0] ), .SUM(PRODUCT[947]) );
  FADDER S2_947_1 ( .CIN(\ab[947][1] ), .IN0(\CARRYB[946][1] ), .IN1(
        \SUMB[946][2] ), .COUT(\CARRYB[947][1] ), .SUM(\SUMB[947][1] ) );
  FADDER S3_947_2 ( .CIN(\ab[947][2] ), .IN0(\CARRYB[946][2] ), .IN1(
        \ab[946][3] ), .COUT(\CARRYB[947][2] ), .SUM(\SUMB[947][2] ) );
  FADDER S1_946_0 ( .CIN(\ab[946][0] ), .IN0(\CARRYB[945][0] ), .IN1(
        \SUMB[945][1] ), .COUT(\CARRYB[946][0] ), .SUM(PRODUCT[946]) );
  FADDER S2_946_1 ( .CIN(\ab[946][1] ), .IN0(\CARRYB[945][1] ), .IN1(
        \SUMB[945][2] ), .COUT(\CARRYB[946][1] ), .SUM(\SUMB[946][1] ) );
  FADDER S3_946_2 ( .CIN(\ab[946][2] ), .IN0(\CARRYB[945][2] ), .IN1(
        \ab[945][3] ), .COUT(\CARRYB[946][2] ), .SUM(\SUMB[946][2] ) );
  FADDER S1_945_0 ( .CIN(\ab[945][0] ), .IN0(\CARRYB[944][0] ), .IN1(
        \SUMB[944][1] ), .COUT(\CARRYB[945][0] ), .SUM(PRODUCT[945]) );
  FADDER S2_945_1 ( .CIN(\ab[945][1] ), .IN0(\CARRYB[944][1] ), .IN1(
        \SUMB[944][2] ), .COUT(\CARRYB[945][1] ), .SUM(\SUMB[945][1] ) );
  FADDER S3_945_2 ( .CIN(\ab[945][2] ), .IN0(\CARRYB[944][2] ), .IN1(
        \ab[944][3] ), .COUT(\CARRYB[945][2] ), .SUM(\SUMB[945][2] ) );
  FADDER S1_944_0 ( .CIN(\ab[944][0] ), .IN0(\CARRYB[943][0] ), .IN1(
        \SUMB[943][1] ), .COUT(\CARRYB[944][0] ), .SUM(PRODUCT[944]) );
  FADDER S2_944_1 ( .CIN(\ab[944][1] ), .IN0(\CARRYB[943][1] ), .IN1(
        \SUMB[943][2] ), .COUT(\CARRYB[944][1] ), .SUM(\SUMB[944][1] ) );
  FADDER S3_944_2 ( .CIN(\ab[944][2] ), .IN0(\CARRYB[943][2] ), .IN1(
        \ab[943][3] ), .COUT(\CARRYB[944][2] ), .SUM(\SUMB[944][2] ) );
  FADDER S1_943_0 ( .CIN(\ab[943][0] ), .IN0(\CARRYB[942][0] ), .IN1(
        \SUMB[942][1] ), .COUT(\CARRYB[943][0] ), .SUM(PRODUCT[943]) );
  FADDER S2_943_1 ( .CIN(\ab[943][1] ), .IN0(\CARRYB[942][1] ), .IN1(
        \SUMB[942][2] ), .COUT(\CARRYB[943][1] ), .SUM(\SUMB[943][1] ) );
  FADDER S3_943_2 ( .CIN(\ab[943][2] ), .IN0(\CARRYB[942][2] ), .IN1(
        \ab[942][3] ), .COUT(\CARRYB[943][2] ), .SUM(\SUMB[943][2] ) );
  FADDER S1_942_0 ( .CIN(\ab[942][0] ), .IN0(\CARRYB[941][0] ), .IN1(
        \SUMB[941][1] ), .COUT(\CARRYB[942][0] ), .SUM(PRODUCT[942]) );
  FADDER S2_942_1 ( .CIN(\ab[942][1] ), .IN0(\CARRYB[941][1] ), .IN1(
        \SUMB[941][2] ), .COUT(\CARRYB[942][1] ), .SUM(\SUMB[942][1] ) );
  FADDER S3_942_2 ( .CIN(\ab[942][2] ), .IN0(\CARRYB[941][2] ), .IN1(
        \ab[941][3] ), .COUT(\CARRYB[942][2] ), .SUM(\SUMB[942][2] ) );
  FADDER S1_941_0 ( .CIN(\ab[941][0] ), .IN0(\CARRYB[940][0] ), .IN1(
        \SUMB[940][1] ), .COUT(\CARRYB[941][0] ), .SUM(PRODUCT[941]) );
  FADDER S2_941_1 ( .CIN(\ab[941][1] ), .IN0(\CARRYB[940][1] ), .IN1(
        \SUMB[940][2] ), .COUT(\CARRYB[941][1] ), .SUM(\SUMB[941][1] ) );
  FADDER S3_941_2 ( .CIN(\ab[941][2] ), .IN0(\CARRYB[940][2] ), .IN1(
        \ab[940][3] ), .COUT(\CARRYB[941][2] ), .SUM(\SUMB[941][2] ) );
  FADDER S1_940_0 ( .CIN(\ab[940][0] ), .IN0(\CARRYB[939][0] ), .IN1(
        \SUMB[939][1] ), .COUT(\CARRYB[940][0] ), .SUM(PRODUCT[940]) );
  FADDER S2_940_1 ( .CIN(\ab[940][1] ), .IN0(\CARRYB[939][1] ), .IN1(
        \SUMB[939][2] ), .COUT(\CARRYB[940][1] ), .SUM(\SUMB[940][1] ) );
  FADDER S3_940_2 ( .CIN(\ab[940][2] ), .IN0(\CARRYB[939][2] ), .IN1(
        \ab[939][3] ), .COUT(\CARRYB[940][2] ), .SUM(\SUMB[940][2] ) );
  FADDER S1_939_0 ( .CIN(\ab[939][0] ), .IN0(\CARRYB[938][0] ), .IN1(
        \SUMB[938][1] ), .COUT(\CARRYB[939][0] ), .SUM(PRODUCT[939]) );
  FADDER S2_939_1 ( .CIN(\ab[939][1] ), .IN0(\CARRYB[938][1] ), .IN1(
        \SUMB[938][2] ), .COUT(\CARRYB[939][1] ), .SUM(\SUMB[939][1] ) );
  FADDER S3_939_2 ( .CIN(\ab[939][2] ), .IN0(\CARRYB[938][2] ), .IN1(
        \ab[938][3] ), .COUT(\CARRYB[939][2] ), .SUM(\SUMB[939][2] ) );
  FADDER S1_938_0 ( .CIN(\ab[938][0] ), .IN0(\CARRYB[937][0] ), .IN1(
        \SUMB[937][1] ), .COUT(\CARRYB[938][0] ), .SUM(PRODUCT[938]) );
  FADDER S2_938_1 ( .CIN(\ab[938][1] ), .IN0(\CARRYB[937][1] ), .IN1(
        \SUMB[937][2] ), .COUT(\CARRYB[938][1] ), .SUM(\SUMB[938][1] ) );
  FADDER S3_938_2 ( .CIN(\ab[938][2] ), .IN0(\CARRYB[937][2] ), .IN1(
        \ab[937][3] ), .COUT(\CARRYB[938][2] ), .SUM(\SUMB[938][2] ) );
  FADDER S1_937_0 ( .CIN(\ab[937][0] ), .IN0(\CARRYB[936][0] ), .IN1(
        \SUMB[936][1] ), .COUT(\CARRYB[937][0] ), .SUM(PRODUCT[937]) );
  FADDER S2_937_1 ( .CIN(\ab[937][1] ), .IN0(\CARRYB[936][1] ), .IN1(
        \SUMB[936][2] ), .COUT(\CARRYB[937][1] ), .SUM(\SUMB[937][1] ) );
  FADDER S3_937_2 ( .CIN(\ab[937][2] ), .IN0(\CARRYB[936][2] ), .IN1(
        \ab[936][3] ), .COUT(\CARRYB[937][2] ), .SUM(\SUMB[937][2] ) );
  FADDER S1_936_0 ( .CIN(\ab[936][0] ), .IN0(\CARRYB[935][0] ), .IN1(
        \SUMB[935][1] ), .COUT(\CARRYB[936][0] ), .SUM(PRODUCT[936]) );
  FADDER S2_936_1 ( .CIN(\ab[936][1] ), .IN0(\CARRYB[935][1] ), .IN1(
        \SUMB[935][2] ), .COUT(\CARRYB[936][1] ), .SUM(\SUMB[936][1] ) );
  FADDER S3_936_2 ( .CIN(\ab[936][2] ), .IN0(\CARRYB[935][2] ), .IN1(
        \ab[935][3] ), .COUT(\CARRYB[936][2] ), .SUM(\SUMB[936][2] ) );
  FADDER S1_935_0 ( .CIN(\ab[935][0] ), .IN0(\CARRYB[934][0] ), .IN1(
        \SUMB[934][1] ), .COUT(\CARRYB[935][0] ), .SUM(PRODUCT[935]) );
  FADDER S2_935_1 ( .CIN(\ab[935][1] ), .IN0(\CARRYB[934][1] ), .IN1(
        \SUMB[934][2] ), .COUT(\CARRYB[935][1] ), .SUM(\SUMB[935][1] ) );
  FADDER S3_935_2 ( .CIN(\ab[935][2] ), .IN0(\CARRYB[934][2] ), .IN1(
        \ab[934][3] ), .COUT(\CARRYB[935][2] ), .SUM(\SUMB[935][2] ) );
  FADDER S1_934_0 ( .CIN(\ab[934][0] ), .IN0(\CARRYB[933][0] ), .IN1(
        \SUMB[933][1] ), .COUT(\CARRYB[934][0] ), .SUM(PRODUCT[934]) );
  FADDER S2_934_1 ( .CIN(\ab[934][1] ), .IN0(\CARRYB[933][1] ), .IN1(
        \SUMB[933][2] ), .COUT(\CARRYB[934][1] ), .SUM(\SUMB[934][1] ) );
  FADDER S3_934_2 ( .CIN(\ab[934][2] ), .IN0(\CARRYB[933][2] ), .IN1(
        \ab[933][3] ), .COUT(\CARRYB[934][2] ), .SUM(\SUMB[934][2] ) );
  FADDER S1_933_0 ( .CIN(\ab[933][0] ), .IN0(\CARRYB[932][0] ), .IN1(
        \SUMB[932][1] ), .COUT(\CARRYB[933][0] ), .SUM(PRODUCT[933]) );
  FADDER S2_933_1 ( .CIN(\ab[933][1] ), .IN0(\CARRYB[932][1] ), .IN1(
        \SUMB[932][2] ), .COUT(\CARRYB[933][1] ), .SUM(\SUMB[933][1] ) );
  FADDER S3_933_2 ( .CIN(\ab[933][2] ), .IN0(\CARRYB[932][2] ), .IN1(
        \ab[932][3] ), .COUT(\CARRYB[933][2] ), .SUM(\SUMB[933][2] ) );
  FADDER S1_932_0 ( .CIN(\ab[932][0] ), .IN0(\CARRYB[931][0] ), .IN1(
        \SUMB[931][1] ), .COUT(\CARRYB[932][0] ), .SUM(PRODUCT[932]) );
  FADDER S2_932_1 ( .CIN(\ab[932][1] ), .IN0(\CARRYB[931][1] ), .IN1(
        \SUMB[931][2] ), .COUT(\CARRYB[932][1] ), .SUM(\SUMB[932][1] ) );
  FADDER S3_932_2 ( .CIN(\ab[932][2] ), .IN0(\CARRYB[931][2] ), .IN1(
        \ab[931][3] ), .COUT(\CARRYB[932][2] ), .SUM(\SUMB[932][2] ) );
  FADDER S1_931_0 ( .CIN(\ab[931][0] ), .IN0(\CARRYB[930][0] ), .IN1(
        \SUMB[930][1] ), .COUT(\CARRYB[931][0] ), .SUM(PRODUCT[931]) );
  FADDER S2_931_1 ( .CIN(\ab[931][1] ), .IN0(\CARRYB[930][1] ), .IN1(
        \SUMB[930][2] ), .COUT(\CARRYB[931][1] ), .SUM(\SUMB[931][1] ) );
  FADDER S3_931_2 ( .CIN(\ab[931][2] ), .IN0(\CARRYB[930][2] ), .IN1(
        \ab[930][3] ), .COUT(\CARRYB[931][2] ), .SUM(\SUMB[931][2] ) );
  FADDER S1_930_0 ( .CIN(\ab[930][0] ), .IN0(\CARRYB[929][0] ), .IN1(
        \SUMB[929][1] ), .COUT(\CARRYB[930][0] ), .SUM(PRODUCT[930]) );
  FADDER S2_930_1 ( .CIN(\ab[930][1] ), .IN0(\CARRYB[929][1] ), .IN1(
        \SUMB[929][2] ), .COUT(\CARRYB[930][1] ), .SUM(\SUMB[930][1] ) );
  FADDER S3_930_2 ( .CIN(\ab[930][2] ), .IN0(\CARRYB[929][2] ), .IN1(
        \ab[929][3] ), .COUT(\CARRYB[930][2] ), .SUM(\SUMB[930][2] ) );
  FADDER S1_929_0 ( .CIN(\ab[929][0] ), .IN0(\CARRYB[928][0] ), .IN1(
        \SUMB[928][1] ), .COUT(\CARRYB[929][0] ), .SUM(PRODUCT[929]) );
  FADDER S2_929_1 ( .CIN(\ab[929][1] ), .IN0(\CARRYB[928][1] ), .IN1(
        \SUMB[928][2] ), .COUT(\CARRYB[929][1] ), .SUM(\SUMB[929][1] ) );
  FADDER S3_929_2 ( .CIN(\ab[929][2] ), .IN0(\CARRYB[928][2] ), .IN1(
        \ab[928][3] ), .COUT(\CARRYB[929][2] ), .SUM(\SUMB[929][2] ) );
  FADDER S1_928_0 ( .CIN(\ab[928][0] ), .IN0(\CARRYB[927][0] ), .IN1(
        \SUMB[927][1] ), .COUT(\CARRYB[928][0] ), .SUM(PRODUCT[928]) );
  FADDER S2_928_1 ( .CIN(\ab[928][1] ), .IN0(\CARRYB[927][1] ), .IN1(
        \SUMB[927][2] ), .COUT(\CARRYB[928][1] ), .SUM(\SUMB[928][1] ) );
  FADDER S3_928_2 ( .CIN(\ab[928][2] ), .IN0(\CARRYB[927][2] ), .IN1(
        \ab[927][3] ), .COUT(\CARRYB[928][2] ), .SUM(\SUMB[928][2] ) );
  FADDER S1_927_0 ( .CIN(\ab[927][0] ), .IN0(\CARRYB[926][0] ), .IN1(
        \SUMB[926][1] ), .COUT(\CARRYB[927][0] ), .SUM(PRODUCT[927]) );
  FADDER S2_927_1 ( .CIN(\ab[927][1] ), .IN0(\CARRYB[926][1] ), .IN1(
        \SUMB[926][2] ), .COUT(\CARRYB[927][1] ), .SUM(\SUMB[927][1] ) );
  FADDER S3_927_2 ( .CIN(\ab[927][2] ), .IN0(\CARRYB[926][2] ), .IN1(
        \ab[926][3] ), .COUT(\CARRYB[927][2] ), .SUM(\SUMB[927][2] ) );
  FADDER S1_926_0 ( .CIN(\ab[926][0] ), .IN0(\CARRYB[925][0] ), .IN1(
        \SUMB[925][1] ), .COUT(\CARRYB[926][0] ), .SUM(PRODUCT[926]) );
  FADDER S2_926_1 ( .CIN(\ab[926][1] ), .IN0(\CARRYB[925][1] ), .IN1(
        \SUMB[925][2] ), .COUT(\CARRYB[926][1] ), .SUM(\SUMB[926][1] ) );
  FADDER S3_926_2 ( .CIN(\ab[926][2] ), .IN0(\CARRYB[925][2] ), .IN1(
        \ab[925][3] ), .COUT(\CARRYB[926][2] ), .SUM(\SUMB[926][2] ) );
  FADDER S1_925_0 ( .CIN(\ab[925][0] ), .IN0(\CARRYB[924][0] ), .IN1(
        \SUMB[924][1] ), .COUT(\CARRYB[925][0] ), .SUM(PRODUCT[925]) );
  FADDER S2_925_1 ( .CIN(\ab[925][1] ), .IN0(\CARRYB[924][1] ), .IN1(
        \SUMB[924][2] ), .COUT(\CARRYB[925][1] ), .SUM(\SUMB[925][1] ) );
  FADDER S3_925_2 ( .CIN(\ab[925][2] ), .IN0(\CARRYB[924][2] ), .IN1(
        \ab[924][3] ), .COUT(\CARRYB[925][2] ), .SUM(\SUMB[925][2] ) );
  FADDER S1_924_0 ( .CIN(\ab[924][0] ), .IN0(\CARRYB[923][0] ), .IN1(
        \SUMB[923][1] ), .COUT(\CARRYB[924][0] ), .SUM(PRODUCT[924]) );
  FADDER S2_924_1 ( .CIN(\ab[924][1] ), .IN0(\CARRYB[923][1] ), .IN1(
        \SUMB[923][2] ), .COUT(\CARRYB[924][1] ), .SUM(\SUMB[924][1] ) );
  FADDER S3_924_2 ( .CIN(\ab[924][2] ), .IN0(\CARRYB[923][2] ), .IN1(
        \ab[923][3] ), .COUT(\CARRYB[924][2] ), .SUM(\SUMB[924][2] ) );
  FADDER S1_923_0 ( .CIN(\ab[923][0] ), .IN0(\CARRYB[922][0] ), .IN1(
        \SUMB[922][1] ), .COUT(\CARRYB[923][0] ), .SUM(PRODUCT[923]) );
  FADDER S2_923_1 ( .CIN(\ab[923][1] ), .IN0(\CARRYB[922][1] ), .IN1(
        \SUMB[922][2] ), .COUT(\CARRYB[923][1] ), .SUM(\SUMB[923][1] ) );
  FADDER S3_923_2 ( .CIN(\ab[923][2] ), .IN0(\CARRYB[922][2] ), .IN1(
        \ab[922][3] ), .COUT(\CARRYB[923][2] ), .SUM(\SUMB[923][2] ) );
  FADDER S1_922_0 ( .CIN(\ab[922][0] ), .IN0(\CARRYB[921][0] ), .IN1(
        \SUMB[921][1] ), .COUT(\CARRYB[922][0] ), .SUM(PRODUCT[922]) );
  FADDER S2_922_1 ( .CIN(\ab[922][1] ), .IN0(\CARRYB[921][1] ), .IN1(
        \SUMB[921][2] ), .COUT(\CARRYB[922][1] ), .SUM(\SUMB[922][1] ) );
  FADDER S3_922_2 ( .CIN(\ab[922][2] ), .IN0(\CARRYB[921][2] ), .IN1(
        \ab[921][3] ), .COUT(\CARRYB[922][2] ), .SUM(\SUMB[922][2] ) );
  FADDER S1_921_0 ( .CIN(\ab[921][0] ), .IN0(\CARRYB[920][0] ), .IN1(
        \SUMB[920][1] ), .COUT(\CARRYB[921][0] ), .SUM(PRODUCT[921]) );
  FADDER S2_921_1 ( .CIN(\ab[921][1] ), .IN0(\CARRYB[920][1] ), .IN1(
        \SUMB[920][2] ), .COUT(\CARRYB[921][1] ), .SUM(\SUMB[921][1] ) );
  FADDER S3_921_2 ( .CIN(\ab[921][2] ), .IN0(\CARRYB[920][2] ), .IN1(
        \ab[920][3] ), .COUT(\CARRYB[921][2] ), .SUM(\SUMB[921][2] ) );
  FADDER S1_920_0 ( .CIN(\ab[920][0] ), .IN0(\CARRYB[919][0] ), .IN1(
        \SUMB[919][1] ), .COUT(\CARRYB[920][0] ), .SUM(PRODUCT[920]) );
  FADDER S2_920_1 ( .CIN(\ab[920][1] ), .IN0(\CARRYB[919][1] ), .IN1(
        \SUMB[919][2] ), .COUT(\CARRYB[920][1] ), .SUM(\SUMB[920][1] ) );
  FADDER S3_920_2 ( .CIN(\ab[920][2] ), .IN0(\CARRYB[919][2] ), .IN1(
        \ab[919][3] ), .COUT(\CARRYB[920][2] ), .SUM(\SUMB[920][2] ) );
  FADDER S1_919_0 ( .CIN(\ab[919][0] ), .IN0(\CARRYB[918][0] ), .IN1(
        \SUMB[918][1] ), .COUT(\CARRYB[919][0] ), .SUM(PRODUCT[919]) );
  FADDER S2_919_1 ( .CIN(\ab[919][1] ), .IN0(\CARRYB[918][1] ), .IN1(
        \SUMB[918][2] ), .COUT(\CARRYB[919][1] ), .SUM(\SUMB[919][1] ) );
  FADDER S3_919_2 ( .CIN(\ab[919][2] ), .IN0(\CARRYB[918][2] ), .IN1(
        \ab[918][3] ), .COUT(\CARRYB[919][2] ), .SUM(\SUMB[919][2] ) );
  FADDER S1_918_0 ( .CIN(\ab[918][0] ), .IN0(\CARRYB[917][0] ), .IN1(
        \SUMB[917][1] ), .COUT(\CARRYB[918][0] ), .SUM(PRODUCT[918]) );
  FADDER S2_918_1 ( .CIN(\ab[918][1] ), .IN0(\CARRYB[917][1] ), .IN1(
        \SUMB[917][2] ), .COUT(\CARRYB[918][1] ), .SUM(\SUMB[918][1] ) );
  FADDER S3_918_2 ( .CIN(\ab[918][2] ), .IN0(\CARRYB[917][2] ), .IN1(
        \ab[917][3] ), .COUT(\CARRYB[918][2] ), .SUM(\SUMB[918][2] ) );
  FADDER S1_917_0 ( .CIN(\ab[917][0] ), .IN0(\CARRYB[916][0] ), .IN1(
        \SUMB[916][1] ), .COUT(\CARRYB[917][0] ), .SUM(PRODUCT[917]) );
  FADDER S2_917_1 ( .CIN(\ab[917][1] ), .IN0(\CARRYB[916][1] ), .IN1(
        \SUMB[916][2] ), .COUT(\CARRYB[917][1] ), .SUM(\SUMB[917][1] ) );
  FADDER S3_917_2 ( .CIN(\ab[917][2] ), .IN0(\CARRYB[916][2] ), .IN1(
        \ab[916][3] ), .COUT(\CARRYB[917][2] ), .SUM(\SUMB[917][2] ) );
  FADDER S1_916_0 ( .CIN(\ab[916][0] ), .IN0(\CARRYB[915][0] ), .IN1(
        \SUMB[915][1] ), .COUT(\CARRYB[916][0] ), .SUM(PRODUCT[916]) );
  FADDER S2_916_1 ( .CIN(\ab[916][1] ), .IN0(\CARRYB[915][1] ), .IN1(
        \SUMB[915][2] ), .COUT(\CARRYB[916][1] ), .SUM(\SUMB[916][1] ) );
  FADDER S3_916_2 ( .CIN(\ab[916][2] ), .IN0(\CARRYB[915][2] ), .IN1(
        \ab[915][3] ), .COUT(\CARRYB[916][2] ), .SUM(\SUMB[916][2] ) );
  FADDER S1_915_0 ( .CIN(\ab[915][0] ), .IN0(\CARRYB[914][0] ), .IN1(
        \SUMB[914][1] ), .COUT(\CARRYB[915][0] ), .SUM(PRODUCT[915]) );
  FADDER S2_915_1 ( .CIN(\ab[915][1] ), .IN0(\CARRYB[914][1] ), .IN1(
        \SUMB[914][2] ), .COUT(\CARRYB[915][1] ), .SUM(\SUMB[915][1] ) );
  FADDER S3_915_2 ( .CIN(\ab[915][2] ), .IN0(\CARRYB[914][2] ), .IN1(
        \ab[914][3] ), .COUT(\CARRYB[915][2] ), .SUM(\SUMB[915][2] ) );
  FADDER S1_914_0 ( .CIN(\ab[914][0] ), .IN0(\CARRYB[913][0] ), .IN1(
        \SUMB[913][1] ), .COUT(\CARRYB[914][0] ), .SUM(PRODUCT[914]) );
  FADDER S2_914_1 ( .CIN(\ab[914][1] ), .IN0(\CARRYB[913][1] ), .IN1(
        \SUMB[913][2] ), .COUT(\CARRYB[914][1] ), .SUM(\SUMB[914][1] ) );
  FADDER S3_914_2 ( .CIN(\ab[914][2] ), .IN0(\CARRYB[913][2] ), .IN1(
        \ab[913][3] ), .COUT(\CARRYB[914][2] ), .SUM(\SUMB[914][2] ) );
  FADDER S1_913_0 ( .CIN(\ab[913][0] ), .IN0(\CARRYB[912][0] ), .IN1(
        \SUMB[912][1] ), .COUT(\CARRYB[913][0] ), .SUM(PRODUCT[913]) );
  FADDER S2_913_1 ( .CIN(\ab[913][1] ), .IN0(\CARRYB[912][1] ), .IN1(
        \SUMB[912][2] ), .COUT(\CARRYB[913][1] ), .SUM(\SUMB[913][1] ) );
  FADDER S3_913_2 ( .CIN(\ab[913][2] ), .IN0(\CARRYB[912][2] ), .IN1(
        \ab[912][3] ), .COUT(\CARRYB[913][2] ), .SUM(\SUMB[913][2] ) );
  FADDER S1_912_0 ( .CIN(\ab[912][0] ), .IN0(\CARRYB[911][0] ), .IN1(
        \SUMB[911][1] ), .COUT(\CARRYB[912][0] ), .SUM(PRODUCT[912]) );
  FADDER S2_912_1 ( .CIN(\ab[912][1] ), .IN0(\CARRYB[911][1] ), .IN1(
        \SUMB[911][2] ), .COUT(\CARRYB[912][1] ), .SUM(\SUMB[912][1] ) );
  FADDER S3_912_2 ( .CIN(\ab[912][2] ), .IN0(\CARRYB[911][2] ), .IN1(
        \ab[911][3] ), .COUT(\CARRYB[912][2] ), .SUM(\SUMB[912][2] ) );
  FADDER S1_911_0 ( .CIN(\ab[911][0] ), .IN0(\CARRYB[910][0] ), .IN1(
        \SUMB[910][1] ), .COUT(\CARRYB[911][0] ), .SUM(PRODUCT[911]) );
  FADDER S2_911_1 ( .CIN(\ab[911][1] ), .IN0(\CARRYB[910][1] ), .IN1(
        \SUMB[910][2] ), .COUT(\CARRYB[911][1] ), .SUM(\SUMB[911][1] ) );
  FADDER S3_911_2 ( .CIN(\ab[911][2] ), .IN0(\CARRYB[910][2] ), .IN1(
        \ab[910][3] ), .COUT(\CARRYB[911][2] ), .SUM(\SUMB[911][2] ) );
  FADDER S1_910_0 ( .CIN(\ab[910][0] ), .IN0(\CARRYB[909][0] ), .IN1(
        \SUMB[909][1] ), .COUT(\CARRYB[910][0] ), .SUM(PRODUCT[910]) );
  FADDER S2_910_1 ( .CIN(\ab[910][1] ), .IN0(\CARRYB[909][1] ), .IN1(
        \SUMB[909][2] ), .COUT(\CARRYB[910][1] ), .SUM(\SUMB[910][1] ) );
  FADDER S3_910_2 ( .CIN(\ab[910][2] ), .IN0(\CARRYB[909][2] ), .IN1(
        \ab[909][3] ), .COUT(\CARRYB[910][2] ), .SUM(\SUMB[910][2] ) );
  FADDER S1_909_0 ( .CIN(\ab[909][0] ), .IN0(\CARRYB[908][0] ), .IN1(
        \SUMB[908][1] ), .COUT(\CARRYB[909][0] ), .SUM(PRODUCT[909]) );
  FADDER S2_909_1 ( .CIN(\ab[909][1] ), .IN0(\CARRYB[908][1] ), .IN1(
        \SUMB[908][2] ), .COUT(\CARRYB[909][1] ), .SUM(\SUMB[909][1] ) );
  FADDER S3_909_2 ( .CIN(\ab[909][2] ), .IN0(\CARRYB[908][2] ), .IN1(
        \ab[908][3] ), .COUT(\CARRYB[909][2] ), .SUM(\SUMB[909][2] ) );
  FADDER S1_908_0 ( .CIN(\ab[908][0] ), .IN0(\CARRYB[907][0] ), .IN1(
        \SUMB[907][1] ), .COUT(\CARRYB[908][0] ), .SUM(PRODUCT[908]) );
  FADDER S2_908_1 ( .CIN(\ab[908][1] ), .IN0(\CARRYB[907][1] ), .IN1(
        \SUMB[907][2] ), .COUT(\CARRYB[908][1] ), .SUM(\SUMB[908][1] ) );
  FADDER S3_908_2 ( .CIN(\ab[908][2] ), .IN0(\CARRYB[907][2] ), .IN1(
        \ab[907][3] ), .COUT(\CARRYB[908][2] ), .SUM(\SUMB[908][2] ) );
  FADDER S1_907_0 ( .CIN(\ab[907][0] ), .IN0(\CARRYB[906][0] ), .IN1(
        \SUMB[906][1] ), .COUT(\CARRYB[907][0] ), .SUM(PRODUCT[907]) );
  FADDER S2_907_1 ( .CIN(\ab[907][1] ), .IN0(\CARRYB[906][1] ), .IN1(
        \SUMB[906][2] ), .COUT(\CARRYB[907][1] ), .SUM(\SUMB[907][1] ) );
  FADDER S3_907_2 ( .CIN(\ab[907][2] ), .IN0(\CARRYB[906][2] ), .IN1(
        \ab[906][3] ), .COUT(\CARRYB[907][2] ), .SUM(\SUMB[907][2] ) );
  FADDER S1_906_0 ( .CIN(\ab[906][0] ), .IN0(\CARRYB[905][0] ), .IN1(
        \SUMB[905][1] ), .COUT(\CARRYB[906][0] ), .SUM(PRODUCT[906]) );
  FADDER S2_906_1 ( .CIN(\ab[906][1] ), .IN0(\CARRYB[905][1] ), .IN1(
        \SUMB[905][2] ), .COUT(\CARRYB[906][1] ), .SUM(\SUMB[906][1] ) );
  FADDER S3_906_2 ( .CIN(\ab[906][2] ), .IN0(\CARRYB[905][2] ), .IN1(
        \ab[905][3] ), .COUT(\CARRYB[906][2] ), .SUM(\SUMB[906][2] ) );
  FADDER S1_905_0 ( .CIN(\ab[905][0] ), .IN0(\CARRYB[904][0] ), .IN1(
        \SUMB[904][1] ), .COUT(\CARRYB[905][0] ), .SUM(PRODUCT[905]) );
  FADDER S2_905_1 ( .CIN(\ab[905][1] ), .IN0(\CARRYB[904][1] ), .IN1(
        \SUMB[904][2] ), .COUT(\CARRYB[905][1] ), .SUM(\SUMB[905][1] ) );
  FADDER S3_905_2 ( .CIN(\ab[905][2] ), .IN0(\CARRYB[904][2] ), .IN1(
        \ab[904][3] ), .COUT(\CARRYB[905][2] ), .SUM(\SUMB[905][2] ) );
  FADDER S1_904_0 ( .CIN(\ab[904][0] ), .IN0(\CARRYB[903][0] ), .IN1(
        \SUMB[903][1] ), .COUT(\CARRYB[904][0] ), .SUM(PRODUCT[904]) );
  FADDER S2_904_1 ( .CIN(\ab[904][1] ), .IN0(\CARRYB[903][1] ), .IN1(
        \SUMB[903][2] ), .COUT(\CARRYB[904][1] ), .SUM(\SUMB[904][1] ) );
  FADDER S3_904_2 ( .CIN(\ab[904][2] ), .IN0(\CARRYB[903][2] ), .IN1(
        \ab[903][3] ), .COUT(\CARRYB[904][2] ), .SUM(\SUMB[904][2] ) );
  FADDER S1_903_0 ( .CIN(\ab[903][0] ), .IN0(\CARRYB[902][0] ), .IN1(
        \SUMB[902][1] ), .COUT(\CARRYB[903][0] ), .SUM(PRODUCT[903]) );
  FADDER S2_903_1 ( .CIN(\ab[903][1] ), .IN0(\CARRYB[902][1] ), .IN1(
        \SUMB[902][2] ), .COUT(\CARRYB[903][1] ), .SUM(\SUMB[903][1] ) );
  FADDER S3_903_2 ( .CIN(\ab[903][2] ), .IN0(\CARRYB[902][2] ), .IN1(
        \ab[902][3] ), .COUT(\CARRYB[903][2] ), .SUM(\SUMB[903][2] ) );
  FADDER S1_902_0 ( .CIN(\ab[902][0] ), .IN0(\CARRYB[901][0] ), .IN1(
        \SUMB[901][1] ), .COUT(\CARRYB[902][0] ), .SUM(PRODUCT[902]) );
  FADDER S2_902_1 ( .CIN(\ab[902][1] ), .IN0(\CARRYB[901][1] ), .IN1(
        \SUMB[901][2] ), .COUT(\CARRYB[902][1] ), .SUM(\SUMB[902][1] ) );
  FADDER S3_902_2 ( .CIN(\ab[902][2] ), .IN0(\CARRYB[901][2] ), .IN1(
        \ab[901][3] ), .COUT(\CARRYB[902][2] ), .SUM(\SUMB[902][2] ) );
  FADDER S1_901_0 ( .CIN(\ab[901][0] ), .IN0(\CARRYB[900][0] ), .IN1(
        \SUMB[900][1] ), .COUT(\CARRYB[901][0] ), .SUM(PRODUCT[901]) );
  FADDER S2_901_1 ( .CIN(\ab[901][1] ), .IN0(\CARRYB[900][1] ), .IN1(
        \SUMB[900][2] ), .COUT(\CARRYB[901][1] ), .SUM(\SUMB[901][1] ) );
  FADDER S3_901_2 ( .CIN(\ab[901][2] ), .IN0(\CARRYB[900][2] ), .IN1(
        \ab[900][3] ), .COUT(\CARRYB[901][2] ), .SUM(\SUMB[901][2] ) );
  FADDER S1_900_0 ( .CIN(\ab[900][0] ), .IN0(\CARRYB[899][0] ), .IN1(
        \SUMB[899][1] ), .COUT(\CARRYB[900][0] ), .SUM(PRODUCT[900]) );
  FADDER S2_900_1 ( .CIN(\ab[900][1] ), .IN0(\CARRYB[899][1] ), .IN1(
        \SUMB[899][2] ), .COUT(\CARRYB[900][1] ), .SUM(\SUMB[900][1] ) );
  FADDER S3_900_2 ( .CIN(\ab[900][2] ), .IN0(\CARRYB[899][2] ), .IN1(
        \ab[899][3] ), .COUT(\CARRYB[900][2] ), .SUM(\SUMB[900][2] ) );
  FADDER S1_899_0 ( .CIN(\ab[899][0] ), .IN0(\CARRYB[898][0] ), .IN1(
        \SUMB[898][1] ), .COUT(\CARRYB[899][0] ), .SUM(PRODUCT[899]) );
  FADDER S2_899_1 ( .CIN(\ab[899][1] ), .IN0(\CARRYB[898][1] ), .IN1(
        \SUMB[898][2] ), .COUT(\CARRYB[899][1] ), .SUM(\SUMB[899][1] ) );
  FADDER S3_899_2 ( .CIN(\ab[899][2] ), .IN0(\CARRYB[898][2] ), .IN1(
        \ab[898][3] ), .COUT(\CARRYB[899][2] ), .SUM(\SUMB[899][2] ) );
  FADDER S1_898_0 ( .CIN(\ab[898][0] ), .IN0(\CARRYB[897][0] ), .IN1(
        \SUMB[897][1] ), .COUT(\CARRYB[898][0] ), .SUM(PRODUCT[898]) );
  FADDER S2_898_1 ( .CIN(\ab[898][1] ), .IN0(\CARRYB[897][1] ), .IN1(
        \SUMB[897][2] ), .COUT(\CARRYB[898][1] ), .SUM(\SUMB[898][1] ) );
  FADDER S3_898_2 ( .CIN(\ab[898][2] ), .IN0(\CARRYB[897][2] ), .IN1(
        \ab[897][3] ), .COUT(\CARRYB[898][2] ), .SUM(\SUMB[898][2] ) );
  FADDER S1_897_0 ( .CIN(\ab[897][0] ), .IN0(\CARRYB[896][0] ), .IN1(
        \SUMB[896][1] ), .COUT(\CARRYB[897][0] ), .SUM(PRODUCT[897]) );
  FADDER S2_897_1 ( .CIN(\ab[897][1] ), .IN0(\CARRYB[896][1] ), .IN1(
        \SUMB[896][2] ), .COUT(\CARRYB[897][1] ), .SUM(\SUMB[897][1] ) );
  FADDER S3_897_2 ( .CIN(\ab[897][2] ), .IN0(\CARRYB[896][2] ), .IN1(
        \ab[896][3] ), .COUT(\CARRYB[897][2] ), .SUM(\SUMB[897][2] ) );
  FADDER S1_896_0 ( .CIN(\ab[896][0] ), .IN0(\CARRYB[895][0] ), .IN1(
        \SUMB[895][1] ), .COUT(\CARRYB[896][0] ), .SUM(PRODUCT[896]) );
  FADDER S2_896_1 ( .CIN(\ab[896][1] ), .IN0(\CARRYB[895][1] ), .IN1(
        \SUMB[895][2] ), .COUT(\CARRYB[896][1] ), .SUM(\SUMB[896][1] ) );
  FADDER S3_896_2 ( .CIN(\ab[896][2] ), .IN0(\CARRYB[895][2] ), .IN1(
        \ab[895][3] ), .COUT(\CARRYB[896][2] ), .SUM(\SUMB[896][2] ) );
  FADDER S1_895_0 ( .CIN(\ab[895][0] ), .IN0(\CARRYB[894][0] ), .IN1(
        \SUMB[894][1] ), .COUT(\CARRYB[895][0] ), .SUM(PRODUCT[895]) );
  FADDER S2_895_1 ( .CIN(\ab[895][1] ), .IN0(\CARRYB[894][1] ), .IN1(
        \SUMB[894][2] ), .COUT(\CARRYB[895][1] ), .SUM(\SUMB[895][1] ) );
  FADDER S3_895_2 ( .CIN(\ab[895][2] ), .IN0(\CARRYB[894][2] ), .IN1(
        \ab[894][3] ), .COUT(\CARRYB[895][2] ), .SUM(\SUMB[895][2] ) );
  FADDER S1_894_0 ( .CIN(\ab[894][0] ), .IN0(\CARRYB[893][0] ), .IN1(
        \SUMB[893][1] ), .COUT(\CARRYB[894][0] ), .SUM(PRODUCT[894]) );
  FADDER S2_894_1 ( .CIN(\ab[894][1] ), .IN0(\CARRYB[893][1] ), .IN1(
        \SUMB[893][2] ), .COUT(\CARRYB[894][1] ), .SUM(\SUMB[894][1] ) );
  FADDER S3_894_2 ( .CIN(\ab[894][2] ), .IN0(\CARRYB[893][2] ), .IN1(
        \ab[893][3] ), .COUT(\CARRYB[894][2] ), .SUM(\SUMB[894][2] ) );
  FADDER S1_893_0 ( .CIN(\ab[893][0] ), .IN0(\CARRYB[892][0] ), .IN1(
        \SUMB[892][1] ), .COUT(\CARRYB[893][0] ), .SUM(PRODUCT[893]) );
  FADDER S2_893_1 ( .CIN(\ab[893][1] ), .IN0(\CARRYB[892][1] ), .IN1(
        \SUMB[892][2] ), .COUT(\CARRYB[893][1] ), .SUM(\SUMB[893][1] ) );
  FADDER S3_893_2 ( .CIN(\ab[893][2] ), .IN0(\CARRYB[892][2] ), .IN1(
        \ab[892][3] ), .COUT(\CARRYB[893][2] ), .SUM(\SUMB[893][2] ) );
  FADDER S1_892_0 ( .CIN(\ab[892][0] ), .IN0(\CARRYB[891][0] ), .IN1(
        \SUMB[891][1] ), .COUT(\CARRYB[892][0] ), .SUM(PRODUCT[892]) );
  FADDER S2_892_1 ( .CIN(\ab[892][1] ), .IN0(\CARRYB[891][1] ), .IN1(
        \SUMB[891][2] ), .COUT(\CARRYB[892][1] ), .SUM(\SUMB[892][1] ) );
  FADDER S3_892_2 ( .CIN(\ab[892][2] ), .IN0(\CARRYB[891][2] ), .IN1(
        \ab[891][3] ), .COUT(\CARRYB[892][2] ), .SUM(\SUMB[892][2] ) );
  FADDER S1_891_0 ( .CIN(\ab[891][0] ), .IN0(\CARRYB[890][0] ), .IN1(
        \SUMB[890][1] ), .COUT(\CARRYB[891][0] ), .SUM(PRODUCT[891]) );
  FADDER S2_891_1 ( .CIN(\ab[891][1] ), .IN0(\CARRYB[890][1] ), .IN1(
        \SUMB[890][2] ), .COUT(\CARRYB[891][1] ), .SUM(\SUMB[891][1] ) );
  FADDER S3_891_2 ( .CIN(\ab[891][2] ), .IN0(\CARRYB[890][2] ), .IN1(
        \ab[890][3] ), .COUT(\CARRYB[891][2] ), .SUM(\SUMB[891][2] ) );
  FADDER S1_890_0 ( .CIN(\ab[890][0] ), .IN0(\CARRYB[889][0] ), .IN1(
        \SUMB[889][1] ), .COUT(\CARRYB[890][0] ), .SUM(PRODUCT[890]) );
  FADDER S2_890_1 ( .CIN(\ab[890][1] ), .IN0(\CARRYB[889][1] ), .IN1(
        \SUMB[889][2] ), .COUT(\CARRYB[890][1] ), .SUM(\SUMB[890][1] ) );
  FADDER S3_890_2 ( .CIN(\ab[890][2] ), .IN0(\CARRYB[889][2] ), .IN1(
        \ab[889][3] ), .COUT(\CARRYB[890][2] ), .SUM(\SUMB[890][2] ) );
  FADDER S1_889_0 ( .CIN(\ab[889][0] ), .IN0(\CARRYB[888][0] ), .IN1(
        \SUMB[888][1] ), .COUT(\CARRYB[889][0] ), .SUM(PRODUCT[889]) );
  FADDER S2_889_1 ( .CIN(\ab[889][1] ), .IN0(\CARRYB[888][1] ), .IN1(
        \SUMB[888][2] ), .COUT(\CARRYB[889][1] ), .SUM(\SUMB[889][1] ) );
  FADDER S3_889_2 ( .CIN(\ab[889][2] ), .IN0(\CARRYB[888][2] ), .IN1(
        \ab[888][3] ), .COUT(\CARRYB[889][2] ), .SUM(\SUMB[889][2] ) );
  FADDER S1_888_0 ( .CIN(\ab[888][0] ), .IN0(\CARRYB[887][0] ), .IN1(
        \SUMB[887][1] ), .COUT(\CARRYB[888][0] ), .SUM(PRODUCT[888]) );
  FADDER S2_888_1 ( .CIN(\ab[888][1] ), .IN0(\CARRYB[887][1] ), .IN1(
        \SUMB[887][2] ), .COUT(\CARRYB[888][1] ), .SUM(\SUMB[888][1] ) );
  FADDER S3_888_2 ( .CIN(\ab[888][2] ), .IN0(\CARRYB[887][2] ), .IN1(
        \ab[887][3] ), .COUT(\CARRYB[888][2] ), .SUM(\SUMB[888][2] ) );
  FADDER S1_887_0 ( .CIN(\ab[887][0] ), .IN0(\CARRYB[886][0] ), .IN1(
        \SUMB[886][1] ), .COUT(\CARRYB[887][0] ), .SUM(PRODUCT[887]) );
  FADDER S2_887_1 ( .CIN(\ab[887][1] ), .IN0(\CARRYB[886][1] ), .IN1(
        \SUMB[886][2] ), .COUT(\CARRYB[887][1] ), .SUM(\SUMB[887][1] ) );
  FADDER S3_887_2 ( .CIN(\ab[887][2] ), .IN0(\CARRYB[886][2] ), .IN1(
        \ab[886][3] ), .COUT(\CARRYB[887][2] ), .SUM(\SUMB[887][2] ) );
  FADDER S1_886_0 ( .CIN(\ab[886][0] ), .IN0(\CARRYB[885][0] ), .IN1(
        \SUMB[885][1] ), .COUT(\CARRYB[886][0] ), .SUM(PRODUCT[886]) );
  FADDER S2_886_1 ( .CIN(\ab[886][1] ), .IN0(\CARRYB[885][1] ), .IN1(
        \SUMB[885][2] ), .COUT(\CARRYB[886][1] ), .SUM(\SUMB[886][1] ) );
  FADDER S3_886_2 ( .CIN(\ab[886][2] ), .IN0(\CARRYB[885][2] ), .IN1(
        \ab[885][3] ), .COUT(\CARRYB[886][2] ), .SUM(\SUMB[886][2] ) );
  FADDER S1_885_0 ( .CIN(\ab[885][0] ), .IN0(\CARRYB[884][0] ), .IN1(
        \SUMB[884][1] ), .COUT(\CARRYB[885][0] ), .SUM(PRODUCT[885]) );
  FADDER S2_885_1 ( .CIN(\ab[885][1] ), .IN0(\CARRYB[884][1] ), .IN1(
        \SUMB[884][2] ), .COUT(\CARRYB[885][1] ), .SUM(\SUMB[885][1] ) );
  FADDER S3_885_2 ( .CIN(\ab[885][2] ), .IN0(\CARRYB[884][2] ), .IN1(
        \ab[884][3] ), .COUT(\CARRYB[885][2] ), .SUM(\SUMB[885][2] ) );
  FADDER S1_884_0 ( .CIN(\ab[884][0] ), .IN0(\CARRYB[883][0] ), .IN1(
        \SUMB[883][1] ), .COUT(\CARRYB[884][0] ), .SUM(PRODUCT[884]) );
  FADDER S2_884_1 ( .CIN(\ab[884][1] ), .IN0(\CARRYB[883][1] ), .IN1(
        \SUMB[883][2] ), .COUT(\CARRYB[884][1] ), .SUM(\SUMB[884][1] ) );
  FADDER S3_884_2 ( .CIN(\ab[884][2] ), .IN0(\CARRYB[883][2] ), .IN1(
        \ab[883][3] ), .COUT(\CARRYB[884][2] ), .SUM(\SUMB[884][2] ) );
  FADDER S1_883_0 ( .CIN(\ab[883][0] ), .IN0(\CARRYB[882][0] ), .IN1(
        \SUMB[882][1] ), .COUT(\CARRYB[883][0] ), .SUM(PRODUCT[883]) );
  FADDER S2_883_1 ( .CIN(\ab[883][1] ), .IN0(\CARRYB[882][1] ), .IN1(
        \SUMB[882][2] ), .COUT(\CARRYB[883][1] ), .SUM(\SUMB[883][1] ) );
  FADDER S3_883_2 ( .CIN(\ab[883][2] ), .IN0(\CARRYB[882][2] ), .IN1(
        \ab[882][3] ), .COUT(\CARRYB[883][2] ), .SUM(\SUMB[883][2] ) );
  FADDER S1_882_0 ( .CIN(\ab[882][0] ), .IN0(\CARRYB[881][0] ), .IN1(
        \SUMB[881][1] ), .COUT(\CARRYB[882][0] ), .SUM(PRODUCT[882]) );
  FADDER S2_882_1 ( .CIN(\ab[882][1] ), .IN0(\CARRYB[881][1] ), .IN1(
        \SUMB[881][2] ), .COUT(\CARRYB[882][1] ), .SUM(\SUMB[882][1] ) );
  FADDER S3_882_2 ( .CIN(\ab[882][2] ), .IN0(\CARRYB[881][2] ), .IN1(
        \ab[881][3] ), .COUT(\CARRYB[882][2] ), .SUM(\SUMB[882][2] ) );
  FADDER S1_881_0 ( .CIN(\ab[881][0] ), .IN0(\CARRYB[880][0] ), .IN1(
        \SUMB[880][1] ), .COUT(\CARRYB[881][0] ), .SUM(PRODUCT[881]) );
  FADDER S2_881_1 ( .CIN(\ab[881][1] ), .IN0(\CARRYB[880][1] ), .IN1(
        \SUMB[880][2] ), .COUT(\CARRYB[881][1] ), .SUM(\SUMB[881][1] ) );
  FADDER S3_881_2 ( .CIN(\ab[881][2] ), .IN0(\CARRYB[880][2] ), .IN1(
        \ab[880][3] ), .COUT(\CARRYB[881][2] ), .SUM(\SUMB[881][2] ) );
  FADDER S1_880_0 ( .CIN(\ab[880][0] ), .IN0(\CARRYB[879][0] ), .IN1(
        \SUMB[879][1] ), .COUT(\CARRYB[880][0] ), .SUM(PRODUCT[880]) );
  FADDER S2_880_1 ( .CIN(\ab[880][1] ), .IN0(\CARRYB[879][1] ), .IN1(
        \SUMB[879][2] ), .COUT(\CARRYB[880][1] ), .SUM(\SUMB[880][1] ) );
  FADDER S3_880_2 ( .CIN(\ab[880][2] ), .IN0(\CARRYB[879][2] ), .IN1(
        \ab[879][3] ), .COUT(\CARRYB[880][2] ), .SUM(\SUMB[880][2] ) );
  FADDER S1_879_0 ( .CIN(\ab[879][0] ), .IN0(\CARRYB[878][0] ), .IN1(
        \SUMB[878][1] ), .COUT(\CARRYB[879][0] ), .SUM(PRODUCT[879]) );
  FADDER S2_879_1 ( .CIN(\ab[879][1] ), .IN0(\CARRYB[878][1] ), .IN1(
        \SUMB[878][2] ), .COUT(\CARRYB[879][1] ), .SUM(\SUMB[879][1] ) );
  FADDER S3_879_2 ( .CIN(\ab[879][2] ), .IN0(\CARRYB[878][2] ), .IN1(
        \ab[878][3] ), .COUT(\CARRYB[879][2] ), .SUM(\SUMB[879][2] ) );
  FADDER S1_878_0 ( .CIN(\ab[878][0] ), .IN0(\CARRYB[877][0] ), .IN1(
        \SUMB[877][1] ), .COUT(\CARRYB[878][0] ), .SUM(PRODUCT[878]) );
  FADDER S2_878_1 ( .CIN(\ab[878][1] ), .IN0(\CARRYB[877][1] ), .IN1(
        \SUMB[877][2] ), .COUT(\CARRYB[878][1] ), .SUM(\SUMB[878][1] ) );
  FADDER S3_878_2 ( .CIN(\ab[878][2] ), .IN0(\CARRYB[877][2] ), .IN1(
        \ab[877][3] ), .COUT(\CARRYB[878][2] ), .SUM(\SUMB[878][2] ) );
  FADDER S1_877_0 ( .CIN(\ab[877][0] ), .IN0(\CARRYB[876][0] ), .IN1(
        \SUMB[876][1] ), .COUT(\CARRYB[877][0] ), .SUM(PRODUCT[877]) );
  FADDER S2_877_1 ( .CIN(\ab[877][1] ), .IN0(\CARRYB[876][1] ), .IN1(
        \SUMB[876][2] ), .COUT(\CARRYB[877][1] ), .SUM(\SUMB[877][1] ) );
  FADDER S3_877_2 ( .CIN(\ab[877][2] ), .IN0(\CARRYB[876][2] ), .IN1(
        \ab[876][3] ), .COUT(\CARRYB[877][2] ), .SUM(\SUMB[877][2] ) );
  FADDER S1_876_0 ( .CIN(\ab[876][0] ), .IN0(\CARRYB[875][0] ), .IN1(
        \SUMB[875][1] ), .COUT(\CARRYB[876][0] ), .SUM(PRODUCT[876]) );
  FADDER S2_876_1 ( .CIN(\ab[876][1] ), .IN0(\CARRYB[875][1] ), .IN1(
        \SUMB[875][2] ), .COUT(\CARRYB[876][1] ), .SUM(\SUMB[876][1] ) );
  FADDER S3_876_2 ( .CIN(\ab[876][2] ), .IN0(\CARRYB[875][2] ), .IN1(
        \ab[875][3] ), .COUT(\CARRYB[876][2] ), .SUM(\SUMB[876][2] ) );
  FADDER S1_875_0 ( .CIN(\ab[875][0] ), .IN0(\CARRYB[874][0] ), .IN1(
        \SUMB[874][1] ), .COUT(\CARRYB[875][0] ), .SUM(PRODUCT[875]) );
  FADDER S2_875_1 ( .CIN(\ab[875][1] ), .IN0(\CARRYB[874][1] ), .IN1(
        \SUMB[874][2] ), .COUT(\CARRYB[875][1] ), .SUM(\SUMB[875][1] ) );
  FADDER S3_875_2 ( .CIN(\ab[875][2] ), .IN0(\CARRYB[874][2] ), .IN1(
        \ab[874][3] ), .COUT(\CARRYB[875][2] ), .SUM(\SUMB[875][2] ) );
  FADDER S1_874_0 ( .CIN(\ab[874][0] ), .IN0(\CARRYB[873][0] ), .IN1(
        \SUMB[873][1] ), .COUT(\CARRYB[874][0] ), .SUM(PRODUCT[874]) );
  FADDER S2_874_1 ( .CIN(\ab[874][1] ), .IN0(\CARRYB[873][1] ), .IN1(
        \SUMB[873][2] ), .COUT(\CARRYB[874][1] ), .SUM(\SUMB[874][1] ) );
  FADDER S3_874_2 ( .CIN(\ab[874][2] ), .IN0(\CARRYB[873][2] ), .IN1(
        \ab[873][3] ), .COUT(\CARRYB[874][2] ), .SUM(\SUMB[874][2] ) );
  FADDER S1_873_0 ( .CIN(\ab[873][0] ), .IN0(\CARRYB[872][0] ), .IN1(
        \SUMB[872][1] ), .COUT(\CARRYB[873][0] ), .SUM(PRODUCT[873]) );
  FADDER S2_873_1 ( .CIN(\ab[873][1] ), .IN0(\CARRYB[872][1] ), .IN1(
        \SUMB[872][2] ), .COUT(\CARRYB[873][1] ), .SUM(\SUMB[873][1] ) );
  FADDER S3_873_2 ( .CIN(\ab[873][2] ), .IN0(\CARRYB[872][2] ), .IN1(
        \ab[872][3] ), .COUT(\CARRYB[873][2] ), .SUM(\SUMB[873][2] ) );
  FADDER S1_872_0 ( .CIN(\ab[872][0] ), .IN0(\CARRYB[871][0] ), .IN1(
        \SUMB[871][1] ), .COUT(\CARRYB[872][0] ), .SUM(PRODUCT[872]) );
  FADDER S2_872_1 ( .CIN(\ab[872][1] ), .IN0(\CARRYB[871][1] ), .IN1(
        \SUMB[871][2] ), .COUT(\CARRYB[872][1] ), .SUM(\SUMB[872][1] ) );
  FADDER S3_872_2 ( .CIN(\ab[872][2] ), .IN0(\CARRYB[871][2] ), .IN1(
        \ab[871][3] ), .COUT(\CARRYB[872][2] ), .SUM(\SUMB[872][2] ) );
  FADDER S1_871_0 ( .CIN(\ab[871][0] ), .IN0(\CARRYB[870][0] ), .IN1(
        \SUMB[870][1] ), .COUT(\CARRYB[871][0] ), .SUM(PRODUCT[871]) );
  FADDER S2_871_1 ( .CIN(\ab[871][1] ), .IN0(\CARRYB[870][1] ), .IN1(
        \SUMB[870][2] ), .COUT(\CARRYB[871][1] ), .SUM(\SUMB[871][1] ) );
  FADDER S3_871_2 ( .CIN(\ab[871][2] ), .IN0(\CARRYB[870][2] ), .IN1(
        \ab[870][3] ), .COUT(\CARRYB[871][2] ), .SUM(\SUMB[871][2] ) );
  FADDER S1_870_0 ( .CIN(\ab[870][0] ), .IN0(\CARRYB[869][0] ), .IN1(
        \SUMB[869][1] ), .COUT(\CARRYB[870][0] ), .SUM(PRODUCT[870]) );
  FADDER S2_870_1 ( .CIN(\ab[870][1] ), .IN0(\CARRYB[869][1] ), .IN1(
        \SUMB[869][2] ), .COUT(\CARRYB[870][1] ), .SUM(\SUMB[870][1] ) );
  FADDER S3_870_2 ( .CIN(\ab[870][2] ), .IN0(\CARRYB[869][2] ), .IN1(
        \ab[869][3] ), .COUT(\CARRYB[870][2] ), .SUM(\SUMB[870][2] ) );
  FADDER S1_869_0 ( .CIN(\ab[869][0] ), .IN0(\CARRYB[868][0] ), .IN1(
        \SUMB[868][1] ), .COUT(\CARRYB[869][0] ), .SUM(PRODUCT[869]) );
  FADDER S2_869_1 ( .CIN(\ab[869][1] ), .IN0(\CARRYB[868][1] ), .IN1(
        \SUMB[868][2] ), .COUT(\CARRYB[869][1] ), .SUM(\SUMB[869][1] ) );
  FADDER S3_869_2 ( .CIN(\ab[869][2] ), .IN0(\CARRYB[868][2] ), .IN1(
        \ab[868][3] ), .COUT(\CARRYB[869][2] ), .SUM(\SUMB[869][2] ) );
  FADDER S1_868_0 ( .CIN(\ab[868][0] ), .IN0(\CARRYB[867][0] ), .IN1(
        \SUMB[867][1] ), .COUT(\CARRYB[868][0] ), .SUM(PRODUCT[868]) );
  FADDER S2_868_1 ( .CIN(\ab[868][1] ), .IN0(\CARRYB[867][1] ), .IN1(
        \SUMB[867][2] ), .COUT(\CARRYB[868][1] ), .SUM(\SUMB[868][1] ) );
  FADDER S3_868_2 ( .CIN(\ab[868][2] ), .IN0(\CARRYB[867][2] ), .IN1(
        \ab[867][3] ), .COUT(\CARRYB[868][2] ), .SUM(\SUMB[868][2] ) );
  FADDER S1_867_0 ( .CIN(\ab[867][0] ), .IN0(\CARRYB[866][0] ), .IN1(
        \SUMB[866][1] ), .COUT(\CARRYB[867][0] ), .SUM(PRODUCT[867]) );
  FADDER S2_867_1 ( .CIN(\ab[867][1] ), .IN0(\CARRYB[866][1] ), .IN1(
        \SUMB[866][2] ), .COUT(\CARRYB[867][1] ), .SUM(\SUMB[867][1] ) );
  FADDER S3_867_2 ( .CIN(\ab[867][2] ), .IN0(\CARRYB[866][2] ), .IN1(
        \ab[866][3] ), .COUT(\CARRYB[867][2] ), .SUM(\SUMB[867][2] ) );
  FADDER S1_866_0 ( .CIN(\ab[866][0] ), .IN0(\CARRYB[865][0] ), .IN1(
        \SUMB[865][1] ), .COUT(\CARRYB[866][0] ), .SUM(PRODUCT[866]) );
  FADDER S2_866_1 ( .CIN(\ab[866][1] ), .IN0(\CARRYB[865][1] ), .IN1(
        \SUMB[865][2] ), .COUT(\CARRYB[866][1] ), .SUM(\SUMB[866][1] ) );
  FADDER S3_866_2 ( .CIN(\ab[866][2] ), .IN0(\CARRYB[865][2] ), .IN1(
        \ab[865][3] ), .COUT(\CARRYB[866][2] ), .SUM(\SUMB[866][2] ) );
  FADDER S1_865_0 ( .CIN(\ab[865][0] ), .IN0(\CARRYB[864][0] ), .IN1(
        \SUMB[864][1] ), .COUT(\CARRYB[865][0] ), .SUM(PRODUCT[865]) );
  FADDER S2_865_1 ( .CIN(\ab[865][1] ), .IN0(\CARRYB[864][1] ), .IN1(
        \SUMB[864][2] ), .COUT(\CARRYB[865][1] ), .SUM(\SUMB[865][1] ) );
  FADDER S3_865_2 ( .CIN(\ab[865][2] ), .IN0(\CARRYB[864][2] ), .IN1(
        \ab[864][3] ), .COUT(\CARRYB[865][2] ), .SUM(\SUMB[865][2] ) );
  FADDER S1_864_0 ( .CIN(\ab[864][0] ), .IN0(\CARRYB[863][0] ), .IN1(
        \SUMB[863][1] ), .COUT(\CARRYB[864][0] ), .SUM(PRODUCT[864]) );
  FADDER S2_864_1 ( .CIN(\ab[864][1] ), .IN0(\CARRYB[863][1] ), .IN1(
        \SUMB[863][2] ), .COUT(\CARRYB[864][1] ), .SUM(\SUMB[864][1] ) );
  FADDER S3_864_2 ( .CIN(\ab[864][2] ), .IN0(\CARRYB[863][2] ), .IN1(
        \ab[863][3] ), .COUT(\CARRYB[864][2] ), .SUM(\SUMB[864][2] ) );
  FADDER S1_863_0 ( .CIN(\ab[863][0] ), .IN0(\CARRYB[862][0] ), .IN1(
        \SUMB[862][1] ), .COUT(\CARRYB[863][0] ), .SUM(PRODUCT[863]) );
  FADDER S2_863_1 ( .CIN(\ab[863][1] ), .IN0(\CARRYB[862][1] ), .IN1(
        \SUMB[862][2] ), .COUT(\CARRYB[863][1] ), .SUM(\SUMB[863][1] ) );
  FADDER S3_863_2 ( .CIN(\ab[863][2] ), .IN0(\CARRYB[862][2] ), .IN1(
        \ab[862][3] ), .COUT(\CARRYB[863][2] ), .SUM(\SUMB[863][2] ) );
  FADDER S1_862_0 ( .CIN(\ab[862][0] ), .IN0(\CARRYB[861][0] ), .IN1(
        \SUMB[861][1] ), .COUT(\CARRYB[862][0] ), .SUM(PRODUCT[862]) );
  FADDER S2_862_1 ( .CIN(\ab[862][1] ), .IN0(\CARRYB[861][1] ), .IN1(
        \SUMB[861][2] ), .COUT(\CARRYB[862][1] ), .SUM(\SUMB[862][1] ) );
  FADDER S3_862_2 ( .CIN(\ab[862][2] ), .IN0(\CARRYB[861][2] ), .IN1(
        \ab[861][3] ), .COUT(\CARRYB[862][2] ), .SUM(\SUMB[862][2] ) );
  FADDER S1_861_0 ( .CIN(\ab[861][0] ), .IN0(\CARRYB[860][0] ), .IN1(
        \SUMB[860][1] ), .COUT(\CARRYB[861][0] ), .SUM(PRODUCT[861]) );
  FADDER S2_861_1 ( .CIN(\ab[861][1] ), .IN0(\CARRYB[860][1] ), .IN1(
        \SUMB[860][2] ), .COUT(\CARRYB[861][1] ), .SUM(\SUMB[861][1] ) );
  FADDER S3_861_2 ( .CIN(\ab[861][2] ), .IN0(\CARRYB[860][2] ), .IN1(
        \ab[860][3] ), .COUT(\CARRYB[861][2] ), .SUM(\SUMB[861][2] ) );
  FADDER S1_860_0 ( .CIN(\ab[860][0] ), .IN0(\CARRYB[859][0] ), .IN1(
        \SUMB[859][1] ), .COUT(\CARRYB[860][0] ), .SUM(PRODUCT[860]) );
  FADDER S2_860_1 ( .CIN(\ab[860][1] ), .IN0(\CARRYB[859][1] ), .IN1(
        \SUMB[859][2] ), .COUT(\CARRYB[860][1] ), .SUM(\SUMB[860][1] ) );
  FADDER S3_860_2 ( .CIN(\ab[860][2] ), .IN0(\CARRYB[859][2] ), .IN1(
        \ab[859][3] ), .COUT(\CARRYB[860][2] ), .SUM(\SUMB[860][2] ) );
  FADDER S1_859_0 ( .CIN(\ab[859][0] ), .IN0(\CARRYB[858][0] ), .IN1(
        \SUMB[858][1] ), .COUT(\CARRYB[859][0] ), .SUM(PRODUCT[859]) );
  FADDER S2_859_1 ( .CIN(\ab[859][1] ), .IN0(\CARRYB[858][1] ), .IN1(
        \SUMB[858][2] ), .COUT(\CARRYB[859][1] ), .SUM(\SUMB[859][1] ) );
  FADDER S3_859_2 ( .CIN(\ab[859][2] ), .IN0(\CARRYB[858][2] ), .IN1(
        \ab[858][3] ), .COUT(\CARRYB[859][2] ), .SUM(\SUMB[859][2] ) );
  FADDER S1_858_0 ( .CIN(\ab[858][0] ), .IN0(\CARRYB[857][0] ), .IN1(
        \SUMB[857][1] ), .COUT(\CARRYB[858][0] ), .SUM(PRODUCT[858]) );
  FADDER S2_858_1 ( .CIN(\ab[858][1] ), .IN0(\CARRYB[857][1] ), .IN1(
        \SUMB[857][2] ), .COUT(\CARRYB[858][1] ), .SUM(\SUMB[858][1] ) );
  FADDER S3_858_2 ( .CIN(\ab[858][2] ), .IN0(\CARRYB[857][2] ), .IN1(
        \ab[857][3] ), .COUT(\CARRYB[858][2] ), .SUM(\SUMB[858][2] ) );
  FADDER S1_857_0 ( .CIN(\ab[857][0] ), .IN0(\CARRYB[856][0] ), .IN1(
        \SUMB[856][1] ), .COUT(\CARRYB[857][0] ), .SUM(PRODUCT[857]) );
  FADDER S2_857_1 ( .CIN(\ab[857][1] ), .IN0(\CARRYB[856][1] ), .IN1(
        \SUMB[856][2] ), .COUT(\CARRYB[857][1] ), .SUM(\SUMB[857][1] ) );
  FADDER S3_857_2 ( .CIN(\ab[857][2] ), .IN0(\CARRYB[856][2] ), .IN1(
        \ab[856][3] ), .COUT(\CARRYB[857][2] ), .SUM(\SUMB[857][2] ) );
  FADDER S1_856_0 ( .CIN(\ab[856][0] ), .IN0(\CARRYB[855][0] ), .IN1(
        \SUMB[855][1] ), .COUT(\CARRYB[856][0] ), .SUM(PRODUCT[856]) );
  FADDER S2_856_1 ( .CIN(\ab[856][1] ), .IN0(\CARRYB[855][1] ), .IN1(
        \SUMB[855][2] ), .COUT(\CARRYB[856][1] ), .SUM(\SUMB[856][1] ) );
  FADDER S3_856_2 ( .CIN(\ab[856][2] ), .IN0(\CARRYB[855][2] ), .IN1(
        \ab[855][3] ), .COUT(\CARRYB[856][2] ), .SUM(\SUMB[856][2] ) );
  FADDER S1_855_0 ( .CIN(\ab[855][0] ), .IN0(\CARRYB[854][0] ), .IN1(
        \SUMB[854][1] ), .COUT(\CARRYB[855][0] ), .SUM(PRODUCT[855]) );
  FADDER S2_855_1 ( .CIN(\ab[855][1] ), .IN0(\CARRYB[854][1] ), .IN1(
        \SUMB[854][2] ), .COUT(\CARRYB[855][1] ), .SUM(\SUMB[855][1] ) );
  FADDER S3_855_2 ( .CIN(\ab[855][2] ), .IN0(\CARRYB[854][2] ), .IN1(
        \ab[854][3] ), .COUT(\CARRYB[855][2] ), .SUM(\SUMB[855][2] ) );
  FADDER S1_854_0 ( .CIN(\ab[854][0] ), .IN0(\CARRYB[853][0] ), .IN1(
        \SUMB[853][1] ), .COUT(\CARRYB[854][0] ), .SUM(PRODUCT[854]) );
  FADDER S2_854_1 ( .CIN(\ab[854][1] ), .IN0(\CARRYB[853][1] ), .IN1(
        \SUMB[853][2] ), .COUT(\CARRYB[854][1] ), .SUM(\SUMB[854][1] ) );
  FADDER S3_854_2 ( .CIN(\ab[854][2] ), .IN0(\CARRYB[853][2] ), .IN1(
        \ab[853][3] ), .COUT(\CARRYB[854][2] ), .SUM(\SUMB[854][2] ) );
  FADDER S1_853_0 ( .CIN(\ab[853][0] ), .IN0(\CARRYB[852][0] ), .IN1(
        \SUMB[852][1] ), .COUT(\CARRYB[853][0] ), .SUM(PRODUCT[853]) );
  FADDER S2_853_1 ( .CIN(\ab[853][1] ), .IN0(\CARRYB[852][1] ), .IN1(
        \SUMB[852][2] ), .COUT(\CARRYB[853][1] ), .SUM(\SUMB[853][1] ) );
  FADDER S3_853_2 ( .CIN(\ab[853][2] ), .IN0(\CARRYB[852][2] ), .IN1(
        \ab[852][3] ), .COUT(\CARRYB[853][2] ), .SUM(\SUMB[853][2] ) );
  FADDER S1_852_0 ( .CIN(\ab[852][0] ), .IN0(\CARRYB[851][0] ), .IN1(
        \SUMB[851][1] ), .COUT(\CARRYB[852][0] ), .SUM(PRODUCT[852]) );
  FADDER S2_852_1 ( .CIN(\ab[852][1] ), .IN0(\CARRYB[851][1] ), .IN1(
        \SUMB[851][2] ), .COUT(\CARRYB[852][1] ), .SUM(\SUMB[852][1] ) );
  FADDER S3_852_2 ( .CIN(\ab[852][2] ), .IN0(\CARRYB[851][2] ), .IN1(
        \ab[851][3] ), .COUT(\CARRYB[852][2] ), .SUM(\SUMB[852][2] ) );
  FADDER S1_851_0 ( .CIN(\ab[851][0] ), .IN0(\CARRYB[850][0] ), .IN1(
        \SUMB[850][1] ), .COUT(\CARRYB[851][0] ), .SUM(PRODUCT[851]) );
  FADDER S2_851_1 ( .CIN(\ab[851][1] ), .IN0(\CARRYB[850][1] ), .IN1(
        \SUMB[850][2] ), .COUT(\CARRYB[851][1] ), .SUM(\SUMB[851][1] ) );
  FADDER S3_851_2 ( .CIN(\ab[851][2] ), .IN0(\CARRYB[850][2] ), .IN1(
        \ab[850][3] ), .COUT(\CARRYB[851][2] ), .SUM(\SUMB[851][2] ) );
  FADDER S1_850_0 ( .CIN(\ab[850][0] ), .IN0(\CARRYB[849][0] ), .IN1(
        \SUMB[849][1] ), .COUT(\CARRYB[850][0] ), .SUM(PRODUCT[850]) );
  FADDER S2_850_1 ( .CIN(\ab[850][1] ), .IN0(\CARRYB[849][1] ), .IN1(
        \SUMB[849][2] ), .COUT(\CARRYB[850][1] ), .SUM(\SUMB[850][1] ) );
  FADDER S3_850_2 ( .CIN(\ab[850][2] ), .IN0(\CARRYB[849][2] ), .IN1(
        \ab[849][3] ), .COUT(\CARRYB[850][2] ), .SUM(\SUMB[850][2] ) );
  FADDER S1_849_0 ( .CIN(\ab[849][0] ), .IN0(\CARRYB[848][0] ), .IN1(
        \SUMB[848][1] ), .COUT(\CARRYB[849][0] ), .SUM(PRODUCT[849]) );
  FADDER S2_849_1 ( .CIN(\ab[849][1] ), .IN0(\CARRYB[848][1] ), .IN1(
        \SUMB[848][2] ), .COUT(\CARRYB[849][1] ), .SUM(\SUMB[849][1] ) );
  FADDER S3_849_2 ( .CIN(\ab[849][2] ), .IN0(\CARRYB[848][2] ), .IN1(
        \ab[848][3] ), .COUT(\CARRYB[849][2] ), .SUM(\SUMB[849][2] ) );
  FADDER S1_848_0 ( .CIN(\ab[848][0] ), .IN0(\CARRYB[847][0] ), .IN1(
        \SUMB[847][1] ), .COUT(\CARRYB[848][0] ), .SUM(PRODUCT[848]) );
  FADDER S2_848_1 ( .CIN(\ab[848][1] ), .IN0(\CARRYB[847][1] ), .IN1(
        \SUMB[847][2] ), .COUT(\CARRYB[848][1] ), .SUM(\SUMB[848][1] ) );
  FADDER S3_848_2 ( .CIN(\ab[848][2] ), .IN0(\CARRYB[847][2] ), .IN1(
        \ab[847][3] ), .COUT(\CARRYB[848][2] ), .SUM(\SUMB[848][2] ) );
  FADDER S1_847_0 ( .CIN(\ab[847][0] ), .IN0(\CARRYB[846][0] ), .IN1(
        \SUMB[846][1] ), .COUT(\CARRYB[847][0] ), .SUM(PRODUCT[847]) );
  FADDER S2_847_1 ( .CIN(\ab[847][1] ), .IN0(\CARRYB[846][1] ), .IN1(
        \SUMB[846][2] ), .COUT(\CARRYB[847][1] ), .SUM(\SUMB[847][1] ) );
  FADDER S3_847_2 ( .CIN(\ab[847][2] ), .IN0(\CARRYB[846][2] ), .IN1(
        \ab[846][3] ), .COUT(\CARRYB[847][2] ), .SUM(\SUMB[847][2] ) );
  FADDER S1_846_0 ( .CIN(\ab[846][0] ), .IN0(\CARRYB[845][0] ), .IN1(
        \SUMB[845][1] ), .COUT(\CARRYB[846][0] ), .SUM(PRODUCT[846]) );
  FADDER S2_846_1 ( .CIN(\ab[846][1] ), .IN0(\CARRYB[845][1] ), .IN1(
        \SUMB[845][2] ), .COUT(\CARRYB[846][1] ), .SUM(\SUMB[846][1] ) );
  FADDER S3_846_2 ( .CIN(\ab[846][2] ), .IN0(\CARRYB[845][2] ), .IN1(
        \ab[845][3] ), .COUT(\CARRYB[846][2] ), .SUM(\SUMB[846][2] ) );
  FADDER S1_845_0 ( .CIN(\ab[845][0] ), .IN0(\CARRYB[844][0] ), .IN1(
        \SUMB[844][1] ), .COUT(\CARRYB[845][0] ), .SUM(PRODUCT[845]) );
  FADDER S2_845_1 ( .CIN(\ab[845][1] ), .IN0(\CARRYB[844][1] ), .IN1(
        \SUMB[844][2] ), .COUT(\CARRYB[845][1] ), .SUM(\SUMB[845][1] ) );
  FADDER S3_845_2 ( .CIN(\ab[845][2] ), .IN0(\CARRYB[844][2] ), .IN1(
        \ab[844][3] ), .COUT(\CARRYB[845][2] ), .SUM(\SUMB[845][2] ) );
  FADDER S1_844_0 ( .CIN(\ab[844][0] ), .IN0(\CARRYB[843][0] ), .IN1(
        \SUMB[843][1] ), .COUT(\CARRYB[844][0] ), .SUM(PRODUCT[844]) );
  FADDER S2_844_1 ( .CIN(\ab[844][1] ), .IN0(\CARRYB[843][1] ), .IN1(
        \SUMB[843][2] ), .COUT(\CARRYB[844][1] ), .SUM(\SUMB[844][1] ) );
  FADDER S3_844_2 ( .CIN(\ab[844][2] ), .IN0(\CARRYB[843][2] ), .IN1(
        \ab[843][3] ), .COUT(\CARRYB[844][2] ), .SUM(\SUMB[844][2] ) );
  FADDER S1_843_0 ( .CIN(\ab[843][0] ), .IN0(\CARRYB[842][0] ), .IN1(
        \SUMB[842][1] ), .COUT(\CARRYB[843][0] ), .SUM(PRODUCT[843]) );
  FADDER S2_843_1 ( .CIN(\ab[843][1] ), .IN0(\CARRYB[842][1] ), .IN1(
        \SUMB[842][2] ), .COUT(\CARRYB[843][1] ), .SUM(\SUMB[843][1] ) );
  FADDER S3_843_2 ( .CIN(\ab[843][2] ), .IN0(\CARRYB[842][2] ), .IN1(
        \ab[842][3] ), .COUT(\CARRYB[843][2] ), .SUM(\SUMB[843][2] ) );
  FADDER S1_842_0 ( .CIN(\ab[842][0] ), .IN0(\CARRYB[841][0] ), .IN1(
        \SUMB[841][1] ), .COUT(\CARRYB[842][0] ), .SUM(PRODUCT[842]) );
  FADDER S2_842_1 ( .CIN(\ab[842][1] ), .IN0(\CARRYB[841][1] ), .IN1(
        \SUMB[841][2] ), .COUT(\CARRYB[842][1] ), .SUM(\SUMB[842][1] ) );
  FADDER S3_842_2 ( .CIN(\ab[842][2] ), .IN0(\CARRYB[841][2] ), .IN1(
        \ab[841][3] ), .COUT(\CARRYB[842][2] ), .SUM(\SUMB[842][2] ) );
  FADDER S1_841_0 ( .CIN(\ab[841][0] ), .IN0(\CARRYB[840][0] ), .IN1(
        \SUMB[840][1] ), .COUT(\CARRYB[841][0] ), .SUM(PRODUCT[841]) );
  FADDER S2_841_1 ( .CIN(\ab[841][1] ), .IN0(\CARRYB[840][1] ), .IN1(
        \SUMB[840][2] ), .COUT(\CARRYB[841][1] ), .SUM(\SUMB[841][1] ) );
  FADDER S3_841_2 ( .CIN(\ab[841][2] ), .IN0(\CARRYB[840][2] ), .IN1(
        \ab[840][3] ), .COUT(\CARRYB[841][2] ), .SUM(\SUMB[841][2] ) );
  FADDER S1_840_0 ( .CIN(\ab[840][0] ), .IN0(\CARRYB[839][0] ), .IN1(
        \SUMB[839][1] ), .COUT(\CARRYB[840][0] ), .SUM(PRODUCT[840]) );
  FADDER S2_840_1 ( .CIN(\ab[840][1] ), .IN0(\CARRYB[839][1] ), .IN1(
        \SUMB[839][2] ), .COUT(\CARRYB[840][1] ), .SUM(\SUMB[840][1] ) );
  FADDER S3_840_2 ( .CIN(\ab[840][2] ), .IN0(\CARRYB[839][2] ), .IN1(
        \ab[839][3] ), .COUT(\CARRYB[840][2] ), .SUM(\SUMB[840][2] ) );
  FADDER S1_839_0 ( .CIN(\ab[839][0] ), .IN0(\CARRYB[838][0] ), .IN1(
        \SUMB[838][1] ), .COUT(\CARRYB[839][0] ), .SUM(PRODUCT[839]) );
  FADDER S2_839_1 ( .CIN(\ab[839][1] ), .IN0(\CARRYB[838][1] ), .IN1(
        \SUMB[838][2] ), .COUT(\CARRYB[839][1] ), .SUM(\SUMB[839][1] ) );
  FADDER S3_839_2 ( .CIN(\ab[839][2] ), .IN0(\CARRYB[838][2] ), .IN1(
        \ab[838][3] ), .COUT(\CARRYB[839][2] ), .SUM(\SUMB[839][2] ) );
  FADDER S1_838_0 ( .CIN(\ab[838][0] ), .IN0(\CARRYB[837][0] ), .IN1(
        \SUMB[837][1] ), .COUT(\CARRYB[838][0] ), .SUM(PRODUCT[838]) );
  FADDER S2_838_1 ( .CIN(\ab[838][1] ), .IN0(\CARRYB[837][1] ), .IN1(
        \SUMB[837][2] ), .COUT(\CARRYB[838][1] ), .SUM(\SUMB[838][1] ) );
  FADDER S3_838_2 ( .CIN(\ab[838][2] ), .IN0(\CARRYB[837][2] ), .IN1(
        \ab[837][3] ), .COUT(\CARRYB[838][2] ), .SUM(\SUMB[838][2] ) );
  FADDER S1_837_0 ( .CIN(\ab[837][0] ), .IN0(\CARRYB[836][0] ), .IN1(
        \SUMB[836][1] ), .COUT(\CARRYB[837][0] ), .SUM(PRODUCT[837]) );
  FADDER S2_837_1 ( .CIN(\ab[837][1] ), .IN0(\CARRYB[836][1] ), .IN1(
        \SUMB[836][2] ), .COUT(\CARRYB[837][1] ), .SUM(\SUMB[837][1] ) );
  FADDER S3_837_2 ( .CIN(\ab[837][2] ), .IN0(\CARRYB[836][2] ), .IN1(
        \ab[836][3] ), .COUT(\CARRYB[837][2] ), .SUM(\SUMB[837][2] ) );
  FADDER S1_836_0 ( .CIN(\ab[836][0] ), .IN0(\CARRYB[835][0] ), .IN1(
        \SUMB[835][1] ), .COUT(\CARRYB[836][0] ), .SUM(PRODUCT[836]) );
  FADDER S2_836_1 ( .CIN(\ab[836][1] ), .IN0(\CARRYB[835][1] ), .IN1(
        \SUMB[835][2] ), .COUT(\CARRYB[836][1] ), .SUM(\SUMB[836][1] ) );
  FADDER S3_836_2 ( .CIN(\ab[836][2] ), .IN0(\CARRYB[835][2] ), .IN1(
        \ab[835][3] ), .COUT(\CARRYB[836][2] ), .SUM(\SUMB[836][2] ) );
  FADDER S1_835_0 ( .CIN(\ab[835][0] ), .IN0(\CARRYB[834][0] ), .IN1(
        \SUMB[834][1] ), .COUT(\CARRYB[835][0] ), .SUM(PRODUCT[835]) );
  FADDER S2_835_1 ( .CIN(\ab[835][1] ), .IN0(\CARRYB[834][1] ), .IN1(
        \SUMB[834][2] ), .COUT(\CARRYB[835][1] ), .SUM(\SUMB[835][1] ) );
  FADDER S3_835_2 ( .CIN(\ab[835][2] ), .IN0(\CARRYB[834][2] ), .IN1(
        \ab[834][3] ), .COUT(\CARRYB[835][2] ), .SUM(\SUMB[835][2] ) );
  FADDER S1_834_0 ( .CIN(\ab[834][0] ), .IN0(\CARRYB[833][0] ), .IN1(
        \SUMB[833][1] ), .COUT(\CARRYB[834][0] ), .SUM(PRODUCT[834]) );
  FADDER S2_834_1 ( .CIN(\ab[834][1] ), .IN0(\CARRYB[833][1] ), .IN1(
        \SUMB[833][2] ), .COUT(\CARRYB[834][1] ), .SUM(\SUMB[834][1] ) );
  FADDER S3_834_2 ( .CIN(\ab[834][2] ), .IN0(\CARRYB[833][2] ), .IN1(
        \ab[833][3] ), .COUT(\CARRYB[834][2] ), .SUM(\SUMB[834][2] ) );
  FADDER S1_833_0 ( .CIN(\ab[833][0] ), .IN0(\CARRYB[832][0] ), .IN1(
        \SUMB[832][1] ), .COUT(\CARRYB[833][0] ), .SUM(PRODUCT[833]) );
  FADDER S2_833_1 ( .CIN(\ab[833][1] ), .IN0(\CARRYB[832][1] ), .IN1(
        \SUMB[832][2] ), .COUT(\CARRYB[833][1] ), .SUM(\SUMB[833][1] ) );
  FADDER S3_833_2 ( .CIN(\ab[833][2] ), .IN0(\CARRYB[832][2] ), .IN1(
        \ab[832][3] ), .COUT(\CARRYB[833][2] ), .SUM(\SUMB[833][2] ) );
  FADDER S1_832_0 ( .CIN(\ab[832][0] ), .IN0(\CARRYB[831][0] ), .IN1(
        \SUMB[831][1] ), .COUT(\CARRYB[832][0] ), .SUM(PRODUCT[832]) );
  FADDER S2_832_1 ( .CIN(\ab[832][1] ), .IN0(\CARRYB[831][1] ), .IN1(
        \SUMB[831][2] ), .COUT(\CARRYB[832][1] ), .SUM(\SUMB[832][1] ) );
  FADDER S3_832_2 ( .CIN(\ab[832][2] ), .IN0(\CARRYB[831][2] ), .IN1(
        \ab[831][3] ), .COUT(\CARRYB[832][2] ), .SUM(\SUMB[832][2] ) );
  FADDER S1_831_0 ( .CIN(\ab[831][0] ), .IN0(\CARRYB[830][0] ), .IN1(
        \SUMB[830][1] ), .COUT(\CARRYB[831][0] ), .SUM(PRODUCT[831]) );
  FADDER S2_831_1 ( .CIN(\ab[831][1] ), .IN0(\CARRYB[830][1] ), .IN1(
        \SUMB[830][2] ), .COUT(\CARRYB[831][1] ), .SUM(\SUMB[831][1] ) );
  FADDER S3_831_2 ( .CIN(\ab[831][2] ), .IN0(\CARRYB[830][2] ), .IN1(
        \ab[830][3] ), .COUT(\CARRYB[831][2] ), .SUM(\SUMB[831][2] ) );
  FADDER S1_830_0 ( .CIN(\ab[830][0] ), .IN0(\CARRYB[829][0] ), .IN1(
        \SUMB[829][1] ), .COUT(\CARRYB[830][0] ), .SUM(PRODUCT[830]) );
  FADDER S2_830_1 ( .CIN(\ab[830][1] ), .IN0(\CARRYB[829][1] ), .IN1(
        \SUMB[829][2] ), .COUT(\CARRYB[830][1] ), .SUM(\SUMB[830][1] ) );
  FADDER S3_830_2 ( .CIN(\ab[830][2] ), .IN0(\CARRYB[829][2] ), .IN1(
        \ab[829][3] ), .COUT(\CARRYB[830][2] ), .SUM(\SUMB[830][2] ) );
  FADDER S1_829_0 ( .CIN(\ab[829][0] ), .IN0(\CARRYB[828][0] ), .IN1(
        \SUMB[828][1] ), .COUT(\CARRYB[829][0] ), .SUM(PRODUCT[829]) );
  FADDER S2_829_1 ( .CIN(\ab[829][1] ), .IN0(\CARRYB[828][1] ), .IN1(
        \SUMB[828][2] ), .COUT(\CARRYB[829][1] ), .SUM(\SUMB[829][1] ) );
  FADDER S3_829_2 ( .CIN(\ab[829][2] ), .IN0(\CARRYB[828][2] ), .IN1(
        \ab[828][3] ), .COUT(\CARRYB[829][2] ), .SUM(\SUMB[829][2] ) );
  FADDER S1_828_0 ( .CIN(\ab[828][0] ), .IN0(\CARRYB[827][0] ), .IN1(
        \SUMB[827][1] ), .COUT(\CARRYB[828][0] ), .SUM(PRODUCT[828]) );
  FADDER S2_828_1 ( .CIN(\ab[828][1] ), .IN0(\CARRYB[827][1] ), .IN1(
        \SUMB[827][2] ), .COUT(\CARRYB[828][1] ), .SUM(\SUMB[828][1] ) );
  FADDER S3_828_2 ( .CIN(\ab[828][2] ), .IN0(\CARRYB[827][2] ), .IN1(
        \ab[827][3] ), .COUT(\CARRYB[828][2] ), .SUM(\SUMB[828][2] ) );
  FADDER S1_827_0 ( .CIN(\ab[827][0] ), .IN0(\CARRYB[826][0] ), .IN1(
        \SUMB[826][1] ), .COUT(\CARRYB[827][0] ), .SUM(PRODUCT[827]) );
  FADDER S2_827_1 ( .CIN(\ab[827][1] ), .IN0(\CARRYB[826][1] ), .IN1(
        \SUMB[826][2] ), .COUT(\CARRYB[827][1] ), .SUM(\SUMB[827][1] ) );
  FADDER S3_827_2 ( .CIN(\ab[827][2] ), .IN0(\CARRYB[826][2] ), .IN1(
        \ab[826][3] ), .COUT(\CARRYB[827][2] ), .SUM(\SUMB[827][2] ) );
  FADDER S1_826_0 ( .CIN(\ab[826][0] ), .IN0(\CARRYB[825][0] ), .IN1(
        \SUMB[825][1] ), .COUT(\CARRYB[826][0] ), .SUM(PRODUCT[826]) );
  FADDER S2_826_1 ( .CIN(\ab[826][1] ), .IN0(\CARRYB[825][1] ), .IN1(
        \SUMB[825][2] ), .COUT(\CARRYB[826][1] ), .SUM(\SUMB[826][1] ) );
  FADDER S3_826_2 ( .CIN(\ab[826][2] ), .IN0(\CARRYB[825][2] ), .IN1(
        \ab[825][3] ), .COUT(\CARRYB[826][2] ), .SUM(\SUMB[826][2] ) );
  FADDER S1_825_0 ( .CIN(\ab[825][0] ), .IN0(\CARRYB[824][0] ), .IN1(
        \SUMB[824][1] ), .COUT(\CARRYB[825][0] ), .SUM(PRODUCT[825]) );
  FADDER S2_825_1 ( .CIN(\ab[825][1] ), .IN0(\CARRYB[824][1] ), .IN1(
        \SUMB[824][2] ), .COUT(\CARRYB[825][1] ), .SUM(\SUMB[825][1] ) );
  FADDER S3_825_2 ( .CIN(\ab[825][2] ), .IN0(\CARRYB[824][2] ), .IN1(
        \ab[824][3] ), .COUT(\CARRYB[825][2] ), .SUM(\SUMB[825][2] ) );
  FADDER S1_824_0 ( .CIN(\ab[824][0] ), .IN0(\CARRYB[823][0] ), .IN1(
        \SUMB[823][1] ), .COUT(\CARRYB[824][0] ), .SUM(PRODUCT[824]) );
  FADDER S2_824_1 ( .CIN(\ab[824][1] ), .IN0(\CARRYB[823][1] ), .IN1(
        \SUMB[823][2] ), .COUT(\CARRYB[824][1] ), .SUM(\SUMB[824][1] ) );
  FADDER S3_824_2 ( .CIN(\ab[824][2] ), .IN0(\CARRYB[823][2] ), .IN1(
        \ab[823][3] ), .COUT(\CARRYB[824][2] ), .SUM(\SUMB[824][2] ) );
  FADDER S1_823_0 ( .CIN(\ab[823][0] ), .IN0(\CARRYB[822][0] ), .IN1(
        \SUMB[822][1] ), .COUT(\CARRYB[823][0] ), .SUM(PRODUCT[823]) );
  FADDER S2_823_1 ( .CIN(\ab[823][1] ), .IN0(\CARRYB[822][1] ), .IN1(
        \SUMB[822][2] ), .COUT(\CARRYB[823][1] ), .SUM(\SUMB[823][1] ) );
  FADDER S3_823_2 ( .CIN(\ab[823][2] ), .IN0(\CARRYB[822][2] ), .IN1(
        \ab[822][3] ), .COUT(\CARRYB[823][2] ), .SUM(\SUMB[823][2] ) );
  FADDER S1_822_0 ( .CIN(\ab[822][0] ), .IN0(\CARRYB[821][0] ), .IN1(
        \SUMB[821][1] ), .COUT(\CARRYB[822][0] ), .SUM(PRODUCT[822]) );
  FADDER S2_822_1 ( .CIN(\ab[822][1] ), .IN0(\CARRYB[821][1] ), .IN1(
        \SUMB[821][2] ), .COUT(\CARRYB[822][1] ), .SUM(\SUMB[822][1] ) );
  FADDER S3_822_2 ( .CIN(\ab[822][2] ), .IN0(\CARRYB[821][2] ), .IN1(
        \ab[821][3] ), .COUT(\CARRYB[822][2] ), .SUM(\SUMB[822][2] ) );
  FADDER S1_821_0 ( .CIN(\ab[821][0] ), .IN0(\CARRYB[820][0] ), .IN1(
        \SUMB[820][1] ), .COUT(\CARRYB[821][0] ), .SUM(PRODUCT[821]) );
  FADDER S2_821_1 ( .CIN(\ab[821][1] ), .IN0(\CARRYB[820][1] ), .IN1(
        \SUMB[820][2] ), .COUT(\CARRYB[821][1] ), .SUM(\SUMB[821][1] ) );
  FADDER S3_821_2 ( .CIN(\ab[821][2] ), .IN0(\CARRYB[820][2] ), .IN1(
        \ab[820][3] ), .COUT(\CARRYB[821][2] ), .SUM(\SUMB[821][2] ) );
  FADDER S1_820_0 ( .CIN(\ab[820][0] ), .IN0(\CARRYB[819][0] ), .IN1(
        \SUMB[819][1] ), .COUT(\CARRYB[820][0] ), .SUM(PRODUCT[820]) );
  FADDER S2_820_1 ( .CIN(\ab[820][1] ), .IN0(\CARRYB[819][1] ), .IN1(
        \SUMB[819][2] ), .COUT(\CARRYB[820][1] ), .SUM(\SUMB[820][1] ) );
  FADDER S3_820_2 ( .CIN(\ab[820][2] ), .IN0(\CARRYB[819][2] ), .IN1(
        \ab[819][3] ), .COUT(\CARRYB[820][2] ), .SUM(\SUMB[820][2] ) );
  FADDER S1_819_0 ( .CIN(\ab[819][0] ), .IN0(\CARRYB[818][0] ), .IN1(
        \SUMB[818][1] ), .COUT(\CARRYB[819][0] ), .SUM(PRODUCT[819]) );
  FADDER S2_819_1 ( .CIN(\ab[819][1] ), .IN0(\CARRYB[818][1] ), .IN1(
        \SUMB[818][2] ), .COUT(\CARRYB[819][1] ), .SUM(\SUMB[819][1] ) );
  FADDER S3_819_2 ( .CIN(\ab[819][2] ), .IN0(\CARRYB[818][2] ), .IN1(
        \ab[818][3] ), .COUT(\CARRYB[819][2] ), .SUM(\SUMB[819][2] ) );
  FADDER S1_818_0 ( .CIN(\ab[818][0] ), .IN0(\CARRYB[817][0] ), .IN1(
        \SUMB[817][1] ), .COUT(\CARRYB[818][0] ), .SUM(PRODUCT[818]) );
  FADDER S2_818_1 ( .CIN(\ab[818][1] ), .IN0(\CARRYB[817][1] ), .IN1(
        \SUMB[817][2] ), .COUT(\CARRYB[818][1] ), .SUM(\SUMB[818][1] ) );
  FADDER S3_818_2 ( .CIN(\ab[818][2] ), .IN0(\CARRYB[817][2] ), .IN1(
        \ab[817][3] ), .COUT(\CARRYB[818][2] ), .SUM(\SUMB[818][2] ) );
  FADDER S1_817_0 ( .CIN(\ab[817][0] ), .IN0(\CARRYB[816][0] ), .IN1(
        \SUMB[816][1] ), .COUT(\CARRYB[817][0] ), .SUM(PRODUCT[817]) );
  FADDER S2_817_1 ( .CIN(\ab[817][1] ), .IN0(\CARRYB[816][1] ), .IN1(
        \SUMB[816][2] ), .COUT(\CARRYB[817][1] ), .SUM(\SUMB[817][1] ) );
  FADDER S3_817_2 ( .CIN(\ab[817][2] ), .IN0(\CARRYB[816][2] ), .IN1(
        \ab[816][3] ), .COUT(\CARRYB[817][2] ), .SUM(\SUMB[817][2] ) );
  FADDER S1_816_0 ( .CIN(\ab[816][0] ), .IN0(\CARRYB[815][0] ), .IN1(
        \SUMB[815][1] ), .COUT(\CARRYB[816][0] ), .SUM(PRODUCT[816]) );
  FADDER S2_816_1 ( .CIN(\ab[816][1] ), .IN0(\CARRYB[815][1] ), .IN1(
        \SUMB[815][2] ), .COUT(\CARRYB[816][1] ), .SUM(\SUMB[816][1] ) );
  FADDER S3_816_2 ( .CIN(\ab[816][2] ), .IN0(\CARRYB[815][2] ), .IN1(
        \ab[815][3] ), .COUT(\CARRYB[816][2] ), .SUM(\SUMB[816][2] ) );
  FADDER S1_815_0 ( .CIN(\ab[815][0] ), .IN0(\CARRYB[814][0] ), .IN1(
        \SUMB[814][1] ), .COUT(\CARRYB[815][0] ), .SUM(PRODUCT[815]) );
  FADDER S2_815_1 ( .CIN(\ab[815][1] ), .IN0(\CARRYB[814][1] ), .IN1(
        \SUMB[814][2] ), .COUT(\CARRYB[815][1] ), .SUM(\SUMB[815][1] ) );
  FADDER S3_815_2 ( .CIN(\ab[815][2] ), .IN0(\CARRYB[814][2] ), .IN1(
        \ab[814][3] ), .COUT(\CARRYB[815][2] ), .SUM(\SUMB[815][2] ) );
  FADDER S1_814_0 ( .CIN(\ab[814][0] ), .IN0(\CARRYB[813][0] ), .IN1(
        \SUMB[813][1] ), .COUT(\CARRYB[814][0] ), .SUM(PRODUCT[814]) );
  FADDER S2_814_1 ( .CIN(\ab[814][1] ), .IN0(\CARRYB[813][1] ), .IN1(
        \SUMB[813][2] ), .COUT(\CARRYB[814][1] ), .SUM(\SUMB[814][1] ) );
  FADDER S3_814_2 ( .CIN(\ab[814][2] ), .IN0(\CARRYB[813][2] ), .IN1(
        \ab[813][3] ), .COUT(\CARRYB[814][2] ), .SUM(\SUMB[814][2] ) );
  FADDER S1_813_0 ( .CIN(\ab[813][0] ), .IN0(\CARRYB[812][0] ), .IN1(
        \SUMB[812][1] ), .COUT(\CARRYB[813][0] ), .SUM(PRODUCT[813]) );
  FADDER S2_813_1 ( .CIN(\ab[813][1] ), .IN0(\CARRYB[812][1] ), .IN1(
        \SUMB[812][2] ), .COUT(\CARRYB[813][1] ), .SUM(\SUMB[813][1] ) );
  FADDER S3_813_2 ( .CIN(\ab[813][2] ), .IN0(\CARRYB[812][2] ), .IN1(
        \ab[812][3] ), .COUT(\CARRYB[813][2] ), .SUM(\SUMB[813][2] ) );
  FADDER S1_812_0 ( .CIN(\ab[812][0] ), .IN0(\CARRYB[811][0] ), .IN1(
        \SUMB[811][1] ), .COUT(\CARRYB[812][0] ), .SUM(PRODUCT[812]) );
  FADDER S2_812_1 ( .CIN(\ab[812][1] ), .IN0(\CARRYB[811][1] ), .IN1(
        \SUMB[811][2] ), .COUT(\CARRYB[812][1] ), .SUM(\SUMB[812][1] ) );
  FADDER S3_812_2 ( .CIN(\ab[812][2] ), .IN0(\CARRYB[811][2] ), .IN1(
        \ab[811][3] ), .COUT(\CARRYB[812][2] ), .SUM(\SUMB[812][2] ) );
  FADDER S1_811_0 ( .CIN(\ab[811][0] ), .IN0(\CARRYB[810][0] ), .IN1(
        \SUMB[810][1] ), .COUT(\CARRYB[811][0] ), .SUM(PRODUCT[811]) );
  FADDER S2_811_1 ( .CIN(\ab[811][1] ), .IN0(\CARRYB[810][1] ), .IN1(
        \SUMB[810][2] ), .COUT(\CARRYB[811][1] ), .SUM(\SUMB[811][1] ) );
  FADDER S3_811_2 ( .CIN(\ab[811][2] ), .IN0(\CARRYB[810][2] ), .IN1(
        \ab[810][3] ), .COUT(\CARRYB[811][2] ), .SUM(\SUMB[811][2] ) );
  FADDER S1_810_0 ( .CIN(\ab[810][0] ), .IN0(\CARRYB[809][0] ), .IN1(
        \SUMB[809][1] ), .COUT(\CARRYB[810][0] ), .SUM(PRODUCT[810]) );
  FADDER S2_810_1 ( .CIN(\ab[810][1] ), .IN0(\CARRYB[809][1] ), .IN1(
        \SUMB[809][2] ), .COUT(\CARRYB[810][1] ), .SUM(\SUMB[810][1] ) );
  FADDER S3_810_2 ( .CIN(\ab[810][2] ), .IN0(\CARRYB[809][2] ), .IN1(
        \ab[809][3] ), .COUT(\CARRYB[810][2] ), .SUM(\SUMB[810][2] ) );
  FADDER S1_809_0 ( .CIN(\ab[809][0] ), .IN0(\CARRYB[808][0] ), .IN1(
        \SUMB[808][1] ), .COUT(\CARRYB[809][0] ), .SUM(PRODUCT[809]) );
  FADDER S2_809_1 ( .CIN(\ab[809][1] ), .IN0(\CARRYB[808][1] ), .IN1(
        \SUMB[808][2] ), .COUT(\CARRYB[809][1] ), .SUM(\SUMB[809][1] ) );
  FADDER S3_809_2 ( .CIN(\ab[809][2] ), .IN0(\CARRYB[808][2] ), .IN1(
        \ab[808][3] ), .COUT(\CARRYB[809][2] ), .SUM(\SUMB[809][2] ) );
  FADDER S1_808_0 ( .CIN(\ab[808][0] ), .IN0(\CARRYB[807][0] ), .IN1(
        \SUMB[807][1] ), .COUT(\CARRYB[808][0] ), .SUM(PRODUCT[808]) );
  FADDER S2_808_1 ( .CIN(\ab[808][1] ), .IN0(\CARRYB[807][1] ), .IN1(
        \SUMB[807][2] ), .COUT(\CARRYB[808][1] ), .SUM(\SUMB[808][1] ) );
  FADDER S3_808_2 ( .CIN(\ab[808][2] ), .IN0(\CARRYB[807][2] ), .IN1(
        \ab[807][3] ), .COUT(\CARRYB[808][2] ), .SUM(\SUMB[808][2] ) );
  FADDER S1_807_0 ( .CIN(\ab[807][0] ), .IN0(\CARRYB[806][0] ), .IN1(
        \SUMB[806][1] ), .COUT(\CARRYB[807][0] ), .SUM(PRODUCT[807]) );
  FADDER S2_807_1 ( .CIN(\ab[807][1] ), .IN0(\CARRYB[806][1] ), .IN1(
        \SUMB[806][2] ), .COUT(\CARRYB[807][1] ), .SUM(\SUMB[807][1] ) );
  FADDER S3_807_2 ( .CIN(\ab[807][2] ), .IN0(\CARRYB[806][2] ), .IN1(
        \ab[806][3] ), .COUT(\CARRYB[807][2] ), .SUM(\SUMB[807][2] ) );
  FADDER S1_806_0 ( .CIN(\ab[806][0] ), .IN0(\CARRYB[805][0] ), .IN1(
        \SUMB[805][1] ), .COUT(\CARRYB[806][0] ), .SUM(PRODUCT[806]) );
  FADDER S2_806_1 ( .CIN(\ab[806][1] ), .IN0(\CARRYB[805][1] ), .IN1(
        \SUMB[805][2] ), .COUT(\CARRYB[806][1] ), .SUM(\SUMB[806][1] ) );
  FADDER S3_806_2 ( .CIN(\ab[806][2] ), .IN0(\CARRYB[805][2] ), .IN1(
        \ab[805][3] ), .COUT(\CARRYB[806][2] ), .SUM(\SUMB[806][2] ) );
  FADDER S1_805_0 ( .CIN(\ab[805][0] ), .IN0(\CARRYB[804][0] ), .IN1(
        \SUMB[804][1] ), .COUT(\CARRYB[805][0] ), .SUM(PRODUCT[805]) );
  FADDER S2_805_1 ( .CIN(\ab[805][1] ), .IN0(\CARRYB[804][1] ), .IN1(
        \SUMB[804][2] ), .COUT(\CARRYB[805][1] ), .SUM(\SUMB[805][1] ) );
  FADDER S3_805_2 ( .CIN(\ab[805][2] ), .IN0(\CARRYB[804][2] ), .IN1(
        \ab[804][3] ), .COUT(\CARRYB[805][2] ), .SUM(\SUMB[805][2] ) );
  FADDER S1_804_0 ( .CIN(\ab[804][0] ), .IN0(\CARRYB[803][0] ), .IN1(
        \SUMB[803][1] ), .COUT(\CARRYB[804][0] ), .SUM(PRODUCT[804]) );
  FADDER S2_804_1 ( .CIN(\ab[804][1] ), .IN0(\CARRYB[803][1] ), .IN1(
        \SUMB[803][2] ), .COUT(\CARRYB[804][1] ), .SUM(\SUMB[804][1] ) );
  FADDER S3_804_2 ( .CIN(\ab[804][2] ), .IN0(\CARRYB[803][2] ), .IN1(
        \ab[803][3] ), .COUT(\CARRYB[804][2] ), .SUM(\SUMB[804][2] ) );
  FADDER S1_803_0 ( .CIN(\ab[803][0] ), .IN0(\CARRYB[802][0] ), .IN1(
        \SUMB[802][1] ), .COUT(\CARRYB[803][0] ), .SUM(PRODUCT[803]) );
  FADDER S2_803_1 ( .CIN(\ab[803][1] ), .IN0(\CARRYB[802][1] ), .IN1(
        \SUMB[802][2] ), .COUT(\CARRYB[803][1] ), .SUM(\SUMB[803][1] ) );
  FADDER S3_803_2 ( .CIN(\ab[803][2] ), .IN0(\CARRYB[802][2] ), .IN1(
        \ab[802][3] ), .COUT(\CARRYB[803][2] ), .SUM(\SUMB[803][2] ) );
  FADDER S1_802_0 ( .CIN(\ab[802][0] ), .IN0(\CARRYB[801][0] ), .IN1(
        \SUMB[801][1] ), .COUT(\CARRYB[802][0] ), .SUM(PRODUCT[802]) );
  FADDER S2_802_1 ( .CIN(\ab[802][1] ), .IN0(\CARRYB[801][1] ), .IN1(
        \SUMB[801][2] ), .COUT(\CARRYB[802][1] ), .SUM(\SUMB[802][1] ) );
  FADDER S3_802_2 ( .CIN(\ab[802][2] ), .IN0(\CARRYB[801][2] ), .IN1(
        \ab[801][3] ), .COUT(\CARRYB[802][2] ), .SUM(\SUMB[802][2] ) );
  FADDER S1_801_0 ( .CIN(\ab[801][0] ), .IN0(\CARRYB[800][0] ), .IN1(
        \SUMB[800][1] ), .COUT(\CARRYB[801][0] ), .SUM(PRODUCT[801]) );
  FADDER S2_801_1 ( .CIN(\ab[801][1] ), .IN0(\CARRYB[800][1] ), .IN1(
        \SUMB[800][2] ), .COUT(\CARRYB[801][1] ), .SUM(\SUMB[801][1] ) );
  FADDER S3_801_2 ( .CIN(\ab[801][2] ), .IN0(\CARRYB[800][2] ), .IN1(
        \ab[800][3] ), .COUT(\CARRYB[801][2] ), .SUM(\SUMB[801][2] ) );
  FADDER S1_800_0 ( .CIN(\ab[800][0] ), .IN0(\CARRYB[799][0] ), .IN1(
        \SUMB[799][1] ), .COUT(\CARRYB[800][0] ), .SUM(PRODUCT[800]) );
  FADDER S2_800_1 ( .CIN(\ab[800][1] ), .IN0(\CARRYB[799][1] ), .IN1(
        \SUMB[799][2] ), .COUT(\CARRYB[800][1] ), .SUM(\SUMB[800][1] ) );
  FADDER S3_800_2 ( .CIN(\ab[800][2] ), .IN0(\CARRYB[799][2] ), .IN1(
        \ab[799][3] ), .COUT(\CARRYB[800][2] ), .SUM(\SUMB[800][2] ) );
  FADDER S1_799_0 ( .CIN(\ab[799][0] ), .IN0(\CARRYB[798][0] ), .IN1(
        \SUMB[798][1] ), .COUT(\CARRYB[799][0] ), .SUM(PRODUCT[799]) );
  FADDER S2_799_1 ( .CIN(\ab[799][1] ), .IN0(\CARRYB[798][1] ), .IN1(
        \SUMB[798][2] ), .COUT(\CARRYB[799][1] ), .SUM(\SUMB[799][1] ) );
  FADDER S3_799_2 ( .CIN(\ab[799][2] ), .IN0(\CARRYB[798][2] ), .IN1(
        \ab[798][3] ), .COUT(\CARRYB[799][2] ), .SUM(\SUMB[799][2] ) );
  FADDER S1_798_0 ( .CIN(\ab[798][0] ), .IN0(\CARRYB[797][0] ), .IN1(
        \SUMB[797][1] ), .COUT(\CARRYB[798][0] ), .SUM(PRODUCT[798]) );
  FADDER S2_798_1 ( .CIN(\ab[798][1] ), .IN0(\CARRYB[797][1] ), .IN1(
        \SUMB[797][2] ), .COUT(\CARRYB[798][1] ), .SUM(\SUMB[798][1] ) );
  FADDER S3_798_2 ( .CIN(\ab[798][2] ), .IN0(\CARRYB[797][2] ), .IN1(
        \ab[797][3] ), .COUT(\CARRYB[798][2] ), .SUM(\SUMB[798][2] ) );
  FADDER S1_797_0 ( .CIN(\ab[797][0] ), .IN0(\CARRYB[796][0] ), .IN1(
        \SUMB[796][1] ), .COUT(\CARRYB[797][0] ), .SUM(PRODUCT[797]) );
  FADDER S2_797_1 ( .CIN(\ab[797][1] ), .IN0(\CARRYB[796][1] ), .IN1(
        \SUMB[796][2] ), .COUT(\CARRYB[797][1] ), .SUM(\SUMB[797][1] ) );
  FADDER S3_797_2 ( .CIN(\ab[797][2] ), .IN0(\CARRYB[796][2] ), .IN1(
        \ab[796][3] ), .COUT(\CARRYB[797][2] ), .SUM(\SUMB[797][2] ) );
  FADDER S1_796_0 ( .CIN(\ab[796][0] ), .IN0(\CARRYB[795][0] ), .IN1(
        \SUMB[795][1] ), .COUT(\CARRYB[796][0] ), .SUM(PRODUCT[796]) );
  FADDER S2_796_1 ( .CIN(\ab[796][1] ), .IN0(\CARRYB[795][1] ), .IN1(
        \SUMB[795][2] ), .COUT(\CARRYB[796][1] ), .SUM(\SUMB[796][1] ) );
  FADDER S3_796_2 ( .CIN(\ab[796][2] ), .IN0(\CARRYB[795][2] ), .IN1(
        \ab[795][3] ), .COUT(\CARRYB[796][2] ), .SUM(\SUMB[796][2] ) );
  FADDER S1_795_0 ( .CIN(\ab[795][0] ), .IN0(\CARRYB[794][0] ), .IN1(
        \SUMB[794][1] ), .COUT(\CARRYB[795][0] ), .SUM(PRODUCT[795]) );
  FADDER S2_795_1 ( .CIN(\ab[795][1] ), .IN0(\CARRYB[794][1] ), .IN1(
        \SUMB[794][2] ), .COUT(\CARRYB[795][1] ), .SUM(\SUMB[795][1] ) );
  FADDER S3_795_2 ( .CIN(\ab[795][2] ), .IN0(\CARRYB[794][2] ), .IN1(
        \ab[794][3] ), .COUT(\CARRYB[795][2] ), .SUM(\SUMB[795][2] ) );
  FADDER S1_794_0 ( .CIN(\ab[794][0] ), .IN0(\CARRYB[793][0] ), .IN1(
        \SUMB[793][1] ), .COUT(\CARRYB[794][0] ), .SUM(PRODUCT[794]) );
  FADDER S2_794_1 ( .CIN(\ab[794][1] ), .IN0(\CARRYB[793][1] ), .IN1(
        \SUMB[793][2] ), .COUT(\CARRYB[794][1] ), .SUM(\SUMB[794][1] ) );
  FADDER S3_794_2 ( .CIN(\ab[794][2] ), .IN0(\CARRYB[793][2] ), .IN1(
        \ab[793][3] ), .COUT(\CARRYB[794][2] ), .SUM(\SUMB[794][2] ) );
  FADDER S1_793_0 ( .CIN(\ab[793][0] ), .IN0(\CARRYB[792][0] ), .IN1(
        \SUMB[792][1] ), .COUT(\CARRYB[793][0] ), .SUM(PRODUCT[793]) );
  FADDER S2_793_1 ( .CIN(\ab[793][1] ), .IN0(\CARRYB[792][1] ), .IN1(
        \SUMB[792][2] ), .COUT(\CARRYB[793][1] ), .SUM(\SUMB[793][1] ) );
  FADDER S3_793_2 ( .CIN(\ab[793][2] ), .IN0(\CARRYB[792][2] ), .IN1(
        \ab[792][3] ), .COUT(\CARRYB[793][2] ), .SUM(\SUMB[793][2] ) );
  FADDER S1_792_0 ( .CIN(\ab[792][0] ), .IN0(\CARRYB[791][0] ), .IN1(
        \SUMB[791][1] ), .COUT(\CARRYB[792][0] ), .SUM(PRODUCT[792]) );
  FADDER S2_792_1 ( .CIN(\ab[792][1] ), .IN0(\CARRYB[791][1] ), .IN1(
        \SUMB[791][2] ), .COUT(\CARRYB[792][1] ), .SUM(\SUMB[792][1] ) );
  FADDER S3_792_2 ( .CIN(\ab[792][2] ), .IN0(\CARRYB[791][2] ), .IN1(
        \ab[791][3] ), .COUT(\CARRYB[792][2] ), .SUM(\SUMB[792][2] ) );
  FADDER S1_791_0 ( .CIN(\ab[791][0] ), .IN0(\CARRYB[790][0] ), .IN1(
        \SUMB[790][1] ), .COUT(\CARRYB[791][0] ), .SUM(PRODUCT[791]) );
  FADDER S2_791_1 ( .CIN(\ab[791][1] ), .IN0(\CARRYB[790][1] ), .IN1(
        \SUMB[790][2] ), .COUT(\CARRYB[791][1] ), .SUM(\SUMB[791][1] ) );
  FADDER S3_791_2 ( .CIN(\ab[791][2] ), .IN0(\CARRYB[790][2] ), .IN1(
        \ab[790][3] ), .COUT(\CARRYB[791][2] ), .SUM(\SUMB[791][2] ) );
  FADDER S1_790_0 ( .CIN(\ab[790][0] ), .IN0(\CARRYB[789][0] ), .IN1(
        \SUMB[789][1] ), .COUT(\CARRYB[790][0] ), .SUM(PRODUCT[790]) );
  FADDER S2_790_1 ( .CIN(\ab[790][1] ), .IN0(\CARRYB[789][1] ), .IN1(
        \SUMB[789][2] ), .COUT(\CARRYB[790][1] ), .SUM(\SUMB[790][1] ) );
  FADDER S3_790_2 ( .CIN(\ab[790][2] ), .IN0(\CARRYB[789][2] ), .IN1(
        \ab[789][3] ), .COUT(\CARRYB[790][2] ), .SUM(\SUMB[790][2] ) );
  FADDER S1_789_0 ( .CIN(\ab[789][0] ), .IN0(\CARRYB[788][0] ), .IN1(
        \SUMB[788][1] ), .COUT(\CARRYB[789][0] ), .SUM(PRODUCT[789]) );
  FADDER S2_789_1 ( .CIN(\ab[789][1] ), .IN0(\CARRYB[788][1] ), .IN1(
        \SUMB[788][2] ), .COUT(\CARRYB[789][1] ), .SUM(\SUMB[789][1] ) );
  FADDER S3_789_2 ( .CIN(\ab[789][2] ), .IN0(\CARRYB[788][2] ), .IN1(
        \ab[788][3] ), .COUT(\CARRYB[789][2] ), .SUM(\SUMB[789][2] ) );
  FADDER S1_788_0 ( .CIN(\ab[788][0] ), .IN0(\CARRYB[787][0] ), .IN1(
        \SUMB[787][1] ), .COUT(\CARRYB[788][0] ), .SUM(PRODUCT[788]) );
  FADDER S2_788_1 ( .CIN(\ab[788][1] ), .IN0(\CARRYB[787][1] ), .IN1(
        \SUMB[787][2] ), .COUT(\CARRYB[788][1] ), .SUM(\SUMB[788][1] ) );
  FADDER S3_788_2 ( .CIN(\ab[788][2] ), .IN0(\CARRYB[787][2] ), .IN1(
        \ab[787][3] ), .COUT(\CARRYB[788][2] ), .SUM(\SUMB[788][2] ) );
  FADDER S1_787_0 ( .CIN(\ab[787][0] ), .IN0(\CARRYB[786][0] ), .IN1(
        \SUMB[786][1] ), .COUT(\CARRYB[787][0] ), .SUM(PRODUCT[787]) );
  FADDER S2_787_1 ( .CIN(\ab[787][1] ), .IN0(\CARRYB[786][1] ), .IN1(
        \SUMB[786][2] ), .COUT(\CARRYB[787][1] ), .SUM(\SUMB[787][1] ) );
  FADDER S3_787_2 ( .CIN(\ab[787][2] ), .IN0(\CARRYB[786][2] ), .IN1(
        \ab[786][3] ), .COUT(\CARRYB[787][2] ), .SUM(\SUMB[787][2] ) );
  FADDER S1_786_0 ( .CIN(\ab[786][0] ), .IN0(\CARRYB[785][0] ), .IN1(
        \SUMB[785][1] ), .COUT(\CARRYB[786][0] ), .SUM(PRODUCT[786]) );
  FADDER S2_786_1 ( .CIN(\ab[786][1] ), .IN0(\CARRYB[785][1] ), .IN1(
        \SUMB[785][2] ), .COUT(\CARRYB[786][1] ), .SUM(\SUMB[786][1] ) );
  FADDER S3_786_2 ( .CIN(\ab[786][2] ), .IN0(\CARRYB[785][2] ), .IN1(
        \ab[785][3] ), .COUT(\CARRYB[786][2] ), .SUM(\SUMB[786][2] ) );
  FADDER S1_785_0 ( .CIN(\ab[785][0] ), .IN0(\CARRYB[784][0] ), .IN1(
        \SUMB[784][1] ), .COUT(\CARRYB[785][0] ), .SUM(PRODUCT[785]) );
  FADDER S2_785_1 ( .CIN(\ab[785][1] ), .IN0(\CARRYB[784][1] ), .IN1(
        \SUMB[784][2] ), .COUT(\CARRYB[785][1] ), .SUM(\SUMB[785][1] ) );
  FADDER S3_785_2 ( .CIN(\ab[785][2] ), .IN0(\CARRYB[784][2] ), .IN1(
        \ab[784][3] ), .COUT(\CARRYB[785][2] ), .SUM(\SUMB[785][2] ) );
  FADDER S1_784_0 ( .CIN(\ab[784][0] ), .IN0(\CARRYB[783][0] ), .IN1(
        \SUMB[783][1] ), .COUT(\CARRYB[784][0] ), .SUM(PRODUCT[784]) );
  FADDER S2_784_1 ( .CIN(\ab[784][1] ), .IN0(\CARRYB[783][1] ), .IN1(
        \SUMB[783][2] ), .COUT(\CARRYB[784][1] ), .SUM(\SUMB[784][1] ) );
  FADDER S3_784_2 ( .CIN(\ab[784][2] ), .IN0(\CARRYB[783][2] ), .IN1(
        \ab[783][3] ), .COUT(\CARRYB[784][2] ), .SUM(\SUMB[784][2] ) );
  FADDER S1_783_0 ( .CIN(\ab[783][0] ), .IN0(\CARRYB[782][0] ), .IN1(
        \SUMB[782][1] ), .COUT(\CARRYB[783][0] ), .SUM(PRODUCT[783]) );
  FADDER S2_783_1 ( .CIN(\ab[783][1] ), .IN0(\CARRYB[782][1] ), .IN1(
        \SUMB[782][2] ), .COUT(\CARRYB[783][1] ), .SUM(\SUMB[783][1] ) );
  FADDER S3_783_2 ( .CIN(\ab[783][2] ), .IN0(\CARRYB[782][2] ), .IN1(
        \ab[782][3] ), .COUT(\CARRYB[783][2] ), .SUM(\SUMB[783][2] ) );
  FADDER S1_782_0 ( .CIN(\ab[782][0] ), .IN0(\CARRYB[781][0] ), .IN1(
        \SUMB[781][1] ), .COUT(\CARRYB[782][0] ), .SUM(PRODUCT[782]) );
  FADDER S2_782_1 ( .CIN(\ab[782][1] ), .IN0(\CARRYB[781][1] ), .IN1(
        \SUMB[781][2] ), .COUT(\CARRYB[782][1] ), .SUM(\SUMB[782][1] ) );
  FADDER S3_782_2 ( .CIN(\ab[782][2] ), .IN0(\CARRYB[781][2] ), .IN1(
        \ab[781][3] ), .COUT(\CARRYB[782][2] ), .SUM(\SUMB[782][2] ) );
  FADDER S1_781_0 ( .CIN(\ab[781][0] ), .IN0(\CARRYB[780][0] ), .IN1(
        \SUMB[780][1] ), .COUT(\CARRYB[781][0] ), .SUM(PRODUCT[781]) );
  FADDER S2_781_1 ( .CIN(\ab[781][1] ), .IN0(\CARRYB[780][1] ), .IN1(
        \SUMB[780][2] ), .COUT(\CARRYB[781][1] ), .SUM(\SUMB[781][1] ) );
  FADDER S3_781_2 ( .CIN(\ab[781][2] ), .IN0(\CARRYB[780][2] ), .IN1(
        \ab[780][3] ), .COUT(\CARRYB[781][2] ), .SUM(\SUMB[781][2] ) );
  FADDER S1_780_0 ( .CIN(\ab[780][0] ), .IN0(\CARRYB[779][0] ), .IN1(
        \SUMB[779][1] ), .COUT(\CARRYB[780][0] ), .SUM(PRODUCT[780]) );
  FADDER S2_780_1 ( .CIN(\ab[780][1] ), .IN0(\CARRYB[779][1] ), .IN1(
        \SUMB[779][2] ), .COUT(\CARRYB[780][1] ), .SUM(\SUMB[780][1] ) );
  FADDER S3_780_2 ( .CIN(\ab[780][2] ), .IN0(\CARRYB[779][2] ), .IN1(
        \ab[779][3] ), .COUT(\CARRYB[780][2] ), .SUM(\SUMB[780][2] ) );
  FADDER S1_779_0 ( .CIN(\ab[779][0] ), .IN0(\CARRYB[778][0] ), .IN1(
        \SUMB[778][1] ), .COUT(\CARRYB[779][0] ), .SUM(PRODUCT[779]) );
  FADDER S2_779_1 ( .CIN(\ab[779][1] ), .IN0(\CARRYB[778][1] ), .IN1(
        \SUMB[778][2] ), .COUT(\CARRYB[779][1] ), .SUM(\SUMB[779][1] ) );
  FADDER S3_779_2 ( .CIN(\ab[779][2] ), .IN0(\CARRYB[778][2] ), .IN1(
        \ab[778][3] ), .COUT(\CARRYB[779][2] ), .SUM(\SUMB[779][2] ) );
  FADDER S1_778_0 ( .CIN(\ab[778][0] ), .IN0(\CARRYB[777][0] ), .IN1(
        \SUMB[777][1] ), .COUT(\CARRYB[778][0] ), .SUM(PRODUCT[778]) );
  FADDER S2_778_1 ( .CIN(\ab[778][1] ), .IN0(\CARRYB[777][1] ), .IN1(
        \SUMB[777][2] ), .COUT(\CARRYB[778][1] ), .SUM(\SUMB[778][1] ) );
  FADDER S3_778_2 ( .CIN(\ab[778][2] ), .IN0(\CARRYB[777][2] ), .IN1(
        \ab[777][3] ), .COUT(\CARRYB[778][2] ), .SUM(\SUMB[778][2] ) );
  FADDER S1_777_0 ( .CIN(\ab[777][0] ), .IN0(\CARRYB[776][0] ), .IN1(
        \SUMB[776][1] ), .COUT(\CARRYB[777][0] ), .SUM(PRODUCT[777]) );
  FADDER S2_777_1 ( .CIN(\ab[777][1] ), .IN0(\CARRYB[776][1] ), .IN1(
        \SUMB[776][2] ), .COUT(\CARRYB[777][1] ), .SUM(\SUMB[777][1] ) );
  FADDER S3_777_2 ( .CIN(\ab[777][2] ), .IN0(\CARRYB[776][2] ), .IN1(
        \ab[776][3] ), .COUT(\CARRYB[777][2] ), .SUM(\SUMB[777][2] ) );
  FADDER S1_776_0 ( .CIN(\ab[776][0] ), .IN0(\CARRYB[775][0] ), .IN1(
        \SUMB[775][1] ), .COUT(\CARRYB[776][0] ), .SUM(PRODUCT[776]) );
  FADDER S2_776_1 ( .CIN(\ab[776][1] ), .IN0(\CARRYB[775][1] ), .IN1(
        \SUMB[775][2] ), .COUT(\CARRYB[776][1] ), .SUM(\SUMB[776][1] ) );
  FADDER S3_776_2 ( .CIN(\ab[776][2] ), .IN0(\CARRYB[775][2] ), .IN1(
        \ab[775][3] ), .COUT(\CARRYB[776][2] ), .SUM(\SUMB[776][2] ) );
  FADDER S1_775_0 ( .CIN(\ab[775][0] ), .IN0(\CARRYB[774][0] ), .IN1(
        \SUMB[774][1] ), .COUT(\CARRYB[775][0] ), .SUM(PRODUCT[775]) );
  FADDER S2_775_1 ( .CIN(\ab[775][1] ), .IN0(\CARRYB[774][1] ), .IN1(
        \SUMB[774][2] ), .COUT(\CARRYB[775][1] ), .SUM(\SUMB[775][1] ) );
  FADDER S3_775_2 ( .CIN(\ab[775][2] ), .IN0(\CARRYB[774][2] ), .IN1(
        \ab[774][3] ), .COUT(\CARRYB[775][2] ), .SUM(\SUMB[775][2] ) );
  FADDER S1_774_0 ( .CIN(\ab[774][0] ), .IN0(\CARRYB[773][0] ), .IN1(
        \SUMB[773][1] ), .COUT(\CARRYB[774][0] ), .SUM(PRODUCT[774]) );
  FADDER S2_774_1 ( .CIN(\ab[774][1] ), .IN0(\CARRYB[773][1] ), .IN1(
        \SUMB[773][2] ), .COUT(\CARRYB[774][1] ), .SUM(\SUMB[774][1] ) );
  FADDER S3_774_2 ( .CIN(\ab[774][2] ), .IN0(\CARRYB[773][2] ), .IN1(
        \ab[773][3] ), .COUT(\CARRYB[774][2] ), .SUM(\SUMB[774][2] ) );
  FADDER S1_773_0 ( .CIN(\ab[773][0] ), .IN0(\CARRYB[772][0] ), .IN1(
        \SUMB[772][1] ), .COUT(\CARRYB[773][0] ), .SUM(PRODUCT[773]) );
  FADDER S2_773_1 ( .CIN(\ab[773][1] ), .IN0(\CARRYB[772][1] ), .IN1(
        \SUMB[772][2] ), .COUT(\CARRYB[773][1] ), .SUM(\SUMB[773][1] ) );
  FADDER S3_773_2 ( .CIN(\ab[773][2] ), .IN0(\CARRYB[772][2] ), .IN1(
        \ab[772][3] ), .COUT(\CARRYB[773][2] ), .SUM(\SUMB[773][2] ) );
  FADDER S1_772_0 ( .CIN(\ab[772][0] ), .IN0(\CARRYB[771][0] ), .IN1(
        \SUMB[771][1] ), .COUT(\CARRYB[772][0] ), .SUM(PRODUCT[772]) );
  FADDER S2_772_1 ( .CIN(\ab[772][1] ), .IN0(\CARRYB[771][1] ), .IN1(
        \SUMB[771][2] ), .COUT(\CARRYB[772][1] ), .SUM(\SUMB[772][1] ) );
  FADDER S3_772_2 ( .CIN(\ab[772][2] ), .IN0(\CARRYB[771][2] ), .IN1(
        \ab[771][3] ), .COUT(\CARRYB[772][2] ), .SUM(\SUMB[772][2] ) );
  FADDER S1_771_0 ( .CIN(\ab[771][0] ), .IN0(\CARRYB[770][0] ), .IN1(
        \SUMB[770][1] ), .COUT(\CARRYB[771][0] ), .SUM(PRODUCT[771]) );
  FADDER S2_771_1 ( .CIN(\ab[771][1] ), .IN0(\CARRYB[770][1] ), .IN1(
        \SUMB[770][2] ), .COUT(\CARRYB[771][1] ), .SUM(\SUMB[771][1] ) );
  FADDER S3_771_2 ( .CIN(\ab[771][2] ), .IN0(\CARRYB[770][2] ), .IN1(
        \ab[770][3] ), .COUT(\CARRYB[771][2] ), .SUM(\SUMB[771][2] ) );
  FADDER S1_770_0 ( .CIN(\ab[770][0] ), .IN0(\CARRYB[769][0] ), .IN1(
        \SUMB[769][1] ), .COUT(\CARRYB[770][0] ), .SUM(PRODUCT[770]) );
  FADDER S2_770_1 ( .CIN(\ab[770][1] ), .IN0(\CARRYB[769][1] ), .IN1(
        \SUMB[769][2] ), .COUT(\CARRYB[770][1] ), .SUM(\SUMB[770][1] ) );
  FADDER S3_770_2 ( .CIN(\ab[770][2] ), .IN0(\CARRYB[769][2] ), .IN1(
        \ab[769][3] ), .COUT(\CARRYB[770][2] ), .SUM(\SUMB[770][2] ) );
  FADDER S1_769_0 ( .CIN(\ab[769][0] ), .IN0(\CARRYB[768][0] ), .IN1(
        \SUMB[768][1] ), .COUT(\CARRYB[769][0] ), .SUM(PRODUCT[769]) );
  FADDER S2_769_1 ( .CIN(\ab[769][1] ), .IN0(\CARRYB[768][1] ), .IN1(
        \SUMB[768][2] ), .COUT(\CARRYB[769][1] ), .SUM(\SUMB[769][1] ) );
  FADDER S3_769_2 ( .CIN(\ab[769][2] ), .IN0(\CARRYB[768][2] ), .IN1(
        \ab[768][3] ), .COUT(\CARRYB[769][2] ), .SUM(\SUMB[769][2] ) );
  FADDER S1_768_0 ( .CIN(\ab[768][0] ), .IN0(\CARRYB[767][0] ), .IN1(
        \SUMB[767][1] ), .COUT(\CARRYB[768][0] ), .SUM(PRODUCT[768]) );
  FADDER S2_768_1 ( .CIN(\ab[768][1] ), .IN0(\CARRYB[767][1] ), .IN1(
        \SUMB[767][2] ), .COUT(\CARRYB[768][1] ), .SUM(\SUMB[768][1] ) );
  FADDER S3_768_2 ( .CIN(\ab[768][2] ), .IN0(\CARRYB[767][2] ), .IN1(
        \ab[767][3] ), .COUT(\CARRYB[768][2] ), .SUM(\SUMB[768][2] ) );
  FADDER S1_767_0 ( .CIN(\ab[767][0] ), .IN0(\CARRYB[766][0] ), .IN1(
        \SUMB[766][1] ), .COUT(\CARRYB[767][0] ), .SUM(PRODUCT[767]) );
  FADDER S2_767_1 ( .CIN(\ab[767][1] ), .IN0(\CARRYB[766][1] ), .IN1(
        \SUMB[766][2] ), .COUT(\CARRYB[767][1] ), .SUM(\SUMB[767][1] ) );
  FADDER S3_767_2 ( .CIN(\ab[767][2] ), .IN0(\CARRYB[766][2] ), .IN1(
        \ab[766][3] ), .COUT(\CARRYB[767][2] ), .SUM(\SUMB[767][2] ) );
  FADDER S1_766_0 ( .CIN(\ab[766][0] ), .IN0(\CARRYB[765][0] ), .IN1(
        \SUMB[765][1] ), .COUT(\CARRYB[766][0] ), .SUM(PRODUCT[766]) );
  FADDER S2_766_1 ( .CIN(\ab[766][1] ), .IN0(\CARRYB[765][1] ), .IN1(
        \SUMB[765][2] ), .COUT(\CARRYB[766][1] ), .SUM(\SUMB[766][1] ) );
  FADDER S3_766_2 ( .CIN(\ab[766][2] ), .IN0(\CARRYB[765][2] ), .IN1(
        \ab[765][3] ), .COUT(\CARRYB[766][2] ), .SUM(\SUMB[766][2] ) );
  FADDER S1_765_0 ( .CIN(\ab[765][0] ), .IN0(\CARRYB[764][0] ), .IN1(
        \SUMB[764][1] ), .COUT(\CARRYB[765][0] ), .SUM(PRODUCT[765]) );
  FADDER S2_765_1 ( .CIN(\ab[765][1] ), .IN0(\CARRYB[764][1] ), .IN1(
        \SUMB[764][2] ), .COUT(\CARRYB[765][1] ), .SUM(\SUMB[765][1] ) );
  FADDER S3_765_2 ( .CIN(\ab[765][2] ), .IN0(\CARRYB[764][2] ), .IN1(
        \ab[764][3] ), .COUT(\CARRYB[765][2] ), .SUM(\SUMB[765][2] ) );
  FADDER S1_764_0 ( .CIN(\ab[764][0] ), .IN0(\CARRYB[763][0] ), .IN1(
        \SUMB[763][1] ), .COUT(\CARRYB[764][0] ), .SUM(PRODUCT[764]) );
  FADDER S2_764_1 ( .CIN(\ab[764][1] ), .IN0(\CARRYB[763][1] ), .IN1(
        \SUMB[763][2] ), .COUT(\CARRYB[764][1] ), .SUM(\SUMB[764][1] ) );
  FADDER S3_764_2 ( .CIN(\ab[764][2] ), .IN0(\CARRYB[763][2] ), .IN1(
        \ab[763][3] ), .COUT(\CARRYB[764][2] ), .SUM(\SUMB[764][2] ) );
  FADDER S1_763_0 ( .CIN(\ab[763][0] ), .IN0(\CARRYB[762][0] ), .IN1(
        \SUMB[762][1] ), .COUT(\CARRYB[763][0] ), .SUM(PRODUCT[763]) );
  FADDER S2_763_1 ( .CIN(\ab[763][1] ), .IN0(\CARRYB[762][1] ), .IN1(
        \SUMB[762][2] ), .COUT(\CARRYB[763][1] ), .SUM(\SUMB[763][1] ) );
  FADDER S3_763_2 ( .CIN(\ab[763][2] ), .IN0(\CARRYB[762][2] ), .IN1(
        \ab[762][3] ), .COUT(\CARRYB[763][2] ), .SUM(\SUMB[763][2] ) );
  FADDER S1_762_0 ( .CIN(\ab[762][0] ), .IN0(\CARRYB[761][0] ), .IN1(
        \SUMB[761][1] ), .COUT(\CARRYB[762][0] ), .SUM(PRODUCT[762]) );
  FADDER S2_762_1 ( .CIN(\ab[762][1] ), .IN0(\CARRYB[761][1] ), .IN1(
        \SUMB[761][2] ), .COUT(\CARRYB[762][1] ), .SUM(\SUMB[762][1] ) );
  FADDER S3_762_2 ( .CIN(\ab[762][2] ), .IN0(\CARRYB[761][2] ), .IN1(
        \ab[761][3] ), .COUT(\CARRYB[762][2] ), .SUM(\SUMB[762][2] ) );
  FADDER S1_761_0 ( .CIN(\ab[761][0] ), .IN0(\CARRYB[760][0] ), .IN1(
        \SUMB[760][1] ), .COUT(\CARRYB[761][0] ), .SUM(PRODUCT[761]) );
  FADDER S2_761_1 ( .CIN(\ab[761][1] ), .IN0(\CARRYB[760][1] ), .IN1(
        \SUMB[760][2] ), .COUT(\CARRYB[761][1] ), .SUM(\SUMB[761][1] ) );
  FADDER S3_761_2 ( .CIN(\ab[761][2] ), .IN0(\CARRYB[760][2] ), .IN1(
        \ab[760][3] ), .COUT(\CARRYB[761][2] ), .SUM(\SUMB[761][2] ) );
  FADDER S1_760_0 ( .CIN(\ab[760][0] ), .IN0(\CARRYB[759][0] ), .IN1(
        \SUMB[759][1] ), .COUT(\CARRYB[760][0] ), .SUM(PRODUCT[760]) );
  FADDER S2_760_1 ( .CIN(\ab[760][1] ), .IN0(\CARRYB[759][1] ), .IN1(
        \SUMB[759][2] ), .COUT(\CARRYB[760][1] ), .SUM(\SUMB[760][1] ) );
  FADDER S3_760_2 ( .CIN(\ab[760][2] ), .IN0(\CARRYB[759][2] ), .IN1(
        \ab[759][3] ), .COUT(\CARRYB[760][2] ), .SUM(\SUMB[760][2] ) );
  FADDER S1_759_0 ( .CIN(\ab[759][0] ), .IN0(\CARRYB[758][0] ), .IN1(
        \SUMB[758][1] ), .COUT(\CARRYB[759][0] ), .SUM(PRODUCT[759]) );
  FADDER S2_759_1 ( .CIN(\ab[759][1] ), .IN0(\CARRYB[758][1] ), .IN1(
        \SUMB[758][2] ), .COUT(\CARRYB[759][1] ), .SUM(\SUMB[759][1] ) );
  FADDER S3_759_2 ( .CIN(\ab[759][2] ), .IN0(\CARRYB[758][2] ), .IN1(
        \ab[758][3] ), .COUT(\CARRYB[759][2] ), .SUM(\SUMB[759][2] ) );
  FADDER S1_758_0 ( .CIN(\ab[758][0] ), .IN0(\CARRYB[757][0] ), .IN1(
        \SUMB[757][1] ), .COUT(\CARRYB[758][0] ), .SUM(PRODUCT[758]) );
  FADDER S2_758_1 ( .CIN(\ab[758][1] ), .IN0(\CARRYB[757][1] ), .IN1(
        \SUMB[757][2] ), .COUT(\CARRYB[758][1] ), .SUM(\SUMB[758][1] ) );
  FADDER S3_758_2 ( .CIN(\ab[758][2] ), .IN0(\CARRYB[757][2] ), .IN1(
        \ab[757][3] ), .COUT(\CARRYB[758][2] ), .SUM(\SUMB[758][2] ) );
  FADDER S1_757_0 ( .CIN(\ab[757][0] ), .IN0(\CARRYB[756][0] ), .IN1(
        \SUMB[756][1] ), .COUT(\CARRYB[757][0] ), .SUM(PRODUCT[757]) );
  FADDER S2_757_1 ( .CIN(\ab[757][1] ), .IN0(\CARRYB[756][1] ), .IN1(
        \SUMB[756][2] ), .COUT(\CARRYB[757][1] ), .SUM(\SUMB[757][1] ) );
  FADDER S3_757_2 ( .CIN(\ab[757][2] ), .IN0(\CARRYB[756][2] ), .IN1(
        \ab[756][3] ), .COUT(\CARRYB[757][2] ), .SUM(\SUMB[757][2] ) );
  FADDER S1_756_0 ( .CIN(\ab[756][0] ), .IN0(\CARRYB[755][0] ), .IN1(
        \SUMB[755][1] ), .COUT(\CARRYB[756][0] ), .SUM(PRODUCT[756]) );
  FADDER S2_756_1 ( .CIN(\ab[756][1] ), .IN0(\CARRYB[755][1] ), .IN1(
        \SUMB[755][2] ), .COUT(\CARRYB[756][1] ), .SUM(\SUMB[756][1] ) );
  FADDER S3_756_2 ( .CIN(\ab[756][2] ), .IN0(\CARRYB[755][2] ), .IN1(
        \ab[755][3] ), .COUT(\CARRYB[756][2] ), .SUM(\SUMB[756][2] ) );
  FADDER S1_755_0 ( .CIN(\ab[755][0] ), .IN0(\CARRYB[754][0] ), .IN1(
        \SUMB[754][1] ), .COUT(\CARRYB[755][0] ), .SUM(PRODUCT[755]) );
  FADDER S2_755_1 ( .CIN(\ab[755][1] ), .IN0(\CARRYB[754][1] ), .IN1(
        \SUMB[754][2] ), .COUT(\CARRYB[755][1] ), .SUM(\SUMB[755][1] ) );
  FADDER S3_755_2 ( .CIN(\ab[755][2] ), .IN0(\CARRYB[754][2] ), .IN1(
        \ab[754][3] ), .COUT(\CARRYB[755][2] ), .SUM(\SUMB[755][2] ) );
  FADDER S1_754_0 ( .CIN(\ab[754][0] ), .IN0(\CARRYB[753][0] ), .IN1(
        \SUMB[753][1] ), .COUT(\CARRYB[754][0] ), .SUM(PRODUCT[754]) );
  FADDER S2_754_1 ( .CIN(\ab[754][1] ), .IN0(\CARRYB[753][1] ), .IN1(
        \SUMB[753][2] ), .COUT(\CARRYB[754][1] ), .SUM(\SUMB[754][1] ) );
  FADDER S3_754_2 ( .CIN(\ab[754][2] ), .IN0(\CARRYB[753][2] ), .IN1(
        \ab[753][3] ), .COUT(\CARRYB[754][2] ), .SUM(\SUMB[754][2] ) );
  FADDER S1_753_0 ( .CIN(\ab[753][0] ), .IN0(\CARRYB[752][0] ), .IN1(
        \SUMB[752][1] ), .COUT(\CARRYB[753][0] ), .SUM(PRODUCT[753]) );
  FADDER S2_753_1 ( .CIN(\ab[753][1] ), .IN0(\CARRYB[752][1] ), .IN1(
        \SUMB[752][2] ), .COUT(\CARRYB[753][1] ), .SUM(\SUMB[753][1] ) );
  FADDER S3_753_2 ( .CIN(\ab[753][2] ), .IN0(\CARRYB[752][2] ), .IN1(
        \ab[752][3] ), .COUT(\CARRYB[753][2] ), .SUM(\SUMB[753][2] ) );
  FADDER S1_752_0 ( .CIN(\ab[752][0] ), .IN0(\CARRYB[751][0] ), .IN1(
        \SUMB[751][1] ), .COUT(\CARRYB[752][0] ), .SUM(PRODUCT[752]) );
  FADDER S2_752_1 ( .CIN(\ab[752][1] ), .IN0(\CARRYB[751][1] ), .IN1(
        \SUMB[751][2] ), .COUT(\CARRYB[752][1] ), .SUM(\SUMB[752][1] ) );
  FADDER S3_752_2 ( .CIN(\ab[752][2] ), .IN0(\CARRYB[751][2] ), .IN1(
        \ab[751][3] ), .COUT(\CARRYB[752][2] ), .SUM(\SUMB[752][2] ) );
  FADDER S1_751_0 ( .CIN(\ab[751][0] ), .IN0(\CARRYB[750][0] ), .IN1(
        \SUMB[750][1] ), .COUT(\CARRYB[751][0] ), .SUM(PRODUCT[751]) );
  FADDER S2_751_1 ( .CIN(\ab[751][1] ), .IN0(\CARRYB[750][1] ), .IN1(
        \SUMB[750][2] ), .COUT(\CARRYB[751][1] ), .SUM(\SUMB[751][1] ) );
  FADDER S3_751_2 ( .CIN(\ab[751][2] ), .IN0(\CARRYB[750][2] ), .IN1(
        \ab[750][3] ), .COUT(\CARRYB[751][2] ), .SUM(\SUMB[751][2] ) );
  FADDER S1_750_0 ( .CIN(\ab[750][0] ), .IN0(\CARRYB[749][0] ), .IN1(
        \SUMB[749][1] ), .COUT(\CARRYB[750][0] ), .SUM(PRODUCT[750]) );
  FADDER S2_750_1 ( .CIN(\ab[750][1] ), .IN0(\CARRYB[749][1] ), .IN1(
        \SUMB[749][2] ), .COUT(\CARRYB[750][1] ), .SUM(\SUMB[750][1] ) );
  FADDER S3_750_2 ( .CIN(\ab[750][2] ), .IN0(\CARRYB[749][2] ), .IN1(
        \ab[749][3] ), .COUT(\CARRYB[750][2] ), .SUM(\SUMB[750][2] ) );
  FADDER S1_749_0 ( .CIN(\ab[749][0] ), .IN0(\CARRYB[748][0] ), .IN1(
        \SUMB[748][1] ), .COUT(\CARRYB[749][0] ), .SUM(PRODUCT[749]) );
  FADDER S2_749_1 ( .CIN(\ab[749][1] ), .IN0(\CARRYB[748][1] ), .IN1(
        \SUMB[748][2] ), .COUT(\CARRYB[749][1] ), .SUM(\SUMB[749][1] ) );
  FADDER S3_749_2 ( .CIN(\ab[749][2] ), .IN0(\CARRYB[748][2] ), .IN1(
        \ab[748][3] ), .COUT(\CARRYB[749][2] ), .SUM(\SUMB[749][2] ) );
  FADDER S1_748_0 ( .CIN(\ab[748][0] ), .IN0(\CARRYB[747][0] ), .IN1(
        \SUMB[747][1] ), .COUT(\CARRYB[748][0] ), .SUM(PRODUCT[748]) );
  FADDER S2_748_1 ( .CIN(\ab[748][1] ), .IN0(\CARRYB[747][1] ), .IN1(
        \SUMB[747][2] ), .COUT(\CARRYB[748][1] ), .SUM(\SUMB[748][1] ) );
  FADDER S3_748_2 ( .CIN(\ab[748][2] ), .IN0(\CARRYB[747][2] ), .IN1(
        \ab[747][3] ), .COUT(\CARRYB[748][2] ), .SUM(\SUMB[748][2] ) );
  FADDER S1_747_0 ( .CIN(\ab[747][0] ), .IN0(\CARRYB[746][0] ), .IN1(
        \SUMB[746][1] ), .COUT(\CARRYB[747][0] ), .SUM(PRODUCT[747]) );
  FADDER S2_747_1 ( .CIN(\ab[747][1] ), .IN0(\CARRYB[746][1] ), .IN1(
        \SUMB[746][2] ), .COUT(\CARRYB[747][1] ), .SUM(\SUMB[747][1] ) );
  FADDER S3_747_2 ( .CIN(\ab[747][2] ), .IN0(\CARRYB[746][2] ), .IN1(
        \ab[746][3] ), .COUT(\CARRYB[747][2] ), .SUM(\SUMB[747][2] ) );
  FADDER S1_746_0 ( .CIN(\ab[746][0] ), .IN0(\CARRYB[745][0] ), .IN1(
        \SUMB[745][1] ), .COUT(\CARRYB[746][0] ), .SUM(PRODUCT[746]) );
  FADDER S2_746_1 ( .CIN(\ab[746][1] ), .IN0(\CARRYB[745][1] ), .IN1(
        \SUMB[745][2] ), .COUT(\CARRYB[746][1] ), .SUM(\SUMB[746][1] ) );
  FADDER S3_746_2 ( .CIN(\ab[746][2] ), .IN0(\CARRYB[745][2] ), .IN1(
        \ab[745][3] ), .COUT(\CARRYB[746][2] ), .SUM(\SUMB[746][2] ) );
  FADDER S1_745_0 ( .CIN(\ab[745][0] ), .IN0(\CARRYB[744][0] ), .IN1(
        \SUMB[744][1] ), .COUT(\CARRYB[745][0] ), .SUM(PRODUCT[745]) );
  FADDER S2_745_1 ( .CIN(\ab[745][1] ), .IN0(\CARRYB[744][1] ), .IN1(
        \SUMB[744][2] ), .COUT(\CARRYB[745][1] ), .SUM(\SUMB[745][1] ) );
  FADDER S3_745_2 ( .CIN(\ab[745][2] ), .IN0(\CARRYB[744][2] ), .IN1(
        \ab[744][3] ), .COUT(\CARRYB[745][2] ), .SUM(\SUMB[745][2] ) );
  FADDER S1_744_0 ( .CIN(\ab[744][0] ), .IN0(\CARRYB[743][0] ), .IN1(
        \SUMB[743][1] ), .COUT(\CARRYB[744][0] ), .SUM(PRODUCT[744]) );
  FADDER S2_744_1 ( .CIN(\ab[744][1] ), .IN0(\CARRYB[743][1] ), .IN1(
        \SUMB[743][2] ), .COUT(\CARRYB[744][1] ), .SUM(\SUMB[744][1] ) );
  FADDER S3_744_2 ( .CIN(\ab[744][2] ), .IN0(\CARRYB[743][2] ), .IN1(
        \ab[743][3] ), .COUT(\CARRYB[744][2] ), .SUM(\SUMB[744][2] ) );
  FADDER S1_743_0 ( .CIN(\ab[743][0] ), .IN0(\CARRYB[742][0] ), .IN1(
        \SUMB[742][1] ), .COUT(\CARRYB[743][0] ), .SUM(PRODUCT[743]) );
  FADDER S2_743_1 ( .CIN(\ab[743][1] ), .IN0(\CARRYB[742][1] ), .IN1(
        \SUMB[742][2] ), .COUT(\CARRYB[743][1] ), .SUM(\SUMB[743][1] ) );
  FADDER S3_743_2 ( .CIN(\ab[743][2] ), .IN0(\CARRYB[742][2] ), .IN1(
        \ab[742][3] ), .COUT(\CARRYB[743][2] ), .SUM(\SUMB[743][2] ) );
  FADDER S1_742_0 ( .CIN(\ab[742][0] ), .IN0(\CARRYB[741][0] ), .IN1(
        \SUMB[741][1] ), .COUT(\CARRYB[742][0] ), .SUM(PRODUCT[742]) );
  FADDER S2_742_1 ( .CIN(\ab[742][1] ), .IN0(\CARRYB[741][1] ), .IN1(
        \SUMB[741][2] ), .COUT(\CARRYB[742][1] ), .SUM(\SUMB[742][1] ) );
  FADDER S3_742_2 ( .CIN(\ab[742][2] ), .IN0(\CARRYB[741][2] ), .IN1(
        \ab[741][3] ), .COUT(\CARRYB[742][2] ), .SUM(\SUMB[742][2] ) );
  FADDER S1_741_0 ( .CIN(\ab[741][0] ), .IN0(\CARRYB[740][0] ), .IN1(
        \SUMB[740][1] ), .COUT(\CARRYB[741][0] ), .SUM(PRODUCT[741]) );
  FADDER S2_741_1 ( .CIN(\ab[741][1] ), .IN0(\CARRYB[740][1] ), .IN1(
        \SUMB[740][2] ), .COUT(\CARRYB[741][1] ), .SUM(\SUMB[741][1] ) );
  FADDER S3_741_2 ( .CIN(\ab[741][2] ), .IN0(\CARRYB[740][2] ), .IN1(
        \ab[740][3] ), .COUT(\CARRYB[741][2] ), .SUM(\SUMB[741][2] ) );
  FADDER S1_740_0 ( .CIN(\ab[740][0] ), .IN0(\CARRYB[739][0] ), .IN1(
        \SUMB[739][1] ), .COUT(\CARRYB[740][0] ), .SUM(PRODUCT[740]) );
  FADDER S2_740_1 ( .CIN(\ab[740][1] ), .IN0(\CARRYB[739][1] ), .IN1(
        \SUMB[739][2] ), .COUT(\CARRYB[740][1] ), .SUM(\SUMB[740][1] ) );
  FADDER S3_740_2 ( .CIN(\ab[740][2] ), .IN0(\CARRYB[739][2] ), .IN1(
        \ab[739][3] ), .COUT(\CARRYB[740][2] ), .SUM(\SUMB[740][2] ) );
  FADDER S1_739_0 ( .CIN(\ab[739][0] ), .IN0(\CARRYB[738][0] ), .IN1(
        \SUMB[738][1] ), .COUT(\CARRYB[739][0] ), .SUM(PRODUCT[739]) );
  FADDER S2_739_1 ( .CIN(\ab[739][1] ), .IN0(\CARRYB[738][1] ), .IN1(
        \SUMB[738][2] ), .COUT(\CARRYB[739][1] ), .SUM(\SUMB[739][1] ) );
  FADDER S3_739_2 ( .CIN(\ab[739][2] ), .IN0(\CARRYB[738][2] ), .IN1(
        \ab[738][3] ), .COUT(\CARRYB[739][2] ), .SUM(\SUMB[739][2] ) );
  FADDER S1_738_0 ( .CIN(\ab[738][0] ), .IN0(\CARRYB[737][0] ), .IN1(
        \SUMB[737][1] ), .COUT(\CARRYB[738][0] ), .SUM(PRODUCT[738]) );
  FADDER S2_738_1 ( .CIN(\ab[738][1] ), .IN0(\CARRYB[737][1] ), .IN1(
        \SUMB[737][2] ), .COUT(\CARRYB[738][1] ), .SUM(\SUMB[738][1] ) );
  FADDER S3_738_2 ( .CIN(\ab[738][2] ), .IN0(\CARRYB[737][2] ), .IN1(
        \ab[737][3] ), .COUT(\CARRYB[738][2] ), .SUM(\SUMB[738][2] ) );
  FADDER S1_737_0 ( .CIN(\ab[737][0] ), .IN0(\CARRYB[736][0] ), .IN1(
        \SUMB[736][1] ), .COUT(\CARRYB[737][0] ), .SUM(PRODUCT[737]) );
  FADDER S2_737_1 ( .CIN(\ab[737][1] ), .IN0(\CARRYB[736][1] ), .IN1(
        \SUMB[736][2] ), .COUT(\CARRYB[737][1] ), .SUM(\SUMB[737][1] ) );
  FADDER S3_737_2 ( .CIN(\ab[737][2] ), .IN0(\CARRYB[736][2] ), .IN1(
        \ab[736][3] ), .COUT(\CARRYB[737][2] ), .SUM(\SUMB[737][2] ) );
  FADDER S1_736_0 ( .CIN(\ab[736][0] ), .IN0(\CARRYB[735][0] ), .IN1(
        \SUMB[735][1] ), .COUT(\CARRYB[736][0] ), .SUM(PRODUCT[736]) );
  FADDER S2_736_1 ( .CIN(\ab[736][1] ), .IN0(\CARRYB[735][1] ), .IN1(
        \SUMB[735][2] ), .COUT(\CARRYB[736][1] ), .SUM(\SUMB[736][1] ) );
  FADDER S3_736_2 ( .CIN(\ab[736][2] ), .IN0(\CARRYB[735][2] ), .IN1(
        \ab[735][3] ), .COUT(\CARRYB[736][2] ), .SUM(\SUMB[736][2] ) );
  FADDER S1_735_0 ( .CIN(\ab[735][0] ), .IN0(\CARRYB[734][0] ), .IN1(
        \SUMB[734][1] ), .COUT(\CARRYB[735][0] ), .SUM(PRODUCT[735]) );
  FADDER S2_735_1 ( .CIN(\ab[735][1] ), .IN0(\CARRYB[734][1] ), .IN1(
        \SUMB[734][2] ), .COUT(\CARRYB[735][1] ), .SUM(\SUMB[735][1] ) );
  FADDER S3_735_2 ( .CIN(\ab[735][2] ), .IN0(\CARRYB[734][2] ), .IN1(
        \ab[734][3] ), .COUT(\CARRYB[735][2] ), .SUM(\SUMB[735][2] ) );
  FADDER S1_734_0 ( .CIN(\ab[734][0] ), .IN0(\CARRYB[733][0] ), .IN1(
        \SUMB[733][1] ), .COUT(\CARRYB[734][0] ), .SUM(PRODUCT[734]) );
  FADDER S2_734_1 ( .CIN(\ab[734][1] ), .IN0(\CARRYB[733][1] ), .IN1(
        \SUMB[733][2] ), .COUT(\CARRYB[734][1] ), .SUM(\SUMB[734][1] ) );
  FADDER S3_734_2 ( .CIN(\ab[734][2] ), .IN0(\CARRYB[733][2] ), .IN1(
        \ab[733][3] ), .COUT(\CARRYB[734][2] ), .SUM(\SUMB[734][2] ) );
  FADDER S1_733_0 ( .CIN(\ab[733][0] ), .IN0(\CARRYB[732][0] ), .IN1(
        \SUMB[732][1] ), .COUT(\CARRYB[733][0] ), .SUM(PRODUCT[733]) );
  FADDER S2_733_1 ( .CIN(\ab[733][1] ), .IN0(\CARRYB[732][1] ), .IN1(
        \SUMB[732][2] ), .COUT(\CARRYB[733][1] ), .SUM(\SUMB[733][1] ) );
  FADDER S3_733_2 ( .CIN(\ab[733][2] ), .IN0(\CARRYB[732][2] ), .IN1(
        \ab[732][3] ), .COUT(\CARRYB[733][2] ), .SUM(\SUMB[733][2] ) );
  FADDER S1_732_0 ( .CIN(\ab[732][0] ), .IN0(\CARRYB[731][0] ), .IN1(
        \SUMB[731][1] ), .COUT(\CARRYB[732][0] ), .SUM(PRODUCT[732]) );
  FADDER S2_732_1 ( .CIN(\ab[732][1] ), .IN0(\CARRYB[731][1] ), .IN1(
        \SUMB[731][2] ), .COUT(\CARRYB[732][1] ), .SUM(\SUMB[732][1] ) );
  FADDER S3_732_2 ( .CIN(\ab[732][2] ), .IN0(\CARRYB[731][2] ), .IN1(
        \ab[731][3] ), .COUT(\CARRYB[732][2] ), .SUM(\SUMB[732][2] ) );
  FADDER S1_731_0 ( .CIN(\ab[731][0] ), .IN0(\CARRYB[730][0] ), .IN1(
        \SUMB[730][1] ), .COUT(\CARRYB[731][0] ), .SUM(PRODUCT[731]) );
  FADDER S2_731_1 ( .CIN(\ab[731][1] ), .IN0(\CARRYB[730][1] ), .IN1(
        \SUMB[730][2] ), .COUT(\CARRYB[731][1] ), .SUM(\SUMB[731][1] ) );
  FADDER S3_731_2 ( .CIN(\ab[731][2] ), .IN0(\CARRYB[730][2] ), .IN1(
        \ab[730][3] ), .COUT(\CARRYB[731][2] ), .SUM(\SUMB[731][2] ) );
  FADDER S1_730_0 ( .CIN(\ab[730][0] ), .IN0(\CARRYB[729][0] ), .IN1(
        \SUMB[729][1] ), .COUT(\CARRYB[730][0] ), .SUM(PRODUCT[730]) );
  FADDER S2_730_1 ( .CIN(\ab[730][1] ), .IN0(\CARRYB[729][1] ), .IN1(
        \SUMB[729][2] ), .COUT(\CARRYB[730][1] ), .SUM(\SUMB[730][1] ) );
  FADDER S3_730_2 ( .CIN(\ab[730][2] ), .IN0(\CARRYB[729][2] ), .IN1(
        \ab[729][3] ), .COUT(\CARRYB[730][2] ), .SUM(\SUMB[730][2] ) );
  FADDER S1_729_0 ( .CIN(\ab[729][0] ), .IN0(\CARRYB[728][0] ), .IN1(
        \SUMB[728][1] ), .COUT(\CARRYB[729][0] ), .SUM(PRODUCT[729]) );
  FADDER S2_729_1 ( .CIN(\ab[729][1] ), .IN0(\CARRYB[728][1] ), .IN1(
        \SUMB[728][2] ), .COUT(\CARRYB[729][1] ), .SUM(\SUMB[729][1] ) );
  FADDER S3_729_2 ( .CIN(\ab[729][2] ), .IN0(\CARRYB[728][2] ), .IN1(
        \ab[728][3] ), .COUT(\CARRYB[729][2] ), .SUM(\SUMB[729][2] ) );
  FADDER S1_728_0 ( .CIN(\ab[728][0] ), .IN0(\CARRYB[727][0] ), .IN1(
        \SUMB[727][1] ), .COUT(\CARRYB[728][0] ), .SUM(PRODUCT[728]) );
  FADDER S2_728_1 ( .CIN(\ab[728][1] ), .IN0(\CARRYB[727][1] ), .IN1(
        \SUMB[727][2] ), .COUT(\CARRYB[728][1] ), .SUM(\SUMB[728][1] ) );
  FADDER S3_728_2 ( .CIN(\ab[728][2] ), .IN0(\CARRYB[727][2] ), .IN1(
        \ab[727][3] ), .COUT(\CARRYB[728][2] ), .SUM(\SUMB[728][2] ) );
  FADDER S1_727_0 ( .CIN(\ab[727][0] ), .IN0(\CARRYB[726][0] ), .IN1(
        \SUMB[726][1] ), .COUT(\CARRYB[727][0] ), .SUM(PRODUCT[727]) );
  FADDER S2_727_1 ( .CIN(\ab[727][1] ), .IN0(\CARRYB[726][1] ), .IN1(
        \SUMB[726][2] ), .COUT(\CARRYB[727][1] ), .SUM(\SUMB[727][1] ) );
  FADDER S3_727_2 ( .CIN(\ab[727][2] ), .IN0(\CARRYB[726][2] ), .IN1(
        \ab[726][3] ), .COUT(\CARRYB[727][2] ), .SUM(\SUMB[727][2] ) );
  FADDER S1_726_0 ( .CIN(\ab[726][0] ), .IN0(\CARRYB[725][0] ), .IN1(
        \SUMB[725][1] ), .COUT(\CARRYB[726][0] ), .SUM(PRODUCT[726]) );
  FADDER S2_726_1 ( .CIN(\ab[726][1] ), .IN0(\CARRYB[725][1] ), .IN1(
        \SUMB[725][2] ), .COUT(\CARRYB[726][1] ), .SUM(\SUMB[726][1] ) );
  FADDER S3_726_2 ( .CIN(\ab[726][2] ), .IN0(\CARRYB[725][2] ), .IN1(
        \ab[725][3] ), .COUT(\CARRYB[726][2] ), .SUM(\SUMB[726][2] ) );
  FADDER S1_725_0 ( .CIN(\ab[725][0] ), .IN0(\CARRYB[724][0] ), .IN1(
        \SUMB[724][1] ), .COUT(\CARRYB[725][0] ), .SUM(PRODUCT[725]) );
  FADDER S2_725_1 ( .CIN(\ab[725][1] ), .IN0(\CARRYB[724][1] ), .IN1(
        \SUMB[724][2] ), .COUT(\CARRYB[725][1] ), .SUM(\SUMB[725][1] ) );
  FADDER S3_725_2 ( .CIN(\ab[725][2] ), .IN0(\CARRYB[724][2] ), .IN1(
        \ab[724][3] ), .COUT(\CARRYB[725][2] ), .SUM(\SUMB[725][2] ) );
  FADDER S1_724_0 ( .CIN(\ab[724][0] ), .IN0(\CARRYB[723][0] ), .IN1(
        \SUMB[723][1] ), .COUT(\CARRYB[724][0] ), .SUM(PRODUCT[724]) );
  FADDER S2_724_1 ( .CIN(\ab[724][1] ), .IN0(\CARRYB[723][1] ), .IN1(
        \SUMB[723][2] ), .COUT(\CARRYB[724][1] ), .SUM(\SUMB[724][1] ) );
  FADDER S3_724_2 ( .CIN(\ab[724][2] ), .IN0(\CARRYB[723][2] ), .IN1(
        \ab[723][3] ), .COUT(\CARRYB[724][2] ), .SUM(\SUMB[724][2] ) );
  FADDER S1_723_0 ( .CIN(\ab[723][0] ), .IN0(\CARRYB[722][0] ), .IN1(
        \SUMB[722][1] ), .COUT(\CARRYB[723][0] ), .SUM(PRODUCT[723]) );
  FADDER S2_723_1 ( .CIN(\ab[723][1] ), .IN0(\CARRYB[722][1] ), .IN1(
        \SUMB[722][2] ), .COUT(\CARRYB[723][1] ), .SUM(\SUMB[723][1] ) );
  FADDER S3_723_2 ( .CIN(\ab[723][2] ), .IN0(\CARRYB[722][2] ), .IN1(
        \ab[722][3] ), .COUT(\CARRYB[723][2] ), .SUM(\SUMB[723][2] ) );
  FADDER S1_722_0 ( .CIN(\ab[722][0] ), .IN0(\CARRYB[721][0] ), .IN1(
        \SUMB[721][1] ), .COUT(\CARRYB[722][0] ), .SUM(PRODUCT[722]) );
  FADDER S2_722_1 ( .CIN(\ab[722][1] ), .IN0(\CARRYB[721][1] ), .IN1(
        \SUMB[721][2] ), .COUT(\CARRYB[722][1] ), .SUM(\SUMB[722][1] ) );
  FADDER S3_722_2 ( .CIN(\ab[722][2] ), .IN0(\CARRYB[721][2] ), .IN1(
        \ab[721][3] ), .COUT(\CARRYB[722][2] ), .SUM(\SUMB[722][2] ) );
  FADDER S1_721_0 ( .CIN(\ab[721][0] ), .IN0(\CARRYB[720][0] ), .IN1(
        \SUMB[720][1] ), .COUT(\CARRYB[721][0] ), .SUM(PRODUCT[721]) );
  FADDER S2_721_1 ( .CIN(\ab[721][1] ), .IN0(\CARRYB[720][1] ), .IN1(
        \SUMB[720][2] ), .COUT(\CARRYB[721][1] ), .SUM(\SUMB[721][1] ) );
  FADDER S3_721_2 ( .CIN(\ab[721][2] ), .IN0(\CARRYB[720][2] ), .IN1(
        \ab[720][3] ), .COUT(\CARRYB[721][2] ), .SUM(\SUMB[721][2] ) );
  FADDER S1_720_0 ( .CIN(\ab[720][0] ), .IN0(\CARRYB[719][0] ), .IN1(
        \SUMB[719][1] ), .COUT(\CARRYB[720][0] ), .SUM(PRODUCT[720]) );
  FADDER S2_720_1 ( .CIN(\ab[720][1] ), .IN0(\CARRYB[719][1] ), .IN1(
        \SUMB[719][2] ), .COUT(\CARRYB[720][1] ), .SUM(\SUMB[720][1] ) );
  FADDER S3_720_2 ( .CIN(\ab[720][2] ), .IN0(\CARRYB[719][2] ), .IN1(
        \ab[719][3] ), .COUT(\CARRYB[720][2] ), .SUM(\SUMB[720][2] ) );
  FADDER S1_719_0 ( .CIN(\ab[719][0] ), .IN0(\CARRYB[718][0] ), .IN1(
        \SUMB[718][1] ), .COUT(\CARRYB[719][0] ), .SUM(PRODUCT[719]) );
  FADDER S2_719_1 ( .CIN(\ab[719][1] ), .IN0(\CARRYB[718][1] ), .IN1(
        \SUMB[718][2] ), .COUT(\CARRYB[719][1] ), .SUM(\SUMB[719][1] ) );
  FADDER S3_719_2 ( .CIN(\ab[719][2] ), .IN0(\CARRYB[718][2] ), .IN1(
        \ab[718][3] ), .COUT(\CARRYB[719][2] ), .SUM(\SUMB[719][2] ) );
  FADDER S1_718_0 ( .CIN(\ab[718][0] ), .IN0(\CARRYB[717][0] ), .IN1(
        \SUMB[717][1] ), .COUT(\CARRYB[718][0] ), .SUM(PRODUCT[718]) );
  FADDER S2_718_1 ( .CIN(\ab[718][1] ), .IN0(\CARRYB[717][1] ), .IN1(
        \SUMB[717][2] ), .COUT(\CARRYB[718][1] ), .SUM(\SUMB[718][1] ) );
  FADDER S3_718_2 ( .CIN(\ab[718][2] ), .IN0(\CARRYB[717][2] ), .IN1(
        \ab[717][3] ), .COUT(\CARRYB[718][2] ), .SUM(\SUMB[718][2] ) );
  FADDER S1_717_0 ( .CIN(\ab[717][0] ), .IN0(\CARRYB[716][0] ), .IN1(
        \SUMB[716][1] ), .COUT(\CARRYB[717][0] ), .SUM(PRODUCT[717]) );
  FADDER S2_717_1 ( .CIN(\ab[717][1] ), .IN0(\CARRYB[716][1] ), .IN1(
        \SUMB[716][2] ), .COUT(\CARRYB[717][1] ), .SUM(\SUMB[717][1] ) );
  FADDER S3_717_2 ( .CIN(\ab[717][2] ), .IN0(\CARRYB[716][2] ), .IN1(
        \ab[716][3] ), .COUT(\CARRYB[717][2] ), .SUM(\SUMB[717][2] ) );
  FADDER S1_716_0 ( .CIN(\ab[716][0] ), .IN0(\CARRYB[715][0] ), .IN1(
        \SUMB[715][1] ), .COUT(\CARRYB[716][0] ), .SUM(PRODUCT[716]) );
  FADDER S2_716_1 ( .CIN(\ab[716][1] ), .IN0(\CARRYB[715][1] ), .IN1(
        \SUMB[715][2] ), .COUT(\CARRYB[716][1] ), .SUM(\SUMB[716][1] ) );
  FADDER S3_716_2 ( .CIN(\ab[716][2] ), .IN0(\CARRYB[715][2] ), .IN1(
        \ab[715][3] ), .COUT(\CARRYB[716][2] ), .SUM(\SUMB[716][2] ) );
  FADDER S1_715_0 ( .CIN(\ab[715][0] ), .IN0(\CARRYB[714][0] ), .IN1(
        \SUMB[714][1] ), .COUT(\CARRYB[715][0] ), .SUM(PRODUCT[715]) );
  FADDER S2_715_1 ( .CIN(\ab[715][1] ), .IN0(\CARRYB[714][1] ), .IN1(
        \SUMB[714][2] ), .COUT(\CARRYB[715][1] ), .SUM(\SUMB[715][1] ) );
  FADDER S3_715_2 ( .CIN(\ab[715][2] ), .IN0(\CARRYB[714][2] ), .IN1(
        \ab[714][3] ), .COUT(\CARRYB[715][2] ), .SUM(\SUMB[715][2] ) );
  FADDER S1_714_0 ( .CIN(\ab[714][0] ), .IN0(\CARRYB[713][0] ), .IN1(
        \SUMB[713][1] ), .COUT(\CARRYB[714][0] ), .SUM(PRODUCT[714]) );
  FADDER S2_714_1 ( .CIN(\ab[714][1] ), .IN0(\CARRYB[713][1] ), .IN1(
        \SUMB[713][2] ), .COUT(\CARRYB[714][1] ), .SUM(\SUMB[714][1] ) );
  FADDER S3_714_2 ( .CIN(\ab[714][2] ), .IN0(\CARRYB[713][2] ), .IN1(
        \ab[713][3] ), .COUT(\CARRYB[714][2] ), .SUM(\SUMB[714][2] ) );
  FADDER S1_713_0 ( .CIN(\ab[713][0] ), .IN0(\CARRYB[712][0] ), .IN1(
        \SUMB[712][1] ), .COUT(\CARRYB[713][0] ), .SUM(PRODUCT[713]) );
  FADDER S2_713_1 ( .CIN(\ab[713][1] ), .IN0(\CARRYB[712][1] ), .IN1(
        \SUMB[712][2] ), .COUT(\CARRYB[713][1] ), .SUM(\SUMB[713][1] ) );
  FADDER S3_713_2 ( .CIN(\ab[713][2] ), .IN0(\CARRYB[712][2] ), .IN1(
        \ab[712][3] ), .COUT(\CARRYB[713][2] ), .SUM(\SUMB[713][2] ) );
  FADDER S1_712_0 ( .CIN(\ab[712][0] ), .IN0(\CARRYB[711][0] ), .IN1(
        \SUMB[711][1] ), .COUT(\CARRYB[712][0] ), .SUM(PRODUCT[712]) );
  FADDER S2_712_1 ( .CIN(\ab[712][1] ), .IN0(\CARRYB[711][1] ), .IN1(
        \SUMB[711][2] ), .COUT(\CARRYB[712][1] ), .SUM(\SUMB[712][1] ) );
  FADDER S3_712_2 ( .CIN(\ab[712][2] ), .IN0(\CARRYB[711][2] ), .IN1(
        \ab[711][3] ), .COUT(\CARRYB[712][2] ), .SUM(\SUMB[712][2] ) );
  FADDER S1_711_0 ( .CIN(\ab[711][0] ), .IN0(\CARRYB[710][0] ), .IN1(
        \SUMB[710][1] ), .COUT(\CARRYB[711][0] ), .SUM(PRODUCT[711]) );
  FADDER S2_711_1 ( .CIN(\ab[711][1] ), .IN0(\CARRYB[710][1] ), .IN1(
        \SUMB[710][2] ), .COUT(\CARRYB[711][1] ), .SUM(\SUMB[711][1] ) );
  FADDER S3_711_2 ( .CIN(\ab[711][2] ), .IN0(\CARRYB[710][2] ), .IN1(
        \ab[710][3] ), .COUT(\CARRYB[711][2] ), .SUM(\SUMB[711][2] ) );
  FADDER S1_710_0 ( .CIN(\ab[710][0] ), .IN0(\CARRYB[709][0] ), .IN1(
        \SUMB[709][1] ), .COUT(\CARRYB[710][0] ), .SUM(PRODUCT[710]) );
  FADDER S2_710_1 ( .CIN(\ab[710][1] ), .IN0(\CARRYB[709][1] ), .IN1(
        \SUMB[709][2] ), .COUT(\CARRYB[710][1] ), .SUM(\SUMB[710][1] ) );
  FADDER S3_710_2 ( .CIN(\ab[710][2] ), .IN0(\CARRYB[709][2] ), .IN1(
        \ab[709][3] ), .COUT(\CARRYB[710][2] ), .SUM(\SUMB[710][2] ) );
  FADDER S1_709_0 ( .CIN(\ab[709][0] ), .IN0(\CARRYB[708][0] ), .IN1(
        \SUMB[708][1] ), .COUT(\CARRYB[709][0] ), .SUM(PRODUCT[709]) );
  FADDER S2_709_1 ( .CIN(\ab[709][1] ), .IN0(\CARRYB[708][1] ), .IN1(
        \SUMB[708][2] ), .COUT(\CARRYB[709][1] ), .SUM(\SUMB[709][1] ) );
  FADDER S3_709_2 ( .CIN(\ab[709][2] ), .IN0(\CARRYB[708][2] ), .IN1(
        \ab[708][3] ), .COUT(\CARRYB[709][2] ), .SUM(\SUMB[709][2] ) );
  FADDER S1_708_0 ( .CIN(\ab[708][0] ), .IN0(\CARRYB[707][0] ), .IN1(
        \SUMB[707][1] ), .COUT(\CARRYB[708][0] ), .SUM(PRODUCT[708]) );
  FADDER S2_708_1 ( .CIN(\ab[708][1] ), .IN0(\CARRYB[707][1] ), .IN1(
        \SUMB[707][2] ), .COUT(\CARRYB[708][1] ), .SUM(\SUMB[708][1] ) );
  FADDER S3_708_2 ( .CIN(\ab[708][2] ), .IN0(\CARRYB[707][2] ), .IN1(
        \ab[707][3] ), .COUT(\CARRYB[708][2] ), .SUM(\SUMB[708][2] ) );
  FADDER S1_707_0 ( .CIN(\ab[707][0] ), .IN0(\CARRYB[706][0] ), .IN1(
        \SUMB[706][1] ), .COUT(\CARRYB[707][0] ), .SUM(PRODUCT[707]) );
  FADDER S2_707_1 ( .CIN(\ab[707][1] ), .IN0(\CARRYB[706][1] ), .IN1(
        \SUMB[706][2] ), .COUT(\CARRYB[707][1] ), .SUM(\SUMB[707][1] ) );
  FADDER S3_707_2 ( .CIN(\ab[707][2] ), .IN0(\CARRYB[706][2] ), .IN1(
        \ab[706][3] ), .COUT(\CARRYB[707][2] ), .SUM(\SUMB[707][2] ) );
  FADDER S1_706_0 ( .CIN(\ab[706][0] ), .IN0(\CARRYB[705][0] ), .IN1(
        \SUMB[705][1] ), .COUT(\CARRYB[706][0] ), .SUM(PRODUCT[706]) );
  FADDER S2_706_1 ( .CIN(\ab[706][1] ), .IN0(\CARRYB[705][1] ), .IN1(
        \SUMB[705][2] ), .COUT(\CARRYB[706][1] ), .SUM(\SUMB[706][1] ) );
  FADDER S3_706_2 ( .CIN(\ab[706][2] ), .IN0(\CARRYB[705][2] ), .IN1(
        \ab[705][3] ), .COUT(\CARRYB[706][2] ), .SUM(\SUMB[706][2] ) );
  FADDER S1_705_0 ( .CIN(\ab[705][0] ), .IN0(\CARRYB[704][0] ), .IN1(
        \SUMB[704][1] ), .COUT(\CARRYB[705][0] ), .SUM(PRODUCT[705]) );
  FADDER S2_705_1 ( .CIN(\ab[705][1] ), .IN0(\CARRYB[704][1] ), .IN1(
        \SUMB[704][2] ), .COUT(\CARRYB[705][1] ), .SUM(\SUMB[705][1] ) );
  FADDER S3_705_2 ( .CIN(\ab[705][2] ), .IN0(\CARRYB[704][2] ), .IN1(
        \ab[704][3] ), .COUT(\CARRYB[705][2] ), .SUM(\SUMB[705][2] ) );
  FADDER S1_704_0 ( .CIN(\ab[704][0] ), .IN0(\CARRYB[703][0] ), .IN1(
        \SUMB[703][1] ), .COUT(\CARRYB[704][0] ), .SUM(PRODUCT[704]) );
  FADDER S2_704_1 ( .CIN(\ab[704][1] ), .IN0(\CARRYB[703][1] ), .IN1(
        \SUMB[703][2] ), .COUT(\CARRYB[704][1] ), .SUM(\SUMB[704][1] ) );
  FADDER S3_704_2 ( .CIN(\ab[704][2] ), .IN0(\CARRYB[703][2] ), .IN1(
        \ab[703][3] ), .COUT(\CARRYB[704][2] ), .SUM(\SUMB[704][2] ) );
  FADDER S1_703_0 ( .CIN(\ab[703][0] ), .IN0(\CARRYB[702][0] ), .IN1(
        \SUMB[702][1] ), .COUT(\CARRYB[703][0] ), .SUM(PRODUCT[703]) );
  FADDER S2_703_1 ( .CIN(\ab[703][1] ), .IN0(\CARRYB[702][1] ), .IN1(
        \SUMB[702][2] ), .COUT(\CARRYB[703][1] ), .SUM(\SUMB[703][1] ) );
  FADDER S3_703_2 ( .CIN(\ab[703][2] ), .IN0(\CARRYB[702][2] ), .IN1(
        \ab[702][3] ), .COUT(\CARRYB[703][2] ), .SUM(\SUMB[703][2] ) );
  FADDER S1_702_0 ( .CIN(\ab[702][0] ), .IN0(\CARRYB[701][0] ), .IN1(
        \SUMB[701][1] ), .COUT(\CARRYB[702][0] ), .SUM(PRODUCT[702]) );
  FADDER S2_702_1 ( .CIN(\ab[702][1] ), .IN0(\CARRYB[701][1] ), .IN1(
        \SUMB[701][2] ), .COUT(\CARRYB[702][1] ), .SUM(\SUMB[702][1] ) );
  FADDER S3_702_2 ( .CIN(\ab[702][2] ), .IN0(\CARRYB[701][2] ), .IN1(
        \ab[701][3] ), .COUT(\CARRYB[702][2] ), .SUM(\SUMB[702][2] ) );
  FADDER S1_701_0 ( .CIN(\ab[701][0] ), .IN0(\CARRYB[700][0] ), .IN1(
        \SUMB[700][1] ), .COUT(\CARRYB[701][0] ), .SUM(PRODUCT[701]) );
  FADDER S2_701_1 ( .CIN(\ab[701][1] ), .IN0(\CARRYB[700][1] ), .IN1(
        \SUMB[700][2] ), .COUT(\CARRYB[701][1] ), .SUM(\SUMB[701][1] ) );
  FADDER S3_701_2 ( .CIN(\ab[701][2] ), .IN0(\CARRYB[700][2] ), .IN1(
        \ab[700][3] ), .COUT(\CARRYB[701][2] ), .SUM(\SUMB[701][2] ) );
  FADDER S1_700_0 ( .CIN(\ab[700][0] ), .IN0(\CARRYB[699][0] ), .IN1(
        \SUMB[699][1] ), .COUT(\CARRYB[700][0] ), .SUM(PRODUCT[700]) );
  FADDER S2_700_1 ( .CIN(\ab[700][1] ), .IN0(\CARRYB[699][1] ), .IN1(
        \SUMB[699][2] ), .COUT(\CARRYB[700][1] ), .SUM(\SUMB[700][1] ) );
  FADDER S3_700_2 ( .CIN(\ab[700][2] ), .IN0(\CARRYB[699][2] ), .IN1(
        \ab[699][3] ), .COUT(\CARRYB[700][2] ), .SUM(\SUMB[700][2] ) );
  FADDER S1_699_0 ( .CIN(\ab[699][0] ), .IN0(\CARRYB[698][0] ), .IN1(
        \SUMB[698][1] ), .COUT(\CARRYB[699][0] ), .SUM(PRODUCT[699]) );
  FADDER S2_699_1 ( .CIN(\ab[699][1] ), .IN0(\CARRYB[698][1] ), .IN1(
        \SUMB[698][2] ), .COUT(\CARRYB[699][1] ), .SUM(\SUMB[699][1] ) );
  FADDER S3_699_2 ( .CIN(\ab[699][2] ), .IN0(\CARRYB[698][2] ), .IN1(
        \ab[698][3] ), .COUT(\CARRYB[699][2] ), .SUM(\SUMB[699][2] ) );
  FADDER S1_698_0 ( .CIN(\ab[698][0] ), .IN0(\CARRYB[697][0] ), .IN1(
        \SUMB[697][1] ), .COUT(\CARRYB[698][0] ), .SUM(PRODUCT[698]) );
  FADDER S2_698_1 ( .CIN(\ab[698][1] ), .IN0(\CARRYB[697][1] ), .IN1(
        \SUMB[697][2] ), .COUT(\CARRYB[698][1] ), .SUM(\SUMB[698][1] ) );
  FADDER S3_698_2 ( .CIN(\ab[698][2] ), .IN0(\CARRYB[697][2] ), .IN1(
        \ab[697][3] ), .COUT(\CARRYB[698][2] ), .SUM(\SUMB[698][2] ) );
  FADDER S1_697_0 ( .CIN(\ab[697][0] ), .IN0(\CARRYB[696][0] ), .IN1(
        \SUMB[696][1] ), .COUT(\CARRYB[697][0] ), .SUM(PRODUCT[697]) );
  FADDER S2_697_1 ( .CIN(\ab[697][1] ), .IN0(\CARRYB[696][1] ), .IN1(
        \SUMB[696][2] ), .COUT(\CARRYB[697][1] ), .SUM(\SUMB[697][1] ) );
  FADDER S3_697_2 ( .CIN(\ab[697][2] ), .IN0(\CARRYB[696][2] ), .IN1(
        \ab[696][3] ), .COUT(\CARRYB[697][2] ), .SUM(\SUMB[697][2] ) );
  FADDER S1_696_0 ( .CIN(\ab[696][0] ), .IN0(\CARRYB[695][0] ), .IN1(
        \SUMB[695][1] ), .COUT(\CARRYB[696][0] ), .SUM(PRODUCT[696]) );
  FADDER S2_696_1 ( .CIN(\ab[696][1] ), .IN0(\CARRYB[695][1] ), .IN1(
        \SUMB[695][2] ), .COUT(\CARRYB[696][1] ), .SUM(\SUMB[696][1] ) );
  FADDER S3_696_2 ( .CIN(\ab[696][2] ), .IN0(\CARRYB[695][2] ), .IN1(
        \ab[695][3] ), .COUT(\CARRYB[696][2] ), .SUM(\SUMB[696][2] ) );
  FADDER S1_695_0 ( .CIN(\ab[695][0] ), .IN0(\CARRYB[694][0] ), .IN1(
        \SUMB[694][1] ), .COUT(\CARRYB[695][0] ), .SUM(PRODUCT[695]) );
  FADDER S2_695_1 ( .CIN(\ab[695][1] ), .IN0(\CARRYB[694][1] ), .IN1(
        \SUMB[694][2] ), .COUT(\CARRYB[695][1] ), .SUM(\SUMB[695][1] ) );
  FADDER S3_695_2 ( .CIN(\ab[695][2] ), .IN0(\CARRYB[694][2] ), .IN1(
        \ab[694][3] ), .COUT(\CARRYB[695][2] ), .SUM(\SUMB[695][2] ) );
  FADDER S1_694_0 ( .CIN(\ab[694][0] ), .IN0(\CARRYB[693][0] ), .IN1(
        \SUMB[693][1] ), .COUT(\CARRYB[694][0] ), .SUM(PRODUCT[694]) );
  FADDER S2_694_1 ( .CIN(\ab[694][1] ), .IN0(\CARRYB[693][1] ), .IN1(
        \SUMB[693][2] ), .COUT(\CARRYB[694][1] ), .SUM(\SUMB[694][1] ) );
  FADDER S3_694_2 ( .CIN(\ab[694][2] ), .IN0(\CARRYB[693][2] ), .IN1(
        \ab[693][3] ), .COUT(\CARRYB[694][2] ), .SUM(\SUMB[694][2] ) );
  FADDER S1_693_0 ( .CIN(\ab[693][0] ), .IN0(\CARRYB[692][0] ), .IN1(
        \SUMB[692][1] ), .COUT(\CARRYB[693][0] ), .SUM(PRODUCT[693]) );
  FADDER S2_693_1 ( .CIN(\ab[693][1] ), .IN0(\CARRYB[692][1] ), .IN1(
        \SUMB[692][2] ), .COUT(\CARRYB[693][1] ), .SUM(\SUMB[693][1] ) );
  FADDER S3_693_2 ( .CIN(\ab[693][2] ), .IN0(\CARRYB[692][2] ), .IN1(
        \ab[692][3] ), .COUT(\CARRYB[693][2] ), .SUM(\SUMB[693][2] ) );
  FADDER S1_692_0 ( .CIN(\ab[692][0] ), .IN0(\CARRYB[691][0] ), .IN1(
        \SUMB[691][1] ), .COUT(\CARRYB[692][0] ), .SUM(PRODUCT[692]) );
  FADDER S2_692_1 ( .CIN(\ab[692][1] ), .IN0(\CARRYB[691][1] ), .IN1(
        \SUMB[691][2] ), .COUT(\CARRYB[692][1] ), .SUM(\SUMB[692][1] ) );
  FADDER S3_692_2 ( .CIN(\ab[692][2] ), .IN0(\CARRYB[691][2] ), .IN1(
        \ab[691][3] ), .COUT(\CARRYB[692][2] ), .SUM(\SUMB[692][2] ) );
  FADDER S1_691_0 ( .CIN(\ab[691][0] ), .IN0(\CARRYB[690][0] ), .IN1(
        \SUMB[690][1] ), .COUT(\CARRYB[691][0] ), .SUM(PRODUCT[691]) );
  FADDER S2_691_1 ( .CIN(\ab[691][1] ), .IN0(\CARRYB[690][1] ), .IN1(
        \SUMB[690][2] ), .COUT(\CARRYB[691][1] ), .SUM(\SUMB[691][1] ) );
  FADDER S3_691_2 ( .CIN(\ab[691][2] ), .IN0(\CARRYB[690][2] ), .IN1(
        \ab[690][3] ), .COUT(\CARRYB[691][2] ), .SUM(\SUMB[691][2] ) );
  FADDER S1_690_0 ( .CIN(\ab[690][0] ), .IN0(\CARRYB[689][0] ), .IN1(
        \SUMB[689][1] ), .COUT(\CARRYB[690][0] ), .SUM(PRODUCT[690]) );
  FADDER S2_690_1 ( .CIN(\ab[690][1] ), .IN0(\CARRYB[689][1] ), .IN1(
        \SUMB[689][2] ), .COUT(\CARRYB[690][1] ), .SUM(\SUMB[690][1] ) );
  FADDER S3_690_2 ( .CIN(\ab[690][2] ), .IN0(\CARRYB[689][2] ), .IN1(
        \ab[689][3] ), .COUT(\CARRYB[690][2] ), .SUM(\SUMB[690][2] ) );
  FADDER S1_689_0 ( .CIN(\ab[689][0] ), .IN0(\CARRYB[688][0] ), .IN1(
        \SUMB[688][1] ), .COUT(\CARRYB[689][0] ), .SUM(PRODUCT[689]) );
  FADDER S2_689_1 ( .CIN(\ab[689][1] ), .IN0(\CARRYB[688][1] ), .IN1(
        \SUMB[688][2] ), .COUT(\CARRYB[689][1] ), .SUM(\SUMB[689][1] ) );
  FADDER S3_689_2 ( .CIN(\ab[689][2] ), .IN0(\CARRYB[688][2] ), .IN1(
        \ab[688][3] ), .COUT(\CARRYB[689][2] ), .SUM(\SUMB[689][2] ) );
  FADDER S1_688_0 ( .CIN(\ab[688][0] ), .IN0(\CARRYB[687][0] ), .IN1(
        \SUMB[687][1] ), .COUT(\CARRYB[688][0] ), .SUM(PRODUCT[688]) );
  FADDER S2_688_1 ( .CIN(\ab[688][1] ), .IN0(\CARRYB[687][1] ), .IN1(
        \SUMB[687][2] ), .COUT(\CARRYB[688][1] ), .SUM(\SUMB[688][1] ) );
  FADDER S3_688_2 ( .CIN(\ab[688][2] ), .IN0(\CARRYB[687][2] ), .IN1(
        \ab[687][3] ), .COUT(\CARRYB[688][2] ), .SUM(\SUMB[688][2] ) );
  FADDER S1_687_0 ( .CIN(\ab[687][0] ), .IN0(\CARRYB[686][0] ), .IN1(
        \SUMB[686][1] ), .COUT(\CARRYB[687][0] ), .SUM(PRODUCT[687]) );
  FADDER S2_687_1 ( .CIN(\ab[687][1] ), .IN0(\CARRYB[686][1] ), .IN1(
        \SUMB[686][2] ), .COUT(\CARRYB[687][1] ), .SUM(\SUMB[687][1] ) );
  FADDER S3_687_2 ( .CIN(\ab[687][2] ), .IN0(\CARRYB[686][2] ), .IN1(
        \ab[686][3] ), .COUT(\CARRYB[687][2] ), .SUM(\SUMB[687][2] ) );
  FADDER S1_686_0 ( .CIN(\ab[686][0] ), .IN0(\CARRYB[685][0] ), .IN1(
        \SUMB[685][1] ), .COUT(\CARRYB[686][0] ), .SUM(PRODUCT[686]) );
  FADDER S2_686_1 ( .CIN(\ab[686][1] ), .IN0(\CARRYB[685][1] ), .IN1(
        \SUMB[685][2] ), .COUT(\CARRYB[686][1] ), .SUM(\SUMB[686][1] ) );
  FADDER S3_686_2 ( .CIN(\ab[686][2] ), .IN0(\CARRYB[685][2] ), .IN1(
        \ab[685][3] ), .COUT(\CARRYB[686][2] ), .SUM(\SUMB[686][2] ) );
  FADDER S1_685_0 ( .CIN(\ab[685][0] ), .IN0(\CARRYB[684][0] ), .IN1(
        \SUMB[684][1] ), .COUT(\CARRYB[685][0] ), .SUM(PRODUCT[685]) );
  FADDER S2_685_1 ( .CIN(\ab[685][1] ), .IN0(\CARRYB[684][1] ), .IN1(
        \SUMB[684][2] ), .COUT(\CARRYB[685][1] ), .SUM(\SUMB[685][1] ) );
  FADDER S3_685_2 ( .CIN(\ab[685][2] ), .IN0(\CARRYB[684][2] ), .IN1(
        \ab[684][3] ), .COUT(\CARRYB[685][2] ), .SUM(\SUMB[685][2] ) );
  FADDER S1_684_0 ( .CIN(\ab[684][0] ), .IN0(\CARRYB[683][0] ), .IN1(
        \SUMB[683][1] ), .COUT(\CARRYB[684][0] ), .SUM(PRODUCT[684]) );
  FADDER S2_684_1 ( .CIN(\ab[684][1] ), .IN0(\CARRYB[683][1] ), .IN1(
        \SUMB[683][2] ), .COUT(\CARRYB[684][1] ), .SUM(\SUMB[684][1] ) );
  FADDER S3_684_2 ( .CIN(\ab[684][2] ), .IN0(\CARRYB[683][2] ), .IN1(
        \ab[683][3] ), .COUT(\CARRYB[684][2] ), .SUM(\SUMB[684][2] ) );
  FADDER S1_683_0 ( .CIN(\ab[683][0] ), .IN0(\CARRYB[682][0] ), .IN1(
        \SUMB[682][1] ), .COUT(\CARRYB[683][0] ), .SUM(PRODUCT[683]) );
  FADDER S2_683_1 ( .CIN(\ab[683][1] ), .IN0(\CARRYB[682][1] ), .IN1(
        \SUMB[682][2] ), .COUT(\CARRYB[683][1] ), .SUM(\SUMB[683][1] ) );
  FADDER S3_683_2 ( .CIN(\ab[683][2] ), .IN0(\CARRYB[682][2] ), .IN1(
        \ab[682][3] ), .COUT(\CARRYB[683][2] ), .SUM(\SUMB[683][2] ) );
  FADDER S1_682_0 ( .CIN(\ab[682][0] ), .IN0(\CARRYB[681][0] ), .IN1(
        \SUMB[681][1] ), .COUT(\CARRYB[682][0] ), .SUM(PRODUCT[682]) );
  FADDER S2_682_1 ( .CIN(\ab[682][1] ), .IN0(\CARRYB[681][1] ), .IN1(
        \SUMB[681][2] ), .COUT(\CARRYB[682][1] ), .SUM(\SUMB[682][1] ) );
  FADDER S3_682_2 ( .CIN(\ab[682][2] ), .IN0(\CARRYB[681][2] ), .IN1(
        \ab[681][3] ), .COUT(\CARRYB[682][2] ), .SUM(\SUMB[682][2] ) );
  FADDER S1_681_0 ( .CIN(\ab[681][0] ), .IN0(\CARRYB[680][0] ), .IN1(
        \SUMB[680][1] ), .COUT(\CARRYB[681][0] ), .SUM(PRODUCT[681]) );
  FADDER S2_681_1 ( .CIN(\ab[681][1] ), .IN0(\CARRYB[680][1] ), .IN1(
        \SUMB[680][2] ), .COUT(\CARRYB[681][1] ), .SUM(\SUMB[681][1] ) );
  FADDER S3_681_2 ( .CIN(\ab[681][2] ), .IN0(\CARRYB[680][2] ), .IN1(
        \ab[680][3] ), .COUT(\CARRYB[681][2] ), .SUM(\SUMB[681][2] ) );
  FADDER S1_680_0 ( .CIN(\ab[680][0] ), .IN0(\CARRYB[679][0] ), .IN1(
        \SUMB[679][1] ), .COUT(\CARRYB[680][0] ), .SUM(PRODUCT[680]) );
  FADDER S2_680_1 ( .CIN(\ab[680][1] ), .IN0(\CARRYB[679][1] ), .IN1(
        \SUMB[679][2] ), .COUT(\CARRYB[680][1] ), .SUM(\SUMB[680][1] ) );
  FADDER S3_680_2 ( .CIN(\ab[680][2] ), .IN0(\CARRYB[679][2] ), .IN1(
        \ab[679][3] ), .COUT(\CARRYB[680][2] ), .SUM(\SUMB[680][2] ) );
  FADDER S1_679_0 ( .CIN(\ab[679][0] ), .IN0(\CARRYB[678][0] ), .IN1(
        \SUMB[678][1] ), .COUT(\CARRYB[679][0] ), .SUM(PRODUCT[679]) );
  FADDER S2_679_1 ( .CIN(\ab[679][1] ), .IN0(\CARRYB[678][1] ), .IN1(
        \SUMB[678][2] ), .COUT(\CARRYB[679][1] ), .SUM(\SUMB[679][1] ) );
  FADDER S3_679_2 ( .CIN(\ab[679][2] ), .IN0(\CARRYB[678][2] ), .IN1(
        \ab[678][3] ), .COUT(\CARRYB[679][2] ), .SUM(\SUMB[679][2] ) );
  FADDER S1_678_0 ( .CIN(\ab[678][0] ), .IN0(\CARRYB[677][0] ), .IN1(
        \SUMB[677][1] ), .COUT(\CARRYB[678][0] ), .SUM(PRODUCT[678]) );
  FADDER S2_678_1 ( .CIN(\ab[678][1] ), .IN0(\CARRYB[677][1] ), .IN1(
        \SUMB[677][2] ), .COUT(\CARRYB[678][1] ), .SUM(\SUMB[678][1] ) );
  FADDER S3_678_2 ( .CIN(\ab[678][2] ), .IN0(\CARRYB[677][2] ), .IN1(
        \ab[677][3] ), .COUT(\CARRYB[678][2] ), .SUM(\SUMB[678][2] ) );
  FADDER S1_677_0 ( .CIN(\ab[677][0] ), .IN0(\CARRYB[676][0] ), .IN1(
        \SUMB[676][1] ), .COUT(\CARRYB[677][0] ), .SUM(PRODUCT[677]) );
  FADDER S2_677_1 ( .CIN(\ab[677][1] ), .IN0(\CARRYB[676][1] ), .IN1(
        \SUMB[676][2] ), .COUT(\CARRYB[677][1] ), .SUM(\SUMB[677][1] ) );
  FADDER S3_677_2 ( .CIN(\ab[677][2] ), .IN0(\CARRYB[676][2] ), .IN1(
        \ab[676][3] ), .COUT(\CARRYB[677][2] ), .SUM(\SUMB[677][2] ) );
  FADDER S1_676_0 ( .CIN(\ab[676][0] ), .IN0(\CARRYB[675][0] ), .IN1(
        \SUMB[675][1] ), .COUT(\CARRYB[676][0] ), .SUM(PRODUCT[676]) );
  FADDER S2_676_1 ( .CIN(\ab[676][1] ), .IN0(\CARRYB[675][1] ), .IN1(
        \SUMB[675][2] ), .COUT(\CARRYB[676][1] ), .SUM(\SUMB[676][1] ) );
  FADDER S3_676_2 ( .CIN(\ab[676][2] ), .IN0(\CARRYB[675][2] ), .IN1(
        \ab[675][3] ), .COUT(\CARRYB[676][2] ), .SUM(\SUMB[676][2] ) );
  FADDER S1_675_0 ( .CIN(\ab[675][0] ), .IN0(\CARRYB[674][0] ), .IN1(
        \SUMB[674][1] ), .COUT(\CARRYB[675][0] ), .SUM(PRODUCT[675]) );
  FADDER S2_675_1 ( .CIN(\ab[675][1] ), .IN0(\CARRYB[674][1] ), .IN1(
        \SUMB[674][2] ), .COUT(\CARRYB[675][1] ), .SUM(\SUMB[675][1] ) );
  FADDER S3_675_2 ( .CIN(\ab[675][2] ), .IN0(\CARRYB[674][2] ), .IN1(
        \ab[674][3] ), .COUT(\CARRYB[675][2] ), .SUM(\SUMB[675][2] ) );
  FADDER S1_674_0 ( .CIN(\ab[674][0] ), .IN0(\CARRYB[673][0] ), .IN1(
        \SUMB[673][1] ), .COUT(\CARRYB[674][0] ), .SUM(PRODUCT[674]) );
  FADDER S2_674_1 ( .CIN(\ab[674][1] ), .IN0(\CARRYB[673][1] ), .IN1(
        \SUMB[673][2] ), .COUT(\CARRYB[674][1] ), .SUM(\SUMB[674][1] ) );
  FADDER S3_674_2 ( .CIN(\ab[674][2] ), .IN0(\CARRYB[673][2] ), .IN1(
        \ab[673][3] ), .COUT(\CARRYB[674][2] ), .SUM(\SUMB[674][2] ) );
  FADDER S1_673_0 ( .CIN(\ab[673][0] ), .IN0(\CARRYB[672][0] ), .IN1(
        \SUMB[672][1] ), .COUT(\CARRYB[673][0] ), .SUM(PRODUCT[673]) );
  FADDER S2_673_1 ( .CIN(\ab[673][1] ), .IN0(\CARRYB[672][1] ), .IN1(
        \SUMB[672][2] ), .COUT(\CARRYB[673][1] ), .SUM(\SUMB[673][1] ) );
  FADDER S3_673_2 ( .CIN(\ab[673][2] ), .IN0(\CARRYB[672][2] ), .IN1(
        \ab[672][3] ), .COUT(\CARRYB[673][2] ), .SUM(\SUMB[673][2] ) );
  FADDER S1_672_0 ( .CIN(\ab[672][0] ), .IN0(\CARRYB[671][0] ), .IN1(
        \SUMB[671][1] ), .COUT(\CARRYB[672][0] ), .SUM(PRODUCT[672]) );
  FADDER S2_672_1 ( .CIN(\ab[672][1] ), .IN0(\CARRYB[671][1] ), .IN1(
        \SUMB[671][2] ), .COUT(\CARRYB[672][1] ), .SUM(\SUMB[672][1] ) );
  FADDER S3_672_2 ( .CIN(\ab[672][2] ), .IN0(\CARRYB[671][2] ), .IN1(
        \ab[671][3] ), .COUT(\CARRYB[672][2] ), .SUM(\SUMB[672][2] ) );
  FADDER S1_671_0 ( .CIN(\ab[671][0] ), .IN0(\CARRYB[670][0] ), .IN1(
        \SUMB[670][1] ), .COUT(\CARRYB[671][0] ), .SUM(PRODUCT[671]) );
  FADDER S2_671_1 ( .CIN(\ab[671][1] ), .IN0(\CARRYB[670][1] ), .IN1(
        \SUMB[670][2] ), .COUT(\CARRYB[671][1] ), .SUM(\SUMB[671][1] ) );
  FADDER S3_671_2 ( .CIN(\ab[671][2] ), .IN0(\CARRYB[670][2] ), .IN1(
        \ab[670][3] ), .COUT(\CARRYB[671][2] ), .SUM(\SUMB[671][2] ) );
  FADDER S1_670_0 ( .CIN(\ab[670][0] ), .IN0(\CARRYB[669][0] ), .IN1(
        \SUMB[669][1] ), .COUT(\CARRYB[670][0] ), .SUM(PRODUCT[670]) );
  FADDER S2_670_1 ( .CIN(\ab[670][1] ), .IN0(\CARRYB[669][1] ), .IN1(
        \SUMB[669][2] ), .COUT(\CARRYB[670][1] ), .SUM(\SUMB[670][1] ) );
  FADDER S3_670_2 ( .CIN(\ab[670][2] ), .IN0(\CARRYB[669][2] ), .IN1(
        \ab[669][3] ), .COUT(\CARRYB[670][2] ), .SUM(\SUMB[670][2] ) );
  FADDER S1_669_0 ( .CIN(\ab[669][0] ), .IN0(\CARRYB[668][0] ), .IN1(
        \SUMB[668][1] ), .COUT(\CARRYB[669][0] ), .SUM(PRODUCT[669]) );
  FADDER S2_669_1 ( .CIN(\ab[669][1] ), .IN0(\CARRYB[668][1] ), .IN1(
        \SUMB[668][2] ), .COUT(\CARRYB[669][1] ), .SUM(\SUMB[669][1] ) );
  FADDER S3_669_2 ( .CIN(\ab[669][2] ), .IN0(\CARRYB[668][2] ), .IN1(
        \ab[668][3] ), .COUT(\CARRYB[669][2] ), .SUM(\SUMB[669][2] ) );
  FADDER S1_668_0 ( .CIN(\ab[668][0] ), .IN0(\CARRYB[667][0] ), .IN1(
        \SUMB[667][1] ), .COUT(\CARRYB[668][0] ), .SUM(PRODUCT[668]) );
  FADDER S2_668_1 ( .CIN(\ab[668][1] ), .IN0(\CARRYB[667][1] ), .IN1(
        \SUMB[667][2] ), .COUT(\CARRYB[668][1] ), .SUM(\SUMB[668][1] ) );
  FADDER S3_668_2 ( .CIN(\ab[668][2] ), .IN0(\CARRYB[667][2] ), .IN1(
        \ab[667][3] ), .COUT(\CARRYB[668][2] ), .SUM(\SUMB[668][2] ) );
  FADDER S1_667_0 ( .CIN(\ab[667][0] ), .IN0(\CARRYB[666][0] ), .IN1(
        \SUMB[666][1] ), .COUT(\CARRYB[667][0] ), .SUM(PRODUCT[667]) );
  FADDER S2_667_1 ( .CIN(\ab[667][1] ), .IN0(\CARRYB[666][1] ), .IN1(
        \SUMB[666][2] ), .COUT(\CARRYB[667][1] ), .SUM(\SUMB[667][1] ) );
  FADDER S3_667_2 ( .CIN(\ab[667][2] ), .IN0(\CARRYB[666][2] ), .IN1(
        \ab[666][3] ), .COUT(\CARRYB[667][2] ), .SUM(\SUMB[667][2] ) );
  FADDER S1_666_0 ( .CIN(\ab[666][0] ), .IN0(\CARRYB[665][0] ), .IN1(
        \SUMB[665][1] ), .COUT(\CARRYB[666][0] ), .SUM(PRODUCT[666]) );
  FADDER S2_666_1 ( .CIN(\ab[666][1] ), .IN0(\CARRYB[665][1] ), .IN1(
        \SUMB[665][2] ), .COUT(\CARRYB[666][1] ), .SUM(\SUMB[666][1] ) );
  FADDER S3_666_2 ( .CIN(\ab[666][2] ), .IN0(\CARRYB[665][2] ), .IN1(
        \ab[665][3] ), .COUT(\CARRYB[666][2] ), .SUM(\SUMB[666][2] ) );
  FADDER S1_665_0 ( .CIN(\ab[665][0] ), .IN0(\CARRYB[664][0] ), .IN1(
        \SUMB[664][1] ), .COUT(\CARRYB[665][0] ), .SUM(PRODUCT[665]) );
  FADDER S2_665_1 ( .CIN(\ab[665][1] ), .IN0(\CARRYB[664][1] ), .IN1(
        \SUMB[664][2] ), .COUT(\CARRYB[665][1] ), .SUM(\SUMB[665][1] ) );
  FADDER S3_665_2 ( .CIN(\ab[665][2] ), .IN0(\CARRYB[664][2] ), .IN1(
        \ab[664][3] ), .COUT(\CARRYB[665][2] ), .SUM(\SUMB[665][2] ) );
  FADDER S1_664_0 ( .CIN(\ab[664][0] ), .IN0(\CARRYB[663][0] ), .IN1(
        \SUMB[663][1] ), .COUT(\CARRYB[664][0] ), .SUM(PRODUCT[664]) );
  FADDER S2_664_1 ( .CIN(\ab[664][1] ), .IN0(\CARRYB[663][1] ), .IN1(
        \SUMB[663][2] ), .COUT(\CARRYB[664][1] ), .SUM(\SUMB[664][1] ) );
  FADDER S3_664_2 ( .CIN(\ab[664][2] ), .IN0(\CARRYB[663][2] ), .IN1(
        \ab[663][3] ), .COUT(\CARRYB[664][2] ), .SUM(\SUMB[664][2] ) );
  FADDER S1_663_0 ( .CIN(\ab[663][0] ), .IN0(\CARRYB[662][0] ), .IN1(
        \SUMB[662][1] ), .COUT(\CARRYB[663][0] ), .SUM(PRODUCT[663]) );
  FADDER S2_663_1 ( .CIN(\ab[663][1] ), .IN0(\CARRYB[662][1] ), .IN1(
        \SUMB[662][2] ), .COUT(\CARRYB[663][1] ), .SUM(\SUMB[663][1] ) );
  FADDER S3_663_2 ( .CIN(\ab[663][2] ), .IN0(\CARRYB[662][2] ), .IN1(
        \ab[662][3] ), .COUT(\CARRYB[663][2] ), .SUM(\SUMB[663][2] ) );
  FADDER S1_662_0 ( .CIN(\ab[662][0] ), .IN0(\CARRYB[661][0] ), .IN1(
        \SUMB[661][1] ), .COUT(\CARRYB[662][0] ), .SUM(PRODUCT[662]) );
  FADDER S2_662_1 ( .CIN(\ab[662][1] ), .IN0(\CARRYB[661][1] ), .IN1(
        \SUMB[661][2] ), .COUT(\CARRYB[662][1] ), .SUM(\SUMB[662][1] ) );
  FADDER S3_662_2 ( .CIN(\ab[662][2] ), .IN0(\CARRYB[661][2] ), .IN1(
        \ab[661][3] ), .COUT(\CARRYB[662][2] ), .SUM(\SUMB[662][2] ) );
  FADDER S1_661_0 ( .CIN(\ab[661][0] ), .IN0(\CARRYB[660][0] ), .IN1(
        \SUMB[660][1] ), .COUT(\CARRYB[661][0] ), .SUM(PRODUCT[661]) );
  FADDER S2_661_1 ( .CIN(\ab[661][1] ), .IN0(\CARRYB[660][1] ), .IN1(
        \SUMB[660][2] ), .COUT(\CARRYB[661][1] ), .SUM(\SUMB[661][1] ) );
  FADDER S3_661_2 ( .CIN(\ab[661][2] ), .IN0(\CARRYB[660][2] ), .IN1(
        \ab[660][3] ), .COUT(\CARRYB[661][2] ), .SUM(\SUMB[661][2] ) );
  FADDER S1_660_0 ( .CIN(\ab[660][0] ), .IN0(\CARRYB[659][0] ), .IN1(
        \SUMB[659][1] ), .COUT(\CARRYB[660][0] ), .SUM(PRODUCT[660]) );
  FADDER S2_660_1 ( .CIN(\ab[660][1] ), .IN0(\CARRYB[659][1] ), .IN1(
        \SUMB[659][2] ), .COUT(\CARRYB[660][1] ), .SUM(\SUMB[660][1] ) );
  FADDER S3_660_2 ( .CIN(\ab[660][2] ), .IN0(\CARRYB[659][2] ), .IN1(
        \ab[659][3] ), .COUT(\CARRYB[660][2] ), .SUM(\SUMB[660][2] ) );
  FADDER S1_659_0 ( .CIN(\ab[659][0] ), .IN0(\CARRYB[658][0] ), .IN1(
        \SUMB[658][1] ), .COUT(\CARRYB[659][0] ), .SUM(PRODUCT[659]) );
  FADDER S2_659_1 ( .CIN(\ab[659][1] ), .IN0(\CARRYB[658][1] ), .IN1(
        \SUMB[658][2] ), .COUT(\CARRYB[659][1] ), .SUM(\SUMB[659][1] ) );
  FADDER S3_659_2 ( .CIN(\ab[659][2] ), .IN0(\CARRYB[658][2] ), .IN1(
        \ab[658][3] ), .COUT(\CARRYB[659][2] ), .SUM(\SUMB[659][2] ) );
  FADDER S1_658_0 ( .CIN(\ab[658][0] ), .IN0(\CARRYB[657][0] ), .IN1(
        \SUMB[657][1] ), .COUT(\CARRYB[658][0] ), .SUM(PRODUCT[658]) );
  FADDER S2_658_1 ( .CIN(\ab[658][1] ), .IN0(\CARRYB[657][1] ), .IN1(
        \SUMB[657][2] ), .COUT(\CARRYB[658][1] ), .SUM(\SUMB[658][1] ) );
  FADDER S3_658_2 ( .CIN(\ab[658][2] ), .IN0(\CARRYB[657][2] ), .IN1(
        \ab[657][3] ), .COUT(\CARRYB[658][2] ), .SUM(\SUMB[658][2] ) );
  FADDER S1_657_0 ( .CIN(\ab[657][0] ), .IN0(\CARRYB[656][0] ), .IN1(
        \SUMB[656][1] ), .COUT(\CARRYB[657][0] ), .SUM(PRODUCT[657]) );
  FADDER S2_657_1 ( .CIN(\ab[657][1] ), .IN0(\CARRYB[656][1] ), .IN1(
        \SUMB[656][2] ), .COUT(\CARRYB[657][1] ), .SUM(\SUMB[657][1] ) );
  FADDER S3_657_2 ( .CIN(\ab[657][2] ), .IN0(\CARRYB[656][2] ), .IN1(
        \ab[656][3] ), .COUT(\CARRYB[657][2] ), .SUM(\SUMB[657][2] ) );
  FADDER S1_656_0 ( .CIN(\ab[656][0] ), .IN0(\CARRYB[655][0] ), .IN1(
        \SUMB[655][1] ), .COUT(\CARRYB[656][0] ), .SUM(PRODUCT[656]) );
  FADDER S2_656_1 ( .CIN(\ab[656][1] ), .IN0(\CARRYB[655][1] ), .IN1(
        \SUMB[655][2] ), .COUT(\CARRYB[656][1] ), .SUM(\SUMB[656][1] ) );
  FADDER S3_656_2 ( .CIN(\ab[656][2] ), .IN0(\CARRYB[655][2] ), .IN1(
        \ab[655][3] ), .COUT(\CARRYB[656][2] ), .SUM(\SUMB[656][2] ) );
  FADDER S1_655_0 ( .CIN(\ab[655][0] ), .IN0(\CARRYB[654][0] ), .IN1(
        \SUMB[654][1] ), .COUT(\CARRYB[655][0] ), .SUM(PRODUCT[655]) );
  FADDER S2_655_1 ( .CIN(\ab[655][1] ), .IN0(\CARRYB[654][1] ), .IN1(
        \SUMB[654][2] ), .COUT(\CARRYB[655][1] ), .SUM(\SUMB[655][1] ) );
  FADDER S3_655_2 ( .CIN(\ab[655][2] ), .IN0(\CARRYB[654][2] ), .IN1(
        \ab[654][3] ), .COUT(\CARRYB[655][2] ), .SUM(\SUMB[655][2] ) );
  FADDER S1_654_0 ( .CIN(\ab[654][0] ), .IN0(\CARRYB[653][0] ), .IN1(
        \SUMB[653][1] ), .COUT(\CARRYB[654][0] ), .SUM(PRODUCT[654]) );
  FADDER S2_654_1 ( .CIN(\ab[654][1] ), .IN0(\CARRYB[653][1] ), .IN1(
        \SUMB[653][2] ), .COUT(\CARRYB[654][1] ), .SUM(\SUMB[654][1] ) );
  FADDER S3_654_2 ( .CIN(\ab[654][2] ), .IN0(\CARRYB[653][2] ), .IN1(
        \ab[653][3] ), .COUT(\CARRYB[654][2] ), .SUM(\SUMB[654][2] ) );
  FADDER S1_653_0 ( .CIN(\ab[653][0] ), .IN0(\CARRYB[652][0] ), .IN1(
        \SUMB[652][1] ), .COUT(\CARRYB[653][0] ), .SUM(PRODUCT[653]) );
  FADDER S2_653_1 ( .CIN(\ab[653][1] ), .IN0(\CARRYB[652][1] ), .IN1(
        \SUMB[652][2] ), .COUT(\CARRYB[653][1] ), .SUM(\SUMB[653][1] ) );
  FADDER S3_653_2 ( .CIN(\ab[653][2] ), .IN0(\CARRYB[652][2] ), .IN1(
        \ab[652][3] ), .COUT(\CARRYB[653][2] ), .SUM(\SUMB[653][2] ) );
  FADDER S1_652_0 ( .CIN(\ab[652][0] ), .IN0(\CARRYB[651][0] ), .IN1(
        \SUMB[651][1] ), .COUT(\CARRYB[652][0] ), .SUM(PRODUCT[652]) );
  FADDER S2_652_1 ( .CIN(\ab[652][1] ), .IN0(\CARRYB[651][1] ), .IN1(
        \SUMB[651][2] ), .COUT(\CARRYB[652][1] ), .SUM(\SUMB[652][1] ) );
  FADDER S3_652_2 ( .CIN(\ab[652][2] ), .IN0(\CARRYB[651][2] ), .IN1(
        \ab[651][3] ), .COUT(\CARRYB[652][2] ), .SUM(\SUMB[652][2] ) );
  FADDER S1_651_0 ( .CIN(\ab[651][0] ), .IN0(\CARRYB[650][0] ), .IN1(
        \SUMB[650][1] ), .COUT(\CARRYB[651][0] ), .SUM(PRODUCT[651]) );
  FADDER S2_651_1 ( .CIN(\ab[651][1] ), .IN0(\CARRYB[650][1] ), .IN1(
        \SUMB[650][2] ), .COUT(\CARRYB[651][1] ), .SUM(\SUMB[651][1] ) );
  FADDER S3_651_2 ( .CIN(\ab[651][2] ), .IN0(\CARRYB[650][2] ), .IN1(
        \ab[650][3] ), .COUT(\CARRYB[651][2] ), .SUM(\SUMB[651][2] ) );
  FADDER S1_650_0 ( .CIN(\ab[650][0] ), .IN0(\CARRYB[649][0] ), .IN1(
        \SUMB[649][1] ), .COUT(\CARRYB[650][0] ), .SUM(PRODUCT[650]) );
  FADDER S2_650_1 ( .CIN(\ab[650][1] ), .IN0(\CARRYB[649][1] ), .IN1(
        \SUMB[649][2] ), .COUT(\CARRYB[650][1] ), .SUM(\SUMB[650][1] ) );
  FADDER S3_650_2 ( .CIN(\ab[650][2] ), .IN0(\CARRYB[649][2] ), .IN1(
        \ab[649][3] ), .COUT(\CARRYB[650][2] ), .SUM(\SUMB[650][2] ) );
  FADDER S1_649_0 ( .CIN(\ab[649][0] ), .IN0(\CARRYB[648][0] ), .IN1(
        \SUMB[648][1] ), .COUT(\CARRYB[649][0] ), .SUM(PRODUCT[649]) );
  FADDER S2_649_1 ( .CIN(\ab[649][1] ), .IN0(\CARRYB[648][1] ), .IN1(
        \SUMB[648][2] ), .COUT(\CARRYB[649][1] ), .SUM(\SUMB[649][1] ) );
  FADDER S3_649_2 ( .CIN(\ab[649][2] ), .IN0(\CARRYB[648][2] ), .IN1(
        \ab[648][3] ), .COUT(\CARRYB[649][2] ), .SUM(\SUMB[649][2] ) );
  FADDER S1_648_0 ( .CIN(\ab[648][0] ), .IN0(\CARRYB[647][0] ), .IN1(
        \SUMB[647][1] ), .COUT(\CARRYB[648][0] ), .SUM(PRODUCT[648]) );
  FADDER S2_648_1 ( .CIN(\ab[648][1] ), .IN0(\CARRYB[647][1] ), .IN1(
        \SUMB[647][2] ), .COUT(\CARRYB[648][1] ), .SUM(\SUMB[648][1] ) );
  FADDER S3_648_2 ( .CIN(\ab[648][2] ), .IN0(\CARRYB[647][2] ), .IN1(
        \ab[647][3] ), .COUT(\CARRYB[648][2] ), .SUM(\SUMB[648][2] ) );
  FADDER S1_647_0 ( .CIN(\ab[647][0] ), .IN0(\CARRYB[646][0] ), .IN1(
        \SUMB[646][1] ), .COUT(\CARRYB[647][0] ), .SUM(PRODUCT[647]) );
  FADDER S2_647_1 ( .CIN(\ab[647][1] ), .IN0(\CARRYB[646][1] ), .IN1(
        \SUMB[646][2] ), .COUT(\CARRYB[647][1] ), .SUM(\SUMB[647][1] ) );
  FADDER S3_647_2 ( .CIN(\ab[647][2] ), .IN0(\CARRYB[646][2] ), .IN1(
        \ab[646][3] ), .COUT(\CARRYB[647][2] ), .SUM(\SUMB[647][2] ) );
  FADDER S1_646_0 ( .CIN(\ab[646][0] ), .IN0(\CARRYB[645][0] ), .IN1(
        \SUMB[645][1] ), .COUT(\CARRYB[646][0] ), .SUM(PRODUCT[646]) );
  FADDER S2_646_1 ( .CIN(\ab[646][1] ), .IN0(\CARRYB[645][1] ), .IN1(
        \SUMB[645][2] ), .COUT(\CARRYB[646][1] ), .SUM(\SUMB[646][1] ) );
  FADDER S3_646_2 ( .CIN(\ab[646][2] ), .IN0(\CARRYB[645][2] ), .IN1(
        \ab[645][3] ), .COUT(\CARRYB[646][2] ), .SUM(\SUMB[646][2] ) );
  FADDER S1_645_0 ( .CIN(\ab[645][0] ), .IN0(\CARRYB[644][0] ), .IN1(
        \SUMB[644][1] ), .COUT(\CARRYB[645][0] ), .SUM(PRODUCT[645]) );
  FADDER S2_645_1 ( .CIN(\ab[645][1] ), .IN0(\CARRYB[644][1] ), .IN1(
        \SUMB[644][2] ), .COUT(\CARRYB[645][1] ), .SUM(\SUMB[645][1] ) );
  FADDER S3_645_2 ( .CIN(\ab[645][2] ), .IN0(\CARRYB[644][2] ), .IN1(
        \ab[644][3] ), .COUT(\CARRYB[645][2] ), .SUM(\SUMB[645][2] ) );
  FADDER S1_644_0 ( .CIN(\ab[644][0] ), .IN0(\CARRYB[643][0] ), .IN1(
        \SUMB[643][1] ), .COUT(\CARRYB[644][0] ), .SUM(PRODUCT[644]) );
  FADDER S2_644_1 ( .CIN(\ab[644][1] ), .IN0(\CARRYB[643][1] ), .IN1(
        \SUMB[643][2] ), .COUT(\CARRYB[644][1] ), .SUM(\SUMB[644][1] ) );
  FADDER S3_644_2 ( .CIN(\ab[644][2] ), .IN0(\CARRYB[643][2] ), .IN1(
        \ab[643][3] ), .COUT(\CARRYB[644][2] ), .SUM(\SUMB[644][2] ) );
  FADDER S1_643_0 ( .CIN(\ab[643][0] ), .IN0(\CARRYB[642][0] ), .IN1(
        \SUMB[642][1] ), .COUT(\CARRYB[643][0] ), .SUM(PRODUCT[643]) );
  FADDER S2_643_1 ( .CIN(\ab[643][1] ), .IN0(\CARRYB[642][1] ), .IN1(
        \SUMB[642][2] ), .COUT(\CARRYB[643][1] ), .SUM(\SUMB[643][1] ) );
  FADDER S3_643_2 ( .CIN(\ab[643][2] ), .IN0(\CARRYB[642][2] ), .IN1(
        \ab[642][3] ), .COUT(\CARRYB[643][2] ), .SUM(\SUMB[643][2] ) );
  FADDER S1_642_0 ( .CIN(\ab[642][0] ), .IN0(\CARRYB[641][0] ), .IN1(
        \SUMB[641][1] ), .COUT(\CARRYB[642][0] ), .SUM(PRODUCT[642]) );
  FADDER S2_642_1 ( .CIN(\ab[642][1] ), .IN0(\CARRYB[641][1] ), .IN1(
        \SUMB[641][2] ), .COUT(\CARRYB[642][1] ), .SUM(\SUMB[642][1] ) );
  FADDER S3_642_2 ( .CIN(\ab[642][2] ), .IN0(\CARRYB[641][2] ), .IN1(
        \ab[641][3] ), .COUT(\CARRYB[642][2] ), .SUM(\SUMB[642][2] ) );
  FADDER S1_641_0 ( .CIN(\ab[641][0] ), .IN0(\CARRYB[640][0] ), .IN1(
        \SUMB[640][1] ), .COUT(\CARRYB[641][0] ), .SUM(PRODUCT[641]) );
  FADDER S2_641_1 ( .CIN(\ab[641][1] ), .IN0(\CARRYB[640][1] ), .IN1(
        \SUMB[640][2] ), .COUT(\CARRYB[641][1] ), .SUM(\SUMB[641][1] ) );
  FADDER S3_641_2 ( .CIN(\ab[641][2] ), .IN0(\CARRYB[640][2] ), .IN1(
        \ab[640][3] ), .COUT(\CARRYB[641][2] ), .SUM(\SUMB[641][2] ) );
  FADDER S1_640_0 ( .CIN(\ab[640][0] ), .IN0(\CARRYB[639][0] ), .IN1(
        \SUMB[639][1] ), .COUT(\CARRYB[640][0] ), .SUM(PRODUCT[640]) );
  FADDER S2_640_1 ( .CIN(\ab[640][1] ), .IN0(\CARRYB[639][1] ), .IN1(
        \SUMB[639][2] ), .COUT(\CARRYB[640][1] ), .SUM(\SUMB[640][1] ) );
  FADDER S3_640_2 ( .CIN(\ab[640][2] ), .IN0(\CARRYB[639][2] ), .IN1(
        \ab[639][3] ), .COUT(\CARRYB[640][2] ), .SUM(\SUMB[640][2] ) );
  FADDER S1_639_0 ( .CIN(\ab[639][0] ), .IN0(\CARRYB[638][0] ), .IN1(
        \SUMB[638][1] ), .COUT(\CARRYB[639][0] ), .SUM(PRODUCT[639]) );
  FADDER S2_639_1 ( .CIN(\ab[639][1] ), .IN0(\CARRYB[638][1] ), .IN1(
        \SUMB[638][2] ), .COUT(\CARRYB[639][1] ), .SUM(\SUMB[639][1] ) );
  FADDER S3_639_2 ( .CIN(\ab[639][2] ), .IN0(\CARRYB[638][2] ), .IN1(
        \ab[638][3] ), .COUT(\CARRYB[639][2] ), .SUM(\SUMB[639][2] ) );
  FADDER S1_638_0 ( .CIN(\ab[638][0] ), .IN0(\CARRYB[637][0] ), .IN1(
        \SUMB[637][1] ), .COUT(\CARRYB[638][0] ), .SUM(PRODUCT[638]) );
  FADDER S2_638_1 ( .CIN(\ab[638][1] ), .IN0(\CARRYB[637][1] ), .IN1(
        \SUMB[637][2] ), .COUT(\CARRYB[638][1] ), .SUM(\SUMB[638][1] ) );
  FADDER S3_638_2 ( .CIN(\ab[638][2] ), .IN0(\CARRYB[637][2] ), .IN1(
        \ab[637][3] ), .COUT(\CARRYB[638][2] ), .SUM(\SUMB[638][2] ) );
  FADDER S1_637_0 ( .CIN(\ab[637][0] ), .IN0(\CARRYB[636][0] ), .IN1(
        \SUMB[636][1] ), .COUT(\CARRYB[637][0] ), .SUM(PRODUCT[637]) );
  FADDER S2_637_1 ( .CIN(\ab[637][1] ), .IN0(\CARRYB[636][1] ), .IN1(
        \SUMB[636][2] ), .COUT(\CARRYB[637][1] ), .SUM(\SUMB[637][1] ) );
  FADDER S3_637_2 ( .CIN(\ab[637][2] ), .IN0(\CARRYB[636][2] ), .IN1(
        \ab[636][3] ), .COUT(\CARRYB[637][2] ), .SUM(\SUMB[637][2] ) );
  FADDER S1_636_0 ( .CIN(\ab[636][0] ), .IN0(\CARRYB[635][0] ), .IN1(
        \SUMB[635][1] ), .COUT(\CARRYB[636][0] ), .SUM(PRODUCT[636]) );
  FADDER S2_636_1 ( .CIN(\ab[636][1] ), .IN0(\CARRYB[635][1] ), .IN1(
        \SUMB[635][2] ), .COUT(\CARRYB[636][1] ), .SUM(\SUMB[636][1] ) );
  FADDER S3_636_2 ( .CIN(\ab[636][2] ), .IN0(\CARRYB[635][2] ), .IN1(
        \ab[635][3] ), .COUT(\CARRYB[636][2] ), .SUM(\SUMB[636][2] ) );
  FADDER S1_635_0 ( .CIN(\ab[635][0] ), .IN0(\CARRYB[634][0] ), .IN1(
        \SUMB[634][1] ), .COUT(\CARRYB[635][0] ), .SUM(PRODUCT[635]) );
  FADDER S2_635_1 ( .CIN(\ab[635][1] ), .IN0(\CARRYB[634][1] ), .IN1(
        \SUMB[634][2] ), .COUT(\CARRYB[635][1] ), .SUM(\SUMB[635][1] ) );
  FADDER S3_635_2 ( .CIN(\ab[635][2] ), .IN0(\CARRYB[634][2] ), .IN1(
        \ab[634][3] ), .COUT(\CARRYB[635][2] ), .SUM(\SUMB[635][2] ) );
  FADDER S1_634_0 ( .CIN(\ab[634][0] ), .IN0(\CARRYB[633][0] ), .IN1(
        \SUMB[633][1] ), .COUT(\CARRYB[634][0] ), .SUM(PRODUCT[634]) );
  FADDER S2_634_1 ( .CIN(\ab[634][1] ), .IN0(\CARRYB[633][1] ), .IN1(
        \SUMB[633][2] ), .COUT(\CARRYB[634][1] ), .SUM(\SUMB[634][1] ) );
  FADDER S3_634_2 ( .CIN(\ab[634][2] ), .IN0(\CARRYB[633][2] ), .IN1(
        \ab[633][3] ), .COUT(\CARRYB[634][2] ), .SUM(\SUMB[634][2] ) );
  FADDER S1_633_0 ( .CIN(\ab[633][0] ), .IN0(\CARRYB[632][0] ), .IN1(
        \SUMB[632][1] ), .COUT(\CARRYB[633][0] ), .SUM(PRODUCT[633]) );
  FADDER S2_633_1 ( .CIN(\ab[633][1] ), .IN0(\CARRYB[632][1] ), .IN1(
        \SUMB[632][2] ), .COUT(\CARRYB[633][1] ), .SUM(\SUMB[633][1] ) );
  FADDER S3_633_2 ( .CIN(\ab[633][2] ), .IN0(\CARRYB[632][2] ), .IN1(
        \ab[632][3] ), .COUT(\CARRYB[633][2] ), .SUM(\SUMB[633][2] ) );
  FADDER S1_632_0 ( .CIN(\ab[632][0] ), .IN0(\CARRYB[631][0] ), .IN1(
        \SUMB[631][1] ), .COUT(\CARRYB[632][0] ), .SUM(PRODUCT[632]) );
  FADDER S2_632_1 ( .CIN(\ab[632][1] ), .IN0(\CARRYB[631][1] ), .IN1(
        \SUMB[631][2] ), .COUT(\CARRYB[632][1] ), .SUM(\SUMB[632][1] ) );
  FADDER S3_632_2 ( .CIN(\ab[632][2] ), .IN0(\CARRYB[631][2] ), .IN1(
        \ab[631][3] ), .COUT(\CARRYB[632][2] ), .SUM(\SUMB[632][2] ) );
  FADDER S1_631_0 ( .CIN(\ab[631][0] ), .IN0(\CARRYB[630][0] ), .IN1(
        \SUMB[630][1] ), .COUT(\CARRYB[631][0] ), .SUM(PRODUCT[631]) );
  FADDER S2_631_1 ( .CIN(\ab[631][1] ), .IN0(\CARRYB[630][1] ), .IN1(
        \SUMB[630][2] ), .COUT(\CARRYB[631][1] ), .SUM(\SUMB[631][1] ) );
  FADDER S3_631_2 ( .CIN(\ab[631][2] ), .IN0(\CARRYB[630][2] ), .IN1(
        \ab[630][3] ), .COUT(\CARRYB[631][2] ), .SUM(\SUMB[631][2] ) );
  FADDER S1_630_0 ( .CIN(\ab[630][0] ), .IN0(\CARRYB[629][0] ), .IN1(
        \SUMB[629][1] ), .COUT(\CARRYB[630][0] ), .SUM(PRODUCT[630]) );
  FADDER S2_630_1 ( .CIN(\ab[630][1] ), .IN0(\CARRYB[629][1] ), .IN1(
        \SUMB[629][2] ), .COUT(\CARRYB[630][1] ), .SUM(\SUMB[630][1] ) );
  FADDER S3_630_2 ( .CIN(\ab[630][2] ), .IN0(\CARRYB[629][2] ), .IN1(
        \ab[629][3] ), .COUT(\CARRYB[630][2] ), .SUM(\SUMB[630][2] ) );
  FADDER S1_629_0 ( .CIN(\ab[629][0] ), .IN0(\CARRYB[628][0] ), .IN1(
        \SUMB[628][1] ), .COUT(\CARRYB[629][0] ), .SUM(PRODUCT[629]) );
  FADDER S2_629_1 ( .CIN(\ab[629][1] ), .IN0(\CARRYB[628][1] ), .IN1(
        \SUMB[628][2] ), .COUT(\CARRYB[629][1] ), .SUM(\SUMB[629][1] ) );
  FADDER S3_629_2 ( .CIN(\ab[629][2] ), .IN0(\CARRYB[628][2] ), .IN1(
        \ab[628][3] ), .COUT(\CARRYB[629][2] ), .SUM(\SUMB[629][2] ) );
  FADDER S1_628_0 ( .CIN(\ab[628][0] ), .IN0(\CARRYB[627][0] ), .IN1(
        \SUMB[627][1] ), .COUT(\CARRYB[628][0] ), .SUM(PRODUCT[628]) );
  FADDER S2_628_1 ( .CIN(\ab[628][1] ), .IN0(\CARRYB[627][1] ), .IN1(
        \SUMB[627][2] ), .COUT(\CARRYB[628][1] ), .SUM(\SUMB[628][1] ) );
  FADDER S3_628_2 ( .CIN(\ab[628][2] ), .IN0(\CARRYB[627][2] ), .IN1(
        \ab[627][3] ), .COUT(\CARRYB[628][2] ), .SUM(\SUMB[628][2] ) );
  FADDER S1_627_0 ( .CIN(\ab[627][0] ), .IN0(\CARRYB[626][0] ), .IN1(
        \SUMB[626][1] ), .COUT(\CARRYB[627][0] ), .SUM(PRODUCT[627]) );
  FADDER S2_627_1 ( .CIN(\ab[627][1] ), .IN0(\CARRYB[626][1] ), .IN1(
        \SUMB[626][2] ), .COUT(\CARRYB[627][1] ), .SUM(\SUMB[627][1] ) );
  FADDER S3_627_2 ( .CIN(\ab[627][2] ), .IN0(\CARRYB[626][2] ), .IN1(
        \ab[626][3] ), .COUT(\CARRYB[627][2] ), .SUM(\SUMB[627][2] ) );
  FADDER S1_626_0 ( .CIN(\ab[626][0] ), .IN0(\CARRYB[625][0] ), .IN1(
        \SUMB[625][1] ), .COUT(\CARRYB[626][0] ), .SUM(PRODUCT[626]) );
  FADDER S2_626_1 ( .CIN(\ab[626][1] ), .IN0(\CARRYB[625][1] ), .IN1(
        \SUMB[625][2] ), .COUT(\CARRYB[626][1] ), .SUM(\SUMB[626][1] ) );
  FADDER S3_626_2 ( .CIN(\ab[626][2] ), .IN0(\CARRYB[625][2] ), .IN1(
        \ab[625][3] ), .COUT(\CARRYB[626][2] ), .SUM(\SUMB[626][2] ) );
  FADDER S1_625_0 ( .CIN(\ab[625][0] ), .IN0(\CARRYB[624][0] ), .IN1(
        \SUMB[624][1] ), .COUT(\CARRYB[625][0] ), .SUM(PRODUCT[625]) );
  FADDER S2_625_1 ( .CIN(\ab[625][1] ), .IN0(\CARRYB[624][1] ), .IN1(
        \SUMB[624][2] ), .COUT(\CARRYB[625][1] ), .SUM(\SUMB[625][1] ) );
  FADDER S3_625_2 ( .CIN(\ab[625][2] ), .IN0(\CARRYB[624][2] ), .IN1(
        \ab[624][3] ), .COUT(\CARRYB[625][2] ), .SUM(\SUMB[625][2] ) );
  FADDER S1_624_0 ( .CIN(\ab[624][0] ), .IN0(\CARRYB[623][0] ), .IN1(
        \SUMB[623][1] ), .COUT(\CARRYB[624][0] ), .SUM(PRODUCT[624]) );
  FADDER S2_624_1 ( .CIN(\ab[624][1] ), .IN0(\CARRYB[623][1] ), .IN1(
        \SUMB[623][2] ), .COUT(\CARRYB[624][1] ), .SUM(\SUMB[624][1] ) );
  FADDER S3_624_2 ( .CIN(\ab[624][2] ), .IN0(\CARRYB[623][2] ), .IN1(
        \ab[623][3] ), .COUT(\CARRYB[624][2] ), .SUM(\SUMB[624][2] ) );
  FADDER S1_623_0 ( .CIN(\ab[623][0] ), .IN0(\CARRYB[622][0] ), .IN1(
        \SUMB[622][1] ), .COUT(\CARRYB[623][0] ), .SUM(PRODUCT[623]) );
  FADDER S2_623_1 ( .CIN(\ab[623][1] ), .IN0(\CARRYB[622][1] ), .IN1(
        \SUMB[622][2] ), .COUT(\CARRYB[623][1] ), .SUM(\SUMB[623][1] ) );
  FADDER S3_623_2 ( .CIN(\ab[623][2] ), .IN0(\CARRYB[622][2] ), .IN1(
        \ab[622][3] ), .COUT(\CARRYB[623][2] ), .SUM(\SUMB[623][2] ) );
  FADDER S1_622_0 ( .CIN(\ab[622][0] ), .IN0(\CARRYB[621][0] ), .IN1(
        \SUMB[621][1] ), .COUT(\CARRYB[622][0] ), .SUM(PRODUCT[622]) );
  FADDER S2_622_1 ( .CIN(\ab[622][1] ), .IN0(\CARRYB[621][1] ), .IN1(
        \SUMB[621][2] ), .COUT(\CARRYB[622][1] ), .SUM(\SUMB[622][1] ) );
  FADDER S3_622_2 ( .CIN(\ab[622][2] ), .IN0(\CARRYB[621][2] ), .IN1(
        \ab[621][3] ), .COUT(\CARRYB[622][2] ), .SUM(\SUMB[622][2] ) );
  FADDER S1_621_0 ( .CIN(\ab[621][0] ), .IN0(\CARRYB[620][0] ), .IN1(
        \SUMB[620][1] ), .COUT(\CARRYB[621][0] ), .SUM(PRODUCT[621]) );
  FADDER S2_621_1 ( .CIN(\ab[621][1] ), .IN0(\CARRYB[620][1] ), .IN1(
        \SUMB[620][2] ), .COUT(\CARRYB[621][1] ), .SUM(\SUMB[621][1] ) );
  FADDER S3_621_2 ( .CIN(\ab[621][2] ), .IN0(\CARRYB[620][2] ), .IN1(
        \ab[620][3] ), .COUT(\CARRYB[621][2] ), .SUM(\SUMB[621][2] ) );
  FADDER S1_620_0 ( .CIN(\ab[620][0] ), .IN0(\CARRYB[619][0] ), .IN1(
        \SUMB[619][1] ), .COUT(\CARRYB[620][0] ), .SUM(PRODUCT[620]) );
  FADDER S2_620_1 ( .CIN(\ab[620][1] ), .IN0(\CARRYB[619][1] ), .IN1(
        \SUMB[619][2] ), .COUT(\CARRYB[620][1] ), .SUM(\SUMB[620][1] ) );
  FADDER S3_620_2 ( .CIN(\ab[620][2] ), .IN0(\CARRYB[619][2] ), .IN1(
        \ab[619][3] ), .COUT(\CARRYB[620][2] ), .SUM(\SUMB[620][2] ) );
  FADDER S1_619_0 ( .CIN(\ab[619][0] ), .IN0(\CARRYB[618][0] ), .IN1(
        \SUMB[618][1] ), .COUT(\CARRYB[619][0] ), .SUM(PRODUCT[619]) );
  FADDER S2_619_1 ( .CIN(\ab[619][1] ), .IN0(\CARRYB[618][1] ), .IN1(
        \SUMB[618][2] ), .COUT(\CARRYB[619][1] ), .SUM(\SUMB[619][1] ) );
  FADDER S3_619_2 ( .CIN(\ab[619][2] ), .IN0(\CARRYB[618][2] ), .IN1(
        \ab[618][3] ), .COUT(\CARRYB[619][2] ), .SUM(\SUMB[619][2] ) );
  FADDER S1_618_0 ( .CIN(\ab[618][0] ), .IN0(\CARRYB[617][0] ), .IN1(
        \SUMB[617][1] ), .COUT(\CARRYB[618][0] ), .SUM(PRODUCT[618]) );
  FADDER S2_618_1 ( .CIN(\ab[618][1] ), .IN0(\CARRYB[617][1] ), .IN1(
        \SUMB[617][2] ), .COUT(\CARRYB[618][1] ), .SUM(\SUMB[618][1] ) );
  FADDER S3_618_2 ( .CIN(\ab[618][2] ), .IN0(\CARRYB[617][2] ), .IN1(
        \ab[617][3] ), .COUT(\CARRYB[618][2] ), .SUM(\SUMB[618][2] ) );
  FADDER S1_617_0 ( .CIN(\ab[617][0] ), .IN0(\CARRYB[616][0] ), .IN1(
        \SUMB[616][1] ), .COUT(\CARRYB[617][0] ), .SUM(PRODUCT[617]) );
  FADDER S2_617_1 ( .CIN(\ab[617][1] ), .IN0(\CARRYB[616][1] ), .IN1(
        \SUMB[616][2] ), .COUT(\CARRYB[617][1] ), .SUM(\SUMB[617][1] ) );
  FADDER S3_617_2 ( .CIN(\ab[617][2] ), .IN0(\CARRYB[616][2] ), .IN1(
        \ab[616][3] ), .COUT(\CARRYB[617][2] ), .SUM(\SUMB[617][2] ) );
  FADDER S1_616_0 ( .CIN(\ab[616][0] ), .IN0(\CARRYB[615][0] ), .IN1(
        \SUMB[615][1] ), .COUT(\CARRYB[616][0] ), .SUM(PRODUCT[616]) );
  FADDER S2_616_1 ( .CIN(\ab[616][1] ), .IN0(\CARRYB[615][1] ), .IN1(
        \SUMB[615][2] ), .COUT(\CARRYB[616][1] ), .SUM(\SUMB[616][1] ) );
  FADDER S3_616_2 ( .CIN(\ab[616][2] ), .IN0(\CARRYB[615][2] ), .IN1(
        \ab[615][3] ), .COUT(\CARRYB[616][2] ), .SUM(\SUMB[616][2] ) );
  FADDER S1_615_0 ( .CIN(\ab[615][0] ), .IN0(\CARRYB[614][0] ), .IN1(
        \SUMB[614][1] ), .COUT(\CARRYB[615][0] ), .SUM(PRODUCT[615]) );
  FADDER S2_615_1 ( .CIN(\ab[615][1] ), .IN0(\CARRYB[614][1] ), .IN1(
        \SUMB[614][2] ), .COUT(\CARRYB[615][1] ), .SUM(\SUMB[615][1] ) );
  FADDER S3_615_2 ( .CIN(\ab[615][2] ), .IN0(\CARRYB[614][2] ), .IN1(
        \ab[614][3] ), .COUT(\CARRYB[615][2] ), .SUM(\SUMB[615][2] ) );
  FADDER S1_614_0 ( .CIN(\ab[614][0] ), .IN0(\CARRYB[613][0] ), .IN1(
        \SUMB[613][1] ), .COUT(\CARRYB[614][0] ), .SUM(PRODUCT[614]) );
  FADDER S2_614_1 ( .CIN(\ab[614][1] ), .IN0(\CARRYB[613][1] ), .IN1(
        \SUMB[613][2] ), .COUT(\CARRYB[614][1] ), .SUM(\SUMB[614][1] ) );
  FADDER S3_614_2 ( .CIN(\ab[614][2] ), .IN0(\CARRYB[613][2] ), .IN1(
        \ab[613][3] ), .COUT(\CARRYB[614][2] ), .SUM(\SUMB[614][2] ) );
  FADDER S1_613_0 ( .CIN(\ab[613][0] ), .IN0(\CARRYB[612][0] ), .IN1(
        \SUMB[612][1] ), .COUT(\CARRYB[613][0] ), .SUM(PRODUCT[613]) );
  FADDER S2_613_1 ( .CIN(\ab[613][1] ), .IN0(\CARRYB[612][1] ), .IN1(
        \SUMB[612][2] ), .COUT(\CARRYB[613][1] ), .SUM(\SUMB[613][1] ) );
  FADDER S3_613_2 ( .CIN(\ab[613][2] ), .IN0(\CARRYB[612][2] ), .IN1(
        \ab[612][3] ), .COUT(\CARRYB[613][2] ), .SUM(\SUMB[613][2] ) );
  FADDER S1_612_0 ( .CIN(\ab[612][0] ), .IN0(\CARRYB[611][0] ), .IN1(
        \SUMB[611][1] ), .COUT(\CARRYB[612][0] ), .SUM(PRODUCT[612]) );
  FADDER S2_612_1 ( .CIN(\ab[612][1] ), .IN0(\CARRYB[611][1] ), .IN1(
        \SUMB[611][2] ), .COUT(\CARRYB[612][1] ), .SUM(\SUMB[612][1] ) );
  FADDER S3_612_2 ( .CIN(\ab[612][2] ), .IN0(\CARRYB[611][2] ), .IN1(
        \ab[611][3] ), .COUT(\CARRYB[612][2] ), .SUM(\SUMB[612][2] ) );
  FADDER S1_611_0 ( .CIN(\ab[611][0] ), .IN0(\CARRYB[610][0] ), .IN1(
        \SUMB[610][1] ), .COUT(\CARRYB[611][0] ), .SUM(PRODUCT[611]) );
  FADDER S2_611_1 ( .CIN(\ab[611][1] ), .IN0(\CARRYB[610][1] ), .IN1(
        \SUMB[610][2] ), .COUT(\CARRYB[611][1] ), .SUM(\SUMB[611][1] ) );
  FADDER S3_611_2 ( .CIN(\ab[611][2] ), .IN0(\CARRYB[610][2] ), .IN1(
        \ab[610][3] ), .COUT(\CARRYB[611][2] ), .SUM(\SUMB[611][2] ) );
  FADDER S1_610_0 ( .CIN(\ab[610][0] ), .IN0(\CARRYB[609][0] ), .IN1(
        \SUMB[609][1] ), .COUT(\CARRYB[610][0] ), .SUM(PRODUCT[610]) );
  FADDER S2_610_1 ( .CIN(\ab[610][1] ), .IN0(\CARRYB[609][1] ), .IN1(
        \SUMB[609][2] ), .COUT(\CARRYB[610][1] ), .SUM(\SUMB[610][1] ) );
  FADDER S3_610_2 ( .CIN(\ab[610][2] ), .IN0(\CARRYB[609][2] ), .IN1(
        \ab[609][3] ), .COUT(\CARRYB[610][2] ), .SUM(\SUMB[610][2] ) );
  FADDER S1_609_0 ( .CIN(\ab[609][0] ), .IN0(\CARRYB[608][0] ), .IN1(
        \SUMB[608][1] ), .COUT(\CARRYB[609][0] ), .SUM(PRODUCT[609]) );
  FADDER S2_609_1 ( .CIN(\ab[609][1] ), .IN0(\CARRYB[608][1] ), .IN1(
        \SUMB[608][2] ), .COUT(\CARRYB[609][1] ), .SUM(\SUMB[609][1] ) );
  FADDER S3_609_2 ( .CIN(\ab[609][2] ), .IN0(\CARRYB[608][2] ), .IN1(
        \ab[608][3] ), .COUT(\CARRYB[609][2] ), .SUM(\SUMB[609][2] ) );
  FADDER S1_608_0 ( .CIN(\ab[608][0] ), .IN0(\CARRYB[607][0] ), .IN1(
        \SUMB[607][1] ), .COUT(\CARRYB[608][0] ), .SUM(PRODUCT[608]) );
  FADDER S2_608_1 ( .CIN(\ab[608][1] ), .IN0(\CARRYB[607][1] ), .IN1(
        \SUMB[607][2] ), .COUT(\CARRYB[608][1] ), .SUM(\SUMB[608][1] ) );
  FADDER S3_608_2 ( .CIN(\ab[608][2] ), .IN0(\CARRYB[607][2] ), .IN1(
        \ab[607][3] ), .COUT(\CARRYB[608][2] ), .SUM(\SUMB[608][2] ) );
  FADDER S1_607_0 ( .CIN(\ab[607][0] ), .IN0(\CARRYB[606][0] ), .IN1(
        \SUMB[606][1] ), .COUT(\CARRYB[607][0] ), .SUM(PRODUCT[607]) );
  FADDER S2_607_1 ( .CIN(\ab[607][1] ), .IN0(\CARRYB[606][1] ), .IN1(
        \SUMB[606][2] ), .COUT(\CARRYB[607][1] ), .SUM(\SUMB[607][1] ) );
  FADDER S3_607_2 ( .CIN(\ab[607][2] ), .IN0(\CARRYB[606][2] ), .IN1(
        \ab[606][3] ), .COUT(\CARRYB[607][2] ), .SUM(\SUMB[607][2] ) );
  FADDER S1_606_0 ( .CIN(\ab[606][0] ), .IN0(\CARRYB[605][0] ), .IN1(
        \SUMB[605][1] ), .COUT(\CARRYB[606][0] ), .SUM(PRODUCT[606]) );
  FADDER S2_606_1 ( .CIN(\ab[606][1] ), .IN0(\CARRYB[605][1] ), .IN1(
        \SUMB[605][2] ), .COUT(\CARRYB[606][1] ), .SUM(\SUMB[606][1] ) );
  FADDER S3_606_2 ( .CIN(\ab[606][2] ), .IN0(\CARRYB[605][2] ), .IN1(
        \ab[605][3] ), .COUT(\CARRYB[606][2] ), .SUM(\SUMB[606][2] ) );
  FADDER S1_605_0 ( .CIN(\ab[605][0] ), .IN0(\CARRYB[604][0] ), .IN1(
        \SUMB[604][1] ), .COUT(\CARRYB[605][0] ), .SUM(PRODUCT[605]) );
  FADDER S2_605_1 ( .CIN(\ab[605][1] ), .IN0(\CARRYB[604][1] ), .IN1(
        \SUMB[604][2] ), .COUT(\CARRYB[605][1] ), .SUM(\SUMB[605][1] ) );
  FADDER S3_605_2 ( .CIN(\ab[605][2] ), .IN0(\CARRYB[604][2] ), .IN1(
        \ab[604][3] ), .COUT(\CARRYB[605][2] ), .SUM(\SUMB[605][2] ) );
  FADDER S1_604_0 ( .CIN(\ab[604][0] ), .IN0(\CARRYB[603][0] ), .IN1(
        \SUMB[603][1] ), .COUT(\CARRYB[604][0] ), .SUM(PRODUCT[604]) );
  FADDER S2_604_1 ( .CIN(\ab[604][1] ), .IN0(\CARRYB[603][1] ), .IN1(
        \SUMB[603][2] ), .COUT(\CARRYB[604][1] ), .SUM(\SUMB[604][1] ) );
  FADDER S3_604_2 ( .CIN(\ab[604][2] ), .IN0(\CARRYB[603][2] ), .IN1(
        \ab[603][3] ), .COUT(\CARRYB[604][2] ), .SUM(\SUMB[604][2] ) );
  FADDER S1_603_0 ( .CIN(\ab[603][0] ), .IN0(\CARRYB[602][0] ), .IN1(
        \SUMB[602][1] ), .COUT(\CARRYB[603][0] ), .SUM(PRODUCT[603]) );
  FADDER S2_603_1 ( .CIN(\ab[603][1] ), .IN0(\CARRYB[602][1] ), .IN1(
        \SUMB[602][2] ), .COUT(\CARRYB[603][1] ), .SUM(\SUMB[603][1] ) );
  FADDER S3_603_2 ( .CIN(\ab[603][2] ), .IN0(\CARRYB[602][2] ), .IN1(
        \ab[602][3] ), .COUT(\CARRYB[603][2] ), .SUM(\SUMB[603][2] ) );
  FADDER S1_602_0 ( .CIN(\ab[602][0] ), .IN0(\CARRYB[601][0] ), .IN1(
        \SUMB[601][1] ), .COUT(\CARRYB[602][0] ), .SUM(PRODUCT[602]) );
  FADDER S2_602_1 ( .CIN(\ab[602][1] ), .IN0(\CARRYB[601][1] ), .IN1(
        \SUMB[601][2] ), .COUT(\CARRYB[602][1] ), .SUM(\SUMB[602][1] ) );
  FADDER S3_602_2 ( .CIN(\ab[602][2] ), .IN0(\CARRYB[601][2] ), .IN1(
        \ab[601][3] ), .COUT(\CARRYB[602][2] ), .SUM(\SUMB[602][2] ) );
  FADDER S1_601_0 ( .CIN(\ab[601][0] ), .IN0(\CARRYB[600][0] ), .IN1(
        \SUMB[600][1] ), .COUT(\CARRYB[601][0] ), .SUM(PRODUCT[601]) );
  FADDER S2_601_1 ( .CIN(\ab[601][1] ), .IN0(\CARRYB[600][1] ), .IN1(
        \SUMB[600][2] ), .COUT(\CARRYB[601][1] ), .SUM(\SUMB[601][1] ) );
  FADDER S3_601_2 ( .CIN(\ab[601][2] ), .IN0(\CARRYB[600][2] ), .IN1(
        \ab[600][3] ), .COUT(\CARRYB[601][2] ), .SUM(\SUMB[601][2] ) );
  FADDER S1_600_0 ( .CIN(\ab[600][0] ), .IN0(\CARRYB[599][0] ), .IN1(
        \SUMB[599][1] ), .COUT(\CARRYB[600][0] ), .SUM(PRODUCT[600]) );
  FADDER S2_600_1 ( .CIN(\ab[600][1] ), .IN0(\CARRYB[599][1] ), .IN1(
        \SUMB[599][2] ), .COUT(\CARRYB[600][1] ), .SUM(\SUMB[600][1] ) );
  FADDER S3_600_2 ( .CIN(\ab[600][2] ), .IN0(\CARRYB[599][2] ), .IN1(
        \ab[599][3] ), .COUT(\CARRYB[600][2] ), .SUM(\SUMB[600][2] ) );
  FADDER S1_599_0 ( .CIN(\ab[599][0] ), .IN0(\CARRYB[598][0] ), .IN1(
        \SUMB[598][1] ), .COUT(\CARRYB[599][0] ), .SUM(PRODUCT[599]) );
  FADDER S2_599_1 ( .CIN(\ab[599][1] ), .IN0(\CARRYB[598][1] ), .IN1(
        \SUMB[598][2] ), .COUT(\CARRYB[599][1] ), .SUM(\SUMB[599][1] ) );
  FADDER S3_599_2 ( .CIN(\ab[599][2] ), .IN0(\CARRYB[598][2] ), .IN1(
        \ab[598][3] ), .COUT(\CARRYB[599][2] ), .SUM(\SUMB[599][2] ) );
  FADDER S1_598_0 ( .CIN(\ab[598][0] ), .IN0(\CARRYB[597][0] ), .IN1(
        \SUMB[597][1] ), .COUT(\CARRYB[598][0] ), .SUM(PRODUCT[598]) );
  FADDER S2_598_1 ( .CIN(\ab[598][1] ), .IN0(\CARRYB[597][1] ), .IN1(
        \SUMB[597][2] ), .COUT(\CARRYB[598][1] ), .SUM(\SUMB[598][1] ) );
  FADDER S3_598_2 ( .CIN(\ab[598][2] ), .IN0(\CARRYB[597][2] ), .IN1(
        \ab[597][3] ), .COUT(\CARRYB[598][2] ), .SUM(\SUMB[598][2] ) );
  FADDER S1_597_0 ( .CIN(\ab[597][0] ), .IN0(\CARRYB[596][0] ), .IN1(
        \SUMB[596][1] ), .COUT(\CARRYB[597][0] ), .SUM(PRODUCT[597]) );
  FADDER S2_597_1 ( .CIN(\ab[597][1] ), .IN0(\CARRYB[596][1] ), .IN1(
        \SUMB[596][2] ), .COUT(\CARRYB[597][1] ), .SUM(\SUMB[597][1] ) );
  FADDER S3_597_2 ( .CIN(\ab[597][2] ), .IN0(\CARRYB[596][2] ), .IN1(
        \ab[596][3] ), .COUT(\CARRYB[597][2] ), .SUM(\SUMB[597][2] ) );
  FADDER S1_596_0 ( .CIN(\ab[596][0] ), .IN0(\CARRYB[595][0] ), .IN1(
        \SUMB[595][1] ), .COUT(\CARRYB[596][0] ), .SUM(PRODUCT[596]) );
  FADDER S2_596_1 ( .CIN(\ab[596][1] ), .IN0(\CARRYB[595][1] ), .IN1(
        \SUMB[595][2] ), .COUT(\CARRYB[596][1] ), .SUM(\SUMB[596][1] ) );
  FADDER S3_596_2 ( .CIN(\ab[596][2] ), .IN0(\CARRYB[595][2] ), .IN1(
        \ab[595][3] ), .COUT(\CARRYB[596][2] ), .SUM(\SUMB[596][2] ) );
  FADDER S1_595_0 ( .CIN(\ab[595][0] ), .IN0(\CARRYB[594][0] ), .IN1(
        \SUMB[594][1] ), .COUT(\CARRYB[595][0] ), .SUM(PRODUCT[595]) );
  FADDER S2_595_1 ( .CIN(\ab[595][1] ), .IN0(\CARRYB[594][1] ), .IN1(
        \SUMB[594][2] ), .COUT(\CARRYB[595][1] ), .SUM(\SUMB[595][1] ) );
  FADDER S3_595_2 ( .CIN(\ab[595][2] ), .IN0(\CARRYB[594][2] ), .IN1(
        \ab[594][3] ), .COUT(\CARRYB[595][2] ), .SUM(\SUMB[595][2] ) );
  FADDER S1_594_0 ( .CIN(\ab[594][0] ), .IN0(\CARRYB[593][0] ), .IN1(
        \SUMB[593][1] ), .COUT(\CARRYB[594][0] ), .SUM(PRODUCT[594]) );
  FADDER S2_594_1 ( .CIN(\ab[594][1] ), .IN0(\CARRYB[593][1] ), .IN1(
        \SUMB[593][2] ), .COUT(\CARRYB[594][1] ), .SUM(\SUMB[594][1] ) );
  FADDER S3_594_2 ( .CIN(\ab[594][2] ), .IN0(\CARRYB[593][2] ), .IN1(
        \ab[593][3] ), .COUT(\CARRYB[594][2] ), .SUM(\SUMB[594][2] ) );
  FADDER S1_593_0 ( .CIN(\ab[593][0] ), .IN0(\CARRYB[592][0] ), .IN1(
        \SUMB[592][1] ), .COUT(\CARRYB[593][0] ), .SUM(PRODUCT[593]) );
  FADDER S2_593_1 ( .CIN(\ab[593][1] ), .IN0(\CARRYB[592][1] ), .IN1(
        \SUMB[592][2] ), .COUT(\CARRYB[593][1] ), .SUM(\SUMB[593][1] ) );
  FADDER S3_593_2 ( .CIN(\ab[593][2] ), .IN0(\CARRYB[592][2] ), .IN1(
        \ab[592][3] ), .COUT(\CARRYB[593][2] ), .SUM(\SUMB[593][2] ) );
  FADDER S1_592_0 ( .CIN(\ab[592][0] ), .IN0(\CARRYB[591][0] ), .IN1(
        \SUMB[591][1] ), .COUT(\CARRYB[592][0] ), .SUM(PRODUCT[592]) );
  FADDER S2_592_1 ( .CIN(\ab[592][1] ), .IN0(\CARRYB[591][1] ), .IN1(
        \SUMB[591][2] ), .COUT(\CARRYB[592][1] ), .SUM(\SUMB[592][1] ) );
  FADDER S3_592_2 ( .CIN(\ab[592][2] ), .IN0(\CARRYB[591][2] ), .IN1(
        \ab[591][3] ), .COUT(\CARRYB[592][2] ), .SUM(\SUMB[592][2] ) );
  FADDER S1_591_0 ( .CIN(\ab[591][0] ), .IN0(\CARRYB[590][0] ), .IN1(
        \SUMB[590][1] ), .COUT(\CARRYB[591][0] ), .SUM(PRODUCT[591]) );
  FADDER S2_591_1 ( .CIN(\ab[591][1] ), .IN0(\CARRYB[590][1] ), .IN1(
        \SUMB[590][2] ), .COUT(\CARRYB[591][1] ), .SUM(\SUMB[591][1] ) );
  FADDER S3_591_2 ( .CIN(\ab[591][2] ), .IN0(\CARRYB[590][2] ), .IN1(
        \ab[590][3] ), .COUT(\CARRYB[591][2] ), .SUM(\SUMB[591][2] ) );
  FADDER S1_590_0 ( .CIN(\ab[590][0] ), .IN0(\CARRYB[589][0] ), .IN1(
        \SUMB[589][1] ), .COUT(\CARRYB[590][0] ), .SUM(PRODUCT[590]) );
  FADDER S2_590_1 ( .CIN(\ab[590][1] ), .IN0(\CARRYB[589][1] ), .IN1(
        \SUMB[589][2] ), .COUT(\CARRYB[590][1] ), .SUM(\SUMB[590][1] ) );
  FADDER S3_590_2 ( .CIN(\ab[590][2] ), .IN0(\CARRYB[589][2] ), .IN1(
        \ab[589][3] ), .COUT(\CARRYB[590][2] ), .SUM(\SUMB[590][2] ) );
  FADDER S1_589_0 ( .CIN(\ab[589][0] ), .IN0(\CARRYB[588][0] ), .IN1(
        \SUMB[588][1] ), .COUT(\CARRYB[589][0] ), .SUM(PRODUCT[589]) );
  FADDER S2_589_1 ( .CIN(\ab[589][1] ), .IN0(\CARRYB[588][1] ), .IN1(
        \SUMB[588][2] ), .COUT(\CARRYB[589][1] ), .SUM(\SUMB[589][1] ) );
  FADDER S3_589_2 ( .CIN(\ab[589][2] ), .IN0(\CARRYB[588][2] ), .IN1(
        \ab[588][3] ), .COUT(\CARRYB[589][2] ), .SUM(\SUMB[589][2] ) );
  FADDER S1_588_0 ( .CIN(\ab[588][0] ), .IN0(\CARRYB[587][0] ), .IN1(
        \SUMB[587][1] ), .COUT(\CARRYB[588][0] ), .SUM(PRODUCT[588]) );
  FADDER S2_588_1 ( .CIN(\ab[588][1] ), .IN0(\CARRYB[587][1] ), .IN1(
        \SUMB[587][2] ), .COUT(\CARRYB[588][1] ), .SUM(\SUMB[588][1] ) );
  FADDER S3_588_2 ( .CIN(\ab[588][2] ), .IN0(\CARRYB[587][2] ), .IN1(
        \ab[587][3] ), .COUT(\CARRYB[588][2] ), .SUM(\SUMB[588][2] ) );
  FADDER S1_587_0 ( .CIN(\ab[587][0] ), .IN0(\CARRYB[586][0] ), .IN1(
        \SUMB[586][1] ), .COUT(\CARRYB[587][0] ), .SUM(PRODUCT[587]) );
  FADDER S2_587_1 ( .CIN(\ab[587][1] ), .IN0(\CARRYB[586][1] ), .IN1(
        \SUMB[586][2] ), .COUT(\CARRYB[587][1] ), .SUM(\SUMB[587][1] ) );
  FADDER S3_587_2 ( .CIN(\ab[587][2] ), .IN0(\CARRYB[586][2] ), .IN1(
        \ab[586][3] ), .COUT(\CARRYB[587][2] ), .SUM(\SUMB[587][2] ) );
  FADDER S1_586_0 ( .CIN(\ab[586][0] ), .IN0(\CARRYB[585][0] ), .IN1(
        \SUMB[585][1] ), .COUT(\CARRYB[586][0] ), .SUM(PRODUCT[586]) );
  FADDER S2_586_1 ( .CIN(\ab[586][1] ), .IN0(\CARRYB[585][1] ), .IN1(
        \SUMB[585][2] ), .COUT(\CARRYB[586][1] ), .SUM(\SUMB[586][1] ) );
  FADDER S3_586_2 ( .CIN(\ab[586][2] ), .IN0(\CARRYB[585][2] ), .IN1(
        \ab[585][3] ), .COUT(\CARRYB[586][2] ), .SUM(\SUMB[586][2] ) );
  FADDER S1_585_0 ( .CIN(\ab[585][0] ), .IN0(\CARRYB[584][0] ), .IN1(
        \SUMB[584][1] ), .COUT(\CARRYB[585][0] ), .SUM(PRODUCT[585]) );
  FADDER S2_585_1 ( .CIN(\ab[585][1] ), .IN0(\CARRYB[584][1] ), .IN1(
        \SUMB[584][2] ), .COUT(\CARRYB[585][1] ), .SUM(\SUMB[585][1] ) );
  FADDER S3_585_2 ( .CIN(\ab[585][2] ), .IN0(\CARRYB[584][2] ), .IN1(
        \ab[584][3] ), .COUT(\CARRYB[585][2] ), .SUM(\SUMB[585][2] ) );
  FADDER S1_584_0 ( .CIN(\ab[584][0] ), .IN0(\CARRYB[583][0] ), .IN1(
        \SUMB[583][1] ), .COUT(\CARRYB[584][0] ), .SUM(PRODUCT[584]) );
  FADDER S2_584_1 ( .CIN(\ab[584][1] ), .IN0(\CARRYB[583][1] ), .IN1(
        \SUMB[583][2] ), .COUT(\CARRYB[584][1] ), .SUM(\SUMB[584][1] ) );
  FADDER S3_584_2 ( .CIN(\ab[584][2] ), .IN0(\CARRYB[583][2] ), .IN1(
        \ab[583][3] ), .COUT(\CARRYB[584][2] ), .SUM(\SUMB[584][2] ) );
  FADDER S1_583_0 ( .CIN(\ab[583][0] ), .IN0(\CARRYB[582][0] ), .IN1(
        \SUMB[582][1] ), .COUT(\CARRYB[583][0] ), .SUM(PRODUCT[583]) );
  FADDER S2_583_1 ( .CIN(\ab[583][1] ), .IN0(\CARRYB[582][1] ), .IN1(
        \SUMB[582][2] ), .COUT(\CARRYB[583][1] ), .SUM(\SUMB[583][1] ) );
  FADDER S3_583_2 ( .CIN(\ab[583][2] ), .IN0(\CARRYB[582][2] ), .IN1(
        \ab[582][3] ), .COUT(\CARRYB[583][2] ), .SUM(\SUMB[583][2] ) );
  FADDER S1_582_0 ( .CIN(\ab[582][0] ), .IN0(\CARRYB[581][0] ), .IN1(
        \SUMB[581][1] ), .COUT(\CARRYB[582][0] ), .SUM(PRODUCT[582]) );
  FADDER S2_582_1 ( .CIN(\ab[582][1] ), .IN0(\CARRYB[581][1] ), .IN1(
        \SUMB[581][2] ), .COUT(\CARRYB[582][1] ), .SUM(\SUMB[582][1] ) );
  FADDER S3_582_2 ( .CIN(\ab[582][2] ), .IN0(\CARRYB[581][2] ), .IN1(
        \ab[581][3] ), .COUT(\CARRYB[582][2] ), .SUM(\SUMB[582][2] ) );
  FADDER S1_581_0 ( .CIN(\ab[581][0] ), .IN0(\CARRYB[580][0] ), .IN1(
        \SUMB[580][1] ), .COUT(\CARRYB[581][0] ), .SUM(PRODUCT[581]) );
  FADDER S2_581_1 ( .CIN(\ab[581][1] ), .IN0(\CARRYB[580][1] ), .IN1(
        \SUMB[580][2] ), .COUT(\CARRYB[581][1] ), .SUM(\SUMB[581][1] ) );
  FADDER S3_581_2 ( .CIN(\ab[581][2] ), .IN0(\CARRYB[580][2] ), .IN1(
        \ab[580][3] ), .COUT(\CARRYB[581][2] ), .SUM(\SUMB[581][2] ) );
  FADDER S1_580_0 ( .CIN(\ab[580][0] ), .IN0(\CARRYB[579][0] ), .IN1(
        \SUMB[579][1] ), .COUT(\CARRYB[580][0] ), .SUM(PRODUCT[580]) );
  FADDER S2_580_1 ( .CIN(\ab[580][1] ), .IN0(\CARRYB[579][1] ), .IN1(
        \SUMB[579][2] ), .COUT(\CARRYB[580][1] ), .SUM(\SUMB[580][1] ) );
  FADDER S3_580_2 ( .CIN(\ab[580][2] ), .IN0(\CARRYB[579][2] ), .IN1(
        \ab[579][3] ), .COUT(\CARRYB[580][2] ), .SUM(\SUMB[580][2] ) );
  FADDER S1_579_0 ( .CIN(\ab[579][0] ), .IN0(\CARRYB[578][0] ), .IN1(
        \SUMB[578][1] ), .COUT(\CARRYB[579][0] ), .SUM(PRODUCT[579]) );
  FADDER S2_579_1 ( .CIN(\ab[579][1] ), .IN0(\CARRYB[578][1] ), .IN1(
        \SUMB[578][2] ), .COUT(\CARRYB[579][1] ), .SUM(\SUMB[579][1] ) );
  FADDER S3_579_2 ( .CIN(\ab[579][2] ), .IN0(\CARRYB[578][2] ), .IN1(
        \ab[578][3] ), .COUT(\CARRYB[579][2] ), .SUM(\SUMB[579][2] ) );
  FADDER S1_578_0 ( .CIN(\ab[578][0] ), .IN0(\CARRYB[577][0] ), .IN1(
        \SUMB[577][1] ), .COUT(\CARRYB[578][0] ), .SUM(PRODUCT[578]) );
  FADDER S2_578_1 ( .CIN(\ab[578][1] ), .IN0(\CARRYB[577][1] ), .IN1(
        \SUMB[577][2] ), .COUT(\CARRYB[578][1] ), .SUM(\SUMB[578][1] ) );
  FADDER S3_578_2 ( .CIN(\ab[578][2] ), .IN0(\CARRYB[577][2] ), .IN1(
        \ab[577][3] ), .COUT(\CARRYB[578][2] ), .SUM(\SUMB[578][2] ) );
  FADDER S1_577_0 ( .CIN(\ab[577][0] ), .IN0(\CARRYB[576][0] ), .IN1(
        \SUMB[576][1] ), .COUT(\CARRYB[577][0] ), .SUM(PRODUCT[577]) );
  FADDER S2_577_1 ( .CIN(\ab[577][1] ), .IN0(\CARRYB[576][1] ), .IN1(
        \SUMB[576][2] ), .COUT(\CARRYB[577][1] ), .SUM(\SUMB[577][1] ) );
  FADDER S3_577_2 ( .CIN(\ab[577][2] ), .IN0(\CARRYB[576][2] ), .IN1(
        \ab[576][3] ), .COUT(\CARRYB[577][2] ), .SUM(\SUMB[577][2] ) );
  FADDER S1_576_0 ( .CIN(\ab[576][0] ), .IN0(\CARRYB[575][0] ), .IN1(
        \SUMB[575][1] ), .COUT(\CARRYB[576][0] ), .SUM(PRODUCT[576]) );
  FADDER S2_576_1 ( .CIN(\ab[576][1] ), .IN0(\CARRYB[575][1] ), .IN1(
        \SUMB[575][2] ), .COUT(\CARRYB[576][1] ), .SUM(\SUMB[576][1] ) );
  FADDER S3_576_2 ( .CIN(\ab[576][2] ), .IN0(\CARRYB[575][2] ), .IN1(
        \ab[575][3] ), .COUT(\CARRYB[576][2] ), .SUM(\SUMB[576][2] ) );
  FADDER S1_575_0 ( .CIN(\ab[575][0] ), .IN0(\CARRYB[574][0] ), .IN1(
        \SUMB[574][1] ), .COUT(\CARRYB[575][0] ), .SUM(PRODUCT[575]) );
  FADDER S2_575_1 ( .CIN(\ab[575][1] ), .IN0(\CARRYB[574][1] ), .IN1(
        \SUMB[574][2] ), .COUT(\CARRYB[575][1] ), .SUM(\SUMB[575][1] ) );
  FADDER S3_575_2 ( .CIN(\ab[575][2] ), .IN0(\CARRYB[574][2] ), .IN1(
        \ab[574][3] ), .COUT(\CARRYB[575][2] ), .SUM(\SUMB[575][2] ) );
  FADDER S1_574_0 ( .CIN(\ab[574][0] ), .IN0(\CARRYB[573][0] ), .IN1(
        \SUMB[573][1] ), .COUT(\CARRYB[574][0] ), .SUM(PRODUCT[574]) );
  FADDER S2_574_1 ( .CIN(\ab[574][1] ), .IN0(\CARRYB[573][1] ), .IN1(
        \SUMB[573][2] ), .COUT(\CARRYB[574][1] ), .SUM(\SUMB[574][1] ) );
  FADDER S3_574_2 ( .CIN(\ab[574][2] ), .IN0(\CARRYB[573][2] ), .IN1(
        \ab[573][3] ), .COUT(\CARRYB[574][2] ), .SUM(\SUMB[574][2] ) );
  FADDER S1_573_0 ( .CIN(\ab[573][0] ), .IN0(\CARRYB[572][0] ), .IN1(
        \SUMB[572][1] ), .COUT(\CARRYB[573][0] ), .SUM(PRODUCT[573]) );
  FADDER S2_573_1 ( .CIN(\ab[573][1] ), .IN0(\CARRYB[572][1] ), .IN1(
        \SUMB[572][2] ), .COUT(\CARRYB[573][1] ), .SUM(\SUMB[573][1] ) );
  FADDER S3_573_2 ( .CIN(\ab[573][2] ), .IN0(\CARRYB[572][2] ), .IN1(
        \ab[572][3] ), .COUT(\CARRYB[573][2] ), .SUM(\SUMB[573][2] ) );
  FADDER S1_572_0 ( .CIN(\ab[572][0] ), .IN0(\CARRYB[571][0] ), .IN1(
        \SUMB[571][1] ), .COUT(\CARRYB[572][0] ), .SUM(PRODUCT[572]) );
  FADDER S2_572_1 ( .CIN(\ab[572][1] ), .IN0(\CARRYB[571][1] ), .IN1(
        \SUMB[571][2] ), .COUT(\CARRYB[572][1] ), .SUM(\SUMB[572][1] ) );
  FADDER S3_572_2 ( .CIN(\ab[572][2] ), .IN0(\CARRYB[571][2] ), .IN1(
        \ab[571][3] ), .COUT(\CARRYB[572][2] ), .SUM(\SUMB[572][2] ) );
  FADDER S1_571_0 ( .CIN(\ab[571][0] ), .IN0(\CARRYB[570][0] ), .IN1(
        \SUMB[570][1] ), .COUT(\CARRYB[571][0] ), .SUM(PRODUCT[571]) );
  FADDER S2_571_1 ( .CIN(\ab[571][1] ), .IN0(\CARRYB[570][1] ), .IN1(
        \SUMB[570][2] ), .COUT(\CARRYB[571][1] ), .SUM(\SUMB[571][1] ) );
  FADDER S3_571_2 ( .CIN(\ab[571][2] ), .IN0(\CARRYB[570][2] ), .IN1(
        \ab[570][3] ), .COUT(\CARRYB[571][2] ), .SUM(\SUMB[571][2] ) );
  FADDER S1_570_0 ( .CIN(\ab[570][0] ), .IN0(\CARRYB[569][0] ), .IN1(
        \SUMB[569][1] ), .COUT(\CARRYB[570][0] ), .SUM(PRODUCT[570]) );
  FADDER S2_570_1 ( .CIN(\ab[570][1] ), .IN0(\CARRYB[569][1] ), .IN1(
        \SUMB[569][2] ), .COUT(\CARRYB[570][1] ), .SUM(\SUMB[570][1] ) );
  FADDER S3_570_2 ( .CIN(\ab[570][2] ), .IN0(\CARRYB[569][2] ), .IN1(
        \ab[569][3] ), .COUT(\CARRYB[570][2] ), .SUM(\SUMB[570][2] ) );
  FADDER S1_569_0 ( .CIN(\ab[569][0] ), .IN0(\CARRYB[568][0] ), .IN1(
        \SUMB[568][1] ), .COUT(\CARRYB[569][0] ), .SUM(PRODUCT[569]) );
  FADDER S2_569_1 ( .CIN(\ab[569][1] ), .IN0(\CARRYB[568][1] ), .IN1(
        \SUMB[568][2] ), .COUT(\CARRYB[569][1] ), .SUM(\SUMB[569][1] ) );
  FADDER S3_569_2 ( .CIN(\ab[569][2] ), .IN0(\CARRYB[568][2] ), .IN1(
        \ab[568][3] ), .COUT(\CARRYB[569][2] ), .SUM(\SUMB[569][2] ) );
  FADDER S1_568_0 ( .CIN(\ab[568][0] ), .IN0(\CARRYB[567][0] ), .IN1(
        \SUMB[567][1] ), .COUT(\CARRYB[568][0] ), .SUM(PRODUCT[568]) );
  FADDER S2_568_1 ( .CIN(\ab[568][1] ), .IN0(\CARRYB[567][1] ), .IN1(
        \SUMB[567][2] ), .COUT(\CARRYB[568][1] ), .SUM(\SUMB[568][1] ) );
  FADDER S3_568_2 ( .CIN(\ab[568][2] ), .IN0(\CARRYB[567][2] ), .IN1(
        \ab[567][3] ), .COUT(\CARRYB[568][2] ), .SUM(\SUMB[568][2] ) );
  FADDER S1_567_0 ( .CIN(\ab[567][0] ), .IN0(\CARRYB[566][0] ), .IN1(
        \SUMB[566][1] ), .COUT(\CARRYB[567][0] ), .SUM(PRODUCT[567]) );
  FADDER S2_567_1 ( .CIN(\ab[567][1] ), .IN0(\CARRYB[566][1] ), .IN1(
        \SUMB[566][2] ), .COUT(\CARRYB[567][1] ), .SUM(\SUMB[567][1] ) );
  FADDER S3_567_2 ( .CIN(\ab[567][2] ), .IN0(\CARRYB[566][2] ), .IN1(
        \ab[566][3] ), .COUT(\CARRYB[567][2] ), .SUM(\SUMB[567][2] ) );
  FADDER S1_566_0 ( .CIN(\ab[566][0] ), .IN0(\CARRYB[565][0] ), .IN1(
        \SUMB[565][1] ), .COUT(\CARRYB[566][0] ), .SUM(PRODUCT[566]) );
  FADDER S2_566_1 ( .CIN(\ab[566][1] ), .IN0(\CARRYB[565][1] ), .IN1(
        \SUMB[565][2] ), .COUT(\CARRYB[566][1] ), .SUM(\SUMB[566][1] ) );
  FADDER S3_566_2 ( .CIN(\ab[566][2] ), .IN0(\CARRYB[565][2] ), .IN1(
        \ab[565][3] ), .COUT(\CARRYB[566][2] ), .SUM(\SUMB[566][2] ) );
  FADDER S1_565_0 ( .CIN(\ab[565][0] ), .IN0(\CARRYB[564][0] ), .IN1(
        \SUMB[564][1] ), .COUT(\CARRYB[565][0] ), .SUM(PRODUCT[565]) );
  FADDER S2_565_1 ( .CIN(\ab[565][1] ), .IN0(\CARRYB[564][1] ), .IN1(
        \SUMB[564][2] ), .COUT(\CARRYB[565][1] ), .SUM(\SUMB[565][1] ) );
  FADDER S3_565_2 ( .CIN(\ab[565][2] ), .IN0(\CARRYB[564][2] ), .IN1(
        \ab[564][3] ), .COUT(\CARRYB[565][2] ), .SUM(\SUMB[565][2] ) );
  FADDER S1_564_0 ( .CIN(\ab[564][0] ), .IN0(\CARRYB[563][0] ), .IN1(
        \SUMB[563][1] ), .COUT(\CARRYB[564][0] ), .SUM(PRODUCT[564]) );
  FADDER S2_564_1 ( .CIN(\ab[564][1] ), .IN0(\CARRYB[563][1] ), .IN1(
        \SUMB[563][2] ), .COUT(\CARRYB[564][1] ), .SUM(\SUMB[564][1] ) );
  FADDER S3_564_2 ( .CIN(\ab[564][2] ), .IN0(\CARRYB[563][2] ), .IN1(
        \ab[563][3] ), .COUT(\CARRYB[564][2] ), .SUM(\SUMB[564][2] ) );
  FADDER S1_563_0 ( .CIN(\ab[563][0] ), .IN0(\CARRYB[562][0] ), .IN1(
        \SUMB[562][1] ), .COUT(\CARRYB[563][0] ), .SUM(PRODUCT[563]) );
  FADDER S2_563_1 ( .CIN(\ab[563][1] ), .IN0(\CARRYB[562][1] ), .IN1(
        \SUMB[562][2] ), .COUT(\CARRYB[563][1] ), .SUM(\SUMB[563][1] ) );
  FADDER S3_563_2 ( .CIN(\ab[563][2] ), .IN0(\CARRYB[562][2] ), .IN1(
        \ab[562][3] ), .COUT(\CARRYB[563][2] ), .SUM(\SUMB[563][2] ) );
  FADDER S1_562_0 ( .CIN(\ab[562][0] ), .IN0(\CARRYB[561][0] ), .IN1(
        \SUMB[561][1] ), .COUT(\CARRYB[562][0] ), .SUM(PRODUCT[562]) );
  FADDER S2_562_1 ( .CIN(\ab[562][1] ), .IN0(\CARRYB[561][1] ), .IN1(
        \SUMB[561][2] ), .COUT(\CARRYB[562][1] ), .SUM(\SUMB[562][1] ) );
  FADDER S3_562_2 ( .CIN(\ab[562][2] ), .IN0(\CARRYB[561][2] ), .IN1(
        \ab[561][3] ), .COUT(\CARRYB[562][2] ), .SUM(\SUMB[562][2] ) );
  FADDER S1_561_0 ( .CIN(\ab[561][0] ), .IN0(\CARRYB[560][0] ), .IN1(
        \SUMB[560][1] ), .COUT(\CARRYB[561][0] ), .SUM(PRODUCT[561]) );
  FADDER S2_561_1 ( .CIN(\ab[561][1] ), .IN0(\CARRYB[560][1] ), .IN1(
        \SUMB[560][2] ), .COUT(\CARRYB[561][1] ), .SUM(\SUMB[561][1] ) );
  FADDER S3_561_2 ( .CIN(\ab[561][2] ), .IN0(\CARRYB[560][2] ), .IN1(
        \ab[560][3] ), .COUT(\CARRYB[561][2] ), .SUM(\SUMB[561][2] ) );
  FADDER S1_560_0 ( .CIN(\ab[560][0] ), .IN0(\CARRYB[559][0] ), .IN1(
        \SUMB[559][1] ), .COUT(\CARRYB[560][0] ), .SUM(PRODUCT[560]) );
  FADDER S2_560_1 ( .CIN(\ab[560][1] ), .IN0(\CARRYB[559][1] ), .IN1(
        \SUMB[559][2] ), .COUT(\CARRYB[560][1] ), .SUM(\SUMB[560][1] ) );
  FADDER S3_560_2 ( .CIN(\ab[560][2] ), .IN0(\CARRYB[559][2] ), .IN1(
        \ab[559][3] ), .COUT(\CARRYB[560][2] ), .SUM(\SUMB[560][2] ) );
  FADDER S1_559_0 ( .CIN(\ab[559][0] ), .IN0(\CARRYB[558][0] ), .IN1(
        \SUMB[558][1] ), .COUT(\CARRYB[559][0] ), .SUM(PRODUCT[559]) );
  FADDER S2_559_1 ( .CIN(\ab[559][1] ), .IN0(\CARRYB[558][1] ), .IN1(
        \SUMB[558][2] ), .COUT(\CARRYB[559][1] ), .SUM(\SUMB[559][1] ) );
  FADDER S3_559_2 ( .CIN(\ab[559][2] ), .IN0(\CARRYB[558][2] ), .IN1(
        \ab[558][3] ), .COUT(\CARRYB[559][2] ), .SUM(\SUMB[559][2] ) );
  FADDER S1_558_0 ( .CIN(\ab[558][0] ), .IN0(\CARRYB[557][0] ), .IN1(
        \SUMB[557][1] ), .COUT(\CARRYB[558][0] ), .SUM(PRODUCT[558]) );
  FADDER S2_558_1 ( .CIN(\ab[558][1] ), .IN0(\CARRYB[557][1] ), .IN1(
        \SUMB[557][2] ), .COUT(\CARRYB[558][1] ), .SUM(\SUMB[558][1] ) );
  FADDER S3_558_2 ( .CIN(\ab[558][2] ), .IN0(\CARRYB[557][2] ), .IN1(
        \ab[557][3] ), .COUT(\CARRYB[558][2] ), .SUM(\SUMB[558][2] ) );
  FADDER S1_557_0 ( .CIN(\ab[557][0] ), .IN0(\CARRYB[556][0] ), .IN1(
        \SUMB[556][1] ), .COUT(\CARRYB[557][0] ), .SUM(PRODUCT[557]) );
  FADDER S2_557_1 ( .CIN(\ab[557][1] ), .IN0(\CARRYB[556][1] ), .IN1(
        \SUMB[556][2] ), .COUT(\CARRYB[557][1] ), .SUM(\SUMB[557][1] ) );
  FADDER S3_557_2 ( .CIN(\ab[557][2] ), .IN0(\CARRYB[556][2] ), .IN1(
        \ab[556][3] ), .COUT(\CARRYB[557][2] ), .SUM(\SUMB[557][2] ) );
  FADDER S1_556_0 ( .CIN(\ab[556][0] ), .IN0(\CARRYB[555][0] ), .IN1(
        \SUMB[555][1] ), .COUT(\CARRYB[556][0] ), .SUM(PRODUCT[556]) );
  FADDER S2_556_1 ( .CIN(\ab[556][1] ), .IN0(\CARRYB[555][1] ), .IN1(
        \SUMB[555][2] ), .COUT(\CARRYB[556][1] ), .SUM(\SUMB[556][1] ) );
  FADDER S3_556_2 ( .CIN(\ab[556][2] ), .IN0(\CARRYB[555][2] ), .IN1(
        \ab[555][3] ), .COUT(\CARRYB[556][2] ), .SUM(\SUMB[556][2] ) );
  FADDER S1_555_0 ( .CIN(\ab[555][0] ), .IN0(\CARRYB[554][0] ), .IN1(
        \SUMB[554][1] ), .COUT(\CARRYB[555][0] ), .SUM(PRODUCT[555]) );
  FADDER S2_555_1 ( .CIN(\ab[555][1] ), .IN0(\CARRYB[554][1] ), .IN1(
        \SUMB[554][2] ), .COUT(\CARRYB[555][1] ), .SUM(\SUMB[555][1] ) );
  FADDER S3_555_2 ( .CIN(\ab[555][2] ), .IN0(\CARRYB[554][2] ), .IN1(
        \ab[554][3] ), .COUT(\CARRYB[555][2] ), .SUM(\SUMB[555][2] ) );
  FADDER S1_554_0 ( .CIN(\ab[554][0] ), .IN0(\CARRYB[553][0] ), .IN1(
        \SUMB[553][1] ), .COUT(\CARRYB[554][0] ), .SUM(PRODUCT[554]) );
  FADDER S2_554_1 ( .CIN(\ab[554][1] ), .IN0(\CARRYB[553][1] ), .IN1(
        \SUMB[553][2] ), .COUT(\CARRYB[554][1] ), .SUM(\SUMB[554][1] ) );
  FADDER S3_554_2 ( .CIN(\ab[554][2] ), .IN0(\CARRYB[553][2] ), .IN1(
        \ab[553][3] ), .COUT(\CARRYB[554][2] ), .SUM(\SUMB[554][2] ) );
  FADDER S1_553_0 ( .CIN(\ab[553][0] ), .IN0(\CARRYB[552][0] ), .IN1(
        \SUMB[552][1] ), .COUT(\CARRYB[553][0] ), .SUM(PRODUCT[553]) );
  FADDER S2_553_1 ( .CIN(\ab[553][1] ), .IN0(\CARRYB[552][1] ), .IN1(
        \SUMB[552][2] ), .COUT(\CARRYB[553][1] ), .SUM(\SUMB[553][1] ) );
  FADDER S3_553_2 ( .CIN(\ab[553][2] ), .IN0(\CARRYB[552][2] ), .IN1(
        \ab[552][3] ), .COUT(\CARRYB[553][2] ), .SUM(\SUMB[553][2] ) );
  FADDER S1_552_0 ( .CIN(\ab[552][0] ), .IN0(\CARRYB[551][0] ), .IN1(
        \SUMB[551][1] ), .COUT(\CARRYB[552][0] ), .SUM(PRODUCT[552]) );
  FADDER S2_552_1 ( .CIN(\ab[552][1] ), .IN0(\CARRYB[551][1] ), .IN1(
        \SUMB[551][2] ), .COUT(\CARRYB[552][1] ), .SUM(\SUMB[552][1] ) );
  FADDER S3_552_2 ( .CIN(\ab[552][2] ), .IN0(\CARRYB[551][2] ), .IN1(
        \ab[551][3] ), .COUT(\CARRYB[552][2] ), .SUM(\SUMB[552][2] ) );
  FADDER S1_551_0 ( .CIN(\ab[551][0] ), .IN0(\CARRYB[550][0] ), .IN1(
        \SUMB[550][1] ), .COUT(\CARRYB[551][0] ), .SUM(PRODUCT[551]) );
  FADDER S2_551_1 ( .CIN(\ab[551][1] ), .IN0(\CARRYB[550][1] ), .IN1(
        \SUMB[550][2] ), .COUT(\CARRYB[551][1] ), .SUM(\SUMB[551][1] ) );
  FADDER S3_551_2 ( .CIN(\ab[551][2] ), .IN0(\CARRYB[550][2] ), .IN1(
        \ab[550][3] ), .COUT(\CARRYB[551][2] ), .SUM(\SUMB[551][2] ) );
  FADDER S1_550_0 ( .CIN(\ab[550][0] ), .IN0(\CARRYB[549][0] ), .IN1(
        \SUMB[549][1] ), .COUT(\CARRYB[550][0] ), .SUM(PRODUCT[550]) );
  FADDER S2_550_1 ( .CIN(\ab[550][1] ), .IN0(\CARRYB[549][1] ), .IN1(
        \SUMB[549][2] ), .COUT(\CARRYB[550][1] ), .SUM(\SUMB[550][1] ) );
  FADDER S3_550_2 ( .CIN(\ab[550][2] ), .IN0(\CARRYB[549][2] ), .IN1(
        \ab[549][3] ), .COUT(\CARRYB[550][2] ), .SUM(\SUMB[550][2] ) );
  FADDER S1_549_0 ( .CIN(\ab[549][0] ), .IN0(\CARRYB[548][0] ), .IN1(
        \SUMB[548][1] ), .COUT(\CARRYB[549][0] ), .SUM(PRODUCT[549]) );
  FADDER S2_549_1 ( .CIN(\ab[549][1] ), .IN0(\CARRYB[548][1] ), .IN1(
        \SUMB[548][2] ), .COUT(\CARRYB[549][1] ), .SUM(\SUMB[549][1] ) );
  FADDER S3_549_2 ( .CIN(\ab[549][2] ), .IN0(\CARRYB[548][2] ), .IN1(
        \ab[548][3] ), .COUT(\CARRYB[549][2] ), .SUM(\SUMB[549][2] ) );
  FADDER S1_548_0 ( .CIN(\ab[548][0] ), .IN0(\CARRYB[547][0] ), .IN1(
        \SUMB[547][1] ), .COUT(\CARRYB[548][0] ), .SUM(PRODUCT[548]) );
  FADDER S2_548_1 ( .CIN(\ab[548][1] ), .IN0(\CARRYB[547][1] ), .IN1(
        \SUMB[547][2] ), .COUT(\CARRYB[548][1] ), .SUM(\SUMB[548][1] ) );
  FADDER S3_548_2 ( .CIN(\ab[548][2] ), .IN0(\CARRYB[547][2] ), .IN1(
        \ab[547][3] ), .COUT(\CARRYB[548][2] ), .SUM(\SUMB[548][2] ) );
  FADDER S1_547_0 ( .CIN(\ab[547][0] ), .IN0(\CARRYB[546][0] ), .IN1(
        \SUMB[546][1] ), .COUT(\CARRYB[547][0] ), .SUM(PRODUCT[547]) );
  FADDER S2_547_1 ( .CIN(\ab[547][1] ), .IN0(\CARRYB[546][1] ), .IN1(
        \SUMB[546][2] ), .COUT(\CARRYB[547][1] ), .SUM(\SUMB[547][1] ) );
  FADDER S3_547_2 ( .CIN(\ab[547][2] ), .IN0(\CARRYB[546][2] ), .IN1(
        \ab[546][3] ), .COUT(\CARRYB[547][2] ), .SUM(\SUMB[547][2] ) );
  FADDER S1_546_0 ( .CIN(\ab[546][0] ), .IN0(\CARRYB[545][0] ), .IN1(
        \SUMB[545][1] ), .COUT(\CARRYB[546][0] ), .SUM(PRODUCT[546]) );
  FADDER S2_546_1 ( .CIN(\ab[546][1] ), .IN0(\CARRYB[545][1] ), .IN1(
        \SUMB[545][2] ), .COUT(\CARRYB[546][1] ), .SUM(\SUMB[546][1] ) );
  FADDER S3_546_2 ( .CIN(\ab[546][2] ), .IN0(\CARRYB[545][2] ), .IN1(
        \ab[545][3] ), .COUT(\CARRYB[546][2] ), .SUM(\SUMB[546][2] ) );
  FADDER S1_545_0 ( .CIN(\ab[545][0] ), .IN0(\CARRYB[544][0] ), .IN1(
        \SUMB[544][1] ), .COUT(\CARRYB[545][0] ), .SUM(PRODUCT[545]) );
  FADDER S2_545_1 ( .CIN(\ab[545][1] ), .IN0(\CARRYB[544][1] ), .IN1(
        \SUMB[544][2] ), .COUT(\CARRYB[545][1] ), .SUM(\SUMB[545][1] ) );
  FADDER S3_545_2 ( .CIN(\ab[545][2] ), .IN0(\CARRYB[544][2] ), .IN1(
        \ab[544][3] ), .COUT(\CARRYB[545][2] ), .SUM(\SUMB[545][2] ) );
  FADDER S1_544_0 ( .CIN(\ab[544][0] ), .IN0(\CARRYB[543][0] ), .IN1(
        \SUMB[543][1] ), .COUT(\CARRYB[544][0] ), .SUM(PRODUCT[544]) );
  FADDER S2_544_1 ( .CIN(\ab[544][1] ), .IN0(\CARRYB[543][1] ), .IN1(
        \SUMB[543][2] ), .COUT(\CARRYB[544][1] ), .SUM(\SUMB[544][1] ) );
  FADDER S3_544_2 ( .CIN(\ab[544][2] ), .IN0(\CARRYB[543][2] ), .IN1(
        \ab[543][3] ), .COUT(\CARRYB[544][2] ), .SUM(\SUMB[544][2] ) );
  FADDER S1_543_0 ( .CIN(\ab[543][0] ), .IN0(\CARRYB[542][0] ), .IN1(
        \SUMB[542][1] ), .COUT(\CARRYB[543][0] ), .SUM(PRODUCT[543]) );
  FADDER S2_543_1 ( .CIN(\ab[543][1] ), .IN0(\CARRYB[542][1] ), .IN1(
        \SUMB[542][2] ), .COUT(\CARRYB[543][1] ), .SUM(\SUMB[543][1] ) );
  FADDER S3_543_2 ( .CIN(\ab[543][2] ), .IN0(\CARRYB[542][2] ), .IN1(
        \ab[542][3] ), .COUT(\CARRYB[543][2] ), .SUM(\SUMB[543][2] ) );
  FADDER S1_542_0 ( .CIN(\ab[542][0] ), .IN0(\CARRYB[541][0] ), .IN1(
        \SUMB[541][1] ), .COUT(\CARRYB[542][0] ), .SUM(PRODUCT[542]) );
  FADDER S2_542_1 ( .CIN(\ab[542][1] ), .IN0(\CARRYB[541][1] ), .IN1(
        \SUMB[541][2] ), .COUT(\CARRYB[542][1] ), .SUM(\SUMB[542][1] ) );
  FADDER S3_542_2 ( .CIN(\ab[542][2] ), .IN0(\CARRYB[541][2] ), .IN1(
        \ab[541][3] ), .COUT(\CARRYB[542][2] ), .SUM(\SUMB[542][2] ) );
  FADDER S1_541_0 ( .CIN(\ab[541][0] ), .IN0(\CARRYB[540][0] ), .IN1(
        \SUMB[540][1] ), .COUT(\CARRYB[541][0] ), .SUM(PRODUCT[541]) );
  FADDER S2_541_1 ( .CIN(\ab[541][1] ), .IN0(\CARRYB[540][1] ), .IN1(
        \SUMB[540][2] ), .COUT(\CARRYB[541][1] ), .SUM(\SUMB[541][1] ) );
  FADDER S3_541_2 ( .CIN(\ab[541][2] ), .IN0(\CARRYB[540][2] ), .IN1(
        \ab[540][3] ), .COUT(\CARRYB[541][2] ), .SUM(\SUMB[541][2] ) );
  FADDER S1_540_0 ( .CIN(\ab[540][0] ), .IN0(\CARRYB[539][0] ), .IN1(
        \SUMB[539][1] ), .COUT(\CARRYB[540][0] ), .SUM(PRODUCT[540]) );
  FADDER S2_540_1 ( .CIN(\ab[540][1] ), .IN0(\CARRYB[539][1] ), .IN1(
        \SUMB[539][2] ), .COUT(\CARRYB[540][1] ), .SUM(\SUMB[540][1] ) );
  FADDER S3_540_2 ( .CIN(\ab[540][2] ), .IN0(\CARRYB[539][2] ), .IN1(
        \ab[539][3] ), .COUT(\CARRYB[540][2] ), .SUM(\SUMB[540][2] ) );
  FADDER S1_539_0 ( .CIN(\ab[539][0] ), .IN0(\CARRYB[538][0] ), .IN1(
        \SUMB[538][1] ), .COUT(\CARRYB[539][0] ), .SUM(PRODUCT[539]) );
  FADDER S2_539_1 ( .CIN(\ab[539][1] ), .IN0(\CARRYB[538][1] ), .IN1(
        \SUMB[538][2] ), .COUT(\CARRYB[539][1] ), .SUM(\SUMB[539][1] ) );
  FADDER S3_539_2 ( .CIN(\ab[539][2] ), .IN0(\CARRYB[538][2] ), .IN1(
        \ab[538][3] ), .COUT(\CARRYB[539][2] ), .SUM(\SUMB[539][2] ) );
  FADDER S1_538_0 ( .CIN(\ab[538][0] ), .IN0(\CARRYB[537][0] ), .IN1(
        \SUMB[537][1] ), .COUT(\CARRYB[538][0] ), .SUM(PRODUCT[538]) );
  FADDER S2_538_1 ( .CIN(\ab[538][1] ), .IN0(\CARRYB[537][1] ), .IN1(
        \SUMB[537][2] ), .COUT(\CARRYB[538][1] ), .SUM(\SUMB[538][1] ) );
  FADDER S3_538_2 ( .CIN(\ab[538][2] ), .IN0(\CARRYB[537][2] ), .IN1(
        \ab[537][3] ), .COUT(\CARRYB[538][2] ), .SUM(\SUMB[538][2] ) );
  FADDER S1_537_0 ( .CIN(\ab[537][0] ), .IN0(\CARRYB[536][0] ), .IN1(
        \SUMB[536][1] ), .COUT(\CARRYB[537][0] ), .SUM(PRODUCT[537]) );
  FADDER S2_537_1 ( .CIN(\ab[537][1] ), .IN0(\CARRYB[536][1] ), .IN1(
        \SUMB[536][2] ), .COUT(\CARRYB[537][1] ), .SUM(\SUMB[537][1] ) );
  FADDER S3_537_2 ( .CIN(\ab[537][2] ), .IN0(\CARRYB[536][2] ), .IN1(
        \ab[536][3] ), .COUT(\CARRYB[537][2] ), .SUM(\SUMB[537][2] ) );
  FADDER S1_536_0 ( .CIN(\ab[536][0] ), .IN0(\CARRYB[535][0] ), .IN1(
        \SUMB[535][1] ), .COUT(\CARRYB[536][0] ), .SUM(PRODUCT[536]) );
  FADDER S2_536_1 ( .CIN(\ab[536][1] ), .IN0(\CARRYB[535][1] ), .IN1(
        \SUMB[535][2] ), .COUT(\CARRYB[536][1] ), .SUM(\SUMB[536][1] ) );
  FADDER S3_536_2 ( .CIN(\ab[536][2] ), .IN0(\CARRYB[535][2] ), .IN1(
        \ab[535][3] ), .COUT(\CARRYB[536][2] ), .SUM(\SUMB[536][2] ) );
  FADDER S1_535_0 ( .CIN(\ab[535][0] ), .IN0(\CARRYB[534][0] ), .IN1(
        \SUMB[534][1] ), .COUT(\CARRYB[535][0] ), .SUM(PRODUCT[535]) );
  FADDER S2_535_1 ( .CIN(\ab[535][1] ), .IN0(\CARRYB[534][1] ), .IN1(
        \SUMB[534][2] ), .COUT(\CARRYB[535][1] ), .SUM(\SUMB[535][1] ) );
  FADDER S3_535_2 ( .CIN(\ab[535][2] ), .IN0(\CARRYB[534][2] ), .IN1(
        \ab[534][3] ), .COUT(\CARRYB[535][2] ), .SUM(\SUMB[535][2] ) );
  FADDER S1_534_0 ( .CIN(\ab[534][0] ), .IN0(\CARRYB[533][0] ), .IN1(
        \SUMB[533][1] ), .COUT(\CARRYB[534][0] ), .SUM(PRODUCT[534]) );
  FADDER S2_534_1 ( .CIN(\ab[534][1] ), .IN0(\CARRYB[533][1] ), .IN1(
        \SUMB[533][2] ), .COUT(\CARRYB[534][1] ), .SUM(\SUMB[534][1] ) );
  FADDER S3_534_2 ( .CIN(\ab[534][2] ), .IN0(\CARRYB[533][2] ), .IN1(
        \ab[533][3] ), .COUT(\CARRYB[534][2] ), .SUM(\SUMB[534][2] ) );
  FADDER S1_533_0 ( .CIN(\ab[533][0] ), .IN0(\CARRYB[532][0] ), .IN1(
        \SUMB[532][1] ), .COUT(\CARRYB[533][0] ), .SUM(PRODUCT[533]) );
  FADDER S2_533_1 ( .CIN(\ab[533][1] ), .IN0(\CARRYB[532][1] ), .IN1(
        \SUMB[532][2] ), .COUT(\CARRYB[533][1] ), .SUM(\SUMB[533][1] ) );
  FADDER S3_533_2 ( .CIN(\ab[533][2] ), .IN0(\CARRYB[532][2] ), .IN1(
        \ab[532][3] ), .COUT(\CARRYB[533][2] ), .SUM(\SUMB[533][2] ) );
  FADDER S1_532_0 ( .CIN(\ab[532][0] ), .IN0(\CARRYB[531][0] ), .IN1(
        \SUMB[531][1] ), .COUT(\CARRYB[532][0] ), .SUM(PRODUCT[532]) );
  FADDER S2_532_1 ( .CIN(\ab[532][1] ), .IN0(\CARRYB[531][1] ), .IN1(
        \SUMB[531][2] ), .COUT(\CARRYB[532][1] ), .SUM(\SUMB[532][1] ) );
  FADDER S3_532_2 ( .CIN(\ab[532][2] ), .IN0(\CARRYB[531][2] ), .IN1(
        \ab[531][3] ), .COUT(\CARRYB[532][2] ), .SUM(\SUMB[532][2] ) );
  FADDER S1_531_0 ( .CIN(\ab[531][0] ), .IN0(\CARRYB[530][0] ), .IN1(
        \SUMB[530][1] ), .COUT(\CARRYB[531][0] ), .SUM(PRODUCT[531]) );
  FADDER S2_531_1 ( .CIN(\ab[531][1] ), .IN0(\CARRYB[530][1] ), .IN1(
        \SUMB[530][2] ), .COUT(\CARRYB[531][1] ), .SUM(\SUMB[531][1] ) );
  FADDER S3_531_2 ( .CIN(\ab[531][2] ), .IN0(\CARRYB[530][2] ), .IN1(
        \ab[530][3] ), .COUT(\CARRYB[531][2] ), .SUM(\SUMB[531][2] ) );
  FADDER S1_530_0 ( .CIN(\ab[530][0] ), .IN0(\CARRYB[529][0] ), .IN1(
        \SUMB[529][1] ), .COUT(\CARRYB[530][0] ), .SUM(PRODUCT[530]) );
  FADDER S2_530_1 ( .CIN(\ab[530][1] ), .IN0(\CARRYB[529][1] ), .IN1(
        \SUMB[529][2] ), .COUT(\CARRYB[530][1] ), .SUM(\SUMB[530][1] ) );
  FADDER S3_530_2 ( .CIN(\ab[530][2] ), .IN0(\CARRYB[529][2] ), .IN1(
        \ab[529][3] ), .COUT(\CARRYB[530][2] ), .SUM(\SUMB[530][2] ) );
  FADDER S1_529_0 ( .CIN(\ab[529][0] ), .IN0(\CARRYB[528][0] ), .IN1(
        \SUMB[528][1] ), .COUT(\CARRYB[529][0] ), .SUM(PRODUCT[529]) );
  FADDER S2_529_1 ( .CIN(\ab[529][1] ), .IN0(\CARRYB[528][1] ), .IN1(
        \SUMB[528][2] ), .COUT(\CARRYB[529][1] ), .SUM(\SUMB[529][1] ) );
  FADDER S3_529_2 ( .CIN(\ab[529][2] ), .IN0(\CARRYB[528][2] ), .IN1(
        \ab[528][3] ), .COUT(\CARRYB[529][2] ), .SUM(\SUMB[529][2] ) );
  FADDER S1_528_0 ( .CIN(\ab[528][0] ), .IN0(\CARRYB[527][0] ), .IN1(
        \SUMB[527][1] ), .COUT(\CARRYB[528][0] ), .SUM(PRODUCT[528]) );
  FADDER S2_528_1 ( .CIN(\ab[528][1] ), .IN0(\CARRYB[527][1] ), .IN1(
        \SUMB[527][2] ), .COUT(\CARRYB[528][1] ), .SUM(\SUMB[528][1] ) );
  FADDER S3_528_2 ( .CIN(\ab[528][2] ), .IN0(\CARRYB[527][2] ), .IN1(
        \ab[527][3] ), .COUT(\CARRYB[528][2] ), .SUM(\SUMB[528][2] ) );
  FADDER S1_527_0 ( .CIN(\ab[527][0] ), .IN0(\CARRYB[526][0] ), .IN1(
        \SUMB[526][1] ), .COUT(\CARRYB[527][0] ), .SUM(PRODUCT[527]) );
  FADDER S2_527_1 ( .CIN(\ab[527][1] ), .IN0(\CARRYB[526][1] ), .IN1(
        \SUMB[526][2] ), .COUT(\CARRYB[527][1] ), .SUM(\SUMB[527][1] ) );
  FADDER S3_527_2 ( .CIN(\ab[527][2] ), .IN0(\CARRYB[526][2] ), .IN1(
        \ab[526][3] ), .COUT(\CARRYB[527][2] ), .SUM(\SUMB[527][2] ) );
  FADDER S1_526_0 ( .CIN(\ab[526][0] ), .IN0(\CARRYB[525][0] ), .IN1(
        \SUMB[525][1] ), .COUT(\CARRYB[526][0] ), .SUM(PRODUCT[526]) );
  FADDER S2_526_1 ( .CIN(\ab[526][1] ), .IN0(\CARRYB[525][1] ), .IN1(
        \SUMB[525][2] ), .COUT(\CARRYB[526][1] ), .SUM(\SUMB[526][1] ) );
  FADDER S3_526_2 ( .CIN(\ab[526][2] ), .IN0(\CARRYB[525][2] ), .IN1(
        \ab[525][3] ), .COUT(\CARRYB[526][2] ), .SUM(\SUMB[526][2] ) );
  FADDER S1_525_0 ( .CIN(\ab[525][0] ), .IN0(\CARRYB[524][0] ), .IN1(
        \SUMB[524][1] ), .COUT(\CARRYB[525][0] ), .SUM(PRODUCT[525]) );
  FADDER S2_525_1 ( .CIN(\ab[525][1] ), .IN0(\CARRYB[524][1] ), .IN1(
        \SUMB[524][2] ), .COUT(\CARRYB[525][1] ), .SUM(\SUMB[525][1] ) );
  FADDER S3_525_2 ( .CIN(\ab[525][2] ), .IN0(\CARRYB[524][2] ), .IN1(
        \ab[524][3] ), .COUT(\CARRYB[525][2] ), .SUM(\SUMB[525][2] ) );
  FADDER S1_524_0 ( .CIN(\ab[524][0] ), .IN0(\CARRYB[523][0] ), .IN1(
        \SUMB[523][1] ), .COUT(\CARRYB[524][0] ), .SUM(PRODUCT[524]) );
  FADDER S2_524_1 ( .CIN(\ab[524][1] ), .IN0(\CARRYB[523][1] ), .IN1(
        \SUMB[523][2] ), .COUT(\CARRYB[524][1] ), .SUM(\SUMB[524][1] ) );
  FADDER S3_524_2 ( .CIN(\ab[524][2] ), .IN0(\CARRYB[523][2] ), .IN1(
        \ab[523][3] ), .COUT(\CARRYB[524][2] ), .SUM(\SUMB[524][2] ) );
  FADDER S1_523_0 ( .CIN(\ab[523][0] ), .IN0(\CARRYB[522][0] ), .IN1(
        \SUMB[522][1] ), .COUT(\CARRYB[523][0] ), .SUM(PRODUCT[523]) );
  FADDER S2_523_1 ( .CIN(\ab[523][1] ), .IN0(\CARRYB[522][1] ), .IN1(
        \SUMB[522][2] ), .COUT(\CARRYB[523][1] ), .SUM(\SUMB[523][1] ) );
  FADDER S3_523_2 ( .CIN(\ab[523][2] ), .IN0(\CARRYB[522][2] ), .IN1(
        \ab[522][3] ), .COUT(\CARRYB[523][2] ), .SUM(\SUMB[523][2] ) );
  FADDER S1_522_0 ( .CIN(\ab[522][0] ), .IN0(\CARRYB[521][0] ), .IN1(
        \SUMB[521][1] ), .COUT(\CARRYB[522][0] ), .SUM(PRODUCT[522]) );
  FADDER S2_522_1 ( .CIN(\ab[522][1] ), .IN0(\CARRYB[521][1] ), .IN1(
        \SUMB[521][2] ), .COUT(\CARRYB[522][1] ), .SUM(\SUMB[522][1] ) );
  FADDER S3_522_2 ( .CIN(\ab[522][2] ), .IN0(\CARRYB[521][2] ), .IN1(
        \ab[521][3] ), .COUT(\CARRYB[522][2] ), .SUM(\SUMB[522][2] ) );
  FADDER S1_521_0 ( .CIN(\ab[521][0] ), .IN0(\CARRYB[520][0] ), .IN1(
        \SUMB[520][1] ), .COUT(\CARRYB[521][0] ), .SUM(PRODUCT[521]) );
  FADDER S2_521_1 ( .CIN(\ab[521][1] ), .IN0(\CARRYB[520][1] ), .IN1(
        \SUMB[520][2] ), .COUT(\CARRYB[521][1] ), .SUM(\SUMB[521][1] ) );
  FADDER S3_521_2 ( .CIN(\ab[521][2] ), .IN0(\CARRYB[520][2] ), .IN1(
        \ab[520][3] ), .COUT(\CARRYB[521][2] ), .SUM(\SUMB[521][2] ) );
  FADDER S1_520_0 ( .CIN(\ab[520][0] ), .IN0(\CARRYB[519][0] ), .IN1(
        \SUMB[519][1] ), .COUT(\CARRYB[520][0] ), .SUM(PRODUCT[520]) );
  FADDER S2_520_1 ( .CIN(\ab[520][1] ), .IN0(\CARRYB[519][1] ), .IN1(
        \SUMB[519][2] ), .COUT(\CARRYB[520][1] ), .SUM(\SUMB[520][1] ) );
  FADDER S3_520_2 ( .CIN(\ab[520][2] ), .IN0(\CARRYB[519][2] ), .IN1(
        \ab[519][3] ), .COUT(\CARRYB[520][2] ), .SUM(\SUMB[520][2] ) );
  FADDER S1_519_0 ( .CIN(\ab[519][0] ), .IN0(\CARRYB[518][0] ), .IN1(
        \SUMB[518][1] ), .COUT(\CARRYB[519][0] ), .SUM(PRODUCT[519]) );
  FADDER S2_519_1 ( .CIN(\ab[519][1] ), .IN0(\CARRYB[518][1] ), .IN1(
        \SUMB[518][2] ), .COUT(\CARRYB[519][1] ), .SUM(\SUMB[519][1] ) );
  FADDER S3_519_2 ( .CIN(\ab[519][2] ), .IN0(\CARRYB[518][2] ), .IN1(
        \ab[518][3] ), .COUT(\CARRYB[519][2] ), .SUM(\SUMB[519][2] ) );
  FADDER S1_518_0 ( .CIN(\ab[518][0] ), .IN0(\CARRYB[517][0] ), .IN1(
        \SUMB[517][1] ), .COUT(\CARRYB[518][0] ), .SUM(PRODUCT[518]) );
  FADDER S2_518_1 ( .CIN(\ab[518][1] ), .IN0(\CARRYB[517][1] ), .IN1(
        \SUMB[517][2] ), .COUT(\CARRYB[518][1] ), .SUM(\SUMB[518][1] ) );
  FADDER S3_518_2 ( .CIN(\ab[518][2] ), .IN0(\CARRYB[517][2] ), .IN1(
        \ab[517][3] ), .COUT(\CARRYB[518][2] ), .SUM(\SUMB[518][2] ) );
  FADDER S1_517_0 ( .CIN(\ab[517][0] ), .IN0(\CARRYB[516][0] ), .IN1(
        \SUMB[516][1] ), .COUT(\CARRYB[517][0] ), .SUM(PRODUCT[517]) );
  FADDER S2_517_1 ( .CIN(\ab[517][1] ), .IN0(\CARRYB[516][1] ), .IN1(
        \SUMB[516][2] ), .COUT(\CARRYB[517][1] ), .SUM(\SUMB[517][1] ) );
  FADDER S3_517_2 ( .CIN(\ab[517][2] ), .IN0(\CARRYB[516][2] ), .IN1(
        \ab[516][3] ), .COUT(\CARRYB[517][2] ), .SUM(\SUMB[517][2] ) );
  FADDER S1_516_0 ( .CIN(\ab[516][0] ), .IN0(\CARRYB[515][0] ), .IN1(
        \SUMB[515][1] ), .COUT(\CARRYB[516][0] ), .SUM(PRODUCT[516]) );
  FADDER S2_516_1 ( .CIN(\ab[516][1] ), .IN0(\CARRYB[515][1] ), .IN1(
        \SUMB[515][2] ), .COUT(\CARRYB[516][1] ), .SUM(\SUMB[516][1] ) );
  FADDER S3_516_2 ( .CIN(\ab[516][2] ), .IN0(\CARRYB[515][2] ), .IN1(
        \ab[515][3] ), .COUT(\CARRYB[516][2] ), .SUM(\SUMB[516][2] ) );
  FADDER S1_515_0 ( .CIN(\ab[515][0] ), .IN0(\CARRYB[514][0] ), .IN1(
        \SUMB[514][1] ), .COUT(\CARRYB[515][0] ), .SUM(PRODUCT[515]) );
  FADDER S2_515_1 ( .CIN(\ab[515][1] ), .IN0(\CARRYB[514][1] ), .IN1(
        \SUMB[514][2] ), .COUT(\CARRYB[515][1] ), .SUM(\SUMB[515][1] ) );
  FADDER S3_515_2 ( .CIN(\ab[515][2] ), .IN0(\CARRYB[514][2] ), .IN1(
        \ab[514][3] ), .COUT(\CARRYB[515][2] ), .SUM(\SUMB[515][2] ) );
  FADDER S1_514_0 ( .CIN(\ab[514][0] ), .IN0(\CARRYB[513][0] ), .IN1(
        \SUMB[513][1] ), .COUT(\CARRYB[514][0] ), .SUM(PRODUCT[514]) );
  FADDER S2_514_1 ( .CIN(\ab[514][1] ), .IN0(\CARRYB[513][1] ), .IN1(
        \SUMB[513][2] ), .COUT(\CARRYB[514][1] ), .SUM(\SUMB[514][1] ) );
  FADDER S3_514_2 ( .CIN(\ab[514][2] ), .IN0(\CARRYB[513][2] ), .IN1(
        \ab[513][3] ), .COUT(\CARRYB[514][2] ), .SUM(\SUMB[514][2] ) );
  FADDER S1_513_0 ( .CIN(\ab[513][0] ), .IN0(\CARRYB[512][0] ), .IN1(
        \SUMB[512][1] ), .COUT(\CARRYB[513][0] ), .SUM(PRODUCT[513]) );
  FADDER S2_513_1 ( .CIN(\ab[513][1] ), .IN0(\CARRYB[512][1] ), .IN1(
        \SUMB[512][2] ), .COUT(\CARRYB[513][1] ), .SUM(\SUMB[513][1] ) );
  FADDER S3_513_2 ( .CIN(\ab[513][2] ), .IN0(\CARRYB[512][2] ), .IN1(
        \ab[512][3] ), .COUT(\CARRYB[513][2] ), .SUM(\SUMB[513][2] ) );
  FADDER S1_512_0 ( .CIN(\ab[512][0] ), .IN0(\CARRYB[511][0] ), .IN1(
        \SUMB[511][1] ), .COUT(\CARRYB[512][0] ), .SUM(PRODUCT[512]) );
  FADDER S2_512_1 ( .CIN(\ab[512][1] ), .IN0(\CARRYB[511][1] ), .IN1(
        \SUMB[511][2] ), .COUT(\CARRYB[512][1] ), .SUM(\SUMB[512][1] ) );
  FADDER S3_512_2 ( .CIN(\ab[512][2] ), .IN0(\CARRYB[511][2] ), .IN1(
        \ab[511][3] ), .COUT(\CARRYB[512][2] ), .SUM(\SUMB[512][2] ) );
  FADDER S1_511_0 ( .CIN(\ab[511][0] ), .IN0(\CARRYB[510][0] ), .IN1(
        \SUMB[510][1] ), .COUT(\CARRYB[511][0] ), .SUM(PRODUCT[511]) );
  FADDER S2_511_1 ( .CIN(\ab[511][1] ), .IN0(\CARRYB[510][1] ), .IN1(
        \SUMB[510][2] ), .COUT(\CARRYB[511][1] ), .SUM(\SUMB[511][1] ) );
  FADDER S3_511_2 ( .CIN(\ab[511][2] ), .IN0(\CARRYB[510][2] ), .IN1(
        \ab[510][3] ), .COUT(\CARRYB[511][2] ), .SUM(\SUMB[511][2] ) );
  FADDER S1_510_0 ( .CIN(\ab[510][0] ), .IN0(\CARRYB[509][0] ), .IN1(
        \SUMB[509][1] ), .COUT(\CARRYB[510][0] ), .SUM(PRODUCT[510]) );
  FADDER S2_510_1 ( .CIN(\ab[510][1] ), .IN0(\CARRYB[509][1] ), .IN1(
        \SUMB[509][2] ), .COUT(\CARRYB[510][1] ), .SUM(\SUMB[510][1] ) );
  FADDER S3_510_2 ( .CIN(\ab[510][2] ), .IN0(\CARRYB[509][2] ), .IN1(
        \ab[509][3] ), .COUT(\CARRYB[510][2] ), .SUM(\SUMB[510][2] ) );
  FADDER S1_509_0 ( .CIN(\ab[509][0] ), .IN0(\CARRYB[508][0] ), .IN1(
        \SUMB[508][1] ), .COUT(\CARRYB[509][0] ), .SUM(PRODUCT[509]) );
  FADDER S2_509_1 ( .CIN(\ab[509][1] ), .IN0(\CARRYB[508][1] ), .IN1(
        \SUMB[508][2] ), .COUT(\CARRYB[509][1] ), .SUM(\SUMB[509][1] ) );
  FADDER S3_509_2 ( .CIN(\ab[509][2] ), .IN0(\CARRYB[508][2] ), .IN1(
        \ab[508][3] ), .COUT(\CARRYB[509][2] ), .SUM(\SUMB[509][2] ) );
  FADDER S1_508_0 ( .CIN(\ab[508][0] ), .IN0(\CARRYB[507][0] ), .IN1(
        \SUMB[507][1] ), .COUT(\CARRYB[508][0] ), .SUM(PRODUCT[508]) );
  FADDER S2_508_1 ( .CIN(\ab[508][1] ), .IN0(\CARRYB[507][1] ), .IN1(
        \SUMB[507][2] ), .COUT(\CARRYB[508][1] ), .SUM(\SUMB[508][1] ) );
  FADDER S3_508_2 ( .CIN(\ab[508][2] ), .IN0(\CARRYB[507][2] ), .IN1(
        \ab[507][3] ), .COUT(\CARRYB[508][2] ), .SUM(\SUMB[508][2] ) );
  FADDER S1_507_0 ( .CIN(\ab[507][0] ), .IN0(\CARRYB[506][0] ), .IN1(
        \SUMB[506][1] ), .COUT(\CARRYB[507][0] ), .SUM(PRODUCT[507]) );
  FADDER S2_507_1 ( .CIN(\ab[507][1] ), .IN0(\CARRYB[506][1] ), .IN1(
        \SUMB[506][2] ), .COUT(\CARRYB[507][1] ), .SUM(\SUMB[507][1] ) );
  FADDER S3_507_2 ( .CIN(\ab[507][2] ), .IN0(\CARRYB[506][2] ), .IN1(
        \ab[506][3] ), .COUT(\CARRYB[507][2] ), .SUM(\SUMB[507][2] ) );
  FADDER S1_506_0 ( .CIN(\ab[506][0] ), .IN0(\CARRYB[505][0] ), .IN1(
        \SUMB[505][1] ), .COUT(\CARRYB[506][0] ), .SUM(PRODUCT[506]) );
  FADDER S2_506_1 ( .CIN(\ab[506][1] ), .IN0(\CARRYB[505][1] ), .IN1(
        \SUMB[505][2] ), .COUT(\CARRYB[506][1] ), .SUM(\SUMB[506][1] ) );
  FADDER S3_506_2 ( .CIN(\ab[506][2] ), .IN0(\CARRYB[505][2] ), .IN1(
        \ab[505][3] ), .COUT(\CARRYB[506][2] ), .SUM(\SUMB[506][2] ) );
  FADDER S1_505_0 ( .CIN(\ab[505][0] ), .IN0(\CARRYB[504][0] ), .IN1(
        \SUMB[504][1] ), .COUT(\CARRYB[505][0] ), .SUM(PRODUCT[505]) );
  FADDER S2_505_1 ( .CIN(\ab[505][1] ), .IN0(\CARRYB[504][1] ), .IN1(
        \SUMB[504][2] ), .COUT(\CARRYB[505][1] ), .SUM(\SUMB[505][1] ) );
  FADDER S3_505_2 ( .CIN(\ab[505][2] ), .IN0(\CARRYB[504][2] ), .IN1(
        \ab[504][3] ), .COUT(\CARRYB[505][2] ), .SUM(\SUMB[505][2] ) );
  FADDER S1_504_0 ( .CIN(\ab[504][0] ), .IN0(\CARRYB[503][0] ), .IN1(
        \SUMB[503][1] ), .COUT(\CARRYB[504][0] ), .SUM(PRODUCT[504]) );
  FADDER S2_504_1 ( .CIN(\ab[504][1] ), .IN0(\CARRYB[503][1] ), .IN1(
        \SUMB[503][2] ), .COUT(\CARRYB[504][1] ), .SUM(\SUMB[504][1] ) );
  FADDER S3_504_2 ( .CIN(\ab[504][2] ), .IN0(\CARRYB[503][2] ), .IN1(
        \ab[503][3] ), .COUT(\CARRYB[504][2] ), .SUM(\SUMB[504][2] ) );
  FADDER S1_503_0 ( .CIN(\ab[503][0] ), .IN0(\CARRYB[502][0] ), .IN1(
        \SUMB[502][1] ), .COUT(\CARRYB[503][0] ), .SUM(PRODUCT[503]) );
  FADDER S2_503_1 ( .CIN(\ab[503][1] ), .IN0(\CARRYB[502][1] ), .IN1(
        \SUMB[502][2] ), .COUT(\CARRYB[503][1] ), .SUM(\SUMB[503][1] ) );
  FADDER S3_503_2 ( .CIN(\ab[503][2] ), .IN0(\CARRYB[502][2] ), .IN1(
        \ab[502][3] ), .COUT(\CARRYB[503][2] ), .SUM(\SUMB[503][2] ) );
  FADDER S1_502_0 ( .CIN(\ab[502][0] ), .IN0(\CARRYB[501][0] ), .IN1(
        \SUMB[501][1] ), .COUT(\CARRYB[502][0] ), .SUM(PRODUCT[502]) );
  FADDER S2_502_1 ( .CIN(\ab[502][1] ), .IN0(\CARRYB[501][1] ), .IN1(
        \SUMB[501][2] ), .COUT(\CARRYB[502][1] ), .SUM(\SUMB[502][1] ) );
  FADDER S3_502_2 ( .CIN(\ab[502][2] ), .IN0(\CARRYB[501][2] ), .IN1(
        \ab[501][3] ), .COUT(\CARRYB[502][2] ), .SUM(\SUMB[502][2] ) );
  FADDER S1_501_0 ( .CIN(\ab[501][0] ), .IN0(\CARRYB[500][0] ), .IN1(
        \SUMB[500][1] ), .COUT(\CARRYB[501][0] ), .SUM(PRODUCT[501]) );
  FADDER S2_501_1 ( .CIN(\ab[501][1] ), .IN0(\CARRYB[500][1] ), .IN1(
        \SUMB[500][2] ), .COUT(\CARRYB[501][1] ), .SUM(\SUMB[501][1] ) );
  FADDER S3_501_2 ( .CIN(\ab[501][2] ), .IN0(\CARRYB[500][2] ), .IN1(
        \ab[500][3] ), .COUT(\CARRYB[501][2] ), .SUM(\SUMB[501][2] ) );
  FADDER S1_500_0 ( .CIN(\ab[500][0] ), .IN0(\CARRYB[499][0] ), .IN1(
        \SUMB[499][1] ), .COUT(\CARRYB[500][0] ), .SUM(PRODUCT[500]) );
  FADDER S2_500_1 ( .CIN(\ab[500][1] ), .IN0(\CARRYB[499][1] ), .IN1(
        \SUMB[499][2] ), .COUT(\CARRYB[500][1] ), .SUM(\SUMB[500][1] ) );
  FADDER S3_500_2 ( .CIN(\ab[500][2] ), .IN0(\CARRYB[499][2] ), .IN1(
        \ab[499][3] ), .COUT(\CARRYB[500][2] ), .SUM(\SUMB[500][2] ) );
  FADDER S1_499_0 ( .CIN(\ab[499][0] ), .IN0(\CARRYB[498][0] ), .IN1(
        \SUMB[498][1] ), .COUT(\CARRYB[499][0] ), .SUM(PRODUCT[499]) );
  FADDER S2_499_1 ( .CIN(\ab[499][1] ), .IN0(\CARRYB[498][1] ), .IN1(
        \SUMB[498][2] ), .COUT(\CARRYB[499][1] ), .SUM(\SUMB[499][1] ) );
  FADDER S3_499_2 ( .CIN(\ab[499][2] ), .IN0(\CARRYB[498][2] ), .IN1(
        \ab[498][3] ), .COUT(\CARRYB[499][2] ), .SUM(\SUMB[499][2] ) );
  FADDER S1_498_0 ( .CIN(\ab[498][0] ), .IN0(\CARRYB[497][0] ), .IN1(
        \SUMB[497][1] ), .COUT(\CARRYB[498][0] ), .SUM(PRODUCT[498]) );
  FADDER S2_498_1 ( .CIN(\ab[498][1] ), .IN0(\CARRYB[497][1] ), .IN1(
        \SUMB[497][2] ), .COUT(\CARRYB[498][1] ), .SUM(\SUMB[498][1] ) );
  FADDER S3_498_2 ( .CIN(\ab[498][2] ), .IN0(\CARRYB[497][2] ), .IN1(
        \ab[497][3] ), .COUT(\CARRYB[498][2] ), .SUM(\SUMB[498][2] ) );
  FADDER S1_497_0 ( .CIN(\ab[497][0] ), .IN0(\CARRYB[496][0] ), .IN1(
        \SUMB[496][1] ), .COUT(\CARRYB[497][0] ), .SUM(PRODUCT[497]) );
  FADDER S2_497_1 ( .CIN(\ab[497][1] ), .IN0(\CARRYB[496][1] ), .IN1(
        \SUMB[496][2] ), .COUT(\CARRYB[497][1] ), .SUM(\SUMB[497][1] ) );
  FADDER S3_497_2 ( .CIN(\ab[497][2] ), .IN0(\CARRYB[496][2] ), .IN1(
        \ab[496][3] ), .COUT(\CARRYB[497][2] ), .SUM(\SUMB[497][2] ) );
  FADDER S1_496_0 ( .CIN(\ab[496][0] ), .IN0(\CARRYB[495][0] ), .IN1(
        \SUMB[495][1] ), .COUT(\CARRYB[496][0] ), .SUM(PRODUCT[496]) );
  FADDER S2_496_1 ( .CIN(\ab[496][1] ), .IN0(\CARRYB[495][1] ), .IN1(
        \SUMB[495][2] ), .COUT(\CARRYB[496][1] ), .SUM(\SUMB[496][1] ) );
  FADDER S3_496_2 ( .CIN(\ab[496][2] ), .IN0(\CARRYB[495][2] ), .IN1(
        \ab[495][3] ), .COUT(\CARRYB[496][2] ), .SUM(\SUMB[496][2] ) );
  FADDER S1_495_0 ( .CIN(\ab[495][0] ), .IN0(\CARRYB[494][0] ), .IN1(
        \SUMB[494][1] ), .COUT(\CARRYB[495][0] ), .SUM(PRODUCT[495]) );
  FADDER S2_495_1 ( .CIN(\ab[495][1] ), .IN0(\CARRYB[494][1] ), .IN1(
        \SUMB[494][2] ), .COUT(\CARRYB[495][1] ), .SUM(\SUMB[495][1] ) );
  FADDER S3_495_2 ( .CIN(\ab[495][2] ), .IN0(\CARRYB[494][2] ), .IN1(
        \ab[494][3] ), .COUT(\CARRYB[495][2] ), .SUM(\SUMB[495][2] ) );
  FADDER S1_494_0 ( .CIN(\ab[494][0] ), .IN0(\CARRYB[493][0] ), .IN1(
        \SUMB[493][1] ), .COUT(\CARRYB[494][0] ), .SUM(PRODUCT[494]) );
  FADDER S2_494_1 ( .CIN(\ab[494][1] ), .IN0(\CARRYB[493][1] ), .IN1(
        \SUMB[493][2] ), .COUT(\CARRYB[494][1] ), .SUM(\SUMB[494][1] ) );
  FADDER S3_494_2 ( .CIN(\ab[494][2] ), .IN0(\CARRYB[493][2] ), .IN1(
        \ab[493][3] ), .COUT(\CARRYB[494][2] ), .SUM(\SUMB[494][2] ) );
  FADDER S1_493_0 ( .CIN(\ab[493][0] ), .IN0(\CARRYB[492][0] ), .IN1(
        \SUMB[492][1] ), .COUT(\CARRYB[493][0] ), .SUM(PRODUCT[493]) );
  FADDER S2_493_1 ( .CIN(\ab[493][1] ), .IN0(\CARRYB[492][1] ), .IN1(
        \SUMB[492][2] ), .COUT(\CARRYB[493][1] ), .SUM(\SUMB[493][1] ) );
  FADDER S3_493_2 ( .CIN(\ab[493][2] ), .IN0(\CARRYB[492][2] ), .IN1(
        \ab[492][3] ), .COUT(\CARRYB[493][2] ), .SUM(\SUMB[493][2] ) );
  FADDER S1_492_0 ( .CIN(\ab[492][0] ), .IN0(\CARRYB[491][0] ), .IN1(
        \SUMB[491][1] ), .COUT(\CARRYB[492][0] ), .SUM(PRODUCT[492]) );
  FADDER S2_492_1 ( .CIN(\ab[492][1] ), .IN0(\CARRYB[491][1] ), .IN1(
        \SUMB[491][2] ), .COUT(\CARRYB[492][1] ), .SUM(\SUMB[492][1] ) );
  FADDER S3_492_2 ( .CIN(\ab[492][2] ), .IN0(\CARRYB[491][2] ), .IN1(
        \ab[491][3] ), .COUT(\CARRYB[492][2] ), .SUM(\SUMB[492][2] ) );
  FADDER S1_491_0 ( .CIN(\ab[491][0] ), .IN0(\CARRYB[490][0] ), .IN1(
        \SUMB[490][1] ), .COUT(\CARRYB[491][0] ), .SUM(PRODUCT[491]) );
  FADDER S2_491_1 ( .CIN(\ab[491][1] ), .IN0(\CARRYB[490][1] ), .IN1(
        \SUMB[490][2] ), .COUT(\CARRYB[491][1] ), .SUM(\SUMB[491][1] ) );
  FADDER S3_491_2 ( .CIN(\ab[491][2] ), .IN0(\CARRYB[490][2] ), .IN1(
        \ab[490][3] ), .COUT(\CARRYB[491][2] ), .SUM(\SUMB[491][2] ) );
  FADDER S1_490_0 ( .CIN(\ab[490][0] ), .IN0(\CARRYB[489][0] ), .IN1(
        \SUMB[489][1] ), .COUT(\CARRYB[490][0] ), .SUM(PRODUCT[490]) );
  FADDER S2_490_1 ( .CIN(\ab[490][1] ), .IN0(\CARRYB[489][1] ), .IN1(
        \SUMB[489][2] ), .COUT(\CARRYB[490][1] ), .SUM(\SUMB[490][1] ) );
  FADDER S3_490_2 ( .CIN(\ab[490][2] ), .IN0(\CARRYB[489][2] ), .IN1(
        \ab[489][3] ), .COUT(\CARRYB[490][2] ), .SUM(\SUMB[490][2] ) );
  FADDER S1_489_0 ( .CIN(\ab[489][0] ), .IN0(\CARRYB[488][0] ), .IN1(
        \SUMB[488][1] ), .COUT(\CARRYB[489][0] ), .SUM(PRODUCT[489]) );
  FADDER S2_489_1 ( .CIN(\ab[489][1] ), .IN0(\CARRYB[488][1] ), .IN1(
        \SUMB[488][2] ), .COUT(\CARRYB[489][1] ), .SUM(\SUMB[489][1] ) );
  FADDER S3_489_2 ( .CIN(\ab[489][2] ), .IN0(\CARRYB[488][2] ), .IN1(
        \ab[488][3] ), .COUT(\CARRYB[489][2] ), .SUM(\SUMB[489][2] ) );
  FADDER S1_488_0 ( .CIN(\ab[488][0] ), .IN0(\CARRYB[487][0] ), .IN1(
        \SUMB[487][1] ), .COUT(\CARRYB[488][0] ), .SUM(PRODUCT[488]) );
  FADDER S2_488_1 ( .CIN(\ab[488][1] ), .IN0(\CARRYB[487][1] ), .IN1(
        \SUMB[487][2] ), .COUT(\CARRYB[488][1] ), .SUM(\SUMB[488][1] ) );
  FADDER S3_488_2 ( .CIN(\ab[488][2] ), .IN0(\CARRYB[487][2] ), .IN1(
        \ab[487][3] ), .COUT(\CARRYB[488][2] ), .SUM(\SUMB[488][2] ) );
  FADDER S1_487_0 ( .CIN(\ab[487][0] ), .IN0(\CARRYB[486][0] ), .IN1(
        \SUMB[486][1] ), .COUT(\CARRYB[487][0] ), .SUM(PRODUCT[487]) );
  FADDER S2_487_1 ( .CIN(\ab[487][1] ), .IN0(\CARRYB[486][1] ), .IN1(
        \SUMB[486][2] ), .COUT(\CARRYB[487][1] ), .SUM(\SUMB[487][1] ) );
  FADDER S3_487_2 ( .CIN(\ab[487][2] ), .IN0(\CARRYB[486][2] ), .IN1(
        \ab[486][3] ), .COUT(\CARRYB[487][2] ), .SUM(\SUMB[487][2] ) );
  FADDER S1_486_0 ( .CIN(\ab[486][0] ), .IN0(\CARRYB[485][0] ), .IN1(
        \SUMB[485][1] ), .COUT(\CARRYB[486][0] ), .SUM(PRODUCT[486]) );
  FADDER S2_486_1 ( .CIN(\ab[486][1] ), .IN0(\CARRYB[485][1] ), .IN1(
        \SUMB[485][2] ), .COUT(\CARRYB[486][1] ), .SUM(\SUMB[486][1] ) );
  FADDER S3_486_2 ( .CIN(\ab[486][2] ), .IN0(\CARRYB[485][2] ), .IN1(
        \ab[485][3] ), .COUT(\CARRYB[486][2] ), .SUM(\SUMB[486][2] ) );
  FADDER S1_485_0 ( .CIN(\ab[485][0] ), .IN0(\CARRYB[484][0] ), .IN1(
        \SUMB[484][1] ), .COUT(\CARRYB[485][0] ), .SUM(PRODUCT[485]) );
  FADDER S2_485_1 ( .CIN(\ab[485][1] ), .IN0(\CARRYB[484][1] ), .IN1(
        \SUMB[484][2] ), .COUT(\CARRYB[485][1] ), .SUM(\SUMB[485][1] ) );
  FADDER S3_485_2 ( .CIN(\ab[485][2] ), .IN0(\CARRYB[484][2] ), .IN1(
        \ab[484][3] ), .COUT(\CARRYB[485][2] ), .SUM(\SUMB[485][2] ) );
  FADDER S1_484_0 ( .CIN(\ab[484][0] ), .IN0(\CARRYB[483][0] ), .IN1(
        \SUMB[483][1] ), .COUT(\CARRYB[484][0] ), .SUM(PRODUCT[484]) );
  FADDER S2_484_1 ( .CIN(\ab[484][1] ), .IN0(\CARRYB[483][1] ), .IN1(
        \SUMB[483][2] ), .COUT(\CARRYB[484][1] ), .SUM(\SUMB[484][1] ) );
  FADDER S3_484_2 ( .CIN(\ab[484][2] ), .IN0(\CARRYB[483][2] ), .IN1(
        \ab[483][3] ), .COUT(\CARRYB[484][2] ), .SUM(\SUMB[484][2] ) );
  FADDER S1_483_0 ( .CIN(\ab[483][0] ), .IN0(\CARRYB[482][0] ), .IN1(
        \SUMB[482][1] ), .COUT(\CARRYB[483][0] ), .SUM(PRODUCT[483]) );
  FADDER S2_483_1 ( .CIN(\ab[483][1] ), .IN0(\CARRYB[482][1] ), .IN1(
        \SUMB[482][2] ), .COUT(\CARRYB[483][1] ), .SUM(\SUMB[483][1] ) );
  FADDER S3_483_2 ( .CIN(\ab[483][2] ), .IN0(\CARRYB[482][2] ), .IN1(
        \ab[482][3] ), .COUT(\CARRYB[483][2] ), .SUM(\SUMB[483][2] ) );
  FADDER S1_482_0 ( .CIN(\ab[482][0] ), .IN0(\CARRYB[481][0] ), .IN1(
        \SUMB[481][1] ), .COUT(\CARRYB[482][0] ), .SUM(PRODUCT[482]) );
  FADDER S2_482_1 ( .CIN(\ab[482][1] ), .IN0(\CARRYB[481][1] ), .IN1(
        \SUMB[481][2] ), .COUT(\CARRYB[482][1] ), .SUM(\SUMB[482][1] ) );
  FADDER S3_482_2 ( .CIN(\ab[482][2] ), .IN0(\CARRYB[481][2] ), .IN1(
        \ab[481][3] ), .COUT(\CARRYB[482][2] ), .SUM(\SUMB[482][2] ) );
  FADDER S1_481_0 ( .CIN(\ab[481][0] ), .IN0(\CARRYB[480][0] ), .IN1(
        \SUMB[480][1] ), .COUT(\CARRYB[481][0] ), .SUM(PRODUCT[481]) );
  FADDER S2_481_1 ( .CIN(\ab[481][1] ), .IN0(\CARRYB[480][1] ), .IN1(
        \SUMB[480][2] ), .COUT(\CARRYB[481][1] ), .SUM(\SUMB[481][1] ) );
  FADDER S3_481_2 ( .CIN(\ab[481][2] ), .IN0(\CARRYB[480][2] ), .IN1(
        \ab[480][3] ), .COUT(\CARRYB[481][2] ), .SUM(\SUMB[481][2] ) );
  FADDER S1_480_0 ( .CIN(\ab[480][0] ), .IN0(\CARRYB[479][0] ), .IN1(
        \SUMB[479][1] ), .COUT(\CARRYB[480][0] ), .SUM(PRODUCT[480]) );
  FADDER S2_480_1 ( .CIN(\ab[480][1] ), .IN0(\CARRYB[479][1] ), .IN1(
        \SUMB[479][2] ), .COUT(\CARRYB[480][1] ), .SUM(\SUMB[480][1] ) );
  FADDER S3_480_2 ( .CIN(\ab[480][2] ), .IN0(\CARRYB[479][2] ), .IN1(
        \ab[479][3] ), .COUT(\CARRYB[480][2] ), .SUM(\SUMB[480][2] ) );
  FADDER S1_479_0 ( .CIN(\ab[479][0] ), .IN0(\CARRYB[478][0] ), .IN1(
        \SUMB[478][1] ), .COUT(\CARRYB[479][0] ), .SUM(PRODUCT[479]) );
  FADDER S2_479_1 ( .CIN(\ab[479][1] ), .IN0(\CARRYB[478][1] ), .IN1(
        \SUMB[478][2] ), .COUT(\CARRYB[479][1] ), .SUM(\SUMB[479][1] ) );
  FADDER S3_479_2 ( .CIN(\ab[479][2] ), .IN0(\CARRYB[478][2] ), .IN1(
        \ab[478][3] ), .COUT(\CARRYB[479][2] ), .SUM(\SUMB[479][2] ) );
  FADDER S1_478_0 ( .CIN(\ab[478][0] ), .IN0(\CARRYB[477][0] ), .IN1(
        \SUMB[477][1] ), .COUT(\CARRYB[478][0] ), .SUM(PRODUCT[478]) );
  FADDER S2_478_1 ( .CIN(\ab[478][1] ), .IN0(\CARRYB[477][1] ), .IN1(
        \SUMB[477][2] ), .COUT(\CARRYB[478][1] ), .SUM(\SUMB[478][1] ) );
  FADDER S3_478_2 ( .CIN(\ab[478][2] ), .IN0(\CARRYB[477][2] ), .IN1(
        \ab[477][3] ), .COUT(\CARRYB[478][2] ), .SUM(\SUMB[478][2] ) );
  FADDER S1_477_0 ( .CIN(\ab[477][0] ), .IN0(\CARRYB[476][0] ), .IN1(
        \SUMB[476][1] ), .COUT(\CARRYB[477][0] ), .SUM(PRODUCT[477]) );
  FADDER S2_477_1 ( .CIN(\ab[477][1] ), .IN0(\CARRYB[476][1] ), .IN1(
        \SUMB[476][2] ), .COUT(\CARRYB[477][1] ), .SUM(\SUMB[477][1] ) );
  FADDER S3_477_2 ( .CIN(\ab[477][2] ), .IN0(\CARRYB[476][2] ), .IN1(
        \ab[476][3] ), .COUT(\CARRYB[477][2] ), .SUM(\SUMB[477][2] ) );
  FADDER S1_476_0 ( .CIN(\ab[476][0] ), .IN0(\CARRYB[475][0] ), .IN1(
        \SUMB[475][1] ), .COUT(\CARRYB[476][0] ), .SUM(PRODUCT[476]) );
  FADDER S2_476_1 ( .CIN(\ab[476][1] ), .IN0(\CARRYB[475][1] ), .IN1(
        \SUMB[475][2] ), .COUT(\CARRYB[476][1] ), .SUM(\SUMB[476][1] ) );
  FADDER S3_476_2 ( .CIN(\ab[476][2] ), .IN0(\CARRYB[475][2] ), .IN1(
        \ab[475][3] ), .COUT(\CARRYB[476][2] ), .SUM(\SUMB[476][2] ) );
  FADDER S1_475_0 ( .CIN(\ab[475][0] ), .IN0(\CARRYB[474][0] ), .IN1(
        \SUMB[474][1] ), .COUT(\CARRYB[475][0] ), .SUM(PRODUCT[475]) );
  FADDER S2_475_1 ( .CIN(\ab[475][1] ), .IN0(\CARRYB[474][1] ), .IN1(
        \SUMB[474][2] ), .COUT(\CARRYB[475][1] ), .SUM(\SUMB[475][1] ) );
  FADDER S3_475_2 ( .CIN(\ab[475][2] ), .IN0(\CARRYB[474][2] ), .IN1(
        \ab[474][3] ), .COUT(\CARRYB[475][2] ), .SUM(\SUMB[475][2] ) );
  FADDER S1_474_0 ( .CIN(\ab[474][0] ), .IN0(\CARRYB[473][0] ), .IN1(
        \SUMB[473][1] ), .COUT(\CARRYB[474][0] ), .SUM(PRODUCT[474]) );
  FADDER S2_474_1 ( .CIN(\ab[474][1] ), .IN0(\CARRYB[473][1] ), .IN1(
        \SUMB[473][2] ), .COUT(\CARRYB[474][1] ), .SUM(\SUMB[474][1] ) );
  FADDER S3_474_2 ( .CIN(\ab[474][2] ), .IN0(\CARRYB[473][2] ), .IN1(
        \ab[473][3] ), .COUT(\CARRYB[474][2] ), .SUM(\SUMB[474][2] ) );
  FADDER S1_473_0 ( .CIN(\ab[473][0] ), .IN0(\CARRYB[472][0] ), .IN1(
        \SUMB[472][1] ), .COUT(\CARRYB[473][0] ), .SUM(PRODUCT[473]) );
  FADDER S2_473_1 ( .CIN(\ab[473][1] ), .IN0(\CARRYB[472][1] ), .IN1(
        \SUMB[472][2] ), .COUT(\CARRYB[473][1] ), .SUM(\SUMB[473][1] ) );
  FADDER S3_473_2 ( .CIN(\ab[473][2] ), .IN0(\CARRYB[472][2] ), .IN1(
        \ab[472][3] ), .COUT(\CARRYB[473][2] ), .SUM(\SUMB[473][2] ) );
  FADDER S1_472_0 ( .CIN(\ab[472][0] ), .IN0(\CARRYB[471][0] ), .IN1(
        \SUMB[471][1] ), .COUT(\CARRYB[472][0] ), .SUM(PRODUCT[472]) );
  FADDER S2_472_1 ( .CIN(\ab[472][1] ), .IN0(\CARRYB[471][1] ), .IN1(
        \SUMB[471][2] ), .COUT(\CARRYB[472][1] ), .SUM(\SUMB[472][1] ) );
  FADDER S3_472_2 ( .CIN(\ab[472][2] ), .IN0(\CARRYB[471][2] ), .IN1(
        \ab[471][3] ), .COUT(\CARRYB[472][2] ), .SUM(\SUMB[472][2] ) );
  FADDER S1_471_0 ( .CIN(\ab[471][0] ), .IN0(\CARRYB[470][0] ), .IN1(
        \SUMB[470][1] ), .COUT(\CARRYB[471][0] ), .SUM(PRODUCT[471]) );
  FADDER S2_471_1 ( .CIN(\ab[471][1] ), .IN0(\CARRYB[470][1] ), .IN1(
        \SUMB[470][2] ), .COUT(\CARRYB[471][1] ), .SUM(\SUMB[471][1] ) );
  FADDER S3_471_2 ( .CIN(\ab[471][2] ), .IN0(\CARRYB[470][2] ), .IN1(
        \ab[470][3] ), .COUT(\CARRYB[471][2] ), .SUM(\SUMB[471][2] ) );
  FADDER S1_470_0 ( .CIN(\ab[470][0] ), .IN0(\CARRYB[469][0] ), .IN1(
        \SUMB[469][1] ), .COUT(\CARRYB[470][0] ), .SUM(PRODUCT[470]) );
  FADDER S2_470_1 ( .CIN(\ab[470][1] ), .IN0(\CARRYB[469][1] ), .IN1(
        \SUMB[469][2] ), .COUT(\CARRYB[470][1] ), .SUM(\SUMB[470][1] ) );
  FADDER S3_470_2 ( .CIN(\ab[470][2] ), .IN0(\CARRYB[469][2] ), .IN1(
        \ab[469][3] ), .COUT(\CARRYB[470][2] ), .SUM(\SUMB[470][2] ) );
  FADDER S1_469_0 ( .CIN(\ab[469][0] ), .IN0(\CARRYB[468][0] ), .IN1(
        \SUMB[468][1] ), .COUT(\CARRYB[469][0] ), .SUM(PRODUCT[469]) );
  FADDER S2_469_1 ( .CIN(\ab[469][1] ), .IN0(\CARRYB[468][1] ), .IN1(
        \SUMB[468][2] ), .COUT(\CARRYB[469][1] ), .SUM(\SUMB[469][1] ) );
  FADDER S3_469_2 ( .CIN(\ab[469][2] ), .IN0(\CARRYB[468][2] ), .IN1(
        \ab[468][3] ), .COUT(\CARRYB[469][2] ), .SUM(\SUMB[469][2] ) );
  FADDER S1_468_0 ( .CIN(\ab[468][0] ), .IN0(\CARRYB[467][0] ), .IN1(
        \SUMB[467][1] ), .COUT(\CARRYB[468][0] ), .SUM(PRODUCT[468]) );
  FADDER S2_468_1 ( .CIN(\ab[468][1] ), .IN0(\CARRYB[467][1] ), .IN1(
        \SUMB[467][2] ), .COUT(\CARRYB[468][1] ), .SUM(\SUMB[468][1] ) );
  FADDER S3_468_2 ( .CIN(\ab[468][2] ), .IN0(\CARRYB[467][2] ), .IN1(
        \ab[467][3] ), .COUT(\CARRYB[468][2] ), .SUM(\SUMB[468][2] ) );
  FADDER S1_467_0 ( .CIN(\ab[467][0] ), .IN0(\CARRYB[466][0] ), .IN1(
        \SUMB[466][1] ), .COUT(\CARRYB[467][0] ), .SUM(PRODUCT[467]) );
  FADDER S2_467_1 ( .CIN(\ab[467][1] ), .IN0(\CARRYB[466][1] ), .IN1(
        \SUMB[466][2] ), .COUT(\CARRYB[467][1] ), .SUM(\SUMB[467][1] ) );
  FADDER S3_467_2 ( .CIN(\ab[467][2] ), .IN0(\CARRYB[466][2] ), .IN1(
        \ab[466][3] ), .COUT(\CARRYB[467][2] ), .SUM(\SUMB[467][2] ) );
  FADDER S1_466_0 ( .CIN(\ab[466][0] ), .IN0(\CARRYB[465][0] ), .IN1(
        \SUMB[465][1] ), .COUT(\CARRYB[466][0] ), .SUM(PRODUCT[466]) );
  FADDER S2_466_1 ( .CIN(\ab[466][1] ), .IN0(\CARRYB[465][1] ), .IN1(
        \SUMB[465][2] ), .COUT(\CARRYB[466][1] ), .SUM(\SUMB[466][1] ) );
  FADDER S3_466_2 ( .CIN(\ab[466][2] ), .IN0(\CARRYB[465][2] ), .IN1(
        \ab[465][3] ), .COUT(\CARRYB[466][2] ), .SUM(\SUMB[466][2] ) );
  FADDER S1_465_0 ( .CIN(\ab[465][0] ), .IN0(\CARRYB[464][0] ), .IN1(
        \SUMB[464][1] ), .COUT(\CARRYB[465][0] ), .SUM(PRODUCT[465]) );
  FADDER S2_465_1 ( .CIN(\ab[465][1] ), .IN0(\CARRYB[464][1] ), .IN1(
        \SUMB[464][2] ), .COUT(\CARRYB[465][1] ), .SUM(\SUMB[465][1] ) );
  FADDER S3_465_2 ( .CIN(\ab[465][2] ), .IN0(\CARRYB[464][2] ), .IN1(
        \ab[464][3] ), .COUT(\CARRYB[465][2] ), .SUM(\SUMB[465][2] ) );
  FADDER S1_464_0 ( .CIN(\ab[464][0] ), .IN0(\CARRYB[463][0] ), .IN1(
        \SUMB[463][1] ), .COUT(\CARRYB[464][0] ), .SUM(PRODUCT[464]) );
  FADDER S2_464_1 ( .CIN(\ab[464][1] ), .IN0(\CARRYB[463][1] ), .IN1(
        \SUMB[463][2] ), .COUT(\CARRYB[464][1] ), .SUM(\SUMB[464][1] ) );
  FADDER S3_464_2 ( .CIN(\ab[464][2] ), .IN0(\CARRYB[463][2] ), .IN1(
        \ab[463][3] ), .COUT(\CARRYB[464][2] ), .SUM(\SUMB[464][2] ) );
  FADDER S1_463_0 ( .CIN(\ab[463][0] ), .IN0(\CARRYB[462][0] ), .IN1(
        \SUMB[462][1] ), .COUT(\CARRYB[463][0] ), .SUM(PRODUCT[463]) );
  FADDER S2_463_1 ( .CIN(\ab[463][1] ), .IN0(\CARRYB[462][1] ), .IN1(
        \SUMB[462][2] ), .COUT(\CARRYB[463][1] ), .SUM(\SUMB[463][1] ) );
  FADDER S3_463_2 ( .CIN(\ab[463][2] ), .IN0(\CARRYB[462][2] ), .IN1(
        \ab[462][3] ), .COUT(\CARRYB[463][2] ), .SUM(\SUMB[463][2] ) );
  FADDER S1_462_0 ( .CIN(\ab[462][0] ), .IN0(\CARRYB[461][0] ), .IN1(
        \SUMB[461][1] ), .COUT(\CARRYB[462][0] ), .SUM(PRODUCT[462]) );
  FADDER S2_462_1 ( .CIN(\ab[462][1] ), .IN0(\CARRYB[461][1] ), .IN1(
        \SUMB[461][2] ), .COUT(\CARRYB[462][1] ), .SUM(\SUMB[462][1] ) );
  FADDER S3_462_2 ( .CIN(\ab[462][2] ), .IN0(\CARRYB[461][2] ), .IN1(
        \ab[461][3] ), .COUT(\CARRYB[462][2] ), .SUM(\SUMB[462][2] ) );
  FADDER S1_461_0 ( .CIN(\ab[461][0] ), .IN0(\CARRYB[460][0] ), .IN1(
        \SUMB[460][1] ), .COUT(\CARRYB[461][0] ), .SUM(PRODUCT[461]) );
  FADDER S2_461_1 ( .CIN(\ab[461][1] ), .IN0(\CARRYB[460][1] ), .IN1(
        \SUMB[460][2] ), .COUT(\CARRYB[461][1] ), .SUM(\SUMB[461][1] ) );
  FADDER S3_461_2 ( .CIN(\ab[461][2] ), .IN0(\CARRYB[460][2] ), .IN1(
        \ab[460][3] ), .COUT(\CARRYB[461][2] ), .SUM(\SUMB[461][2] ) );
  FADDER S1_460_0 ( .CIN(\ab[460][0] ), .IN0(\CARRYB[459][0] ), .IN1(
        \SUMB[459][1] ), .COUT(\CARRYB[460][0] ), .SUM(PRODUCT[460]) );
  FADDER S2_460_1 ( .CIN(\ab[460][1] ), .IN0(\CARRYB[459][1] ), .IN1(
        \SUMB[459][2] ), .COUT(\CARRYB[460][1] ), .SUM(\SUMB[460][1] ) );
  FADDER S3_460_2 ( .CIN(\ab[460][2] ), .IN0(\CARRYB[459][2] ), .IN1(
        \ab[459][3] ), .COUT(\CARRYB[460][2] ), .SUM(\SUMB[460][2] ) );
  FADDER S1_459_0 ( .CIN(\ab[459][0] ), .IN0(\CARRYB[458][0] ), .IN1(
        \SUMB[458][1] ), .COUT(\CARRYB[459][0] ), .SUM(PRODUCT[459]) );
  FADDER S2_459_1 ( .CIN(\ab[459][1] ), .IN0(\CARRYB[458][1] ), .IN1(
        \SUMB[458][2] ), .COUT(\CARRYB[459][1] ), .SUM(\SUMB[459][1] ) );
  FADDER S3_459_2 ( .CIN(\ab[459][2] ), .IN0(\CARRYB[458][2] ), .IN1(
        \ab[458][3] ), .COUT(\CARRYB[459][2] ), .SUM(\SUMB[459][2] ) );
  FADDER S1_458_0 ( .CIN(\ab[458][0] ), .IN0(\CARRYB[457][0] ), .IN1(
        \SUMB[457][1] ), .COUT(\CARRYB[458][0] ), .SUM(PRODUCT[458]) );
  FADDER S2_458_1 ( .CIN(\ab[458][1] ), .IN0(\CARRYB[457][1] ), .IN1(
        \SUMB[457][2] ), .COUT(\CARRYB[458][1] ), .SUM(\SUMB[458][1] ) );
  FADDER S3_458_2 ( .CIN(\ab[458][2] ), .IN0(\CARRYB[457][2] ), .IN1(
        \ab[457][3] ), .COUT(\CARRYB[458][2] ), .SUM(\SUMB[458][2] ) );
  FADDER S1_457_0 ( .CIN(\ab[457][0] ), .IN0(\CARRYB[456][0] ), .IN1(
        \SUMB[456][1] ), .COUT(\CARRYB[457][0] ), .SUM(PRODUCT[457]) );
  FADDER S2_457_1 ( .CIN(\ab[457][1] ), .IN0(\CARRYB[456][1] ), .IN1(
        \SUMB[456][2] ), .COUT(\CARRYB[457][1] ), .SUM(\SUMB[457][1] ) );
  FADDER S3_457_2 ( .CIN(\ab[457][2] ), .IN0(\CARRYB[456][2] ), .IN1(
        \ab[456][3] ), .COUT(\CARRYB[457][2] ), .SUM(\SUMB[457][2] ) );
  FADDER S1_456_0 ( .CIN(\ab[456][0] ), .IN0(\CARRYB[455][0] ), .IN1(
        \SUMB[455][1] ), .COUT(\CARRYB[456][0] ), .SUM(PRODUCT[456]) );
  FADDER S2_456_1 ( .CIN(\ab[456][1] ), .IN0(\CARRYB[455][1] ), .IN1(
        \SUMB[455][2] ), .COUT(\CARRYB[456][1] ), .SUM(\SUMB[456][1] ) );
  FADDER S3_456_2 ( .CIN(\ab[456][2] ), .IN0(\CARRYB[455][2] ), .IN1(
        \ab[455][3] ), .COUT(\CARRYB[456][2] ), .SUM(\SUMB[456][2] ) );
  FADDER S1_455_0 ( .CIN(\ab[455][0] ), .IN0(\CARRYB[454][0] ), .IN1(
        \SUMB[454][1] ), .COUT(\CARRYB[455][0] ), .SUM(PRODUCT[455]) );
  FADDER S2_455_1 ( .CIN(\ab[455][1] ), .IN0(\CARRYB[454][1] ), .IN1(
        \SUMB[454][2] ), .COUT(\CARRYB[455][1] ), .SUM(\SUMB[455][1] ) );
  FADDER S3_455_2 ( .CIN(\ab[455][2] ), .IN0(\CARRYB[454][2] ), .IN1(
        \ab[454][3] ), .COUT(\CARRYB[455][2] ), .SUM(\SUMB[455][2] ) );
  FADDER S1_454_0 ( .CIN(\ab[454][0] ), .IN0(\CARRYB[453][0] ), .IN1(
        \SUMB[453][1] ), .COUT(\CARRYB[454][0] ), .SUM(PRODUCT[454]) );
  FADDER S2_454_1 ( .CIN(\ab[454][1] ), .IN0(\CARRYB[453][1] ), .IN1(
        \SUMB[453][2] ), .COUT(\CARRYB[454][1] ), .SUM(\SUMB[454][1] ) );
  FADDER S3_454_2 ( .CIN(\ab[454][2] ), .IN0(\CARRYB[453][2] ), .IN1(
        \ab[453][3] ), .COUT(\CARRYB[454][2] ), .SUM(\SUMB[454][2] ) );
  FADDER S1_453_0 ( .CIN(\ab[453][0] ), .IN0(\CARRYB[452][0] ), .IN1(
        \SUMB[452][1] ), .COUT(\CARRYB[453][0] ), .SUM(PRODUCT[453]) );
  FADDER S2_453_1 ( .CIN(\ab[453][1] ), .IN0(\CARRYB[452][1] ), .IN1(
        \SUMB[452][2] ), .COUT(\CARRYB[453][1] ), .SUM(\SUMB[453][1] ) );
  FADDER S3_453_2 ( .CIN(\ab[453][2] ), .IN0(\CARRYB[452][2] ), .IN1(
        \ab[452][3] ), .COUT(\CARRYB[453][2] ), .SUM(\SUMB[453][2] ) );
  FADDER S1_452_0 ( .CIN(\ab[452][0] ), .IN0(\CARRYB[451][0] ), .IN1(
        \SUMB[451][1] ), .COUT(\CARRYB[452][0] ), .SUM(PRODUCT[452]) );
  FADDER S2_452_1 ( .CIN(\ab[452][1] ), .IN0(\CARRYB[451][1] ), .IN1(
        \SUMB[451][2] ), .COUT(\CARRYB[452][1] ), .SUM(\SUMB[452][1] ) );
  FADDER S3_452_2 ( .CIN(\ab[452][2] ), .IN0(\CARRYB[451][2] ), .IN1(
        \ab[451][3] ), .COUT(\CARRYB[452][2] ), .SUM(\SUMB[452][2] ) );
  FADDER S1_451_0 ( .CIN(\ab[451][0] ), .IN0(\CARRYB[450][0] ), .IN1(
        \SUMB[450][1] ), .COUT(\CARRYB[451][0] ), .SUM(PRODUCT[451]) );
  FADDER S2_451_1 ( .CIN(\ab[451][1] ), .IN0(\CARRYB[450][1] ), .IN1(
        \SUMB[450][2] ), .COUT(\CARRYB[451][1] ), .SUM(\SUMB[451][1] ) );
  FADDER S3_451_2 ( .CIN(\ab[451][2] ), .IN0(\CARRYB[450][2] ), .IN1(
        \ab[450][3] ), .COUT(\CARRYB[451][2] ), .SUM(\SUMB[451][2] ) );
  FADDER S1_450_0 ( .CIN(\ab[450][0] ), .IN0(\CARRYB[449][0] ), .IN1(
        \SUMB[449][1] ), .COUT(\CARRYB[450][0] ), .SUM(PRODUCT[450]) );
  FADDER S2_450_1 ( .CIN(\ab[450][1] ), .IN0(\CARRYB[449][1] ), .IN1(
        \SUMB[449][2] ), .COUT(\CARRYB[450][1] ), .SUM(\SUMB[450][1] ) );
  FADDER S3_450_2 ( .CIN(\ab[450][2] ), .IN0(\CARRYB[449][2] ), .IN1(
        \ab[449][3] ), .COUT(\CARRYB[450][2] ), .SUM(\SUMB[450][2] ) );
  FADDER S1_449_0 ( .CIN(\ab[449][0] ), .IN0(\CARRYB[448][0] ), .IN1(
        \SUMB[448][1] ), .COUT(\CARRYB[449][0] ), .SUM(PRODUCT[449]) );
  FADDER S2_449_1 ( .CIN(\ab[449][1] ), .IN0(\CARRYB[448][1] ), .IN1(
        \SUMB[448][2] ), .COUT(\CARRYB[449][1] ), .SUM(\SUMB[449][1] ) );
  FADDER S3_449_2 ( .CIN(\ab[449][2] ), .IN0(\CARRYB[448][2] ), .IN1(
        \ab[448][3] ), .COUT(\CARRYB[449][2] ), .SUM(\SUMB[449][2] ) );
  FADDER S1_448_0 ( .CIN(\ab[448][0] ), .IN0(\CARRYB[447][0] ), .IN1(
        \SUMB[447][1] ), .COUT(\CARRYB[448][0] ), .SUM(PRODUCT[448]) );
  FADDER S2_448_1 ( .CIN(\ab[448][1] ), .IN0(\CARRYB[447][1] ), .IN1(
        \SUMB[447][2] ), .COUT(\CARRYB[448][1] ), .SUM(\SUMB[448][1] ) );
  FADDER S3_448_2 ( .CIN(\ab[448][2] ), .IN0(\CARRYB[447][2] ), .IN1(
        \ab[447][3] ), .COUT(\CARRYB[448][2] ), .SUM(\SUMB[448][2] ) );
  FADDER S1_447_0 ( .CIN(\ab[447][0] ), .IN0(\CARRYB[446][0] ), .IN1(
        \SUMB[446][1] ), .COUT(\CARRYB[447][0] ), .SUM(PRODUCT[447]) );
  FADDER S2_447_1 ( .CIN(\ab[447][1] ), .IN0(\CARRYB[446][1] ), .IN1(
        \SUMB[446][2] ), .COUT(\CARRYB[447][1] ), .SUM(\SUMB[447][1] ) );
  FADDER S3_447_2 ( .CIN(\ab[447][2] ), .IN0(\CARRYB[446][2] ), .IN1(
        \ab[446][3] ), .COUT(\CARRYB[447][2] ), .SUM(\SUMB[447][2] ) );
  FADDER S1_446_0 ( .CIN(\ab[446][0] ), .IN0(\CARRYB[445][0] ), .IN1(
        \SUMB[445][1] ), .COUT(\CARRYB[446][0] ), .SUM(PRODUCT[446]) );
  FADDER S2_446_1 ( .CIN(\ab[446][1] ), .IN0(\CARRYB[445][1] ), .IN1(
        \SUMB[445][2] ), .COUT(\CARRYB[446][1] ), .SUM(\SUMB[446][1] ) );
  FADDER S3_446_2 ( .CIN(\ab[446][2] ), .IN0(\CARRYB[445][2] ), .IN1(
        \ab[445][3] ), .COUT(\CARRYB[446][2] ), .SUM(\SUMB[446][2] ) );
  FADDER S1_445_0 ( .CIN(\ab[445][0] ), .IN0(\CARRYB[444][0] ), .IN1(
        \SUMB[444][1] ), .COUT(\CARRYB[445][0] ), .SUM(PRODUCT[445]) );
  FADDER S2_445_1 ( .CIN(\ab[445][1] ), .IN0(\CARRYB[444][1] ), .IN1(
        \SUMB[444][2] ), .COUT(\CARRYB[445][1] ), .SUM(\SUMB[445][1] ) );
  FADDER S3_445_2 ( .CIN(\ab[445][2] ), .IN0(\CARRYB[444][2] ), .IN1(
        \ab[444][3] ), .COUT(\CARRYB[445][2] ), .SUM(\SUMB[445][2] ) );
  FADDER S1_444_0 ( .CIN(\ab[444][0] ), .IN0(\CARRYB[443][0] ), .IN1(
        \SUMB[443][1] ), .COUT(\CARRYB[444][0] ), .SUM(PRODUCT[444]) );
  FADDER S2_444_1 ( .CIN(\ab[444][1] ), .IN0(\CARRYB[443][1] ), .IN1(
        \SUMB[443][2] ), .COUT(\CARRYB[444][1] ), .SUM(\SUMB[444][1] ) );
  FADDER S3_444_2 ( .CIN(\ab[444][2] ), .IN0(\CARRYB[443][2] ), .IN1(
        \ab[443][3] ), .COUT(\CARRYB[444][2] ), .SUM(\SUMB[444][2] ) );
  FADDER S1_443_0 ( .CIN(\ab[443][0] ), .IN0(\CARRYB[442][0] ), .IN1(
        \SUMB[442][1] ), .COUT(\CARRYB[443][0] ), .SUM(PRODUCT[443]) );
  FADDER S2_443_1 ( .CIN(\ab[443][1] ), .IN0(\CARRYB[442][1] ), .IN1(
        \SUMB[442][2] ), .COUT(\CARRYB[443][1] ), .SUM(\SUMB[443][1] ) );
  FADDER S3_443_2 ( .CIN(\ab[443][2] ), .IN0(\CARRYB[442][2] ), .IN1(
        \ab[442][3] ), .COUT(\CARRYB[443][2] ), .SUM(\SUMB[443][2] ) );
  FADDER S1_442_0 ( .CIN(\ab[442][0] ), .IN0(\CARRYB[441][0] ), .IN1(
        \SUMB[441][1] ), .COUT(\CARRYB[442][0] ), .SUM(PRODUCT[442]) );
  FADDER S2_442_1 ( .CIN(\ab[442][1] ), .IN0(\CARRYB[441][1] ), .IN1(
        \SUMB[441][2] ), .COUT(\CARRYB[442][1] ), .SUM(\SUMB[442][1] ) );
  FADDER S3_442_2 ( .CIN(\ab[442][2] ), .IN0(\CARRYB[441][2] ), .IN1(
        \ab[441][3] ), .COUT(\CARRYB[442][2] ), .SUM(\SUMB[442][2] ) );
  FADDER S1_441_0 ( .CIN(\ab[441][0] ), .IN0(\CARRYB[440][0] ), .IN1(
        \SUMB[440][1] ), .COUT(\CARRYB[441][0] ), .SUM(PRODUCT[441]) );
  FADDER S2_441_1 ( .CIN(\ab[441][1] ), .IN0(\CARRYB[440][1] ), .IN1(
        \SUMB[440][2] ), .COUT(\CARRYB[441][1] ), .SUM(\SUMB[441][1] ) );
  FADDER S3_441_2 ( .CIN(\ab[441][2] ), .IN0(\CARRYB[440][2] ), .IN1(
        \ab[440][3] ), .COUT(\CARRYB[441][2] ), .SUM(\SUMB[441][2] ) );
  FADDER S1_440_0 ( .CIN(\ab[440][0] ), .IN0(\CARRYB[439][0] ), .IN1(
        \SUMB[439][1] ), .COUT(\CARRYB[440][0] ), .SUM(PRODUCT[440]) );
  FADDER S2_440_1 ( .CIN(\ab[440][1] ), .IN0(\CARRYB[439][1] ), .IN1(
        \SUMB[439][2] ), .COUT(\CARRYB[440][1] ), .SUM(\SUMB[440][1] ) );
  FADDER S3_440_2 ( .CIN(\ab[440][2] ), .IN0(\CARRYB[439][2] ), .IN1(
        \ab[439][3] ), .COUT(\CARRYB[440][2] ), .SUM(\SUMB[440][2] ) );
  FADDER S1_439_0 ( .CIN(\ab[439][0] ), .IN0(\CARRYB[438][0] ), .IN1(
        \SUMB[438][1] ), .COUT(\CARRYB[439][0] ), .SUM(PRODUCT[439]) );
  FADDER S2_439_1 ( .CIN(\ab[439][1] ), .IN0(\CARRYB[438][1] ), .IN1(
        \SUMB[438][2] ), .COUT(\CARRYB[439][1] ), .SUM(\SUMB[439][1] ) );
  FADDER S3_439_2 ( .CIN(\ab[439][2] ), .IN0(\CARRYB[438][2] ), .IN1(
        \ab[438][3] ), .COUT(\CARRYB[439][2] ), .SUM(\SUMB[439][2] ) );
  FADDER S1_438_0 ( .CIN(\ab[438][0] ), .IN0(\CARRYB[437][0] ), .IN1(
        \SUMB[437][1] ), .COUT(\CARRYB[438][0] ), .SUM(PRODUCT[438]) );
  FADDER S2_438_1 ( .CIN(\ab[438][1] ), .IN0(\CARRYB[437][1] ), .IN1(
        \SUMB[437][2] ), .COUT(\CARRYB[438][1] ), .SUM(\SUMB[438][1] ) );
  FADDER S3_438_2 ( .CIN(\ab[438][2] ), .IN0(\CARRYB[437][2] ), .IN1(
        \ab[437][3] ), .COUT(\CARRYB[438][2] ), .SUM(\SUMB[438][2] ) );
  FADDER S1_437_0 ( .CIN(\ab[437][0] ), .IN0(\CARRYB[436][0] ), .IN1(
        \SUMB[436][1] ), .COUT(\CARRYB[437][0] ), .SUM(PRODUCT[437]) );
  FADDER S2_437_1 ( .CIN(\ab[437][1] ), .IN0(\CARRYB[436][1] ), .IN1(
        \SUMB[436][2] ), .COUT(\CARRYB[437][1] ), .SUM(\SUMB[437][1] ) );
  FADDER S3_437_2 ( .CIN(\ab[437][2] ), .IN0(\CARRYB[436][2] ), .IN1(
        \ab[436][3] ), .COUT(\CARRYB[437][2] ), .SUM(\SUMB[437][2] ) );
  FADDER S1_436_0 ( .CIN(\ab[436][0] ), .IN0(\CARRYB[435][0] ), .IN1(
        \SUMB[435][1] ), .COUT(\CARRYB[436][0] ), .SUM(PRODUCT[436]) );
  FADDER S2_436_1 ( .CIN(\ab[436][1] ), .IN0(\CARRYB[435][1] ), .IN1(
        \SUMB[435][2] ), .COUT(\CARRYB[436][1] ), .SUM(\SUMB[436][1] ) );
  FADDER S3_436_2 ( .CIN(\ab[436][2] ), .IN0(\CARRYB[435][2] ), .IN1(
        \ab[435][3] ), .COUT(\CARRYB[436][2] ), .SUM(\SUMB[436][2] ) );
  FADDER S1_435_0 ( .CIN(\ab[435][0] ), .IN0(\CARRYB[434][0] ), .IN1(
        \SUMB[434][1] ), .COUT(\CARRYB[435][0] ), .SUM(PRODUCT[435]) );
  FADDER S2_435_1 ( .CIN(\ab[435][1] ), .IN0(\CARRYB[434][1] ), .IN1(
        \SUMB[434][2] ), .COUT(\CARRYB[435][1] ), .SUM(\SUMB[435][1] ) );
  FADDER S3_435_2 ( .CIN(\ab[435][2] ), .IN0(\CARRYB[434][2] ), .IN1(
        \ab[434][3] ), .COUT(\CARRYB[435][2] ), .SUM(\SUMB[435][2] ) );
  FADDER S1_434_0 ( .CIN(\ab[434][0] ), .IN0(\CARRYB[433][0] ), .IN1(
        \SUMB[433][1] ), .COUT(\CARRYB[434][0] ), .SUM(PRODUCT[434]) );
  FADDER S2_434_1 ( .CIN(\ab[434][1] ), .IN0(\CARRYB[433][1] ), .IN1(
        \SUMB[433][2] ), .COUT(\CARRYB[434][1] ), .SUM(\SUMB[434][1] ) );
  FADDER S3_434_2 ( .CIN(\ab[434][2] ), .IN0(\CARRYB[433][2] ), .IN1(
        \ab[433][3] ), .COUT(\CARRYB[434][2] ), .SUM(\SUMB[434][2] ) );
  FADDER S1_433_0 ( .CIN(\ab[433][0] ), .IN0(\CARRYB[432][0] ), .IN1(
        \SUMB[432][1] ), .COUT(\CARRYB[433][0] ), .SUM(PRODUCT[433]) );
  FADDER S2_433_1 ( .CIN(\ab[433][1] ), .IN0(\CARRYB[432][1] ), .IN1(
        \SUMB[432][2] ), .COUT(\CARRYB[433][1] ), .SUM(\SUMB[433][1] ) );
  FADDER S3_433_2 ( .CIN(\ab[433][2] ), .IN0(\CARRYB[432][2] ), .IN1(
        \ab[432][3] ), .COUT(\CARRYB[433][2] ), .SUM(\SUMB[433][2] ) );
  FADDER S1_432_0 ( .CIN(\ab[432][0] ), .IN0(\CARRYB[431][0] ), .IN1(
        \SUMB[431][1] ), .COUT(\CARRYB[432][0] ), .SUM(PRODUCT[432]) );
  FADDER S2_432_1 ( .CIN(\ab[432][1] ), .IN0(\CARRYB[431][1] ), .IN1(
        \SUMB[431][2] ), .COUT(\CARRYB[432][1] ), .SUM(\SUMB[432][1] ) );
  FADDER S3_432_2 ( .CIN(\ab[432][2] ), .IN0(\CARRYB[431][2] ), .IN1(
        \ab[431][3] ), .COUT(\CARRYB[432][2] ), .SUM(\SUMB[432][2] ) );
  FADDER S1_431_0 ( .CIN(\ab[431][0] ), .IN0(\CARRYB[430][0] ), .IN1(
        \SUMB[430][1] ), .COUT(\CARRYB[431][0] ), .SUM(PRODUCT[431]) );
  FADDER S2_431_1 ( .CIN(\ab[431][1] ), .IN0(\CARRYB[430][1] ), .IN1(
        \SUMB[430][2] ), .COUT(\CARRYB[431][1] ), .SUM(\SUMB[431][1] ) );
  FADDER S3_431_2 ( .CIN(\ab[431][2] ), .IN0(\CARRYB[430][2] ), .IN1(
        \ab[430][3] ), .COUT(\CARRYB[431][2] ), .SUM(\SUMB[431][2] ) );
  FADDER S1_430_0 ( .CIN(\ab[430][0] ), .IN0(\CARRYB[429][0] ), .IN1(
        \SUMB[429][1] ), .COUT(\CARRYB[430][0] ), .SUM(PRODUCT[430]) );
  FADDER S2_430_1 ( .CIN(\ab[430][1] ), .IN0(\CARRYB[429][1] ), .IN1(
        \SUMB[429][2] ), .COUT(\CARRYB[430][1] ), .SUM(\SUMB[430][1] ) );
  FADDER S3_430_2 ( .CIN(\ab[430][2] ), .IN0(\CARRYB[429][2] ), .IN1(
        \ab[429][3] ), .COUT(\CARRYB[430][2] ), .SUM(\SUMB[430][2] ) );
  FADDER S1_429_0 ( .CIN(\ab[429][0] ), .IN0(\CARRYB[428][0] ), .IN1(
        \SUMB[428][1] ), .COUT(\CARRYB[429][0] ), .SUM(PRODUCT[429]) );
  FADDER S2_429_1 ( .CIN(\ab[429][1] ), .IN0(\CARRYB[428][1] ), .IN1(
        \SUMB[428][2] ), .COUT(\CARRYB[429][1] ), .SUM(\SUMB[429][1] ) );
  FADDER S3_429_2 ( .CIN(\ab[429][2] ), .IN0(\CARRYB[428][2] ), .IN1(
        \ab[428][3] ), .COUT(\CARRYB[429][2] ), .SUM(\SUMB[429][2] ) );
  FADDER S1_428_0 ( .CIN(\ab[428][0] ), .IN0(\CARRYB[427][0] ), .IN1(
        \SUMB[427][1] ), .COUT(\CARRYB[428][0] ), .SUM(PRODUCT[428]) );
  FADDER S2_428_1 ( .CIN(\ab[428][1] ), .IN0(\CARRYB[427][1] ), .IN1(
        \SUMB[427][2] ), .COUT(\CARRYB[428][1] ), .SUM(\SUMB[428][1] ) );
  FADDER S3_428_2 ( .CIN(\ab[428][2] ), .IN0(\CARRYB[427][2] ), .IN1(
        \ab[427][3] ), .COUT(\CARRYB[428][2] ), .SUM(\SUMB[428][2] ) );
  FADDER S1_427_0 ( .CIN(\ab[427][0] ), .IN0(\CARRYB[426][0] ), .IN1(
        \SUMB[426][1] ), .COUT(\CARRYB[427][0] ), .SUM(PRODUCT[427]) );
  FADDER S2_427_1 ( .CIN(\ab[427][1] ), .IN0(\CARRYB[426][1] ), .IN1(
        \SUMB[426][2] ), .COUT(\CARRYB[427][1] ), .SUM(\SUMB[427][1] ) );
  FADDER S3_427_2 ( .CIN(\ab[427][2] ), .IN0(\CARRYB[426][2] ), .IN1(
        \ab[426][3] ), .COUT(\CARRYB[427][2] ), .SUM(\SUMB[427][2] ) );
  FADDER S1_426_0 ( .CIN(\ab[426][0] ), .IN0(\CARRYB[425][0] ), .IN1(
        \SUMB[425][1] ), .COUT(\CARRYB[426][0] ), .SUM(PRODUCT[426]) );
  FADDER S2_426_1 ( .CIN(\ab[426][1] ), .IN0(\CARRYB[425][1] ), .IN1(
        \SUMB[425][2] ), .COUT(\CARRYB[426][1] ), .SUM(\SUMB[426][1] ) );
  FADDER S3_426_2 ( .CIN(\ab[426][2] ), .IN0(\CARRYB[425][2] ), .IN1(
        \ab[425][3] ), .COUT(\CARRYB[426][2] ), .SUM(\SUMB[426][2] ) );
  FADDER S1_425_0 ( .CIN(\ab[425][0] ), .IN0(\CARRYB[424][0] ), .IN1(
        \SUMB[424][1] ), .COUT(\CARRYB[425][0] ), .SUM(PRODUCT[425]) );
  FADDER S2_425_1 ( .CIN(\ab[425][1] ), .IN0(\CARRYB[424][1] ), .IN1(
        \SUMB[424][2] ), .COUT(\CARRYB[425][1] ), .SUM(\SUMB[425][1] ) );
  FADDER S3_425_2 ( .CIN(\ab[425][2] ), .IN0(\CARRYB[424][2] ), .IN1(
        \ab[424][3] ), .COUT(\CARRYB[425][2] ), .SUM(\SUMB[425][2] ) );
  FADDER S1_424_0 ( .CIN(\ab[424][0] ), .IN0(\CARRYB[423][0] ), .IN1(
        \SUMB[423][1] ), .COUT(\CARRYB[424][0] ), .SUM(PRODUCT[424]) );
  FADDER S2_424_1 ( .CIN(\ab[424][1] ), .IN0(\CARRYB[423][1] ), .IN1(
        \SUMB[423][2] ), .COUT(\CARRYB[424][1] ), .SUM(\SUMB[424][1] ) );
  FADDER S3_424_2 ( .CIN(\ab[424][2] ), .IN0(\CARRYB[423][2] ), .IN1(
        \ab[423][3] ), .COUT(\CARRYB[424][2] ), .SUM(\SUMB[424][2] ) );
  FADDER S1_423_0 ( .CIN(\ab[423][0] ), .IN0(\CARRYB[422][0] ), .IN1(
        \SUMB[422][1] ), .COUT(\CARRYB[423][0] ), .SUM(PRODUCT[423]) );
  FADDER S2_423_1 ( .CIN(\ab[423][1] ), .IN0(\CARRYB[422][1] ), .IN1(
        \SUMB[422][2] ), .COUT(\CARRYB[423][1] ), .SUM(\SUMB[423][1] ) );
  FADDER S3_423_2 ( .CIN(\ab[423][2] ), .IN0(\CARRYB[422][2] ), .IN1(
        \ab[422][3] ), .COUT(\CARRYB[423][2] ), .SUM(\SUMB[423][2] ) );
  FADDER S1_422_0 ( .CIN(\ab[422][0] ), .IN0(\CARRYB[421][0] ), .IN1(
        \SUMB[421][1] ), .COUT(\CARRYB[422][0] ), .SUM(PRODUCT[422]) );
  FADDER S2_422_1 ( .CIN(\ab[422][1] ), .IN0(\CARRYB[421][1] ), .IN1(
        \SUMB[421][2] ), .COUT(\CARRYB[422][1] ), .SUM(\SUMB[422][1] ) );
  FADDER S3_422_2 ( .CIN(\ab[422][2] ), .IN0(\CARRYB[421][2] ), .IN1(
        \ab[421][3] ), .COUT(\CARRYB[422][2] ), .SUM(\SUMB[422][2] ) );
  FADDER S1_421_0 ( .CIN(\ab[421][0] ), .IN0(\CARRYB[420][0] ), .IN1(
        \SUMB[420][1] ), .COUT(\CARRYB[421][0] ), .SUM(PRODUCT[421]) );
  FADDER S2_421_1 ( .CIN(\ab[421][1] ), .IN0(\CARRYB[420][1] ), .IN1(
        \SUMB[420][2] ), .COUT(\CARRYB[421][1] ), .SUM(\SUMB[421][1] ) );
  FADDER S3_421_2 ( .CIN(\ab[421][2] ), .IN0(\CARRYB[420][2] ), .IN1(
        \ab[420][3] ), .COUT(\CARRYB[421][2] ), .SUM(\SUMB[421][2] ) );
  FADDER S1_420_0 ( .CIN(\ab[420][0] ), .IN0(\CARRYB[419][0] ), .IN1(
        \SUMB[419][1] ), .COUT(\CARRYB[420][0] ), .SUM(PRODUCT[420]) );
  FADDER S2_420_1 ( .CIN(\ab[420][1] ), .IN0(\CARRYB[419][1] ), .IN1(
        \SUMB[419][2] ), .COUT(\CARRYB[420][1] ), .SUM(\SUMB[420][1] ) );
  FADDER S3_420_2 ( .CIN(\ab[420][2] ), .IN0(\CARRYB[419][2] ), .IN1(
        \ab[419][3] ), .COUT(\CARRYB[420][2] ), .SUM(\SUMB[420][2] ) );
  FADDER S1_419_0 ( .CIN(\ab[419][0] ), .IN0(\CARRYB[418][0] ), .IN1(
        \SUMB[418][1] ), .COUT(\CARRYB[419][0] ), .SUM(PRODUCT[419]) );
  FADDER S2_419_1 ( .CIN(\ab[419][1] ), .IN0(\CARRYB[418][1] ), .IN1(
        \SUMB[418][2] ), .COUT(\CARRYB[419][1] ), .SUM(\SUMB[419][1] ) );
  FADDER S3_419_2 ( .CIN(\ab[419][2] ), .IN0(\CARRYB[418][2] ), .IN1(
        \ab[418][3] ), .COUT(\CARRYB[419][2] ), .SUM(\SUMB[419][2] ) );
  FADDER S1_418_0 ( .CIN(\ab[418][0] ), .IN0(\CARRYB[417][0] ), .IN1(
        \SUMB[417][1] ), .COUT(\CARRYB[418][0] ), .SUM(PRODUCT[418]) );
  FADDER S2_418_1 ( .CIN(\ab[418][1] ), .IN0(\CARRYB[417][1] ), .IN1(
        \SUMB[417][2] ), .COUT(\CARRYB[418][1] ), .SUM(\SUMB[418][1] ) );
  FADDER S3_418_2 ( .CIN(\ab[418][2] ), .IN0(\CARRYB[417][2] ), .IN1(
        \ab[417][3] ), .COUT(\CARRYB[418][2] ), .SUM(\SUMB[418][2] ) );
  FADDER S1_417_0 ( .CIN(\ab[417][0] ), .IN0(\CARRYB[416][0] ), .IN1(
        \SUMB[416][1] ), .COUT(\CARRYB[417][0] ), .SUM(PRODUCT[417]) );
  FADDER S2_417_1 ( .CIN(\ab[417][1] ), .IN0(\CARRYB[416][1] ), .IN1(
        \SUMB[416][2] ), .COUT(\CARRYB[417][1] ), .SUM(\SUMB[417][1] ) );
  FADDER S3_417_2 ( .CIN(\ab[417][2] ), .IN0(\CARRYB[416][2] ), .IN1(
        \ab[416][3] ), .COUT(\CARRYB[417][2] ), .SUM(\SUMB[417][2] ) );
  FADDER S1_416_0 ( .CIN(\ab[416][0] ), .IN0(\CARRYB[415][0] ), .IN1(
        \SUMB[415][1] ), .COUT(\CARRYB[416][0] ), .SUM(PRODUCT[416]) );
  FADDER S2_416_1 ( .CIN(\ab[416][1] ), .IN0(\CARRYB[415][1] ), .IN1(
        \SUMB[415][2] ), .COUT(\CARRYB[416][1] ), .SUM(\SUMB[416][1] ) );
  FADDER S3_416_2 ( .CIN(\ab[416][2] ), .IN0(\CARRYB[415][2] ), .IN1(
        \ab[415][3] ), .COUT(\CARRYB[416][2] ), .SUM(\SUMB[416][2] ) );
  FADDER S1_415_0 ( .CIN(\ab[415][0] ), .IN0(\CARRYB[414][0] ), .IN1(
        \SUMB[414][1] ), .COUT(\CARRYB[415][0] ), .SUM(PRODUCT[415]) );
  FADDER S2_415_1 ( .CIN(\ab[415][1] ), .IN0(\CARRYB[414][1] ), .IN1(
        \SUMB[414][2] ), .COUT(\CARRYB[415][1] ), .SUM(\SUMB[415][1] ) );
  FADDER S3_415_2 ( .CIN(\ab[415][2] ), .IN0(\CARRYB[414][2] ), .IN1(
        \ab[414][3] ), .COUT(\CARRYB[415][2] ), .SUM(\SUMB[415][2] ) );
  FADDER S1_414_0 ( .CIN(\ab[414][0] ), .IN0(\CARRYB[413][0] ), .IN1(
        \SUMB[413][1] ), .COUT(\CARRYB[414][0] ), .SUM(PRODUCT[414]) );
  FADDER S2_414_1 ( .CIN(\ab[414][1] ), .IN0(\CARRYB[413][1] ), .IN1(
        \SUMB[413][2] ), .COUT(\CARRYB[414][1] ), .SUM(\SUMB[414][1] ) );
  FADDER S3_414_2 ( .CIN(\ab[414][2] ), .IN0(\CARRYB[413][2] ), .IN1(
        \ab[413][3] ), .COUT(\CARRYB[414][2] ), .SUM(\SUMB[414][2] ) );
  FADDER S1_413_0 ( .CIN(\ab[413][0] ), .IN0(\CARRYB[412][0] ), .IN1(
        \SUMB[412][1] ), .COUT(\CARRYB[413][0] ), .SUM(PRODUCT[413]) );
  FADDER S2_413_1 ( .CIN(\ab[413][1] ), .IN0(\CARRYB[412][1] ), .IN1(
        \SUMB[412][2] ), .COUT(\CARRYB[413][1] ), .SUM(\SUMB[413][1] ) );
  FADDER S3_413_2 ( .CIN(\ab[413][2] ), .IN0(\CARRYB[412][2] ), .IN1(
        \ab[412][3] ), .COUT(\CARRYB[413][2] ), .SUM(\SUMB[413][2] ) );
  FADDER S1_412_0 ( .CIN(\ab[412][0] ), .IN0(\CARRYB[411][0] ), .IN1(
        \SUMB[411][1] ), .COUT(\CARRYB[412][0] ), .SUM(PRODUCT[412]) );
  FADDER S2_412_1 ( .CIN(\ab[412][1] ), .IN0(\CARRYB[411][1] ), .IN1(
        \SUMB[411][2] ), .COUT(\CARRYB[412][1] ), .SUM(\SUMB[412][1] ) );
  FADDER S3_412_2 ( .CIN(\ab[412][2] ), .IN0(\CARRYB[411][2] ), .IN1(
        \ab[411][3] ), .COUT(\CARRYB[412][2] ), .SUM(\SUMB[412][2] ) );
  FADDER S1_411_0 ( .CIN(\ab[411][0] ), .IN0(\CARRYB[410][0] ), .IN1(
        \SUMB[410][1] ), .COUT(\CARRYB[411][0] ), .SUM(PRODUCT[411]) );
  FADDER S2_411_1 ( .CIN(\ab[411][1] ), .IN0(\CARRYB[410][1] ), .IN1(
        \SUMB[410][2] ), .COUT(\CARRYB[411][1] ), .SUM(\SUMB[411][1] ) );
  FADDER S3_411_2 ( .CIN(\ab[411][2] ), .IN0(\CARRYB[410][2] ), .IN1(
        \ab[410][3] ), .COUT(\CARRYB[411][2] ), .SUM(\SUMB[411][2] ) );
  FADDER S1_410_0 ( .CIN(\ab[410][0] ), .IN0(\CARRYB[409][0] ), .IN1(
        \SUMB[409][1] ), .COUT(\CARRYB[410][0] ), .SUM(PRODUCT[410]) );
  FADDER S2_410_1 ( .CIN(\ab[410][1] ), .IN0(\CARRYB[409][1] ), .IN1(
        \SUMB[409][2] ), .COUT(\CARRYB[410][1] ), .SUM(\SUMB[410][1] ) );
  FADDER S3_410_2 ( .CIN(\ab[410][2] ), .IN0(\CARRYB[409][2] ), .IN1(
        \ab[409][3] ), .COUT(\CARRYB[410][2] ), .SUM(\SUMB[410][2] ) );
  FADDER S1_409_0 ( .CIN(\ab[409][0] ), .IN0(\CARRYB[408][0] ), .IN1(
        \SUMB[408][1] ), .COUT(\CARRYB[409][0] ), .SUM(PRODUCT[409]) );
  FADDER S2_409_1 ( .CIN(\ab[409][1] ), .IN0(\CARRYB[408][1] ), .IN1(
        \SUMB[408][2] ), .COUT(\CARRYB[409][1] ), .SUM(\SUMB[409][1] ) );
  FADDER S3_409_2 ( .CIN(\ab[409][2] ), .IN0(\CARRYB[408][2] ), .IN1(
        \ab[408][3] ), .COUT(\CARRYB[409][2] ), .SUM(\SUMB[409][2] ) );
  FADDER S1_408_0 ( .CIN(\ab[408][0] ), .IN0(\CARRYB[407][0] ), .IN1(
        \SUMB[407][1] ), .COUT(\CARRYB[408][0] ), .SUM(PRODUCT[408]) );
  FADDER S2_408_1 ( .CIN(\ab[408][1] ), .IN0(\CARRYB[407][1] ), .IN1(
        \SUMB[407][2] ), .COUT(\CARRYB[408][1] ), .SUM(\SUMB[408][1] ) );
  FADDER S3_408_2 ( .CIN(\ab[408][2] ), .IN0(\CARRYB[407][2] ), .IN1(
        \ab[407][3] ), .COUT(\CARRYB[408][2] ), .SUM(\SUMB[408][2] ) );
  FADDER S1_407_0 ( .CIN(\ab[407][0] ), .IN0(\CARRYB[406][0] ), .IN1(
        \SUMB[406][1] ), .COUT(\CARRYB[407][0] ), .SUM(PRODUCT[407]) );
  FADDER S2_407_1 ( .CIN(\ab[407][1] ), .IN0(\CARRYB[406][1] ), .IN1(
        \SUMB[406][2] ), .COUT(\CARRYB[407][1] ), .SUM(\SUMB[407][1] ) );
  FADDER S3_407_2 ( .CIN(\ab[407][2] ), .IN0(\CARRYB[406][2] ), .IN1(
        \ab[406][3] ), .COUT(\CARRYB[407][2] ), .SUM(\SUMB[407][2] ) );
  FADDER S1_406_0 ( .CIN(\ab[406][0] ), .IN0(\CARRYB[405][0] ), .IN1(
        \SUMB[405][1] ), .COUT(\CARRYB[406][0] ), .SUM(PRODUCT[406]) );
  FADDER S2_406_1 ( .CIN(\ab[406][1] ), .IN0(\CARRYB[405][1] ), .IN1(
        \SUMB[405][2] ), .COUT(\CARRYB[406][1] ), .SUM(\SUMB[406][1] ) );
  FADDER S3_406_2 ( .CIN(\ab[406][2] ), .IN0(\CARRYB[405][2] ), .IN1(
        \ab[405][3] ), .COUT(\CARRYB[406][2] ), .SUM(\SUMB[406][2] ) );
  FADDER S1_405_0 ( .CIN(\ab[405][0] ), .IN0(\CARRYB[404][0] ), .IN1(
        \SUMB[404][1] ), .COUT(\CARRYB[405][0] ), .SUM(PRODUCT[405]) );
  FADDER S2_405_1 ( .CIN(\ab[405][1] ), .IN0(\CARRYB[404][1] ), .IN1(
        \SUMB[404][2] ), .COUT(\CARRYB[405][1] ), .SUM(\SUMB[405][1] ) );
  FADDER S3_405_2 ( .CIN(\ab[405][2] ), .IN0(\CARRYB[404][2] ), .IN1(
        \ab[404][3] ), .COUT(\CARRYB[405][2] ), .SUM(\SUMB[405][2] ) );
  FADDER S1_404_0 ( .CIN(\ab[404][0] ), .IN0(\CARRYB[403][0] ), .IN1(
        \SUMB[403][1] ), .COUT(\CARRYB[404][0] ), .SUM(PRODUCT[404]) );
  FADDER S2_404_1 ( .CIN(\ab[404][1] ), .IN0(\CARRYB[403][1] ), .IN1(
        \SUMB[403][2] ), .COUT(\CARRYB[404][1] ), .SUM(\SUMB[404][1] ) );
  FADDER S3_404_2 ( .CIN(\ab[404][2] ), .IN0(\CARRYB[403][2] ), .IN1(
        \ab[403][3] ), .COUT(\CARRYB[404][2] ), .SUM(\SUMB[404][2] ) );
  FADDER S1_403_0 ( .CIN(\ab[403][0] ), .IN0(\CARRYB[402][0] ), .IN1(
        \SUMB[402][1] ), .COUT(\CARRYB[403][0] ), .SUM(PRODUCT[403]) );
  FADDER S2_403_1 ( .CIN(\ab[403][1] ), .IN0(\CARRYB[402][1] ), .IN1(
        \SUMB[402][2] ), .COUT(\CARRYB[403][1] ), .SUM(\SUMB[403][1] ) );
  FADDER S3_403_2 ( .CIN(\ab[403][2] ), .IN0(\CARRYB[402][2] ), .IN1(
        \ab[402][3] ), .COUT(\CARRYB[403][2] ), .SUM(\SUMB[403][2] ) );
  FADDER S1_402_0 ( .CIN(\ab[402][0] ), .IN0(\CARRYB[401][0] ), .IN1(
        \SUMB[401][1] ), .COUT(\CARRYB[402][0] ), .SUM(PRODUCT[402]) );
  FADDER S2_402_1 ( .CIN(\ab[402][1] ), .IN0(\CARRYB[401][1] ), .IN1(
        \SUMB[401][2] ), .COUT(\CARRYB[402][1] ), .SUM(\SUMB[402][1] ) );
  FADDER S3_402_2 ( .CIN(\ab[402][2] ), .IN0(\CARRYB[401][2] ), .IN1(
        \ab[401][3] ), .COUT(\CARRYB[402][2] ), .SUM(\SUMB[402][2] ) );
  FADDER S1_401_0 ( .CIN(\ab[401][0] ), .IN0(\CARRYB[400][0] ), .IN1(
        \SUMB[400][1] ), .COUT(\CARRYB[401][0] ), .SUM(PRODUCT[401]) );
  FADDER S2_401_1 ( .CIN(\ab[401][1] ), .IN0(\CARRYB[400][1] ), .IN1(
        \SUMB[400][2] ), .COUT(\CARRYB[401][1] ), .SUM(\SUMB[401][1] ) );
  FADDER S3_401_2 ( .CIN(\ab[401][2] ), .IN0(\CARRYB[400][2] ), .IN1(
        \ab[400][3] ), .COUT(\CARRYB[401][2] ), .SUM(\SUMB[401][2] ) );
  FADDER S1_400_0 ( .CIN(\ab[400][0] ), .IN0(\CARRYB[399][0] ), .IN1(
        \SUMB[399][1] ), .COUT(\CARRYB[400][0] ), .SUM(PRODUCT[400]) );
  FADDER S2_400_1 ( .CIN(\ab[400][1] ), .IN0(\CARRYB[399][1] ), .IN1(
        \SUMB[399][2] ), .COUT(\CARRYB[400][1] ), .SUM(\SUMB[400][1] ) );
  FADDER S3_400_2 ( .CIN(\ab[400][2] ), .IN0(\CARRYB[399][2] ), .IN1(
        \ab[399][3] ), .COUT(\CARRYB[400][2] ), .SUM(\SUMB[400][2] ) );
  FADDER S1_399_0 ( .CIN(\ab[399][0] ), .IN0(\CARRYB[398][0] ), .IN1(
        \SUMB[398][1] ), .COUT(\CARRYB[399][0] ), .SUM(PRODUCT[399]) );
  FADDER S2_399_1 ( .CIN(\ab[399][1] ), .IN0(\CARRYB[398][1] ), .IN1(
        \SUMB[398][2] ), .COUT(\CARRYB[399][1] ), .SUM(\SUMB[399][1] ) );
  FADDER S3_399_2 ( .CIN(\ab[399][2] ), .IN0(\CARRYB[398][2] ), .IN1(
        \ab[398][3] ), .COUT(\CARRYB[399][2] ), .SUM(\SUMB[399][2] ) );
  FADDER S1_398_0 ( .CIN(\ab[398][0] ), .IN0(\CARRYB[397][0] ), .IN1(
        \SUMB[397][1] ), .COUT(\CARRYB[398][0] ), .SUM(PRODUCT[398]) );
  FADDER S2_398_1 ( .CIN(\ab[398][1] ), .IN0(\CARRYB[397][1] ), .IN1(
        \SUMB[397][2] ), .COUT(\CARRYB[398][1] ), .SUM(\SUMB[398][1] ) );
  FADDER S3_398_2 ( .CIN(\ab[398][2] ), .IN0(\CARRYB[397][2] ), .IN1(
        \ab[397][3] ), .COUT(\CARRYB[398][2] ), .SUM(\SUMB[398][2] ) );
  FADDER S1_397_0 ( .CIN(\ab[397][0] ), .IN0(\CARRYB[396][0] ), .IN1(
        \SUMB[396][1] ), .COUT(\CARRYB[397][0] ), .SUM(PRODUCT[397]) );
  FADDER S2_397_1 ( .CIN(\ab[397][1] ), .IN0(\CARRYB[396][1] ), .IN1(
        \SUMB[396][2] ), .COUT(\CARRYB[397][1] ), .SUM(\SUMB[397][1] ) );
  FADDER S3_397_2 ( .CIN(\ab[397][2] ), .IN0(\CARRYB[396][2] ), .IN1(
        \ab[396][3] ), .COUT(\CARRYB[397][2] ), .SUM(\SUMB[397][2] ) );
  FADDER S1_396_0 ( .CIN(\ab[396][0] ), .IN0(\CARRYB[395][0] ), .IN1(
        \SUMB[395][1] ), .COUT(\CARRYB[396][0] ), .SUM(PRODUCT[396]) );
  FADDER S2_396_1 ( .CIN(\ab[396][1] ), .IN0(\CARRYB[395][1] ), .IN1(
        \SUMB[395][2] ), .COUT(\CARRYB[396][1] ), .SUM(\SUMB[396][1] ) );
  FADDER S3_396_2 ( .CIN(\ab[396][2] ), .IN0(\CARRYB[395][2] ), .IN1(
        \ab[395][3] ), .COUT(\CARRYB[396][2] ), .SUM(\SUMB[396][2] ) );
  FADDER S1_395_0 ( .CIN(\ab[395][0] ), .IN0(\CARRYB[394][0] ), .IN1(
        \SUMB[394][1] ), .COUT(\CARRYB[395][0] ), .SUM(PRODUCT[395]) );
  FADDER S2_395_1 ( .CIN(\ab[395][1] ), .IN0(\CARRYB[394][1] ), .IN1(
        \SUMB[394][2] ), .COUT(\CARRYB[395][1] ), .SUM(\SUMB[395][1] ) );
  FADDER S3_395_2 ( .CIN(\ab[395][2] ), .IN0(\CARRYB[394][2] ), .IN1(
        \ab[394][3] ), .COUT(\CARRYB[395][2] ), .SUM(\SUMB[395][2] ) );
  FADDER S1_394_0 ( .CIN(\ab[394][0] ), .IN0(\CARRYB[393][0] ), .IN1(
        \SUMB[393][1] ), .COUT(\CARRYB[394][0] ), .SUM(PRODUCT[394]) );
  FADDER S2_394_1 ( .CIN(\ab[394][1] ), .IN0(\CARRYB[393][1] ), .IN1(
        \SUMB[393][2] ), .COUT(\CARRYB[394][1] ), .SUM(\SUMB[394][1] ) );
  FADDER S3_394_2 ( .CIN(\ab[394][2] ), .IN0(\CARRYB[393][2] ), .IN1(
        \ab[393][3] ), .COUT(\CARRYB[394][2] ), .SUM(\SUMB[394][2] ) );
  FADDER S1_393_0 ( .CIN(\ab[393][0] ), .IN0(\CARRYB[392][0] ), .IN1(
        \SUMB[392][1] ), .COUT(\CARRYB[393][0] ), .SUM(PRODUCT[393]) );
  FADDER S2_393_1 ( .CIN(\ab[393][1] ), .IN0(\CARRYB[392][1] ), .IN1(
        \SUMB[392][2] ), .COUT(\CARRYB[393][1] ), .SUM(\SUMB[393][1] ) );
  FADDER S3_393_2 ( .CIN(\ab[393][2] ), .IN0(\CARRYB[392][2] ), .IN1(
        \ab[392][3] ), .COUT(\CARRYB[393][2] ), .SUM(\SUMB[393][2] ) );
  FADDER S1_392_0 ( .CIN(\ab[392][0] ), .IN0(\CARRYB[391][0] ), .IN1(
        \SUMB[391][1] ), .COUT(\CARRYB[392][0] ), .SUM(PRODUCT[392]) );
  FADDER S2_392_1 ( .CIN(\ab[392][1] ), .IN0(\CARRYB[391][1] ), .IN1(
        \SUMB[391][2] ), .COUT(\CARRYB[392][1] ), .SUM(\SUMB[392][1] ) );
  FADDER S3_392_2 ( .CIN(\ab[392][2] ), .IN0(\CARRYB[391][2] ), .IN1(
        \ab[391][3] ), .COUT(\CARRYB[392][2] ), .SUM(\SUMB[392][2] ) );
  FADDER S1_391_0 ( .CIN(\ab[391][0] ), .IN0(\CARRYB[390][0] ), .IN1(
        \SUMB[390][1] ), .COUT(\CARRYB[391][0] ), .SUM(PRODUCT[391]) );
  FADDER S2_391_1 ( .CIN(\ab[391][1] ), .IN0(\CARRYB[390][1] ), .IN1(
        \SUMB[390][2] ), .COUT(\CARRYB[391][1] ), .SUM(\SUMB[391][1] ) );
  FADDER S3_391_2 ( .CIN(\ab[391][2] ), .IN0(\CARRYB[390][2] ), .IN1(
        \ab[390][3] ), .COUT(\CARRYB[391][2] ), .SUM(\SUMB[391][2] ) );
  FADDER S1_390_0 ( .CIN(\ab[390][0] ), .IN0(\CARRYB[389][0] ), .IN1(
        \SUMB[389][1] ), .COUT(\CARRYB[390][0] ), .SUM(PRODUCT[390]) );
  FADDER S2_390_1 ( .CIN(\ab[390][1] ), .IN0(\CARRYB[389][1] ), .IN1(
        \SUMB[389][2] ), .COUT(\CARRYB[390][1] ), .SUM(\SUMB[390][1] ) );
  FADDER S3_390_2 ( .CIN(\ab[390][2] ), .IN0(\CARRYB[389][2] ), .IN1(
        \ab[389][3] ), .COUT(\CARRYB[390][2] ), .SUM(\SUMB[390][2] ) );
  FADDER S1_389_0 ( .CIN(\ab[389][0] ), .IN0(\CARRYB[388][0] ), .IN1(
        \SUMB[388][1] ), .COUT(\CARRYB[389][0] ), .SUM(PRODUCT[389]) );
  FADDER S2_389_1 ( .CIN(\ab[389][1] ), .IN0(\CARRYB[388][1] ), .IN1(
        \SUMB[388][2] ), .COUT(\CARRYB[389][1] ), .SUM(\SUMB[389][1] ) );
  FADDER S3_389_2 ( .CIN(\ab[389][2] ), .IN0(\CARRYB[388][2] ), .IN1(
        \ab[388][3] ), .COUT(\CARRYB[389][2] ), .SUM(\SUMB[389][2] ) );
  FADDER S1_388_0 ( .CIN(\ab[388][0] ), .IN0(\CARRYB[387][0] ), .IN1(
        \SUMB[387][1] ), .COUT(\CARRYB[388][0] ), .SUM(PRODUCT[388]) );
  FADDER S2_388_1 ( .CIN(\ab[388][1] ), .IN0(\CARRYB[387][1] ), .IN1(
        \SUMB[387][2] ), .COUT(\CARRYB[388][1] ), .SUM(\SUMB[388][1] ) );
  FADDER S3_388_2 ( .CIN(\ab[388][2] ), .IN0(\CARRYB[387][2] ), .IN1(
        \ab[387][3] ), .COUT(\CARRYB[388][2] ), .SUM(\SUMB[388][2] ) );
  FADDER S1_387_0 ( .CIN(\ab[387][0] ), .IN0(\CARRYB[386][0] ), .IN1(
        \SUMB[386][1] ), .COUT(\CARRYB[387][0] ), .SUM(PRODUCT[387]) );
  FADDER S2_387_1 ( .CIN(\ab[387][1] ), .IN0(\CARRYB[386][1] ), .IN1(
        \SUMB[386][2] ), .COUT(\CARRYB[387][1] ), .SUM(\SUMB[387][1] ) );
  FADDER S3_387_2 ( .CIN(\ab[387][2] ), .IN0(\CARRYB[386][2] ), .IN1(
        \ab[386][3] ), .COUT(\CARRYB[387][2] ), .SUM(\SUMB[387][2] ) );
  FADDER S1_386_0 ( .CIN(\ab[386][0] ), .IN0(\CARRYB[385][0] ), .IN1(
        \SUMB[385][1] ), .COUT(\CARRYB[386][0] ), .SUM(PRODUCT[386]) );
  FADDER S2_386_1 ( .CIN(\ab[386][1] ), .IN0(\CARRYB[385][1] ), .IN1(
        \SUMB[385][2] ), .COUT(\CARRYB[386][1] ), .SUM(\SUMB[386][1] ) );
  FADDER S3_386_2 ( .CIN(\ab[386][2] ), .IN0(\CARRYB[385][2] ), .IN1(
        \ab[385][3] ), .COUT(\CARRYB[386][2] ), .SUM(\SUMB[386][2] ) );
  FADDER S1_385_0 ( .CIN(\ab[385][0] ), .IN0(\CARRYB[384][0] ), .IN1(
        \SUMB[384][1] ), .COUT(\CARRYB[385][0] ), .SUM(PRODUCT[385]) );
  FADDER S2_385_1 ( .CIN(\ab[385][1] ), .IN0(\CARRYB[384][1] ), .IN1(
        \SUMB[384][2] ), .COUT(\CARRYB[385][1] ), .SUM(\SUMB[385][1] ) );
  FADDER S3_385_2 ( .CIN(\ab[385][2] ), .IN0(\CARRYB[384][2] ), .IN1(
        \ab[384][3] ), .COUT(\CARRYB[385][2] ), .SUM(\SUMB[385][2] ) );
  FADDER S1_384_0 ( .CIN(\ab[384][0] ), .IN0(\CARRYB[383][0] ), .IN1(
        \SUMB[383][1] ), .COUT(\CARRYB[384][0] ), .SUM(PRODUCT[384]) );
  FADDER S2_384_1 ( .CIN(\ab[384][1] ), .IN0(\CARRYB[383][1] ), .IN1(
        \SUMB[383][2] ), .COUT(\CARRYB[384][1] ), .SUM(\SUMB[384][1] ) );
  FADDER S3_384_2 ( .CIN(\ab[384][2] ), .IN0(\CARRYB[383][2] ), .IN1(
        \ab[383][3] ), .COUT(\CARRYB[384][2] ), .SUM(\SUMB[384][2] ) );
  FADDER S1_383_0 ( .CIN(\ab[383][0] ), .IN0(\CARRYB[382][0] ), .IN1(
        \SUMB[382][1] ), .COUT(\CARRYB[383][0] ), .SUM(PRODUCT[383]) );
  FADDER S2_383_1 ( .CIN(\ab[383][1] ), .IN0(\CARRYB[382][1] ), .IN1(
        \SUMB[382][2] ), .COUT(\CARRYB[383][1] ), .SUM(\SUMB[383][1] ) );
  FADDER S3_383_2 ( .CIN(\ab[383][2] ), .IN0(\CARRYB[382][2] ), .IN1(
        \ab[382][3] ), .COUT(\CARRYB[383][2] ), .SUM(\SUMB[383][2] ) );
  FADDER S1_382_0 ( .CIN(\ab[382][0] ), .IN0(\CARRYB[381][0] ), .IN1(
        \SUMB[381][1] ), .COUT(\CARRYB[382][0] ), .SUM(PRODUCT[382]) );
  FADDER S2_382_1 ( .CIN(\ab[382][1] ), .IN0(\CARRYB[381][1] ), .IN1(
        \SUMB[381][2] ), .COUT(\CARRYB[382][1] ), .SUM(\SUMB[382][1] ) );
  FADDER S3_382_2 ( .CIN(\ab[382][2] ), .IN0(\CARRYB[381][2] ), .IN1(
        \ab[381][3] ), .COUT(\CARRYB[382][2] ), .SUM(\SUMB[382][2] ) );
  FADDER S1_381_0 ( .CIN(\ab[381][0] ), .IN0(\CARRYB[380][0] ), .IN1(
        \SUMB[380][1] ), .COUT(\CARRYB[381][0] ), .SUM(PRODUCT[381]) );
  FADDER S2_381_1 ( .CIN(\ab[381][1] ), .IN0(\CARRYB[380][1] ), .IN1(
        \SUMB[380][2] ), .COUT(\CARRYB[381][1] ), .SUM(\SUMB[381][1] ) );
  FADDER S3_381_2 ( .CIN(\ab[381][2] ), .IN0(\CARRYB[380][2] ), .IN1(
        \ab[380][3] ), .COUT(\CARRYB[381][2] ), .SUM(\SUMB[381][2] ) );
  FADDER S1_380_0 ( .CIN(\ab[380][0] ), .IN0(\CARRYB[379][0] ), .IN1(
        \SUMB[379][1] ), .COUT(\CARRYB[380][0] ), .SUM(PRODUCT[380]) );
  FADDER S2_380_1 ( .CIN(\ab[380][1] ), .IN0(\CARRYB[379][1] ), .IN1(
        \SUMB[379][2] ), .COUT(\CARRYB[380][1] ), .SUM(\SUMB[380][1] ) );
  FADDER S3_380_2 ( .CIN(\ab[380][2] ), .IN0(\CARRYB[379][2] ), .IN1(
        \ab[379][3] ), .COUT(\CARRYB[380][2] ), .SUM(\SUMB[380][2] ) );
  FADDER S1_379_0 ( .CIN(\ab[379][0] ), .IN0(\CARRYB[378][0] ), .IN1(
        \SUMB[378][1] ), .COUT(\CARRYB[379][0] ), .SUM(PRODUCT[379]) );
  FADDER S2_379_1 ( .CIN(\ab[379][1] ), .IN0(\CARRYB[378][1] ), .IN1(
        \SUMB[378][2] ), .COUT(\CARRYB[379][1] ), .SUM(\SUMB[379][1] ) );
  FADDER S3_379_2 ( .CIN(\ab[379][2] ), .IN0(\CARRYB[378][2] ), .IN1(
        \ab[378][3] ), .COUT(\CARRYB[379][2] ), .SUM(\SUMB[379][2] ) );
  FADDER S1_378_0 ( .CIN(\ab[378][0] ), .IN0(\CARRYB[377][0] ), .IN1(
        \SUMB[377][1] ), .COUT(\CARRYB[378][0] ), .SUM(PRODUCT[378]) );
  FADDER S2_378_1 ( .CIN(\ab[378][1] ), .IN0(\CARRYB[377][1] ), .IN1(
        \SUMB[377][2] ), .COUT(\CARRYB[378][1] ), .SUM(\SUMB[378][1] ) );
  FADDER S3_378_2 ( .CIN(\ab[378][2] ), .IN0(\CARRYB[377][2] ), .IN1(
        \ab[377][3] ), .COUT(\CARRYB[378][2] ), .SUM(\SUMB[378][2] ) );
  FADDER S1_377_0 ( .CIN(\ab[377][0] ), .IN0(\CARRYB[376][0] ), .IN1(
        \SUMB[376][1] ), .COUT(\CARRYB[377][0] ), .SUM(PRODUCT[377]) );
  FADDER S2_377_1 ( .CIN(\ab[377][1] ), .IN0(\CARRYB[376][1] ), .IN1(
        \SUMB[376][2] ), .COUT(\CARRYB[377][1] ), .SUM(\SUMB[377][1] ) );
  FADDER S3_377_2 ( .CIN(\ab[377][2] ), .IN0(\CARRYB[376][2] ), .IN1(
        \ab[376][3] ), .COUT(\CARRYB[377][2] ), .SUM(\SUMB[377][2] ) );
  FADDER S1_376_0 ( .CIN(\ab[376][0] ), .IN0(\CARRYB[375][0] ), .IN1(
        \SUMB[375][1] ), .COUT(\CARRYB[376][0] ), .SUM(PRODUCT[376]) );
  FADDER S2_376_1 ( .CIN(\ab[376][1] ), .IN0(\CARRYB[375][1] ), .IN1(
        \SUMB[375][2] ), .COUT(\CARRYB[376][1] ), .SUM(\SUMB[376][1] ) );
  FADDER S3_376_2 ( .CIN(\ab[376][2] ), .IN0(\CARRYB[375][2] ), .IN1(
        \ab[375][3] ), .COUT(\CARRYB[376][2] ), .SUM(\SUMB[376][2] ) );
  FADDER S1_375_0 ( .CIN(\ab[375][0] ), .IN0(\CARRYB[374][0] ), .IN1(
        \SUMB[374][1] ), .COUT(\CARRYB[375][0] ), .SUM(PRODUCT[375]) );
  FADDER S2_375_1 ( .CIN(\ab[375][1] ), .IN0(\CARRYB[374][1] ), .IN1(
        \SUMB[374][2] ), .COUT(\CARRYB[375][1] ), .SUM(\SUMB[375][1] ) );
  FADDER S3_375_2 ( .CIN(\ab[375][2] ), .IN0(\CARRYB[374][2] ), .IN1(
        \ab[374][3] ), .COUT(\CARRYB[375][2] ), .SUM(\SUMB[375][2] ) );
  FADDER S1_374_0 ( .CIN(\ab[374][0] ), .IN0(\CARRYB[373][0] ), .IN1(
        \SUMB[373][1] ), .COUT(\CARRYB[374][0] ), .SUM(PRODUCT[374]) );
  FADDER S2_374_1 ( .CIN(\ab[374][1] ), .IN0(\CARRYB[373][1] ), .IN1(
        \SUMB[373][2] ), .COUT(\CARRYB[374][1] ), .SUM(\SUMB[374][1] ) );
  FADDER S3_374_2 ( .CIN(\ab[374][2] ), .IN0(\CARRYB[373][2] ), .IN1(
        \ab[373][3] ), .COUT(\CARRYB[374][2] ), .SUM(\SUMB[374][2] ) );
  FADDER S1_373_0 ( .CIN(\ab[373][0] ), .IN0(\CARRYB[372][0] ), .IN1(
        \SUMB[372][1] ), .COUT(\CARRYB[373][0] ), .SUM(PRODUCT[373]) );
  FADDER S2_373_1 ( .CIN(\ab[373][1] ), .IN0(\CARRYB[372][1] ), .IN1(
        \SUMB[372][2] ), .COUT(\CARRYB[373][1] ), .SUM(\SUMB[373][1] ) );
  FADDER S3_373_2 ( .CIN(\ab[373][2] ), .IN0(\CARRYB[372][2] ), .IN1(
        \ab[372][3] ), .COUT(\CARRYB[373][2] ), .SUM(\SUMB[373][2] ) );
  FADDER S1_372_0 ( .CIN(\ab[372][0] ), .IN0(\CARRYB[371][0] ), .IN1(
        \SUMB[371][1] ), .COUT(\CARRYB[372][0] ), .SUM(PRODUCT[372]) );
  FADDER S2_372_1 ( .CIN(\ab[372][1] ), .IN0(\CARRYB[371][1] ), .IN1(
        \SUMB[371][2] ), .COUT(\CARRYB[372][1] ), .SUM(\SUMB[372][1] ) );
  FADDER S3_372_2 ( .CIN(\ab[372][2] ), .IN0(\CARRYB[371][2] ), .IN1(
        \ab[371][3] ), .COUT(\CARRYB[372][2] ), .SUM(\SUMB[372][2] ) );
  FADDER S1_371_0 ( .CIN(\ab[371][0] ), .IN0(\CARRYB[370][0] ), .IN1(
        \SUMB[370][1] ), .COUT(\CARRYB[371][0] ), .SUM(PRODUCT[371]) );
  FADDER S2_371_1 ( .CIN(\ab[371][1] ), .IN0(\CARRYB[370][1] ), .IN1(
        \SUMB[370][2] ), .COUT(\CARRYB[371][1] ), .SUM(\SUMB[371][1] ) );
  FADDER S3_371_2 ( .CIN(\ab[371][2] ), .IN0(\CARRYB[370][2] ), .IN1(
        \ab[370][3] ), .COUT(\CARRYB[371][2] ), .SUM(\SUMB[371][2] ) );
  FADDER S1_370_0 ( .CIN(\ab[370][0] ), .IN0(\CARRYB[369][0] ), .IN1(
        \SUMB[369][1] ), .COUT(\CARRYB[370][0] ), .SUM(PRODUCT[370]) );
  FADDER S2_370_1 ( .CIN(\ab[370][1] ), .IN0(\CARRYB[369][1] ), .IN1(
        \SUMB[369][2] ), .COUT(\CARRYB[370][1] ), .SUM(\SUMB[370][1] ) );
  FADDER S3_370_2 ( .CIN(\ab[370][2] ), .IN0(\CARRYB[369][2] ), .IN1(
        \ab[369][3] ), .COUT(\CARRYB[370][2] ), .SUM(\SUMB[370][2] ) );
  FADDER S1_369_0 ( .CIN(\ab[369][0] ), .IN0(\CARRYB[368][0] ), .IN1(
        \SUMB[368][1] ), .COUT(\CARRYB[369][0] ), .SUM(PRODUCT[369]) );
  FADDER S2_369_1 ( .CIN(\ab[369][1] ), .IN0(\CARRYB[368][1] ), .IN1(
        \SUMB[368][2] ), .COUT(\CARRYB[369][1] ), .SUM(\SUMB[369][1] ) );
  FADDER S3_369_2 ( .CIN(\ab[369][2] ), .IN0(\CARRYB[368][2] ), .IN1(
        \ab[368][3] ), .COUT(\CARRYB[369][2] ), .SUM(\SUMB[369][2] ) );
  FADDER S1_368_0 ( .CIN(\ab[368][0] ), .IN0(\CARRYB[367][0] ), .IN1(
        \SUMB[367][1] ), .COUT(\CARRYB[368][0] ), .SUM(PRODUCT[368]) );
  FADDER S2_368_1 ( .CIN(\ab[368][1] ), .IN0(\CARRYB[367][1] ), .IN1(
        \SUMB[367][2] ), .COUT(\CARRYB[368][1] ), .SUM(\SUMB[368][1] ) );
  FADDER S3_368_2 ( .CIN(\ab[368][2] ), .IN0(\CARRYB[367][2] ), .IN1(
        \ab[367][3] ), .COUT(\CARRYB[368][2] ), .SUM(\SUMB[368][2] ) );
  FADDER S1_367_0 ( .CIN(\ab[367][0] ), .IN0(\CARRYB[366][0] ), .IN1(
        \SUMB[366][1] ), .COUT(\CARRYB[367][0] ), .SUM(PRODUCT[367]) );
  FADDER S2_367_1 ( .CIN(\ab[367][1] ), .IN0(\CARRYB[366][1] ), .IN1(
        \SUMB[366][2] ), .COUT(\CARRYB[367][1] ), .SUM(\SUMB[367][1] ) );
  FADDER S3_367_2 ( .CIN(\ab[367][2] ), .IN0(\CARRYB[366][2] ), .IN1(
        \ab[366][3] ), .COUT(\CARRYB[367][2] ), .SUM(\SUMB[367][2] ) );
  FADDER S1_366_0 ( .CIN(\ab[366][0] ), .IN0(\CARRYB[365][0] ), .IN1(
        \SUMB[365][1] ), .COUT(\CARRYB[366][0] ), .SUM(PRODUCT[366]) );
  FADDER S2_366_1 ( .CIN(\ab[366][1] ), .IN0(\CARRYB[365][1] ), .IN1(
        \SUMB[365][2] ), .COUT(\CARRYB[366][1] ), .SUM(\SUMB[366][1] ) );
  FADDER S3_366_2 ( .CIN(\ab[366][2] ), .IN0(\CARRYB[365][2] ), .IN1(
        \ab[365][3] ), .COUT(\CARRYB[366][2] ), .SUM(\SUMB[366][2] ) );
  FADDER S1_365_0 ( .CIN(\ab[365][0] ), .IN0(\CARRYB[364][0] ), .IN1(
        \SUMB[364][1] ), .COUT(\CARRYB[365][0] ), .SUM(PRODUCT[365]) );
  FADDER S2_365_1 ( .CIN(\ab[365][1] ), .IN0(\CARRYB[364][1] ), .IN1(
        \SUMB[364][2] ), .COUT(\CARRYB[365][1] ), .SUM(\SUMB[365][1] ) );
  FADDER S3_365_2 ( .CIN(\ab[365][2] ), .IN0(\CARRYB[364][2] ), .IN1(
        \ab[364][3] ), .COUT(\CARRYB[365][2] ), .SUM(\SUMB[365][2] ) );
  FADDER S1_364_0 ( .CIN(\ab[364][0] ), .IN0(\CARRYB[363][0] ), .IN1(
        \SUMB[363][1] ), .COUT(\CARRYB[364][0] ), .SUM(PRODUCT[364]) );
  FADDER S2_364_1 ( .CIN(\ab[364][1] ), .IN0(\CARRYB[363][1] ), .IN1(
        \SUMB[363][2] ), .COUT(\CARRYB[364][1] ), .SUM(\SUMB[364][1] ) );
  FADDER S3_364_2 ( .CIN(\ab[364][2] ), .IN0(\CARRYB[363][2] ), .IN1(
        \ab[363][3] ), .COUT(\CARRYB[364][2] ), .SUM(\SUMB[364][2] ) );
  FADDER S1_363_0 ( .CIN(\ab[363][0] ), .IN0(\CARRYB[362][0] ), .IN1(
        \SUMB[362][1] ), .COUT(\CARRYB[363][0] ), .SUM(PRODUCT[363]) );
  FADDER S2_363_1 ( .CIN(\ab[363][1] ), .IN0(\CARRYB[362][1] ), .IN1(
        \SUMB[362][2] ), .COUT(\CARRYB[363][1] ), .SUM(\SUMB[363][1] ) );
  FADDER S3_363_2 ( .CIN(\ab[363][2] ), .IN0(\CARRYB[362][2] ), .IN1(
        \ab[362][3] ), .COUT(\CARRYB[363][2] ), .SUM(\SUMB[363][2] ) );
  FADDER S1_362_0 ( .CIN(\ab[362][0] ), .IN0(\CARRYB[361][0] ), .IN1(
        \SUMB[361][1] ), .COUT(\CARRYB[362][0] ), .SUM(PRODUCT[362]) );
  FADDER S2_362_1 ( .CIN(\ab[362][1] ), .IN0(\CARRYB[361][1] ), .IN1(
        \SUMB[361][2] ), .COUT(\CARRYB[362][1] ), .SUM(\SUMB[362][1] ) );
  FADDER S3_362_2 ( .CIN(\ab[362][2] ), .IN0(\CARRYB[361][2] ), .IN1(
        \ab[361][3] ), .COUT(\CARRYB[362][2] ), .SUM(\SUMB[362][2] ) );
  FADDER S1_361_0 ( .CIN(\ab[361][0] ), .IN0(\CARRYB[360][0] ), .IN1(
        \SUMB[360][1] ), .COUT(\CARRYB[361][0] ), .SUM(PRODUCT[361]) );
  FADDER S2_361_1 ( .CIN(\ab[361][1] ), .IN0(\CARRYB[360][1] ), .IN1(
        \SUMB[360][2] ), .COUT(\CARRYB[361][1] ), .SUM(\SUMB[361][1] ) );
  FADDER S3_361_2 ( .CIN(\ab[361][2] ), .IN0(\CARRYB[360][2] ), .IN1(
        \ab[360][3] ), .COUT(\CARRYB[361][2] ), .SUM(\SUMB[361][2] ) );
  FADDER S1_360_0 ( .CIN(\ab[360][0] ), .IN0(\CARRYB[359][0] ), .IN1(
        \SUMB[359][1] ), .COUT(\CARRYB[360][0] ), .SUM(PRODUCT[360]) );
  FADDER S2_360_1 ( .CIN(\ab[360][1] ), .IN0(\CARRYB[359][1] ), .IN1(
        \SUMB[359][2] ), .COUT(\CARRYB[360][1] ), .SUM(\SUMB[360][1] ) );
  FADDER S3_360_2 ( .CIN(\ab[360][2] ), .IN0(\CARRYB[359][2] ), .IN1(
        \ab[359][3] ), .COUT(\CARRYB[360][2] ), .SUM(\SUMB[360][2] ) );
  FADDER S1_359_0 ( .CIN(\ab[359][0] ), .IN0(\CARRYB[358][0] ), .IN1(
        \SUMB[358][1] ), .COUT(\CARRYB[359][0] ), .SUM(PRODUCT[359]) );
  FADDER S2_359_1 ( .CIN(\ab[359][1] ), .IN0(\CARRYB[358][1] ), .IN1(
        \SUMB[358][2] ), .COUT(\CARRYB[359][1] ), .SUM(\SUMB[359][1] ) );
  FADDER S3_359_2 ( .CIN(\ab[359][2] ), .IN0(\CARRYB[358][2] ), .IN1(
        \ab[358][3] ), .COUT(\CARRYB[359][2] ), .SUM(\SUMB[359][2] ) );
  FADDER S1_358_0 ( .CIN(\ab[358][0] ), .IN0(\CARRYB[357][0] ), .IN1(
        \SUMB[357][1] ), .COUT(\CARRYB[358][0] ), .SUM(PRODUCT[358]) );
  FADDER S2_358_1 ( .CIN(\ab[358][1] ), .IN0(\CARRYB[357][1] ), .IN1(
        \SUMB[357][2] ), .COUT(\CARRYB[358][1] ), .SUM(\SUMB[358][1] ) );
  FADDER S3_358_2 ( .CIN(\ab[358][2] ), .IN0(\CARRYB[357][2] ), .IN1(
        \ab[357][3] ), .COUT(\CARRYB[358][2] ), .SUM(\SUMB[358][2] ) );
  FADDER S1_357_0 ( .CIN(\ab[357][0] ), .IN0(\CARRYB[356][0] ), .IN1(
        \SUMB[356][1] ), .COUT(\CARRYB[357][0] ), .SUM(PRODUCT[357]) );
  FADDER S2_357_1 ( .CIN(\ab[357][1] ), .IN0(\CARRYB[356][1] ), .IN1(
        \SUMB[356][2] ), .COUT(\CARRYB[357][1] ), .SUM(\SUMB[357][1] ) );
  FADDER S3_357_2 ( .CIN(\ab[357][2] ), .IN0(\CARRYB[356][2] ), .IN1(
        \ab[356][3] ), .COUT(\CARRYB[357][2] ), .SUM(\SUMB[357][2] ) );
  FADDER S1_356_0 ( .CIN(\ab[356][0] ), .IN0(\CARRYB[355][0] ), .IN1(
        \SUMB[355][1] ), .COUT(\CARRYB[356][0] ), .SUM(PRODUCT[356]) );
  FADDER S2_356_1 ( .CIN(\ab[356][1] ), .IN0(\CARRYB[355][1] ), .IN1(
        \SUMB[355][2] ), .COUT(\CARRYB[356][1] ), .SUM(\SUMB[356][1] ) );
  FADDER S3_356_2 ( .CIN(\ab[356][2] ), .IN0(\CARRYB[355][2] ), .IN1(
        \ab[355][3] ), .COUT(\CARRYB[356][2] ), .SUM(\SUMB[356][2] ) );
  FADDER S1_355_0 ( .CIN(\ab[355][0] ), .IN0(\CARRYB[354][0] ), .IN1(
        \SUMB[354][1] ), .COUT(\CARRYB[355][0] ), .SUM(PRODUCT[355]) );
  FADDER S2_355_1 ( .CIN(\ab[355][1] ), .IN0(\CARRYB[354][1] ), .IN1(
        \SUMB[354][2] ), .COUT(\CARRYB[355][1] ), .SUM(\SUMB[355][1] ) );
  FADDER S3_355_2 ( .CIN(\ab[355][2] ), .IN0(\CARRYB[354][2] ), .IN1(
        \ab[354][3] ), .COUT(\CARRYB[355][2] ), .SUM(\SUMB[355][2] ) );
  FADDER S1_354_0 ( .CIN(\ab[354][0] ), .IN0(\CARRYB[353][0] ), .IN1(
        \SUMB[353][1] ), .COUT(\CARRYB[354][0] ), .SUM(PRODUCT[354]) );
  FADDER S2_354_1 ( .CIN(\ab[354][1] ), .IN0(\CARRYB[353][1] ), .IN1(
        \SUMB[353][2] ), .COUT(\CARRYB[354][1] ), .SUM(\SUMB[354][1] ) );
  FADDER S3_354_2 ( .CIN(\ab[354][2] ), .IN0(\CARRYB[353][2] ), .IN1(
        \ab[353][3] ), .COUT(\CARRYB[354][2] ), .SUM(\SUMB[354][2] ) );
  FADDER S1_353_0 ( .CIN(\ab[353][0] ), .IN0(\CARRYB[352][0] ), .IN1(
        \SUMB[352][1] ), .COUT(\CARRYB[353][0] ), .SUM(PRODUCT[353]) );
  FADDER S2_353_1 ( .CIN(\ab[353][1] ), .IN0(\CARRYB[352][1] ), .IN1(
        \SUMB[352][2] ), .COUT(\CARRYB[353][1] ), .SUM(\SUMB[353][1] ) );
  FADDER S3_353_2 ( .CIN(\ab[353][2] ), .IN0(\CARRYB[352][2] ), .IN1(
        \ab[352][3] ), .COUT(\CARRYB[353][2] ), .SUM(\SUMB[353][2] ) );
  FADDER S1_352_0 ( .CIN(\ab[352][0] ), .IN0(\CARRYB[351][0] ), .IN1(
        \SUMB[351][1] ), .COUT(\CARRYB[352][0] ), .SUM(PRODUCT[352]) );
  FADDER S2_352_1 ( .CIN(\ab[352][1] ), .IN0(\CARRYB[351][1] ), .IN1(
        \SUMB[351][2] ), .COUT(\CARRYB[352][1] ), .SUM(\SUMB[352][1] ) );
  FADDER S3_352_2 ( .CIN(\ab[352][2] ), .IN0(\CARRYB[351][2] ), .IN1(
        \ab[351][3] ), .COUT(\CARRYB[352][2] ), .SUM(\SUMB[352][2] ) );
  FADDER S1_351_0 ( .CIN(\ab[351][0] ), .IN0(\CARRYB[350][0] ), .IN1(
        \SUMB[350][1] ), .COUT(\CARRYB[351][0] ), .SUM(PRODUCT[351]) );
  FADDER S2_351_1 ( .CIN(\ab[351][1] ), .IN0(\CARRYB[350][1] ), .IN1(
        \SUMB[350][2] ), .COUT(\CARRYB[351][1] ), .SUM(\SUMB[351][1] ) );
  FADDER S3_351_2 ( .CIN(\ab[351][2] ), .IN0(\CARRYB[350][2] ), .IN1(
        \ab[350][3] ), .COUT(\CARRYB[351][2] ), .SUM(\SUMB[351][2] ) );
  FADDER S1_350_0 ( .CIN(\ab[350][0] ), .IN0(\CARRYB[349][0] ), .IN1(
        \SUMB[349][1] ), .COUT(\CARRYB[350][0] ), .SUM(PRODUCT[350]) );
  FADDER S2_350_1 ( .CIN(\ab[350][1] ), .IN0(\CARRYB[349][1] ), .IN1(
        \SUMB[349][2] ), .COUT(\CARRYB[350][1] ), .SUM(\SUMB[350][1] ) );
  FADDER S3_350_2 ( .CIN(\ab[350][2] ), .IN0(\CARRYB[349][2] ), .IN1(
        \ab[349][3] ), .COUT(\CARRYB[350][2] ), .SUM(\SUMB[350][2] ) );
  FADDER S1_349_0 ( .CIN(\ab[349][0] ), .IN0(\CARRYB[348][0] ), .IN1(
        \SUMB[348][1] ), .COUT(\CARRYB[349][0] ), .SUM(PRODUCT[349]) );
  FADDER S2_349_1 ( .CIN(\ab[349][1] ), .IN0(\CARRYB[348][1] ), .IN1(
        \SUMB[348][2] ), .COUT(\CARRYB[349][1] ), .SUM(\SUMB[349][1] ) );
  FADDER S3_349_2 ( .CIN(\ab[349][2] ), .IN0(\CARRYB[348][2] ), .IN1(
        \ab[348][3] ), .COUT(\CARRYB[349][2] ), .SUM(\SUMB[349][2] ) );
  FADDER S1_348_0 ( .CIN(\ab[348][0] ), .IN0(\CARRYB[347][0] ), .IN1(
        \SUMB[347][1] ), .COUT(\CARRYB[348][0] ), .SUM(PRODUCT[348]) );
  FADDER S2_348_1 ( .CIN(\ab[348][1] ), .IN0(\CARRYB[347][1] ), .IN1(
        \SUMB[347][2] ), .COUT(\CARRYB[348][1] ), .SUM(\SUMB[348][1] ) );
  FADDER S3_348_2 ( .CIN(\ab[348][2] ), .IN0(\CARRYB[347][2] ), .IN1(
        \ab[347][3] ), .COUT(\CARRYB[348][2] ), .SUM(\SUMB[348][2] ) );
  FADDER S1_347_0 ( .CIN(\ab[347][0] ), .IN0(\CARRYB[346][0] ), .IN1(
        \SUMB[346][1] ), .COUT(\CARRYB[347][0] ), .SUM(PRODUCT[347]) );
  FADDER S2_347_1 ( .CIN(\ab[347][1] ), .IN0(\CARRYB[346][1] ), .IN1(
        \SUMB[346][2] ), .COUT(\CARRYB[347][1] ), .SUM(\SUMB[347][1] ) );
  FADDER S3_347_2 ( .CIN(\ab[347][2] ), .IN0(\CARRYB[346][2] ), .IN1(
        \ab[346][3] ), .COUT(\CARRYB[347][2] ), .SUM(\SUMB[347][2] ) );
  FADDER S1_346_0 ( .CIN(\ab[346][0] ), .IN0(\CARRYB[345][0] ), .IN1(
        \SUMB[345][1] ), .COUT(\CARRYB[346][0] ), .SUM(PRODUCT[346]) );
  FADDER S2_346_1 ( .CIN(\ab[346][1] ), .IN0(\CARRYB[345][1] ), .IN1(
        \SUMB[345][2] ), .COUT(\CARRYB[346][1] ), .SUM(\SUMB[346][1] ) );
  FADDER S3_346_2 ( .CIN(\ab[346][2] ), .IN0(\CARRYB[345][2] ), .IN1(
        \ab[345][3] ), .COUT(\CARRYB[346][2] ), .SUM(\SUMB[346][2] ) );
  FADDER S1_345_0 ( .CIN(\ab[345][0] ), .IN0(\CARRYB[344][0] ), .IN1(
        \SUMB[344][1] ), .COUT(\CARRYB[345][0] ), .SUM(PRODUCT[345]) );
  FADDER S2_345_1 ( .CIN(\ab[345][1] ), .IN0(\CARRYB[344][1] ), .IN1(
        \SUMB[344][2] ), .COUT(\CARRYB[345][1] ), .SUM(\SUMB[345][1] ) );
  FADDER S3_345_2 ( .CIN(\ab[345][2] ), .IN0(\CARRYB[344][2] ), .IN1(
        \ab[344][3] ), .COUT(\CARRYB[345][2] ), .SUM(\SUMB[345][2] ) );
  FADDER S1_344_0 ( .CIN(\ab[344][0] ), .IN0(\CARRYB[343][0] ), .IN1(
        \SUMB[343][1] ), .COUT(\CARRYB[344][0] ), .SUM(PRODUCT[344]) );
  FADDER S2_344_1 ( .CIN(\ab[344][1] ), .IN0(\CARRYB[343][1] ), .IN1(
        \SUMB[343][2] ), .COUT(\CARRYB[344][1] ), .SUM(\SUMB[344][1] ) );
  FADDER S3_344_2 ( .CIN(\ab[344][2] ), .IN0(\CARRYB[343][2] ), .IN1(
        \ab[343][3] ), .COUT(\CARRYB[344][2] ), .SUM(\SUMB[344][2] ) );
  FADDER S1_343_0 ( .CIN(\ab[343][0] ), .IN0(\CARRYB[342][0] ), .IN1(
        \SUMB[342][1] ), .COUT(\CARRYB[343][0] ), .SUM(PRODUCT[343]) );
  FADDER S2_343_1 ( .CIN(\ab[343][1] ), .IN0(\CARRYB[342][1] ), .IN1(
        \SUMB[342][2] ), .COUT(\CARRYB[343][1] ), .SUM(\SUMB[343][1] ) );
  FADDER S3_343_2 ( .CIN(\ab[343][2] ), .IN0(\CARRYB[342][2] ), .IN1(
        \ab[342][3] ), .COUT(\CARRYB[343][2] ), .SUM(\SUMB[343][2] ) );
  FADDER S1_342_0 ( .CIN(\ab[342][0] ), .IN0(\CARRYB[341][0] ), .IN1(
        \SUMB[341][1] ), .COUT(\CARRYB[342][0] ), .SUM(PRODUCT[342]) );
  FADDER S2_342_1 ( .CIN(\ab[342][1] ), .IN0(\CARRYB[341][1] ), .IN1(
        \SUMB[341][2] ), .COUT(\CARRYB[342][1] ), .SUM(\SUMB[342][1] ) );
  FADDER S3_342_2 ( .CIN(\ab[342][2] ), .IN0(\CARRYB[341][2] ), .IN1(
        \ab[341][3] ), .COUT(\CARRYB[342][2] ), .SUM(\SUMB[342][2] ) );
  FADDER S1_341_0 ( .CIN(\ab[341][0] ), .IN0(\CARRYB[340][0] ), .IN1(
        \SUMB[340][1] ), .COUT(\CARRYB[341][0] ), .SUM(PRODUCT[341]) );
  FADDER S2_341_1 ( .CIN(\ab[341][1] ), .IN0(\CARRYB[340][1] ), .IN1(
        \SUMB[340][2] ), .COUT(\CARRYB[341][1] ), .SUM(\SUMB[341][1] ) );
  FADDER S3_341_2 ( .CIN(\ab[341][2] ), .IN0(\CARRYB[340][2] ), .IN1(
        \ab[340][3] ), .COUT(\CARRYB[341][2] ), .SUM(\SUMB[341][2] ) );
  FADDER S1_340_0 ( .CIN(\ab[340][0] ), .IN0(\CARRYB[339][0] ), .IN1(
        \SUMB[339][1] ), .COUT(\CARRYB[340][0] ), .SUM(PRODUCT[340]) );
  FADDER S2_340_1 ( .CIN(\ab[340][1] ), .IN0(\CARRYB[339][1] ), .IN1(
        \SUMB[339][2] ), .COUT(\CARRYB[340][1] ), .SUM(\SUMB[340][1] ) );
  FADDER S3_340_2 ( .CIN(\ab[340][2] ), .IN0(\CARRYB[339][2] ), .IN1(
        \ab[339][3] ), .COUT(\CARRYB[340][2] ), .SUM(\SUMB[340][2] ) );
  FADDER S1_339_0 ( .CIN(\ab[339][0] ), .IN0(\CARRYB[338][0] ), .IN1(
        \SUMB[338][1] ), .COUT(\CARRYB[339][0] ), .SUM(PRODUCT[339]) );
  FADDER S2_339_1 ( .CIN(\ab[339][1] ), .IN0(\CARRYB[338][1] ), .IN1(
        \SUMB[338][2] ), .COUT(\CARRYB[339][1] ), .SUM(\SUMB[339][1] ) );
  FADDER S3_339_2 ( .CIN(\ab[339][2] ), .IN0(\CARRYB[338][2] ), .IN1(
        \ab[338][3] ), .COUT(\CARRYB[339][2] ), .SUM(\SUMB[339][2] ) );
  FADDER S1_338_0 ( .CIN(\ab[338][0] ), .IN0(\CARRYB[337][0] ), .IN1(
        \SUMB[337][1] ), .COUT(\CARRYB[338][0] ), .SUM(PRODUCT[338]) );
  FADDER S2_338_1 ( .CIN(\ab[338][1] ), .IN0(\CARRYB[337][1] ), .IN1(
        \SUMB[337][2] ), .COUT(\CARRYB[338][1] ), .SUM(\SUMB[338][1] ) );
  FADDER S3_338_2 ( .CIN(\ab[338][2] ), .IN0(\CARRYB[337][2] ), .IN1(
        \ab[337][3] ), .COUT(\CARRYB[338][2] ), .SUM(\SUMB[338][2] ) );
  FADDER S1_337_0 ( .CIN(\ab[337][0] ), .IN0(\CARRYB[336][0] ), .IN1(
        \SUMB[336][1] ), .COUT(\CARRYB[337][0] ), .SUM(PRODUCT[337]) );
  FADDER S2_337_1 ( .CIN(\ab[337][1] ), .IN0(\CARRYB[336][1] ), .IN1(
        \SUMB[336][2] ), .COUT(\CARRYB[337][1] ), .SUM(\SUMB[337][1] ) );
  FADDER S3_337_2 ( .CIN(\ab[337][2] ), .IN0(\CARRYB[336][2] ), .IN1(
        \ab[336][3] ), .COUT(\CARRYB[337][2] ), .SUM(\SUMB[337][2] ) );
  FADDER S1_336_0 ( .CIN(\ab[336][0] ), .IN0(\CARRYB[335][0] ), .IN1(
        \SUMB[335][1] ), .COUT(\CARRYB[336][0] ), .SUM(PRODUCT[336]) );
  FADDER S2_336_1 ( .CIN(\ab[336][1] ), .IN0(\CARRYB[335][1] ), .IN1(
        \SUMB[335][2] ), .COUT(\CARRYB[336][1] ), .SUM(\SUMB[336][1] ) );
  FADDER S3_336_2 ( .CIN(\ab[336][2] ), .IN0(\CARRYB[335][2] ), .IN1(
        \ab[335][3] ), .COUT(\CARRYB[336][2] ), .SUM(\SUMB[336][2] ) );
  FADDER S1_335_0 ( .CIN(\ab[335][0] ), .IN0(\CARRYB[334][0] ), .IN1(
        \SUMB[334][1] ), .COUT(\CARRYB[335][0] ), .SUM(PRODUCT[335]) );
  FADDER S2_335_1 ( .CIN(\ab[335][1] ), .IN0(\CARRYB[334][1] ), .IN1(
        \SUMB[334][2] ), .COUT(\CARRYB[335][1] ), .SUM(\SUMB[335][1] ) );
  FADDER S3_335_2 ( .CIN(\ab[335][2] ), .IN0(\CARRYB[334][2] ), .IN1(
        \ab[334][3] ), .COUT(\CARRYB[335][2] ), .SUM(\SUMB[335][2] ) );
  FADDER S1_334_0 ( .CIN(\ab[334][0] ), .IN0(\CARRYB[333][0] ), .IN1(
        \SUMB[333][1] ), .COUT(\CARRYB[334][0] ), .SUM(PRODUCT[334]) );
  FADDER S2_334_1 ( .CIN(\ab[334][1] ), .IN0(\CARRYB[333][1] ), .IN1(
        \SUMB[333][2] ), .COUT(\CARRYB[334][1] ), .SUM(\SUMB[334][1] ) );
  FADDER S3_334_2 ( .CIN(\ab[334][2] ), .IN0(\CARRYB[333][2] ), .IN1(
        \ab[333][3] ), .COUT(\CARRYB[334][2] ), .SUM(\SUMB[334][2] ) );
  FADDER S1_333_0 ( .CIN(\ab[333][0] ), .IN0(\CARRYB[332][0] ), .IN1(
        \SUMB[332][1] ), .COUT(\CARRYB[333][0] ), .SUM(PRODUCT[333]) );
  FADDER S2_333_1 ( .CIN(\ab[333][1] ), .IN0(\CARRYB[332][1] ), .IN1(
        \SUMB[332][2] ), .COUT(\CARRYB[333][1] ), .SUM(\SUMB[333][1] ) );
  FADDER S3_333_2 ( .CIN(\ab[333][2] ), .IN0(\CARRYB[332][2] ), .IN1(
        \ab[332][3] ), .COUT(\CARRYB[333][2] ), .SUM(\SUMB[333][2] ) );
  FADDER S1_332_0 ( .CIN(\ab[332][0] ), .IN0(\CARRYB[331][0] ), .IN1(
        \SUMB[331][1] ), .COUT(\CARRYB[332][0] ), .SUM(PRODUCT[332]) );
  FADDER S2_332_1 ( .CIN(\ab[332][1] ), .IN0(\CARRYB[331][1] ), .IN1(
        \SUMB[331][2] ), .COUT(\CARRYB[332][1] ), .SUM(\SUMB[332][1] ) );
  FADDER S3_332_2 ( .CIN(\ab[332][2] ), .IN0(\CARRYB[331][2] ), .IN1(
        \ab[331][3] ), .COUT(\CARRYB[332][2] ), .SUM(\SUMB[332][2] ) );
  FADDER S1_331_0 ( .CIN(\ab[331][0] ), .IN0(\CARRYB[330][0] ), .IN1(
        \SUMB[330][1] ), .COUT(\CARRYB[331][0] ), .SUM(PRODUCT[331]) );
  FADDER S2_331_1 ( .CIN(\ab[331][1] ), .IN0(\CARRYB[330][1] ), .IN1(
        \SUMB[330][2] ), .COUT(\CARRYB[331][1] ), .SUM(\SUMB[331][1] ) );
  FADDER S3_331_2 ( .CIN(\ab[331][2] ), .IN0(\CARRYB[330][2] ), .IN1(
        \ab[330][3] ), .COUT(\CARRYB[331][2] ), .SUM(\SUMB[331][2] ) );
  FADDER S1_330_0 ( .CIN(\ab[330][0] ), .IN0(\CARRYB[329][0] ), .IN1(
        \SUMB[329][1] ), .COUT(\CARRYB[330][0] ), .SUM(PRODUCT[330]) );
  FADDER S2_330_1 ( .CIN(\ab[330][1] ), .IN0(\CARRYB[329][1] ), .IN1(
        \SUMB[329][2] ), .COUT(\CARRYB[330][1] ), .SUM(\SUMB[330][1] ) );
  FADDER S3_330_2 ( .CIN(\ab[330][2] ), .IN0(\CARRYB[329][2] ), .IN1(
        \ab[329][3] ), .COUT(\CARRYB[330][2] ), .SUM(\SUMB[330][2] ) );
  FADDER S1_329_0 ( .CIN(\ab[329][0] ), .IN0(\CARRYB[328][0] ), .IN1(
        \SUMB[328][1] ), .COUT(\CARRYB[329][0] ), .SUM(PRODUCT[329]) );
  FADDER S2_329_1 ( .CIN(\ab[329][1] ), .IN0(\CARRYB[328][1] ), .IN1(
        \SUMB[328][2] ), .COUT(\CARRYB[329][1] ), .SUM(\SUMB[329][1] ) );
  FADDER S3_329_2 ( .CIN(\ab[329][2] ), .IN0(\CARRYB[328][2] ), .IN1(
        \ab[328][3] ), .COUT(\CARRYB[329][2] ), .SUM(\SUMB[329][2] ) );
  FADDER S1_328_0 ( .CIN(\ab[328][0] ), .IN0(\CARRYB[327][0] ), .IN1(
        \SUMB[327][1] ), .COUT(\CARRYB[328][0] ), .SUM(PRODUCT[328]) );
  FADDER S2_328_1 ( .CIN(\ab[328][1] ), .IN0(\CARRYB[327][1] ), .IN1(
        \SUMB[327][2] ), .COUT(\CARRYB[328][1] ), .SUM(\SUMB[328][1] ) );
  FADDER S3_328_2 ( .CIN(\ab[328][2] ), .IN0(\CARRYB[327][2] ), .IN1(
        \ab[327][3] ), .COUT(\CARRYB[328][2] ), .SUM(\SUMB[328][2] ) );
  FADDER S1_327_0 ( .CIN(\ab[327][0] ), .IN0(\CARRYB[326][0] ), .IN1(
        \SUMB[326][1] ), .COUT(\CARRYB[327][0] ), .SUM(PRODUCT[327]) );
  FADDER S2_327_1 ( .CIN(\ab[327][1] ), .IN0(\CARRYB[326][1] ), .IN1(
        \SUMB[326][2] ), .COUT(\CARRYB[327][1] ), .SUM(\SUMB[327][1] ) );
  FADDER S3_327_2 ( .CIN(\ab[327][2] ), .IN0(\CARRYB[326][2] ), .IN1(
        \ab[326][3] ), .COUT(\CARRYB[327][2] ), .SUM(\SUMB[327][2] ) );
  FADDER S1_326_0 ( .CIN(\ab[326][0] ), .IN0(\CARRYB[325][0] ), .IN1(
        \SUMB[325][1] ), .COUT(\CARRYB[326][0] ), .SUM(PRODUCT[326]) );
  FADDER S2_326_1 ( .CIN(\ab[326][1] ), .IN0(\CARRYB[325][1] ), .IN1(
        \SUMB[325][2] ), .COUT(\CARRYB[326][1] ), .SUM(\SUMB[326][1] ) );
  FADDER S3_326_2 ( .CIN(\ab[326][2] ), .IN0(\CARRYB[325][2] ), .IN1(
        \ab[325][3] ), .COUT(\CARRYB[326][2] ), .SUM(\SUMB[326][2] ) );
  FADDER S1_325_0 ( .CIN(\ab[325][0] ), .IN0(\CARRYB[324][0] ), .IN1(
        \SUMB[324][1] ), .COUT(\CARRYB[325][0] ), .SUM(PRODUCT[325]) );
  FADDER S2_325_1 ( .CIN(\ab[325][1] ), .IN0(\CARRYB[324][1] ), .IN1(
        \SUMB[324][2] ), .COUT(\CARRYB[325][1] ), .SUM(\SUMB[325][1] ) );
  FADDER S3_325_2 ( .CIN(\ab[325][2] ), .IN0(\CARRYB[324][2] ), .IN1(
        \ab[324][3] ), .COUT(\CARRYB[325][2] ), .SUM(\SUMB[325][2] ) );
  FADDER S1_324_0 ( .CIN(\ab[324][0] ), .IN0(\CARRYB[323][0] ), .IN1(
        \SUMB[323][1] ), .COUT(\CARRYB[324][0] ), .SUM(PRODUCT[324]) );
  FADDER S2_324_1 ( .CIN(\ab[324][1] ), .IN0(\CARRYB[323][1] ), .IN1(
        \SUMB[323][2] ), .COUT(\CARRYB[324][1] ), .SUM(\SUMB[324][1] ) );
  FADDER S3_324_2 ( .CIN(\ab[324][2] ), .IN0(\CARRYB[323][2] ), .IN1(
        \ab[323][3] ), .COUT(\CARRYB[324][2] ), .SUM(\SUMB[324][2] ) );
  FADDER S1_323_0 ( .CIN(\ab[323][0] ), .IN0(\CARRYB[322][0] ), .IN1(
        \SUMB[322][1] ), .COUT(\CARRYB[323][0] ), .SUM(PRODUCT[323]) );
  FADDER S2_323_1 ( .CIN(\ab[323][1] ), .IN0(\CARRYB[322][1] ), .IN1(
        \SUMB[322][2] ), .COUT(\CARRYB[323][1] ), .SUM(\SUMB[323][1] ) );
  FADDER S3_323_2 ( .CIN(\ab[323][2] ), .IN0(\CARRYB[322][2] ), .IN1(
        \ab[322][3] ), .COUT(\CARRYB[323][2] ), .SUM(\SUMB[323][2] ) );
  FADDER S1_322_0 ( .CIN(\ab[322][0] ), .IN0(\CARRYB[321][0] ), .IN1(
        \SUMB[321][1] ), .COUT(\CARRYB[322][0] ), .SUM(PRODUCT[322]) );
  FADDER S2_322_1 ( .CIN(\ab[322][1] ), .IN0(\CARRYB[321][1] ), .IN1(
        \SUMB[321][2] ), .COUT(\CARRYB[322][1] ), .SUM(\SUMB[322][1] ) );
  FADDER S3_322_2 ( .CIN(\ab[322][2] ), .IN0(\CARRYB[321][2] ), .IN1(
        \ab[321][3] ), .COUT(\CARRYB[322][2] ), .SUM(\SUMB[322][2] ) );
  FADDER S1_321_0 ( .CIN(\ab[321][0] ), .IN0(\CARRYB[320][0] ), .IN1(
        \SUMB[320][1] ), .COUT(\CARRYB[321][0] ), .SUM(PRODUCT[321]) );
  FADDER S2_321_1 ( .CIN(\ab[321][1] ), .IN0(\CARRYB[320][1] ), .IN1(
        \SUMB[320][2] ), .COUT(\CARRYB[321][1] ), .SUM(\SUMB[321][1] ) );
  FADDER S3_321_2 ( .CIN(\ab[321][2] ), .IN0(\CARRYB[320][2] ), .IN1(
        \ab[320][3] ), .COUT(\CARRYB[321][2] ), .SUM(\SUMB[321][2] ) );
  FADDER S1_320_0 ( .CIN(\ab[320][0] ), .IN0(\CARRYB[319][0] ), .IN1(
        \SUMB[319][1] ), .COUT(\CARRYB[320][0] ), .SUM(PRODUCT[320]) );
  FADDER S2_320_1 ( .CIN(\ab[320][1] ), .IN0(\CARRYB[319][1] ), .IN1(
        \SUMB[319][2] ), .COUT(\CARRYB[320][1] ), .SUM(\SUMB[320][1] ) );
  FADDER S3_320_2 ( .CIN(\ab[320][2] ), .IN0(\CARRYB[319][2] ), .IN1(
        \ab[319][3] ), .COUT(\CARRYB[320][2] ), .SUM(\SUMB[320][2] ) );
  FADDER S1_319_0 ( .CIN(\ab[319][0] ), .IN0(\CARRYB[318][0] ), .IN1(
        \SUMB[318][1] ), .COUT(\CARRYB[319][0] ), .SUM(PRODUCT[319]) );
  FADDER S2_319_1 ( .CIN(\ab[319][1] ), .IN0(\CARRYB[318][1] ), .IN1(
        \SUMB[318][2] ), .COUT(\CARRYB[319][1] ), .SUM(\SUMB[319][1] ) );
  FADDER S3_319_2 ( .CIN(\ab[319][2] ), .IN0(\CARRYB[318][2] ), .IN1(
        \ab[318][3] ), .COUT(\CARRYB[319][2] ), .SUM(\SUMB[319][2] ) );
  FADDER S1_318_0 ( .CIN(\ab[318][0] ), .IN0(\CARRYB[317][0] ), .IN1(
        \SUMB[317][1] ), .COUT(\CARRYB[318][0] ), .SUM(PRODUCT[318]) );
  FADDER S2_318_1 ( .CIN(\ab[318][1] ), .IN0(\CARRYB[317][1] ), .IN1(
        \SUMB[317][2] ), .COUT(\CARRYB[318][1] ), .SUM(\SUMB[318][1] ) );
  FADDER S3_318_2 ( .CIN(\ab[318][2] ), .IN0(\CARRYB[317][2] ), .IN1(
        \ab[317][3] ), .COUT(\CARRYB[318][2] ), .SUM(\SUMB[318][2] ) );
  FADDER S1_317_0 ( .CIN(\ab[317][0] ), .IN0(\CARRYB[316][0] ), .IN1(
        \SUMB[316][1] ), .COUT(\CARRYB[317][0] ), .SUM(PRODUCT[317]) );
  FADDER S2_317_1 ( .CIN(\ab[317][1] ), .IN0(\CARRYB[316][1] ), .IN1(
        \SUMB[316][2] ), .COUT(\CARRYB[317][1] ), .SUM(\SUMB[317][1] ) );
  FADDER S3_317_2 ( .CIN(\ab[317][2] ), .IN0(\CARRYB[316][2] ), .IN1(
        \ab[316][3] ), .COUT(\CARRYB[317][2] ), .SUM(\SUMB[317][2] ) );
  FADDER S1_316_0 ( .CIN(\ab[316][0] ), .IN0(\CARRYB[315][0] ), .IN1(
        \SUMB[315][1] ), .COUT(\CARRYB[316][0] ), .SUM(PRODUCT[316]) );
  FADDER S2_316_1 ( .CIN(\ab[316][1] ), .IN0(\CARRYB[315][1] ), .IN1(
        \SUMB[315][2] ), .COUT(\CARRYB[316][1] ), .SUM(\SUMB[316][1] ) );
  FADDER S3_316_2 ( .CIN(\ab[316][2] ), .IN0(\CARRYB[315][2] ), .IN1(
        \ab[315][3] ), .COUT(\CARRYB[316][2] ), .SUM(\SUMB[316][2] ) );
  FADDER S1_315_0 ( .CIN(\ab[315][0] ), .IN0(\CARRYB[314][0] ), .IN1(
        \SUMB[314][1] ), .COUT(\CARRYB[315][0] ), .SUM(PRODUCT[315]) );
  FADDER S2_315_1 ( .CIN(\ab[315][1] ), .IN0(\CARRYB[314][1] ), .IN1(
        \SUMB[314][2] ), .COUT(\CARRYB[315][1] ), .SUM(\SUMB[315][1] ) );
  FADDER S3_315_2 ( .CIN(\ab[315][2] ), .IN0(\CARRYB[314][2] ), .IN1(
        \ab[314][3] ), .COUT(\CARRYB[315][2] ), .SUM(\SUMB[315][2] ) );
  FADDER S1_314_0 ( .CIN(\ab[314][0] ), .IN0(\CARRYB[313][0] ), .IN1(
        \SUMB[313][1] ), .COUT(\CARRYB[314][0] ), .SUM(PRODUCT[314]) );
  FADDER S2_314_1 ( .CIN(\ab[314][1] ), .IN0(\CARRYB[313][1] ), .IN1(
        \SUMB[313][2] ), .COUT(\CARRYB[314][1] ), .SUM(\SUMB[314][1] ) );
  FADDER S3_314_2 ( .CIN(\ab[314][2] ), .IN0(\CARRYB[313][2] ), .IN1(
        \ab[313][3] ), .COUT(\CARRYB[314][2] ), .SUM(\SUMB[314][2] ) );
  FADDER S1_313_0 ( .CIN(\ab[313][0] ), .IN0(\CARRYB[312][0] ), .IN1(
        \SUMB[312][1] ), .COUT(\CARRYB[313][0] ), .SUM(PRODUCT[313]) );
  FADDER S2_313_1 ( .CIN(\ab[313][1] ), .IN0(\CARRYB[312][1] ), .IN1(
        \SUMB[312][2] ), .COUT(\CARRYB[313][1] ), .SUM(\SUMB[313][1] ) );
  FADDER S3_313_2 ( .CIN(\ab[313][2] ), .IN0(\CARRYB[312][2] ), .IN1(
        \ab[312][3] ), .COUT(\CARRYB[313][2] ), .SUM(\SUMB[313][2] ) );
  FADDER S1_312_0 ( .CIN(\ab[312][0] ), .IN0(\CARRYB[311][0] ), .IN1(
        \SUMB[311][1] ), .COUT(\CARRYB[312][0] ), .SUM(PRODUCT[312]) );
  FADDER S2_312_1 ( .CIN(\ab[312][1] ), .IN0(\CARRYB[311][1] ), .IN1(
        \SUMB[311][2] ), .COUT(\CARRYB[312][1] ), .SUM(\SUMB[312][1] ) );
  FADDER S3_312_2 ( .CIN(\ab[312][2] ), .IN0(\CARRYB[311][2] ), .IN1(
        \ab[311][3] ), .COUT(\CARRYB[312][2] ), .SUM(\SUMB[312][2] ) );
  FADDER S1_311_0 ( .CIN(\ab[311][0] ), .IN0(\CARRYB[310][0] ), .IN1(
        \SUMB[310][1] ), .COUT(\CARRYB[311][0] ), .SUM(PRODUCT[311]) );
  FADDER S2_311_1 ( .CIN(\ab[311][1] ), .IN0(\CARRYB[310][1] ), .IN1(
        \SUMB[310][2] ), .COUT(\CARRYB[311][1] ), .SUM(\SUMB[311][1] ) );
  FADDER S3_311_2 ( .CIN(\ab[311][2] ), .IN0(\CARRYB[310][2] ), .IN1(
        \ab[310][3] ), .COUT(\CARRYB[311][2] ), .SUM(\SUMB[311][2] ) );
  FADDER S1_310_0 ( .CIN(\ab[310][0] ), .IN0(\CARRYB[309][0] ), .IN1(
        \SUMB[309][1] ), .COUT(\CARRYB[310][0] ), .SUM(PRODUCT[310]) );
  FADDER S2_310_1 ( .CIN(\ab[310][1] ), .IN0(\CARRYB[309][1] ), .IN1(
        \SUMB[309][2] ), .COUT(\CARRYB[310][1] ), .SUM(\SUMB[310][1] ) );
  FADDER S3_310_2 ( .CIN(\ab[310][2] ), .IN0(\CARRYB[309][2] ), .IN1(
        \ab[309][3] ), .COUT(\CARRYB[310][2] ), .SUM(\SUMB[310][2] ) );
  FADDER S1_309_0 ( .CIN(\ab[309][0] ), .IN0(\CARRYB[308][0] ), .IN1(
        \SUMB[308][1] ), .COUT(\CARRYB[309][0] ), .SUM(PRODUCT[309]) );
  FADDER S2_309_1 ( .CIN(\ab[309][1] ), .IN0(\CARRYB[308][1] ), .IN1(
        \SUMB[308][2] ), .COUT(\CARRYB[309][1] ), .SUM(\SUMB[309][1] ) );
  FADDER S3_309_2 ( .CIN(\ab[309][2] ), .IN0(\CARRYB[308][2] ), .IN1(
        \ab[308][3] ), .COUT(\CARRYB[309][2] ), .SUM(\SUMB[309][2] ) );
  FADDER S1_308_0 ( .CIN(\ab[308][0] ), .IN0(\CARRYB[307][0] ), .IN1(
        \SUMB[307][1] ), .COUT(\CARRYB[308][0] ), .SUM(PRODUCT[308]) );
  FADDER S2_308_1 ( .CIN(\ab[308][1] ), .IN0(\CARRYB[307][1] ), .IN1(
        \SUMB[307][2] ), .COUT(\CARRYB[308][1] ), .SUM(\SUMB[308][1] ) );
  FADDER S3_308_2 ( .CIN(\ab[308][2] ), .IN0(\CARRYB[307][2] ), .IN1(
        \ab[307][3] ), .COUT(\CARRYB[308][2] ), .SUM(\SUMB[308][2] ) );
  FADDER S1_307_0 ( .CIN(\ab[307][0] ), .IN0(\CARRYB[306][0] ), .IN1(
        \SUMB[306][1] ), .COUT(\CARRYB[307][0] ), .SUM(PRODUCT[307]) );
  FADDER S2_307_1 ( .CIN(\ab[307][1] ), .IN0(\CARRYB[306][1] ), .IN1(
        \SUMB[306][2] ), .COUT(\CARRYB[307][1] ), .SUM(\SUMB[307][1] ) );
  FADDER S3_307_2 ( .CIN(\ab[307][2] ), .IN0(\CARRYB[306][2] ), .IN1(
        \ab[306][3] ), .COUT(\CARRYB[307][2] ), .SUM(\SUMB[307][2] ) );
  FADDER S1_306_0 ( .CIN(\ab[306][0] ), .IN0(\CARRYB[305][0] ), .IN1(
        \SUMB[305][1] ), .COUT(\CARRYB[306][0] ), .SUM(PRODUCT[306]) );
  FADDER S2_306_1 ( .CIN(\ab[306][1] ), .IN0(\CARRYB[305][1] ), .IN1(
        \SUMB[305][2] ), .COUT(\CARRYB[306][1] ), .SUM(\SUMB[306][1] ) );
  FADDER S3_306_2 ( .CIN(\ab[306][2] ), .IN0(\CARRYB[305][2] ), .IN1(
        \ab[305][3] ), .COUT(\CARRYB[306][2] ), .SUM(\SUMB[306][2] ) );
  FADDER S1_305_0 ( .CIN(\ab[305][0] ), .IN0(\CARRYB[304][0] ), .IN1(
        \SUMB[304][1] ), .COUT(\CARRYB[305][0] ), .SUM(PRODUCT[305]) );
  FADDER S2_305_1 ( .CIN(\ab[305][1] ), .IN0(\CARRYB[304][1] ), .IN1(
        \SUMB[304][2] ), .COUT(\CARRYB[305][1] ), .SUM(\SUMB[305][1] ) );
  FADDER S3_305_2 ( .CIN(\ab[305][2] ), .IN0(\CARRYB[304][2] ), .IN1(
        \ab[304][3] ), .COUT(\CARRYB[305][2] ), .SUM(\SUMB[305][2] ) );
  FADDER S1_304_0 ( .CIN(\ab[304][0] ), .IN0(\CARRYB[303][0] ), .IN1(
        \SUMB[303][1] ), .COUT(\CARRYB[304][0] ), .SUM(PRODUCT[304]) );
  FADDER S2_304_1 ( .CIN(\ab[304][1] ), .IN0(\CARRYB[303][1] ), .IN1(
        \SUMB[303][2] ), .COUT(\CARRYB[304][1] ), .SUM(\SUMB[304][1] ) );
  FADDER S3_304_2 ( .CIN(\ab[304][2] ), .IN0(\CARRYB[303][2] ), .IN1(
        \ab[303][3] ), .COUT(\CARRYB[304][2] ), .SUM(\SUMB[304][2] ) );
  FADDER S1_303_0 ( .CIN(\ab[303][0] ), .IN0(\CARRYB[302][0] ), .IN1(
        \SUMB[302][1] ), .COUT(\CARRYB[303][0] ), .SUM(PRODUCT[303]) );
  FADDER S2_303_1 ( .CIN(\ab[303][1] ), .IN0(\CARRYB[302][1] ), .IN1(
        \SUMB[302][2] ), .COUT(\CARRYB[303][1] ), .SUM(\SUMB[303][1] ) );
  FADDER S3_303_2 ( .CIN(\ab[303][2] ), .IN0(\CARRYB[302][2] ), .IN1(
        \ab[302][3] ), .COUT(\CARRYB[303][2] ), .SUM(\SUMB[303][2] ) );
  FADDER S1_302_0 ( .CIN(\ab[302][0] ), .IN0(\CARRYB[301][0] ), .IN1(
        \SUMB[301][1] ), .COUT(\CARRYB[302][0] ), .SUM(PRODUCT[302]) );
  FADDER S2_302_1 ( .CIN(\ab[302][1] ), .IN0(\CARRYB[301][1] ), .IN1(
        \SUMB[301][2] ), .COUT(\CARRYB[302][1] ), .SUM(\SUMB[302][1] ) );
  FADDER S3_302_2 ( .CIN(\ab[302][2] ), .IN0(\CARRYB[301][2] ), .IN1(
        \ab[301][3] ), .COUT(\CARRYB[302][2] ), .SUM(\SUMB[302][2] ) );
  FADDER S1_301_0 ( .CIN(\ab[301][0] ), .IN0(\CARRYB[300][0] ), .IN1(
        \SUMB[300][1] ), .COUT(\CARRYB[301][0] ), .SUM(PRODUCT[301]) );
  FADDER S2_301_1 ( .CIN(\ab[301][1] ), .IN0(\CARRYB[300][1] ), .IN1(
        \SUMB[300][2] ), .COUT(\CARRYB[301][1] ), .SUM(\SUMB[301][1] ) );
  FADDER S3_301_2 ( .CIN(\ab[301][2] ), .IN0(\CARRYB[300][2] ), .IN1(
        \ab[300][3] ), .COUT(\CARRYB[301][2] ), .SUM(\SUMB[301][2] ) );
  FADDER S1_300_0 ( .CIN(\ab[300][0] ), .IN0(\CARRYB[299][0] ), .IN1(
        \SUMB[299][1] ), .COUT(\CARRYB[300][0] ), .SUM(PRODUCT[300]) );
  FADDER S2_300_1 ( .CIN(\ab[300][1] ), .IN0(\CARRYB[299][1] ), .IN1(
        \SUMB[299][2] ), .COUT(\CARRYB[300][1] ), .SUM(\SUMB[300][1] ) );
  FADDER S3_300_2 ( .CIN(\ab[300][2] ), .IN0(\CARRYB[299][2] ), .IN1(
        \ab[299][3] ), .COUT(\CARRYB[300][2] ), .SUM(\SUMB[300][2] ) );
  FADDER S1_299_0 ( .CIN(\ab[299][0] ), .IN0(\CARRYB[298][0] ), .IN1(
        \SUMB[298][1] ), .COUT(\CARRYB[299][0] ), .SUM(PRODUCT[299]) );
  FADDER S2_299_1 ( .CIN(\ab[299][1] ), .IN0(\CARRYB[298][1] ), .IN1(
        \SUMB[298][2] ), .COUT(\CARRYB[299][1] ), .SUM(\SUMB[299][1] ) );
  FADDER S3_299_2 ( .CIN(\ab[299][2] ), .IN0(\CARRYB[298][2] ), .IN1(
        \ab[298][3] ), .COUT(\CARRYB[299][2] ), .SUM(\SUMB[299][2] ) );
  FADDER S1_298_0 ( .CIN(\ab[298][0] ), .IN0(\CARRYB[297][0] ), .IN1(
        \SUMB[297][1] ), .COUT(\CARRYB[298][0] ), .SUM(PRODUCT[298]) );
  FADDER S2_298_1 ( .CIN(\ab[298][1] ), .IN0(\CARRYB[297][1] ), .IN1(
        \SUMB[297][2] ), .COUT(\CARRYB[298][1] ), .SUM(\SUMB[298][1] ) );
  FADDER S3_298_2 ( .CIN(\ab[298][2] ), .IN0(\CARRYB[297][2] ), .IN1(
        \ab[297][3] ), .COUT(\CARRYB[298][2] ), .SUM(\SUMB[298][2] ) );
  FADDER S1_297_0 ( .CIN(\ab[297][0] ), .IN0(\CARRYB[296][0] ), .IN1(
        \SUMB[296][1] ), .COUT(\CARRYB[297][0] ), .SUM(PRODUCT[297]) );
  FADDER S2_297_1 ( .CIN(\ab[297][1] ), .IN0(\CARRYB[296][1] ), .IN1(
        \SUMB[296][2] ), .COUT(\CARRYB[297][1] ), .SUM(\SUMB[297][1] ) );
  FADDER S3_297_2 ( .CIN(\ab[297][2] ), .IN0(\CARRYB[296][2] ), .IN1(
        \ab[296][3] ), .COUT(\CARRYB[297][2] ), .SUM(\SUMB[297][2] ) );
  FADDER S1_296_0 ( .CIN(\ab[296][0] ), .IN0(\CARRYB[295][0] ), .IN1(
        \SUMB[295][1] ), .COUT(\CARRYB[296][0] ), .SUM(PRODUCT[296]) );
  FADDER S2_296_1 ( .CIN(\ab[296][1] ), .IN0(\CARRYB[295][1] ), .IN1(
        \SUMB[295][2] ), .COUT(\CARRYB[296][1] ), .SUM(\SUMB[296][1] ) );
  FADDER S3_296_2 ( .CIN(\ab[296][2] ), .IN0(\CARRYB[295][2] ), .IN1(
        \ab[295][3] ), .COUT(\CARRYB[296][2] ), .SUM(\SUMB[296][2] ) );
  FADDER S1_295_0 ( .CIN(\ab[295][0] ), .IN0(\CARRYB[294][0] ), .IN1(
        \SUMB[294][1] ), .COUT(\CARRYB[295][0] ), .SUM(PRODUCT[295]) );
  FADDER S2_295_1 ( .CIN(\ab[295][1] ), .IN0(\CARRYB[294][1] ), .IN1(
        \SUMB[294][2] ), .COUT(\CARRYB[295][1] ), .SUM(\SUMB[295][1] ) );
  FADDER S3_295_2 ( .CIN(\ab[295][2] ), .IN0(\CARRYB[294][2] ), .IN1(
        \ab[294][3] ), .COUT(\CARRYB[295][2] ), .SUM(\SUMB[295][2] ) );
  FADDER S1_294_0 ( .CIN(\ab[294][0] ), .IN0(\CARRYB[293][0] ), .IN1(
        \SUMB[293][1] ), .COUT(\CARRYB[294][0] ), .SUM(PRODUCT[294]) );
  FADDER S2_294_1 ( .CIN(\ab[294][1] ), .IN0(\CARRYB[293][1] ), .IN1(
        \SUMB[293][2] ), .COUT(\CARRYB[294][1] ), .SUM(\SUMB[294][1] ) );
  FADDER S3_294_2 ( .CIN(\ab[294][2] ), .IN0(\CARRYB[293][2] ), .IN1(
        \ab[293][3] ), .COUT(\CARRYB[294][2] ), .SUM(\SUMB[294][2] ) );
  FADDER S1_293_0 ( .CIN(\ab[293][0] ), .IN0(\CARRYB[292][0] ), .IN1(
        \SUMB[292][1] ), .COUT(\CARRYB[293][0] ), .SUM(PRODUCT[293]) );
  FADDER S2_293_1 ( .CIN(\ab[293][1] ), .IN0(\CARRYB[292][1] ), .IN1(
        \SUMB[292][2] ), .COUT(\CARRYB[293][1] ), .SUM(\SUMB[293][1] ) );
  FADDER S3_293_2 ( .CIN(\ab[293][2] ), .IN0(\CARRYB[292][2] ), .IN1(
        \ab[292][3] ), .COUT(\CARRYB[293][2] ), .SUM(\SUMB[293][2] ) );
  FADDER S1_292_0 ( .CIN(\ab[292][0] ), .IN0(\CARRYB[291][0] ), .IN1(
        \SUMB[291][1] ), .COUT(\CARRYB[292][0] ), .SUM(PRODUCT[292]) );
  FADDER S2_292_1 ( .CIN(\ab[292][1] ), .IN0(\CARRYB[291][1] ), .IN1(
        \SUMB[291][2] ), .COUT(\CARRYB[292][1] ), .SUM(\SUMB[292][1] ) );
  FADDER S3_292_2 ( .CIN(\ab[292][2] ), .IN0(\CARRYB[291][2] ), .IN1(
        \ab[291][3] ), .COUT(\CARRYB[292][2] ), .SUM(\SUMB[292][2] ) );
  FADDER S1_291_0 ( .CIN(\ab[291][0] ), .IN0(\CARRYB[290][0] ), .IN1(
        \SUMB[290][1] ), .COUT(\CARRYB[291][0] ), .SUM(PRODUCT[291]) );
  FADDER S2_291_1 ( .CIN(\ab[291][1] ), .IN0(\CARRYB[290][1] ), .IN1(
        \SUMB[290][2] ), .COUT(\CARRYB[291][1] ), .SUM(\SUMB[291][1] ) );
  FADDER S3_291_2 ( .CIN(\ab[291][2] ), .IN0(\CARRYB[290][2] ), .IN1(
        \ab[290][3] ), .COUT(\CARRYB[291][2] ), .SUM(\SUMB[291][2] ) );
  FADDER S1_290_0 ( .CIN(\ab[290][0] ), .IN0(\CARRYB[289][0] ), .IN1(
        \SUMB[289][1] ), .COUT(\CARRYB[290][0] ), .SUM(PRODUCT[290]) );
  FADDER S2_290_1 ( .CIN(\ab[290][1] ), .IN0(\CARRYB[289][1] ), .IN1(
        \SUMB[289][2] ), .COUT(\CARRYB[290][1] ), .SUM(\SUMB[290][1] ) );
  FADDER S3_290_2 ( .CIN(\ab[290][2] ), .IN0(\CARRYB[289][2] ), .IN1(
        \ab[289][3] ), .COUT(\CARRYB[290][2] ), .SUM(\SUMB[290][2] ) );
  FADDER S1_289_0 ( .CIN(\ab[289][0] ), .IN0(\CARRYB[288][0] ), .IN1(
        \SUMB[288][1] ), .COUT(\CARRYB[289][0] ), .SUM(PRODUCT[289]) );
  FADDER S2_289_1 ( .CIN(\ab[289][1] ), .IN0(\CARRYB[288][1] ), .IN1(
        \SUMB[288][2] ), .COUT(\CARRYB[289][1] ), .SUM(\SUMB[289][1] ) );
  FADDER S3_289_2 ( .CIN(\ab[289][2] ), .IN0(\CARRYB[288][2] ), .IN1(
        \ab[288][3] ), .COUT(\CARRYB[289][2] ), .SUM(\SUMB[289][2] ) );
  FADDER S1_288_0 ( .CIN(\ab[288][0] ), .IN0(\CARRYB[287][0] ), .IN1(
        \SUMB[287][1] ), .COUT(\CARRYB[288][0] ), .SUM(PRODUCT[288]) );
  FADDER S2_288_1 ( .CIN(\ab[288][1] ), .IN0(\CARRYB[287][1] ), .IN1(
        \SUMB[287][2] ), .COUT(\CARRYB[288][1] ), .SUM(\SUMB[288][1] ) );
  FADDER S3_288_2 ( .CIN(\ab[288][2] ), .IN0(\CARRYB[287][2] ), .IN1(
        \ab[287][3] ), .COUT(\CARRYB[288][2] ), .SUM(\SUMB[288][2] ) );
  FADDER S1_287_0 ( .CIN(\ab[287][0] ), .IN0(\CARRYB[286][0] ), .IN1(
        \SUMB[286][1] ), .COUT(\CARRYB[287][0] ), .SUM(PRODUCT[287]) );
  FADDER S2_287_1 ( .CIN(\ab[287][1] ), .IN0(\CARRYB[286][1] ), .IN1(
        \SUMB[286][2] ), .COUT(\CARRYB[287][1] ), .SUM(\SUMB[287][1] ) );
  FADDER S3_287_2 ( .CIN(\ab[287][2] ), .IN0(\CARRYB[286][2] ), .IN1(
        \ab[286][3] ), .COUT(\CARRYB[287][2] ), .SUM(\SUMB[287][2] ) );
  FADDER S1_286_0 ( .CIN(\ab[286][0] ), .IN0(\CARRYB[285][0] ), .IN1(
        \SUMB[285][1] ), .COUT(\CARRYB[286][0] ), .SUM(PRODUCT[286]) );
  FADDER S2_286_1 ( .CIN(\ab[286][1] ), .IN0(\CARRYB[285][1] ), .IN1(
        \SUMB[285][2] ), .COUT(\CARRYB[286][1] ), .SUM(\SUMB[286][1] ) );
  FADDER S3_286_2 ( .CIN(\ab[286][2] ), .IN0(\CARRYB[285][2] ), .IN1(
        \ab[285][3] ), .COUT(\CARRYB[286][2] ), .SUM(\SUMB[286][2] ) );
  FADDER S1_285_0 ( .CIN(\ab[285][0] ), .IN0(\CARRYB[284][0] ), .IN1(
        \SUMB[284][1] ), .COUT(\CARRYB[285][0] ), .SUM(PRODUCT[285]) );
  FADDER S2_285_1 ( .CIN(\ab[285][1] ), .IN0(\CARRYB[284][1] ), .IN1(
        \SUMB[284][2] ), .COUT(\CARRYB[285][1] ), .SUM(\SUMB[285][1] ) );
  FADDER S3_285_2 ( .CIN(\ab[285][2] ), .IN0(\CARRYB[284][2] ), .IN1(
        \ab[284][3] ), .COUT(\CARRYB[285][2] ), .SUM(\SUMB[285][2] ) );
  FADDER S1_284_0 ( .CIN(\ab[284][0] ), .IN0(\CARRYB[283][0] ), .IN1(
        \SUMB[283][1] ), .COUT(\CARRYB[284][0] ), .SUM(PRODUCT[284]) );
  FADDER S2_284_1 ( .CIN(\ab[284][1] ), .IN0(\CARRYB[283][1] ), .IN1(
        \SUMB[283][2] ), .COUT(\CARRYB[284][1] ), .SUM(\SUMB[284][1] ) );
  FADDER S3_284_2 ( .CIN(\ab[284][2] ), .IN0(\CARRYB[283][2] ), .IN1(
        \ab[283][3] ), .COUT(\CARRYB[284][2] ), .SUM(\SUMB[284][2] ) );
  FADDER S1_283_0 ( .CIN(\ab[283][0] ), .IN0(\CARRYB[282][0] ), .IN1(
        \SUMB[282][1] ), .COUT(\CARRYB[283][0] ), .SUM(PRODUCT[283]) );
  FADDER S2_283_1 ( .CIN(\ab[283][1] ), .IN0(\CARRYB[282][1] ), .IN1(
        \SUMB[282][2] ), .COUT(\CARRYB[283][1] ), .SUM(\SUMB[283][1] ) );
  FADDER S3_283_2 ( .CIN(\ab[283][2] ), .IN0(\CARRYB[282][2] ), .IN1(
        \ab[282][3] ), .COUT(\CARRYB[283][2] ), .SUM(\SUMB[283][2] ) );
  FADDER S1_282_0 ( .CIN(\ab[282][0] ), .IN0(\CARRYB[281][0] ), .IN1(
        \SUMB[281][1] ), .COUT(\CARRYB[282][0] ), .SUM(PRODUCT[282]) );
  FADDER S2_282_1 ( .CIN(\ab[282][1] ), .IN0(\CARRYB[281][1] ), .IN1(
        \SUMB[281][2] ), .COUT(\CARRYB[282][1] ), .SUM(\SUMB[282][1] ) );
  FADDER S3_282_2 ( .CIN(\ab[282][2] ), .IN0(\CARRYB[281][2] ), .IN1(
        \ab[281][3] ), .COUT(\CARRYB[282][2] ), .SUM(\SUMB[282][2] ) );
  FADDER S1_281_0 ( .CIN(\ab[281][0] ), .IN0(\CARRYB[280][0] ), .IN1(
        \SUMB[280][1] ), .COUT(\CARRYB[281][0] ), .SUM(PRODUCT[281]) );
  FADDER S2_281_1 ( .CIN(\ab[281][1] ), .IN0(\CARRYB[280][1] ), .IN1(
        \SUMB[280][2] ), .COUT(\CARRYB[281][1] ), .SUM(\SUMB[281][1] ) );
  FADDER S3_281_2 ( .CIN(\ab[281][2] ), .IN0(\CARRYB[280][2] ), .IN1(
        \ab[280][3] ), .COUT(\CARRYB[281][2] ), .SUM(\SUMB[281][2] ) );
  FADDER S1_280_0 ( .CIN(\ab[280][0] ), .IN0(\CARRYB[279][0] ), .IN1(
        \SUMB[279][1] ), .COUT(\CARRYB[280][0] ), .SUM(PRODUCT[280]) );
  FADDER S2_280_1 ( .CIN(\ab[280][1] ), .IN0(\CARRYB[279][1] ), .IN1(
        \SUMB[279][2] ), .COUT(\CARRYB[280][1] ), .SUM(\SUMB[280][1] ) );
  FADDER S3_280_2 ( .CIN(\ab[280][2] ), .IN0(\CARRYB[279][2] ), .IN1(
        \ab[279][3] ), .COUT(\CARRYB[280][2] ), .SUM(\SUMB[280][2] ) );
  FADDER S1_279_0 ( .CIN(\ab[279][0] ), .IN0(\CARRYB[278][0] ), .IN1(
        \SUMB[278][1] ), .COUT(\CARRYB[279][0] ), .SUM(PRODUCT[279]) );
  FADDER S2_279_1 ( .CIN(\ab[279][1] ), .IN0(\CARRYB[278][1] ), .IN1(
        \SUMB[278][2] ), .COUT(\CARRYB[279][1] ), .SUM(\SUMB[279][1] ) );
  FADDER S3_279_2 ( .CIN(\ab[279][2] ), .IN0(\CARRYB[278][2] ), .IN1(
        \ab[278][3] ), .COUT(\CARRYB[279][2] ), .SUM(\SUMB[279][2] ) );
  FADDER S1_278_0 ( .CIN(\ab[278][0] ), .IN0(\CARRYB[277][0] ), .IN1(
        \SUMB[277][1] ), .COUT(\CARRYB[278][0] ), .SUM(PRODUCT[278]) );
  FADDER S2_278_1 ( .CIN(\ab[278][1] ), .IN0(\CARRYB[277][1] ), .IN1(
        \SUMB[277][2] ), .COUT(\CARRYB[278][1] ), .SUM(\SUMB[278][1] ) );
  FADDER S3_278_2 ( .CIN(\ab[278][2] ), .IN0(\CARRYB[277][2] ), .IN1(
        \ab[277][3] ), .COUT(\CARRYB[278][2] ), .SUM(\SUMB[278][2] ) );
  FADDER S1_277_0 ( .CIN(\ab[277][0] ), .IN0(\CARRYB[276][0] ), .IN1(
        \SUMB[276][1] ), .COUT(\CARRYB[277][0] ), .SUM(PRODUCT[277]) );
  FADDER S2_277_1 ( .CIN(\ab[277][1] ), .IN0(\CARRYB[276][1] ), .IN1(
        \SUMB[276][2] ), .COUT(\CARRYB[277][1] ), .SUM(\SUMB[277][1] ) );
  FADDER S3_277_2 ( .CIN(\ab[277][2] ), .IN0(\CARRYB[276][2] ), .IN1(
        \ab[276][3] ), .COUT(\CARRYB[277][2] ), .SUM(\SUMB[277][2] ) );
  FADDER S1_276_0 ( .CIN(\ab[276][0] ), .IN0(\CARRYB[275][0] ), .IN1(
        \SUMB[275][1] ), .COUT(\CARRYB[276][0] ), .SUM(PRODUCT[276]) );
  FADDER S2_276_1 ( .CIN(\ab[276][1] ), .IN0(\CARRYB[275][1] ), .IN1(
        \SUMB[275][2] ), .COUT(\CARRYB[276][1] ), .SUM(\SUMB[276][1] ) );
  FADDER S3_276_2 ( .CIN(\ab[276][2] ), .IN0(\CARRYB[275][2] ), .IN1(
        \ab[275][3] ), .COUT(\CARRYB[276][2] ), .SUM(\SUMB[276][2] ) );
  FADDER S1_275_0 ( .CIN(\ab[275][0] ), .IN0(\CARRYB[274][0] ), .IN1(
        \SUMB[274][1] ), .COUT(\CARRYB[275][0] ), .SUM(PRODUCT[275]) );
  FADDER S2_275_1 ( .CIN(\ab[275][1] ), .IN0(\CARRYB[274][1] ), .IN1(
        \SUMB[274][2] ), .COUT(\CARRYB[275][1] ), .SUM(\SUMB[275][1] ) );
  FADDER S3_275_2 ( .CIN(\ab[275][2] ), .IN0(\CARRYB[274][2] ), .IN1(
        \ab[274][3] ), .COUT(\CARRYB[275][2] ), .SUM(\SUMB[275][2] ) );
  FADDER S1_274_0 ( .CIN(\ab[274][0] ), .IN0(\CARRYB[273][0] ), .IN1(
        \SUMB[273][1] ), .COUT(\CARRYB[274][0] ), .SUM(PRODUCT[274]) );
  FADDER S2_274_1 ( .CIN(\ab[274][1] ), .IN0(\CARRYB[273][1] ), .IN1(
        \SUMB[273][2] ), .COUT(\CARRYB[274][1] ), .SUM(\SUMB[274][1] ) );
  FADDER S3_274_2 ( .CIN(\ab[274][2] ), .IN0(\CARRYB[273][2] ), .IN1(
        \ab[273][3] ), .COUT(\CARRYB[274][2] ), .SUM(\SUMB[274][2] ) );
  FADDER S1_273_0 ( .CIN(\ab[273][0] ), .IN0(\CARRYB[272][0] ), .IN1(
        \SUMB[272][1] ), .COUT(\CARRYB[273][0] ), .SUM(PRODUCT[273]) );
  FADDER S2_273_1 ( .CIN(\ab[273][1] ), .IN0(\CARRYB[272][1] ), .IN1(
        \SUMB[272][2] ), .COUT(\CARRYB[273][1] ), .SUM(\SUMB[273][1] ) );
  FADDER S3_273_2 ( .CIN(\ab[273][2] ), .IN0(\CARRYB[272][2] ), .IN1(
        \ab[272][3] ), .COUT(\CARRYB[273][2] ), .SUM(\SUMB[273][2] ) );
  FADDER S1_272_0 ( .CIN(\ab[272][0] ), .IN0(\CARRYB[271][0] ), .IN1(
        \SUMB[271][1] ), .COUT(\CARRYB[272][0] ), .SUM(PRODUCT[272]) );
  FADDER S2_272_1 ( .CIN(\ab[272][1] ), .IN0(\CARRYB[271][1] ), .IN1(
        \SUMB[271][2] ), .COUT(\CARRYB[272][1] ), .SUM(\SUMB[272][1] ) );
  FADDER S3_272_2 ( .CIN(\ab[272][2] ), .IN0(\CARRYB[271][2] ), .IN1(
        \ab[271][3] ), .COUT(\CARRYB[272][2] ), .SUM(\SUMB[272][2] ) );
  FADDER S1_271_0 ( .CIN(\ab[271][0] ), .IN0(\CARRYB[270][0] ), .IN1(
        \SUMB[270][1] ), .COUT(\CARRYB[271][0] ), .SUM(PRODUCT[271]) );
  FADDER S2_271_1 ( .CIN(\ab[271][1] ), .IN0(\CARRYB[270][1] ), .IN1(
        \SUMB[270][2] ), .COUT(\CARRYB[271][1] ), .SUM(\SUMB[271][1] ) );
  FADDER S3_271_2 ( .CIN(\ab[271][2] ), .IN0(\CARRYB[270][2] ), .IN1(
        \ab[270][3] ), .COUT(\CARRYB[271][2] ), .SUM(\SUMB[271][2] ) );
  FADDER S1_270_0 ( .CIN(\ab[270][0] ), .IN0(\CARRYB[269][0] ), .IN1(
        \SUMB[269][1] ), .COUT(\CARRYB[270][0] ), .SUM(PRODUCT[270]) );
  FADDER S2_270_1 ( .CIN(\ab[270][1] ), .IN0(\CARRYB[269][1] ), .IN1(
        \SUMB[269][2] ), .COUT(\CARRYB[270][1] ), .SUM(\SUMB[270][1] ) );
  FADDER S3_270_2 ( .CIN(\ab[270][2] ), .IN0(\CARRYB[269][2] ), .IN1(
        \ab[269][3] ), .COUT(\CARRYB[270][2] ), .SUM(\SUMB[270][2] ) );
  FADDER S1_269_0 ( .CIN(\ab[269][0] ), .IN0(\CARRYB[268][0] ), .IN1(
        \SUMB[268][1] ), .COUT(\CARRYB[269][0] ), .SUM(PRODUCT[269]) );
  FADDER S2_269_1 ( .CIN(\ab[269][1] ), .IN0(\CARRYB[268][1] ), .IN1(
        \SUMB[268][2] ), .COUT(\CARRYB[269][1] ), .SUM(\SUMB[269][1] ) );
  FADDER S3_269_2 ( .CIN(\ab[269][2] ), .IN0(\CARRYB[268][2] ), .IN1(
        \ab[268][3] ), .COUT(\CARRYB[269][2] ), .SUM(\SUMB[269][2] ) );
  FADDER S1_268_0 ( .CIN(\ab[268][0] ), .IN0(\CARRYB[267][0] ), .IN1(
        \SUMB[267][1] ), .COUT(\CARRYB[268][0] ), .SUM(PRODUCT[268]) );
  FADDER S2_268_1 ( .CIN(\ab[268][1] ), .IN0(\CARRYB[267][1] ), .IN1(
        \SUMB[267][2] ), .COUT(\CARRYB[268][1] ), .SUM(\SUMB[268][1] ) );
  FADDER S3_268_2 ( .CIN(\ab[268][2] ), .IN0(\CARRYB[267][2] ), .IN1(
        \ab[267][3] ), .COUT(\CARRYB[268][2] ), .SUM(\SUMB[268][2] ) );
  FADDER S1_267_0 ( .CIN(\ab[267][0] ), .IN0(\CARRYB[266][0] ), .IN1(
        \SUMB[266][1] ), .COUT(\CARRYB[267][0] ), .SUM(PRODUCT[267]) );
  FADDER S2_267_1 ( .CIN(\ab[267][1] ), .IN0(\CARRYB[266][1] ), .IN1(
        \SUMB[266][2] ), .COUT(\CARRYB[267][1] ), .SUM(\SUMB[267][1] ) );
  FADDER S3_267_2 ( .CIN(\ab[267][2] ), .IN0(\CARRYB[266][2] ), .IN1(
        \ab[266][3] ), .COUT(\CARRYB[267][2] ), .SUM(\SUMB[267][2] ) );
  FADDER S1_266_0 ( .CIN(\ab[266][0] ), .IN0(\CARRYB[265][0] ), .IN1(
        \SUMB[265][1] ), .COUT(\CARRYB[266][0] ), .SUM(PRODUCT[266]) );
  FADDER S2_266_1 ( .CIN(\ab[266][1] ), .IN0(\CARRYB[265][1] ), .IN1(
        \SUMB[265][2] ), .COUT(\CARRYB[266][1] ), .SUM(\SUMB[266][1] ) );
  FADDER S3_266_2 ( .CIN(\ab[266][2] ), .IN0(\CARRYB[265][2] ), .IN1(
        \ab[265][3] ), .COUT(\CARRYB[266][2] ), .SUM(\SUMB[266][2] ) );
  FADDER S1_265_0 ( .CIN(\ab[265][0] ), .IN0(\CARRYB[264][0] ), .IN1(
        \SUMB[264][1] ), .COUT(\CARRYB[265][0] ), .SUM(PRODUCT[265]) );
  FADDER S2_265_1 ( .CIN(\ab[265][1] ), .IN0(\CARRYB[264][1] ), .IN1(
        \SUMB[264][2] ), .COUT(\CARRYB[265][1] ), .SUM(\SUMB[265][1] ) );
  FADDER S3_265_2 ( .CIN(\ab[265][2] ), .IN0(\CARRYB[264][2] ), .IN1(
        \ab[264][3] ), .COUT(\CARRYB[265][2] ), .SUM(\SUMB[265][2] ) );
  FADDER S1_264_0 ( .CIN(\ab[264][0] ), .IN0(\CARRYB[263][0] ), .IN1(
        \SUMB[263][1] ), .COUT(\CARRYB[264][0] ), .SUM(PRODUCT[264]) );
  FADDER S2_264_1 ( .CIN(\ab[264][1] ), .IN0(\CARRYB[263][1] ), .IN1(
        \SUMB[263][2] ), .COUT(\CARRYB[264][1] ), .SUM(\SUMB[264][1] ) );
  FADDER S3_264_2 ( .CIN(\ab[264][2] ), .IN0(\CARRYB[263][2] ), .IN1(
        \ab[263][3] ), .COUT(\CARRYB[264][2] ), .SUM(\SUMB[264][2] ) );
  FADDER S1_263_0 ( .CIN(\ab[263][0] ), .IN0(\CARRYB[262][0] ), .IN1(
        \SUMB[262][1] ), .COUT(\CARRYB[263][0] ), .SUM(PRODUCT[263]) );
  FADDER S2_263_1 ( .CIN(\ab[263][1] ), .IN0(\CARRYB[262][1] ), .IN1(
        \SUMB[262][2] ), .COUT(\CARRYB[263][1] ), .SUM(\SUMB[263][1] ) );
  FADDER S3_263_2 ( .CIN(\ab[263][2] ), .IN0(\CARRYB[262][2] ), .IN1(
        \ab[262][3] ), .COUT(\CARRYB[263][2] ), .SUM(\SUMB[263][2] ) );
  FADDER S1_262_0 ( .CIN(\ab[262][0] ), .IN0(\CARRYB[261][0] ), .IN1(
        \SUMB[261][1] ), .COUT(\CARRYB[262][0] ), .SUM(PRODUCT[262]) );
  FADDER S2_262_1 ( .CIN(\ab[262][1] ), .IN0(\CARRYB[261][1] ), .IN1(
        \SUMB[261][2] ), .COUT(\CARRYB[262][1] ), .SUM(\SUMB[262][1] ) );
  FADDER S3_262_2 ( .CIN(\ab[262][2] ), .IN0(\CARRYB[261][2] ), .IN1(
        \ab[261][3] ), .COUT(\CARRYB[262][2] ), .SUM(\SUMB[262][2] ) );
  FADDER S1_261_0 ( .CIN(\ab[261][0] ), .IN0(\CARRYB[260][0] ), .IN1(
        \SUMB[260][1] ), .COUT(\CARRYB[261][0] ), .SUM(PRODUCT[261]) );
  FADDER S2_261_1 ( .CIN(\ab[261][1] ), .IN0(\CARRYB[260][1] ), .IN1(
        \SUMB[260][2] ), .COUT(\CARRYB[261][1] ), .SUM(\SUMB[261][1] ) );
  FADDER S3_261_2 ( .CIN(\ab[261][2] ), .IN0(\CARRYB[260][2] ), .IN1(
        \ab[260][3] ), .COUT(\CARRYB[261][2] ), .SUM(\SUMB[261][2] ) );
  FADDER S1_260_0 ( .CIN(\ab[260][0] ), .IN0(\CARRYB[259][0] ), .IN1(
        \SUMB[259][1] ), .COUT(\CARRYB[260][0] ), .SUM(PRODUCT[260]) );
  FADDER S2_260_1 ( .CIN(\ab[260][1] ), .IN0(\CARRYB[259][1] ), .IN1(
        \SUMB[259][2] ), .COUT(\CARRYB[260][1] ), .SUM(\SUMB[260][1] ) );
  FADDER S3_260_2 ( .CIN(\ab[260][2] ), .IN0(\CARRYB[259][2] ), .IN1(
        \ab[259][3] ), .COUT(\CARRYB[260][2] ), .SUM(\SUMB[260][2] ) );
  FADDER S1_259_0 ( .CIN(\ab[259][0] ), .IN0(\CARRYB[258][0] ), .IN1(
        \SUMB[258][1] ), .COUT(\CARRYB[259][0] ), .SUM(PRODUCT[259]) );
  FADDER S2_259_1 ( .CIN(\ab[259][1] ), .IN0(\CARRYB[258][1] ), .IN1(
        \SUMB[258][2] ), .COUT(\CARRYB[259][1] ), .SUM(\SUMB[259][1] ) );
  FADDER S3_259_2 ( .CIN(\ab[259][2] ), .IN0(\CARRYB[258][2] ), .IN1(
        \ab[258][3] ), .COUT(\CARRYB[259][2] ), .SUM(\SUMB[259][2] ) );
  FADDER S1_258_0 ( .CIN(\ab[258][0] ), .IN0(\CARRYB[257][0] ), .IN1(
        \SUMB[257][1] ), .COUT(\CARRYB[258][0] ), .SUM(PRODUCT[258]) );
  FADDER S2_258_1 ( .CIN(\ab[258][1] ), .IN0(\CARRYB[257][1] ), .IN1(
        \SUMB[257][2] ), .COUT(\CARRYB[258][1] ), .SUM(\SUMB[258][1] ) );
  FADDER S3_258_2 ( .CIN(\ab[258][2] ), .IN0(\CARRYB[257][2] ), .IN1(
        \ab[257][3] ), .COUT(\CARRYB[258][2] ), .SUM(\SUMB[258][2] ) );
  FADDER S1_257_0 ( .CIN(\ab[257][0] ), .IN0(\CARRYB[256][0] ), .IN1(
        \SUMB[256][1] ), .COUT(\CARRYB[257][0] ), .SUM(PRODUCT[257]) );
  FADDER S2_257_1 ( .CIN(\ab[257][1] ), .IN0(\CARRYB[256][1] ), .IN1(
        \SUMB[256][2] ), .COUT(\CARRYB[257][1] ), .SUM(\SUMB[257][1] ) );
  FADDER S3_257_2 ( .CIN(\ab[257][2] ), .IN0(\CARRYB[256][2] ), .IN1(
        \ab[256][3] ), .COUT(\CARRYB[257][2] ), .SUM(\SUMB[257][2] ) );
  FADDER S1_256_0 ( .CIN(\ab[256][0] ), .IN0(\CARRYB[255][0] ), .IN1(
        \SUMB[255][1] ), .COUT(\CARRYB[256][0] ), .SUM(PRODUCT[256]) );
  FADDER S2_256_1 ( .CIN(\ab[256][1] ), .IN0(\CARRYB[255][1] ), .IN1(
        \SUMB[255][2] ), .COUT(\CARRYB[256][1] ), .SUM(\SUMB[256][1] ) );
  FADDER S3_256_2 ( .CIN(\ab[256][2] ), .IN0(\CARRYB[255][2] ), .IN1(
        \ab[255][3] ), .COUT(\CARRYB[256][2] ), .SUM(\SUMB[256][2] ) );
  FADDER S1_255_0 ( .CIN(\ab[255][0] ), .IN0(\CARRYB[254][0] ), .IN1(
        \SUMB[254][1] ), .COUT(\CARRYB[255][0] ), .SUM(PRODUCT[255]) );
  FADDER S2_255_1 ( .CIN(\ab[255][1] ), .IN0(\CARRYB[254][1] ), .IN1(
        \SUMB[254][2] ), .COUT(\CARRYB[255][1] ), .SUM(\SUMB[255][1] ) );
  FADDER S3_255_2 ( .CIN(\ab[255][2] ), .IN0(\CARRYB[254][2] ), .IN1(
        \ab[254][3] ), .COUT(\CARRYB[255][2] ), .SUM(\SUMB[255][2] ) );
  FADDER S1_254_0 ( .CIN(\ab[254][0] ), .IN0(\CARRYB[253][0] ), .IN1(
        \SUMB[253][1] ), .COUT(\CARRYB[254][0] ), .SUM(PRODUCT[254]) );
  FADDER S2_254_1 ( .CIN(\ab[254][1] ), .IN0(\CARRYB[253][1] ), .IN1(
        \SUMB[253][2] ), .COUT(\CARRYB[254][1] ), .SUM(\SUMB[254][1] ) );
  FADDER S3_254_2 ( .CIN(\ab[254][2] ), .IN0(\CARRYB[253][2] ), .IN1(
        \ab[253][3] ), .COUT(\CARRYB[254][2] ), .SUM(\SUMB[254][2] ) );
  FADDER S1_253_0 ( .CIN(\ab[253][0] ), .IN0(\CARRYB[252][0] ), .IN1(
        \SUMB[252][1] ), .COUT(\CARRYB[253][0] ), .SUM(PRODUCT[253]) );
  FADDER S2_253_1 ( .CIN(\ab[253][1] ), .IN0(\CARRYB[252][1] ), .IN1(
        \SUMB[252][2] ), .COUT(\CARRYB[253][1] ), .SUM(\SUMB[253][1] ) );
  FADDER S3_253_2 ( .CIN(\ab[253][2] ), .IN0(\CARRYB[252][2] ), .IN1(
        \ab[252][3] ), .COUT(\CARRYB[253][2] ), .SUM(\SUMB[253][2] ) );
  FADDER S1_252_0 ( .CIN(\ab[252][0] ), .IN0(\CARRYB[251][0] ), .IN1(
        \SUMB[251][1] ), .COUT(\CARRYB[252][0] ), .SUM(PRODUCT[252]) );
  FADDER S2_252_1 ( .CIN(\ab[252][1] ), .IN0(\CARRYB[251][1] ), .IN1(
        \SUMB[251][2] ), .COUT(\CARRYB[252][1] ), .SUM(\SUMB[252][1] ) );
  FADDER S3_252_2 ( .CIN(\ab[252][2] ), .IN0(\CARRYB[251][2] ), .IN1(
        \ab[251][3] ), .COUT(\CARRYB[252][2] ), .SUM(\SUMB[252][2] ) );
  FADDER S1_251_0 ( .CIN(\ab[251][0] ), .IN0(\CARRYB[250][0] ), .IN1(
        \SUMB[250][1] ), .COUT(\CARRYB[251][0] ), .SUM(PRODUCT[251]) );
  FADDER S2_251_1 ( .CIN(\ab[251][1] ), .IN0(\CARRYB[250][1] ), .IN1(
        \SUMB[250][2] ), .COUT(\CARRYB[251][1] ), .SUM(\SUMB[251][1] ) );
  FADDER S3_251_2 ( .CIN(\ab[251][2] ), .IN0(\CARRYB[250][2] ), .IN1(
        \ab[250][3] ), .COUT(\CARRYB[251][2] ), .SUM(\SUMB[251][2] ) );
  FADDER S1_250_0 ( .CIN(\ab[250][0] ), .IN0(\CARRYB[249][0] ), .IN1(
        \SUMB[249][1] ), .COUT(\CARRYB[250][0] ), .SUM(PRODUCT[250]) );
  FADDER S2_250_1 ( .CIN(\ab[250][1] ), .IN0(\CARRYB[249][1] ), .IN1(
        \SUMB[249][2] ), .COUT(\CARRYB[250][1] ), .SUM(\SUMB[250][1] ) );
  FADDER S3_250_2 ( .CIN(\ab[250][2] ), .IN0(\CARRYB[249][2] ), .IN1(
        \ab[249][3] ), .COUT(\CARRYB[250][2] ), .SUM(\SUMB[250][2] ) );
  FADDER S1_249_0 ( .CIN(\ab[249][0] ), .IN0(\CARRYB[248][0] ), .IN1(
        \SUMB[248][1] ), .COUT(\CARRYB[249][0] ), .SUM(PRODUCT[249]) );
  FADDER S2_249_1 ( .CIN(\ab[249][1] ), .IN0(\CARRYB[248][1] ), .IN1(
        \SUMB[248][2] ), .COUT(\CARRYB[249][1] ), .SUM(\SUMB[249][1] ) );
  FADDER S3_249_2 ( .CIN(\ab[249][2] ), .IN0(\CARRYB[248][2] ), .IN1(
        \ab[248][3] ), .COUT(\CARRYB[249][2] ), .SUM(\SUMB[249][2] ) );
  FADDER S1_248_0 ( .CIN(\ab[248][0] ), .IN0(\CARRYB[247][0] ), .IN1(
        \SUMB[247][1] ), .COUT(\CARRYB[248][0] ), .SUM(PRODUCT[248]) );
  FADDER S2_248_1 ( .CIN(\ab[248][1] ), .IN0(\CARRYB[247][1] ), .IN1(
        \SUMB[247][2] ), .COUT(\CARRYB[248][1] ), .SUM(\SUMB[248][1] ) );
  FADDER S3_248_2 ( .CIN(\ab[248][2] ), .IN0(\CARRYB[247][2] ), .IN1(
        \ab[247][3] ), .COUT(\CARRYB[248][2] ), .SUM(\SUMB[248][2] ) );
  FADDER S1_247_0 ( .CIN(\ab[247][0] ), .IN0(\CARRYB[246][0] ), .IN1(
        \SUMB[246][1] ), .COUT(\CARRYB[247][0] ), .SUM(PRODUCT[247]) );
  FADDER S2_247_1 ( .CIN(\ab[247][1] ), .IN0(\CARRYB[246][1] ), .IN1(
        \SUMB[246][2] ), .COUT(\CARRYB[247][1] ), .SUM(\SUMB[247][1] ) );
  FADDER S3_247_2 ( .CIN(\ab[247][2] ), .IN0(\CARRYB[246][2] ), .IN1(
        \ab[246][3] ), .COUT(\CARRYB[247][2] ), .SUM(\SUMB[247][2] ) );
  FADDER S1_246_0 ( .CIN(\ab[246][0] ), .IN0(\CARRYB[245][0] ), .IN1(
        \SUMB[245][1] ), .COUT(\CARRYB[246][0] ), .SUM(PRODUCT[246]) );
  FADDER S2_246_1 ( .CIN(\ab[246][1] ), .IN0(\CARRYB[245][1] ), .IN1(
        \SUMB[245][2] ), .COUT(\CARRYB[246][1] ), .SUM(\SUMB[246][1] ) );
  FADDER S3_246_2 ( .CIN(\ab[246][2] ), .IN0(\CARRYB[245][2] ), .IN1(
        \ab[245][3] ), .COUT(\CARRYB[246][2] ), .SUM(\SUMB[246][2] ) );
  FADDER S1_245_0 ( .CIN(\ab[245][0] ), .IN0(\CARRYB[244][0] ), .IN1(
        \SUMB[244][1] ), .COUT(\CARRYB[245][0] ), .SUM(PRODUCT[245]) );
  FADDER S2_245_1 ( .CIN(\ab[245][1] ), .IN0(\CARRYB[244][1] ), .IN1(
        \SUMB[244][2] ), .COUT(\CARRYB[245][1] ), .SUM(\SUMB[245][1] ) );
  FADDER S3_245_2 ( .CIN(\ab[245][2] ), .IN0(\CARRYB[244][2] ), .IN1(
        \ab[244][3] ), .COUT(\CARRYB[245][2] ), .SUM(\SUMB[245][2] ) );
  FADDER S1_244_0 ( .CIN(\ab[244][0] ), .IN0(\CARRYB[243][0] ), .IN1(
        \SUMB[243][1] ), .COUT(\CARRYB[244][0] ), .SUM(PRODUCT[244]) );
  FADDER S2_244_1 ( .CIN(\ab[244][1] ), .IN0(\CARRYB[243][1] ), .IN1(
        \SUMB[243][2] ), .COUT(\CARRYB[244][1] ), .SUM(\SUMB[244][1] ) );
  FADDER S3_244_2 ( .CIN(\ab[244][2] ), .IN0(\CARRYB[243][2] ), .IN1(
        \ab[243][3] ), .COUT(\CARRYB[244][2] ), .SUM(\SUMB[244][2] ) );
  FADDER S1_243_0 ( .CIN(\ab[243][0] ), .IN0(\CARRYB[242][0] ), .IN1(
        \SUMB[242][1] ), .COUT(\CARRYB[243][0] ), .SUM(PRODUCT[243]) );
  FADDER S2_243_1 ( .CIN(\ab[243][1] ), .IN0(\CARRYB[242][1] ), .IN1(
        \SUMB[242][2] ), .COUT(\CARRYB[243][1] ), .SUM(\SUMB[243][1] ) );
  FADDER S3_243_2 ( .CIN(\ab[243][2] ), .IN0(\CARRYB[242][2] ), .IN1(
        \ab[242][3] ), .COUT(\CARRYB[243][2] ), .SUM(\SUMB[243][2] ) );
  FADDER S1_242_0 ( .CIN(\ab[242][0] ), .IN0(\CARRYB[241][0] ), .IN1(
        \SUMB[241][1] ), .COUT(\CARRYB[242][0] ), .SUM(PRODUCT[242]) );
  FADDER S2_242_1 ( .CIN(\ab[242][1] ), .IN0(\CARRYB[241][1] ), .IN1(
        \SUMB[241][2] ), .COUT(\CARRYB[242][1] ), .SUM(\SUMB[242][1] ) );
  FADDER S3_242_2 ( .CIN(\ab[242][2] ), .IN0(\CARRYB[241][2] ), .IN1(
        \ab[241][3] ), .COUT(\CARRYB[242][2] ), .SUM(\SUMB[242][2] ) );
  FADDER S1_241_0 ( .CIN(\ab[241][0] ), .IN0(\CARRYB[240][0] ), .IN1(
        \SUMB[240][1] ), .COUT(\CARRYB[241][0] ), .SUM(PRODUCT[241]) );
  FADDER S2_241_1 ( .CIN(\ab[241][1] ), .IN0(\CARRYB[240][1] ), .IN1(
        \SUMB[240][2] ), .COUT(\CARRYB[241][1] ), .SUM(\SUMB[241][1] ) );
  FADDER S3_241_2 ( .CIN(\ab[241][2] ), .IN0(\CARRYB[240][2] ), .IN1(
        \ab[240][3] ), .COUT(\CARRYB[241][2] ), .SUM(\SUMB[241][2] ) );
  FADDER S1_240_0 ( .CIN(\ab[240][0] ), .IN0(\CARRYB[239][0] ), .IN1(
        \SUMB[239][1] ), .COUT(\CARRYB[240][0] ), .SUM(PRODUCT[240]) );
  FADDER S2_240_1 ( .CIN(\ab[240][1] ), .IN0(\CARRYB[239][1] ), .IN1(
        \SUMB[239][2] ), .COUT(\CARRYB[240][1] ), .SUM(\SUMB[240][1] ) );
  FADDER S3_240_2 ( .CIN(\ab[240][2] ), .IN0(\CARRYB[239][2] ), .IN1(
        \ab[239][3] ), .COUT(\CARRYB[240][2] ), .SUM(\SUMB[240][2] ) );
  FADDER S1_239_0 ( .CIN(\ab[239][0] ), .IN0(\CARRYB[238][0] ), .IN1(
        \SUMB[238][1] ), .COUT(\CARRYB[239][0] ), .SUM(PRODUCT[239]) );
  FADDER S2_239_1 ( .CIN(\ab[239][1] ), .IN0(\CARRYB[238][1] ), .IN1(
        \SUMB[238][2] ), .COUT(\CARRYB[239][1] ), .SUM(\SUMB[239][1] ) );
  FADDER S3_239_2 ( .CIN(\ab[239][2] ), .IN0(\CARRYB[238][2] ), .IN1(
        \ab[238][3] ), .COUT(\CARRYB[239][2] ), .SUM(\SUMB[239][2] ) );
  FADDER S1_238_0 ( .CIN(\ab[238][0] ), .IN0(\CARRYB[237][0] ), .IN1(
        \SUMB[237][1] ), .COUT(\CARRYB[238][0] ), .SUM(PRODUCT[238]) );
  FADDER S2_238_1 ( .CIN(\ab[238][1] ), .IN0(\CARRYB[237][1] ), .IN1(
        \SUMB[237][2] ), .COUT(\CARRYB[238][1] ), .SUM(\SUMB[238][1] ) );
  FADDER S3_238_2 ( .CIN(\ab[238][2] ), .IN0(\CARRYB[237][2] ), .IN1(
        \ab[237][3] ), .COUT(\CARRYB[238][2] ), .SUM(\SUMB[238][2] ) );
  FADDER S1_237_0 ( .CIN(\ab[237][0] ), .IN0(\CARRYB[236][0] ), .IN1(
        \SUMB[236][1] ), .COUT(\CARRYB[237][0] ), .SUM(PRODUCT[237]) );
  FADDER S2_237_1 ( .CIN(\ab[237][1] ), .IN0(\CARRYB[236][1] ), .IN1(
        \SUMB[236][2] ), .COUT(\CARRYB[237][1] ), .SUM(\SUMB[237][1] ) );
  FADDER S3_237_2 ( .CIN(\ab[237][2] ), .IN0(\CARRYB[236][2] ), .IN1(
        \ab[236][3] ), .COUT(\CARRYB[237][2] ), .SUM(\SUMB[237][2] ) );
  FADDER S1_236_0 ( .CIN(\ab[236][0] ), .IN0(\CARRYB[235][0] ), .IN1(
        \SUMB[235][1] ), .COUT(\CARRYB[236][0] ), .SUM(PRODUCT[236]) );
  FADDER S2_236_1 ( .CIN(\ab[236][1] ), .IN0(\CARRYB[235][1] ), .IN1(
        \SUMB[235][2] ), .COUT(\CARRYB[236][1] ), .SUM(\SUMB[236][1] ) );
  FADDER S3_236_2 ( .CIN(\ab[236][2] ), .IN0(\CARRYB[235][2] ), .IN1(
        \ab[235][3] ), .COUT(\CARRYB[236][2] ), .SUM(\SUMB[236][2] ) );
  FADDER S1_235_0 ( .CIN(\ab[235][0] ), .IN0(\CARRYB[234][0] ), .IN1(
        \SUMB[234][1] ), .COUT(\CARRYB[235][0] ), .SUM(PRODUCT[235]) );
  FADDER S2_235_1 ( .CIN(\ab[235][1] ), .IN0(\CARRYB[234][1] ), .IN1(
        \SUMB[234][2] ), .COUT(\CARRYB[235][1] ), .SUM(\SUMB[235][1] ) );
  FADDER S3_235_2 ( .CIN(\ab[235][2] ), .IN0(\CARRYB[234][2] ), .IN1(
        \ab[234][3] ), .COUT(\CARRYB[235][2] ), .SUM(\SUMB[235][2] ) );
  FADDER S1_234_0 ( .CIN(\ab[234][0] ), .IN0(\CARRYB[233][0] ), .IN1(
        \SUMB[233][1] ), .COUT(\CARRYB[234][0] ), .SUM(PRODUCT[234]) );
  FADDER S2_234_1 ( .CIN(\ab[234][1] ), .IN0(\CARRYB[233][1] ), .IN1(
        \SUMB[233][2] ), .COUT(\CARRYB[234][1] ), .SUM(\SUMB[234][1] ) );
  FADDER S3_234_2 ( .CIN(\ab[234][2] ), .IN0(\CARRYB[233][2] ), .IN1(
        \ab[233][3] ), .COUT(\CARRYB[234][2] ), .SUM(\SUMB[234][2] ) );
  FADDER S1_233_0 ( .CIN(\ab[233][0] ), .IN0(\CARRYB[232][0] ), .IN1(
        \SUMB[232][1] ), .COUT(\CARRYB[233][0] ), .SUM(PRODUCT[233]) );
  FADDER S2_233_1 ( .CIN(\ab[233][1] ), .IN0(\CARRYB[232][1] ), .IN1(
        \SUMB[232][2] ), .COUT(\CARRYB[233][1] ), .SUM(\SUMB[233][1] ) );
  FADDER S3_233_2 ( .CIN(\ab[233][2] ), .IN0(\CARRYB[232][2] ), .IN1(
        \ab[232][3] ), .COUT(\CARRYB[233][2] ), .SUM(\SUMB[233][2] ) );
  FADDER S1_232_0 ( .CIN(\ab[232][0] ), .IN0(\CARRYB[231][0] ), .IN1(
        \SUMB[231][1] ), .COUT(\CARRYB[232][0] ), .SUM(PRODUCT[232]) );
  FADDER S2_232_1 ( .CIN(\ab[232][1] ), .IN0(\CARRYB[231][1] ), .IN1(
        \SUMB[231][2] ), .COUT(\CARRYB[232][1] ), .SUM(\SUMB[232][1] ) );
  FADDER S3_232_2 ( .CIN(\ab[232][2] ), .IN0(\CARRYB[231][2] ), .IN1(
        \ab[231][3] ), .COUT(\CARRYB[232][2] ), .SUM(\SUMB[232][2] ) );
  FADDER S1_231_0 ( .CIN(\ab[231][0] ), .IN0(\CARRYB[230][0] ), .IN1(
        \SUMB[230][1] ), .COUT(\CARRYB[231][0] ), .SUM(PRODUCT[231]) );
  FADDER S2_231_1 ( .CIN(\ab[231][1] ), .IN0(\CARRYB[230][1] ), .IN1(
        \SUMB[230][2] ), .COUT(\CARRYB[231][1] ), .SUM(\SUMB[231][1] ) );
  FADDER S3_231_2 ( .CIN(\ab[231][2] ), .IN0(\CARRYB[230][2] ), .IN1(
        \ab[230][3] ), .COUT(\CARRYB[231][2] ), .SUM(\SUMB[231][2] ) );
  FADDER S1_230_0 ( .CIN(\ab[230][0] ), .IN0(\CARRYB[229][0] ), .IN1(
        \SUMB[229][1] ), .COUT(\CARRYB[230][0] ), .SUM(PRODUCT[230]) );
  FADDER S2_230_1 ( .CIN(\ab[230][1] ), .IN0(\CARRYB[229][1] ), .IN1(
        \SUMB[229][2] ), .COUT(\CARRYB[230][1] ), .SUM(\SUMB[230][1] ) );
  FADDER S3_230_2 ( .CIN(\ab[230][2] ), .IN0(\CARRYB[229][2] ), .IN1(
        \ab[229][3] ), .COUT(\CARRYB[230][2] ), .SUM(\SUMB[230][2] ) );
  FADDER S1_229_0 ( .CIN(\ab[229][0] ), .IN0(\CARRYB[228][0] ), .IN1(
        \SUMB[228][1] ), .COUT(\CARRYB[229][0] ), .SUM(PRODUCT[229]) );
  FADDER S2_229_1 ( .CIN(\ab[229][1] ), .IN0(\CARRYB[228][1] ), .IN1(
        \SUMB[228][2] ), .COUT(\CARRYB[229][1] ), .SUM(\SUMB[229][1] ) );
  FADDER S3_229_2 ( .CIN(\ab[229][2] ), .IN0(\CARRYB[228][2] ), .IN1(
        \ab[228][3] ), .COUT(\CARRYB[229][2] ), .SUM(\SUMB[229][2] ) );
  FADDER S1_228_0 ( .CIN(\ab[228][0] ), .IN0(\CARRYB[227][0] ), .IN1(
        \SUMB[227][1] ), .COUT(\CARRYB[228][0] ), .SUM(PRODUCT[228]) );
  FADDER S2_228_1 ( .CIN(\ab[228][1] ), .IN0(\CARRYB[227][1] ), .IN1(
        \SUMB[227][2] ), .COUT(\CARRYB[228][1] ), .SUM(\SUMB[228][1] ) );
  FADDER S3_228_2 ( .CIN(\ab[228][2] ), .IN0(\CARRYB[227][2] ), .IN1(
        \ab[227][3] ), .COUT(\CARRYB[228][2] ), .SUM(\SUMB[228][2] ) );
  FADDER S1_227_0 ( .CIN(\ab[227][0] ), .IN0(\CARRYB[226][0] ), .IN1(
        \SUMB[226][1] ), .COUT(\CARRYB[227][0] ), .SUM(PRODUCT[227]) );
  FADDER S2_227_1 ( .CIN(\ab[227][1] ), .IN0(\CARRYB[226][1] ), .IN1(
        \SUMB[226][2] ), .COUT(\CARRYB[227][1] ), .SUM(\SUMB[227][1] ) );
  FADDER S3_227_2 ( .CIN(\ab[227][2] ), .IN0(\CARRYB[226][2] ), .IN1(
        \ab[226][3] ), .COUT(\CARRYB[227][2] ), .SUM(\SUMB[227][2] ) );
  FADDER S1_226_0 ( .CIN(\ab[226][0] ), .IN0(\CARRYB[225][0] ), .IN1(
        \SUMB[225][1] ), .COUT(\CARRYB[226][0] ), .SUM(PRODUCT[226]) );
  FADDER S2_226_1 ( .CIN(\ab[226][1] ), .IN0(\CARRYB[225][1] ), .IN1(
        \SUMB[225][2] ), .COUT(\CARRYB[226][1] ), .SUM(\SUMB[226][1] ) );
  FADDER S3_226_2 ( .CIN(\ab[226][2] ), .IN0(\CARRYB[225][2] ), .IN1(
        \ab[225][3] ), .COUT(\CARRYB[226][2] ), .SUM(\SUMB[226][2] ) );
  FADDER S1_225_0 ( .CIN(\ab[225][0] ), .IN0(\CARRYB[224][0] ), .IN1(
        \SUMB[224][1] ), .COUT(\CARRYB[225][0] ), .SUM(PRODUCT[225]) );
  FADDER S2_225_1 ( .CIN(\ab[225][1] ), .IN0(\CARRYB[224][1] ), .IN1(
        \SUMB[224][2] ), .COUT(\CARRYB[225][1] ), .SUM(\SUMB[225][1] ) );
  FADDER S3_225_2 ( .CIN(\ab[225][2] ), .IN0(\CARRYB[224][2] ), .IN1(
        \ab[224][3] ), .COUT(\CARRYB[225][2] ), .SUM(\SUMB[225][2] ) );
  FADDER S1_224_0 ( .CIN(\ab[224][0] ), .IN0(\CARRYB[223][0] ), .IN1(
        \SUMB[223][1] ), .COUT(\CARRYB[224][0] ), .SUM(PRODUCT[224]) );
  FADDER S2_224_1 ( .CIN(\ab[224][1] ), .IN0(\CARRYB[223][1] ), .IN1(
        \SUMB[223][2] ), .COUT(\CARRYB[224][1] ), .SUM(\SUMB[224][1] ) );
  FADDER S3_224_2 ( .CIN(\ab[224][2] ), .IN0(\CARRYB[223][2] ), .IN1(
        \ab[223][3] ), .COUT(\CARRYB[224][2] ), .SUM(\SUMB[224][2] ) );
  FADDER S1_223_0 ( .CIN(\ab[223][0] ), .IN0(\CARRYB[222][0] ), .IN1(
        \SUMB[222][1] ), .COUT(\CARRYB[223][0] ), .SUM(PRODUCT[223]) );
  FADDER S2_223_1 ( .CIN(\ab[223][1] ), .IN0(\CARRYB[222][1] ), .IN1(
        \SUMB[222][2] ), .COUT(\CARRYB[223][1] ), .SUM(\SUMB[223][1] ) );
  FADDER S3_223_2 ( .CIN(\ab[223][2] ), .IN0(\CARRYB[222][2] ), .IN1(
        \ab[222][3] ), .COUT(\CARRYB[223][2] ), .SUM(\SUMB[223][2] ) );
  FADDER S1_222_0 ( .CIN(\ab[222][0] ), .IN0(\CARRYB[221][0] ), .IN1(
        \SUMB[221][1] ), .COUT(\CARRYB[222][0] ), .SUM(PRODUCT[222]) );
  FADDER S2_222_1 ( .CIN(\ab[222][1] ), .IN0(\CARRYB[221][1] ), .IN1(
        \SUMB[221][2] ), .COUT(\CARRYB[222][1] ), .SUM(\SUMB[222][1] ) );
  FADDER S3_222_2 ( .CIN(\ab[222][2] ), .IN0(\CARRYB[221][2] ), .IN1(
        \ab[221][3] ), .COUT(\CARRYB[222][2] ), .SUM(\SUMB[222][2] ) );
  FADDER S1_221_0 ( .CIN(\ab[221][0] ), .IN0(\CARRYB[220][0] ), .IN1(
        \SUMB[220][1] ), .COUT(\CARRYB[221][0] ), .SUM(PRODUCT[221]) );
  FADDER S2_221_1 ( .CIN(\ab[221][1] ), .IN0(\CARRYB[220][1] ), .IN1(
        \SUMB[220][2] ), .COUT(\CARRYB[221][1] ), .SUM(\SUMB[221][1] ) );
  FADDER S3_221_2 ( .CIN(\ab[221][2] ), .IN0(\CARRYB[220][2] ), .IN1(
        \ab[220][3] ), .COUT(\CARRYB[221][2] ), .SUM(\SUMB[221][2] ) );
  FADDER S1_220_0 ( .CIN(\ab[220][0] ), .IN0(\CARRYB[219][0] ), .IN1(
        \SUMB[219][1] ), .COUT(\CARRYB[220][0] ), .SUM(PRODUCT[220]) );
  FADDER S2_220_1 ( .CIN(\ab[220][1] ), .IN0(\CARRYB[219][1] ), .IN1(
        \SUMB[219][2] ), .COUT(\CARRYB[220][1] ), .SUM(\SUMB[220][1] ) );
  FADDER S3_220_2 ( .CIN(\ab[220][2] ), .IN0(\CARRYB[219][2] ), .IN1(
        \ab[219][3] ), .COUT(\CARRYB[220][2] ), .SUM(\SUMB[220][2] ) );
  FADDER S1_219_0 ( .CIN(\ab[219][0] ), .IN0(\CARRYB[218][0] ), .IN1(
        \SUMB[218][1] ), .COUT(\CARRYB[219][0] ), .SUM(PRODUCT[219]) );
  FADDER S2_219_1 ( .CIN(\ab[219][1] ), .IN0(\CARRYB[218][1] ), .IN1(
        \SUMB[218][2] ), .COUT(\CARRYB[219][1] ), .SUM(\SUMB[219][1] ) );
  FADDER S3_219_2 ( .CIN(\ab[219][2] ), .IN0(\CARRYB[218][2] ), .IN1(
        \ab[218][3] ), .COUT(\CARRYB[219][2] ), .SUM(\SUMB[219][2] ) );
  FADDER S1_218_0 ( .CIN(\ab[218][0] ), .IN0(\CARRYB[217][0] ), .IN1(
        \SUMB[217][1] ), .COUT(\CARRYB[218][0] ), .SUM(PRODUCT[218]) );
  FADDER S2_218_1 ( .CIN(\ab[218][1] ), .IN0(\CARRYB[217][1] ), .IN1(
        \SUMB[217][2] ), .COUT(\CARRYB[218][1] ), .SUM(\SUMB[218][1] ) );
  FADDER S3_218_2 ( .CIN(\ab[218][2] ), .IN0(\CARRYB[217][2] ), .IN1(
        \ab[217][3] ), .COUT(\CARRYB[218][2] ), .SUM(\SUMB[218][2] ) );
  FADDER S1_217_0 ( .CIN(\ab[217][0] ), .IN0(\CARRYB[216][0] ), .IN1(
        \SUMB[216][1] ), .COUT(\CARRYB[217][0] ), .SUM(PRODUCT[217]) );
  FADDER S2_217_1 ( .CIN(\ab[217][1] ), .IN0(\CARRYB[216][1] ), .IN1(
        \SUMB[216][2] ), .COUT(\CARRYB[217][1] ), .SUM(\SUMB[217][1] ) );
  FADDER S3_217_2 ( .CIN(\ab[217][2] ), .IN0(\CARRYB[216][2] ), .IN1(
        \ab[216][3] ), .COUT(\CARRYB[217][2] ), .SUM(\SUMB[217][2] ) );
  FADDER S1_216_0 ( .CIN(\ab[216][0] ), .IN0(\CARRYB[215][0] ), .IN1(
        \SUMB[215][1] ), .COUT(\CARRYB[216][0] ), .SUM(PRODUCT[216]) );
  FADDER S2_216_1 ( .CIN(\ab[216][1] ), .IN0(\CARRYB[215][1] ), .IN1(
        \SUMB[215][2] ), .COUT(\CARRYB[216][1] ), .SUM(\SUMB[216][1] ) );
  FADDER S3_216_2 ( .CIN(\ab[216][2] ), .IN0(\CARRYB[215][2] ), .IN1(
        \ab[215][3] ), .COUT(\CARRYB[216][2] ), .SUM(\SUMB[216][2] ) );
  FADDER S1_215_0 ( .CIN(\ab[215][0] ), .IN0(\CARRYB[214][0] ), .IN1(
        \SUMB[214][1] ), .COUT(\CARRYB[215][0] ), .SUM(PRODUCT[215]) );
  FADDER S2_215_1 ( .CIN(\ab[215][1] ), .IN0(\CARRYB[214][1] ), .IN1(
        \SUMB[214][2] ), .COUT(\CARRYB[215][1] ), .SUM(\SUMB[215][1] ) );
  FADDER S3_215_2 ( .CIN(\ab[215][2] ), .IN0(\CARRYB[214][2] ), .IN1(
        \ab[214][3] ), .COUT(\CARRYB[215][2] ), .SUM(\SUMB[215][2] ) );
  FADDER S1_214_0 ( .CIN(\ab[214][0] ), .IN0(\CARRYB[213][0] ), .IN1(
        \SUMB[213][1] ), .COUT(\CARRYB[214][0] ), .SUM(PRODUCT[214]) );
  FADDER S2_214_1 ( .CIN(\ab[214][1] ), .IN0(\CARRYB[213][1] ), .IN1(
        \SUMB[213][2] ), .COUT(\CARRYB[214][1] ), .SUM(\SUMB[214][1] ) );
  FADDER S3_214_2 ( .CIN(\ab[214][2] ), .IN0(\CARRYB[213][2] ), .IN1(
        \ab[213][3] ), .COUT(\CARRYB[214][2] ), .SUM(\SUMB[214][2] ) );
  FADDER S1_213_0 ( .CIN(\ab[213][0] ), .IN0(\CARRYB[212][0] ), .IN1(
        \SUMB[212][1] ), .COUT(\CARRYB[213][0] ), .SUM(PRODUCT[213]) );
  FADDER S2_213_1 ( .CIN(\ab[213][1] ), .IN0(\CARRYB[212][1] ), .IN1(
        \SUMB[212][2] ), .COUT(\CARRYB[213][1] ), .SUM(\SUMB[213][1] ) );
  FADDER S3_213_2 ( .CIN(\ab[213][2] ), .IN0(\CARRYB[212][2] ), .IN1(
        \ab[212][3] ), .COUT(\CARRYB[213][2] ), .SUM(\SUMB[213][2] ) );
  FADDER S1_212_0 ( .CIN(\ab[212][0] ), .IN0(\CARRYB[211][0] ), .IN1(
        \SUMB[211][1] ), .COUT(\CARRYB[212][0] ), .SUM(PRODUCT[212]) );
  FADDER S2_212_1 ( .CIN(\ab[212][1] ), .IN0(\CARRYB[211][1] ), .IN1(
        \SUMB[211][2] ), .COUT(\CARRYB[212][1] ), .SUM(\SUMB[212][1] ) );
  FADDER S3_212_2 ( .CIN(\ab[212][2] ), .IN0(\CARRYB[211][2] ), .IN1(
        \ab[211][3] ), .COUT(\CARRYB[212][2] ), .SUM(\SUMB[212][2] ) );
  FADDER S1_211_0 ( .CIN(\ab[211][0] ), .IN0(\CARRYB[210][0] ), .IN1(
        \SUMB[210][1] ), .COUT(\CARRYB[211][0] ), .SUM(PRODUCT[211]) );
  FADDER S2_211_1 ( .CIN(\ab[211][1] ), .IN0(\CARRYB[210][1] ), .IN1(
        \SUMB[210][2] ), .COUT(\CARRYB[211][1] ), .SUM(\SUMB[211][1] ) );
  FADDER S3_211_2 ( .CIN(\ab[211][2] ), .IN0(\CARRYB[210][2] ), .IN1(
        \ab[210][3] ), .COUT(\CARRYB[211][2] ), .SUM(\SUMB[211][2] ) );
  FADDER S1_210_0 ( .CIN(\ab[210][0] ), .IN0(\CARRYB[209][0] ), .IN1(
        \SUMB[209][1] ), .COUT(\CARRYB[210][0] ), .SUM(PRODUCT[210]) );
  FADDER S2_210_1 ( .CIN(\ab[210][1] ), .IN0(\CARRYB[209][1] ), .IN1(
        \SUMB[209][2] ), .COUT(\CARRYB[210][1] ), .SUM(\SUMB[210][1] ) );
  FADDER S3_210_2 ( .CIN(\ab[210][2] ), .IN0(\CARRYB[209][2] ), .IN1(
        \ab[209][3] ), .COUT(\CARRYB[210][2] ), .SUM(\SUMB[210][2] ) );
  FADDER S1_209_0 ( .CIN(\ab[209][0] ), .IN0(\CARRYB[208][0] ), .IN1(
        \SUMB[208][1] ), .COUT(\CARRYB[209][0] ), .SUM(PRODUCT[209]) );
  FADDER S2_209_1 ( .CIN(\ab[209][1] ), .IN0(\CARRYB[208][1] ), .IN1(
        \SUMB[208][2] ), .COUT(\CARRYB[209][1] ), .SUM(\SUMB[209][1] ) );
  FADDER S3_209_2 ( .CIN(\ab[209][2] ), .IN0(\CARRYB[208][2] ), .IN1(
        \ab[208][3] ), .COUT(\CARRYB[209][2] ), .SUM(\SUMB[209][2] ) );
  FADDER S1_208_0 ( .CIN(\ab[208][0] ), .IN0(\CARRYB[207][0] ), .IN1(
        \SUMB[207][1] ), .COUT(\CARRYB[208][0] ), .SUM(PRODUCT[208]) );
  FADDER S2_208_1 ( .CIN(\ab[208][1] ), .IN0(\CARRYB[207][1] ), .IN1(
        \SUMB[207][2] ), .COUT(\CARRYB[208][1] ), .SUM(\SUMB[208][1] ) );
  FADDER S3_208_2 ( .CIN(\ab[208][2] ), .IN0(\CARRYB[207][2] ), .IN1(
        \ab[207][3] ), .COUT(\CARRYB[208][2] ), .SUM(\SUMB[208][2] ) );
  FADDER S1_207_0 ( .CIN(\ab[207][0] ), .IN0(\CARRYB[206][0] ), .IN1(
        \SUMB[206][1] ), .COUT(\CARRYB[207][0] ), .SUM(PRODUCT[207]) );
  FADDER S2_207_1 ( .CIN(\ab[207][1] ), .IN0(\CARRYB[206][1] ), .IN1(
        \SUMB[206][2] ), .COUT(\CARRYB[207][1] ), .SUM(\SUMB[207][1] ) );
  FADDER S3_207_2 ( .CIN(\ab[207][2] ), .IN0(\CARRYB[206][2] ), .IN1(
        \ab[206][3] ), .COUT(\CARRYB[207][2] ), .SUM(\SUMB[207][2] ) );
  FADDER S1_206_0 ( .CIN(\ab[206][0] ), .IN0(\CARRYB[205][0] ), .IN1(
        \SUMB[205][1] ), .COUT(\CARRYB[206][0] ), .SUM(PRODUCT[206]) );
  FADDER S2_206_1 ( .CIN(\ab[206][1] ), .IN0(\CARRYB[205][1] ), .IN1(
        \SUMB[205][2] ), .COUT(\CARRYB[206][1] ), .SUM(\SUMB[206][1] ) );
  FADDER S3_206_2 ( .CIN(\ab[206][2] ), .IN0(\CARRYB[205][2] ), .IN1(
        \ab[205][3] ), .COUT(\CARRYB[206][2] ), .SUM(\SUMB[206][2] ) );
  FADDER S1_205_0 ( .CIN(\ab[205][0] ), .IN0(\CARRYB[204][0] ), .IN1(
        \SUMB[204][1] ), .COUT(\CARRYB[205][0] ), .SUM(PRODUCT[205]) );
  FADDER S2_205_1 ( .CIN(\ab[205][1] ), .IN0(\CARRYB[204][1] ), .IN1(
        \SUMB[204][2] ), .COUT(\CARRYB[205][1] ), .SUM(\SUMB[205][1] ) );
  FADDER S3_205_2 ( .CIN(\ab[205][2] ), .IN0(\CARRYB[204][2] ), .IN1(
        \ab[204][3] ), .COUT(\CARRYB[205][2] ), .SUM(\SUMB[205][2] ) );
  FADDER S1_204_0 ( .CIN(\ab[204][0] ), .IN0(\CARRYB[203][0] ), .IN1(
        \SUMB[203][1] ), .COUT(\CARRYB[204][0] ), .SUM(PRODUCT[204]) );
  FADDER S2_204_1 ( .CIN(\ab[204][1] ), .IN0(\CARRYB[203][1] ), .IN1(
        \SUMB[203][2] ), .COUT(\CARRYB[204][1] ), .SUM(\SUMB[204][1] ) );
  FADDER S3_204_2 ( .CIN(\ab[204][2] ), .IN0(\CARRYB[203][2] ), .IN1(
        \ab[203][3] ), .COUT(\CARRYB[204][2] ), .SUM(\SUMB[204][2] ) );
  FADDER S1_203_0 ( .CIN(\ab[203][0] ), .IN0(\CARRYB[202][0] ), .IN1(
        \SUMB[202][1] ), .COUT(\CARRYB[203][0] ), .SUM(PRODUCT[203]) );
  FADDER S2_203_1 ( .CIN(\ab[203][1] ), .IN0(\CARRYB[202][1] ), .IN1(
        \SUMB[202][2] ), .COUT(\CARRYB[203][1] ), .SUM(\SUMB[203][1] ) );
  FADDER S3_203_2 ( .CIN(\ab[203][2] ), .IN0(\CARRYB[202][2] ), .IN1(
        \ab[202][3] ), .COUT(\CARRYB[203][2] ), .SUM(\SUMB[203][2] ) );
  FADDER S1_202_0 ( .CIN(\ab[202][0] ), .IN0(\CARRYB[201][0] ), .IN1(
        \SUMB[201][1] ), .COUT(\CARRYB[202][0] ), .SUM(PRODUCT[202]) );
  FADDER S2_202_1 ( .CIN(\ab[202][1] ), .IN0(\CARRYB[201][1] ), .IN1(
        \SUMB[201][2] ), .COUT(\CARRYB[202][1] ), .SUM(\SUMB[202][1] ) );
  FADDER S3_202_2 ( .CIN(\ab[202][2] ), .IN0(\CARRYB[201][2] ), .IN1(
        \ab[201][3] ), .COUT(\CARRYB[202][2] ), .SUM(\SUMB[202][2] ) );
  FADDER S1_201_0 ( .CIN(\ab[201][0] ), .IN0(\CARRYB[200][0] ), .IN1(
        \SUMB[200][1] ), .COUT(\CARRYB[201][0] ), .SUM(PRODUCT[201]) );
  FADDER S2_201_1 ( .CIN(\ab[201][1] ), .IN0(\CARRYB[200][1] ), .IN1(
        \SUMB[200][2] ), .COUT(\CARRYB[201][1] ), .SUM(\SUMB[201][1] ) );
  FADDER S3_201_2 ( .CIN(\ab[201][2] ), .IN0(\CARRYB[200][2] ), .IN1(
        \ab[200][3] ), .COUT(\CARRYB[201][2] ), .SUM(\SUMB[201][2] ) );
  FADDER S1_200_0 ( .CIN(\ab[200][0] ), .IN0(\CARRYB[199][0] ), .IN1(
        \SUMB[199][1] ), .COUT(\CARRYB[200][0] ), .SUM(PRODUCT[200]) );
  FADDER S2_200_1 ( .CIN(\ab[200][1] ), .IN0(\CARRYB[199][1] ), .IN1(
        \SUMB[199][2] ), .COUT(\CARRYB[200][1] ), .SUM(\SUMB[200][1] ) );
  FADDER S3_200_2 ( .CIN(\ab[200][2] ), .IN0(\CARRYB[199][2] ), .IN1(
        \ab[199][3] ), .COUT(\CARRYB[200][2] ), .SUM(\SUMB[200][2] ) );
  FADDER S1_199_0 ( .CIN(\ab[199][0] ), .IN0(\CARRYB[198][0] ), .IN1(
        \SUMB[198][1] ), .COUT(\CARRYB[199][0] ), .SUM(PRODUCT[199]) );
  FADDER S2_199_1 ( .CIN(\ab[199][1] ), .IN0(\CARRYB[198][1] ), .IN1(
        \SUMB[198][2] ), .COUT(\CARRYB[199][1] ), .SUM(\SUMB[199][1] ) );
  FADDER S3_199_2 ( .CIN(\ab[199][2] ), .IN0(\CARRYB[198][2] ), .IN1(
        \ab[198][3] ), .COUT(\CARRYB[199][2] ), .SUM(\SUMB[199][2] ) );
  FADDER S1_198_0 ( .CIN(\ab[198][0] ), .IN0(\CARRYB[197][0] ), .IN1(
        \SUMB[197][1] ), .COUT(\CARRYB[198][0] ), .SUM(PRODUCT[198]) );
  FADDER S2_198_1 ( .CIN(\ab[198][1] ), .IN0(\CARRYB[197][1] ), .IN1(
        \SUMB[197][2] ), .COUT(\CARRYB[198][1] ), .SUM(\SUMB[198][1] ) );
  FADDER S3_198_2 ( .CIN(\ab[198][2] ), .IN0(\CARRYB[197][2] ), .IN1(
        \ab[197][3] ), .COUT(\CARRYB[198][2] ), .SUM(\SUMB[198][2] ) );
  FADDER S1_197_0 ( .CIN(\ab[197][0] ), .IN0(\CARRYB[196][0] ), .IN1(
        \SUMB[196][1] ), .COUT(\CARRYB[197][0] ), .SUM(PRODUCT[197]) );
  FADDER S2_197_1 ( .CIN(\ab[197][1] ), .IN0(\CARRYB[196][1] ), .IN1(
        \SUMB[196][2] ), .COUT(\CARRYB[197][1] ), .SUM(\SUMB[197][1] ) );
  FADDER S3_197_2 ( .CIN(\ab[197][2] ), .IN0(\CARRYB[196][2] ), .IN1(
        \ab[196][3] ), .COUT(\CARRYB[197][2] ), .SUM(\SUMB[197][2] ) );
  FADDER S1_196_0 ( .CIN(\ab[196][0] ), .IN0(\CARRYB[195][0] ), .IN1(
        \SUMB[195][1] ), .COUT(\CARRYB[196][0] ), .SUM(PRODUCT[196]) );
  FADDER S2_196_1 ( .CIN(\ab[196][1] ), .IN0(\CARRYB[195][1] ), .IN1(
        \SUMB[195][2] ), .COUT(\CARRYB[196][1] ), .SUM(\SUMB[196][1] ) );
  FADDER S3_196_2 ( .CIN(\ab[196][2] ), .IN0(\CARRYB[195][2] ), .IN1(
        \ab[195][3] ), .COUT(\CARRYB[196][2] ), .SUM(\SUMB[196][2] ) );
  FADDER S1_195_0 ( .CIN(\ab[195][0] ), .IN0(\CARRYB[194][0] ), .IN1(
        \SUMB[194][1] ), .COUT(\CARRYB[195][0] ), .SUM(PRODUCT[195]) );
  FADDER S2_195_1 ( .CIN(\ab[195][1] ), .IN0(\CARRYB[194][1] ), .IN1(
        \SUMB[194][2] ), .COUT(\CARRYB[195][1] ), .SUM(\SUMB[195][1] ) );
  FADDER S3_195_2 ( .CIN(\ab[195][2] ), .IN0(\CARRYB[194][2] ), .IN1(
        \ab[194][3] ), .COUT(\CARRYB[195][2] ), .SUM(\SUMB[195][2] ) );
  FADDER S1_194_0 ( .CIN(\ab[194][0] ), .IN0(\CARRYB[193][0] ), .IN1(
        \SUMB[193][1] ), .COUT(\CARRYB[194][0] ), .SUM(PRODUCT[194]) );
  FADDER S2_194_1 ( .CIN(\ab[194][1] ), .IN0(\CARRYB[193][1] ), .IN1(
        \SUMB[193][2] ), .COUT(\CARRYB[194][1] ), .SUM(\SUMB[194][1] ) );
  FADDER S3_194_2 ( .CIN(\ab[194][2] ), .IN0(\CARRYB[193][2] ), .IN1(
        \ab[193][3] ), .COUT(\CARRYB[194][2] ), .SUM(\SUMB[194][2] ) );
  FADDER S1_193_0 ( .CIN(\ab[193][0] ), .IN0(\CARRYB[192][0] ), .IN1(
        \SUMB[192][1] ), .COUT(\CARRYB[193][0] ), .SUM(PRODUCT[193]) );
  FADDER S2_193_1 ( .CIN(\ab[193][1] ), .IN0(\CARRYB[192][1] ), .IN1(
        \SUMB[192][2] ), .COUT(\CARRYB[193][1] ), .SUM(\SUMB[193][1] ) );
  FADDER S3_193_2 ( .CIN(\ab[193][2] ), .IN0(\CARRYB[192][2] ), .IN1(
        \ab[192][3] ), .COUT(\CARRYB[193][2] ), .SUM(\SUMB[193][2] ) );
  FADDER S1_192_0 ( .CIN(\ab[192][0] ), .IN0(\CARRYB[191][0] ), .IN1(
        \SUMB[191][1] ), .COUT(\CARRYB[192][0] ), .SUM(PRODUCT[192]) );
  FADDER S2_192_1 ( .CIN(\ab[192][1] ), .IN0(\CARRYB[191][1] ), .IN1(
        \SUMB[191][2] ), .COUT(\CARRYB[192][1] ), .SUM(\SUMB[192][1] ) );
  FADDER S3_192_2 ( .CIN(\ab[192][2] ), .IN0(\CARRYB[191][2] ), .IN1(
        \ab[191][3] ), .COUT(\CARRYB[192][2] ), .SUM(\SUMB[192][2] ) );
  FADDER S1_191_0 ( .CIN(\ab[191][0] ), .IN0(\CARRYB[190][0] ), .IN1(
        \SUMB[190][1] ), .COUT(\CARRYB[191][0] ), .SUM(PRODUCT[191]) );
  FADDER S2_191_1 ( .CIN(\ab[191][1] ), .IN0(\CARRYB[190][1] ), .IN1(
        \SUMB[190][2] ), .COUT(\CARRYB[191][1] ), .SUM(\SUMB[191][1] ) );
  FADDER S3_191_2 ( .CIN(\ab[191][2] ), .IN0(\CARRYB[190][2] ), .IN1(
        \ab[190][3] ), .COUT(\CARRYB[191][2] ), .SUM(\SUMB[191][2] ) );
  FADDER S1_190_0 ( .CIN(\ab[190][0] ), .IN0(\CARRYB[189][0] ), .IN1(
        \SUMB[189][1] ), .COUT(\CARRYB[190][0] ), .SUM(PRODUCT[190]) );
  FADDER S2_190_1 ( .CIN(\ab[190][1] ), .IN0(\CARRYB[189][1] ), .IN1(
        \SUMB[189][2] ), .COUT(\CARRYB[190][1] ), .SUM(\SUMB[190][1] ) );
  FADDER S3_190_2 ( .CIN(\ab[190][2] ), .IN0(\CARRYB[189][2] ), .IN1(
        \ab[189][3] ), .COUT(\CARRYB[190][2] ), .SUM(\SUMB[190][2] ) );
  FADDER S1_189_0 ( .CIN(\ab[189][0] ), .IN0(\CARRYB[188][0] ), .IN1(
        \SUMB[188][1] ), .COUT(\CARRYB[189][0] ), .SUM(PRODUCT[189]) );
  FADDER S2_189_1 ( .CIN(\ab[189][1] ), .IN0(\CARRYB[188][1] ), .IN1(
        \SUMB[188][2] ), .COUT(\CARRYB[189][1] ), .SUM(\SUMB[189][1] ) );
  FADDER S3_189_2 ( .CIN(\ab[189][2] ), .IN0(\CARRYB[188][2] ), .IN1(
        \ab[188][3] ), .COUT(\CARRYB[189][2] ), .SUM(\SUMB[189][2] ) );
  FADDER S1_188_0 ( .CIN(\ab[188][0] ), .IN0(\CARRYB[187][0] ), .IN1(
        \SUMB[187][1] ), .COUT(\CARRYB[188][0] ), .SUM(PRODUCT[188]) );
  FADDER S2_188_1 ( .CIN(\ab[188][1] ), .IN0(\CARRYB[187][1] ), .IN1(
        \SUMB[187][2] ), .COUT(\CARRYB[188][1] ), .SUM(\SUMB[188][1] ) );
  FADDER S3_188_2 ( .CIN(\ab[188][2] ), .IN0(\CARRYB[187][2] ), .IN1(
        \ab[187][3] ), .COUT(\CARRYB[188][2] ), .SUM(\SUMB[188][2] ) );
  FADDER S1_187_0 ( .CIN(\ab[187][0] ), .IN0(\CARRYB[186][0] ), .IN1(
        \SUMB[186][1] ), .COUT(\CARRYB[187][0] ), .SUM(PRODUCT[187]) );
  FADDER S2_187_1 ( .CIN(\ab[187][1] ), .IN0(\CARRYB[186][1] ), .IN1(
        \SUMB[186][2] ), .COUT(\CARRYB[187][1] ), .SUM(\SUMB[187][1] ) );
  FADDER S3_187_2 ( .CIN(\ab[187][2] ), .IN0(\CARRYB[186][2] ), .IN1(
        \ab[186][3] ), .COUT(\CARRYB[187][2] ), .SUM(\SUMB[187][2] ) );
  FADDER S1_186_0 ( .CIN(\ab[186][0] ), .IN0(\CARRYB[185][0] ), .IN1(
        \SUMB[185][1] ), .COUT(\CARRYB[186][0] ), .SUM(PRODUCT[186]) );
  FADDER S2_186_1 ( .CIN(\ab[186][1] ), .IN0(\CARRYB[185][1] ), .IN1(
        \SUMB[185][2] ), .COUT(\CARRYB[186][1] ), .SUM(\SUMB[186][1] ) );
  FADDER S3_186_2 ( .CIN(\ab[186][2] ), .IN0(\CARRYB[185][2] ), .IN1(
        \ab[185][3] ), .COUT(\CARRYB[186][2] ), .SUM(\SUMB[186][2] ) );
  FADDER S1_185_0 ( .CIN(\ab[185][0] ), .IN0(\CARRYB[184][0] ), .IN1(
        \SUMB[184][1] ), .COUT(\CARRYB[185][0] ), .SUM(PRODUCT[185]) );
  FADDER S2_185_1 ( .CIN(\ab[185][1] ), .IN0(\CARRYB[184][1] ), .IN1(
        \SUMB[184][2] ), .COUT(\CARRYB[185][1] ), .SUM(\SUMB[185][1] ) );
  FADDER S3_185_2 ( .CIN(\ab[185][2] ), .IN0(\CARRYB[184][2] ), .IN1(
        \ab[184][3] ), .COUT(\CARRYB[185][2] ), .SUM(\SUMB[185][2] ) );
  FADDER S1_184_0 ( .CIN(\ab[184][0] ), .IN0(\CARRYB[183][0] ), .IN1(
        \SUMB[183][1] ), .COUT(\CARRYB[184][0] ), .SUM(PRODUCT[184]) );
  FADDER S2_184_1 ( .CIN(\ab[184][1] ), .IN0(\CARRYB[183][1] ), .IN1(
        \SUMB[183][2] ), .COUT(\CARRYB[184][1] ), .SUM(\SUMB[184][1] ) );
  FADDER S3_184_2 ( .CIN(\ab[184][2] ), .IN0(\CARRYB[183][2] ), .IN1(
        \ab[183][3] ), .COUT(\CARRYB[184][2] ), .SUM(\SUMB[184][2] ) );
  FADDER S1_183_0 ( .CIN(\ab[183][0] ), .IN0(\CARRYB[182][0] ), .IN1(
        \SUMB[182][1] ), .COUT(\CARRYB[183][0] ), .SUM(PRODUCT[183]) );
  FADDER S2_183_1 ( .CIN(\ab[183][1] ), .IN0(\CARRYB[182][1] ), .IN1(
        \SUMB[182][2] ), .COUT(\CARRYB[183][1] ), .SUM(\SUMB[183][1] ) );
  FADDER S3_183_2 ( .CIN(\ab[183][2] ), .IN0(\CARRYB[182][2] ), .IN1(
        \ab[182][3] ), .COUT(\CARRYB[183][2] ), .SUM(\SUMB[183][2] ) );
  FADDER S1_182_0 ( .CIN(\ab[182][0] ), .IN0(\CARRYB[181][0] ), .IN1(
        \SUMB[181][1] ), .COUT(\CARRYB[182][0] ), .SUM(PRODUCT[182]) );
  FADDER S2_182_1 ( .CIN(\ab[182][1] ), .IN0(\CARRYB[181][1] ), .IN1(
        \SUMB[181][2] ), .COUT(\CARRYB[182][1] ), .SUM(\SUMB[182][1] ) );
  FADDER S3_182_2 ( .CIN(\ab[182][2] ), .IN0(\CARRYB[181][2] ), .IN1(
        \ab[181][3] ), .COUT(\CARRYB[182][2] ), .SUM(\SUMB[182][2] ) );
  FADDER S1_181_0 ( .CIN(\ab[181][0] ), .IN0(\CARRYB[180][0] ), .IN1(
        \SUMB[180][1] ), .COUT(\CARRYB[181][0] ), .SUM(PRODUCT[181]) );
  FADDER S2_181_1 ( .CIN(\ab[181][1] ), .IN0(\CARRYB[180][1] ), .IN1(
        \SUMB[180][2] ), .COUT(\CARRYB[181][1] ), .SUM(\SUMB[181][1] ) );
  FADDER S3_181_2 ( .CIN(\ab[181][2] ), .IN0(\CARRYB[180][2] ), .IN1(
        \ab[180][3] ), .COUT(\CARRYB[181][2] ), .SUM(\SUMB[181][2] ) );
  FADDER S1_180_0 ( .CIN(\ab[180][0] ), .IN0(\CARRYB[179][0] ), .IN1(
        \SUMB[179][1] ), .COUT(\CARRYB[180][0] ), .SUM(PRODUCT[180]) );
  FADDER S2_180_1 ( .CIN(\ab[180][1] ), .IN0(\CARRYB[179][1] ), .IN1(
        \SUMB[179][2] ), .COUT(\CARRYB[180][1] ), .SUM(\SUMB[180][1] ) );
  FADDER S3_180_2 ( .CIN(\ab[180][2] ), .IN0(\CARRYB[179][2] ), .IN1(
        \ab[179][3] ), .COUT(\CARRYB[180][2] ), .SUM(\SUMB[180][2] ) );
  FADDER S1_179_0 ( .CIN(\ab[179][0] ), .IN0(\CARRYB[178][0] ), .IN1(
        \SUMB[178][1] ), .COUT(\CARRYB[179][0] ), .SUM(PRODUCT[179]) );
  FADDER S2_179_1 ( .CIN(\ab[179][1] ), .IN0(\CARRYB[178][1] ), .IN1(
        \SUMB[178][2] ), .COUT(\CARRYB[179][1] ), .SUM(\SUMB[179][1] ) );
  FADDER S3_179_2 ( .CIN(\ab[179][2] ), .IN0(\CARRYB[178][2] ), .IN1(
        \ab[178][3] ), .COUT(\CARRYB[179][2] ), .SUM(\SUMB[179][2] ) );
  FADDER S1_178_0 ( .CIN(\ab[178][0] ), .IN0(\CARRYB[177][0] ), .IN1(
        \SUMB[177][1] ), .COUT(\CARRYB[178][0] ), .SUM(PRODUCT[178]) );
  FADDER S2_178_1 ( .CIN(\ab[178][1] ), .IN0(\CARRYB[177][1] ), .IN1(
        \SUMB[177][2] ), .COUT(\CARRYB[178][1] ), .SUM(\SUMB[178][1] ) );
  FADDER S3_178_2 ( .CIN(\ab[178][2] ), .IN0(\CARRYB[177][2] ), .IN1(
        \ab[177][3] ), .COUT(\CARRYB[178][2] ), .SUM(\SUMB[178][2] ) );
  FADDER S1_177_0 ( .CIN(\ab[177][0] ), .IN0(\CARRYB[176][0] ), .IN1(
        \SUMB[176][1] ), .COUT(\CARRYB[177][0] ), .SUM(PRODUCT[177]) );
  FADDER S2_177_1 ( .CIN(\ab[177][1] ), .IN0(\CARRYB[176][1] ), .IN1(
        \SUMB[176][2] ), .COUT(\CARRYB[177][1] ), .SUM(\SUMB[177][1] ) );
  FADDER S3_177_2 ( .CIN(\ab[177][2] ), .IN0(\CARRYB[176][2] ), .IN1(
        \ab[176][3] ), .COUT(\CARRYB[177][2] ), .SUM(\SUMB[177][2] ) );
  FADDER S1_176_0 ( .CIN(\ab[176][0] ), .IN0(\CARRYB[175][0] ), .IN1(
        \SUMB[175][1] ), .COUT(\CARRYB[176][0] ), .SUM(PRODUCT[176]) );
  FADDER S2_176_1 ( .CIN(\ab[176][1] ), .IN0(\CARRYB[175][1] ), .IN1(
        \SUMB[175][2] ), .COUT(\CARRYB[176][1] ), .SUM(\SUMB[176][1] ) );
  FADDER S3_176_2 ( .CIN(\ab[176][2] ), .IN0(\CARRYB[175][2] ), .IN1(
        \ab[175][3] ), .COUT(\CARRYB[176][2] ), .SUM(\SUMB[176][2] ) );
  FADDER S1_175_0 ( .CIN(\ab[175][0] ), .IN0(\CARRYB[174][0] ), .IN1(
        \SUMB[174][1] ), .COUT(\CARRYB[175][0] ), .SUM(PRODUCT[175]) );
  FADDER S2_175_1 ( .CIN(\ab[175][1] ), .IN0(\CARRYB[174][1] ), .IN1(
        \SUMB[174][2] ), .COUT(\CARRYB[175][1] ), .SUM(\SUMB[175][1] ) );
  FADDER S3_175_2 ( .CIN(\ab[175][2] ), .IN0(\CARRYB[174][2] ), .IN1(
        \ab[174][3] ), .COUT(\CARRYB[175][2] ), .SUM(\SUMB[175][2] ) );
  FADDER S1_174_0 ( .CIN(\ab[174][0] ), .IN0(\CARRYB[173][0] ), .IN1(
        \SUMB[173][1] ), .COUT(\CARRYB[174][0] ), .SUM(PRODUCT[174]) );
  FADDER S2_174_1 ( .CIN(\ab[174][1] ), .IN0(\CARRYB[173][1] ), .IN1(
        \SUMB[173][2] ), .COUT(\CARRYB[174][1] ), .SUM(\SUMB[174][1] ) );
  FADDER S3_174_2 ( .CIN(\ab[174][2] ), .IN0(\CARRYB[173][2] ), .IN1(
        \ab[173][3] ), .COUT(\CARRYB[174][2] ), .SUM(\SUMB[174][2] ) );
  FADDER S1_173_0 ( .CIN(\ab[173][0] ), .IN0(\CARRYB[172][0] ), .IN1(
        \SUMB[172][1] ), .COUT(\CARRYB[173][0] ), .SUM(PRODUCT[173]) );
  FADDER S2_173_1 ( .CIN(\ab[173][1] ), .IN0(\CARRYB[172][1] ), .IN1(
        \SUMB[172][2] ), .COUT(\CARRYB[173][1] ), .SUM(\SUMB[173][1] ) );
  FADDER S3_173_2 ( .CIN(\ab[173][2] ), .IN0(\CARRYB[172][2] ), .IN1(
        \ab[172][3] ), .COUT(\CARRYB[173][2] ), .SUM(\SUMB[173][2] ) );
  FADDER S1_172_0 ( .CIN(\ab[172][0] ), .IN0(\CARRYB[171][0] ), .IN1(
        \SUMB[171][1] ), .COUT(\CARRYB[172][0] ), .SUM(PRODUCT[172]) );
  FADDER S2_172_1 ( .CIN(\ab[172][1] ), .IN0(\CARRYB[171][1] ), .IN1(
        \SUMB[171][2] ), .COUT(\CARRYB[172][1] ), .SUM(\SUMB[172][1] ) );
  FADDER S3_172_2 ( .CIN(\ab[172][2] ), .IN0(\CARRYB[171][2] ), .IN1(
        \ab[171][3] ), .COUT(\CARRYB[172][2] ), .SUM(\SUMB[172][2] ) );
  FADDER S1_171_0 ( .CIN(\ab[171][0] ), .IN0(\CARRYB[170][0] ), .IN1(
        \SUMB[170][1] ), .COUT(\CARRYB[171][0] ), .SUM(PRODUCT[171]) );
  FADDER S2_171_1 ( .CIN(\ab[171][1] ), .IN0(\CARRYB[170][1] ), .IN1(
        \SUMB[170][2] ), .COUT(\CARRYB[171][1] ), .SUM(\SUMB[171][1] ) );
  FADDER S3_171_2 ( .CIN(\ab[171][2] ), .IN0(\CARRYB[170][2] ), .IN1(
        \ab[170][3] ), .COUT(\CARRYB[171][2] ), .SUM(\SUMB[171][2] ) );
  FADDER S1_170_0 ( .CIN(\ab[170][0] ), .IN0(\CARRYB[169][0] ), .IN1(
        \SUMB[169][1] ), .COUT(\CARRYB[170][0] ), .SUM(PRODUCT[170]) );
  FADDER S2_170_1 ( .CIN(\ab[170][1] ), .IN0(\CARRYB[169][1] ), .IN1(
        \SUMB[169][2] ), .COUT(\CARRYB[170][1] ), .SUM(\SUMB[170][1] ) );
  FADDER S3_170_2 ( .CIN(\ab[170][2] ), .IN0(\CARRYB[169][2] ), .IN1(
        \ab[169][3] ), .COUT(\CARRYB[170][2] ), .SUM(\SUMB[170][2] ) );
  FADDER S1_169_0 ( .CIN(\ab[169][0] ), .IN0(\CARRYB[168][0] ), .IN1(
        \SUMB[168][1] ), .COUT(\CARRYB[169][0] ), .SUM(PRODUCT[169]) );
  FADDER S2_169_1 ( .CIN(\ab[169][1] ), .IN0(\CARRYB[168][1] ), .IN1(
        \SUMB[168][2] ), .COUT(\CARRYB[169][1] ), .SUM(\SUMB[169][1] ) );
  FADDER S3_169_2 ( .CIN(\ab[169][2] ), .IN0(\CARRYB[168][2] ), .IN1(
        \ab[168][3] ), .COUT(\CARRYB[169][2] ), .SUM(\SUMB[169][2] ) );
  FADDER S1_168_0 ( .CIN(\ab[168][0] ), .IN0(\CARRYB[167][0] ), .IN1(
        \SUMB[167][1] ), .COUT(\CARRYB[168][0] ), .SUM(PRODUCT[168]) );
  FADDER S2_168_1 ( .CIN(\ab[168][1] ), .IN0(\CARRYB[167][1] ), .IN1(
        \SUMB[167][2] ), .COUT(\CARRYB[168][1] ), .SUM(\SUMB[168][1] ) );
  FADDER S3_168_2 ( .CIN(\ab[168][2] ), .IN0(\CARRYB[167][2] ), .IN1(
        \ab[167][3] ), .COUT(\CARRYB[168][2] ), .SUM(\SUMB[168][2] ) );
  FADDER S1_167_0 ( .CIN(\ab[167][0] ), .IN0(\CARRYB[166][0] ), .IN1(
        \SUMB[166][1] ), .COUT(\CARRYB[167][0] ), .SUM(PRODUCT[167]) );
  FADDER S2_167_1 ( .CIN(\ab[167][1] ), .IN0(\CARRYB[166][1] ), .IN1(
        \SUMB[166][2] ), .COUT(\CARRYB[167][1] ), .SUM(\SUMB[167][1] ) );
  FADDER S3_167_2 ( .CIN(\ab[167][2] ), .IN0(\CARRYB[166][2] ), .IN1(
        \ab[166][3] ), .COUT(\CARRYB[167][2] ), .SUM(\SUMB[167][2] ) );
  FADDER S1_166_0 ( .CIN(\ab[166][0] ), .IN0(\CARRYB[165][0] ), .IN1(
        \SUMB[165][1] ), .COUT(\CARRYB[166][0] ), .SUM(PRODUCT[166]) );
  FADDER S2_166_1 ( .CIN(\ab[166][1] ), .IN0(\CARRYB[165][1] ), .IN1(
        \SUMB[165][2] ), .COUT(\CARRYB[166][1] ), .SUM(\SUMB[166][1] ) );
  FADDER S3_166_2 ( .CIN(\ab[166][2] ), .IN0(\CARRYB[165][2] ), .IN1(
        \ab[165][3] ), .COUT(\CARRYB[166][2] ), .SUM(\SUMB[166][2] ) );
  FADDER S1_165_0 ( .CIN(\ab[165][0] ), .IN0(\CARRYB[164][0] ), .IN1(
        \SUMB[164][1] ), .COUT(\CARRYB[165][0] ), .SUM(PRODUCT[165]) );
  FADDER S2_165_1 ( .CIN(\ab[165][1] ), .IN0(\CARRYB[164][1] ), .IN1(
        \SUMB[164][2] ), .COUT(\CARRYB[165][1] ), .SUM(\SUMB[165][1] ) );
  FADDER S3_165_2 ( .CIN(\ab[165][2] ), .IN0(\CARRYB[164][2] ), .IN1(
        \ab[164][3] ), .COUT(\CARRYB[165][2] ), .SUM(\SUMB[165][2] ) );
  FADDER S1_164_0 ( .CIN(\ab[164][0] ), .IN0(\CARRYB[163][0] ), .IN1(
        \SUMB[163][1] ), .COUT(\CARRYB[164][0] ), .SUM(PRODUCT[164]) );
  FADDER S2_164_1 ( .CIN(\ab[164][1] ), .IN0(\CARRYB[163][1] ), .IN1(
        \SUMB[163][2] ), .COUT(\CARRYB[164][1] ), .SUM(\SUMB[164][1] ) );
  FADDER S3_164_2 ( .CIN(\ab[164][2] ), .IN0(\CARRYB[163][2] ), .IN1(
        \ab[163][3] ), .COUT(\CARRYB[164][2] ), .SUM(\SUMB[164][2] ) );
  FADDER S1_163_0 ( .CIN(\ab[163][0] ), .IN0(\CARRYB[162][0] ), .IN1(
        \SUMB[162][1] ), .COUT(\CARRYB[163][0] ), .SUM(PRODUCT[163]) );
  FADDER S2_163_1 ( .CIN(\ab[163][1] ), .IN0(\CARRYB[162][1] ), .IN1(
        \SUMB[162][2] ), .COUT(\CARRYB[163][1] ), .SUM(\SUMB[163][1] ) );
  FADDER S3_163_2 ( .CIN(\ab[163][2] ), .IN0(\CARRYB[162][2] ), .IN1(
        \ab[162][3] ), .COUT(\CARRYB[163][2] ), .SUM(\SUMB[163][2] ) );
  FADDER S1_162_0 ( .CIN(\ab[162][0] ), .IN0(\CARRYB[161][0] ), .IN1(
        \SUMB[161][1] ), .COUT(\CARRYB[162][0] ), .SUM(PRODUCT[162]) );
  FADDER S2_162_1 ( .CIN(\ab[162][1] ), .IN0(\CARRYB[161][1] ), .IN1(
        \SUMB[161][2] ), .COUT(\CARRYB[162][1] ), .SUM(\SUMB[162][1] ) );
  FADDER S3_162_2 ( .CIN(\ab[162][2] ), .IN0(\CARRYB[161][2] ), .IN1(
        \ab[161][3] ), .COUT(\CARRYB[162][2] ), .SUM(\SUMB[162][2] ) );
  FADDER S1_161_0 ( .CIN(\ab[161][0] ), .IN0(\CARRYB[160][0] ), .IN1(
        \SUMB[160][1] ), .COUT(\CARRYB[161][0] ), .SUM(PRODUCT[161]) );
  FADDER S2_161_1 ( .CIN(\ab[161][1] ), .IN0(\CARRYB[160][1] ), .IN1(
        \SUMB[160][2] ), .COUT(\CARRYB[161][1] ), .SUM(\SUMB[161][1] ) );
  FADDER S3_161_2 ( .CIN(\ab[161][2] ), .IN0(\CARRYB[160][2] ), .IN1(
        \ab[160][3] ), .COUT(\CARRYB[161][2] ), .SUM(\SUMB[161][2] ) );
  FADDER S1_160_0 ( .CIN(\ab[160][0] ), .IN0(\CARRYB[159][0] ), .IN1(
        \SUMB[159][1] ), .COUT(\CARRYB[160][0] ), .SUM(PRODUCT[160]) );
  FADDER S2_160_1 ( .CIN(\ab[160][1] ), .IN0(\CARRYB[159][1] ), .IN1(
        \SUMB[159][2] ), .COUT(\CARRYB[160][1] ), .SUM(\SUMB[160][1] ) );
  FADDER S3_160_2 ( .CIN(\ab[160][2] ), .IN0(\CARRYB[159][2] ), .IN1(
        \ab[159][3] ), .COUT(\CARRYB[160][2] ), .SUM(\SUMB[160][2] ) );
  FADDER S1_159_0 ( .CIN(\ab[159][0] ), .IN0(\CARRYB[158][0] ), .IN1(
        \SUMB[158][1] ), .COUT(\CARRYB[159][0] ), .SUM(PRODUCT[159]) );
  FADDER S2_159_1 ( .CIN(\ab[159][1] ), .IN0(\CARRYB[158][1] ), .IN1(
        \SUMB[158][2] ), .COUT(\CARRYB[159][1] ), .SUM(\SUMB[159][1] ) );
  FADDER S3_159_2 ( .CIN(\ab[159][2] ), .IN0(\CARRYB[158][2] ), .IN1(
        \ab[158][3] ), .COUT(\CARRYB[159][2] ), .SUM(\SUMB[159][2] ) );
  FADDER S1_158_0 ( .CIN(\ab[158][0] ), .IN0(\CARRYB[157][0] ), .IN1(
        \SUMB[157][1] ), .COUT(\CARRYB[158][0] ), .SUM(PRODUCT[158]) );
  FADDER S2_158_1 ( .CIN(\ab[158][1] ), .IN0(\CARRYB[157][1] ), .IN1(
        \SUMB[157][2] ), .COUT(\CARRYB[158][1] ), .SUM(\SUMB[158][1] ) );
  FADDER S3_158_2 ( .CIN(\ab[158][2] ), .IN0(\CARRYB[157][2] ), .IN1(
        \ab[157][3] ), .COUT(\CARRYB[158][2] ), .SUM(\SUMB[158][2] ) );
  FADDER S1_157_0 ( .CIN(\ab[157][0] ), .IN0(\CARRYB[156][0] ), .IN1(
        \SUMB[156][1] ), .COUT(\CARRYB[157][0] ), .SUM(PRODUCT[157]) );
  FADDER S2_157_1 ( .CIN(\ab[157][1] ), .IN0(\CARRYB[156][1] ), .IN1(
        \SUMB[156][2] ), .COUT(\CARRYB[157][1] ), .SUM(\SUMB[157][1] ) );
  FADDER S3_157_2 ( .CIN(\ab[157][2] ), .IN0(\CARRYB[156][2] ), .IN1(
        \ab[156][3] ), .COUT(\CARRYB[157][2] ), .SUM(\SUMB[157][2] ) );
  FADDER S1_156_0 ( .CIN(\ab[156][0] ), .IN0(\CARRYB[155][0] ), .IN1(
        \SUMB[155][1] ), .COUT(\CARRYB[156][0] ), .SUM(PRODUCT[156]) );
  FADDER S2_156_1 ( .CIN(\ab[156][1] ), .IN0(\CARRYB[155][1] ), .IN1(
        \SUMB[155][2] ), .COUT(\CARRYB[156][1] ), .SUM(\SUMB[156][1] ) );
  FADDER S3_156_2 ( .CIN(\ab[156][2] ), .IN0(\CARRYB[155][2] ), .IN1(
        \ab[155][3] ), .COUT(\CARRYB[156][2] ), .SUM(\SUMB[156][2] ) );
  FADDER S1_155_0 ( .CIN(\ab[155][0] ), .IN0(\CARRYB[154][0] ), .IN1(
        \SUMB[154][1] ), .COUT(\CARRYB[155][0] ), .SUM(PRODUCT[155]) );
  FADDER S2_155_1 ( .CIN(\ab[155][1] ), .IN0(\CARRYB[154][1] ), .IN1(
        \SUMB[154][2] ), .COUT(\CARRYB[155][1] ), .SUM(\SUMB[155][1] ) );
  FADDER S3_155_2 ( .CIN(\ab[155][2] ), .IN0(\CARRYB[154][2] ), .IN1(
        \ab[154][3] ), .COUT(\CARRYB[155][2] ), .SUM(\SUMB[155][2] ) );
  FADDER S1_154_0 ( .CIN(\ab[154][0] ), .IN0(\CARRYB[153][0] ), .IN1(
        \SUMB[153][1] ), .COUT(\CARRYB[154][0] ), .SUM(PRODUCT[154]) );
  FADDER S2_154_1 ( .CIN(\ab[154][1] ), .IN0(\CARRYB[153][1] ), .IN1(
        \SUMB[153][2] ), .COUT(\CARRYB[154][1] ), .SUM(\SUMB[154][1] ) );
  FADDER S3_154_2 ( .CIN(\ab[154][2] ), .IN0(\CARRYB[153][2] ), .IN1(
        \ab[153][3] ), .COUT(\CARRYB[154][2] ), .SUM(\SUMB[154][2] ) );
  FADDER S1_153_0 ( .CIN(\ab[153][0] ), .IN0(\CARRYB[152][0] ), .IN1(
        \SUMB[152][1] ), .COUT(\CARRYB[153][0] ), .SUM(PRODUCT[153]) );
  FADDER S2_153_1 ( .CIN(\ab[153][1] ), .IN0(\CARRYB[152][1] ), .IN1(
        \SUMB[152][2] ), .COUT(\CARRYB[153][1] ), .SUM(\SUMB[153][1] ) );
  FADDER S3_153_2 ( .CIN(\ab[153][2] ), .IN0(\CARRYB[152][2] ), .IN1(
        \ab[152][3] ), .COUT(\CARRYB[153][2] ), .SUM(\SUMB[153][2] ) );
  FADDER S1_152_0 ( .CIN(\ab[152][0] ), .IN0(\CARRYB[151][0] ), .IN1(
        \SUMB[151][1] ), .COUT(\CARRYB[152][0] ), .SUM(PRODUCT[152]) );
  FADDER S2_152_1 ( .CIN(\ab[152][1] ), .IN0(\CARRYB[151][1] ), .IN1(
        \SUMB[151][2] ), .COUT(\CARRYB[152][1] ), .SUM(\SUMB[152][1] ) );
  FADDER S3_152_2 ( .CIN(\ab[152][2] ), .IN0(\CARRYB[151][2] ), .IN1(
        \ab[151][3] ), .COUT(\CARRYB[152][2] ), .SUM(\SUMB[152][2] ) );
  FADDER S1_151_0 ( .CIN(\ab[151][0] ), .IN0(\CARRYB[150][0] ), .IN1(
        \SUMB[150][1] ), .COUT(\CARRYB[151][0] ), .SUM(PRODUCT[151]) );
  FADDER S2_151_1 ( .CIN(\ab[151][1] ), .IN0(\CARRYB[150][1] ), .IN1(
        \SUMB[150][2] ), .COUT(\CARRYB[151][1] ), .SUM(\SUMB[151][1] ) );
  FADDER S3_151_2 ( .CIN(\ab[151][2] ), .IN0(\CARRYB[150][2] ), .IN1(
        \ab[150][3] ), .COUT(\CARRYB[151][2] ), .SUM(\SUMB[151][2] ) );
  FADDER S1_150_0 ( .CIN(\ab[150][0] ), .IN0(\CARRYB[149][0] ), .IN1(
        \SUMB[149][1] ), .COUT(\CARRYB[150][0] ), .SUM(PRODUCT[150]) );
  FADDER S2_150_1 ( .CIN(\ab[150][1] ), .IN0(\CARRYB[149][1] ), .IN1(
        \SUMB[149][2] ), .COUT(\CARRYB[150][1] ), .SUM(\SUMB[150][1] ) );
  FADDER S3_150_2 ( .CIN(\ab[150][2] ), .IN0(\CARRYB[149][2] ), .IN1(
        \ab[149][3] ), .COUT(\CARRYB[150][2] ), .SUM(\SUMB[150][2] ) );
  FADDER S1_149_0 ( .CIN(\ab[149][0] ), .IN0(\CARRYB[148][0] ), .IN1(
        \SUMB[148][1] ), .COUT(\CARRYB[149][0] ), .SUM(PRODUCT[149]) );
  FADDER S2_149_1 ( .CIN(\ab[149][1] ), .IN0(\CARRYB[148][1] ), .IN1(
        \SUMB[148][2] ), .COUT(\CARRYB[149][1] ), .SUM(\SUMB[149][1] ) );
  FADDER S3_149_2 ( .CIN(\ab[149][2] ), .IN0(\CARRYB[148][2] ), .IN1(
        \ab[148][3] ), .COUT(\CARRYB[149][2] ), .SUM(\SUMB[149][2] ) );
  FADDER S1_148_0 ( .CIN(\ab[148][0] ), .IN0(\CARRYB[147][0] ), .IN1(
        \SUMB[147][1] ), .COUT(\CARRYB[148][0] ), .SUM(PRODUCT[148]) );
  FADDER S2_148_1 ( .CIN(\ab[148][1] ), .IN0(\CARRYB[147][1] ), .IN1(
        \SUMB[147][2] ), .COUT(\CARRYB[148][1] ), .SUM(\SUMB[148][1] ) );
  FADDER S3_148_2 ( .CIN(\ab[148][2] ), .IN0(\CARRYB[147][2] ), .IN1(
        \ab[147][3] ), .COUT(\CARRYB[148][2] ), .SUM(\SUMB[148][2] ) );
  FADDER S1_147_0 ( .CIN(\ab[147][0] ), .IN0(\CARRYB[146][0] ), .IN1(
        \SUMB[146][1] ), .COUT(\CARRYB[147][0] ), .SUM(PRODUCT[147]) );
  FADDER S2_147_1 ( .CIN(\ab[147][1] ), .IN0(\CARRYB[146][1] ), .IN1(
        \SUMB[146][2] ), .COUT(\CARRYB[147][1] ), .SUM(\SUMB[147][1] ) );
  FADDER S3_147_2 ( .CIN(\ab[147][2] ), .IN0(\CARRYB[146][2] ), .IN1(
        \ab[146][3] ), .COUT(\CARRYB[147][2] ), .SUM(\SUMB[147][2] ) );
  FADDER S1_146_0 ( .CIN(\ab[146][0] ), .IN0(\CARRYB[145][0] ), .IN1(
        \SUMB[145][1] ), .COUT(\CARRYB[146][0] ), .SUM(PRODUCT[146]) );
  FADDER S2_146_1 ( .CIN(\ab[146][1] ), .IN0(\CARRYB[145][1] ), .IN1(
        \SUMB[145][2] ), .COUT(\CARRYB[146][1] ), .SUM(\SUMB[146][1] ) );
  FADDER S3_146_2 ( .CIN(\ab[146][2] ), .IN0(\CARRYB[145][2] ), .IN1(
        \ab[145][3] ), .COUT(\CARRYB[146][2] ), .SUM(\SUMB[146][2] ) );
  FADDER S1_145_0 ( .CIN(\ab[145][0] ), .IN0(\CARRYB[144][0] ), .IN1(
        \SUMB[144][1] ), .COUT(\CARRYB[145][0] ), .SUM(PRODUCT[145]) );
  FADDER S2_145_1 ( .CIN(\ab[145][1] ), .IN0(\CARRYB[144][1] ), .IN1(
        \SUMB[144][2] ), .COUT(\CARRYB[145][1] ), .SUM(\SUMB[145][1] ) );
  FADDER S3_145_2 ( .CIN(\ab[145][2] ), .IN0(\CARRYB[144][2] ), .IN1(
        \ab[144][3] ), .COUT(\CARRYB[145][2] ), .SUM(\SUMB[145][2] ) );
  FADDER S1_144_0 ( .CIN(\ab[144][0] ), .IN0(\CARRYB[143][0] ), .IN1(
        \SUMB[143][1] ), .COUT(\CARRYB[144][0] ), .SUM(PRODUCT[144]) );
  FADDER S2_144_1 ( .CIN(\ab[144][1] ), .IN0(\CARRYB[143][1] ), .IN1(
        \SUMB[143][2] ), .COUT(\CARRYB[144][1] ), .SUM(\SUMB[144][1] ) );
  FADDER S3_144_2 ( .CIN(\ab[144][2] ), .IN0(\CARRYB[143][2] ), .IN1(
        \ab[143][3] ), .COUT(\CARRYB[144][2] ), .SUM(\SUMB[144][2] ) );
  FADDER S1_143_0 ( .CIN(\ab[143][0] ), .IN0(\CARRYB[142][0] ), .IN1(
        \SUMB[142][1] ), .COUT(\CARRYB[143][0] ), .SUM(PRODUCT[143]) );
  FADDER S2_143_1 ( .CIN(\ab[143][1] ), .IN0(\CARRYB[142][1] ), .IN1(
        \SUMB[142][2] ), .COUT(\CARRYB[143][1] ), .SUM(\SUMB[143][1] ) );
  FADDER S3_143_2 ( .CIN(\ab[143][2] ), .IN0(\CARRYB[142][2] ), .IN1(
        \ab[142][3] ), .COUT(\CARRYB[143][2] ), .SUM(\SUMB[143][2] ) );
  FADDER S1_142_0 ( .CIN(\ab[142][0] ), .IN0(\CARRYB[141][0] ), .IN1(
        \SUMB[141][1] ), .COUT(\CARRYB[142][0] ), .SUM(PRODUCT[142]) );
  FADDER S2_142_1 ( .CIN(\ab[142][1] ), .IN0(\CARRYB[141][1] ), .IN1(
        \SUMB[141][2] ), .COUT(\CARRYB[142][1] ), .SUM(\SUMB[142][1] ) );
  FADDER S3_142_2 ( .CIN(\ab[142][2] ), .IN0(\CARRYB[141][2] ), .IN1(
        \ab[141][3] ), .COUT(\CARRYB[142][2] ), .SUM(\SUMB[142][2] ) );
  FADDER S1_141_0 ( .CIN(\ab[141][0] ), .IN0(\CARRYB[140][0] ), .IN1(
        \SUMB[140][1] ), .COUT(\CARRYB[141][0] ), .SUM(PRODUCT[141]) );
  FADDER S2_141_1 ( .CIN(\ab[141][1] ), .IN0(\CARRYB[140][1] ), .IN1(
        \SUMB[140][2] ), .COUT(\CARRYB[141][1] ), .SUM(\SUMB[141][1] ) );
  FADDER S3_141_2 ( .CIN(\ab[141][2] ), .IN0(\CARRYB[140][2] ), .IN1(
        \ab[140][3] ), .COUT(\CARRYB[141][2] ), .SUM(\SUMB[141][2] ) );
  FADDER S1_140_0 ( .CIN(\ab[140][0] ), .IN0(\CARRYB[139][0] ), .IN1(
        \SUMB[139][1] ), .COUT(\CARRYB[140][0] ), .SUM(PRODUCT[140]) );
  FADDER S2_140_1 ( .CIN(\ab[140][1] ), .IN0(\CARRYB[139][1] ), .IN1(
        \SUMB[139][2] ), .COUT(\CARRYB[140][1] ), .SUM(\SUMB[140][1] ) );
  FADDER S3_140_2 ( .CIN(\ab[140][2] ), .IN0(\CARRYB[139][2] ), .IN1(
        \ab[139][3] ), .COUT(\CARRYB[140][2] ), .SUM(\SUMB[140][2] ) );
  FADDER S1_139_0 ( .CIN(\ab[139][0] ), .IN0(\CARRYB[138][0] ), .IN1(
        \SUMB[138][1] ), .COUT(\CARRYB[139][0] ), .SUM(PRODUCT[139]) );
  FADDER S2_139_1 ( .CIN(\ab[139][1] ), .IN0(\CARRYB[138][1] ), .IN1(
        \SUMB[138][2] ), .COUT(\CARRYB[139][1] ), .SUM(\SUMB[139][1] ) );
  FADDER S3_139_2 ( .CIN(\ab[139][2] ), .IN0(\CARRYB[138][2] ), .IN1(
        \ab[138][3] ), .COUT(\CARRYB[139][2] ), .SUM(\SUMB[139][2] ) );
  FADDER S1_138_0 ( .CIN(\ab[138][0] ), .IN0(\CARRYB[137][0] ), .IN1(
        \SUMB[137][1] ), .COUT(\CARRYB[138][0] ), .SUM(PRODUCT[138]) );
  FADDER S2_138_1 ( .CIN(\ab[138][1] ), .IN0(\CARRYB[137][1] ), .IN1(
        \SUMB[137][2] ), .COUT(\CARRYB[138][1] ), .SUM(\SUMB[138][1] ) );
  FADDER S3_138_2 ( .CIN(\ab[138][2] ), .IN0(\CARRYB[137][2] ), .IN1(
        \ab[137][3] ), .COUT(\CARRYB[138][2] ), .SUM(\SUMB[138][2] ) );
  FADDER S1_137_0 ( .CIN(\ab[137][0] ), .IN0(\CARRYB[136][0] ), .IN1(
        \SUMB[136][1] ), .COUT(\CARRYB[137][0] ), .SUM(PRODUCT[137]) );
  FADDER S2_137_1 ( .CIN(\ab[137][1] ), .IN0(\CARRYB[136][1] ), .IN1(
        \SUMB[136][2] ), .COUT(\CARRYB[137][1] ), .SUM(\SUMB[137][1] ) );
  FADDER S3_137_2 ( .CIN(\ab[137][2] ), .IN0(\CARRYB[136][2] ), .IN1(
        \ab[136][3] ), .COUT(\CARRYB[137][2] ), .SUM(\SUMB[137][2] ) );
  FADDER S1_136_0 ( .CIN(\ab[136][0] ), .IN0(\CARRYB[135][0] ), .IN1(
        \SUMB[135][1] ), .COUT(\CARRYB[136][0] ), .SUM(PRODUCT[136]) );
  FADDER S2_136_1 ( .CIN(\ab[136][1] ), .IN0(\CARRYB[135][1] ), .IN1(
        \SUMB[135][2] ), .COUT(\CARRYB[136][1] ), .SUM(\SUMB[136][1] ) );
  FADDER S3_136_2 ( .CIN(\ab[136][2] ), .IN0(\CARRYB[135][2] ), .IN1(
        \ab[135][3] ), .COUT(\CARRYB[136][2] ), .SUM(\SUMB[136][2] ) );
  FADDER S1_135_0 ( .CIN(\ab[135][0] ), .IN0(\CARRYB[134][0] ), .IN1(
        \SUMB[134][1] ), .COUT(\CARRYB[135][0] ), .SUM(PRODUCT[135]) );
  FADDER S2_135_1 ( .CIN(\ab[135][1] ), .IN0(\CARRYB[134][1] ), .IN1(
        \SUMB[134][2] ), .COUT(\CARRYB[135][1] ), .SUM(\SUMB[135][1] ) );
  FADDER S3_135_2 ( .CIN(\ab[135][2] ), .IN0(\CARRYB[134][2] ), .IN1(
        \ab[134][3] ), .COUT(\CARRYB[135][2] ), .SUM(\SUMB[135][2] ) );
  FADDER S1_134_0 ( .CIN(\ab[134][0] ), .IN0(\CARRYB[133][0] ), .IN1(
        \SUMB[133][1] ), .COUT(\CARRYB[134][0] ), .SUM(PRODUCT[134]) );
  FADDER S2_134_1 ( .CIN(\ab[134][1] ), .IN0(\CARRYB[133][1] ), .IN1(
        \SUMB[133][2] ), .COUT(\CARRYB[134][1] ), .SUM(\SUMB[134][1] ) );
  FADDER S3_134_2 ( .CIN(\ab[134][2] ), .IN0(\CARRYB[133][2] ), .IN1(
        \ab[133][3] ), .COUT(\CARRYB[134][2] ), .SUM(\SUMB[134][2] ) );
  FADDER S1_133_0 ( .CIN(\ab[133][0] ), .IN0(\CARRYB[132][0] ), .IN1(
        \SUMB[132][1] ), .COUT(\CARRYB[133][0] ), .SUM(PRODUCT[133]) );
  FADDER S2_133_1 ( .CIN(\ab[133][1] ), .IN0(\CARRYB[132][1] ), .IN1(
        \SUMB[132][2] ), .COUT(\CARRYB[133][1] ), .SUM(\SUMB[133][1] ) );
  FADDER S3_133_2 ( .CIN(\ab[133][2] ), .IN0(\CARRYB[132][2] ), .IN1(
        \ab[132][3] ), .COUT(\CARRYB[133][2] ), .SUM(\SUMB[133][2] ) );
  FADDER S1_132_0 ( .CIN(\ab[132][0] ), .IN0(\CARRYB[131][0] ), .IN1(
        \SUMB[131][1] ), .COUT(\CARRYB[132][0] ), .SUM(PRODUCT[132]) );
  FADDER S2_132_1 ( .CIN(\ab[132][1] ), .IN0(\CARRYB[131][1] ), .IN1(
        \SUMB[131][2] ), .COUT(\CARRYB[132][1] ), .SUM(\SUMB[132][1] ) );
  FADDER S3_132_2 ( .CIN(\ab[132][2] ), .IN0(\CARRYB[131][2] ), .IN1(
        \ab[131][3] ), .COUT(\CARRYB[132][2] ), .SUM(\SUMB[132][2] ) );
  FADDER S1_131_0 ( .CIN(\ab[131][0] ), .IN0(\CARRYB[130][0] ), .IN1(
        \SUMB[130][1] ), .COUT(\CARRYB[131][0] ), .SUM(PRODUCT[131]) );
  FADDER S2_131_1 ( .CIN(\ab[131][1] ), .IN0(\CARRYB[130][1] ), .IN1(
        \SUMB[130][2] ), .COUT(\CARRYB[131][1] ), .SUM(\SUMB[131][1] ) );
  FADDER S3_131_2 ( .CIN(\ab[131][2] ), .IN0(\CARRYB[130][2] ), .IN1(
        \ab[130][3] ), .COUT(\CARRYB[131][2] ), .SUM(\SUMB[131][2] ) );
  FADDER S1_130_0 ( .CIN(\ab[130][0] ), .IN0(\CARRYB[129][0] ), .IN1(
        \SUMB[129][1] ), .COUT(\CARRYB[130][0] ), .SUM(PRODUCT[130]) );
  FADDER S2_130_1 ( .CIN(\ab[130][1] ), .IN0(\CARRYB[129][1] ), .IN1(
        \SUMB[129][2] ), .COUT(\CARRYB[130][1] ), .SUM(\SUMB[130][1] ) );
  FADDER S3_130_2 ( .CIN(\ab[130][2] ), .IN0(\CARRYB[129][2] ), .IN1(
        \ab[129][3] ), .COUT(\CARRYB[130][2] ), .SUM(\SUMB[130][2] ) );
  FADDER S1_129_0 ( .CIN(\ab[129][0] ), .IN0(\CARRYB[128][0] ), .IN1(
        \SUMB[128][1] ), .COUT(\CARRYB[129][0] ), .SUM(PRODUCT[129]) );
  FADDER S2_129_1 ( .CIN(\ab[129][1] ), .IN0(\CARRYB[128][1] ), .IN1(
        \SUMB[128][2] ), .COUT(\CARRYB[129][1] ), .SUM(\SUMB[129][1] ) );
  FADDER S3_129_2 ( .CIN(\ab[129][2] ), .IN0(\CARRYB[128][2] ), .IN1(
        \ab[128][3] ), .COUT(\CARRYB[129][2] ), .SUM(\SUMB[129][2] ) );
  FADDER S1_128_0 ( .CIN(\ab[128][0] ), .IN0(\CARRYB[127][0] ), .IN1(
        \SUMB[127][1] ), .COUT(\CARRYB[128][0] ), .SUM(PRODUCT[128]) );
  FADDER S2_128_1 ( .CIN(\ab[128][1] ), .IN0(\CARRYB[127][1] ), .IN1(
        \SUMB[127][2] ), .COUT(\CARRYB[128][1] ), .SUM(\SUMB[128][1] ) );
  FADDER S3_128_2 ( .CIN(\ab[128][2] ), .IN0(\CARRYB[127][2] ), .IN1(
        \ab[127][3] ), .COUT(\CARRYB[128][2] ), .SUM(\SUMB[128][2] ) );
  FADDER S1_127_0 ( .CIN(\ab[127][0] ), .IN0(\CARRYB[126][0] ), .IN1(
        \SUMB[126][1] ), .COUT(\CARRYB[127][0] ), .SUM(PRODUCT[127]) );
  FADDER S2_127_1 ( .CIN(\ab[127][1] ), .IN0(\CARRYB[126][1] ), .IN1(
        \SUMB[126][2] ), .COUT(\CARRYB[127][1] ), .SUM(\SUMB[127][1] ) );
  FADDER S3_127_2 ( .CIN(\ab[127][2] ), .IN0(\CARRYB[126][2] ), .IN1(
        \ab[126][3] ), .COUT(\CARRYB[127][2] ), .SUM(\SUMB[127][2] ) );
  FADDER S1_126_0 ( .CIN(\ab[126][0] ), .IN0(\CARRYB[125][0] ), .IN1(
        \SUMB[125][1] ), .COUT(\CARRYB[126][0] ), .SUM(PRODUCT[126]) );
  FADDER S2_126_1 ( .CIN(\ab[126][1] ), .IN0(\CARRYB[125][1] ), .IN1(
        \SUMB[125][2] ), .COUT(\CARRYB[126][1] ), .SUM(\SUMB[126][1] ) );
  FADDER S3_126_2 ( .CIN(\ab[126][2] ), .IN0(\CARRYB[125][2] ), .IN1(
        \ab[125][3] ), .COUT(\CARRYB[126][2] ), .SUM(\SUMB[126][2] ) );
  FADDER S1_125_0 ( .CIN(\ab[125][0] ), .IN0(\CARRYB[124][0] ), .IN1(
        \SUMB[124][1] ), .COUT(\CARRYB[125][0] ), .SUM(PRODUCT[125]) );
  FADDER S2_125_1 ( .CIN(\ab[125][1] ), .IN0(\CARRYB[124][1] ), .IN1(
        \SUMB[124][2] ), .COUT(\CARRYB[125][1] ), .SUM(\SUMB[125][1] ) );
  FADDER S3_125_2 ( .CIN(\ab[125][2] ), .IN0(\CARRYB[124][2] ), .IN1(
        \ab[124][3] ), .COUT(\CARRYB[125][2] ), .SUM(\SUMB[125][2] ) );
  FADDER S1_124_0 ( .CIN(\ab[124][0] ), .IN0(\CARRYB[123][0] ), .IN1(
        \SUMB[123][1] ), .COUT(\CARRYB[124][0] ), .SUM(PRODUCT[124]) );
  FADDER S2_124_1 ( .CIN(\ab[124][1] ), .IN0(\CARRYB[123][1] ), .IN1(
        \SUMB[123][2] ), .COUT(\CARRYB[124][1] ), .SUM(\SUMB[124][1] ) );
  FADDER S3_124_2 ( .CIN(\ab[124][2] ), .IN0(\CARRYB[123][2] ), .IN1(
        \ab[123][3] ), .COUT(\CARRYB[124][2] ), .SUM(\SUMB[124][2] ) );
  FADDER S1_123_0 ( .CIN(\ab[123][0] ), .IN0(\CARRYB[122][0] ), .IN1(
        \SUMB[122][1] ), .COUT(\CARRYB[123][0] ), .SUM(PRODUCT[123]) );
  FADDER S2_123_1 ( .CIN(\ab[123][1] ), .IN0(\CARRYB[122][1] ), .IN1(
        \SUMB[122][2] ), .COUT(\CARRYB[123][1] ), .SUM(\SUMB[123][1] ) );
  FADDER S3_123_2 ( .CIN(\ab[123][2] ), .IN0(\CARRYB[122][2] ), .IN1(
        \ab[122][3] ), .COUT(\CARRYB[123][2] ), .SUM(\SUMB[123][2] ) );
  FADDER S1_122_0 ( .CIN(\ab[122][0] ), .IN0(\CARRYB[121][0] ), .IN1(
        \SUMB[121][1] ), .COUT(\CARRYB[122][0] ), .SUM(PRODUCT[122]) );
  FADDER S2_122_1 ( .CIN(\ab[122][1] ), .IN0(\CARRYB[121][1] ), .IN1(
        \SUMB[121][2] ), .COUT(\CARRYB[122][1] ), .SUM(\SUMB[122][1] ) );
  FADDER S3_122_2 ( .CIN(\ab[122][2] ), .IN0(\CARRYB[121][2] ), .IN1(
        \ab[121][3] ), .COUT(\CARRYB[122][2] ), .SUM(\SUMB[122][2] ) );
  FADDER S1_121_0 ( .CIN(\ab[121][0] ), .IN0(\CARRYB[120][0] ), .IN1(
        \SUMB[120][1] ), .COUT(\CARRYB[121][0] ), .SUM(PRODUCT[121]) );
  FADDER S2_121_1 ( .CIN(\ab[121][1] ), .IN0(\CARRYB[120][1] ), .IN1(
        \SUMB[120][2] ), .COUT(\CARRYB[121][1] ), .SUM(\SUMB[121][1] ) );
  FADDER S3_121_2 ( .CIN(\ab[121][2] ), .IN0(\CARRYB[120][2] ), .IN1(
        \ab[120][3] ), .COUT(\CARRYB[121][2] ), .SUM(\SUMB[121][2] ) );
  FADDER S1_120_0 ( .CIN(\ab[120][0] ), .IN0(\CARRYB[119][0] ), .IN1(
        \SUMB[119][1] ), .COUT(\CARRYB[120][0] ), .SUM(PRODUCT[120]) );
  FADDER S2_120_1 ( .CIN(\ab[120][1] ), .IN0(\CARRYB[119][1] ), .IN1(
        \SUMB[119][2] ), .COUT(\CARRYB[120][1] ), .SUM(\SUMB[120][1] ) );
  FADDER S3_120_2 ( .CIN(\ab[120][2] ), .IN0(\CARRYB[119][2] ), .IN1(
        \ab[119][3] ), .COUT(\CARRYB[120][2] ), .SUM(\SUMB[120][2] ) );
  FADDER S1_119_0 ( .CIN(\ab[119][0] ), .IN0(\CARRYB[118][0] ), .IN1(
        \SUMB[118][1] ), .COUT(\CARRYB[119][0] ), .SUM(PRODUCT[119]) );
  FADDER S2_119_1 ( .CIN(\ab[119][1] ), .IN0(\CARRYB[118][1] ), .IN1(
        \SUMB[118][2] ), .COUT(\CARRYB[119][1] ), .SUM(\SUMB[119][1] ) );
  FADDER S3_119_2 ( .CIN(\ab[119][2] ), .IN0(\CARRYB[118][2] ), .IN1(
        \ab[118][3] ), .COUT(\CARRYB[119][2] ), .SUM(\SUMB[119][2] ) );
  FADDER S1_118_0 ( .CIN(\ab[118][0] ), .IN0(\CARRYB[117][0] ), .IN1(
        \SUMB[117][1] ), .COUT(\CARRYB[118][0] ), .SUM(PRODUCT[118]) );
  FADDER S2_118_1 ( .CIN(\ab[118][1] ), .IN0(\CARRYB[117][1] ), .IN1(
        \SUMB[117][2] ), .COUT(\CARRYB[118][1] ), .SUM(\SUMB[118][1] ) );
  FADDER S3_118_2 ( .CIN(\ab[118][2] ), .IN0(\CARRYB[117][2] ), .IN1(
        \ab[117][3] ), .COUT(\CARRYB[118][2] ), .SUM(\SUMB[118][2] ) );
  FADDER S1_117_0 ( .CIN(\ab[117][0] ), .IN0(\CARRYB[116][0] ), .IN1(
        \SUMB[116][1] ), .COUT(\CARRYB[117][0] ), .SUM(PRODUCT[117]) );
  FADDER S2_117_1 ( .CIN(\ab[117][1] ), .IN0(\CARRYB[116][1] ), .IN1(
        \SUMB[116][2] ), .COUT(\CARRYB[117][1] ), .SUM(\SUMB[117][1] ) );
  FADDER S3_117_2 ( .CIN(\ab[117][2] ), .IN0(\CARRYB[116][2] ), .IN1(
        \ab[116][3] ), .COUT(\CARRYB[117][2] ), .SUM(\SUMB[117][2] ) );
  FADDER S1_116_0 ( .CIN(\ab[116][0] ), .IN0(\CARRYB[115][0] ), .IN1(
        \SUMB[115][1] ), .COUT(\CARRYB[116][0] ), .SUM(PRODUCT[116]) );
  FADDER S2_116_1 ( .CIN(\ab[116][1] ), .IN0(\CARRYB[115][1] ), .IN1(
        \SUMB[115][2] ), .COUT(\CARRYB[116][1] ), .SUM(\SUMB[116][1] ) );
  FADDER S3_116_2 ( .CIN(\ab[116][2] ), .IN0(\CARRYB[115][2] ), .IN1(
        \ab[115][3] ), .COUT(\CARRYB[116][2] ), .SUM(\SUMB[116][2] ) );
  FADDER S1_115_0 ( .CIN(\ab[115][0] ), .IN0(\CARRYB[114][0] ), .IN1(
        \SUMB[114][1] ), .COUT(\CARRYB[115][0] ), .SUM(PRODUCT[115]) );
  FADDER S2_115_1 ( .CIN(\ab[115][1] ), .IN0(\CARRYB[114][1] ), .IN1(
        \SUMB[114][2] ), .COUT(\CARRYB[115][1] ), .SUM(\SUMB[115][1] ) );
  FADDER S3_115_2 ( .CIN(\ab[115][2] ), .IN0(\CARRYB[114][2] ), .IN1(
        \ab[114][3] ), .COUT(\CARRYB[115][2] ), .SUM(\SUMB[115][2] ) );
  FADDER S1_114_0 ( .CIN(\ab[114][0] ), .IN0(\CARRYB[113][0] ), .IN1(
        \SUMB[113][1] ), .COUT(\CARRYB[114][0] ), .SUM(PRODUCT[114]) );
  FADDER S2_114_1 ( .CIN(\ab[114][1] ), .IN0(\CARRYB[113][1] ), .IN1(
        \SUMB[113][2] ), .COUT(\CARRYB[114][1] ), .SUM(\SUMB[114][1] ) );
  FADDER S3_114_2 ( .CIN(\ab[114][2] ), .IN0(\CARRYB[113][2] ), .IN1(
        \ab[113][3] ), .COUT(\CARRYB[114][2] ), .SUM(\SUMB[114][2] ) );
  FADDER S1_113_0 ( .CIN(\ab[113][0] ), .IN0(\CARRYB[112][0] ), .IN1(
        \SUMB[112][1] ), .COUT(\CARRYB[113][0] ), .SUM(PRODUCT[113]) );
  FADDER S2_113_1 ( .CIN(\ab[113][1] ), .IN0(\CARRYB[112][1] ), .IN1(
        \SUMB[112][2] ), .COUT(\CARRYB[113][1] ), .SUM(\SUMB[113][1] ) );
  FADDER S3_113_2 ( .CIN(\ab[113][2] ), .IN0(\CARRYB[112][2] ), .IN1(
        \ab[112][3] ), .COUT(\CARRYB[113][2] ), .SUM(\SUMB[113][2] ) );
  FADDER S1_112_0 ( .CIN(\ab[112][0] ), .IN0(\CARRYB[111][0] ), .IN1(
        \SUMB[111][1] ), .COUT(\CARRYB[112][0] ), .SUM(PRODUCT[112]) );
  FADDER S2_112_1 ( .CIN(\ab[112][1] ), .IN0(\CARRYB[111][1] ), .IN1(
        \SUMB[111][2] ), .COUT(\CARRYB[112][1] ), .SUM(\SUMB[112][1] ) );
  FADDER S3_112_2 ( .CIN(\ab[112][2] ), .IN0(\CARRYB[111][2] ), .IN1(
        \ab[111][3] ), .COUT(\CARRYB[112][2] ), .SUM(\SUMB[112][2] ) );
  FADDER S1_111_0 ( .CIN(\ab[111][0] ), .IN0(\CARRYB[110][0] ), .IN1(
        \SUMB[110][1] ), .COUT(\CARRYB[111][0] ), .SUM(PRODUCT[111]) );
  FADDER S2_111_1 ( .CIN(\ab[111][1] ), .IN0(\CARRYB[110][1] ), .IN1(
        \SUMB[110][2] ), .COUT(\CARRYB[111][1] ), .SUM(\SUMB[111][1] ) );
  FADDER S3_111_2 ( .CIN(\ab[111][2] ), .IN0(\CARRYB[110][2] ), .IN1(
        \ab[110][3] ), .COUT(\CARRYB[111][2] ), .SUM(\SUMB[111][2] ) );
  FADDER S1_110_0 ( .CIN(\ab[110][0] ), .IN0(\CARRYB[109][0] ), .IN1(
        \SUMB[109][1] ), .COUT(\CARRYB[110][0] ), .SUM(PRODUCT[110]) );
  FADDER S2_110_1 ( .CIN(\ab[110][1] ), .IN0(\CARRYB[109][1] ), .IN1(
        \SUMB[109][2] ), .COUT(\CARRYB[110][1] ), .SUM(\SUMB[110][1] ) );
  FADDER S3_110_2 ( .CIN(\ab[110][2] ), .IN0(\CARRYB[109][2] ), .IN1(
        \ab[109][3] ), .COUT(\CARRYB[110][2] ), .SUM(\SUMB[110][2] ) );
  FADDER S1_109_0 ( .CIN(\ab[109][0] ), .IN0(\CARRYB[108][0] ), .IN1(
        \SUMB[108][1] ), .COUT(\CARRYB[109][0] ), .SUM(PRODUCT[109]) );
  FADDER S2_109_1 ( .CIN(\ab[109][1] ), .IN0(\CARRYB[108][1] ), .IN1(
        \SUMB[108][2] ), .COUT(\CARRYB[109][1] ), .SUM(\SUMB[109][1] ) );
  FADDER S3_109_2 ( .CIN(\ab[109][2] ), .IN0(\CARRYB[108][2] ), .IN1(
        \ab[108][3] ), .COUT(\CARRYB[109][2] ), .SUM(\SUMB[109][2] ) );
  FADDER S1_108_0 ( .CIN(\ab[108][0] ), .IN0(\CARRYB[107][0] ), .IN1(
        \SUMB[107][1] ), .COUT(\CARRYB[108][0] ), .SUM(PRODUCT[108]) );
  FADDER S2_108_1 ( .CIN(\ab[108][1] ), .IN0(\CARRYB[107][1] ), .IN1(
        \SUMB[107][2] ), .COUT(\CARRYB[108][1] ), .SUM(\SUMB[108][1] ) );
  FADDER S3_108_2 ( .CIN(\ab[108][2] ), .IN0(\CARRYB[107][2] ), .IN1(
        \ab[107][3] ), .COUT(\CARRYB[108][2] ), .SUM(\SUMB[108][2] ) );
  FADDER S1_107_0 ( .CIN(\ab[107][0] ), .IN0(\CARRYB[106][0] ), .IN1(
        \SUMB[106][1] ), .COUT(\CARRYB[107][0] ), .SUM(PRODUCT[107]) );
  FADDER S2_107_1 ( .CIN(\ab[107][1] ), .IN0(\CARRYB[106][1] ), .IN1(
        \SUMB[106][2] ), .COUT(\CARRYB[107][1] ), .SUM(\SUMB[107][1] ) );
  FADDER S3_107_2 ( .CIN(\ab[107][2] ), .IN0(\CARRYB[106][2] ), .IN1(
        \ab[106][3] ), .COUT(\CARRYB[107][2] ), .SUM(\SUMB[107][2] ) );
  FADDER S1_106_0 ( .CIN(\ab[106][0] ), .IN0(\CARRYB[105][0] ), .IN1(
        \SUMB[105][1] ), .COUT(\CARRYB[106][0] ), .SUM(PRODUCT[106]) );
  FADDER S2_106_1 ( .CIN(\ab[106][1] ), .IN0(\CARRYB[105][1] ), .IN1(
        \SUMB[105][2] ), .COUT(\CARRYB[106][1] ), .SUM(\SUMB[106][1] ) );
  FADDER S3_106_2 ( .CIN(\ab[106][2] ), .IN0(\CARRYB[105][2] ), .IN1(
        \ab[105][3] ), .COUT(\CARRYB[106][2] ), .SUM(\SUMB[106][2] ) );
  FADDER S1_105_0 ( .CIN(\ab[105][0] ), .IN0(\CARRYB[104][0] ), .IN1(
        \SUMB[104][1] ), .COUT(\CARRYB[105][0] ), .SUM(PRODUCT[105]) );
  FADDER S2_105_1 ( .CIN(\ab[105][1] ), .IN0(\CARRYB[104][1] ), .IN1(
        \SUMB[104][2] ), .COUT(\CARRYB[105][1] ), .SUM(\SUMB[105][1] ) );
  FADDER S3_105_2 ( .CIN(\ab[105][2] ), .IN0(\CARRYB[104][2] ), .IN1(
        \ab[104][3] ), .COUT(\CARRYB[105][2] ), .SUM(\SUMB[105][2] ) );
  FADDER S1_104_0 ( .CIN(\ab[104][0] ), .IN0(\CARRYB[103][0] ), .IN1(
        \SUMB[103][1] ), .COUT(\CARRYB[104][0] ), .SUM(PRODUCT[104]) );
  FADDER S2_104_1 ( .CIN(\ab[104][1] ), .IN0(\CARRYB[103][1] ), .IN1(
        \SUMB[103][2] ), .COUT(\CARRYB[104][1] ), .SUM(\SUMB[104][1] ) );
  FADDER S3_104_2 ( .CIN(\ab[104][2] ), .IN0(\CARRYB[103][2] ), .IN1(
        \ab[103][3] ), .COUT(\CARRYB[104][2] ), .SUM(\SUMB[104][2] ) );
  FADDER S1_103_0 ( .CIN(\ab[103][0] ), .IN0(\CARRYB[102][0] ), .IN1(
        \SUMB[102][1] ), .COUT(\CARRYB[103][0] ), .SUM(PRODUCT[103]) );
  FADDER S2_103_1 ( .CIN(\ab[103][1] ), .IN0(\CARRYB[102][1] ), .IN1(
        \SUMB[102][2] ), .COUT(\CARRYB[103][1] ), .SUM(\SUMB[103][1] ) );
  FADDER S3_103_2 ( .CIN(\ab[103][2] ), .IN0(\CARRYB[102][2] ), .IN1(
        \ab[102][3] ), .COUT(\CARRYB[103][2] ), .SUM(\SUMB[103][2] ) );
  FADDER S1_102_0 ( .CIN(\ab[102][0] ), .IN0(\CARRYB[101][0] ), .IN1(
        \SUMB[101][1] ), .COUT(\CARRYB[102][0] ), .SUM(PRODUCT[102]) );
  FADDER S2_102_1 ( .CIN(\ab[102][1] ), .IN0(\CARRYB[101][1] ), .IN1(
        \SUMB[101][2] ), .COUT(\CARRYB[102][1] ), .SUM(\SUMB[102][1] ) );
  FADDER S3_102_2 ( .CIN(\ab[102][2] ), .IN0(\CARRYB[101][2] ), .IN1(
        \ab[101][3] ), .COUT(\CARRYB[102][2] ), .SUM(\SUMB[102][2] ) );
  FADDER S1_101_0 ( .CIN(\ab[101][0] ), .IN0(\CARRYB[100][0] ), .IN1(
        \SUMB[100][1] ), .COUT(\CARRYB[101][0] ), .SUM(PRODUCT[101]) );
  FADDER S2_101_1 ( .CIN(\ab[101][1] ), .IN0(\CARRYB[100][1] ), .IN1(
        \SUMB[100][2] ), .COUT(\CARRYB[101][1] ), .SUM(\SUMB[101][1] ) );
  FADDER S3_101_2 ( .CIN(\ab[101][2] ), .IN0(\CARRYB[100][2] ), .IN1(
        \ab[100][3] ), .COUT(\CARRYB[101][2] ), .SUM(\SUMB[101][2] ) );
  FADDER S1_100_0 ( .CIN(\ab[100][0] ), .IN0(\CARRYB[99][0] ), .IN1(
        \SUMB[99][1] ), .COUT(\CARRYB[100][0] ), .SUM(PRODUCT[100]) );
  FADDER S2_100_1 ( .CIN(\ab[100][1] ), .IN0(\CARRYB[99][1] ), .IN1(
        \SUMB[99][2] ), .COUT(\CARRYB[100][1] ), .SUM(\SUMB[100][1] ) );
  FADDER S3_100_2 ( .CIN(\ab[100][2] ), .IN0(\CARRYB[99][2] ), .IN1(
        \ab[99][3] ), .COUT(\CARRYB[100][2] ), .SUM(\SUMB[100][2] ) );
  FADDER S1_99_0 ( .CIN(\ab[99][0] ), .IN0(\CARRYB[98][0] ), .IN1(
        \SUMB[98][1] ), .COUT(\CARRYB[99][0] ), .SUM(PRODUCT[99]) );
  FADDER S2_99_1 ( .CIN(\ab[99][1] ), .IN0(\CARRYB[98][1] ), .IN1(
        \SUMB[98][2] ), .COUT(\CARRYB[99][1] ), .SUM(\SUMB[99][1] ) );
  FADDER S3_99_2 ( .CIN(\ab[99][2] ), .IN0(\CARRYB[98][2] ), .IN1(\ab[98][3] ), 
        .COUT(\CARRYB[99][2] ), .SUM(\SUMB[99][2] ) );
  FADDER S1_98_0 ( .CIN(\ab[98][0] ), .IN0(\CARRYB[97][0] ), .IN1(
        \SUMB[97][1] ), .COUT(\CARRYB[98][0] ), .SUM(PRODUCT[98]) );
  FADDER S2_98_1 ( .CIN(\ab[98][1] ), .IN0(\CARRYB[97][1] ), .IN1(
        \SUMB[97][2] ), .COUT(\CARRYB[98][1] ), .SUM(\SUMB[98][1] ) );
  FADDER S3_98_2 ( .CIN(\ab[98][2] ), .IN0(\CARRYB[97][2] ), .IN1(\ab[97][3] ), 
        .COUT(\CARRYB[98][2] ), .SUM(\SUMB[98][2] ) );
  FADDER S1_97_0 ( .CIN(\ab[97][0] ), .IN0(\CARRYB[96][0] ), .IN1(
        \SUMB[96][1] ), .COUT(\CARRYB[97][0] ), .SUM(PRODUCT[97]) );
  FADDER S2_97_1 ( .CIN(\ab[97][1] ), .IN0(\CARRYB[96][1] ), .IN1(
        \SUMB[96][2] ), .COUT(\CARRYB[97][1] ), .SUM(\SUMB[97][1] ) );
  FADDER S3_97_2 ( .CIN(\ab[97][2] ), .IN0(\CARRYB[96][2] ), .IN1(\ab[96][3] ), 
        .COUT(\CARRYB[97][2] ), .SUM(\SUMB[97][2] ) );
  FADDER S1_96_0 ( .CIN(\ab[96][0] ), .IN0(\CARRYB[95][0] ), .IN1(
        \SUMB[95][1] ), .COUT(\CARRYB[96][0] ), .SUM(PRODUCT[96]) );
  FADDER S2_96_1 ( .CIN(\ab[96][1] ), .IN0(\CARRYB[95][1] ), .IN1(
        \SUMB[95][2] ), .COUT(\CARRYB[96][1] ), .SUM(\SUMB[96][1] ) );
  FADDER S3_96_2 ( .CIN(\ab[96][2] ), .IN0(\CARRYB[95][2] ), .IN1(\ab[95][3] ), 
        .COUT(\CARRYB[96][2] ), .SUM(\SUMB[96][2] ) );
  FADDER S1_95_0 ( .CIN(\ab[95][0] ), .IN0(\CARRYB[94][0] ), .IN1(
        \SUMB[94][1] ), .COUT(\CARRYB[95][0] ), .SUM(PRODUCT[95]) );
  FADDER S2_95_1 ( .CIN(\ab[95][1] ), .IN0(\CARRYB[94][1] ), .IN1(
        \SUMB[94][2] ), .COUT(\CARRYB[95][1] ), .SUM(\SUMB[95][1] ) );
  FADDER S3_95_2 ( .CIN(\ab[95][2] ), .IN0(\CARRYB[94][2] ), .IN1(\ab[94][3] ), 
        .COUT(\CARRYB[95][2] ), .SUM(\SUMB[95][2] ) );
  FADDER S1_94_0 ( .CIN(\ab[94][0] ), .IN0(\CARRYB[93][0] ), .IN1(
        \SUMB[93][1] ), .COUT(\CARRYB[94][0] ), .SUM(PRODUCT[94]) );
  FADDER S2_94_1 ( .CIN(\ab[94][1] ), .IN0(\CARRYB[93][1] ), .IN1(
        \SUMB[93][2] ), .COUT(\CARRYB[94][1] ), .SUM(\SUMB[94][1] ) );
  FADDER S3_94_2 ( .CIN(\ab[94][2] ), .IN0(\CARRYB[93][2] ), .IN1(\ab[93][3] ), 
        .COUT(\CARRYB[94][2] ), .SUM(\SUMB[94][2] ) );
  FADDER S1_93_0 ( .CIN(\ab[93][0] ), .IN0(\CARRYB[92][0] ), .IN1(
        \SUMB[92][1] ), .COUT(\CARRYB[93][0] ), .SUM(PRODUCT[93]) );
  FADDER S2_93_1 ( .CIN(\ab[93][1] ), .IN0(\CARRYB[92][1] ), .IN1(
        \SUMB[92][2] ), .COUT(\CARRYB[93][1] ), .SUM(\SUMB[93][1] ) );
  FADDER S3_93_2 ( .CIN(\ab[93][2] ), .IN0(\CARRYB[92][2] ), .IN1(\ab[92][3] ), 
        .COUT(\CARRYB[93][2] ), .SUM(\SUMB[93][2] ) );
  FADDER S1_92_0 ( .CIN(\ab[92][0] ), .IN0(\CARRYB[91][0] ), .IN1(
        \SUMB[91][1] ), .COUT(\CARRYB[92][0] ), .SUM(PRODUCT[92]) );
  FADDER S2_92_1 ( .CIN(\ab[92][1] ), .IN0(\CARRYB[91][1] ), .IN1(
        \SUMB[91][2] ), .COUT(\CARRYB[92][1] ), .SUM(\SUMB[92][1] ) );
  FADDER S3_92_2 ( .CIN(\ab[92][2] ), .IN0(\CARRYB[91][2] ), .IN1(\ab[91][3] ), 
        .COUT(\CARRYB[92][2] ), .SUM(\SUMB[92][2] ) );
  FADDER S1_91_0 ( .CIN(\ab[91][0] ), .IN0(\CARRYB[90][0] ), .IN1(
        \SUMB[90][1] ), .COUT(\CARRYB[91][0] ), .SUM(PRODUCT[91]) );
  FADDER S2_91_1 ( .CIN(\ab[91][1] ), .IN0(\CARRYB[90][1] ), .IN1(
        \SUMB[90][2] ), .COUT(\CARRYB[91][1] ), .SUM(\SUMB[91][1] ) );
  FADDER S3_91_2 ( .CIN(\ab[91][2] ), .IN0(\CARRYB[90][2] ), .IN1(\ab[90][3] ), 
        .COUT(\CARRYB[91][2] ), .SUM(\SUMB[91][2] ) );
  FADDER S1_90_0 ( .CIN(\ab[90][0] ), .IN0(\CARRYB[89][0] ), .IN1(
        \SUMB[89][1] ), .COUT(\CARRYB[90][0] ), .SUM(PRODUCT[90]) );
  FADDER S2_90_1 ( .CIN(\ab[90][1] ), .IN0(\CARRYB[89][1] ), .IN1(
        \SUMB[89][2] ), .COUT(\CARRYB[90][1] ), .SUM(\SUMB[90][1] ) );
  FADDER S3_90_2 ( .CIN(\ab[90][2] ), .IN0(\CARRYB[89][2] ), .IN1(\ab[89][3] ), 
        .COUT(\CARRYB[90][2] ), .SUM(\SUMB[90][2] ) );
  FADDER S1_89_0 ( .CIN(\ab[89][0] ), .IN0(\CARRYB[88][0] ), .IN1(
        \SUMB[88][1] ), .COUT(\CARRYB[89][0] ), .SUM(PRODUCT[89]) );
  FADDER S2_89_1 ( .CIN(\ab[89][1] ), .IN0(\CARRYB[88][1] ), .IN1(
        \SUMB[88][2] ), .COUT(\CARRYB[89][1] ), .SUM(\SUMB[89][1] ) );
  FADDER S3_89_2 ( .CIN(\ab[89][2] ), .IN0(\CARRYB[88][2] ), .IN1(\ab[88][3] ), 
        .COUT(\CARRYB[89][2] ), .SUM(\SUMB[89][2] ) );
  FADDER S1_88_0 ( .CIN(\ab[88][0] ), .IN0(\CARRYB[87][0] ), .IN1(
        \SUMB[87][1] ), .COUT(\CARRYB[88][0] ), .SUM(PRODUCT[88]) );
  FADDER S2_88_1 ( .CIN(\ab[88][1] ), .IN0(\CARRYB[87][1] ), .IN1(
        \SUMB[87][2] ), .COUT(\CARRYB[88][1] ), .SUM(\SUMB[88][1] ) );
  FADDER S3_88_2 ( .CIN(\ab[88][2] ), .IN0(\CARRYB[87][2] ), .IN1(\ab[87][3] ), 
        .COUT(\CARRYB[88][2] ), .SUM(\SUMB[88][2] ) );
  FADDER S1_87_0 ( .CIN(\ab[87][0] ), .IN0(\CARRYB[86][0] ), .IN1(
        \SUMB[86][1] ), .COUT(\CARRYB[87][0] ), .SUM(PRODUCT[87]) );
  FADDER S2_87_1 ( .CIN(\ab[87][1] ), .IN0(\CARRYB[86][1] ), .IN1(
        \SUMB[86][2] ), .COUT(\CARRYB[87][1] ), .SUM(\SUMB[87][1] ) );
  FADDER S3_87_2 ( .CIN(\ab[87][2] ), .IN0(\CARRYB[86][2] ), .IN1(\ab[86][3] ), 
        .COUT(\CARRYB[87][2] ), .SUM(\SUMB[87][2] ) );
  FADDER S1_86_0 ( .CIN(\ab[86][0] ), .IN0(\CARRYB[85][0] ), .IN1(
        \SUMB[85][1] ), .COUT(\CARRYB[86][0] ), .SUM(PRODUCT[86]) );
  FADDER S2_86_1 ( .CIN(\ab[86][1] ), .IN0(\CARRYB[85][1] ), .IN1(
        \SUMB[85][2] ), .COUT(\CARRYB[86][1] ), .SUM(\SUMB[86][1] ) );
  FADDER S3_86_2 ( .CIN(\ab[86][2] ), .IN0(\CARRYB[85][2] ), .IN1(\ab[85][3] ), 
        .COUT(\CARRYB[86][2] ), .SUM(\SUMB[86][2] ) );
  FADDER S1_85_0 ( .CIN(\ab[85][0] ), .IN0(\CARRYB[84][0] ), .IN1(
        \SUMB[84][1] ), .COUT(\CARRYB[85][0] ), .SUM(PRODUCT[85]) );
  FADDER S2_85_1 ( .CIN(\ab[85][1] ), .IN0(\CARRYB[84][1] ), .IN1(
        \SUMB[84][2] ), .COUT(\CARRYB[85][1] ), .SUM(\SUMB[85][1] ) );
  FADDER S3_85_2 ( .CIN(\ab[85][2] ), .IN0(\CARRYB[84][2] ), .IN1(\ab[84][3] ), 
        .COUT(\CARRYB[85][2] ), .SUM(\SUMB[85][2] ) );
  FADDER S1_84_0 ( .CIN(\ab[84][0] ), .IN0(\CARRYB[83][0] ), .IN1(
        \SUMB[83][1] ), .COUT(\CARRYB[84][0] ), .SUM(PRODUCT[84]) );
  FADDER S2_84_1 ( .CIN(\ab[84][1] ), .IN0(\CARRYB[83][1] ), .IN1(
        \SUMB[83][2] ), .COUT(\CARRYB[84][1] ), .SUM(\SUMB[84][1] ) );
  FADDER S3_84_2 ( .CIN(\ab[84][2] ), .IN0(\CARRYB[83][2] ), .IN1(\ab[83][3] ), 
        .COUT(\CARRYB[84][2] ), .SUM(\SUMB[84][2] ) );
  FADDER S1_83_0 ( .CIN(\ab[83][0] ), .IN0(\CARRYB[82][0] ), .IN1(
        \SUMB[82][1] ), .COUT(\CARRYB[83][0] ), .SUM(PRODUCT[83]) );
  FADDER S2_83_1 ( .CIN(\ab[83][1] ), .IN0(\CARRYB[82][1] ), .IN1(
        \SUMB[82][2] ), .COUT(\CARRYB[83][1] ), .SUM(\SUMB[83][1] ) );
  FADDER S3_83_2 ( .CIN(\ab[83][2] ), .IN0(\CARRYB[82][2] ), .IN1(\ab[82][3] ), 
        .COUT(\CARRYB[83][2] ), .SUM(\SUMB[83][2] ) );
  FADDER S1_82_0 ( .CIN(\ab[82][0] ), .IN0(\CARRYB[81][0] ), .IN1(
        \SUMB[81][1] ), .COUT(\CARRYB[82][0] ), .SUM(PRODUCT[82]) );
  FADDER S2_82_1 ( .CIN(\ab[82][1] ), .IN0(\CARRYB[81][1] ), .IN1(
        \SUMB[81][2] ), .COUT(\CARRYB[82][1] ), .SUM(\SUMB[82][1] ) );
  FADDER S3_82_2 ( .CIN(\ab[82][2] ), .IN0(\CARRYB[81][2] ), .IN1(\ab[81][3] ), 
        .COUT(\CARRYB[82][2] ), .SUM(\SUMB[82][2] ) );
  FADDER S1_81_0 ( .CIN(\ab[81][0] ), .IN0(\CARRYB[80][0] ), .IN1(
        \SUMB[80][1] ), .COUT(\CARRYB[81][0] ), .SUM(PRODUCT[81]) );
  FADDER S2_81_1 ( .CIN(\ab[81][1] ), .IN0(\CARRYB[80][1] ), .IN1(
        \SUMB[80][2] ), .COUT(\CARRYB[81][1] ), .SUM(\SUMB[81][1] ) );
  FADDER S3_81_2 ( .CIN(\ab[81][2] ), .IN0(\CARRYB[80][2] ), .IN1(\ab[80][3] ), 
        .COUT(\CARRYB[81][2] ), .SUM(\SUMB[81][2] ) );
  FADDER S1_80_0 ( .CIN(\ab[80][0] ), .IN0(\CARRYB[79][0] ), .IN1(
        \SUMB[79][1] ), .COUT(\CARRYB[80][0] ), .SUM(PRODUCT[80]) );
  FADDER S2_80_1 ( .CIN(\ab[80][1] ), .IN0(\CARRYB[79][1] ), .IN1(
        \SUMB[79][2] ), .COUT(\CARRYB[80][1] ), .SUM(\SUMB[80][1] ) );
  FADDER S3_80_2 ( .CIN(\ab[80][2] ), .IN0(\CARRYB[79][2] ), .IN1(\ab[79][3] ), 
        .COUT(\CARRYB[80][2] ), .SUM(\SUMB[80][2] ) );
  FADDER S1_79_0 ( .CIN(\ab[79][0] ), .IN0(\CARRYB[78][0] ), .IN1(
        \SUMB[78][1] ), .COUT(\CARRYB[79][0] ), .SUM(PRODUCT[79]) );
  FADDER S2_79_1 ( .CIN(\ab[79][1] ), .IN0(\CARRYB[78][1] ), .IN1(
        \SUMB[78][2] ), .COUT(\CARRYB[79][1] ), .SUM(\SUMB[79][1] ) );
  FADDER S3_79_2 ( .CIN(\ab[79][2] ), .IN0(\CARRYB[78][2] ), .IN1(\ab[78][3] ), 
        .COUT(\CARRYB[79][2] ), .SUM(\SUMB[79][2] ) );
  FADDER S1_78_0 ( .CIN(\ab[78][0] ), .IN0(\CARRYB[77][0] ), .IN1(
        \SUMB[77][1] ), .COUT(\CARRYB[78][0] ), .SUM(PRODUCT[78]) );
  FADDER S2_78_1 ( .CIN(\ab[78][1] ), .IN0(\CARRYB[77][1] ), .IN1(
        \SUMB[77][2] ), .COUT(\CARRYB[78][1] ), .SUM(\SUMB[78][1] ) );
  FADDER S3_78_2 ( .CIN(\ab[78][2] ), .IN0(\CARRYB[77][2] ), .IN1(\ab[77][3] ), 
        .COUT(\CARRYB[78][2] ), .SUM(\SUMB[78][2] ) );
  FADDER S1_77_0 ( .CIN(\ab[77][0] ), .IN0(\CARRYB[76][0] ), .IN1(
        \SUMB[76][1] ), .COUT(\CARRYB[77][0] ), .SUM(PRODUCT[77]) );
  FADDER S2_77_1 ( .CIN(\ab[77][1] ), .IN0(\CARRYB[76][1] ), .IN1(
        \SUMB[76][2] ), .COUT(\CARRYB[77][1] ), .SUM(\SUMB[77][1] ) );
  FADDER S3_77_2 ( .CIN(\ab[77][2] ), .IN0(\CARRYB[76][2] ), .IN1(\ab[76][3] ), 
        .COUT(\CARRYB[77][2] ), .SUM(\SUMB[77][2] ) );
  FADDER S1_76_0 ( .CIN(\ab[76][0] ), .IN0(\CARRYB[75][0] ), .IN1(
        \SUMB[75][1] ), .COUT(\CARRYB[76][0] ), .SUM(PRODUCT[76]) );
  FADDER S2_76_1 ( .CIN(\ab[76][1] ), .IN0(\CARRYB[75][1] ), .IN1(
        \SUMB[75][2] ), .COUT(\CARRYB[76][1] ), .SUM(\SUMB[76][1] ) );
  FADDER S3_76_2 ( .CIN(\ab[76][2] ), .IN0(\CARRYB[75][2] ), .IN1(\ab[75][3] ), 
        .COUT(\CARRYB[76][2] ), .SUM(\SUMB[76][2] ) );
  FADDER S1_75_0 ( .CIN(\ab[75][0] ), .IN0(\CARRYB[74][0] ), .IN1(
        \SUMB[74][1] ), .COUT(\CARRYB[75][0] ), .SUM(PRODUCT[75]) );
  FADDER S2_75_1 ( .CIN(\ab[75][1] ), .IN0(\CARRYB[74][1] ), .IN1(
        \SUMB[74][2] ), .COUT(\CARRYB[75][1] ), .SUM(\SUMB[75][1] ) );
  FADDER S3_75_2 ( .CIN(\ab[75][2] ), .IN0(\CARRYB[74][2] ), .IN1(\ab[74][3] ), 
        .COUT(\CARRYB[75][2] ), .SUM(\SUMB[75][2] ) );
  FADDER S1_74_0 ( .CIN(\ab[74][0] ), .IN0(\CARRYB[73][0] ), .IN1(
        \SUMB[73][1] ), .COUT(\CARRYB[74][0] ), .SUM(PRODUCT[74]) );
  FADDER S2_74_1 ( .CIN(\ab[74][1] ), .IN0(\CARRYB[73][1] ), .IN1(
        \SUMB[73][2] ), .COUT(\CARRYB[74][1] ), .SUM(\SUMB[74][1] ) );
  FADDER S3_74_2 ( .CIN(\ab[74][2] ), .IN0(\CARRYB[73][2] ), .IN1(\ab[73][3] ), 
        .COUT(\CARRYB[74][2] ), .SUM(\SUMB[74][2] ) );
  FADDER S1_73_0 ( .CIN(\ab[73][0] ), .IN0(\CARRYB[72][0] ), .IN1(
        \SUMB[72][1] ), .COUT(\CARRYB[73][0] ), .SUM(PRODUCT[73]) );
  FADDER S2_73_1 ( .CIN(\ab[73][1] ), .IN0(\CARRYB[72][1] ), .IN1(
        \SUMB[72][2] ), .COUT(\CARRYB[73][1] ), .SUM(\SUMB[73][1] ) );
  FADDER S3_73_2 ( .CIN(\ab[73][2] ), .IN0(\CARRYB[72][2] ), .IN1(\ab[72][3] ), 
        .COUT(\CARRYB[73][2] ), .SUM(\SUMB[73][2] ) );
  FADDER S1_72_0 ( .CIN(\ab[72][0] ), .IN0(\CARRYB[71][0] ), .IN1(
        \SUMB[71][1] ), .COUT(\CARRYB[72][0] ), .SUM(PRODUCT[72]) );
  FADDER S2_72_1 ( .CIN(\ab[72][1] ), .IN0(\CARRYB[71][1] ), .IN1(
        \SUMB[71][2] ), .COUT(\CARRYB[72][1] ), .SUM(\SUMB[72][1] ) );
  FADDER S3_72_2 ( .CIN(\ab[72][2] ), .IN0(\CARRYB[71][2] ), .IN1(\ab[71][3] ), 
        .COUT(\CARRYB[72][2] ), .SUM(\SUMB[72][2] ) );
  FADDER S1_71_0 ( .CIN(\ab[71][0] ), .IN0(\CARRYB[70][0] ), .IN1(
        \SUMB[70][1] ), .COUT(\CARRYB[71][0] ), .SUM(PRODUCT[71]) );
  FADDER S2_71_1 ( .CIN(\ab[71][1] ), .IN0(\CARRYB[70][1] ), .IN1(
        \SUMB[70][2] ), .COUT(\CARRYB[71][1] ), .SUM(\SUMB[71][1] ) );
  FADDER S3_71_2 ( .CIN(\ab[71][2] ), .IN0(\CARRYB[70][2] ), .IN1(\ab[70][3] ), 
        .COUT(\CARRYB[71][2] ), .SUM(\SUMB[71][2] ) );
  FADDER S1_70_0 ( .CIN(\ab[70][0] ), .IN0(\CARRYB[69][0] ), .IN1(
        \SUMB[69][1] ), .COUT(\CARRYB[70][0] ), .SUM(PRODUCT[70]) );
  FADDER S2_70_1 ( .CIN(\ab[70][1] ), .IN0(\CARRYB[69][1] ), .IN1(
        \SUMB[69][2] ), .COUT(\CARRYB[70][1] ), .SUM(\SUMB[70][1] ) );
  FADDER S3_70_2 ( .CIN(\ab[70][2] ), .IN0(\CARRYB[69][2] ), .IN1(\ab[69][3] ), 
        .COUT(\CARRYB[70][2] ), .SUM(\SUMB[70][2] ) );
  FADDER S1_69_0 ( .CIN(\ab[69][0] ), .IN0(\CARRYB[68][0] ), .IN1(
        \SUMB[68][1] ), .COUT(\CARRYB[69][0] ), .SUM(PRODUCT[69]) );
  FADDER S2_69_1 ( .CIN(\ab[69][1] ), .IN0(\CARRYB[68][1] ), .IN1(
        \SUMB[68][2] ), .COUT(\CARRYB[69][1] ), .SUM(\SUMB[69][1] ) );
  FADDER S3_69_2 ( .CIN(\ab[69][2] ), .IN0(\CARRYB[68][2] ), .IN1(\ab[68][3] ), 
        .COUT(\CARRYB[69][2] ), .SUM(\SUMB[69][2] ) );
  FADDER S1_68_0 ( .CIN(\ab[68][0] ), .IN0(\CARRYB[67][0] ), .IN1(
        \SUMB[67][1] ), .COUT(\CARRYB[68][0] ), .SUM(PRODUCT[68]) );
  FADDER S2_68_1 ( .CIN(\ab[68][1] ), .IN0(\CARRYB[67][1] ), .IN1(
        \SUMB[67][2] ), .COUT(\CARRYB[68][1] ), .SUM(\SUMB[68][1] ) );
  FADDER S3_68_2 ( .CIN(\ab[68][2] ), .IN0(\CARRYB[67][2] ), .IN1(\ab[67][3] ), 
        .COUT(\CARRYB[68][2] ), .SUM(\SUMB[68][2] ) );
  FADDER S1_67_0 ( .CIN(\ab[67][0] ), .IN0(\CARRYB[66][0] ), .IN1(
        \SUMB[66][1] ), .COUT(\CARRYB[67][0] ), .SUM(PRODUCT[67]) );
  FADDER S2_67_1 ( .CIN(\ab[67][1] ), .IN0(\CARRYB[66][1] ), .IN1(
        \SUMB[66][2] ), .COUT(\CARRYB[67][1] ), .SUM(\SUMB[67][1] ) );
  FADDER S3_67_2 ( .CIN(\ab[67][2] ), .IN0(\CARRYB[66][2] ), .IN1(\ab[66][3] ), 
        .COUT(\CARRYB[67][2] ), .SUM(\SUMB[67][2] ) );
  FADDER S1_66_0 ( .CIN(\ab[66][0] ), .IN0(\CARRYB[65][0] ), .IN1(
        \SUMB[65][1] ), .COUT(\CARRYB[66][0] ), .SUM(PRODUCT[66]) );
  FADDER S2_66_1 ( .CIN(\ab[66][1] ), .IN0(\CARRYB[65][1] ), .IN1(
        \SUMB[65][2] ), .COUT(\CARRYB[66][1] ), .SUM(\SUMB[66][1] ) );
  FADDER S3_66_2 ( .CIN(\ab[66][2] ), .IN0(\CARRYB[65][2] ), .IN1(\ab[65][3] ), 
        .COUT(\CARRYB[66][2] ), .SUM(\SUMB[66][2] ) );
  FADDER S1_65_0 ( .CIN(\ab[65][0] ), .IN0(\CARRYB[64][0] ), .IN1(
        \SUMB[64][1] ), .COUT(\CARRYB[65][0] ), .SUM(PRODUCT[65]) );
  FADDER S2_65_1 ( .CIN(\ab[65][1] ), .IN0(\CARRYB[64][1] ), .IN1(
        \SUMB[64][2] ), .COUT(\CARRYB[65][1] ), .SUM(\SUMB[65][1] ) );
  FADDER S3_65_2 ( .CIN(\ab[65][2] ), .IN0(\CARRYB[64][2] ), .IN1(\ab[64][3] ), 
        .COUT(\CARRYB[65][2] ), .SUM(\SUMB[65][2] ) );
  FADDER S1_64_0 ( .CIN(\ab[64][0] ), .IN0(\CARRYB[63][0] ), .IN1(
        \SUMB[63][1] ), .COUT(\CARRYB[64][0] ), .SUM(PRODUCT[64]) );
  FADDER S2_64_1 ( .CIN(\ab[64][1] ), .IN0(\CARRYB[63][1] ), .IN1(
        \SUMB[63][2] ), .COUT(\CARRYB[64][1] ), .SUM(\SUMB[64][1] ) );
  FADDER S3_64_2 ( .CIN(\ab[64][2] ), .IN0(\CARRYB[63][2] ), .IN1(\ab[63][3] ), 
        .COUT(\CARRYB[64][2] ), .SUM(\SUMB[64][2] ) );
  FADDER S1_63_0 ( .CIN(\ab[63][0] ), .IN0(\CARRYB[62][0] ), .IN1(
        \SUMB[62][1] ), .COUT(\CARRYB[63][0] ), .SUM(PRODUCT[63]) );
  FADDER S2_63_1 ( .CIN(\ab[63][1] ), .IN0(\CARRYB[62][1] ), .IN1(
        \SUMB[62][2] ), .COUT(\CARRYB[63][1] ), .SUM(\SUMB[63][1] ) );
  FADDER S3_63_2 ( .CIN(\ab[63][2] ), .IN0(\CARRYB[62][2] ), .IN1(\ab[62][3] ), 
        .COUT(\CARRYB[63][2] ), .SUM(\SUMB[63][2] ) );
  FADDER S1_62_0 ( .CIN(\ab[62][0] ), .IN0(\CARRYB[61][0] ), .IN1(
        \SUMB[61][1] ), .COUT(\CARRYB[62][0] ), .SUM(PRODUCT[62]) );
  FADDER S2_62_1 ( .CIN(\ab[62][1] ), .IN0(\CARRYB[61][1] ), .IN1(
        \SUMB[61][2] ), .COUT(\CARRYB[62][1] ), .SUM(\SUMB[62][1] ) );
  FADDER S3_62_2 ( .CIN(\ab[62][2] ), .IN0(\CARRYB[61][2] ), .IN1(\ab[61][3] ), 
        .COUT(\CARRYB[62][2] ), .SUM(\SUMB[62][2] ) );
  FADDER S1_61_0 ( .CIN(\ab[61][0] ), .IN0(\CARRYB[60][0] ), .IN1(
        \SUMB[60][1] ), .COUT(\CARRYB[61][0] ), .SUM(PRODUCT[61]) );
  FADDER S2_61_1 ( .CIN(\ab[61][1] ), .IN0(\CARRYB[60][1] ), .IN1(
        \SUMB[60][2] ), .COUT(\CARRYB[61][1] ), .SUM(\SUMB[61][1] ) );
  FADDER S3_61_2 ( .CIN(\ab[61][2] ), .IN0(\CARRYB[60][2] ), .IN1(\ab[60][3] ), 
        .COUT(\CARRYB[61][2] ), .SUM(\SUMB[61][2] ) );
  FADDER S1_60_0 ( .CIN(\ab[60][0] ), .IN0(\CARRYB[59][0] ), .IN1(
        \SUMB[59][1] ), .COUT(\CARRYB[60][0] ), .SUM(PRODUCT[60]) );
  FADDER S2_60_1 ( .CIN(\ab[60][1] ), .IN0(\CARRYB[59][1] ), .IN1(
        \SUMB[59][2] ), .COUT(\CARRYB[60][1] ), .SUM(\SUMB[60][1] ) );
  FADDER S3_60_2 ( .CIN(\ab[60][2] ), .IN0(\CARRYB[59][2] ), .IN1(\ab[59][3] ), 
        .COUT(\CARRYB[60][2] ), .SUM(\SUMB[60][2] ) );
  FADDER S1_59_0 ( .CIN(\ab[59][0] ), .IN0(\CARRYB[58][0] ), .IN1(
        \SUMB[58][1] ), .COUT(\CARRYB[59][0] ), .SUM(PRODUCT[59]) );
  FADDER S2_59_1 ( .CIN(\ab[59][1] ), .IN0(\CARRYB[58][1] ), .IN1(
        \SUMB[58][2] ), .COUT(\CARRYB[59][1] ), .SUM(\SUMB[59][1] ) );
  FADDER S3_59_2 ( .CIN(\ab[59][2] ), .IN0(\CARRYB[58][2] ), .IN1(\ab[58][3] ), 
        .COUT(\CARRYB[59][2] ), .SUM(\SUMB[59][2] ) );
  FADDER S1_58_0 ( .CIN(\ab[58][0] ), .IN0(\CARRYB[57][0] ), .IN1(
        \SUMB[57][1] ), .COUT(\CARRYB[58][0] ), .SUM(PRODUCT[58]) );
  FADDER S2_58_1 ( .CIN(\ab[58][1] ), .IN0(\CARRYB[57][1] ), .IN1(
        \SUMB[57][2] ), .COUT(\CARRYB[58][1] ), .SUM(\SUMB[58][1] ) );
  FADDER S3_58_2 ( .CIN(\ab[58][2] ), .IN0(\CARRYB[57][2] ), .IN1(\ab[57][3] ), 
        .COUT(\CARRYB[58][2] ), .SUM(\SUMB[58][2] ) );
  FADDER S1_57_0 ( .CIN(\ab[57][0] ), .IN0(\CARRYB[56][0] ), .IN1(
        \SUMB[56][1] ), .COUT(\CARRYB[57][0] ), .SUM(PRODUCT[57]) );
  FADDER S2_57_1 ( .CIN(\ab[57][1] ), .IN0(\CARRYB[56][1] ), .IN1(
        \SUMB[56][2] ), .COUT(\CARRYB[57][1] ), .SUM(\SUMB[57][1] ) );
  FADDER S3_57_2 ( .CIN(\ab[57][2] ), .IN0(\CARRYB[56][2] ), .IN1(\ab[56][3] ), 
        .COUT(\CARRYB[57][2] ), .SUM(\SUMB[57][2] ) );
  FADDER S1_56_0 ( .CIN(\ab[56][0] ), .IN0(\CARRYB[55][0] ), .IN1(
        \SUMB[55][1] ), .COUT(\CARRYB[56][0] ), .SUM(PRODUCT[56]) );
  FADDER S2_56_1 ( .CIN(\ab[56][1] ), .IN0(\CARRYB[55][1] ), .IN1(
        \SUMB[55][2] ), .COUT(\CARRYB[56][1] ), .SUM(\SUMB[56][1] ) );
  FADDER S3_56_2 ( .CIN(\ab[56][2] ), .IN0(\CARRYB[55][2] ), .IN1(\ab[55][3] ), 
        .COUT(\CARRYB[56][2] ), .SUM(\SUMB[56][2] ) );
  FADDER S1_55_0 ( .CIN(\ab[55][0] ), .IN0(\CARRYB[54][0] ), .IN1(
        \SUMB[54][1] ), .COUT(\CARRYB[55][0] ), .SUM(PRODUCT[55]) );
  FADDER S2_55_1 ( .CIN(\ab[55][1] ), .IN0(\CARRYB[54][1] ), .IN1(
        \SUMB[54][2] ), .COUT(\CARRYB[55][1] ), .SUM(\SUMB[55][1] ) );
  FADDER S3_55_2 ( .CIN(\ab[55][2] ), .IN0(\CARRYB[54][2] ), .IN1(\ab[54][3] ), 
        .COUT(\CARRYB[55][2] ), .SUM(\SUMB[55][2] ) );
  FADDER S1_54_0 ( .CIN(\ab[54][0] ), .IN0(\CARRYB[53][0] ), .IN1(
        \SUMB[53][1] ), .COUT(\CARRYB[54][0] ), .SUM(PRODUCT[54]) );
  FADDER S2_54_1 ( .CIN(\ab[54][1] ), .IN0(\CARRYB[53][1] ), .IN1(
        \SUMB[53][2] ), .COUT(\CARRYB[54][1] ), .SUM(\SUMB[54][1] ) );
  FADDER S3_54_2 ( .CIN(\ab[54][2] ), .IN0(\CARRYB[53][2] ), .IN1(\ab[53][3] ), 
        .COUT(\CARRYB[54][2] ), .SUM(\SUMB[54][2] ) );
  FADDER S1_53_0 ( .CIN(\ab[53][0] ), .IN0(\CARRYB[52][0] ), .IN1(
        \SUMB[52][1] ), .COUT(\CARRYB[53][0] ), .SUM(PRODUCT[53]) );
  FADDER S2_53_1 ( .CIN(\ab[53][1] ), .IN0(\CARRYB[52][1] ), .IN1(
        \SUMB[52][2] ), .COUT(\CARRYB[53][1] ), .SUM(\SUMB[53][1] ) );
  FADDER S3_53_2 ( .CIN(\ab[53][2] ), .IN0(\CARRYB[52][2] ), .IN1(\ab[52][3] ), 
        .COUT(\CARRYB[53][2] ), .SUM(\SUMB[53][2] ) );
  FADDER S1_52_0 ( .CIN(\ab[52][0] ), .IN0(\CARRYB[51][0] ), .IN1(
        \SUMB[51][1] ), .COUT(\CARRYB[52][0] ), .SUM(PRODUCT[52]) );
  FADDER S2_52_1 ( .CIN(\ab[52][1] ), .IN0(\CARRYB[51][1] ), .IN1(
        \SUMB[51][2] ), .COUT(\CARRYB[52][1] ), .SUM(\SUMB[52][1] ) );
  FADDER S3_52_2 ( .CIN(\ab[52][2] ), .IN0(\CARRYB[51][2] ), .IN1(\ab[51][3] ), 
        .COUT(\CARRYB[52][2] ), .SUM(\SUMB[52][2] ) );
  FADDER S1_51_0 ( .CIN(\ab[51][0] ), .IN0(\CARRYB[50][0] ), .IN1(
        \SUMB[50][1] ), .COUT(\CARRYB[51][0] ), .SUM(PRODUCT[51]) );
  FADDER S2_51_1 ( .CIN(\ab[51][1] ), .IN0(\CARRYB[50][1] ), .IN1(
        \SUMB[50][2] ), .COUT(\CARRYB[51][1] ), .SUM(\SUMB[51][1] ) );
  FADDER S3_51_2 ( .CIN(\ab[51][2] ), .IN0(\CARRYB[50][2] ), .IN1(\ab[50][3] ), 
        .COUT(\CARRYB[51][2] ), .SUM(\SUMB[51][2] ) );
  FADDER S1_50_0 ( .CIN(\ab[50][0] ), .IN0(\CARRYB[49][0] ), .IN1(
        \SUMB[49][1] ), .COUT(\CARRYB[50][0] ), .SUM(PRODUCT[50]) );
  FADDER S2_50_1 ( .CIN(\ab[50][1] ), .IN0(\CARRYB[49][1] ), .IN1(
        \SUMB[49][2] ), .COUT(\CARRYB[50][1] ), .SUM(\SUMB[50][1] ) );
  FADDER S3_50_2 ( .CIN(\ab[50][2] ), .IN0(\CARRYB[49][2] ), .IN1(\ab[49][3] ), 
        .COUT(\CARRYB[50][2] ), .SUM(\SUMB[50][2] ) );
  FADDER S1_49_0 ( .CIN(\ab[49][0] ), .IN0(\CARRYB[48][0] ), .IN1(
        \SUMB[48][1] ), .COUT(\CARRYB[49][0] ), .SUM(PRODUCT[49]) );
  FADDER S2_49_1 ( .CIN(\ab[49][1] ), .IN0(\CARRYB[48][1] ), .IN1(
        \SUMB[48][2] ), .COUT(\CARRYB[49][1] ), .SUM(\SUMB[49][1] ) );
  FADDER S3_49_2 ( .CIN(\ab[49][2] ), .IN0(\CARRYB[48][2] ), .IN1(\ab[48][3] ), 
        .COUT(\CARRYB[49][2] ), .SUM(\SUMB[49][2] ) );
  FADDER S1_48_0 ( .CIN(\ab[48][0] ), .IN0(\CARRYB[47][0] ), .IN1(
        \SUMB[47][1] ), .COUT(\CARRYB[48][0] ), .SUM(PRODUCT[48]) );
  FADDER S2_48_1 ( .CIN(\ab[48][1] ), .IN0(\CARRYB[47][1] ), .IN1(
        \SUMB[47][2] ), .COUT(\CARRYB[48][1] ), .SUM(\SUMB[48][1] ) );
  FADDER S3_48_2 ( .CIN(\ab[48][2] ), .IN0(\CARRYB[47][2] ), .IN1(\ab[47][3] ), 
        .COUT(\CARRYB[48][2] ), .SUM(\SUMB[48][2] ) );
  FADDER S1_47_0 ( .CIN(\ab[47][0] ), .IN0(\CARRYB[46][0] ), .IN1(
        \SUMB[46][1] ), .COUT(\CARRYB[47][0] ), .SUM(PRODUCT[47]) );
  FADDER S2_47_1 ( .CIN(\ab[47][1] ), .IN0(\CARRYB[46][1] ), .IN1(
        \SUMB[46][2] ), .COUT(\CARRYB[47][1] ), .SUM(\SUMB[47][1] ) );
  FADDER S3_47_2 ( .CIN(\ab[47][2] ), .IN0(\CARRYB[46][2] ), .IN1(\ab[46][3] ), 
        .COUT(\CARRYB[47][2] ), .SUM(\SUMB[47][2] ) );
  FADDER S1_46_0 ( .CIN(\ab[46][0] ), .IN0(\CARRYB[45][0] ), .IN1(
        \SUMB[45][1] ), .COUT(\CARRYB[46][0] ), .SUM(PRODUCT[46]) );
  FADDER S2_46_1 ( .CIN(\ab[46][1] ), .IN0(\CARRYB[45][1] ), .IN1(
        \SUMB[45][2] ), .COUT(\CARRYB[46][1] ), .SUM(\SUMB[46][1] ) );
  FADDER S3_46_2 ( .CIN(\ab[46][2] ), .IN0(\CARRYB[45][2] ), .IN1(\ab[45][3] ), 
        .COUT(\CARRYB[46][2] ), .SUM(\SUMB[46][2] ) );
  FADDER S1_45_0 ( .CIN(\ab[45][0] ), .IN0(\CARRYB[44][0] ), .IN1(
        \SUMB[44][1] ), .COUT(\CARRYB[45][0] ), .SUM(PRODUCT[45]) );
  FADDER S2_45_1 ( .CIN(\ab[45][1] ), .IN0(\CARRYB[44][1] ), .IN1(
        \SUMB[44][2] ), .COUT(\CARRYB[45][1] ), .SUM(\SUMB[45][1] ) );
  FADDER S3_45_2 ( .CIN(\ab[45][2] ), .IN0(\CARRYB[44][2] ), .IN1(\ab[44][3] ), 
        .COUT(\CARRYB[45][2] ), .SUM(\SUMB[45][2] ) );
  FADDER S1_44_0 ( .CIN(\ab[44][0] ), .IN0(\CARRYB[43][0] ), .IN1(
        \SUMB[43][1] ), .COUT(\CARRYB[44][0] ), .SUM(PRODUCT[44]) );
  FADDER S2_44_1 ( .CIN(\ab[44][1] ), .IN0(\CARRYB[43][1] ), .IN1(
        \SUMB[43][2] ), .COUT(\CARRYB[44][1] ), .SUM(\SUMB[44][1] ) );
  FADDER S3_44_2 ( .CIN(\ab[44][2] ), .IN0(\CARRYB[43][2] ), .IN1(\ab[43][3] ), 
        .COUT(\CARRYB[44][2] ), .SUM(\SUMB[44][2] ) );
  FADDER S1_43_0 ( .CIN(\ab[43][0] ), .IN0(\CARRYB[42][0] ), .IN1(
        \SUMB[42][1] ), .COUT(\CARRYB[43][0] ), .SUM(PRODUCT[43]) );
  FADDER S2_43_1 ( .CIN(\ab[43][1] ), .IN0(\CARRYB[42][1] ), .IN1(
        \SUMB[42][2] ), .COUT(\CARRYB[43][1] ), .SUM(\SUMB[43][1] ) );
  FADDER S3_43_2 ( .CIN(\ab[43][2] ), .IN0(\CARRYB[42][2] ), .IN1(\ab[42][3] ), 
        .COUT(\CARRYB[43][2] ), .SUM(\SUMB[43][2] ) );
  FADDER S1_42_0 ( .CIN(\ab[42][0] ), .IN0(\CARRYB[41][0] ), .IN1(
        \SUMB[41][1] ), .COUT(\CARRYB[42][0] ), .SUM(PRODUCT[42]) );
  FADDER S2_42_1 ( .CIN(\ab[42][1] ), .IN0(\CARRYB[41][1] ), .IN1(
        \SUMB[41][2] ), .COUT(\CARRYB[42][1] ), .SUM(\SUMB[42][1] ) );
  FADDER S3_42_2 ( .CIN(\ab[42][2] ), .IN0(\CARRYB[41][2] ), .IN1(\ab[41][3] ), 
        .COUT(\CARRYB[42][2] ), .SUM(\SUMB[42][2] ) );
  FADDER S1_41_0 ( .CIN(\ab[41][0] ), .IN0(\CARRYB[40][0] ), .IN1(
        \SUMB[40][1] ), .COUT(\CARRYB[41][0] ), .SUM(PRODUCT[41]) );
  FADDER S2_41_1 ( .CIN(\ab[41][1] ), .IN0(\CARRYB[40][1] ), .IN1(
        \SUMB[40][2] ), .COUT(\CARRYB[41][1] ), .SUM(\SUMB[41][1] ) );
  FADDER S3_41_2 ( .CIN(\ab[41][2] ), .IN0(\CARRYB[40][2] ), .IN1(\ab[40][3] ), 
        .COUT(\CARRYB[41][2] ), .SUM(\SUMB[41][2] ) );
  FADDER S1_40_0 ( .CIN(\ab[40][0] ), .IN0(\CARRYB[39][0] ), .IN1(
        \SUMB[39][1] ), .COUT(\CARRYB[40][0] ), .SUM(PRODUCT[40]) );
  FADDER S2_40_1 ( .CIN(\ab[40][1] ), .IN0(\CARRYB[39][1] ), .IN1(
        \SUMB[39][2] ), .COUT(\CARRYB[40][1] ), .SUM(\SUMB[40][1] ) );
  FADDER S3_40_2 ( .CIN(\ab[40][2] ), .IN0(\CARRYB[39][2] ), .IN1(\ab[39][3] ), 
        .COUT(\CARRYB[40][2] ), .SUM(\SUMB[40][2] ) );
  FADDER S1_39_0 ( .CIN(\ab[39][0] ), .IN0(\CARRYB[38][0] ), .IN1(
        \SUMB[38][1] ), .COUT(\CARRYB[39][0] ), .SUM(PRODUCT[39]) );
  FADDER S2_39_1 ( .CIN(\ab[39][1] ), .IN0(\CARRYB[38][1] ), .IN1(
        \SUMB[38][2] ), .COUT(\CARRYB[39][1] ), .SUM(\SUMB[39][1] ) );
  FADDER S3_39_2 ( .CIN(\ab[39][2] ), .IN0(\CARRYB[38][2] ), .IN1(\ab[38][3] ), 
        .COUT(\CARRYB[39][2] ), .SUM(\SUMB[39][2] ) );
  FADDER S1_38_0 ( .CIN(\ab[38][0] ), .IN0(\CARRYB[37][0] ), .IN1(
        \SUMB[37][1] ), .COUT(\CARRYB[38][0] ), .SUM(PRODUCT[38]) );
  FADDER S2_38_1 ( .CIN(\ab[38][1] ), .IN0(\CARRYB[37][1] ), .IN1(
        \SUMB[37][2] ), .COUT(\CARRYB[38][1] ), .SUM(\SUMB[38][1] ) );
  FADDER S3_38_2 ( .CIN(\ab[38][2] ), .IN0(\CARRYB[37][2] ), .IN1(\ab[37][3] ), 
        .COUT(\CARRYB[38][2] ), .SUM(\SUMB[38][2] ) );
  FADDER S1_37_0 ( .CIN(\ab[37][0] ), .IN0(\CARRYB[36][0] ), .IN1(
        \SUMB[36][1] ), .COUT(\CARRYB[37][0] ), .SUM(PRODUCT[37]) );
  FADDER S2_37_1 ( .CIN(\ab[37][1] ), .IN0(\CARRYB[36][1] ), .IN1(
        \SUMB[36][2] ), .COUT(\CARRYB[37][1] ), .SUM(\SUMB[37][1] ) );
  FADDER S3_37_2 ( .CIN(\ab[37][2] ), .IN0(\CARRYB[36][2] ), .IN1(\ab[36][3] ), 
        .COUT(\CARRYB[37][2] ), .SUM(\SUMB[37][2] ) );
  FADDER S1_36_0 ( .CIN(\ab[36][0] ), .IN0(\CARRYB[35][0] ), .IN1(
        \SUMB[35][1] ), .COUT(\CARRYB[36][0] ), .SUM(PRODUCT[36]) );
  FADDER S2_36_1 ( .CIN(\ab[36][1] ), .IN0(\CARRYB[35][1] ), .IN1(
        \SUMB[35][2] ), .COUT(\CARRYB[36][1] ), .SUM(\SUMB[36][1] ) );
  FADDER S3_36_2 ( .CIN(\ab[36][2] ), .IN0(\CARRYB[35][2] ), .IN1(\ab[35][3] ), 
        .COUT(\CARRYB[36][2] ), .SUM(\SUMB[36][2] ) );
  FADDER S1_35_0 ( .CIN(\ab[35][0] ), .IN0(\CARRYB[34][0] ), .IN1(
        \SUMB[34][1] ), .COUT(\CARRYB[35][0] ), .SUM(PRODUCT[35]) );
  FADDER S2_35_1 ( .CIN(\ab[35][1] ), .IN0(\CARRYB[34][1] ), .IN1(
        \SUMB[34][2] ), .COUT(\CARRYB[35][1] ), .SUM(\SUMB[35][1] ) );
  FADDER S3_35_2 ( .CIN(\ab[35][2] ), .IN0(\CARRYB[34][2] ), .IN1(\ab[34][3] ), 
        .COUT(\CARRYB[35][2] ), .SUM(\SUMB[35][2] ) );
  FADDER S1_34_0 ( .CIN(\ab[34][0] ), .IN0(\CARRYB[33][0] ), .IN1(
        \SUMB[33][1] ), .COUT(\CARRYB[34][0] ), .SUM(PRODUCT[34]) );
  FADDER S2_34_1 ( .CIN(\ab[34][1] ), .IN0(\CARRYB[33][1] ), .IN1(
        \SUMB[33][2] ), .COUT(\CARRYB[34][1] ), .SUM(\SUMB[34][1] ) );
  FADDER S3_34_2 ( .CIN(\ab[34][2] ), .IN0(\CARRYB[33][2] ), .IN1(\ab[33][3] ), 
        .COUT(\CARRYB[34][2] ), .SUM(\SUMB[34][2] ) );
  FADDER S1_33_0 ( .CIN(\ab[33][0] ), .IN0(\CARRYB[32][0] ), .IN1(
        \SUMB[32][1] ), .COUT(\CARRYB[33][0] ), .SUM(PRODUCT[33]) );
  FADDER S2_33_1 ( .CIN(\ab[33][1] ), .IN0(\CARRYB[32][1] ), .IN1(
        \SUMB[32][2] ), .COUT(\CARRYB[33][1] ), .SUM(\SUMB[33][1] ) );
  FADDER S3_33_2 ( .CIN(\ab[33][2] ), .IN0(\CARRYB[32][2] ), .IN1(\ab[32][3] ), 
        .COUT(\CARRYB[33][2] ), .SUM(\SUMB[33][2] ) );
  FADDER S1_32_0 ( .CIN(\ab[32][0] ), .IN0(\CARRYB[31][0] ), .IN1(
        \SUMB[31][1] ), .COUT(\CARRYB[32][0] ), .SUM(PRODUCT[32]) );
  FADDER S2_32_1 ( .CIN(\ab[32][1] ), .IN0(\CARRYB[31][1] ), .IN1(
        \SUMB[31][2] ), .COUT(\CARRYB[32][1] ), .SUM(\SUMB[32][1] ) );
  FADDER S3_32_2 ( .CIN(\ab[32][2] ), .IN0(\CARRYB[31][2] ), .IN1(\ab[31][3] ), 
        .COUT(\CARRYB[32][2] ), .SUM(\SUMB[32][2] ) );
  FADDER S1_31_0 ( .CIN(\ab[31][0] ), .IN0(\CARRYB[30][0] ), .IN1(
        \SUMB[30][1] ), .COUT(\CARRYB[31][0] ), .SUM(PRODUCT[31]) );
  FADDER S2_31_1 ( .CIN(\ab[31][1] ), .IN0(\CARRYB[30][1] ), .IN1(
        \SUMB[30][2] ), .COUT(\CARRYB[31][1] ), .SUM(\SUMB[31][1] ) );
  FADDER S3_31_2 ( .CIN(\ab[31][2] ), .IN0(\CARRYB[30][2] ), .IN1(\ab[30][3] ), 
        .COUT(\CARRYB[31][2] ), .SUM(\SUMB[31][2] ) );
  FADDER S1_30_0 ( .CIN(\ab[30][0] ), .IN0(\CARRYB[29][0] ), .IN1(
        \SUMB[29][1] ), .COUT(\CARRYB[30][0] ), .SUM(PRODUCT[30]) );
  FADDER S2_30_1 ( .CIN(\ab[30][1] ), .IN0(\CARRYB[29][1] ), .IN1(
        \SUMB[29][2] ), .COUT(\CARRYB[30][1] ), .SUM(\SUMB[30][1] ) );
  FADDER S3_30_2 ( .CIN(\ab[30][2] ), .IN0(\CARRYB[29][2] ), .IN1(\ab[29][3] ), 
        .COUT(\CARRYB[30][2] ), .SUM(\SUMB[30][2] ) );
  FADDER S1_29_0 ( .CIN(\ab[29][0] ), .IN0(\CARRYB[28][0] ), .IN1(
        \SUMB[28][1] ), .COUT(\CARRYB[29][0] ), .SUM(PRODUCT[29]) );
  FADDER S2_29_1 ( .CIN(\ab[29][1] ), .IN0(\CARRYB[28][1] ), .IN1(
        \SUMB[28][2] ), .COUT(\CARRYB[29][1] ), .SUM(\SUMB[29][1] ) );
  FADDER S3_29_2 ( .CIN(\ab[29][2] ), .IN0(\CARRYB[28][2] ), .IN1(\ab[28][3] ), 
        .COUT(\CARRYB[29][2] ), .SUM(\SUMB[29][2] ) );
  FADDER S1_28_0 ( .CIN(\ab[28][0] ), .IN0(\CARRYB[27][0] ), .IN1(
        \SUMB[27][1] ), .COUT(\CARRYB[28][0] ), .SUM(PRODUCT[28]) );
  FADDER S2_28_1 ( .CIN(\ab[28][1] ), .IN0(\CARRYB[27][1] ), .IN1(
        \SUMB[27][2] ), .COUT(\CARRYB[28][1] ), .SUM(\SUMB[28][1] ) );
  FADDER S3_28_2 ( .CIN(\ab[28][2] ), .IN0(\CARRYB[27][2] ), .IN1(\ab[27][3] ), 
        .COUT(\CARRYB[28][2] ), .SUM(\SUMB[28][2] ) );
  FADDER S1_27_0 ( .CIN(\ab[27][0] ), .IN0(\CARRYB[26][0] ), .IN1(
        \SUMB[26][1] ), .COUT(\CARRYB[27][0] ), .SUM(PRODUCT[27]) );
  FADDER S2_27_1 ( .CIN(\ab[27][1] ), .IN0(\CARRYB[26][1] ), .IN1(
        \SUMB[26][2] ), .COUT(\CARRYB[27][1] ), .SUM(\SUMB[27][1] ) );
  FADDER S3_27_2 ( .CIN(\ab[27][2] ), .IN0(\CARRYB[26][2] ), .IN1(\ab[26][3] ), 
        .COUT(\CARRYB[27][2] ), .SUM(\SUMB[27][2] ) );
  FADDER S1_26_0 ( .CIN(\ab[26][0] ), .IN0(\CARRYB[25][0] ), .IN1(
        \SUMB[25][1] ), .COUT(\CARRYB[26][0] ), .SUM(PRODUCT[26]) );
  FADDER S2_26_1 ( .CIN(\ab[26][1] ), .IN0(\CARRYB[25][1] ), .IN1(
        \SUMB[25][2] ), .COUT(\CARRYB[26][1] ), .SUM(\SUMB[26][1] ) );
  FADDER S3_26_2 ( .CIN(\ab[26][2] ), .IN0(\CARRYB[25][2] ), .IN1(\ab[25][3] ), 
        .COUT(\CARRYB[26][2] ), .SUM(\SUMB[26][2] ) );
  FADDER S1_25_0 ( .CIN(\ab[25][0] ), .IN0(\CARRYB[24][0] ), .IN1(
        \SUMB[24][1] ), .COUT(\CARRYB[25][0] ), .SUM(PRODUCT[25]) );
  FADDER S2_25_1 ( .CIN(\ab[25][1] ), .IN0(\CARRYB[24][1] ), .IN1(
        \SUMB[24][2] ), .COUT(\CARRYB[25][1] ), .SUM(\SUMB[25][1] ) );
  FADDER S3_25_2 ( .CIN(\ab[25][2] ), .IN0(\CARRYB[24][2] ), .IN1(\ab[24][3] ), 
        .COUT(\CARRYB[25][2] ), .SUM(\SUMB[25][2] ) );
  FADDER S1_24_0 ( .CIN(\ab[24][0] ), .IN0(\CARRYB[23][0] ), .IN1(
        \SUMB[23][1] ), .COUT(\CARRYB[24][0] ), .SUM(PRODUCT[24]) );
  FADDER S2_24_1 ( .CIN(\ab[24][1] ), .IN0(\CARRYB[23][1] ), .IN1(
        \SUMB[23][2] ), .COUT(\CARRYB[24][1] ), .SUM(\SUMB[24][1] ) );
  FADDER S3_24_2 ( .CIN(\ab[24][2] ), .IN0(\CARRYB[23][2] ), .IN1(\ab[23][3] ), 
        .COUT(\CARRYB[24][2] ), .SUM(\SUMB[24][2] ) );
  FADDER S1_23_0 ( .CIN(\ab[23][0] ), .IN0(\CARRYB[22][0] ), .IN1(
        \SUMB[22][1] ), .COUT(\CARRYB[23][0] ), .SUM(PRODUCT[23]) );
  FADDER S2_23_1 ( .CIN(\ab[23][1] ), .IN0(\CARRYB[22][1] ), .IN1(
        \SUMB[22][2] ), .COUT(\CARRYB[23][1] ), .SUM(\SUMB[23][1] ) );
  FADDER S3_23_2 ( .CIN(\ab[23][2] ), .IN0(\CARRYB[22][2] ), .IN1(\ab[22][3] ), 
        .COUT(\CARRYB[23][2] ), .SUM(\SUMB[23][2] ) );
  FADDER S1_22_0 ( .CIN(\ab[22][0] ), .IN0(\CARRYB[21][0] ), .IN1(
        \SUMB[21][1] ), .COUT(\CARRYB[22][0] ), .SUM(PRODUCT[22]) );
  FADDER S2_22_1 ( .CIN(\ab[22][1] ), .IN0(\CARRYB[21][1] ), .IN1(
        \SUMB[21][2] ), .COUT(\CARRYB[22][1] ), .SUM(\SUMB[22][1] ) );
  FADDER S3_22_2 ( .CIN(\ab[22][2] ), .IN0(\CARRYB[21][2] ), .IN1(\ab[21][3] ), 
        .COUT(\CARRYB[22][2] ), .SUM(\SUMB[22][2] ) );
  FADDER S1_21_0 ( .CIN(\ab[21][0] ), .IN0(\CARRYB[20][0] ), .IN1(
        \SUMB[20][1] ), .COUT(\CARRYB[21][0] ), .SUM(PRODUCT[21]) );
  FADDER S2_21_1 ( .CIN(\ab[21][1] ), .IN0(\CARRYB[20][1] ), .IN1(
        \SUMB[20][2] ), .COUT(\CARRYB[21][1] ), .SUM(\SUMB[21][1] ) );
  FADDER S3_21_2 ( .CIN(\ab[21][2] ), .IN0(\CARRYB[20][2] ), .IN1(\ab[20][3] ), 
        .COUT(\CARRYB[21][2] ), .SUM(\SUMB[21][2] ) );
  FADDER S1_20_0 ( .CIN(\ab[20][0] ), .IN0(\CARRYB[19][0] ), .IN1(
        \SUMB[19][1] ), .COUT(\CARRYB[20][0] ), .SUM(PRODUCT[20]) );
  FADDER S2_20_1 ( .CIN(\ab[20][1] ), .IN0(\CARRYB[19][1] ), .IN1(
        \SUMB[19][2] ), .COUT(\CARRYB[20][1] ), .SUM(\SUMB[20][1] ) );
  FADDER S3_20_2 ( .CIN(\ab[20][2] ), .IN0(\CARRYB[19][2] ), .IN1(\ab[19][3] ), 
        .COUT(\CARRYB[20][2] ), .SUM(\SUMB[20][2] ) );
  FADDER S1_19_0 ( .CIN(\ab[19][0] ), .IN0(\CARRYB[18][0] ), .IN1(
        \SUMB[18][1] ), .COUT(\CARRYB[19][0] ), .SUM(PRODUCT[19]) );
  FADDER S2_19_1 ( .CIN(\ab[19][1] ), .IN0(\CARRYB[18][1] ), .IN1(
        \SUMB[18][2] ), .COUT(\CARRYB[19][1] ), .SUM(\SUMB[19][1] ) );
  FADDER S3_19_2 ( .CIN(\ab[19][2] ), .IN0(\CARRYB[18][2] ), .IN1(\ab[18][3] ), 
        .COUT(\CARRYB[19][2] ), .SUM(\SUMB[19][2] ) );
  FADDER S1_18_0 ( .CIN(\ab[18][0] ), .IN0(\CARRYB[17][0] ), .IN1(
        \SUMB[17][1] ), .COUT(\CARRYB[18][0] ), .SUM(PRODUCT[18]) );
  FADDER S2_18_1 ( .CIN(\ab[18][1] ), .IN0(\CARRYB[17][1] ), .IN1(
        \SUMB[17][2] ), .COUT(\CARRYB[18][1] ), .SUM(\SUMB[18][1] ) );
  FADDER S3_18_2 ( .CIN(\ab[18][2] ), .IN0(\CARRYB[17][2] ), .IN1(\ab[17][3] ), 
        .COUT(\CARRYB[18][2] ), .SUM(\SUMB[18][2] ) );
  FADDER S1_17_0 ( .CIN(\ab[17][0] ), .IN0(\CARRYB[16][0] ), .IN1(
        \SUMB[16][1] ), .COUT(\CARRYB[17][0] ), .SUM(PRODUCT[17]) );
  FADDER S2_17_1 ( .CIN(\ab[17][1] ), .IN0(\CARRYB[16][1] ), .IN1(
        \SUMB[16][2] ), .COUT(\CARRYB[17][1] ), .SUM(\SUMB[17][1] ) );
  FADDER S3_17_2 ( .CIN(\ab[17][2] ), .IN0(\CARRYB[16][2] ), .IN1(\ab[16][3] ), 
        .COUT(\CARRYB[17][2] ), .SUM(\SUMB[17][2] ) );
  FADDER S1_16_0 ( .CIN(\ab[16][0] ), .IN0(\CARRYB[15][0] ), .IN1(
        \SUMB[15][1] ), .COUT(\CARRYB[16][0] ), .SUM(PRODUCT[16]) );
  FADDER S2_16_1 ( .CIN(\ab[16][1] ), .IN0(\CARRYB[15][1] ), .IN1(
        \SUMB[15][2] ), .COUT(\CARRYB[16][1] ), .SUM(\SUMB[16][1] ) );
  FADDER S3_16_2 ( .CIN(\ab[16][2] ), .IN0(\CARRYB[15][2] ), .IN1(\ab[15][3] ), 
        .COUT(\CARRYB[16][2] ), .SUM(\SUMB[16][2] ) );
  FADDER S1_15_0 ( .CIN(\ab[15][0] ), .IN0(\CARRYB[14][0] ), .IN1(
        \SUMB[14][1] ), .COUT(\CARRYB[15][0] ), .SUM(PRODUCT[15]) );
  FADDER S2_15_1 ( .CIN(\ab[15][1] ), .IN0(\CARRYB[14][1] ), .IN1(
        \SUMB[14][2] ), .COUT(\CARRYB[15][1] ), .SUM(\SUMB[15][1] ) );
  FADDER S3_15_2 ( .CIN(\ab[15][2] ), .IN0(\CARRYB[14][2] ), .IN1(\ab[14][3] ), 
        .COUT(\CARRYB[15][2] ), .SUM(\SUMB[15][2] ) );
  FADDER S1_14_0 ( .CIN(\ab[14][0] ), .IN0(\CARRYB[13][0] ), .IN1(
        \SUMB[13][1] ), .COUT(\CARRYB[14][0] ), .SUM(PRODUCT[14]) );
  FADDER S2_14_1 ( .CIN(\ab[14][1] ), .IN0(\CARRYB[13][1] ), .IN1(
        \SUMB[13][2] ), .COUT(\CARRYB[14][1] ), .SUM(\SUMB[14][1] ) );
  FADDER S3_14_2 ( .CIN(\ab[14][2] ), .IN0(\CARRYB[13][2] ), .IN1(\ab[13][3] ), 
        .COUT(\CARRYB[14][2] ), .SUM(\SUMB[14][2] ) );
  FADDER S1_13_0 ( .CIN(\ab[13][0] ), .IN0(\CARRYB[12][0] ), .IN1(
        \SUMB[12][1] ), .COUT(\CARRYB[13][0] ), .SUM(PRODUCT[13]) );
  FADDER S2_13_1 ( .CIN(\ab[13][1] ), .IN0(\CARRYB[12][1] ), .IN1(
        \SUMB[12][2] ), .COUT(\CARRYB[13][1] ), .SUM(\SUMB[13][1] ) );
  FADDER S3_13_2 ( .CIN(\ab[13][2] ), .IN0(\CARRYB[12][2] ), .IN1(\ab[12][3] ), 
        .COUT(\CARRYB[13][2] ), .SUM(\SUMB[13][2] ) );
  FADDER S1_12_0 ( .CIN(\ab[12][0] ), .IN0(\CARRYB[11][0] ), .IN1(
        \SUMB[11][1] ), .COUT(\CARRYB[12][0] ), .SUM(PRODUCT[12]) );
  FADDER S2_12_1 ( .CIN(\ab[12][1] ), .IN0(\CARRYB[11][1] ), .IN1(
        \SUMB[11][2] ), .COUT(\CARRYB[12][1] ), .SUM(\SUMB[12][1] ) );
  FADDER S3_12_2 ( .CIN(\ab[12][2] ), .IN0(\CARRYB[11][2] ), .IN1(\ab[11][3] ), 
        .COUT(\CARRYB[12][2] ), .SUM(\SUMB[12][2] ) );
  FADDER S1_11_0 ( .CIN(\ab[11][0] ), .IN0(\CARRYB[10][0] ), .IN1(
        \SUMB[10][1] ), .COUT(\CARRYB[11][0] ), .SUM(PRODUCT[11]) );
  FADDER S2_11_1 ( .CIN(\ab[11][1] ), .IN0(\CARRYB[10][1] ), .IN1(
        \SUMB[10][2] ), .COUT(\CARRYB[11][1] ), .SUM(\SUMB[11][1] ) );
  FADDER S3_11_2 ( .CIN(\ab[11][2] ), .IN0(\CARRYB[10][2] ), .IN1(\ab[10][3] ), 
        .COUT(\CARRYB[11][2] ), .SUM(\SUMB[11][2] ) );
  FADDER S1_10_0 ( .CIN(\ab[10][0] ), .IN0(\CARRYB[9][0] ), .IN1(\SUMB[9][1] ), 
        .COUT(\CARRYB[10][0] ), .SUM(PRODUCT[10]) );
  FADDER S2_10_1 ( .CIN(\ab[10][1] ), .IN0(\CARRYB[9][1] ), .IN1(\SUMB[9][2] ), 
        .COUT(\CARRYB[10][1] ), .SUM(\SUMB[10][1] ) );
  FADDER S3_10_2 ( .CIN(\ab[10][2] ), .IN0(\CARRYB[9][2] ), .IN1(\ab[9][3] ), 
        .COUT(\CARRYB[10][2] ), .SUM(\SUMB[10][2] ) );
  FADDER S1_9_0 ( .CIN(\ab[9][0] ), .IN0(\CARRYB[8][0] ), .IN1(\SUMB[8][1] ), 
        .COUT(\CARRYB[9][0] ), .SUM(PRODUCT[9]) );
  FADDER S2_9_1 ( .CIN(\ab[9][1] ), .IN0(\CARRYB[8][1] ), .IN1(\SUMB[8][2] ), 
        .COUT(\CARRYB[9][1] ), .SUM(\SUMB[9][1] ) );
  FADDER S3_9_2 ( .CIN(\ab[9][2] ), .IN0(\CARRYB[8][2] ), .IN1(\ab[8][3] ), 
        .COUT(\CARRYB[9][2] ), .SUM(\SUMB[9][2] ) );
  FADDER S1_8_0 ( .CIN(\ab[8][0] ), .IN0(\CARRYB[7][0] ), .IN1(\SUMB[7][1] ), 
        .COUT(\CARRYB[8][0] ), .SUM(PRODUCT[8]) );
  FADDER S2_8_1 ( .CIN(\ab[8][1] ), .IN0(\CARRYB[7][1] ), .IN1(\SUMB[7][2] ), 
        .COUT(\CARRYB[8][1] ), .SUM(\SUMB[8][1] ) );
  FADDER S3_8_2 ( .CIN(\ab[8][2] ), .IN0(\CARRYB[7][2] ), .IN1(\ab[7][3] ), 
        .COUT(\CARRYB[8][2] ), .SUM(\SUMB[8][2] ) );
  FADDER S1_7_0 ( .CIN(\ab[7][0] ), .IN0(\CARRYB[6][0] ), .IN1(\SUMB[6][1] ), 
        .COUT(\CARRYB[7][0] ), .SUM(PRODUCT[7]) );
  FADDER S2_7_1 ( .CIN(\ab[7][1] ), .IN0(\CARRYB[6][1] ), .IN1(\SUMB[6][2] ), 
        .COUT(\CARRYB[7][1] ), .SUM(\SUMB[7][1] ) );
  FADDER S3_7_2 ( .CIN(\ab[7][2] ), .IN0(\CARRYB[6][2] ), .IN1(\ab[6][3] ), 
        .COUT(\CARRYB[7][2] ), .SUM(\SUMB[7][2] ) );
  FADDER S1_6_0 ( .CIN(\ab[6][0] ), .IN0(\CARRYB[5][0] ), .IN1(\SUMB[5][1] ), 
        .COUT(\CARRYB[6][0] ), .SUM(PRODUCT[6]) );
  FADDER S2_6_1 ( .CIN(\ab[6][1] ), .IN0(\CARRYB[5][1] ), .IN1(\SUMB[5][2] ), 
        .COUT(\CARRYB[6][1] ), .SUM(\SUMB[6][1] ) );
  FADDER S3_6_2 ( .CIN(\ab[6][2] ), .IN0(\CARRYB[5][2] ), .IN1(\ab[5][3] ), 
        .COUT(\CARRYB[6][2] ), .SUM(\SUMB[6][2] ) );
  FADDER S1_5_0 ( .CIN(\ab[5][0] ), .IN0(\CARRYB[4][0] ), .IN1(\SUMB[4][1] ), 
        .COUT(\CARRYB[5][0] ), .SUM(PRODUCT[5]) );
  FADDER S2_5_1 ( .CIN(\ab[5][1] ), .IN0(\CARRYB[4][1] ), .IN1(\SUMB[4][2] ), 
        .COUT(\CARRYB[5][1] ), .SUM(\SUMB[5][1] ) );
  FADDER S3_5_2 ( .CIN(\ab[5][2] ), .IN0(\CARRYB[4][2] ), .IN1(\ab[4][3] ), 
        .COUT(\CARRYB[5][2] ), .SUM(\SUMB[5][2] ) );
  FADDER S1_4_0 ( .CIN(\ab[4][0] ), .IN0(\CARRYB[3][0] ), .IN1(\SUMB[3][1] ), 
        .COUT(\CARRYB[4][0] ), .SUM(PRODUCT[4]) );
  FADDER S2_4_1 ( .CIN(\ab[4][1] ), .IN0(\CARRYB[3][1] ), .IN1(\SUMB[3][2] ), 
        .COUT(\CARRYB[4][1] ), .SUM(\SUMB[4][1] ) );
  FADDER S3_4_2 ( .CIN(\ab[4][2] ), .IN0(\CARRYB[3][2] ), .IN1(\ab[3][3] ), 
        .COUT(\CARRYB[4][2] ), .SUM(\SUMB[4][2] ) );
  FADDER S1_3_0 ( .CIN(\ab[3][0] ), .IN0(\CARRYB[2][0] ), .IN1(\SUMB[2][1] ), 
        .COUT(\CARRYB[3][0] ), .SUM(PRODUCT[3]) );
  FADDER S2_3_1 ( .CIN(\ab[3][1] ), .IN0(\CARRYB[2][1] ), .IN1(\SUMB[2][2] ), 
        .COUT(\CARRYB[3][1] ), .SUM(\SUMB[3][1] ) );
  FADDER S3_3_2 ( .CIN(\ab[3][2] ), .IN0(\CARRYB[2][2] ), .IN1(\ab[2][3] ), 
        .COUT(\CARRYB[3][2] ), .SUM(\SUMB[3][2] ) );
  FADDER S1_2_0 ( .CIN(\ab[2][0] ), .IN0(\CARRYB[1][0] ), .IN1(\SUMB[1][1] ), 
        .COUT(\CARRYB[2][0] ), .SUM(PRODUCT[2]) );
  FADDER S2_2_1 ( .CIN(\ab[2][1] ), .IN0(\CARRYB[1][1] ), .IN1(\SUMB[1][2] ), 
        .COUT(\CARRYB[2][1] ), .SUM(\SUMB[2][1] ) );
  FADDER S3_2_2 ( .CIN(\ab[2][2] ), .IN0(\CARRYB[1][2] ), .IN1(\ab[1][3] ), 
        .COUT(\CARRYB[2][2] ), .SUM(\SUMB[2][2] ) );
  AND U2 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(\CARRYB[1][0] ) );
  XOR U3 ( .A(\ab[0][1] ), .B(\ab[1][0] ), .Z(PRODUCT[1]) );
  AND U4 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\CARRYB[1][1] ) );
  XOR U5 ( .A(\ab[0][2] ), .B(\ab[1][1] ), .Z(\SUMB[1][1] ) );
  AND U6 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\CARRYB[1][2] ) );
  XOR U7 ( .A(\ab[0][3] ), .B(\ab[1][2] ), .Z(\SUMB[1][2] ) );
  AND U8 ( .A(A[9]), .B(B[3]), .Z(\ab[9][3] ) );
  AND U9 ( .A(A[9]), .B(B[2]), .Z(\ab[9][2] ) );
  AND U10 ( .A(A[9]), .B(B[1]), .Z(\ab[9][1] ) );
  AND U11 ( .A(A[9]), .B(B[0]), .Z(\ab[9][0] ) );
  AND U12 ( .A(B[3]), .B(A[99]), .Z(\ab[99][3] ) );
  AND U13 ( .A(B[2]), .B(A[99]), .Z(\ab[99][2] ) );
  AND U14 ( .A(B[1]), .B(A[99]), .Z(\ab[99][1] ) );
  AND U15 ( .A(A[99]), .B(B[0]), .Z(\ab[99][0] ) );
  AND U16 ( .A(B[3]), .B(A[999]), .Z(\ab[999][3] ) );
  AND U17 ( .A(B[2]), .B(A[999]), .Z(\ab[999][2] ) );
  AND U18 ( .A(B[1]), .B(A[999]), .Z(\ab[999][1] ) );
  AND U19 ( .A(A[999]), .B(B[0]), .Z(\ab[999][0] ) );
  AND U20 ( .A(B[3]), .B(A[998]), .Z(\ab[998][3] ) );
  AND U21 ( .A(B[2]), .B(A[998]), .Z(\ab[998][2] ) );
  AND U22 ( .A(B[1]), .B(A[998]), .Z(\ab[998][1] ) );
  AND U23 ( .A(A[998]), .B(B[0]), .Z(\ab[998][0] ) );
  AND U24 ( .A(B[3]), .B(A[997]), .Z(\ab[997][3] ) );
  AND U25 ( .A(B[2]), .B(A[997]), .Z(\ab[997][2] ) );
  AND U26 ( .A(B[1]), .B(A[997]), .Z(\ab[997][1] ) );
  AND U27 ( .A(A[997]), .B(B[0]), .Z(\ab[997][0] ) );
  AND U28 ( .A(B[3]), .B(A[996]), .Z(\ab[996][3] ) );
  AND U29 ( .A(B[2]), .B(A[996]), .Z(\ab[996][2] ) );
  AND U30 ( .A(B[1]), .B(A[996]), .Z(\ab[996][1] ) );
  AND U31 ( .A(A[996]), .B(B[0]), .Z(\ab[996][0] ) );
  AND U32 ( .A(B[3]), .B(A[995]), .Z(\ab[995][3] ) );
  AND U33 ( .A(B[2]), .B(A[995]), .Z(\ab[995][2] ) );
  AND U34 ( .A(B[1]), .B(A[995]), .Z(\ab[995][1] ) );
  AND U35 ( .A(A[995]), .B(B[0]), .Z(\ab[995][0] ) );
  AND U36 ( .A(B[3]), .B(A[994]), .Z(\ab[994][3] ) );
  AND U37 ( .A(B[2]), .B(A[994]), .Z(\ab[994][2] ) );
  AND U38 ( .A(B[1]), .B(A[994]), .Z(\ab[994][1] ) );
  AND U39 ( .A(A[994]), .B(B[0]), .Z(\ab[994][0] ) );
  AND U40 ( .A(B[3]), .B(A[993]), .Z(\ab[993][3] ) );
  AND U41 ( .A(B[2]), .B(A[993]), .Z(\ab[993][2] ) );
  AND U42 ( .A(B[1]), .B(A[993]), .Z(\ab[993][1] ) );
  AND U43 ( .A(A[993]), .B(B[0]), .Z(\ab[993][0] ) );
  AND U44 ( .A(B[3]), .B(A[992]), .Z(\ab[992][3] ) );
  AND U45 ( .A(B[2]), .B(A[992]), .Z(\ab[992][2] ) );
  AND U46 ( .A(B[1]), .B(A[992]), .Z(\ab[992][1] ) );
  AND U47 ( .A(A[992]), .B(B[0]), .Z(\ab[992][0] ) );
  AND U48 ( .A(B[3]), .B(A[991]), .Z(\ab[991][3] ) );
  AND U49 ( .A(B[2]), .B(A[991]), .Z(\ab[991][2] ) );
  AND U50 ( .A(B[1]), .B(A[991]), .Z(\ab[991][1] ) );
  AND U51 ( .A(A[991]), .B(B[0]), .Z(\ab[991][0] ) );
  AND U52 ( .A(B[3]), .B(A[990]), .Z(\ab[990][3] ) );
  AND U53 ( .A(B[2]), .B(A[990]), .Z(\ab[990][2] ) );
  AND U54 ( .A(B[1]), .B(A[990]), .Z(\ab[990][1] ) );
  AND U55 ( .A(A[990]), .B(B[0]), .Z(\ab[990][0] ) );
  AND U56 ( .A(B[3]), .B(A[98]), .Z(\ab[98][3] ) );
  AND U57 ( .A(B[2]), .B(A[98]), .Z(\ab[98][2] ) );
  AND U58 ( .A(B[1]), .B(A[98]), .Z(\ab[98][1] ) );
  AND U59 ( .A(A[98]), .B(B[0]), .Z(\ab[98][0] ) );
  AND U60 ( .A(B[3]), .B(A[989]), .Z(\ab[989][3] ) );
  AND U61 ( .A(B[2]), .B(A[989]), .Z(\ab[989][2] ) );
  AND U62 ( .A(B[1]), .B(A[989]), .Z(\ab[989][1] ) );
  AND U63 ( .A(A[989]), .B(B[0]), .Z(\ab[989][0] ) );
  AND U64 ( .A(B[3]), .B(A[988]), .Z(\ab[988][3] ) );
  AND U65 ( .A(B[2]), .B(A[988]), .Z(\ab[988][2] ) );
  AND U66 ( .A(B[1]), .B(A[988]), .Z(\ab[988][1] ) );
  AND U67 ( .A(A[988]), .B(B[0]), .Z(\ab[988][0] ) );
  AND U68 ( .A(B[3]), .B(A[987]), .Z(\ab[987][3] ) );
  AND U69 ( .A(B[2]), .B(A[987]), .Z(\ab[987][2] ) );
  AND U70 ( .A(B[1]), .B(A[987]), .Z(\ab[987][1] ) );
  AND U71 ( .A(A[987]), .B(B[0]), .Z(\ab[987][0] ) );
  AND U72 ( .A(B[3]), .B(A[986]), .Z(\ab[986][3] ) );
  AND U73 ( .A(B[2]), .B(A[986]), .Z(\ab[986][2] ) );
  AND U74 ( .A(B[1]), .B(A[986]), .Z(\ab[986][1] ) );
  AND U75 ( .A(A[986]), .B(B[0]), .Z(\ab[986][0] ) );
  AND U76 ( .A(B[3]), .B(A[985]), .Z(\ab[985][3] ) );
  AND U77 ( .A(B[2]), .B(A[985]), .Z(\ab[985][2] ) );
  AND U78 ( .A(B[1]), .B(A[985]), .Z(\ab[985][1] ) );
  AND U79 ( .A(A[985]), .B(B[0]), .Z(\ab[985][0] ) );
  AND U80 ( .A(B[3]), .B(A[984]), .Z(\ab[984][3] ) );
  AND U81 ( .A(B[2]), .B(A[984]), .Z(\ab[984][2] ) );
  AND U82 ( .A(B[1]), .B(A[984]), .Z(\ab[984][1] ) );
  AND U83 ( .A(A[984]), .B(B[0]), .Z(\ab[984][0] ) );
  AND U84 ( .A(B[3]), .B(A[983]), .Z(\ab[983][3] ) );
  AND U85 ( .A(B[2]), .B(A[983]), .Z(\ab[983][2] ) );
  AND U86 ( .A(B[1]), .B(A[983]), .Z(\ab[983][1] ) );
  AND U87 ( .A(A[983]), .B(B[0]), .Z(\ab[983][0] ) );
  AND U88 ( .A(B[3]), .B(A[982]), .Z(\ab[982][3] ) );
  AND U89 ( .A(B[2]), .B(A[982]), .Z(\ab[982][2] ) );
  AND U90 ( .A(B[1]), .B(A[982]), .Z(\ab[982][1] ) );
  AND U91 ( .A(A[982]), .B(B[0]), .Z(\ab[982][0] ) );
  AND U92 ( .A(B[3]), .B(A[981]), .Z(\ab[981][3] ) );
  AND U93 ( .A(B[2]), .B(A[981]), .Z(\ab[981][2] ) );
  AND U94 ( .A(B[1]), .B(A[981]), .Z(\ab[981][1] ) );
  AND U95 ( .A(A[981]), .B(B[0]), .Z(\ab[981][0] ) );
  AND U96 ( .A(B[3]), .B(A[980]), .Z(\ab[980][3] ) );
  AND U97 ( .A(B[2]), .B(A[980]), .Z(\ab[980][2] ) );
  AND U98 ( .A(B[1]), .B(A[980]), .Z(\ab[980][1] ) );
  AND U99 ( .A(A[980]), .B(B[0]), .Z(\ab[980][0] ) );
  AND U100 ( .A(B[3]), .B(A[97]), .Z(\ab[97][3] ) );
  AND U101 ( .A(B[2]), .B(A[97]), .Z(\ab[97][2] ) );
  AND U102 ( .A(B[1]), .B(A[97]), .Z(\ab[97][1] ) );
  AND U103 ( .A(A[97]), .B(B[0]), .Z(\ab[97][0] ) );
  AND U104 ( .A(B[3]), .B(A[979]), .Z(\ab[979][3] ) );
  AND U105 ( .A(B[2]), .B(A[979]), .Z(\ab[979][2] ) );
  AND U106 ( .A(B[1]), .B(A[979]), .Z(\ab[979][1] ) );
  AND U107 ( .A(A[979]), .B(B[0]), .Z(\ab[979][0] ) );
  AND U108 ( .A(B[3]), .B(A[978]), .Z(\ab[978][3] ) );
  AND U109 ( .A(B[2]), .B(A[978]), .Z(\ab[978][2] ) );
  AND U110 ( .A(B[1]), .B(A[978]), .Z(\ab[978][1] ) );
  AND U111 ( .A(A[978]), .B(B[0]), .Z(\ab[978][0] ) );
  AND U112 ( .A(B[3]), .B(A[977]), .Z(\ab[977][3] ) );
  AND U113 ( .A(B[2]), .B(A[977]), .Z(\ab[977][2] ) );
  AND U114 ( .A(B[1]), .B(A[977]), .Z(\ab[977][1] ) );
  AND U115 ( .A(A[977]), .B(B[0]), .Z(\ab[977][0] ) );
  AND U116 ( .A(B[3]), .B(A[976]), .Z(\ab[976][3] ) );
  AND U117 ( .A(B[2]), .B(A[976]), .Z(\ab[976][2] ) );
  AND U118 ( .A(B[1]), .B(A[976]), .Z(\ab[976][1] ) );
  AND U119 ( .A(A[976]), .B(B[0]), .Z(\ab[976][0] ) );
  AND U120 ( .A(B[3]), .B(A[975]), .Z(\ab[975][3] ) );
  AND U121 ( .A(B[2]), .B(A[975]), .Z(\ab[975][2] ) );
  AND U122 ( .A(B[1]), .B(A[975]), .Z(\ab[975][1] ) );
  AND U123 ( .A(A[975]), .B(B[0]), .Z(\ab[975][0] ) );
  AND U124 ( .A(B[3]), .B(A[974]), .Z(\ab[974][3] ) );
  AND U125 ( .A(B[2]), .B(A[974]), .Z(\ab[974][2] ) );
  AND U126 ( .A(B[1]), .B(A[974]), .Z(\ab[974][1] ) );
  AND U127 ( .A(A[974]), .B(B[0]), .Z(\ab[974][0] ) );
  AND U128 ( .A(B[3]), .B(A[973]), .Z(\ab[973][3] ) );
  AND U129 ( .A(B[2]), .B(A[973]), .Z(\ab[973][2] ) );
  AND U130 ( .A(B[1]), .B(A[973]), .Z(\ab[973][1] ) );
  AND U131 ( .A(A[973]), .B(B[0]), .Z(\ab[973][0] ) );
  AND U132 ( .A(B[3]), .B(A[972]), .Z(\ab[972][3] ) );
  AND U133 ( .A(B[2]), .B(A[972]), .Z(\ab[972][2] ) );
  AND U134 ( .A(B[1]), .B(A[972]), .Z(\ab[972][1] ) );
  AND U135 ( .A(A[972]), .B(B[0]), .Z(\ab[972][0] ) );
  AND U136 ( .A(B[3]), .B(A[971]), .Z(\ab[971][3] ) );
  AND U137 ( .A(B[2]), .B(A[971]), .Z(\ab[971][2] ) );
  AND U138 ( .A(B[1]), .B(A[971]), .Z(\ab[971][1] ) );
  AND U139 ( .A(A[971]), .B(B[0]), .Z(\ab[971][0] ) );
  AND U140 ( .A(B[3]), .B(A[970]), .Z(\ab[970][3] ) );
  AND U141 ( .A(B[2]), .B(A[970]), .Z(\ab[970][2] ) );
  AND U142 ( .A(B[1]), .B(A[970]), .Z(\ab[970][1] ) );
  AND U143 ( .A(A[970]), .B(B[0]), .Z(\ab[970][0] ) );
  AND U144 ( .A(B[3]), .B(A[96]), .Z(\ab[96][3] ) );
  AND U145 ( .A(B[2]), .B(A[96]), .Z(\ab[96][2] ) );
  AND U146 ( .A(B[1]), .B(A[96]), .Z(\ab[96][1] ) );
  AND U147 ( .A(A[96]), .B(B[0]), .Z(\ab[96][0] ) );
  AND U148 ( .A(B[3]), .B(A[969]), .Z(\ab[969][3] ) );
  AND U149 ( .A(B[2]), .B(A[969]), .Z(\ab[969][2] ) );
  AND U150 ( .A(B[1]), .B(A[969]), .Z(\ab[969][1] ) );
  AND U151 ( .A(A[969]), .B(B[0]), .Z(\ab[969][0] ) );
  AND U152 ( .A(B[3]), .B(A[968]), .Z(\ab[968][3] ) );
  AND U153 ( .A(B[2]), .B(A[968]), .Z(\ab[968][2] ) );
  AND U154 ( .A(B[1]), .B(A[968]), .Z(\ab[968][1] ) );
  AND U155 ( .A(A[968]), .B(B[0]), .Z(\ab[968][0] ) );
  AND U156 ( .A(B[3]), .B(A[967]), .Z(\ab[967][3] ) );
  AND U157 ( .A(B[2]), .B(A[967]), .Z(\ab[967][2] ) );
  AND U158 ( .A(B[1]), .B(A[967]), .Z(\ab[967][1] ) );
  AND U159 ( .A(A[967]), .B(B[0]), .Z(\ab[967][0] ) );
  AND U160 ( .A(B[3]), .B(A[966]), .Z(\ab[966][3] ) );
  AND U161 ( .A(B[2]), .B(A[966]), .Z(\ab[966][2] ) );
  AND U162 ( .A(B[1]), .B(A[966]), .Z(\ab[966][1] ) );
  AND U163 ( .A(A[966]), .B(B[0]), .Z(\ab[966][0] ) );
  AND U164 ( .A(B[3]), .B(A[965]), .Z(\ab[965][3] ) );
  AND U165 ( .A(B[2]), .B(A[965]), .Z(\ab[965][2] ) );
  AND U166 ( .A(B[1]), .B(A[965]), .Z(\ab[965][1] ) );
  AND U167 ( .A(A[965]), .B(B[0]), .Z(\ab[965][0] ) );
  AND U168 ( .A(B[3]), .B(A[964]), .Z(\ab[964][3] ) );
  AND U169 ( .A(B[2]), .B(A[964]), .Z(\ab[964][2] ) );
  AND U170 ( .A(B[1]), .B(A[964]), .Z(\ab[964][1] ) );
  AND U171 ( .A(A[964]), .B(B[0]), .Z(\ab[964][0] ) );
  AND U172 ( .A(B[3]), .B(A[963]), .Z(\ab[963][3] ) );
  AND U173 ( .A(B[2]), .B(A[963]), .Z(\ab[963][2] ) );
  AND U174 ( .A(B[1]), .B(A[963]), .Z(\ab[963][1] ) );
  AND U175 ( .A(A[963]), .B(B[0]), .Z(\ab[963][0] ) );
  AND U176 ( .A(B[3]), .B(A[962]), .Z(\ab[962][3] ) );
  AND U177 ( .A(B[2]), .B(A[962]), .Z(\ab[962][2] ) );
  AND U178 ( .A(B[1]), .B(A[962]), .Z(\ab[962][1] ) );
  AND U179 ( .A(A[962]), .B(B[0]), .Z(\ab[962][0] ) );
  AND U180 ( .A(B[3]), .B(A[961]), .Z(\ab[961][3] ) );
  AND U181 ( .A(B[2]), .B(A[961]), .Z(\ab[961][2] ) );
  AND U182 ( .A(B[1]), .B(A[961]), .Z(\ab[961][1] ) );
  AND U183 ( .A(A[961]), .B(B[0]), .Z(\ab[961][0] ) );
  AND U184 ( .A(B[3]), .B(A[960]), .Z(\ab[960][3] ) );
  AND U185 ( .A(B[2]), .B(A[960]), .Z(\ab[960][2] ) );
  AND U186 ( .A(B[1]), .B(A[960]), .Z(\ab[960][1] ) );
  AND U187 ( .A(A[960]), .B(B[0]), .Z(\ab[960][0] ) );
  AND U188 ( .A(B[3]), .B(A[95]), .Z(\ab[95][3] ) );
  AND U189 ( .A(B[2]), .B(A[95]), .Z(\ab[95][2] ) );
  AND U190 ( .A(B[1]), .B(A[95]), .Z(\ab[95][1] ) );
  AND U191 ( .A(A[95]), .B(B[0]), .Z(\ab[95][0] ) );
  AND U192 ( .A(B[3]), .B(A[959]), .Z(\ab[959][3] ) );
  AND U193 ( .A(B[2]), .B(A[959]), .Z(\ab[959][2] ) );
  AND U194 ( .A(B[1]), .B(A[959]), .Z(\ab[959][1] ) );
  AND U195 ( .A(A[959]), .B(B[0]), .Z(\ab[959][0] ) );
  AND U196 ( .A(B[3]), .B(A[958]), .Z(\ab[958][3] ) );
  AND U197 ( .A(B[2]), .B(A[958]), .Z(\ab[958][2] ) );
  AND U198 ( .A(B[1]), .B(A[958]), .Z(\ab[958][1] ) );
  AND U199 ( .A(A[958]), .B(B[0]), .Z(\ab[958][0] ) );
  AND U200 ( .A(B[3]), .B(A[957]), .Z(\ab[957][3] ) );
  AND U201 ( .A(B[2]), .B(A[957]), .Z(\ab[957][2] ) );
  AND U202 ( .A(B[1]), .B(A[957]), .Z(\ab[957][1] ) );
  AND U203 ( .A(A[957]), .B(B[0]), .Z(\ab[957][0] ) );
  AND U204 ( .A(B[3]), .B(A[956]), .Z(\ab[956][3] ) );
  AND U205 ( .A(B[2]), .B(A[956]), .Z(\ab[956][2] ) );
  AND U206 ( .A(B[1]), .B(A[956]), .Z(\ab[956][1] ) );
  AND U207 ( .A(A[956]), .B(B[0]), .Z(\ab[956][0] ) );
  AND U208 ( .A(B[3]), .B(A[955]), .Z(\ab[955][3] ) );
  AND U209 ( .A(B[2]), .B(A[955]), .Z(\ab[955][2] ) );
  AND U210 ( .A(B[1]), .B(A[955]), .Z(\ab[955][1] ) );
  AND U211 ( .A(A[955]), .B(B[0]), .Z(\ab[955][0] ) );
  AND U212 ( .A(B[3]), .B(A[954]), .Z(\ab[954][3] ) );
  AND U213 ( .A(B[2]), .B(A[954]), .Z(\ab[954][2] ) );
  AND U214 ( .A(B[1]), .B(A[954]), .Z(\ab[954][1] ) );
  AND U215 ( .A(A[954]), .B(B[0]), .Z(\ab[954][0] ) );
  AND U216 ( .A(B[3]), .B(A[953]), .Z(\ab[953][3] ) );
  AND U217 ( .A(B[2]), .B(A[953]), .Z(\ab[953][2] ) );
  AND U218 ( .A(B[1]), .B(A[953]), .Z(\ab[953][1] ) );
  AND U219 ( .A(A[953]), .B(B[0]), .Z(\ab[953][0] ) );
  AND U220 ( .A(B[3]), .B(A[952]), .Z(\ab[952][3] ) );
  AND U221 ( .A(B[2]), .B(A[952]), .Z(\ab[952][2] ) );
  AND U222 ( .A(B[1]), .B(A[952]), .Z(\ab[952][1] ) );
  AND U223 ( .A(A[952]), .B(B[0]), .Z(\ab[952][0] ) );
  AND U224 ( .A(B[3]), .B(A[951]), .Z(\ab[951][3] ) );
  AND U225 ( .A(B[2]), .B(A[951]), .Z(\ab[951][2] ) );
  AND U226 ( .A(B[1]), .B(A[951]), .Z(\ab[951][1] ) );
  AND U227 ( .A(A[951]), .B(B[0]), .Z(\ab[951][0] ) );
  AND U228 ( .A(B[3]), .B(A[950]), .Z(\ab[950][3] ) );
  AND U229 ( .A(B[2]), .B(A[950]), .Z(\ab[950][2] ) );
  AND U230 ( .A(B[1]), .B(A[950]), .Z(\ab[950][1] ) );
  AND U231 ( .A(A[950]), .B(B[0]), .Z(\ab[950][0] ) );
  AND U232 ( .A(B[3]), .B(A[94]), .Z(\ab[94][3] ) );
  AND U233 ( .A(B[2]), .B(A[94]), .Z(\ab[94][2] ) );
  AND U234 ( .A(B[1]), .B(A[94]), .Z(\ab[94][1] ) );
  AND U235 ( .A(A[94]), .B(B[0]), .Z(\ab[94][0] ) );
  AND U236 ( .A(B[3]), .B(A[949]), .Z(\ab[949][3] ) );
  AND U237 ( .A(B[2]), .B(A[949]), .Z(\ab[949][2] ) );
  AND U238 ( .A(B[1]), .B(A[949]), .Z(\ab[949][1] ) );
  AND U239 ( .A(A[949]), .B(B[0]), .Z(\ab[949][0] ) );
  AND U240 ( .A(B[3]), .B(A[948]), .Z(\ab[948][3] ) );
  AND U241 ( .A(B[2]), .B(A[948]), .Z(\ab[948][2] ) );
  AND U242 ( .A(B[1]), .B(A[948]), .Z(\ab[948][1] ) );
  AND U243 ( .A(A[948]), .B(B[0]), .Z(\ab[948][0] ) );
  AND U244 ( .A(B[3]), .B(A[947]), .Z(\ab[947][3] ) );
  AND U245 ( .A(B[2]), .B(A[947]), .Z(\ab[947][2] ) );
  AND U246 ( .A(B[1]), .B(A[947]), .Z(\ab[947][1] ) );
  AND U247 ( .A(A[947]), .B(B[0]), .Z(\ab[947][0] ) );
  AND U248 ( .A(B[3]), .B(A[946]), .Z(\ab[946][3] ) );
  AND U249 ( .A(B[2]), .B(A[946]), .Z(\ab[946][2] ) );
  AND U250 ( .A(B[1]), .B(A[946]), .Z(\ab[946][1] ) );
  AND U251 ( .A(A[946]), .B(B[0]), .Z(\ab[946][0] ) );
  AND U252 ( .A(B[3]), .B(A[945]), .Z(\ab[945][3] ) );
  AND U253 ( .A(B[2]), .B(A[945]), .Z(\ab[945][2] ) );
  AND U254 ( .A(B[1]), .B(A[945]), .Z(\ab[945][1] ) );
  AND U255 ( .A(A[945]), .B(B[0]), .Z(\ab[945][0] ) );
  AND U256 ( .A(B[3]), .B(A[944]), .Z(\ab[944][3] ) );
  AND U257 ( .A(B[2]), .B(A[944]), .Z(\ab[944][2] ) );
  AND U258 ( .A(B[1]), .B(A[944]), .Z(\ab[944][1] ) );
  AND U259 ( .A(A[944]), .B(B[0]), .Z(\ab[944][0] ) );
  AND U260 ( .A(B[3]), .B(A[943]), .Z(\ab[943][3] ) );
  AND U261 ( .A(B[2]), .B(A[943]), .Z(\ab[943][2] ) );
  AND U262 ( .A(B[1]), .B(A[943]), .Z(\ab[943][1] ) );
  AND U263 ( .A(A[943]), .B(B[0]), .Z(\ab[943][0] ) );
  AND U264 ( .A(B[3]), .B(A[942]), .Z(\ab[942][3] ) );
  AND U265 ( .A(B[2]), .B(A[942]), .Z(\ab[942][2] ) );
  AND U266 ( .A(B[1]), .B(A[942]), .Z(\ab[942][1] ) );
  AND U267 ( .A(A[942]), .B(B[0]), .Z(\ab[942][0] ) );
  AND U268 ( .A(B[3]), .B(A[941]), .Z(\ab[941][3] ) );
  AND U269 ( .A(B[2]), .B(A[941]), .Z(\ab[941][2] ) );
  AND U270 ( .A(B[1]), .B(A[941]), .Z(\ab[941][1] ) );
  AND U271 ( .A(A[941]), .B(B[0]), .Z(\ab[941][0] ) );
  AND U272 ( .A(B[3]), .B(A[940]), .Z(\ab[940][3] ) );
  AND U273 ( .A(B[2]), .B(A[940]), .Z(\ab[940][2] ) );
  AND U274 ( .A(B[1]), .B(A[940]), .Z(\ab[940][1] ) );
  AND U275 ( .A(A[940]), .B(B[0]), .Z(\ab[940][0] ) );
  AND U276 ( .A(B[3]), .B(A[93]), .Z(\ab[93][3] ) );
  AND U277 ( .A(B[2]), .B(A[93]), .Z(\ab[93][2] ) );
  AND U278 ( .A(B[1]), .B(A[93]), .Z(\ab[93][1] ) );
  AND U279 ( .A(A[93]), .B(B[0]), .Z(\ab[93][0] ) );
  AND U280 ( .A(B[3]), .B(A[939]), .Z(\ab[939][3] ) );
  AND U281 ( .A(B[2]), .B(A[939]), .Z(\ab[939][2] ) );
  AND U282 ( .A(B[1]), .B(A[939]), .Z(\ab[939][1] ) );
  AND U283 ( .A(A[939]), .B(B[0]), .Z(\ab[939][0] ) );
  AND U284 ( .A(B[3]), .B(A[938]), .Z(\ab[938][3] ) );
  AND U285 ( .A(B[2]), .B(A[938]), .Z(\ab[938][2] ) );
  AND U286 ( .A(B[1]), .B(A[938]), .Z(\ab[938][1] ) );
  AND U287 ( .A(A[938]), .B(B[0]), .Z(\ab[938][0] ) );
  AND U288 ( .A(B[3]), .B(A[937]), .Z(\ab[937][3] ) );
  AND U289 ( .A(B[2]), .B(A[937]), .Z(\ab[937][2] ) );
  AND U290 ( .A(B[1]), .B(A[937]), .Z(\ab[937][1] ) );
  AND U291 ( .A(A[937]), .B(B[0]), .Z(\ab[937][0] ) );
  AND U292 ( .A(B[3]), .B(A[936]), .Z(\ab[936][3] ) );
  AND U293 ( .A(B[2]), .B(A[936]), .Z(\ab[936][2] ) );
  AND U294 ( .A(B[1]), .B(A[936]), .Z(\ab[936][1] ) );
  AND U295 ( .A(A[936]), .B(B[0]), .Z(\ab[936][0] ) );
  AND U296 ( .A(B[3]), .B(A[935]), .Z(\ab[935][3] ) );
  AND U297 ( .A(B[2]), .B(A[935]), .Z(\ab[935][2] ) );
  AND U298 ( .A(B[1]), .B(A[935]), .Z(\ab[935][1] ) );
  AND U299 ( .A(A[935]), .B(B[0]), .Z(\ab[935][0] ) );
  AND U300 ( .A(B[3]), .B(A[934]), .Z(\ab[934][3] ) );
  AND U301 ( .A(B[2]), .B(A[934]), .Z(\ab[934][2] ) );
  AND U302 ( .A(B[1]), .B(A[934]), .Z(\ab[934][1] ) );
  AND U303 ( .A(A[934]), .B(B[0]), .Z(\ab[934][0] ) );
  AND U304 ( .A(B[3]), .B(A[933]), .Z(\ab[933][3] ) );
  AND U305 ( .A(B[2]), .B(A[933]), .Z(\ab[933][2] ) );
  AND U306 ( .A(B[1]), .B(A[933]), .Z(\ab[933][1] ) );
  AND U307 ( .A(A[933]), .B(B[0]), .Z(\ab[933][0] ) );
  AND U308 ( .A(B[3]), .B(A[932]), .Z(\ab[932][3] ) );
  AND U309 ( .A(B[2]), .B(A[932]), .Z(\ab[932][2] ) );
  AND U310 ( .A(B[1]), .B(A[932]), .Z(\ab[932][1] ) );
  AND U311 ( .A(A[932]), .B(B[0]), .Z(\ab[932][0] ) );
  AND U312 ( .A(B[3]), .B(A[931]), .Z(\ab[931][3] ) );
  AND U313 ( .A(B[2]), .B(A[931]), .Z(\ab[931][2] ) );
  AND U314 ( .A(B[1]), .B(A[931]), .Z(\ab[931][1] ) );
  AND U315 ( .A(A[931]), .B(B[0]), .Z(\ab[931][0] ) );
  AND U316 ( .A(B[3]), .B(A[930]), .Z(\ab[930][3] ) );
  AND U317 ( .A(B[2]), .B(A[930]), .Z(\ab[930][2] ) );
  AND U318 ( .A(B[1]), .B(A[930]), .Z(\ab[930][1] ) );
  AND U319 ( .A(A[930]), .B(B[0]), .Z(\ab[930][0] ) );
  AND U320 ( .A(B[3]), .B(A[92]), .Z(\ab[92][3] ) );
  AND U321 ( .A(B[2]), .B(A[92]), .Z(\ab[92][2] ) );
  AND U322 ( .A(B[1]), .B(A[92]), .Z(\ab[92][1] ) );
  AND U323 ( .A(A[92]), .B(B[0]), .Z(\ab[92][0] ) );
  AND U324 ( .A(B[3]), .B(A[929]), .Z(\ab[929][3] ) );
  AND U325 ( .A(B[2]), .B(A[929]), .Z(\ab[929][2] ) );
  AND U326 ( .A(B[1]), .B(A[929]), .Z(\ab[929][1] ) );
  AND U327 ( .A(A[929]), .B(B[0]), .Z(\ab[929][0] ) );
  AND U328 ( .A(B[3]), .B(A[928]), .Z(\ab[928][3] ) );
  AND U329 ( .A(B[2]), .B(A[928]), .Z(\ab[928][2] ) );
  AND U330 ( .A(B[1]), .B(A[928]), .Z(\ab[928][1] ) );
  AND U331 ( .A(A[928]), .B(B[0]), .Z(\ab[928][0] ) );
  AND U332 ( .A(B[3]), .B(A[927]), .Z(\ab[927][3] ) );
  AND U333 ( .A(B[2]), .B(A[927]), .Z(\ab[927][2] ) );
  AND U334 ( .A(B[1]), .B(A[927]), .Z(\ab[927][1] ) );
  AND U335 ( .A(A[927]), .B(B[0]), .Z(\ab[927][0] ) );
  AND U336 ( .A(B[3]), .B(A[926]), .Z(\ab[926][3] ) );
  AND U337 ( .A(B[2]), .B(A[926]), .Z(\ab[926][2] ) );
  AND U338 ( .A(B[1]), .B(A[926]), .Z(\ab[926][1] ) );
  AND U339 ( .A(A[926]), .B(B[0]), .Z(\ab[926][0] ) );
  AND U340 ( .A(B[3]), .B(A[925]), .Z(\ab[925][3] ) );
  AND U341 ( .A(B[2]), .B(A[925]), .Z(\ab[925][2] ) );
  AND U342 ( .A(B[1]), .B(A[925]), .Z(\ab[925][1] ) );
  AND U343 ( .A(A[925]), .B(B[0]), .Z(\ab[925][0] ) );
  AND U344 ( .A(B[3]), .B(A[924]), .Z(\ab[924][3] ) );
  AND U345 ( .A(B[2]), .B(A[924]), .Z(\ab[924][2] ) );
  AND U346 ( .A(B[1]), .B(A[924]), .Z(\ab[924][1] ) );
  AND U347 ( .A(A[924]), .B(B[0]), .Z(\ab[924][0] ) );
  AND U348 ( .A(B[3]), .B(A[923]), .Z(\ab[923][3] ) );
  AND U349 ( .A(B[2]), .B(A[923]), .Z(\ab[923][2] ) );
  AND U350 ( .A(B[1]), .B(A[923]), .Z(\ab[923][1] ) );
  AND U351 ( .A(A[923]), .B(B[0]), .Z(\ab[923][0] ) );
  AND U352 ( .A(B[3]), .B(A[922]), .Z(\ab[922][3] ) );
  AND U353 ( .A(B[2]), .B(A[922]), .Z(\ab[922][2] ) );
  AND U354 ( .A(B[1]), .B(A[922]), .Z(\ab[922][1] ) );
  AND U355 ( .A(A[922]), .B(B[0]), .Z(\ab[922][0] ) );
  AND U356 ( .A(B[3]), .B(A[921]), .Z(\ab[921][3] ) );
  AND U357 ( .A(B[2]), .B(A[921]), .Z(\ab[921][2] ) );
  AND U358 ( .A(B[1]), .B(A[921]), .Z(\ab[921][1] ) );
  AND U359 ( .A(A[921]), .B(B[0]), .Z(\ab[921][0] ) );
  AND U360 ( .A(B[3]), .B(A[920]), .Z(\ab[920][3] ) );
  AND U361 ( .A(B[2]), .B(A[920]), .Z(\ab[920][2] ) );
  AND U362 ( .A(B[1]), .B(A[920]), .Z(\ab[920][1] ) );
  AND U363 ( .A(A[920]), .B(B[0]), .Z(\ab[920][0] ) );
  AND U364 ( .A(B[3]), .B(A[91]), .Z(\ab[91][3] ) );
  AND U365 ( .A(B[2]), .B(A[91]), .Z(\ab[91][2] ) );
  AND U366 ( .A(B[1]), .B(A[91]), .Z(\ab[91][1] ) );
  AND U367 ( .A(A[91]), .B(B[0]), .Z(\ab[91][0] ) );
  AND U368 ( .A(B[3]), .B(A[919]), .Z(\ab[919][3] ) );
  AND U369 ( .A(B[2]), .B(A[919]), .Z(\ab[919][2] ) );
  AND U370 ( .A(B[1]), .B(A[919]), .Z(\ab[919][1] ) );
  AND U371 ( .A(A[919]), .B(B[0]), .Z(\ab[919][0] ) );
  AND U372 ( .A(B[3]), .B(A[918]), .Z(\ab[918][3] ) );
  AND U373 ( .A(B[2]), .B(A[918]), .Z(\ab[918][2] ) );
  AND U374 ( .A(B[1]), .B(A[918]), .Z(\ab[918][1] ) );
  AND U375 ( .A(A[918]), .B(B[0]), .Z(\ab[918][0] ) );
  AND U376 ( .A(B[3]), .B(A[917]), .Z(\ab[917][3] ) );
  AND U377 ( .A(B[2]), .B(A[917]), .Z(\ab[917][2] ) );
  AND U378 ( .A(B[1]), .B(A[917]), .Z(\ab[917][1] ) );
  AND U379 ( .A(A[917]), .B(B[0]), .Z(\ab[917][0] ) );
  AND U380 ( .A(B[3]), .B(A[916]), .Z(\ab[916][3] ) );
  AND U381 ( .A(B[2]), .B(A[916]), .Z(\ab[916][2] ) );
  AND U382 ( .A(B[1]), .B(A[916]), .Z(\ab[916][1] ) );
  AND U383 ( .A(A[916]), .B(B[0]), .Z(\ab[916][0] ) );
  AND U384 ( .A(B[3]), .B(A[915]), .Z(\ab[915][3] ) );
  AND U385 ( .A(B[2]), .B(A[915]), .Z(\ab[915][2] ) );
  AND U386 ( .A(B[1]), .B(A[915]), .Z(\ab[915][1] ) );
  AND U387 ( .A(A[915]), .B(B[0]), .Z(\ab[915][0] ) );
  AND U388 ( .A(B[3]), .B(A[914]), .Z(\ab[914][3] ) );
  AND U389 ( .A(B[2]), .B(A[914]), .Z(\ab[914][2] ) );
  AND U390 ( .A(B[1]), .B(A[914]), .Z(\ab[914][1] ) );
  AND U391 ( .A(A[914]), .B(B[0]), .Z(\ab[914][0] ) );
  AND U392 ( .A(B[3]), .B(A[913]), .Z(\ab[913][3] ) );
  AND U393 ( .A(B[2]), .B(A[913]), .Z(\ab[913][2] ) );
  AND U394 ( .A(B[1]), .B(A[913]), .Z(\ab[913][1] ) );
  AND U395 ( .A(A[913]), .B(B[0]), .Z(\ab[913][0] ) );
  AND U396 ( .A(B[3]), .B(A[912]), .Z(\ab[912][3] ) );
  AND U397 ( .A(B[2]), .B(A[912]), .Z(\ab[912][2] ) );
  AND U398 ( .A(B[1]), .B(A[912]), .Z(\ab[912][1] ) );
  AND U399 ( .A(A[912]), .B(B[0]), .Z(\ab[912][0] ) );
  AND U400 ( .A(B[3]), .B(A[911]), .Z(\ab[911][3] ) );
  AND U401 ( .A(B[2]), .B(A[911]), .Z(\ab[911][2] ) );
  AND U402 ( .A(B[1]), .B(A[911]), .Z(\ab[911][1] ) );
  AND U403 ( .A(A[911]), .B(B[0]), .Z(\ab[911][0] ) );
  AND U404 ( .A(B[3]), .B(A[910]), .Z(\ab[910][3] ) );
  AND U405 ( .A(B[2]), .B(A[910]), .Z(\ab[910][2] ) );
  AND U406 ( .A(B[1]), .B(A[910]), .Z(\ab[910][1] ) );
  AND U407 ( .A(A[910]), .B(B[0]), .Z(\ab[910][0] ) );
  AND U408 ( .A(B[3]), .B(A[90]), .Z(\ab[90][3] ) );
  AND U409 ( .A(B[2]), .B(A[90]), .Z(\ab[90][2] ) );
  AND U410 ( .A(B[1]), .B(A[90]), .Z(\ab[90][1] ) );
  AND U411 ( .A(A[90]), .B(B[0]), .Z(\ab[90][0] ) );
  AND U412 ( .A(B[3]), .B(A[909]), .Z(\ab[909][3] ) );
  AND U413 ( .A(B[2]), .B(A[909]), .Z(\ab[909][2] ) );
  AND U414 ( .A(B[1]), .B(A[909]), .Z(\ab[909][1] ) );
  AND U415 ( .A(A[909]), .B(B[0]), .Z(\ab[909][0] ) );
  AND U416 ( .A(B[3]), .B(A[908]), .Z(\ab[908][3] ) );
  AND U417 ( .A(B[2]), .B(A[908]), .Z(\ab[908][2] ) );
  AND U418 ( .A(B[1]), .B(A[908]), .Z(\ab[908][1] ) );
  AND U419 ( .A(A[908]), .B(B[0]), .Z(\ab[908][0] ) );
  AND U420 ( .A(B[3]), .B(A[907]), .Z(\ab[907][3] ) );
  AND U421 ( .A(B[2]), .B(A[907]), .Z(\ab[907][2] ) );
  AND U422 ( .A(B[1]), .B(A[907]), .Z(\ab[907][1] ) );
  AND U423 ( .A(A[907]), .B(B[0]), .Z(\ab[907][0] ) );
  AND U424 ( .A(B[3]), .B(A[906]), .Z(\ab[906][3] ) );
  AND U425 ( .A(B[2]), .B(A[906]), .Z(\ab[906][2] ) );
  AND U426 ( .A(B[1]), .B(A[906]), .Z(\ab[906][1] ) );
  AND U427 ( .A(A[906]), .B(B[0]), .Z(\ab[906][0] ) );
  AND U428 ( .A(B[3]), .B(A[905]), .Z(\ab[905][3] ) );
  AND U429 ( .A(B[2]), .B(A[905]), .Z(\ab[905][2] ) );
  AND U430 ( .A(B[1]), .B(A[905]), .Z(\ab[905][1] ) );
  AND U431 ( .A(A[905]), .B(B[0]), .Z(\ab[905][0] ) );
  AND U432 ( .A(B[3]), .B(A[904]), .Z(\ab[904][3] ) );
  AND U433 ( .A(B[2]), .B(A[904]), .Z(\ab[904][2] ) );
  AND U434 ( .A(B[1]), .B(A[904]), .Z(\ab[904][1] ) );
  AND U435 ( .A(A[904]), .B(B[0]), .Z(\ab[904][0] ) );
  AND U436 ( .A(B[3]), .B(A[903]), .Z(\ab[903][3] ) );
  AND U437 ( .A(B[2]), .B(A[903]), .Z(\ab[903][2] ) );
  AND U438 ( .A(B[1]), .B(A[903]), .Z(\ab[903][1] ) );
  AND U439 ( .A(A[903]), .B(B[0]), .Z(\ab[903][0] ) );
  AND U440 ( .A(B[3]), .B(A[902]), .Z(\ab[902][3] ) );
  AND U441 ( .A(B[2]), .B(A[902]), .Z(\ab[902][2] ) );
  AND U442 ( .A(B[1]), .B(A[902]), .Z(\ab[902][1] ) );
  AND U443 ( .A(A[902]), .B(B[0]), .Z(\ab[902][0] ) );
  AND U444 ( .A(B[3]), .B(A[901]), .Z(\ab[901][3] ) );
  AND U445 ( .A(B[2]), .B(A[901]), .Z(\ab[901][2] ) );
  AND U446 ( .A(B[1]), .B(A[901]), .Z(\ab[901][1] ) );
  AND U447 ( .A(A[901]), .B(B[0]), .Z(\ab[901][0] ) );
  AND U448 ( .A(B[3]), .B(A[900]), .Z(\ab[900][3] ) );
  AND U449 ( .A(B[2]), .B(A[900]), .Z(\ab[900][2] ) );
  AND U450 ( .A(B[1]), .B(A[900]), .Z(\ab[900][1] ) );
  AND U451 ( .A(A[900]), .B(B[0]), .Z(\ab[900][0] ) );
  AND U452 ( .A(B[3]), .B(A[8]), .Z(\ab[8][3] ) );
  AND U453 ( .A(B[2]), .B(A[8]), .Z(\ab[8][2] ) );
  AND U454 ( .A(B[1]), .B(A[8]), .Z(\ab[8][1] ) );
  AND U455 ( .A(A[8]), .B(B[0]), .Z(\ab[8][0] ) );
  AND U456 ( .A(B[3]), .B(A[89]), .Z(\ab[89][3] ) );
  AND U457 ( .A(B[2]), .B(A[89]), .Z(\ab[89][2] ) );
  AND U458 ( .A(B[1]), .B(A[89]), .Z(\ab[89][1] ) );
  AND U459 ( .A(A[89]), .B(B[0]), .Z(\ab[89][0] ) );
  AND U460 ( .A(B[3]), .B(A[899]), .Z(\ab[899][3] ) );
  AND U461 ( .A(B[2]), .B(A[899]), .Z(\ab[899][2] ) );
  AND U462 ( .A(B[1]), .B(A[899]), .Z(\ab[899][1] ) );
  AND U463 ( .A(A[899]), .B(B[0]), .Z(\ab[899][0] ) );
  AND U464 ( .A(B[3]), .B(A[898]), .Z(\ab[898][3] ) );
  AND U465 ( .A(B[2]), .B(A[898]), .Z(\ab[898][2] ) );
  AND U466 ( .A(B[1]), .B(A[898]), .Z(\ab[898][1] ) );
  AND U467 ( .A(A[898]), .B(B[0]), .Z(\ab[898][0] ) );
  AND U468 ( .A(B[3]), .B(A[897]), .Z(\ab[897][3] ) );
  AND U469 ( .A(B[2]), .B(A[897]), .Z(\ab[897][2] ) );
  AND U470 ( .A(B[1]), .B(A[897]), .Z(\ab[897][1] ) );
  AND U471 ( .A(A[897]), .B(B[0]), .Z(\ab[897][0] ) );
  AND U472 ( .A(B[3]), .B(A[896]), .Z(\ab[896][3] ) );
  AND U473 ( .A(B[2]), .B(A[896]), .Z(\ab[896][2] ) );
  AND U474 ( .A(B[1]), .B(A[896]), .Z(\ab[896][1] ) );
  AND U475 ( .A(A[896]), .B(B[0]), .Z(\ab[896][0] ) );
  AND U476 ( .A(B[3]), .B(A[895]), .Z(\ab[895][3] ) );
  AND U477 ( .A(B[2]), .B(A[895]), .Z(\ab[895][2] ) );
  AND U478 ( .A(B[1]), .B(A[895]), .Z(\ab[895][1] ) );
  AND U479 ( .A(A[895]), .B(B[0]), .Z(\ab[895][0] ) );
  AND U480 ( .A(B[3]), .B(A[894]), .Z(\ab[894][3] ) );
  AND U481 ( .A(B[2]), .B(A[894]), .Z(\ab[894][2] ) );
  AND U482 ( .A(B[1]), .B(A[894]), .Z(\ab[894][1] ) );
  AND U483 ( .A(A[894]), .B(B[0]), .Z(\ab[894][0] ) );
  AND U484 ( .A(B[3]), .B(A[893]), .Z(\ab[893][3] ) );
  AND U485 ( .A(B[2]), .B(A[893]), .Z(\ab[893][2] ) );
  AND U486 ( .A(B[1]), .B(A[893]), .Z(\ab[893][1] ) );
  AND U487 ( .A(A[893]), .B(B[0]), .Z(\ab[893][0] ) );
  AND U488 ( .A(B[3]), .B(A[892]), .Z(\ab[892][3] ) );
  AND U489 ( .A(B[2]), .B(A[892]), .Z(\ab[892][2] ) );
  AND U490 ( .A(B[1]), .B(A[892]), .Z(\ab[892][1] ) );
  AND U491 ( .A(A[892]), .B(B[0]), .Z(\ab[892][0] ) );
  AND U492 ( .A(B[3]), .B(A[891]), .Z(\ab[891][3] ) );
  AND U493 ( .A(B[2]), .B(A[891]), .Z(\ab[891][2] ) );
  AND U494 ( .A(B[1]), .B(A[891]), .Z(\ab[891][1] ) );
  AND U495 ( .A(A[891]), .B(B[0]), .Z(\ab[891][0] ) );
  AND U496 ( .A(B[3]), .B(A[890]), .Z(\ab[890][3] ) );
  AND U497 ( .A(B[2]), .B(A[890]), .Z(\ab[890][2] ) );
  AND U498 ( .A(B[1]), .B(A[890]), .Z(\ab[890][1] ) );
  AND U499 ( .A(A[890]), .B(B[0]), .Z(\ab[890][0] ) );
  AND U500 ( .A(B[3]), .B(A[88]), .Z(\ab[88][3] ) );
  AND U501 ( .A(B[2]), .B(A[88]), .Z(\ab[88][2] ) );
  AND U502 ( .A(B[1]), .B(A[88]), .Z(\ab[88][1] ) );
  AND U503 ( .A(A[88]), .B(B[0]), .Z(\ab[88][0] ) );
  AND U504 ( .A(B[3]), .B(A[889]), .Z(\ab[889][3] ) );
  AND U505 ( .A(B[2]), .B(A[889]), .Z(\ab[889][2] ) );
  AND U506 ( .A(B[1]), .B(A[889]), .Z(\ab[889][1] ) );
  AND U507 ( .A(A[889]), .B(B[0]), .Z(\ab[889][0] ) );
  AND U508 ( .A(B[3]), .B(A[888]), .Z(\ab[888][3] ) );
  AND U509 ( .A(B[2]), .B(A[888]), .Z(\ab[888][2] ) );
  AND U510 ( .A(B[1]), .B(A[888]), .Z(\ab[888][1] ) );
  AND U511 ( .A(A[888]), .B(B[0]), .Z(\ab[888][0] ) );
  AND U512 ( .A(B[3]), .B(A[887]), .Z(\ab[887][3] ) );
  AND U513 ( .A(B[2]), .B(A[887]), .Z(\ab[887][2] ) );
  AND U514 ( .A(B[1]), .B(A[887]), .Z(\ab[887][1] ) );
  AND U515 ( .A(A[887]), .B(B[0]), .Z(\ab[887][0] ) );
  AND U516 ( .A(B[3]), .B(A[886]), .Z(\ab[886][3] ) );
  AND U517 ( .A(B[2]), .B(A[886]), .Z(\ab[886][2] ) );
  AND U518 ( .A(B[1]), .B(A[886]), .Z(\ab[886][1] ) );
  AND U519 ( .A(A[886]), .B(B[0]), .Z(\ab[886][0] ) );
  AND U520 ( .A(B[3]), .B(A[885]), .Z(\ab[885][3] ) );
  AND U521 ( .A(B[2]), .B(A[885]), .Z(\ab[885][2] ) );
  AND U522 ( .A(B[1]), .B(A[885]), .Z(\ab[885][1] ) );
  AND U523 ( .A(A[885]), .B(B[0]), .Z(\ab[885][0] ) );
  AND U524 ( .A(B[3]), .B(A[884]), .Z(\ab[884][3] ) );
  AND U525 ( .A(B[2]), .B(A[884]), .Z(\ab[884][2] ) );
  AND U526 ( .A(B[1]), .B(A[884]), .Z(\ab[884][1] ) );
  AND U527 ( .A(A[884]), .B(B[0]), .Z(\ab[884][0] ) );
  AND U528 ( .A(B[3]), .B(A[883]), .Z(\ab[883][3] ) );
  AND U529 ( .A(B[2]), .B(A[883]), .Z(\ab[883][2] ) );
  AND U530 ( .A(B[1]), .B(A[883]), .Z(\ab[883][1] ) );
  AND U531 ( .A(A[883]), .B(B[0]), .Z(\ab[883][0] ) );
  AND U532 ( .A(B[3]), .B(A[882]), .Z(\ab[882][3] ) );
  AND U533 ( .A(B[2]), .B(A[882]), .Z(\ab[882][2] ) );
  AND U534 ( .A(B[1]), .B(A[882]), .Z(\ab[882][1] ) );
  AND U535 ( .A(A[882]), .B(B[0]), .Z(\ab[882][0] ) );
  AND U536 ( .A(B[3]), .B(A[881]), .Z(\ab[881][3] ) );
  AND U537 ( .A(B[2]), .B(A[881]), .Z(\ab[881][2] ) );
  AND U538 ( .A(B[1]), .B(A[881]), .Z(\ab[881][1] ) );
  AND U539 ( .A(A[881]), .B(B[0]), .Z(\ab[881][0] ) );
  AND U540 ( .A(B[3]), .B(A[880]), .Z(\ab[880][3] ) );
  AND U541 ( .A(B[2]), .B(A[880]), .Z(\ab[880][2] ) );
  AND U542 ( .A(B[1]), .B(A[880]), .Z(\ab[880][1] ) );
  AND U543 ( .A(A[880]), .B(B[0]), .Z(\ab[880][0] ) );
  AND U544 ( .A(B[3]), .B(A[87]), .Z(\ab[87][3] ) );
  AND U545 ( .A(B[2]), .B(A[87]), .Z(\ab[87][2] ) );
  AND U546 ( .A(B[1]), .B(A[87]), .Z(\ab[87][1] ) );
  AND U547 ( .A(A[87]), .B(B[0]), .Z(\ab[87][0] ) );
  AND U548 ( .A(B[3]), .B(A[879]), .Z(\ab[879][3] ) );
  AND U549 ( .A(B[2]), .B(A[879]), .Z(\ab[879][2] ) );
  AND U550 ( .A(B[1]), .B(A[879]), .Z(\ab[879][1] ) );
  AND U551 ( .A(A[879]), .B(B[0]), .Z(\ab[879][0] ) );
  AND U552 ( .A(B[3]), .B(A[878]), .Z(\ab[878][3] ) );
  AND U553 ( .A(B[2]), .B(A[878]), .Z(\ab[878][2] ) );
  AND U554 ( .A(B[1]), .B(A[878]), .Z(\ab[878][1] ) );
  AND U555 ( .A(A[878]), .B(B[0]), .Z(\ab[878][0] ) );
  AND U556 ( .A(B[3]), .B(A[877]), .Z(\ab[877][3] ) );
  AND U557 ( .A(B[2]), .B(A[877]), .Z(\ab[877][2] ) );
  AND U558 ( .A(B[1]), .B(A[877]), .Z(\ab[877][1] ) );
  AND U559 ( .A(A[877]), .B(B[0]), .Z(\ab[877][0] ) );
  AND U560 ( .A(B[3]), .B(A[876]), .Z(\ab[876][3] ) );
  AND U561 ( .A(B[2]), .B(A[876]), .Z(\ab[876][2] ) );
  AND U562 ( .A(B[1]), .B(A[876]), .Z(\ab[876][1] ) );
  AND U563 ( .A(A[876]), .B(B[0]), .Z(\ab[876][0] ) );
  AND U564 ( .A(B[3]), .B(A[875]), .Z(\ab[875][3] ) );
  AND U565 ( .A(B[2]), .B(A[875]), .Z(\ab[875][2] ) );
  AND U566 ( .A(B[1]), .B(A[875]), .Z(\ab[875][1] ) );
  AND U567 ( .A(A[875]), .B(B[0]), .Z(\ab[875][0] ) );
  AND U568 ( .A(B[3]), .B(A[874]), .Z(\ab[874][3] ) );
  AND U569 ( .A(B[2]), .B(A[874]), .Z(\ab[874][2] ) );
  AND U570 ( .A(B[1]), .B(A[874]), .Z(\ab[874][1] ) );
  AND U571 ( .A(A[874]), .B(B[0]), .Z(\ab[874][0] ) );
  AND U572 ( .A(B[3]), .B(A[873]), .Z(\ab[873][3] ) );
  AND U573 ( .A(B[2]), .B(A[873]), .Z(\ab[873][2] ) );
  AND U574 ( .A(B[1]), .B(A[873]), .Z(\ab[873][1] ) );
  AND U575 ( .A(A[873]), .B(B[0]), .Z(\ab[873][0] ) );
  AND U576 ( .A(B[3]), .B(A[872]), .Z(\ab[872][3] ) );
  AND U577 ( .A(B[2]), .B(A[872]), .Z(\ab[872][2] ) );
  AND U578 ( .A(B[1]), .B(A[872]), .Z(\ab[872][1] ) );
  AND U579 ( .A(A[872]), .B(B[0]), .Z(\ab[872][0] ) );
  AND U580 ( .A(B[3]), .B(A[871]), .Z(\ab[871][3] ) );
  AND U581 ( .A(B[2]), .B(A[871]), .Z(\ab[871][2] ) );
  AND U582 ( .A(B[1]), .B(A[871]), .Z(\ab[871][1] ) );
  AND U583 ( .A(A[871]), .B(B[0]), .Z(\ab[871][0] ) );
  AND U584 ( .A(B[3]), .B(A[870]), .Z(\ab[870][3] ) );
  AND U585 ( .A(B[2]), .B(A[870]), .Z(\ab[870][2] ) );
  AND U586 ( .A(B[1]), .B(A[870]), .Z(\ab[870][1] ) );
  AND U587 ( .A(A[870]), .B(B[0]), .Z(\ab[870][0] ) );
  AND U588 ( .A(B[3]), .B(A[86]), .Z(\ab[86][3] ) );
  AND U589 ( .A(B[2]), .B(A[86]), .Z(\ab[86][2] ) );
  AND U590 ( .A(B[1]), .B(A[86]), .Z(\ab[86][1] ) );
  AND U591 ( .A(A[86]), .B(B[0]), .Z(\ab[86][0] ) );
  AND U592 ( .A(B[3]), .B(A[869]), .Z(\ab[869][3] ) );
  AND U593 ( .A(B[2]), .B(A[869]), .Z(\ab[869][2] ) );
  AND U594 ( .A(B[1]), .B(A[869]), .Z(\ab[869][1] ) );
  AND U595 ( .A(A[869]), .B(B[0]), .Z(\ab[869][0] ) );
  AND U596 ( .A(B[3]), .B(A[868]), .Z(\ab[868][3] ) );
  AND U597 ( .A(B[2]), .B(A[868]), .Z(\ab[868][2] ) );
  AND U598 ( .A(B[1]), .B(A[868]), .Z(\ab[868][1] ) );
  AND U599 ( .A(A[868]), .B(B[0]), .Z(\ab[868][0] ) );
  AND U600 ( .A(B[3]), .B(A[867]), .Z(\ab[867][3] ) );
  AND U601 ( .A(B[2]), .B(A[867]), .Z(\ab[867][2] ) );
  AND U602 ( .A(B[1]), .B(A[867]), .Z(\ab[867][1] ) );
  AND U603 ( .A(A[867]), .B(B[0]), .Z(\ab[867][0] ) );
  AND U604 ( .A(B[3]), .B(A[866]), .Z(\ab[866][3] ) );
  AND U605 ( .A(B[2]), .B(A[866]), .Z(\ab[866][2] ) );
  AND U606 ( .A(B[1]), .B(A[866]), .Z(\ab[866][1] ) );
  AND U607 ( .A(A[866]), .B(B[0]), .Z(\ab[866][0] ) );
  AND U608 ( .A(B[3]), .B(A[865]), .Z(\ab[865][3] ) );
  AND U609 ( .A(B[2]), .B(A[865]), .Z(\ab[865][2] ) );
  AND U610 ( .A(B[1]), .B(A[865]), .Z(\ab[865][1] ) );
  AND U611 ( .A(A[865]), .B(B[0]), .Z(\ab[865][0] ) );
  AND U612 ( .A(B[3]), .B(A[864]), .Z(\ab[864][3] ) );
  AND U613 ( .A(B[2]), .B(A[864]), .Z(\ab[864][2] ) );
  AND U614 ( .A(B[1]), .B(A[864]), .Z(\ab[864][1] ) );
  AND U615 ( .A(A[864]), .B(B[0]), .Z(\ab[864][0] ) );
  AND U616 ( .A(B[3]), .B(A[863]), .Z(\ab[863][3] ) );
  AND U617 ( .A(B[2]), .B(A[863]), .Z(\ab[863][2] ) );
  AND U618 ( .A(B[1]), .B(A[863]), .Z(\ab[863][1] ) );
  AND U619 ( .A(A[863]), .B(B[0]), .Z(\ab[863][0] ) );
  AND U620 ( .A(B[3]), .B(A[862]), .Z(\ab[862][3] ) );
  AND U621 ( .A(B[2]), .B(A[862]), .Z(\ab[862][2] ) );
  AND U622 ( .A(B[1]), .B(A[862]), .Z(\ab[862][1] ) );
  AND U623 ( .A(A[862]), .B(B[0]), .Z(\ab[862][0] ) );
  AND U624 ( .A(B[3]), .B(A[861]), .Z(\ab[861][3] ) );
  AND U625 ( .A(B[2]), .B(A[861]), .Z(\ab[861][2] ) );
  AND U626 ( .A(B[1]), .B(A[861]), .Z(\ab[861][1] ) );
  AND U627 ( .A(A[861]), .B(B[0]), .Z(\ab[861][0] ) );
  AND U628 ( .A(B[3]), .B(A[860]), .Z(\ab[860][3] ) );
  AND U629 ( .A(B[2]), .B(A[860]), .Z(\ab[860][2] ) );
  AND U630 ( .A(B[1]), .B(A[860]), .Z(\ab[860][1] ) );
  AND U631 ( .A(A[860]), .B(B[0]), .Z(\ab[860][0] ) );
  AND U632 ( .A(B[3]), .B(A[85]), .Z(\ab[85][3] ) );
  AND U633 ( .A(B[2]), .B(A[85]), .Z(\ab[85][2] ) );
  AND U634 ( .A(B[1]), .B(A[85]), .Z(\ab[85][1] ) );
  AND U635 ( .A(A[85]), .B(B[0]), .Z(\ab[85][0] ) );
  AND U636 ( .A(B[3]), .B(A[859]), .Z(\ab[859][3] ) );
  AND U637 ( .A(B[2]), .B(A[859]), .Z(\ab[859][2] ) );
  AND U638 ( .A(B[1]), .B(A[859]), .Z(\ab[859][1] ) );
  AND U639 ( .A(A[859]), .B(B[0]), .Z(\ab[859][0] ) );
  AND U640 ( .A(B[3]), .B(A[858]), .Z(\ab[858][3] ) );
  AND U641 ( .A(B[2]), .B(A[858]), .Z(\ab[858][2] ) );
  AND U642 ( .A(B[1]), .B(A[858]), .Z(\ab[858][1] ) );
  AND U643 ( .A(A[858]), .B(B[0]), .Z(\ab[858][0] ) );
  AND U644 ( .A(B[3]), .B(A[857]), .Z(\ab[857][3] ) );
  AND U645 ( .A(B[2]), .B(A[857]), .Z(\ab[857][2] ) );
  AND U646 ( .A(B[1]), .B(A[857]), .Z(\ab[857][1] ) );
  AND U647 ( .A(A[857]), .B(B[0]), .Z(\ab[857][0] ) );
  AND U648 ( .A(B[3]), .B(A[856]), .Z(\ab[856][3] ) );
  AND U649 ( .A(B[2]), .B(A[856]), .Z(\ab[856][2] ) );
  AND U650 ( .A(B[1]), .B(A[856]), .Z(\ab[856][1] ) );
  AND U651 ( .A(A[856]), .B(B[0]), .Z(\ab[856][0] ) );
  AND U652 ( .A(B[3]), .B(A[855]), .Z(\ab[855][3] ) );
  AND U653 ( .A(B[2]), .B(A[855]), .Z(\ab[855][2] ) );
  AND U654 ( .A(B[1]), .B(A[855]), .Z(\ab[855][1] ) );
  AND U655 ( .A(A[855]), .B(B[0]), .Z(\ab[855][0] ) );
  AND U656 ( .A(B[3]), .B(A[854]), .Z(\ab[854][3] ) );
  AND U657 ( .A(B[2]), .B(A[854]), .Z(\ab[854][2] ) );
  AND U658 ( .A(B[1]), .B(A[854]), .Z(\ab[854][1] ) );
  AND U659 ( .A(A[854]), .B(B[0]), .Z(\ab[854][0] ) );
  AND U660 ( .A(B[3]), .B(A[853]), .Z(\ab[853][3] ) );
  AND U661 ( .A(B[2]), .B(A[853]), .Z(\ab[853][2] ) );
  AND U662 ( .A(B[1]), .B(A[853]), .Z(\ab[853][1] ) );
  AND U663 ( .A(A[853]), .B(B[0]), .Z(\ab[853][0] ) );
  AND U664 ( .A(B[3]), .B(A[852]), .Z(\ab[852][3] ) );
  AND U665 ( .A(B[2]), .B(A[852]), .Z(\ab[852][2] ) );
  AND U666 ( .A(B[1]), .B(A[852]), .Z(\ab[852][1] ) );
  AND U667 ( .A(A[852]), .B(B[0]), .Z(\ab[852][0] ) );
  AND U668 ( .A(B[3]), .B(A[851]), .Z(\ab[851][3] ) );
  AND U669 ( .A(B[2]), .B(A[851]), .Z(\ab[851][2] ) );
  AND U670 ( .A(B[1]), .B(A[851]), .Z(\ab[851][1] ) );
  AND U671 ( .A(A[851]), .B(B[0]), .Z(\ab[851][0] ) );
  AND U672 ( .A(B[3]), .B(A[850]), .Z(\ab[850][3] ) );
  AND U673 ( .A(B[2]), .B(A[850]), .Z(\ab[850][2] ) );
  AND U674 ( .A(B[1]), .B(A[850]), .Z(\ab[850][1] ) );
  AND U675 ( .A(A[850]), .B(B[0]), .Z(\ab[850][0] ) );
  AND U676 ( .A(B[3]), .B(A[84]), .Z(\ab[84][3] ) );
  AND U677 ( .A(B[2]), .B(A[84]), .Z(\ab[84][2] ) );
  AND U678 ( .A(B[1]), .B(A[84]), .Z(\ab[84][1] ) );
  AND U679 ( .A(A[84]), .B(B[0]), .Z(\ab[84][0] ) );
  AND U680 ( .A(B[3]), .B(A[849]), .Z(\ab[849][3] ) );
  AND U681 ( .A(B[2]), .B(A[849]), .Z(\ab[849][2] ) );
  AND U682 ( .A(B[1]), .B(A[849]), .Z(\ab[849][1] ) );
  AND U683 ( .A(A[849]), .B(B[0]), .Z(\ab[849][0] ) );
  AND U684 ( .A(B[3]), .B(A[848]), .Z(\ab[848][3] ) );
  AND U685 ( .A(B[2]), .B(A[848]), .Z(\ab[848][2] ) );
  AND U686 ( .A(B[1]), .B(A[848]), .Z(\ab[848][1] ) );
  AND U687 ( .A(A[848]), .B(B[0]), .Z(\ab[848][0] ) );
  AND U688 ( .A(B[3]), .B(A[847]), .Z(\ab[847][3] ) );
  AND U689 ( .A(B[2]), .B(A[847]), .Z(\ab[847][2] ) );
  AND U690 ( .A(B[1]), .B(A[847]), .Z(\ab[847][1] ) );
  AND U691 ( .A(A[847]), .B(B[0]), .Z(\ab[847][0] ) );
  AND U692 ( .A(B[3]), .B(A[846]), .Z(\ab[846][3] ) );
  AND U693 ( .A(B[2]), .B(A[846]), .Z(\ab[846][2] ) );
  AND U694 ( .A(B[1]), .B(A[846]), .Z(\ab[846][1] ) );
  AND U695 ( .A(A[846]), .B(B[0]), .Z(\ab[846][0] ) );
  AND U696 ( .A(B[3]), .B(A[845]), .Z(\ab[845][3] ) );
  AND U697 ( .A(B[2]), .B(A[845]), .Z(\ab[845][2] ) );
  AND U698 ( .A(B[1]), .B(A[845]), .Z(\ab[845][1] ) );
  AND U699 ( .A(A[845]), .B(B[0]), .Z(\ab[845][0] ) );
  AND U700 ( .A(B[3]), .B(A[844]), .Z(\ab[844][3] ) );
  AND U701 ( .A(B[2]), .B(A[844]), .Z(\ab[844][2] ) );
  AND U702 ( .A(B[1]), .B(A[844]), .Z(\ab[844][1] ) );
  AND U703 ( .A(A[844]), .B(B[0]), .Z(\ab[844][0] ) );
  AND U704 ( .A(B[3]), .B(A[843]), .Z(\ab[843][3] ) );
  AND U705 ( .A(B[2]), .B(A[843]), .Z(\ab[843][2] ) );
  AND U706 ( .A(B[1]), .B(A[843]), .Z(\ab[843][1] ) );
  AND U707 ( .A(A[843]), .B(B[0]), .Z(\ab[843][0] ) );
  AND U708 ( .A(B[3]), .B(A[842]), .Z(\ab[842][3] ) );
  AND U709 ( .A(B[2]), .B(A[842]), .Z(\ab[842][2] ) );
  AND U710 ( .A(B[1]), .B(A[842]), .Z(\ab[842][1] ) );
  AND U711 ( .A(A[842]), .B(B[0]), .Z(\ab[842][0] ) );
  AND U712 ( .A(B[3]), .B(A[841]), .Z(\ab[841][3] ) );
  AND U713 ( .A(B[2]), .B(A[841]), .Z(\ab[841][2] ) );
  AND U714 ( .A(B[1]), .B(A[841]), .Z(\ab[841][1] ) );
  AND U715 ( .A(A[841]), .B(B[0]), .Z(\ab[841][0] ) );
  AND U716 ( .A(B[3]), .B(A[840]), .Z(\ab[840][3] ) );
  AND U717 ( .A(B[2]), .B(A[840]), .Z(\ab[840][2] ) );
  AND U718 ( .A(B[1]), .B(A[840]), .Z(\ab[840][1] ) );
  AND U719 ( .A(A[840]), .B(B[0]), .Z(\ab[840][0] ) );
  AND U720 ( .A(B[3]), .B(A[83]), .Z(\ab[83][3] ) );
  AND U721 ( .A(B[2]), .B(A[83]), .Z(\ab[83][2] ) );
  AND U722 ( .A(B[1]), .B(A[83]), .Z(\ab[83][1] ) );
  AND U723 ( .A(A[83]), .B(B[0]), .Z(\ab[83][0] ) );
  AND U724 ( .A(B[3]), .B(A[839]), .Z(\ab[839][3] ) );
  AND U725 ( .A(B[2]), .B(A[839]), .Z(\ab[839][2] ) );
  AND U726 ( .A(B[1]), .B(A[839]), .Z(\ab[839][1] ) );
  AND U727 ( .A(A[839]), .B(B[0]), .Z(\ab[839][0] ) );
  AND U728 ( .A(B[3]), .B(A[838]), .Z(\ab[838][3] ) );
  AND U729 ( .A(B[2]), .B(A[838]), .Z(\ab[838][2] ) );
  AND U730 ( .A(B[1]), .B(A[838]), .Z(\ab[838][1] ) );
  AND U731 ( .A(A[838]), .B(B[0]), .Z(\ab[838][0] ) );
  AND U732 ( .A(B[3]), .B(A[837]), .Z(\ab[837][3] ) );
  AND U733 ( .A(B[2]), .B(A[837]), .Z(\ab[837][2] ) );
  AND U734 ( .A(B[1]), .B(A[837]), .Z(\ab[837][1] ) );
  AND U735 ( .A(A[837]), .B(B[0]), .Z(\ab[837][0] ) );
  AND U736 ( .A(B[3]), .B(A[836]), .Z(\ab[836][3] ) );
  AND U737 ( .A(B[2]), .B(A[836]), .Z(\ab[836][2] ) );
  AND U738 ( .A(B[1]), .B(A[836]), .Z(\ab[836][1] ) );
  AND U739 ( .A(A[836]), .B(B[0]), .Z(\ab[836][0] ) );
  AND U740 ( .A(B[3]), .B(A[835]), .Z(\ab[835][3] ) );
  AND U741 ( .A(B[2]), .B(A[835]), .Z(\ab[835][2] ) );
  AND U742 ( .A(B[1]), .B(A[835]), .Z(\ab[835][1] ) );
  AND U743 ( .A(A[835]), .B(B[0]), .Z(\ab[835][0] ) );
  AND U744 ( .A(B[3]), .B(A[834]), .Z(\ab[834][3] ) );
  AND U745 ( .A(B[2]), .B(A[834]), .Z(\ab[834][2] ) );
  AND U746 ( .A(B[1]), .B(A[834]), .Z(\ab[834][1] ) );
  AND U747 ( .A(A[834]), .B(B[0]), .Z(\ab[834][0] ) );
  AND U748 ( .A(B[3]), .B(A[833]), .Z(\ab[833][3] ) );
  AND U749 ( .A(B[2]), .B(A[833]), .Z(\ab[833][2] ) );
  AND U750 ( .A(B[1]), .B(A[833]), .Z(\ab[833][1] ) );
  AND U751 ( .A(A[833]), .B(B[0]), .Z(\ab[833][0] ) );
  AND U752 ( .A(B[3]), .B(A[832]), .Z(\ab[832][3] ) );
  AND U753 ( .A(B[2]), .B(A[832]), .Z(\ab[832][2] ) );
  AND U754 ( .A(B[1]), .B(A[832]), .Z(\ab[832][1] ) );
  AND U755 ( .A(A[832]), .B(B[0]), .Z(\ab[832][0] ) );
  AND U756 ( .A(B[3]), .B(A[831]), .Z(\ab[831][3] ) );
  AND U757 ( .A(B[2]), .B(A[831]), .Z(\ab[831][2] ) );
  AND U758 ( .A(B[1]), .B(A[831]), .Z(\ab[831][1] ) );
  AND U759 ( .A(A[831]), .B(B[0]), .Z(\ab[831][0] ) );
  AND U760 ( .A(B[3]), .B(A[830]), .Z(\ab[830][3] ) );
  AND U761 ( .A(B[2]), .B(A[830]), .Z(\ab[830][2] ) );
  AND U762 ( .A(B[1]), .B(A[830]), .Z(\ab[830][1] ) );
  AND U763 ( .A(A[830]), .B(B[0]), .Z(\ab[830][0] ) );
  AND U764 ( .A(B[3]), .B(A[82]), .Z(\ab[82][3] ) );
  AND U765 ( .A(B[2]), .B(A[82]), .Z(\ab[82][2] ) );
  AND U766 ( .A(B[1]), .B(A[82]), .Z(\ab[82][1] ) );
  AND U767 ( .A(A[82]), .B(B[0]), .Z(\ab[82][0] ) );
  AND U768 ( .A(B[3]), .B(A[829]), .Z(\ab[829][3] ) );
  AND U769 ( .A(B[2]), .B(A[829]), .Z(\ab[829][2] ) );
  AND U770 ( .A(B[1]), .B(A[829]), .Z(\ab[829][1] ) );
  AND U771 ( .A(A[829]), .B(B[0]), .Z(\ab[829][0] ) );
  AND U772 ( .A(B[3]), .B(A[828]), .Z(\ab[828][3] ) );
  AND U773 ( .A(B[2]), .B(A[828]), .Z(\ab[828][2] ) );
  AND U774 ( .A(B[1]), .B(A[828]), .Z(\ab[828][1] ) );
  AND U775 ( .A(A[828]), .B(B[0]), .Z(\ab[828][0] ) );
  AND U776 ( .A(B[3]), .B(A[827]), .Z(\ab[827][3] ) );
  AND U777 ( .A(B[2]), .B(A[827]), .Z(\ab[827][2] ) );
  AND U778 ( .A(B[1]), .B(A[827]), .Z(\ab[827][1] ) );
  AND U779 ( .A(A[827]), .B(B[0]), .Z(\ab[827][0] ) );
  AND U780 ( .A(B[3]), .B(A[826]), .Z(\ab[826][3] ) );
  AND U781 ( .A(B[2]), .B(A[826]), .Z(\ab[826][2] ) );
  AND U782 ( .A(B[1]), .B(A[826]), .Z(\ab[826][1] ) );
  AND U783 ( .A(A[826]), .B(B[0]), .Z(\ab[826][0] ) );
  AND U784 ( .A(B[3]), .B(A[825]), .Z(\ab[825][3] ) );
  AND U785 ( .A(B[2]), .B(A[825]), .Z(\ab[825][2] ) );
  AND U786 ( .A(B[1]), .B(A[825]), .Z(\ab[825][1] ) );
  AND U787 ( .A(A[825]), .B(B[0]), .Z(\ab[825][0] ) );
  AND U788 ( .A(B[3]), .B(A[824]), .Z(\ab[824][3] ) );
  AND U789 ( .A(B[2]), .B(A[824]), .Z(\ab[824][2] ) );
  AND U790 ( .A(B[1]), .B(A[824]), .Z(\ab[824][1] ) );
  AND U791 ( .A(A[824]), .B(B[0]), .Z(\ab[824][0] ) );
  AND U792 ( .A(B[3]), .B(A[823]), .Z(\ab[823][3] ) );
  AND U793 ( .A(B[2]), .B(A[823]), .Z(\ab[823][2] ) );
  AND U794 ( .A(B[1]), .B(A[823]), .Z(\ab[823][1] ) );
  AND U795 ( .A(A[823]), .B(B[0]), .Z(\ab[823][0] ) );
  AND U796 ( .A(B[3]), .B(A[822]), .Z(\ab[822][3] ) );
  AND U797 ( .A(B[2]), .B(A[822]), .Z(\ab[822][2] ) );
  AND U798 ( .A(B[1]), .B(A[822]), .Z(\ab[822][1] ) );
  AND U799 ( .A(A[822]), .B(B[0]), .Z(\ab[822][0] ) );
  AND U800 ( .A(B[3]), .B(A[821]), .Z(\ab[821][3] ) );
  AND U801 ( .A(B[2]), .B(A[821]), .Z(\ab[821][2] ) );
  AND U802 ( .A(B[1]), .B(A[821]), .Z(\ab[821][1] ) );
  AND U803 ( .A(A[821]), .B(B[0]), .Z(\ab[821][0] ) );
  AND U804 ( .A(B[3]), .B(A[820]), .Z(\ab[820][3] ) );
  AND U805 ( .A(B[2]), .B(A[820]), .Z(\ab[820][2] ) );
  AND U806 ( .A(B[1]), .B(A[820]), .Z(\ab[820][1] ) );
  AND U807 ( .A(A[820]), .B(B[0]), .Z(\ab[820][0] ) );
  AND U808 ( .A(B[3]), .B(A[81]), .Z(\ab[81][3] ) );
  AND U809 ( .A(B[2]), .B(A[81]), .Z(\ab[81][2] ) );
  AND U810 ( .A(B[1]), .B(A[81]), .Z(\ab[81][1] ) );
  AND U811 ( .A(A[81]), .B(B[0]), .Z(\ab[81][0] ) );
  AND U812 ( .A(B[3]), .B(A[819]), .Z(\ab[819][3] ) );
  AND U813 ( .A(B[2]), .B(A[819]), .Z(\ab[819][2] ) );
  AND U814 ( .A(B[1]), .B(A[819]), .Z(\ab[819][1] ) );
  AND U815 ( .A(A[819]), .B(B[0]), .Z(\ab[819][0] ) );
  AND U816 ( .A(B[3]), .B(A[818]), .Z(\ab[818][3] ) );
  AND U817 ( .A(B[2]), .B(A[818]), .Z(\ab[818][2] ) );
  AND U818 ( .A(B[1]), .B(A[818]), .Z(\ab[818][1] ) );
  AND U819 ( .A(A[818]), .B(B[0]), .Z(\ab[818][0] ) );
  AND U820 ( .A(B[3]), .B(A[817]), .Z(\ab[817][3] ) );
  AND U821 ( .A(B[2]), .B(A[817]), .Z(\ab[817][2] ) );
  AND U822 ( .A(B[1]), .B(A[817]), .Z(\ab[817][1] ) );
  AND U823 ( .A(A[817]), .B(B[0]), .Z(\ab[817][0] ) );
  AND U824 ( .A(B[3]), .B(A[816]), .Z(\ab[816][3] ) );
  AND U825 ( .A(B[2]), .B(A[816]), .Z(\ab[816][2] ) );
  AND U826 ( .A(B[1]), .B(A[816]), .Z(\ab[816][1] ) );
  AND U827 ( .A(A[816]), .B(B[0]), .Z(\ab[816][0] ) );
  AND U828 ( .A(B[3]), .B(A[815]), .Z(\ab[815][3] ) );
  AND U829 ( .A(B[2]), .B(A[815]), .Z(\ab[815][2] ) );
  AND U830 ( .A(B[1]), .B(A[815]), .Z(\ab[815][1] ) );
  AND U831 ( .A(A[815]), .B(B[0]), .Z(\ab[815][0] ) );
  AND U832 ( .A(B[3]), .B(A[814]), .Z(\ab[814][3] ) );
  AND U833 ( .A(B[2]), .B(A[814]), .Z(\ab[814][2] ) );
  AND U834 ( .A(B[1]), .B(A[814]), .Z(\ab[814][1] ) );
  AND U835 ( .A(A[814]), .B(B[0]), .Z(\ab[814][0] ) );
  AND U836 ( .A(B[3]), .B(A[813]), .Z(\ab[813][3] ) );
  AND U837 ( .A(B[2]), .B(A[813]), .Z(\ab[813][2] ) );
  AND U838 ( .A(B[1]), .B(A[813]), .Z(\ab[813][1] ) );
  AND U839 ( .A(A[813]), .B(B[0]), .Z(\ab[813][0] ) );
  AND U840 ( .A(B[3]), .B(A[812]), .Z(\ab[812][3] ) );
  AND U841 ( .A(B[2]), .B(A[812]), .Z(\ab[812][2] ) );
  AND U842 ( .A(B[1]), .B(A[812]), .Z(\ab[812][1] ) );
  AND U843 ( .A(A[812]), .B(B[0]), .Z(\ab[812][0] ) );
  AND U844 ( .A(B[3]), .B(A[811]), .Z(\ab[811][3] ) );
  AND U845 ( .A(B[2]), .B(A[811]), .Z(\ab[811][2] ) );
  AND U846 ( .A(B[1]), .B(A[811]), .Z(\ab[811][1] ) );
  AND U847 ( .A(A[811]), .B(B[0]), .Z(\ab[811][0] ) );
  AND U848 ( .A(B[3]), .B(A[810]), .Z(\ab[810][3] ) );
  AND U849 ( .A(B[2]), .B(A[810]), .Z(\ab[810][2] ) );
  AND U850 ( .A(B[1]), .B(A[810]), .Z(\ab[810][1] ) );
  AND U851 ( .A(A[810]), .B(B[0]), .Z(\ab[810][0] ) );
  AND U852 ( .A(B[3]), .B(A[80]), .Z(\ab[80][3] ) );
  AND U853 ( .A(B[2]), .B(A[80]), .Z(\ab[80][2] ) );
  AND U854 ( .A(B[1]), .B(A[80]), .Z(\ab[80][1] ) );
  AND U855 ( .A(A[80]), .B(B[0]), .Z(\ab[80][0] ) );
  AND U856 ( .A(B[3]), .B(A[809]), .Z(\ab[809][3] ) );
  AND U857 ( .A(B[2]), .B(A[809]), .Z(\ab[809][2] ) );
  AND U858 ( .A(B[1]), .B(A[809]), .Z(\ab[809][1] ) );
  AND U859 ( .A(A[809]), .B(B[0]), .Z(\ab[809][0] ) );
  AND U860 ( .A(B[3]), .B(A[808]), .Z(\ab[808][3] ) );
  AND U861 ( .A(B[2]), .B(A[808]), .Z(\ab[808][2] ) );
  AND U862 ( .A(B[1]), .B(A[808]), .Z(\ab[808][1] ) );
  AND U863 ( .A(A[808]), .B(B[0]), .Z(\ab[808][0] ) );
  AND U864 ( .A(B[3]), .B(A[807]), .Z(\ab[807][3] ) );
  AND U865 ( .A(B[2]), .B(A[807]), .Z(\ab[807][2] ) );
  AND U866 ( .A(B[1]), .B(A[807]), .Z(\ab[807][1] ) );
  AND U867 ( .A(A[807]), .B(B[0]), .Z(\ab[807][0] ) );
  AND U868 ( .A(B[3]), .B(A[806]), .Z(\ab[806][3] ) );
  AND U869 ( .A(B[2]), .B(A[806]), .Z(\ab[806][2] ) );
  AND U870 ( .A(B[1]), .B(A[806]), .Z(\ab[806][1] ) );
  AND U871 ( .A(A[806]), .B(B[0]), .Z(\ab[806][0] ) );
  AND U872 ( .A(B[3]), .B(A[805]), .Z(\ab[805][3] ) );
  AND U873 ( .A(B[2]), .B(A[805]), .Z(\ab[805][2] ) );
  AND U874 ( .A(B[1]), .B(A[805]), .Z(\ab[805][1] ) );
  AND U875 ( .A(A[805]), .B(B[0]), .Z(\ab[805][0] ) );
  AND U876 ( .A(B[3]), .B(A[804]), .Z(\ab[804][3] ) );
  AND U877 ( .A(B[2]), .B(A[804]), .Z(\ab[804][2] ) );
  AND U878 ( .A(B[1]), .B(A[804]), .Z(\ab[804][1] ) );
  AND U879 ( .A(A[804]), .B(B[0]), .Z(\ab[804][0] ) );
  AND U880 ( .A(B[3]), .B(A[803]), .Z(\ab[803][3] ) );
  AND U881 ( .A(B[2]), .B(A[803]), .Z(\ab[803][2] ) );
  AND U882 ( .A(B[1]), .B(A[803]), .Z(\ab[803][1] ) );
  AND U883 ( .A(A[803]), .B(B[0]), .Z(\ab[803][0] ) );
  AND U884 ( .A(B[3]), .B(A[802]), .Z(\ab[802][3] ) );
  AND U885 ( .A(B[2]), .B(A[802]), .Z(\ab[802][2] ) );
  AND U886 ( .A(B[1]), .B(A[802]), .Z(\ab[802][1] ) );
  AND U887 ( .A(A[802]), .B(B[0]), .Z(\ab[802][0] ) );
  AND U888 ( .A(B[3]), .B(A[801]), .Z(\ab[801][3] ) );
  AND U889 ( .A(B[2]), .B(A[801]), .Z(\ab[801][2] ) );
  AND U890 ( .A(B[1]), .B(A[801]), .Z(\ab[801][1] ) );
  AND U891 ( .A(A[801]), .B(B[0]), .Z(\ab[801][0] ) );
  AND U892 ( .A(B[3]), .B(A[800]), .Z(\ab[800][3] ) );
  AND U893 ( .A(B[2]), .B(A[800]), .Z(\ab[800][2] ) );
  AND U894 ( .A(B[1]), .B(A[800]), .Z(\ab[800][1] ) );
  AND U895 ( .A(A[800]), .B(B[0]), .Z(\ab[800][0] ) );
  AND U896 ( .A(B[3]), .B(A[7]), .Z(\ab[7][3] ) );
  AND U897 ( .A(B[2]), .B(A[7]), .Z(\ab[7][2] ) );
  AND U898 ( .A(B[1]), .B(A[7]), .Z(\ab[7][1] ) );
  AND U899 ( .A(A[7]), .B(B[0]), .Z(\ab[7][0] ) );
  AND U900 ( .A(B[3]), .B(A[79]), .Z(\ab[79][3] ) );
  AND U901 ( .A(B[2]), .B(A[79]), .Z(\ab[79][2] ) );
  AND U902 ( .A(B[1]), .B(A[79]), .Z(\ab[79][1] ) );
  AND U903 ( .A(A[79]), .B(B[0]), .Z(\ab[79][0] ) );
  AND U904 ( .A(B[3]), .B(A[799]), .Z(\ab[799][3] ) );
  AND U905 ( .A(B[2]), .B(A[799]), .Z(\ab[799][2] ) );
  AND U906 ( .A(B[1]), .B(A[799]), .Z(\ab[799][1] ) );
  AND U907 ( .A(A[799]), .B(B[0]), .Z(\ab[799][0] ) );
  AND U908 ( .A(B[3]), .B(A[798]), .Z(\ab[798][3] ) );
  AND U909 ( .A(B[2]), .B(A[798]), .Z(\ab[798][2] ) );
  AND U910 ( .A(B[1]), .B(A[798]), .Z(\ab[798][1] ) );
  AND U911 ( .A(A[798]), .B(B[0]), .Z(\ab[798][0] ) );
  AND U912 ( .A(B[3]), .B(A[797]), .Z(\ab[797][3] ) );
  AND U913 ( .A(B[2]), .B(A[797]), .Z(\ab[797][2] ) );
  AND U914 ( .A(B[1]), .B(A[797]), .Z(\ab[797][1] ) );
  AND U915 ( .A(A[797]), .B(B[0]), .Z(\ab[797][0] ) );
  AND U916 ( .A(B[3]), .B(A[796]), .Z(\ab[796][3] ) );
  AND U917 ( .A(B[2]), .B(A[796]), .Z(\ab[796][2] ) );
  AND U918 ( .A(B[1]), .B(A[796]), .Z(\ab[796][1] ) );
  AND U919 ( .A(A[796]), .B(B[0]), .Z(\ab[796][0] ) );
  AND U920 ( .A(B[3]), .B(A[795]), .Z(\ab[795][3] ) );
  AND U921 ( .A(B[2]), .B(A[795]), .Z(\ab[795][2] ) );
  AND U922 ( .A(B[1]), .B(A[795]), .Z(\ab[795][1] ) );
  AND U923 ( .A(A[795]), .B(B[0]), .Z(\ab[795][0] ) );
  AND U924 ( .A(B[3]), .B(A[794]), .Z(\ab[794][3] ) );
  AND U925 ( .A(B[2]), .B(A[794]), .Z(\ab[794][2] ) );
  AND U926 ( .A(B[1]), .B(A[794]), .Z(\ab[794][1] ) );
  AND U927 ( .A(A[794]), .B(B[0]), .Z(\ab[794][0] ) );
  AND U928 ( .A(B[3]), .B(A[793]), .Z(\ab[793][3] ) );
  AND U929 ( .A(B[2]), .B(A[793]), .Z(\ab[793][2] ) );
  AND U930 ( .A(B[1]), .B(A[793]), .Z(\ab[793][1] ) );
  AND U931 ( .A(A[793]), .B(B[0]), .Z(\ab[793][0] ) );
  AND U932 ( .A(B[3]), .B(A[792]), .Z(\ab[792][3] ) );
  AND U933 ( .A(B[2]), .B(A[792]), .Z(\ab[792][2] ) );
  AND U934 ( .A(B[1]), .B(A[792]), .Z(\ab[792][1] ) );
  AND U935 ( .A(A[792]), .B(B[0]), .Z(\ab[792][0] ) );
  AND U936 ( .A(B[3]), .B(A[791]), .Z(\ab[791][3] ) );
  AND U937 ( .A(B[2]), .B(A[791]), .Z(\ab[791][2] ) );
  AND U938 ( .A(B[1]), .B(A[791]), .Z(\ab[791][1] ) );
  AND U939 ( .A(A[791]), .B(B[0]), .Z(\ab[791][0] ) );
  AND U940 ( .A(B[3]), .B(A[790]), .Z(\ab[790][3] ) );
  AND U941 ( .A(B[2]), .B(A[790]), .Z(\ab[790][2] ) );
  AND U942 ( .A(B[1]), .B(A[790]), .Z(\ab[790][1] ) );
  AND U943 ( .A(A[790]), .B(B[0]), .Z(\ab[790][0] ) );
  AND U944 ( .A(B[3]), .B(A[78]), .Z(\ab[78][3] ) );
  AND U945 ( .A(B[2]), .B(A[78]), .Z(\ab[78][2] ) );
  AND U946 ( .A(B[1]), .B(A[78]), .Z(\ab[78][1] ) );
  AND U947 ( .A(A[78]), .B(B[0]), .Z(\ab[78][0] ) );
  AND U948 ( .A(B[3]), .B(A[789]), .Z(\ab[789][3] ) );
  AND U949 ( .A(B[2]), .B(A[789]), .Z(\ab[789][2] ) );
  AND U950 ( .A(B[1]), .B(A[789]), .Z(\ab[789][1] ) );
  AND U951 ( .A(A[789]), .B(B[0]), .Z(\ab[789][0] ) );
  AND U952 ( .A(B[3]), .B(A[788]), .Z(\ab[788][3] ) );
  AND U953 ( .A(B[2]), .B(A[788]), .Z(\ab[788][2] ) );
  AND U954 ( .A(B[1]), .B(A[788]), .Z(\ab[788][1] ) );
  AND U955 ( .A(A[788]), .B(B[0]), .Z(\ab[788][0] ) );
  AND U956 ( .A(B[3]), .B(A[787]), .Z(\ab[787][3] ) );
  AND U957 ( .A(B[2]), .B(A[787]), .Z(\ab[787][2] ) );
  AND U958 ( .A(B[1]), .B(A[787]), .Z(\ab[787][1] ) );
  AND U959 ( .A(A[787]), .B(B[0]), .Z(\ab[787][0] ) );
  AND U960 ( .A(B[3]), .B(A[786]), .Z(\ab[786][3] ) );
  AND U961 ( .A(B[2]), .B(A[786]), .Z(\ab[786][2] ) );
  AND U962 ( .A(B[1]), .B(A[786]), .Z(\ab[786][1] ) );
  AND U963 ( .A(A[786]), .B(B[0]), .Z(\ab[786][0] ) );
  AND U964 ( .A(B[3]), .B(A[785]), .Z(\ab[785][3] ) );
  AND U965 ( .A(B[2]), .B(A[785]), .Z(\ab[785][2] ) );
  AND U966 ( .A(B[1]), .B(A[785]), .Z(\ab[785][1] ) );
  AND U967 ( .A(A[785]), .B(B[0]), .Z(\ab[785][0] ) );
  AND U968 ( .A(B[3]), .B(A[784]), .Z(\ab[784][3] ) );
  AND U969 ( .A(B[2]), .B(A[784]), .Z(\ab[784][2] ) );
  AND U970 ( .A(B[1]), .B(A[784]), .Z(\ab[784][1] ) );
  AND U971 ( .A(A[784]), .B(B[0]), .Z(\ab[784][0] ) );
  AND U972 ( .A(B[3]), .B(A[783]), .Z(\ab[783][3] ) );
  AND U973 ( .A(B[2]), .B(A[783]), .Z(\ab[783][2] ) );
  AND U974 ( .A(B[1]), .B(A[783]), .Z(\ab[783][1] ) );
  AND U975 ( .A(A[783]), .B(B[0]), .Z(\ab[783][0] ) );
  AND U976 ( .A(B[3]), .B(A[782]), .Z(\ab[782][3] ) );
  AND U977 ( .A(B[2]), .B(A[782]), .Z(\ab[782][2] ) );
  AND U978 ( .A(B[1]), .B(A[782]), .Z(\ab[782][1] ) );
  AND U979 ( .A(A[782]), .B(B[0]), .Z(\ab[782][0] ) );
  AND U980 ( .A(B[3]), .B(A[781]), .Z(\ab[781][3] ) );
  AND U981 ( .A(B[2]), .B(A[781]), .Z(\ab[781][2] ) );
  AND U982 ( .A(B[1]), .B(A[781]), .Z(\ab[781][1] ) );
  AND U983 ( .A(A[781]), .B(B[0]), .Z(\ab[781][0] ) );
  AND U984 ( .A(B[3]), .B(A[780]), .Z(\ab[780][3] ) );
  AND U985 ( .A(B[2]), .B(A[780]), .Z(\ab[780][2] ) );
  AND U986 ( .A(B[1]), .B(A[780]), .Z(\ab[780][1] ) );
  AND U987 ( .A(A[780]), .B(B[0]), .Z(\ab[780][0] ) );
  AND U988 ( .A(B[3]), .B(A[77]), .Z(\ab[77][3] ) );
  AND U989 ( .A(B[2]), .B(A[77]), .Z(\ab[77][2] ) );
  AND U990 ( .A(B[1]), .B(A[77]), .Z(\ab[77][1] ) );
  AND U991 ( .A(A[77]), .B(B[0]), .Z(\ab[77][0] ) );
  AND U992 ( .A(B[3]), .B(A[779]), .Z(\ab[779][3] ) );
  AND U993 ( .A(B[2]), .B(A[779]), .Z(\ab[779][2] ) );
  AND U994 ( .A(B[1]), .B(A[779]), .Z(\ab[779][1] ) );
  AND U995 ( .A(A[779]), .B(B[0]), .Z(\ab[779][0] ) );
  AND U996 ( .A(B[3]), .B(A[778]), .Z(\ab[778][3] ) );
  AND U997 ( .A(B[2]), .B(A[778]), .Z(\ab[778][2] ) );
  AND U998 ( .A(B[1]), .B(A[778]), .Z(\ab[778][1] ) );
  AND U999 ( .A(A[778]), .B(B[0]), .Z(\ab[778][0] ) );
  AND U1000 ( .A(B[3]), .B(A[777]), .Z(\ab[777][3] ) );
  AND U1001 ( .A(B[2]), .B(A[777]), .Z(\ab[777][2] ) );
  AND U1002 ( .A(B[1]), .B(A[777]), .Z(\ab[777][1] ) );
  AND U1003 ( .A(A[777]), .B(B[0]), .Z(\ab[777][0] ) );
  AND U1004 ( .A(B[3]), .B(A[776]), .Z(\ab[776][3] ) );
  AND U1005 ( .A(B[2]), .B(A[776]), .Z(\ab[776][2] ) );
  AND U1006 ( .A(B[1]), .B(A[776]), .Z(\ab[776][1] ) );
  AND U1007 ( .A(A[776]), .B(B[0]), .Z(\ab[776][0] ) );
  AND U1008 ( .A(B[3]), .B(A[775]), .Z(\ab[775][3] ) );
  AND U1009 ( .A(B[2]), .B(A[775]), .Z(\ab[775][2] ) );
  AND U1010 ( .A(B[1]), .B(A[775]), .Z(\ab[775][1] ) );
  AND U1011 ( .A(A[775]), .B(B[0]), .Z(\ab[775][0] ) );
  AND U1012 ( .A(B[3]), .B(A[774]), .Z(\ab[774][3] ) );
  AND U1013 ( .A(B[2]), .B(A[774]), .Z(\ab[774][2] ) );
  AND U1014 ( .A(B[1]), .B(A[774]), .Z(\ab[774][1] ) );
  AND U1015 ( .A(A[774]), .B(B[0]), .Z(\ab[774][0] ) );
  AND U1016 ( .A(B[3]), .B(A[773]), .Z(\ab[773][3] ) );
  AND U1017 ( .A(B[2]), .B(A[773]), .Z(\ab[773][2] ) );
  AND U1018 ( .A(B[1]), .B(A[773]), .Z(\ab[773][1] ) );
  AND U1019 ( .A(A[773]), .B(B[0]), .Z(\ab[773][0] ) );
  AND U1020 ( .A(B[3]), .B(A[772]), .Z(\ab[772][3] ) );
  AND U1021 ( .A(B[2]), .B(A[772]), .Z(\ab[772][2] ) );
  AND U1022 ( .A(B[1]), .B(A[772]), .Z(\ab[772][1] ) );
  AND U1023 ( .A(A[772]), .B(B[0]), .Z(\ab[772][0] ) );
  AND U1024 ( .A(B[3]), .B(A[771]), .Z(\ab[771][3] ) );
  AND U1025 ( .A(B[2]), .B(A[771]), .Z(\ab[771][2] ) );
  AND U1026 ( .A(B[1]), .B(A[771]), .Z(\ab[771][1] ) );
  AND U1027 ( .A(A[771]), .B(B[0]), .Z(\ab[771][0] ) );
  AND U1028 ( .A(B[3]), .B(A[770]), .Z(\ab[770][3] ) );
  AND U1029 ( .A(B[2]), .B(A[770]), .Z(\ab[770][2] ) );
  AND U1030 ( .A(B[1]), .B(A[770]), .Z(\ab[770][1] ) );
  AND U1031 ( .A(A[770]), .B(B[0]), .Z(\ab[770][0] ) );
  AND U1032 ( .A(B[3]), .B(A[76]), .Z(\ab[76][3] ) );
  AND U1033 ( .A(B[2]), .B(A[76]), .Z(\ab[76][2] ) );
  AND U1034 ( .A(B[1]), .B(A[76]), .Z(\ab[76][1] ) );
  AND U1035 ( .A(A[76]), .B(B[0]), .Z(\ab[76][0] ) );
  AND U1036 ( .A(B[3]), .B(A[769]), .Z(\ab[769][3] ) );
  AND U1037 ( .A(B[2]), .B(A[769]), .Z(\ab[769][2] ) );
  AND U1038 ( .A(B[1]), .B(A[769]), .Z(\ab[769][1] ) );
  AND U1039 ( .A(A[769]), .B(B[0]), .Z(\ab[769][0] ) );
  AND U1040 ( .A(B[3]), .B(A[768]), .Z(\ab[768][3] ) );
  AND U1041 ( .A(B[2]), .B(A[768]), .Z(\ab[768][2] ) );
  AND U1042 ( .A(B[1]), .B(A[768]), .Z(\ab[768][1] ) );
  AND U1043 ( .A(A[768]), .B(B[0]), .Z(\ab[768][0] ) );
  AND U1044 ( .A(B[3]), .B(A[767]), .Z(\ab[767][3] ) );
  AND U1045 ( .A(B[2]), .B(A[767]), .Z(\ab[767][2] ) );
  AND U1046 ( .A(B[1]), .B(A[767]), .Z(\ab[767][1] ) );
  AND U1047 ( .A(A[767]), .B(B[0]), .Z(\ab[767][0] ) );
  AND U1048 ( .A(B[3]), .B(A[766]), .Z(\ab[766][3] ) );
  AND U1049 ( .A(B[2]), .B(A[766]), .Z(\ab[766][2] ) );
  AND U1050 ( .A(B[1]), .B(A[766]), .Z(\ab[766][1] ) );
  AND U1051 ( .A(A[766]), .B(B[0]), .Z(\ab[766][0] ) );
  AND U1052 ( .A(B[3]), .B(A[765]), .Z(\ab[765][3] ) );
  AND U1053 ( .A(B[2]), .B(A[765]), .Z(\ab[765][2] ) );
  AND U1054 ( .A(B[1]), .B(A[765]), .Z(\ab[765][1] ) );
  AND U1055 ( .A(A[765]), .B(B[0]), .Z(\ab[765][0] ) );
  AND U1056 ( .A(B[3]), .B(A[764]), .Z(\ab[764][3] ) );
  AND U1057 ( .A(B[2]), .B(A[764]), .Z(\ab[764][2] ) );
  AND U1058 ( .A(B[1]), .B(A[764]), .Z(\ab[764][1] ) );
  AND U1059 ( .A(A[764]), .B(B[0]), .Z(\ab[764][0] ) );
  AND U1060 ( .A(B[3]), .B(A[763]), .Z(\ab[763][3] ) );
  AND U1061 ( .A(B[2]), .B(A[763]), .Z(\ab[763][2] ) );
  AND U1062 ( .A(B[1]), .B(A[763]), .Z(\ab[763][1] ) );
  AND U1063 ( .A(A[763]), .B(B[0]), .Z(\ab[763][0] ) );
  AND U1064 ( .A(B[3]), .B(A[762]), .Z(\ab[762][3] ) );
  AND U1065 ( .A(B[2]), .B(A[762]), .Z(\ab[762][2] ) );
  AND U1066 ( .A(B[1]), .B(A[762]), .Z(\ab[762][1] ) );
  AND U1067 ( .A(A[762]), .B(B[0]), .Z(\ab[762][0] ) );
  AND U1068 ( .A(B[3]), .B(A[761]), .Z(\ab[761][3] ) );
  AND U1069 ( .A(B[2]), .B(A[761]), .Z(\ab[761][2] ) );
  AND U1070 ( .A(B[1]), .B(A[761]), .Z(\ab[761][1] ) );
  AND U1071 ( .A(A[761]), .B(B[0]), .Z(\ab[761][0] ) );
  AND U1072 ( .A(B[3]), .B(A[760]), .Z(\ab[760][3] ) );
  AND U1073 ( .A(B[2]), .B(A[760]), .Z(\ab[760][2] ) );
  AND U1074 ( .A(B[1]), .B(A[760]), .Z(\ab[760][1] ) );
  AND U1075 ( .A(A[760]), .B(B[0]), .Z(\ab[760][0] ) );
  AND U1076 ( .A(B[3]), .B(A[75]), .Z(\ab[75][3] ) );
  AND U1077 ( .A(B[2]), .B(A[75]), .Z(\ab[75][2] ) );
  AND U1078 ( .A(B[1]), .B(A[75]), .Z(\ab[75][1] ) );
  AND U1079 ( .A(A[75]), .B(B[0]), .Z(\ab[75][0] ) );
  AND U1080 ( .A(B[3]), .B(A[759]), .Z(\ab[759][3] ) );
  AND U1081 ( .A(B[2]), .B(A[759]), .Z(\ab[759][2] ) );
  AND U1082 ( .A(B[1]), .B(A[759]), .Z(\ab[759][1] ) );
  AND U1083 ( .A(A[759]), .B(B[0]), .Z(\ab[759][0] ) );
  AND U1084 ( .A(B[3]), .B(A[758]), .Z(\ab[758][3] ) );
  AND U1085 ( .A(B[2]), .B(A[758]), .Z(\ab[758][2] ) );
  AND U1086 ( .A(B[1]), .B(A[758]), .Z(\ab[758][1] ) );
  AND U1087 ( .A(A[758]), .B(B[0]), .Z(\ab[758][0] ) );
  AND U1088 ( .A(B[3]), .B(A[757]), .Z(\ab[757][3] ) );
  AND U1089 ( .A(B[2]), .B(A[757]), .Z(\ab[757][2] ) );
  AND U1090 ( .A(B[1]), .B(A[757]), .Z(\ab[757][1] ) );
  AND U1091 ( .A(A[757]), .B(B[0]), .Z(\ab[757][0] ) );
  AND U1092 ( .A(B[3]), .B(A[756]), .Z(\ab[756][3] ) );
  AND U1093 ( .A(B[2]), .B(A[756]), .Z(\ab[756][2] ) );
  AND U1094 ( .A(B[1]), .B(A[756]), .Z(\ab[756][1] ) );
  AND U1095 ( .A(A[756]), .B(B[0]), .Z(\ab[756][0] ) );
  AND U1096 ( .A(B[3]), .B(A[755]), .Z(\ab[755][3] ) );
  AND U1097 ( .A(B[2]), .B(A[755]), .Z(\ab[755][2] ) );
  AND U1098 ( .A(B[1]), .B(A[755]), .Z(\ab[755][1] ) );
  AND U1099 ( .A(A[755]), .B(B[0]), .Z(\ab[755][0] ) );
  AND U1100 ( .A(B[3]), .B(A[754]), .Z(\ab[754][3] ) );
  AND U1101 ( .A(B[2]), .B(A[754]), .Z(\ab[754][2] ) );
  AND U1102 ( .A(B[1]), .B(A[754]), .Z(\ab[754][1] ) );
  AND U1103 ( .A(A[754]), .B(B[0]), .Z(\ab[754][0] ) );
  AND U1104 ( .A(B[3]), .B(A[753]), .Z(\ab[753][3] ) );
  AND U1105 ( .A(B[2]), .B(A[753]), .Z(\ab[753][2] ) );
  AND U1106 ( .A(B[1]), .B(A[753]), .Z(\ab[753][1] ) );
  AND U1107 ( .A(A[753]), .B(B[0]), .Z(\ab[753][0] ) );
  AND U1108 ( .A(B[3]), .B(A[752]), .Z(\ab[752][3] ) );
  AND U1109 ( .A(B[2]), .B(A[752]), .Z(\ab[752][2] ) );
  AND U1110 ( .A(B[1]), .B(A[752]), .Z(\ab[752][1] ) );
  AND U1111 ( .A(A[752]), .B(B[0]), .Z(\ab[752][0] ) );
  AND U1112 ( .A(B[3]), .B(A[751]), .Z(\ab[751][3] ) );
  AND U1113 ( .A(B[2]), .B(A[751]), .Z(\ab[751][2] ) );
  AND U1114 ( .A(B[1]), .B(A[751]), .Z(\ab[751][1] ) );
  AND U1115 ( .A(A[751]), .B(B[0]), .Z(\ab[751][0] ) );
  AND U1116 ( .A(B[3]), .B(A[750]), .Z(\ab[750][3] ) );
  AND U1117 ( .A(B[2]), .B(A[750]), .Z(\ab[750][2] ) );
  AND U1118 ( .A(B[1]), .B(A[750]), .Z(\ab[750][1] ) );
  AND U1119 ( .A(A[750]), .B(B[0]), .Z(\ab[750][0] ) );
  AND U1120 ( .A(B[3]), .B(A[74]), .Z(\ab[74][3] ) );
  AND U1121 ( .A(B[2]), .B(A[74]), .Z(\ab[74][2] ) );
  AND U1122 ( .A(B[1]), .B(A[74]), .Z(\ab[74][1] ) );
  AND U1123 ( .A(A[74]), .B(B[0]), .Z(\ab[74][0] ) );
  AND U1124 ( .A(B[3]), .B(A[749]), .Z(\ab[749][3] ) );
  AND U1125 ( .A(B[2]), .B(A[749]), .Z(\ab[749][2] ) );
  AND U1126 ( .A(B[1]), .B(A[749]), .Z(\ab[749][1] ) );
  AND U1127 ( .A(A[749]), .B(B[0]), .Z(\ab[749][0] ) );
  AND U1128 ( .A(B[3]), .B(A[748]), .Z(\ab[748][3] ) );
  AND U1129 ( .A(B[2]), .B(A[748]), .Z(\ab[748][2] ) );
  AND U1130 ( .A(B[1]), .B(A[748]), .Z(\ab[748][1] ) );
  AND U1131 ( .A(A[748]), .B(B[0]), .Z(\ab[748][0] ) );
  AND U1132 ( .A(B[3]), .B(A[747]), .Z(\ab[747][3] ) );
  AND U1133 ( .A(B[2]), .B(A[747]), .Z(\ab[747][2] ) );
  AND U1134 ( .A(B[1]), .B(A[747]), .Z(\ab[747][1] ) );
  AND U1135 ( .A(A[747]), .B(B[0]), .Z(\ab[747][0] ) );
  AND U1136 ( .A(B[3]), .B(A[746]), .Z(\ab[746][3] ) );
  AND U1137 ( .A(B[2]), .B(A[746]), .Z(\ab[746][2] ) );
  AND U1138 ( .A(B[1]), .B(A[746]), .Z(\ab[746][1] ) );
  AND U1139 ( .A(A[746]), .B(B[0]), .Z(\ab[746][0] ) );
  AND U1140 ( .A(B[3]), .B(A[745]), .Z(\ab[745][3] ) );
  AND U1141 ( .A(B[2]), .B(A[745]), .Z(\ab[745][2] ) );
  AND U1142 ( .A(B[1]), .B(A[745]), .Z(\ab[745][1] ) );
  AND U1143 ( .A(A[745]), .B(B[0]), .Z(\ab[745][0] ) );
  AND U1144 ( .A(B[3]), .B(A[744]), .Z(\ab[744][3] ) );
  AND U1145 ( .A(B[2]), .B(A[744]), .Z(\ab[744][2] ) );
  AND U1146 ( .A(B[1]), .B(A[744]), .Z(\ab[744][1] ) );
  AND U1147 ( .A(A[744]), .B(B[0]), .Z(\ab[744][0] ) );
  AND U1148 ( .A(B[3]), .B(A[743]), .Z(\ab[743][3] ) );
  AND U1149 ( .A(B[2]), .B(A[743]), .Z(\ab[743][2] ) );
  AND U1150 ( .A(B[1]), .B(A[743]), .Z(\ab[743][1] ) );
  AND U1151 ( .A(A[743]), .B(B[0]), .Z(\ab[743][0] ) );
  AND U1152 ( .A(B[3]), .B(A[742]), .Z(\ab[742][3] ) );
  AND U1153 ( .A(B[2]), .B(A[742]), .Z(\ab[742][2] ) );
  AND U1154 ( .A(B[1]), .B(A[742]), .Z(\ab[742][1] ) );
  AND U1155 ( .A(A[742]), .B(B[0]), .Z(\ab[742][0] ) );
  AND U1156 ( .A(B[3]), .B(A[741]), .Z(\ab[741][3] ) );
  AND U1157 ( .A(B[2]), .B(A[741]), .Z(\ab[741][2] ) );
  AND U1158 ( .A(B[1]), .B(A[741]), .Z(\ab[741][1] ) );
  AND U1159 ( .A(A[741]), .B(B[0]), .Z(\ab[741][0] ) );
  AND U1160 ( .A(B[3]), .B(A[740]), .Z(\ab[740][3] ) );
  AND U1161 ( .A(B[2]), .B(A[740]), .Z(\ab[740][2] ) );
  AND U1162 ( .A(B[1]), .B(A[740]), .Z(\ab[740][1] ) );
  AND U1163 ( .A(A[740]), .B(B[0]), .Z(\ab[740][0] ) );
  AND U1164 ( .A(B[3]), .B(A[73]), .Z(\ab[73][3] ) );
  AND U1165 ( .A(B[2]), .B(A[73]), .Z(\ab[73][2] ) );
  AND U1166 ( .A(B[1]), .B(A[73]), .Z(\ab[73][1] ) );
  AND U1167 ( .A(A[73]), .B(B[0]), .Z(\ab[73][0] ) );
  AND U1168 ( .A(B[3]), .B(A[739]), .Z(\ab[739][3] ) );
  AND U1169 ( .A(B[2]), .B(A[739]), .Z(\ab[739][2] ) );
  AND U1170 ( .A(B[1]), .B(A[739]), .Z(\ab[739][1] ) );
  AND U1171 ( .A(A[739]), .B(B[0]), .Z(\ab[739][0] ) );
  AND U1172 ( .A(B[3]), .B(A[738]), .Z(\ab[738][3] ) );
  AND U1173 ( .A(B[2]), .B(A[738]), .Z(\ab[738][2] ) );
  AND U1174 ( .A(B[1]), .B(A[738]), .Z(\ab[738][1] ) );
  AND U1175 ( .A(A[738]), .B(B[0]), .Z(\ab[738][0] ) );
  AND U1176 ( .A(B[3]), .B(A[737]), .Z(\ab[737][3] ) );
  AND U1177 ( .A(B[2]), .B(A[737]), .Z(\ab[737][2] ) );
  AND U1178 ( .A(B[1]), .B(A[737]), .Z(\ab[737][1] ) );
  AND U1179 ( .A(A[737]), .B(B[0]), .Z(\ab[737][0] ) );
  AND U1180 ( .A(B[3]), .B(A[736]), .Z(\ab[736][3] ) );
  AND U1181 ( .A(B[2]), .B(A[736]), .Z(\ab[736][2] ) );
  AND U1182 ( .A(B[1]), .B(A[736]), .Z(\ab[736][1] ) );
  AND U1183 ( .A(A[736]), .B(B[0]), .Z(\ab[736][0] ) );
  AND U1184 ( .A(B[3]), .B(A[735]), .Z(\ab[735][3] ) );
  AND U1185 ( .A(B[2]), .B(A[735]), .Z(\ab[735][2] ) );
  AND U1186 ( .A(B[1]), .B(A[735]), .Z(\ab[735][1] ) );
  AND U1187 ( .A(A[735]), .B(B[0]), .Z(\ab[735][0] ) );
  AND U1188 ( .A(B[3]), .B(A[734]), .Z(\ab[734][3] ) );
  AND U1189 ( .A(B[2]), .B(A[734]), .Z(\ab[734][2] ) );
  AND U1190 ( .A(B[1]), .B(A[734]), .Z(\ab[734][1] ) );
  AND U1191 ( .A(A[734]), .B(B[0]), .Z(\ab[734][0] ) );
  AND U1192 ( .A(B[3]), .B(A[733]), .Z(\ab[733][3] ) );
  AND U1193 ( .A(B[2]), .B(A[733]), .Z(\ab[733][2] ) );
  AND U1194 ( .A(B[1]), .B(A[733]), .Z(\ab[733][1] ) );
  AND U1195 ( .A(A[733]), .B(B[0]), .Z(\ab[733][0] ) );
  AND U1196 ( .A(B[3]), .B(A[732]), .Z(\ab[732][3] ) );
  AND U1197 ( .A(B[2]), .B(A[732]), .Z(\ab[732][2] ) );
  AND U1198 ( .A(B[1]), .B(A[732]), .Z(\ab[732][1] ) );
  AND U1199 ( .A(A[732]), .B(B[0]), .Z(\ab[732][0] ) );
  AND U1200 ( .A(B[3]), .B(A[731]), .Z(\ab[731][3] ) );
  AND U1201 ( .A(B[2]), .B(A[731]), .Z(\ab[731][2] ) );
  AND U1202 ( .A(B[1]), .B(A[731]), .Z(\ab[731][1] ) );
  AND U1203 ( .A(A[731]), .B(B[0]), .Z(\ab[731][0] ) );
  AND U1204 ( .A(B[3]), .B(A[730]), .Z(\ab[730][3] ) );
  AND U1205 ( .A(B[2]), .B(A[730]), .Z(\ab[730][2] ) );
  AND U1206 ( .A(B[1]), .B(A[730]), .Z(\ab[730][1] ) );
  AND U1207 ( .A(A[730]), .B(B[0]), .Z(\ab[730][0] ) );
  AND U1208 ( .A(B[3]), .B(A[72]), .Z(\ab[72][3] ) );
  AND U1209 ( .A(B[2]), .B(A[72]), .Z(\ab[72][2] ) );
  AND U1210 ( .A(B[1]), .B(A[72]), .Z(\ab[72][1] ) );
  AND U1211 ( .A(A[72]), .B(B[0]), .Z(\ab[72][0] ) );
  AND U1212 ( .A(B[3]), .B(A[729]), .Z(\ab[729][3] ) );
  AND U1213 ( .A(B[2]), .B(A[729]), .Z(\ab[729][2] ) );
  AND U1214 ( .A(B[1]), .B(A[729]), .Z(\ab[729][1] ) );
  AND U1215 ( .A(A[729]), .B(B[0]), .Z(\ab[729][0] ) );
  AND U1216 ( .A(B[3]), .B(A[728]), .Z(\ab[728][3] ) );
  AND U1217 ( .A(B[2]), .B(A[728]), .Z(\ab[728][2] ) );
  AND U1218 ( .A(B[1]), .B(A[728]), .Z(\ab[728][1] ) );
  AND U1219 ( .A(A[728]), .B(B[0]), .Z(\ab[728][0] ) );
  AND U1220 ( .A(B[3]), .B(A[727]), .Z(\ab[727][3] ) );
  AND U1221 ( .A(B[2]), .B(A[727]), .Z(\ab[727][2] ) );
  AND U1222 ( .A(B[1]), .B(A[727]), .Z(\ab[727][1] ) );
  AND U1223 ( .A(A[727]), .B(B[0]), .Z(\ab[727][0] ) );
  AND U1224 ( .A(B[3]), .B(A[726]), .Z(\ab[726][3] ) );
  AND U1225 ( .A(B[2]), .B(A[726]), .Z(\ab[726][2] ) );
  AND U1226 ( .A(B[1]), .B(A[726]), .Z(\ab[726][1] ) );
  AND U1227 ( .A(A[726]), .B(B[0]), .Z(\ab[726][0] ) );
  AND U1228 ( .A(B[3]), .B(A[725]), .Z(\ab[725][3] ) );
  AND U1229 ( .A(B[2]), .B(A[725]), .Z(\ab[725][2] ) );
  AND U1230 ( .A(B[1]), .B(A[725]), .Z(\ab[725][1] ) );
  AND U1231 ( .A(A[725]), .B(B[0]), .Z(\ab[725][0] ) );
  AND U1232 ( .A(B[3]), .B(A[724]), .Z(\ab[724][3] ) );
  AND U1233 ( .A(B[2]), .B(A[724]), .Z(\ab[724][2] ) );
  AND U1234 ( .A(B[1]), .B(A[724]), .Z(\ab[724][1] ) );
  AND U1235 ( .A(A[724]), .B(B[0]), .Z(\ab[724][0] ) );
  AND U1236 ( .A(B[3]), .B(A[723]), .Z(\ab[723][3] ) );
  AND U1237 ( .A(B[2]), .B(A[723]), .Z(\ab[723][2] ) );
  AND U1238 ( .A(B[1]), .B(A[723]), .Z(\ab[723][1] ) );
  AND U1239 ( .A(A[723]), .B(B[0]), .Z(\ab[723][0] ) );
  AND U1240 ( .A(B[3]), .B(A[722]), .Z(\ab[722][3] ) );
  AND U1241 ( .A(B[2]), .B(A[722]), .Z(\ab[722][2] ) );
  AND U1242 ( .A(B[1]), .B(A[722]), .Z(\ab[722][1] ) );
  AND U1243 ( .A(A[722]), .B(B[0]), .Z(\ab[722][0] ) );
  AND U1244 ( .A(B[3]), .B(A[721]), .Z(\ab[721][3] ) );
  AND U1245 ( .A(B[2]), .B(A[721]), .Z(\ab[721][2] ) );
  AND U1246 ( .A(B[1]), .B(A[721]), .Z(\ab[721][1] ) );
  AND U1247 ( .A(A[721]), .B(B[0]), .Z(\ab[721][0] ) );
  AND U1248 ( .A(B[3]), .B(A[720]), .Z(\ab[720][3] ) );
  AND U1249 ( .A(B[2]), .B(A[720]), .Z(\ab[720][2] ) );
  AND U1250 ( .A(B[1]), .B(A[720]), .Z(\ab[720][1] ) );
  AND U1251 ( .A(A[720]), .B(B[0]), .Z(\ab[720][0] ) );
  AND U1252 ( .A(B[3]), .B(A[71]), .Z(\ab[71][3] ) );
  AND U1253 ( .A(B[2]), .B(A[71]), .Z(\ab[71][2] ) );
  AND U1254 ( .A(B[1]), .B(A[71]), .Z(\ab[71][1] ) );
  AND U1255 ( .A(A[71]), .B(B[0]), .Z(\ab[71][0] ) );
  AND U1256 ( .A(B[3]), .B(A[719]), .Z(\ab[719][3] ) );
  AND U1257 ( .A(B[2]), .B(A[719]), .Z(\ab[719][2] ) );
  AND U1258 ( .A(B[1]), .B(A[719]), .Z(\ab[719][1] ) );
  AND U1259 ( .A(A[719]), .B(B[0]), .Z(\ab[719][0] ) );
  AND U1260 ( .A(B[3]), .B(A[718]), .Z(\ab[718][3] ) );
  AND U1261 ( .A(B[2]), .B(A[718]), .Z(\ab[718][2] ) );
  AND U1262 ( .A(B[1]), .B(A[718]), .Z(\ab[718][1] ) );
  AND U1263 ( .A(A[718]), .B(B[0]), .Z(\ab[718][0] ) );
  AND U1264 ( .A(B[3]), .B(A[717]), .Z(\ab[717][3] ) );
  AND U1265 ( .A(B[2]), .B(A[717]), .Z(\ab[717][2] ) );
  AND U1266 ( .A(B[1]), .B(A[717]), .Z(\ab[717][1] ) );
  AND U1267 ( .A(A[717]), .B(B[0]), .Z(\ab[717][0] ) );
  AND U1268 ( .A(B[3]), .B(A[716]), .Z(\ab[716][3] ) );
  AND U1269 ( .A(B[2]), .B(A[716]), .Z(\ab[716][2] ) );
  AND U1270 ( .A(B[1]), .B(A[716]), .Z(\ab[716][1] ) );
  AND U1271 ( .A(A[716]), .B(B[0]), .Z(\ab[716][0] ) );
  AND U1272 ( .A(B[3]), .B(A[715]), .Z(\ab[715][3] ) );
  AND U1273 ( .A(B[2]), .B(A[715]), .Z(\ab[715][2] ) );
  AND U1274 ( .A(B[1]), .B(A[715]), .Z(\ab[715][1] ) );
  AND U1275 ( .A(A[715]), .B(B[0]), .Z(\ab[715][0] ) );
  AND U1276 ( .A(B[3]), .B(A[714]), .Z(\ab[714][3] ) );
  AND U1277 ( .A(B[2]), .B(A[714]), .Z(\ab[714][2] ) );
  AND U1278 ( .A(B[1]), .B(A[714]), .Z(\ab[714][1] ) );
  AND U1279 ( .A(A[714]), .B(B[0]), .Z(\ab[714][0] ) );
  AND U1280 ( .A(B[3]), .B(A[713]), .Z(\ab[713][3] ) );
  AND U1281 ( .A(B[2]), .B(A[713]), .Z(\ab[713][2] ) );
  AND U1282 ( .A(B[1]), .B(A[713]), .Z(\ab[713][1] ) );
  AND U1283 ( .A(A[713]), .B(B[0]), .Z(\ab[713][0] ) );
  AND U1284 ( .A(B[3]), .B(A[712]), .Z(\ab[712][3] ) );
  AND U1285 ( .A(B[2]), .B(A[712]), .Z(\ab[712][2] ) );
  AND U1286 ( .A(B[1]), .B(A[712]), .Z(\ab[712][1] ) );
  AND U1287 ( .A(A[712]), .B(B[0]), .Z(\ab[712][0] ) );
  AND U1288 ( .A(B[3]), .B(A[711]), .Z(\ab[711][3] ) );
  AND U1289 ( .A(B[2]), .B(A[711]), .Z(\ab[711][2] ) );
  AND U1290 ( .A(B[1]), .B(A[711]), .Z(\ab[711][1] ) );
  AND U1291 ( .A(A[711]), .B(B[0]), .Z(\ab[711][0] ) );
  AND U1292 ( .A(B[3]), .B(A[710]), .Z(\ab[710][3] ) );
  AND U1293 ( .A(B[2]), .B(A[710]), .Z(\ab[710][2] ) );
  AND U1294 ( .A(B[1]), .B(A[710]), .Z(\ab[710][1] ) );
  AND U1295 ( .A(A[710]), .B(B[0]), .Z(\ab[710][0] ) );
  AND U1296 ( .A(B[3]), .B(A[70]), .Z(\ab[70][3] ) );
  AND U1297 ( .A(B[2]), .B(A[70]), .Z(\ab[70][2] ) );
  AND U1298 ( .A(B[1]), .B(A[70]), .Z(\ab[70][1] ) );
  AND U1299 ( .A(A[70]), .B(B[0]), .Z(\ab[70][0] ) );
  AND U1300 ( .A(B[3]), .B(A[709]), .Z(\ab[709][3] ) );
  AND U1301 ( .A(B[2]), .B(A[709]), .Z(\ab[709][2] ) );
  AND U1302 ( .A(B[1]), .B(A[709]), .Z(\ab[709][1] ) );
  AND U1303 ( .A(A[709]), .B(B[0]), .Z(\ab[709][0] ) );
  AND U1304 ( .A(B[3]), .B(A[708]), .Z(\ab[708][3] ) );
  AND U1305 ( .A(B[2]), .B(A[708]), .Z(\ab[708][2] ) );
  AND U1306 ( .A(B[1]), .B(A[708]), .Z(\ab[708][1] ) );
  AND U1307 ( .A(A[708]), .B(B[0]), .Z(\ab[708][0] ) );
  AND U1308 ( .A(B[3]), .B(A[707]), .Z(\ab[707][3] ) );
  AND U1309 ( .A(B[2]), .B(A[707]), .Z(\ab[707][2] ) );
  AND U1310 ( .A(B[1]), .B(A[707]), .Z(\ab[707][1] ) );
  AND U1311 ( .A(A[707]), .B(B[0]), .Z(\ab[707][0] ) );
  AND U1312 ( .A(B[3]), .B(A[706]), .Z(\ab[706][3] ) );
  AND U1313 ( .A(B[2]), .B(A[706]), .Z(\ab[706][2] ) );
  AND U1314 ( .A(B[1]), .B(A[706]), .Z(\ab[706][1] ) );
  AND U1315 ( .A(A[706]), .B(B[0]), .Z(\ab[706][0] ) );
  AND U1316 ( .A(B[3]), .B(A[705]), .Z(\ab[705][3] ) );
  AND U1317 ( .A(B[2]), .B(A[705]), .Z(\ab[705][2] ) );
  AND U1318 ( .A(B[1]), .B(A[705]), .Z(\ab[705][1] ) );
  AND U1319 ( .A(A[705]), .B(B[0]), .Z(\ab[705][0] ) );
  AND U1320 ( .A(B[3]), .B(A[704]), .Z(\ab[704][3] ) );
  AND U1321 ( .A(B[2]), .B(A[704]), .Z(\ab[704][2] ) );
  AND U1322 ( .A(B[1]), .B(A[704]), .Z(\ab[704][1] ) );
  AND U1323 ( .A(A[704]), .B(B[0]), .Z(\ab[704][0] ) );
  AND U1324 ( .A(B[3]), .B(A[703]), .Z(\ab[703][3] ) );
  AND U1325 ( .A(B[2]), .B(A[703]), .Z(\ab[703][2] ) );
  AND U1326 ( .A(B[1]), .B(A[703]), .Z(\ab[703][1] ) );
  AND U1327 ( .A(A[703]), .B(B[0]), .Z(\ab[703][0] ) );
  AND U1328 ( .A(B[3]), .B(A[702]), .Z(\ab[702][3] ) );
  AND U1329 ( .A(B[2]), .B(A[702]), .Z(\ab[702][2] ) );
  AND U1330 ( .A(B[1]), .B(A[702]), .Z(\ab[702][1] ) );
  AND U1331 ( .A(A[702]), .B(B[0]), .Z(\ab[702][0] ) );
  AND U1332 ( .A(B[3]), .B(A[701]), .Z(\ab[701][3] ) );
  AND U1333 ( .A(B[2]), .B(A[701]), .Z(\ab[701][2] ) );
  AND U1334 ( .A(B[1]), .B(A[701]), .Z(\ab[701][1] ) );
  AND U1335 ( .A(A[701]), .B(B[0]), .Z(\ab[701][0] ) );
  AND U1336 ( .A(B[3]), .B(A[700]), .Z(\ab[700][3] ) );
  AND U1337 ( .A(B[2]), .B(A[700]), .Z(\ab[700][2] ) );
  AND U1338 ( .A(B[1]), .B(A[700]), .Z(\ab[700][1] ) );
  AND U1339 ( .A(A[700]), .B(B[0]), .Z(\ab[700][0] ) );
  AND U1340 ( .A(B[3]), .B(A[6]), .Z(\ab[6][3] ) );
  AND U1341 ( .A(B[2]), .B(A[6]), .Z(\ab[6][2] ) );
  AND U1342 ( .A(B[1]), .B(A[6]), .Z(\ab[6][1] ) );
  AND U1343 ( .A(A[6]), .B(B[0]), .Z(\ab[6][0] ) );
  AND U1344 ( .A(B[3]), .B(A[69]), .Z(\ab[69][3] ) );
  AND U1345 ( .A(B[2]), .B(A[69]), .Z(\ab[69][2] ) );
  AND U1346 ( .A(B[1]), .B(A[69]), .Z(\ab[69][1] ) );
  AND U1347 ( .A(A[69]), .B(B[0]), .Z(\ab[69][0] ) );
  AND U1348 ( .A(B[3]), .B(A[699]), .Z(\ab[699][3] ) );
  AND U1349 ( .A(B[2]), .B(A[699]), .Z(\ab[699][2] ) );
  AND U1350 ( .A(B[1]), .B(A[699]), .Z(\ab[699][1] ) );
  AND U1351 ( .A(A[699]), .B(B[0]), .Z(\ab[699][0] ) );
  AND U1352 ( .A(B[3]), .B(A[698]), .Z(\ab[698][3] ) );
  AND U1353 ( .A(B[2]), .B(A[698]), .Z(\ab[698][2] ) );
  AND U1354 ( .A(B[1]), .B(A[698]), .Z(\ab[698][1] ) );
  AND U1355 ( .A(A[698]), .B(B[0]), .Z(\ab[698][0] ) );
  AND U1356 ( .A(B[3]), .B(A[697]), .Z(\ab[697][3] ) );
  AND U1357 ( .A(B[2]), .B(A[697]), .Z(\ab[697][2] ) );
  AND U1358 ( .A(B[1]), .B(A[697]), .Z(\ab[697][1] ) );
  AND U1359 ( .A(A[697]), .B(B[0]), .Z(\ab[697][0] ) );
  AND U1360 ( .A(B[3]), .B(A[696]), .Z(\ab[696][3] ) );
  AND U1361 ( .A(B[2]), .B(A[696]), .Z(\ab[696][2] ) );
  AND U1362 ( .A(B[1]), .B(A[696]), .Z(\ab[696][1] ) );
  AND U1363 ( .A(A[696]), .B(B[0]), .Z(\ab[696][0] ) );
  AND U1364 ( .A(B[3]), .B(A[695]), .Z(\ab[695][3] ) );
  AND U1365 ( .A(B[2]), .B(A[695]), .Z(\ab[695][2] ) );
  AND U1366 ( .A(B[1]), .B(A[695]), .Z(\ab[695][1] ) );
  AND U1367 ( .A(A[695]), .B(B[0]), .Z(\ab[695][0] ) );
  AND U1368 ( .A(B[3]), .B(A[694]), .Z(\ab[694][3] ) );
  AND U1369 ( .A(B[2]), .B(A[694]), .Z(\ab[694][2] ) );
  AND U1370 ( .A(B[1]), .B(A[694]), .Z(\ab[694][1] ) );
  AND U1371 ( .A(A[694]), .B(B[0]), .Z(\ab[694][0] ) );
  AND U1372 ( .A(B[3]), .B(A[693]), .Z(\ab[693][3] ) );
  AND U1373 ( .A(B[2]), .B(A[693]), .Z(\ab[693][2] ) );
  AND U1374 ( .A(B[1]), .B(A[693]), .Z(\ab[693][1] ) );
  AND U1375 ( .A(A[693]), .B(B[0]), .Z(\ab[693][0] ) );
  AND U1376 ( .A(B[3]), .B(A[692]), .Z(\ab[692][3] ) );
  AND U1377 ( .A(B[2]), .B(A[692]), .Z(\ab[692][2] ) );
  AND U1378 ( .A(B[1]), .B(A[692]), .Z(\ab[692][1] ) );
  AND U1379 ( .A(A[692]), .B(B[0]), .Z(\ab[692][0] ) );
  AND U1380 ( .A(B[3]), .B(A[691]), .Z(\ab[691][3] ) );
  AND U1381 ( .A(B[2]), .B(A[691]), .Z(\ab[691][2] ) );
  AND U1382 ( .A(B[1]), .B(A[691]), .Z(\ab[691][1] ) );
  AND U1383 ( .A(A[691]), .B(B[0]), .Z(\ab[691][0] ) );
  AND U1384 ( .A(B[3]), .B(A[690]), .Z(\ab[690][3] ) );
  AND U1385 ( .A(B[2]), .B(A[690]), .Z(\ab[690][2] ) );
  AND U1386 ( .A(B[1]), .B(A[690]), .Z(\ab[690][1] ) );
  AND U1387 ( .A(A[690]), .B(B[0]), .Z(\ab[690][0] ) );
  AND U1388 ( .A(B[3]), .B(A[68]), .Z(\ab[68][3] ) );
  AND U1389 ( .A(B[2]), .B(A[68]), .Z(\ab[68][2] ) );
  AND U1390 ( .A(B[1]), .B(A[68]), .Z(\ab[68][1] ) );
  AND U1391 ( .A(A[68]), .B(B[0]), .Z(\ab[68][0] ) );
  AND U1392 ( .A(B[3]), .B(A[689]), .Z(\ab[689][3] ) );
  AND U1393 ( .A(B[2]), .B(A[689]), .Z(\ab[689][2] ) );
  AND U1394 ( .A(B[1]), .B(A[689]), .Z(\ab[689][1] ) );
  AND U1395 ( .A(A[689]), .B(B[0]), .Z(\ab[689][0] ) );
  AND U1396 ( .A(B[3]), .B(A[688]), .Z(\ab[688][3] ) );
  AND U1397 ( .A(B[2]), .B(A[688]), .Z(\ab[688][2] ) );
  AND U1398 ( .A(B[1]), .B(A[688]), .Z(\ab[688][1] ) );
  AND U1399 ( .A(A[688]), .B(B[0]), .Z(\ab[688][0] ) );
  AND U1400 ( .A(B[3]), .B(A[687]), .Z(\ab[687][3] ) );
  AND U1401 ( .A(B[2]), .B(A[687]), .Z(\ab[687][2] ) );
  AND U1402 ( .A(B[1]), .B(A[687]), .Z(\ab[687][1] ) );
  AND U1403 ( .A(A[687]), .B(B[0]), .Z(\ab[687][0] ) );
  AND U1404 ( .A(B[3]), .B(A[686]), .Z(\ab[686][3] ) );
  AND U1405 ( .A(B[2]), .B(A[686]), .Z(\ab[686][2] ) );
  AND U1406 ( .A(B[1]), .B(A[686]), .Z(\ab[686][1] ) );
  AND U1407 ( .A(A[686]), .B(B[0]), .Z(\ab[686][0] ) );
  AND U1408 ( .A(B[3]), .B(A[685]), .Z(\ab[685][3] ) );
  AND U1409 ( .A(B[2]), .B(A[685]), .Z(\ab[685][2] ) );
  AND U1410 ( .A(B[1]), .B(A[685]), .Z(\ab[685][1] ) );
  AND U1411 ( .A(A[685]), .B(B[0]), .Z(\ab[685][0] ) );
  AND U1412 ( .A(B[3]), .B(A[684]), .Z(\ab[684][3] ) );
  AND U1413 ( .A(B[2]), .B(A[684]), .Z(\ab[684][2] ) );
  AND U1414 ( .A(B[1]), .B(A[684]), .Z(\ab[684][1] ) );
  AND U1415 ( .A(A[684]), .B(B[0]), .Z(\ab[684][0] ) );
  AND U1416 ( .A(B[3]), .B(A[683]), .Z(\ab[683][3] ) );
  AND U1417 ( .A(B[2]), .B(A[683]), .Z(\ab[683][2] ) );
  AND U1418 ( .A(B[1]), .B(A[683]), .Z(\ab[683][1] ) );
  AND U1419 ( .A(A[683]), .B(B[0]), .Z(\ab[683][0] ) );
  AND U1420 ( .A(B[3]), .B(A[682]), .Z(\ab[682][3] ) );
  AND U1421 ( .A(B[2]), .B(A[682]), .Z(\ab[682][2] ) );
  AND U1422 ( .A(B[1]), .B(A[682]), .Z(\ab[682][1] ) );
  AND U1423 ( .A(A[682]), .B(B[0]), .Z(\ab[682][0] ) );
  AND U1424 ( .A(B[3]), .B(A[681]), .Z(\ab[681][3] ) );
  AND U1425 ( .A(B[2]), .B(A[681]), .Z(\ab[681][2] ) );
  AND U1426 ( .A(B[1]), .B(A[681]), .Z(\ab[681][1] ) );
  AND U1427 ( .A(A[681]), .B(B[0]), .Z(\ab[681][0] ) );
  AND U1428 ( .A(B[3]), .B(A[680]), .Z(\ab[680][3] ) );
  AND U1429 ( .A(B[2]), .B(A[680]), .Z(\ab[680][2] ) );
  AND U1430 ( .A(B[1]), .B(A[680]), .Z(\ab[680][1] ) );
  AND U1431 ( .A(A[680]), .B(B[0]), .Z(\ab[680][0] ) );
  AND U1432 ( .A(B[3]), .B(A[67]), .Z(\ab[67][3] ) );
  AND U1433 ( .A(B[2]), .B(A[67]), .Z(\ab[67][2] ) );
  AND U1434 ( .A(B[1]), .B(A[67]), .Z(\ab[67][1] ) );
  AND U1435 ( .A(A[67]), .B(B[0]), .Z(\ab[67][0] ) );
  AND U1436 ( .A(B[3]), .B(A[679]), .Z(\ab[679][3] ) );
  AND U1437 ( .A(B[2]), .B(A[679]), .Z(\ab[679][2] ) );
  AND U1438 ( .A(B[1]), .B(A[679]), .Z(\ab[679][1] ) );
  AND U1439 ( .A(A[679]), .B(B[0]), .Z(\ab[679][0] ) );
  AND U1440 ( .A(B[3]), .B(A[678]), .Z(\ab[678][3] ) );
  AND U1441 ( .A(B[2]), .B(A[678]), .Z(\ab[678][2] ) );
  AND U1442 ( .A(B[1]), .B(A[678]), .Z(\ab[678][1] ) );
  AND U1443 ( .A(A[678]), .B(B[0]), .Z(\ab[678][0] ) );
  AND U1444 ( .A(B[3]), .B(A[677]), .Z(\ab[677][3] ) );
  AND U1445 ( .A(B[2]), .B(A[677]), .Z(\ab[677][2] ) );
  AND U1446 ( .A(B[1]), .B(A[677]), .Z(\ab[677][1] ) );
  AND U1447 ( .A(A[677]), .B(B[0]), .Z(\ab[677][0] ) );
  AND U1448 ( .A(B[3]), .B(A[676]), .Z(\ab[676][3] ) );
  AND U1449 ( .A(B[2]), .B(A[676]), .Z(\ab[676][2] ) );
  AND U1450 ( .A(B[1]), .B(A[676]), .Z(\ab[676][1] ) );
  AND U1451 ( .A(A[676]), .B(B[0]), .Z(\ab[676][0] ) );
  AND U1452 ( .A(B[3]), .B(A[675]), .Z(\ab[675][3] ) );
  AND U1453 ( .A(B[2]), .B(A[675]), .Z(\ab[675][2] ) );
  AND U1454 ( .A(B[1]), .B(A[675]), .Z(\ab[675][1] ) );
  AND U1455 ( .A(A[675]), .B(B[0]), .Z(\ab[675][0] ) );
  AND U1456 ( .A(B[3]), .B(A[674]), .Z(\ab[674][3] ) );
  AND U1457 ( .A(B[2]), .B(A[674]), .Z(\ab[674][2] ) );
  AND U1458 ( .A(B[1]), .B(A[674]), .Z(\ab[674][1] ) );
  AND U1459 ( .A(A[674]), .B(B[0]), .Z(\ab[674][0] ) );
  AND U1460 ( .A(B[3]), .B(A[673]), .Z(\ab[673][3] ) );
  AND U1461 ( .A(B[2]), .B(A[673]), .Z(\ab[673][2] ) );
  AND U1462 ( .A(B[1]), .B(A[673]), .Z(\ab[673][1] ) );
  AND U1463 ( .A(A[673]), .B(B[0]), .Z(\ab[673][0] ) );
  AND U1464 ( .A(B[3]), .B(A[672]), .Z(\ab[672][3] ) );
  AND U1465 ( .A(B[2]), .B(A[672]), .Z(\ab[672][2] ) );
  AND U1466 ( .A(B[1]), .B(A[672]), .Z(\ab[672][1] ) );
  AND U1467 ( .A(A[672]), .B(B[0]), .Z(\ab[672][0] ) );
  AND U1468 ( .A(B[3]), .B(A[671]), .Z(\ab[671][3] ) );
  AND U1469 ( .A(B[2]), .B(A[671]), .Z(\ab[671][2] ) );
  AND U1470 ( .A(B[1]), .B(A[671]), .Z(\ab[671][1] ) );
  AND U1471 ( .A(A[671]), .B(B[0]), .Z(\ab[671][0] ) );
  AND U1472 ( .A(B[3]), .B(A[670]), .Z(\ab[670][3] ) );
  AND U1473 ( .A(B[2]), .B(A[670]), .Z(\ab[670][2] ) );
  AND U1474 ( .A(B[1]), .B(A[670]), .Z(\ab[670][1] ) );
  AND U1475 ( .A(A[670]), .B(B[0]), .Z(\ab[670][0] ) );
  AND U1476 ( .A(B[3]), .B(A[66]), .Z(\ab[66][3] ) );
  AND U1477 ( .A(B[2]), .B(A[66]), .Z(\ab[66][2] ) );
  AND U1478 ( .A(B[1]), .B(A[66]), .Z(\ab[66][1] ) );
  AND U1479 ( .A(A[66]), .B(B[0]), .Z(\ab[66][0] ) );
  AND U1480 ( .A(B[3]), .B(A[669]), .Z(\ab[669][3] ) );
  AND U1481 ( .A(B[2]), .B(A[669]), .Z(\ab[669][2] ) );
  AND U1482 ( .A(B[1]), .B(A[669]), .Z(\ab[669][1] ) );
  AND U1483 ( .A(A[669]), .B(B[0]), .Z(\ab[669][0] ) );
  AND U1484 ( .A(B[3]), .B(A[668]), .Z(\ab[668][3] ) );
  AND U1485 ( .A(B[2]), .B(A[668]), .Z(\ab[668][2] ) );
  AND U1486 ( .A(B[1]), .B(A[668]), .Z(\ab[668][1] ) );
  AND U1487 ( .A(A[668]), .B(B[0]), .Z(\ab[668][0] ) );
  AND U1488 ( .A(B[3]), .B(A[667]), .Z(\ab[667][3] ) );
  AND U1489 ( .A(B[2]), .B(A[667]), .Z(\ab[667][2] ) );
  AND U1490 ( .A(B[1]), .B(A[667]), .Z(\ab[667][1] ) );
  AND U1491 ( .A(A[667]), .B(B[0]), .Z(\ab[667][0] ) );
  AND U1492 ( .A(B[3]), .B(A[666]), .Z(\ab[666][3] ) );
  AND U1493 ( .A(B[2]), .B(A[666]), .Z(\ab[666][2] ) );
  AND U1494 ( .A(B[1]), .B(A[666]), .Z(\ab[666][1] ) );
  AND U1495 ( .A(A[666]), .B(B[0]), .Z(\ab[666][0] ) );
  AND U1496 ( .A(B[3]), .B(A[665]), .Z(\ab[665][3] ) );
  AND U1497 ( .A(B[2]), .B(A[665]), .Z(\ab[665][2] ) );
  AND U1498 ( .A(B[1]), .B(A[665]), .Z(\ab[665][1] ) );
  AND U1499 ( .A(A[665]), .B(B[0]), .Z(\ab[665][0] ) );
  AND U1500 ( .A(B[3]), .B(A[664]), .Z(\ab[664][3] ) );
  AND U1501 ( .A(B[2]), .B(A[664]), .Z(\ab[664][2] ) );
  AND U1502 ( .A(B[1]), .B(A[664]), .Z(\ab[664][1] ) );
  AND U1503 ( .A(A[664]), .B(B[0]), .Z(\ab[664][0] ) );
  AND U1504 ( .A(B[3]), .B(A[663]), .Z(\ab[663][3] ) );
  AND U1505 ( .A(B[2]), .B(A[663]), .Z(\ab[663][2] ) );
  AND U1506 ( .A(B[1]), .B(A[663]), .Z(\ab[663][1] ) );
  AND U1507 ( .A(A[663]), .B(B[0]), .Z(\ab[663][0] ) );
  AND U1508 ( .A(B[3]), .B(A[662]), .Z(\ab[662][3] ) );
  AND U1509 ( .A(B[2]), .B(A[662]), .Z(\ab[662][2] ) );
  AND U1510 ( .A(B[1]), .B(A[662]), .Z(\ab[662][1] ) );
  AND U1511 ( .A(A[662]), .B(B[0]), .Z(\ab[662][0] ) );
  AND U1512 ( .A(B[3]), .B(A[661]), .Z(\ab[661][3] ) );
  AND U1513 ( .A(B[2]), .B(A[661]), .Z(\ab[661][2] ) );
  AND U1514 ( .A(B[1]), .B(A[661]), .Z(\ab[661][1] ) );
  AND U1515 ( .A(A[661]), .B(B[0]), .Z(\ab[661][0] ) );
  AND U1516 ( .A(B[3]), .B(A[660]), .Z(\ab[660][3] ) );
  AND U1517 ( .A(B[2]), .B(A[660]), .Z(\ab[660][2] ) );
  AND U1518 ( .A(B[1]), .B(A[660]), .Z(\ab[660][1] ) );
  AND U1519 ( .A(A[660]), .B(B[0]), .Z(\ab[660][0] ) );
  AND U1520 ( .A(B[3]), .B(A[65]), .Z(\ab[65][3] ) );
  AND U1521 ( .A(B[2]), .B(A[65]), .Z(\ab[65][2] ) );
  AND U1522 ( .A(B[1]), .B(A[65]), .Z(\ab[65][1] ) );
  AND U1523 ( .A(A[65]), .B(B[0]), .Z(\ab[65][0] ) );
  AND U1524 ( .A(B[3]), .B(A[659]), .Z(\ab[659][3] ) );
  AND U1525 ( .A(B[2]), .B(A[659]), .Z(\ab[659][2] ) );
  AND U1526 ( .A(B[1]), .B(A[659]), .Z(\ab[659][1] ) );
  AND U1527 ( .A(A[659]), .B(B[0]), .Z(\ab[659][0] ) );
  AND U1528 ( .A(B[3]), .B(A[658]), .Z(\ab[658][3] ) );
  AND U1529 ( .A(B[2]), .B(A[658]), .Z(\ab[658][2] ) );
  AND U1530 ( .A(B[1]), .B(A[658]), .Z(\ab[658][1] ) );
  AND U1531 ( .A(A[658]), .B(B[0]), .Z(\ab[658][0] ) );
  AND U1532 ( .A(B[3]), .B(A[657]), .Z(\ab[657][3] ) );
  AND U1533 ( .A(B[2]), .B(A[657]), .Z(\ab[657][2] ) );
  AND U1534 ( .A(B[1]), .B(A[657]), .Z(\ab[657][1] ) );
  AND U1535 ( .A(A[657]), .B(B[0]), .Z(\ab[657][0] ) );
  AND U1536 ( .A(B[3]), .B(A[656]), .Z(\ab[656][3] ) );
  AND U1537 ( .A(B[2]), .B(A[656]), .Z(\ab[656][2] ) );
  AND U1538 ( .A(B[1]), .B(A[656]), .Z(\ab[656][1] ) );
  AND U1539 ( .A(A[656]), .B(B[0]), .Z(\ab[656][0] ) );
  AND U1540 ( .A(B[3]), .B(A[655]), .Z(\ab[655][3] ) );
  AND U1541 ( .A(B[2]), .B(A[655]), .Z(\ab[655][2] ) );
  AND U1542 ( .A(B[1]), .B(A[655]), .Z(\ab[655][1] ) );
  AND U1543 ( .A(A[655]), .B(B[0]), .Z(\ab[655][0] ) );
  AND U1544 ( .A(B[3]), .B(A[654]), .Z(\ab[654][3] ) );
  AND U1545 ( .A(B[2]), .B(A[654]), .Z(\ab[654][2] ) );
  AND U1546 ( .A(B[1]), .B(A[654]), .Z(\ab[654][1] ) );
  AND U1547 ( .A(A[654]), .B(B[0]), .Z(\ab[654][0] ) );
  AND U1548 ( .A(B[3]), .B(A[653]), .Z(\ab[653][3] ) );
  AND U1549 ( .A(B[2]), .B(A[653]), .Z(\ab[653][2] ) );
  AND U1550 ( .A(B[1]), .B(A[653]), .Z(\ab[653][1] ) );
  AND U1551 ( .A(A[653]), .B(B[0]), .Z(\ab[653][0] ) );
  AND U1552 ( .A(B[3]), .B(A[652]), .Z(\ab[652][3] ) );
  AND U1553 ( .A(B[2]), .B(A[652]), .Z(\ab[652][2] ) );
  AND U1554 ( .A(B[1]), .B(A[652]), .Z(\ab[652][1] ) );
  AND U1555 ( .A(A[652]), .B(B[0]), .Z(\ab[652][0] ) );
  AND U1556 ( .A(B[3]), .B(A[651]), .Z(\ab[651][3] ) );
  AND U1557 ( .A(B[2]), .B(A[651]), .Z(\ab[651][2] ) );
  AND U1558 ( .A(B[1]), .B(A[651]), .Z(\ab[651][1] ) );
  AND U1559 ( .A(A[651]), .B(B[0]), .Z(\ab[651][0] ) );
  AND U1560 ( .A(B[3]), .B(A[650]), .Z(\ab[650][3] ) );
  AND U1561 ( .A(B[2]), .B(A[650]), .Z(\ab[650][2] ) );
  AND U1562 ( .A(B[1]), .B(A[650]), .Z(\ab[650][1] ) );
  AND U1563 ( .A(A[650]), .B(B[0]), .Z(\ab[650][0] ) );
  AND U1564 ( .A(B[3]), .B(A[64]), .Z(\ab[64][3] ) );
  AND U1565 ( .A(B[2]), .B(A[64]), .Z(\ab[64][2] ) );
  AND U1566 ( .A(B[1]), .B(A[64]), .Z(\ab[64][1] ) );
  AND U1567 ( .A(A[64]), .B(B[0]), .Z(\ab[64][0] ) );
  AND U1568 ( .A(B[3]), .B(A[649]), .Z(\ab[649][3] ) );
  AND U1569 ( .A(B[2]), .B(A[649]), .Z(\ab[649][2] ) );
  AND U1570 ( .A(B[1]), .B(A[649]), .Z(\ab[649][1] ) );
  AND U1571 ( .A(A[649]), .B(B[0]), .Z(\ab[649][0] ) );
  AND U1572 ( .A(B[3]), .B(A[648]), .Z(\ab[648][3] ) );
  AND U1573 ( .A(B[2]), .B(A[648]), .Z(\ab[648][2] ) );
  AND U1574 ( .A(B[1]), .B(A[648]), .Z(\ab[648][1] ) );
  AND U1575 ( .A(A[648]), .B(B[0]), .Z(\ab[648][0] ) );
  AND U1576 ( .A(B[3]), .B(A[647]), .Z(\ab[647][3] ) );
  AND U1577 ( .A(B[2]), .B(A[647]), .Z(\ab[647][2] ) );
  AND U1578 ( .A(B[1]), .B(A[647]), .Z(\ab[647][1] ) );
  AND U1579 ( .A(A[647]), .B(B[0]), .Z(\ab[647][0] ) );
  AND U1580 ( .A(B[3]), .B(A[646]), .Z(\ab[646][3] ) );
  AND U1581 ( .A(B[2]), .B(A[646]), .Z(\ab[646][2] ) );
  AND U1582 ( .A(B[1]), .B(A[646]), .Z(\ab[646][1] ) );
  AND U1583 ( .A(A[646]), .B(B[0]), .Z(\ab[646][0] ) );
  AND U1584 ( .A(B[3]), .B(A[645]), .Z(\ab[645][3] ) );
  AND U1585 ( .A(B[2]), .B(A[645]), .Z(\ab[645][2] ) );
  AND U1586 ( .A(B[1]), .B(A[645]), .Z(\ab[645][1] ) );
  AND U1587 ( .A(A[645]), .B(B[0]), .Z(\ab[645][0] ) );
  AND U1588 ( .A(B[3]), .B(A[644]), .Z(\ab[644][3] ) );
  AND U1589 ( .A(B[2]), .B(A[644]), .Z(\ab[644][2] ) );
  AND U1590 ( .A(B[1]), .B(A[644]), .Z(\ab[644][1] ) );
  AND U1591 ( .A(A[644]), .B(B[0]), .Z(\ab[644][0] ) );
  AND U1592 ( .A(B[3]), .B(A[643]), .Z(\ab[643][3] ) );
  AND U1593 ( .A(B[2]), .B(A[643]), .Z(\ab[643][2] ) );
  AND U1594 ( .A(B[1]), .B(A[643]), .Z(\ab[643][1] ) );
  AND U1595 ( .A(A[643]), .B(B[0]), .Z(\ab[643][0] ) );
  AND U1596 ( .A(B[3]), .B(A[642]), .Z(\ab[642][3] ) );
  AND U1597 ( .A(B[2]), .B(A[642]), .Z(\ab[642][2] ) );
  AND U1598 ( .A(B[1]), .B(A[642]), .Z(\ab[642][1] ) );
  AND U1599 ( .A(A[642]), .B(B[0]), .Z(\ab[642][0] ) );
  AND U1600 ( .A(B[3]), .B(A[641]), .Z(\ab[641][3] ) );
  AND U1601 ( .A(B[2]), .B(A[641]), .Z(\ab[641][2] ) );
  AND U1602 ( .A(B[1]), .B(A[641]), .Z(\ab[641][1] ) );
  AND U1603 ( .A(A[641]), .B(B[0]), .Z(\ab[641][0] ) );
  AND U1604 ( .A(B[3]), .B(A[640]), .Z(\ab[640][3] ) );
  AND U1605 ( .A(B[2]), .B(A[640]), .Z(\ab[640][2] ) );
  AND U1606 ( .A(B[1]), .B(A[640]), .Z(\ab[640][1] ) );
  AND U1607 ( .A(A[640]), .B(B[0]), .Z(\ab[640][0] ) );
  AND U1608 ( .A(B[3]), .B(A[63]), .Z(\ab[63][3] ) );
  AND U1609 ( .A(B[2]), .B(A[63]), .Z(\ab[63][2] ) );
  AND U1610 ( .A(B[1]), .B(A[63]), .Z(\ab[63][1] ) );
  AND U1611 ( .A(A[63]), .B(B[0]), .Z(\ab[63][0] ) );
  AND U1612 ( .A(B[3]), .B(A[639]), .Z(\ab[639][3] ) );
  AND U1613 ( .A(B[2]), .B(A[639]), .Z(\ab[639][2] ) );
  AND U1614 ( .A(B[1]), .B(A[639]), .Z(\ab[639][1] ) );
  AND U1615 ( .A(A[639]), .B(B[0]), .Z(\ab[639][0] ) );
  AND U1616 ( .A(B[3]), .B(A[638]), .Z(\ab[638][3] ) );
  AND U1617 ( .A(B[2]), .B(A[638]), .Z(\ab[638][2] ) );
  AND U1618 ( .A(B[1]), .B(A[638]), .Z(\ab[638][1] ) );
  AND U1619 ( .A(A[638]), .B(B[0]), .Z(\ab[638][0] ) );
  AND U1620 ( .A(B[3]), .B(A[637]), .Z(\ab[637][3] ) );
  AND U1621 ( .A(B[2]), .B(A[637]), .Z(\ab[637][2] ) );
  AND U1622 ( .A(B[1]), .B(A[637]), .Z(\ab[637][1] ) );
  AND U1623 ( .A(A[637]), .B(B[0]), .Z(\ab[637][0] ) );
  AND U1624 ( .A(B[3]), .B(A[636]), .Z(\ab[636][3] ) );
  AND U1625 ( .A(B[2]), .B(A[636]), .Z(\ab[636][2] ) );
  AND U1626 ( .A(B[1]), .B(A[636]), .Z(\ab[636][1] ) );
  AND U1627 ( .A(A[636]), .B(B[0]), .Z(\ab[636][0] ) );
  AND U1628 ( .A(B[3]), .B(A[635]), .Z(\ab[635][3] ) );
  AND U1629 ( .A(B[2]), .B(A[635]), .Z(\ab[635][2] ) );
  AND U1630 ( .A(B[1]), .B(A[635]), .Z(\ab[635][1] ) );
  AND U1631 ( .A(A[635]), .B(B[0]), .Z(\ab[635][0] ) );
  AND U1632 ( .A(B[3]), .B(A[634]), .Z(\ab[634][3] ) );
  AND U1633 ( .A(B[2]), .B(A[634]), .Z(\ab[634][2] ) );
  AND U1634 ( .A(B[1]), .B(A[634]), .Z(\ab[634][1] ) );
  AND U1635 ( .A(A[634]), .B(B[0]), .Z(\ab[634][0] ) );
  AND U1636 ( .A(B[3]), .B(A[633]), .Z(\ab[633][3] ) );
  AND U1637 ( .A(B[2]), .B(A[633]), .Z(\ab[633][2] ) );
  AND U1638 ( .A(B[1]), .B(A[633]), .Z(\ab[633][1] ) );
  AND U1639 ( .A(A[633]), .B(B[0]), .Z(\ab[633][0] ) );
  AND U1640 ( .A(B[3]), .B(A[632]), .Z(\ab[632][3] ) );
  AND U1641 ( .A(B[2]), .B(A[632]), .Z(\ab[632][2] ) );
  AND U1642 ( .A(B[1]), .B(A[632]), .Z(\ab[632][1] ) );
  AND U1643 ( .A(A[632]), .B(B[0]), .Z(\ab[632][0] ) );
  AND U1644 ( .A(B[3]), .B(A[631]), .Z(\ab[631][3] ) );
  AND U1645 ( .A(B[2]), .B(A[631]), .Z(\ab[631][2] ) );
  AND U1646 ( .A(B[1]), .B(A[631]), .Z(\ab[631][1] ) );
  AND U1647 ( .A(A[631]), .B(B[0]), .Z(\ab[631][0] ) );
  AND U1648 ( .A(B[3]), .B(A[630]), .Z(\ab[630][3] ) );
  AND U1649 ( .A(B[2]), .B(A[630]), .Z(\ab[630][2] ) );
  AND U1650 ( .A(B[1]), .B(A[630]), .Z(\ab[630][1] ) );
  AND U1651 ( .A(A[630]), .B(B[0]), .Z(\ab[630][0] ) );
  AND U1652 ( .A(B[3]), .B(A[62]), .Z(\ab[62][3] ) );
  AND U1653 ( .A(B[2]), .B(A[62]), .Z(\ab[62][2] ) );
  AND U1654 ( .A(B[1]), .B(A[62]), .Z(\ab[62][1] ) );
  AND U1655 ( .A(A[62]), .B(B[0]), .Z(\ab[62][0] ) );
  AND U1656 ( .A(B[3]), .B(A[629]), .Z(\ab[629][3] ) );
  AND U1657 ( .A(B[2]), .B(A[629]), .Z(\ab[629][2] ) );
  AND U1658 ( .A(B[1]), .B(A[629]), .Z(\ab[629][1] ) );
  AND U1659 ( .A(A[629]), .B(B[0]), .Z(\ab[629][0] ) );
  AND U1660 ( .A(B[3]), .B(A[628]), .Z(\ab[628][3] ) );
  AND U1661 ( .A(B[2]), .B(A[628]), .Z(\ab[628][2] ) );
  AND U1662 ( .A(B[1]), .B(A[628]), .Z(\ab[628][1] ) );
  AND U1663 ( .A(A[628]), .B(B[0]), .Z(\ab[628][0] ) );
  AND U1664 ( .A(B[3]), .B(A[627]), .Z(\ab[627][3] ) );
  AND U1665 ( .A(B[2]), .B(A[627]), .Z(\ab[627][2] ) );
  AND U1666 ( .A(B[1]), .B(A[627]), .Z(\ab[627][1] ) );
  AND U1667 ( .A(A[627]), .B(B[0]), .Z(\ab[627][0] ) );
  AND U1668 ( .A(B[3]), .B(A[626]), .Z(\ab[626][3] ) );
  AND U1669 ( .A(B[2]), .B(A[626]), .Z(\ab[626][2] ) );
  AND U1670 ( .A(B[1]), .B(A[626]), .Z(\ab[626][1] ) );
  AND U1671 ( .A(A[626]), .B(B[0]), .Z(\ab[626][0] ) );
  AND U1672 ( .A(B[3]), .B(A[625]), .Z(\ab[625][3] ) );
  AND U1673 ( .A(B[2]), .B(A[625]), .Z(\ab[625][2] ) );
  AND U1674 ( .A(B[1]), .B(A[625]), .Z(\ab[625][1] ) );
  AND U1675 ( .A(A[625]), .B(B[0]), .Z(\ab[625][0] ) );
  AND U1676 ( .A(B[3]), .B(A[624]), .Z(\ab[624][3] ) );
  AND U1677 ( .A(B[2]), .B(A[624]), .Z(\ab[624][2] ) );
  AND U1678 ( .A(B[1]), .B(A[624]), .Z(\ab[624][1] ) );
  AND U1679 ( .A(A[624]), .B(B[0]), .Z(\ab[624][0] ) );
  AND U1680 ( .A(B[3]), .B(A[623]), .Z(\ab[623][3] ) );
  AND U1681 ( .A(B[2]), .B(A[623]), .Z(\ab[623][2] ) );
  AND U1682 ( .A(B[1]), .B(A[623]), .Z(\ab[623][1] ) );
  AND U1683 ( .A(A[623]), .B(B[0]), .Z(\ab[623][0] ) );
  AND U1684 ( .A(B[3]), .B(A[622]), .Z(\ab[622][3] ) );
  AND U1685 ( .A(B[2]), .B(A[622]), .Z(\ab[622][2] ) );
  AND U1686 ( .A(B[1]), .B(A[622]), .Z(\ab[622][1] ) );
  AND U1687 ( .A(A[622]), .B(B[0]), .Z(\ab[622][0] ) );
  AND U1688 ( .A(B[3]), .B(A[621]), .Z(\ab[621][3] ) );
  AND U1689 ( .A(B[2]), .B(A[621]), .Z(\ab[621][2] ) );
  AND U1690 ( .A(B[1]), .B(A[621]), .Z(\ab[621][1] ) );
  AND U1691 ( .A(A[621]), .B(B[0]), .Z(\ab[621][0] ) );
  AND U1692 ( .A(B[3]), .B(A[620]), .Z(\ab[620][3] ) );
  AND U1693 ( .A(B[2]), .B(A[620]), .Z(\ab[620][2] ) );
  AND U1694 ( .A(B[1]), .B(A[620]), .Z(\ab[620][1] ) );
  AND U1695 ( .A(A[620]), .B(B[0]), .Z(\ab[620][0] ) );
  AND U1696 ( .A(B[3]), .B(A[61]), .Z(\ab[61][3] ) );
  AND U1697 ( .A(B[2]), .B(A[61]), .Z(\ab[61][2] ) );
  AND U1698 ( .A(B[1]), .B(A[61]), .Z(\ab[61][1] ) );
  AND U1699 ( .A(A[61]), .B(B[0]), .Z(\ab[61][0] ) );
  AND U1700 ( .A(B[3]), .B(A[619]), .Z(\ab[619][3] ) );
  AND U1701 ( .A(B[2]), .B(A[619]), .Z(\ab[619][2] ) );
  AND U1702 ( .A(B[1]), .B(A[619]), .Z(\ab[619][1] ) );
  AND U1703 ( .A(A[619]), .B(B[0]), .Z(\ab[619][0] ) );
  AND U1704 ( .A(B[3]), .B(A[618]), .Z(\ab[618][3] ) );
  AND U1705 ( .A(B[2]), .B(A[618]), .Z(\ab[618][2] ) );
  AND U1706 ( .A(B[1]), .B(A[618]), .Z(\ab[618][1] ) );
  AND U1707 ( .A(A[618]), .B(B[0]), .Z(\ab[618][0] ) );
  AND U1708 ( .A(B[3]), .B(A[617]), .Z(\ab[617][3] ) );
  AND U1709 ( .A(B[2]), .B(A[617]), .Z(\ab[617][2] ) );
  AND U1710 ( .A(B[1]), .B(A[617]), .Z(\ab[617][1] ) );
  AND U1711 ( .A(A[617]), .B(B[0]), .Z(\ab[617][0] ) );
  AND U1712 ( .A(B[3]), .B(A[616]), .Z(\ab[616][3] ) );
  AND U1713 ( .A(B[2]), .B(A[616]), .Z(\ab[616][2] ) );
  AND U1714 ( .A(B[1]), .B(A[616]), .Z(\ab[616][1] ) );
  AND U1715 ( .A(A[616]), .B(B[0]), .Z(\ab[616][0] ) );
  AND U1716 ( .A(B[3]), .B(A[615]), .Z(\ab[615][3] ) );
  AND U1717 ( .A(B[2]), .B(A[615]), .Z(\ab[615][2] ) );
  AND U1718 ( .A(B[1]), .B(A[615]), .Z(\ab[615][1] ) );
  AND U1719 ( .A(A[615]), .B(B[0]), .Z(\ab[615][0] ) );
  AND U1720 ( .A(B[3]), .B(A[614]), .Z(\ab[614][3] ) );
  AND U1721 ( .A(B[2]), .B(A[614]), .Z(\ab[614][2] ) );
  AND U1722 ( .A(B[1]), .B(A[614]), .Z(\ab[614][1] ) );
  AND U1723 ( .A(A[614]), .B(B[0]), .Z(\ab[614][0] ) );
  AND U1724 ( .A(B[3]), .B(A[613]), .Z(\ab[613][3] ) );
  AND U1725 ( .A(B[2]), .B(A[613]), .Z(\ab[613][2] ) );
  AND U1726 ( .A(B[1]), .B(A[613]), .Z(\ab[613][1] ) );
  AND U1727 ( .A(A[613]), .B(B[0]), .Z(\ab[613][0] ) );
  AND U1728 ( .A(B[3]), .B(A[612]), .Z(\ab[612][3] ) );
  AND U1729 ( .A(B[2]), .B(A[612]), .Z(\ab[612][2] ) );
  AND U1730 ( .A(B[1]), .B(A[612]), .Z(\ab[612][1] ) );
  AND U1731 ( .A(A[612]), .B(B[0]), .Z(\ab[612][0] ) );
  AND U1732 ( .A(B[3]), .B(A[611]), .Z(\ab[611][3] ) );
  AND U1733 ( .A(B[2]), .B(A[611]), .Z(\ab[611][2] ) );
  AND U1734 ( .A(B[1]), .B(A[611]), .Z(\ab[611][1] ) );
  AND U1735 ( .A(A[611]), .B(B[0]), .Z(\ab[611][0] ) );
  AND U1736 ( .A(B[3]), .B(A[610]), .Z(\ab[610][3] ) );
  AND U1737 ( .A(B[2]), .B(A[610]), .Z(\ab[610][2] ) );
  AND U1738 ( .A(B[1]), .B(A[610]), .Z(\ab[610][1] ) );
  AND U1739 ( .A(A[610]), .B(B[0]), .Z(\ab[610][0] ) );
  AND U1740 ( .A(B[3]), .B(A[60]), .Z(\ab[60][3] ) );
  AND U1741 ( .A(B[2]), .B(A[60]), .Z(\ab[60][2] ) );
  AND U1742 ( .A(B[1]), .B(A[60]), .Z(\ab[60][1] ) );
  AND U1743 ( .A(A[60]), .B(B[0]), .Z(\ab[60][0] ) );
  AND U1744 ( .A(B[3]), .B(A[609]), .Z(\ab[609][3] ) );
  AND U1745 ( .A(B[2]), .B(A[609]), .Z(\ab[609][2] ) );
  AND U1746 ( .A(B[1]), .B(A[609]), .Z(\ab[609][1] ) );
  AND U1747 ( .A(A[609]), .B(B[0]), .Z(\ab[609][0] ) );
  AND U1748 ( .A(B[3]), .B(A[608]), .Z(\ab[608][3] ) );
  AND U1749 ( .A(B[2]), .B(A[608]), .Z(\ab[608][2] ) );
  AND U1750 ( .A(B[1]), .B(A[608]), .Z(\ab[608][1] ) );
  AND U1751 ( .A(A[608]), .B(B[0]), .Z(\ab[608][0] ) );
  AND U1752 ( .A(B[3]), .B(A[607]), .Z(\ab[607][3] ) );
  AND U1753 ( .A(B[2]), .B(A[607]), .Z(\ab[607][2] ) );
  AND U1754 ( .A(B[1]), .B(A[607]), .Z(\ab[607][1] ) );
  AND U1755 ( .A(A[607]), .B(B[0]), .Z(\ab[607][0] ) );
  AND U1756 ( .A(B[3]), .B(A[606]), .Z(\ab[606][3] ) );
  AND U1757 ( .A(B[2]), .B(A[606]), .Z(\ab[606][2] ) );
  AND U1758 ( .A(B[1]), .B(A[606]), .Z(\ab[606][1] ) );
  AND U1759 ( .A(A[606]), .B(B[0]), .Z(\ab[606][0] ) );
  AND U1760 ( .A(B[3]), .B(A[605]), .Z(\ab[605][3] ) );
  AND U1761 ( .A(B[2]), .B(A[605]), .Z(\ab[605][2] ) );
  AND U1762 ( .A(B[1]), .B(A[605]), .Z(\ab[605][1] ) );
  AND U1763 ( .A(A[605]), .B(B[0]), .Z(\ab[605][0] ) );
  AND U1764 ( .A(B[3]), .B(A[604]), .Z(\ab[604][3] ) );
  AND U1765 ( .A(B[2]), .B(A[604]), .Z(\ab[604][2] ) );
  AND U1766 ( .A(B[1]), .B(A[604]), .Z(\ab[604][1] ) );
  AND U1767 ( .A(A[604]), .B(B[0]), .Z(\ab[604][0] ) );
  AND U1768 ( .A(B[3]), .B(A[603]), .Z(\ab[603][3] ) );
  AND U1769 ( .A(B[2]), .B(A[603]), .Z(\ab[603][2] ) );
  AND U1770 ( .A(B[1]), .B(A[603]), .Z(\ab[603][1] ) );
  AND U1771 ( .A(A[603]), .B(B[0]), .Z(\ab[603][0] ) );
  AND U1772 ( .A(B[3]), .B(A[602]), .Z(\ab[602][3] ) );
  AND U1773 ( .A(B[2]), .B(A[602]), .Z(\ab[602][2] ) );
  AND U1774 ( .A(B[1]), .B(A[602]), .Z(\ab[602][1] ) );
  AND U1775 ( .A(A[602]), .B(B[0]), .Z(\ab[602][0] ) );
  AND U1776 ( .A(B[3]), .B(A[601]), .Z(\ab[601][3] ) );
  AND U1777 ( .A(B[2]), .B(A[601]), .Z(\ab[601][2] ) );
  AND U1778 ( .A(B[1]), .B(A[601]), .Z(\ab[601][1] ) );
  AND U1779 ( .A(A[601]), .B(B[0]), .Z(\ab[601][0] ) );
  AND U1780 ( .A(B[3]), .B(A[600]), .Z(\ab[600][3] ) );
  AND U1781 ( .A(B[2]), .B(A[600]), .Z(\ab[600][2] ) );
  AND U1782 ( .A(B[1]), .B(A[600]), .Z(\ab[600][1] ) );
  AND U1783 ( .A(A[600]), .B(B[0]), .Z(\ab[600][0] ) );
  AND U1784 ( .A(B[3]), .B(A[5]), .Z(\ab[5][3] ) );
  AND U1785 ( .A(B[2]), .B(A[5]), .Z(\ab[5][2] ) );
  AND U1786 ( .A(B[1]), .B(A[5]), .Z(\ab[5][1] ) );
  AND U1787 ( .A(A[5]), .B(B[0]), .Z(\ab[5][0] ) );
  AND U1788 ( .A(B[3]), .B(A[59]), .Z(\ab[59][3] ) );
  AND U1789 ( .A(B[2]), .B(A[59]), .Z(\ab[59][2] ) );
  AND U1790 ( .A(B[1]), .B(A[59]), .Z(\ab[59][1] ) );
  AND U1791 ( .A(A[59]), .B(B[0]), .Z(\ab[59][0] ) );
  AND U1792 ( .A(B[3]), .B(A[599]), .Z(\ab[599][3] ) );
  AND U1793 ( .A(B[2]), .B(A[599]), .Z(\ab[599][2] ) );
  AND U1794 ( .A(B[1]), .B(A[599]), .Z(\ab[599][1] ) );
  AND U1795 ( .A(A[599]), .B(B[0]), .Z(\ab[599][0] ) );
  AND U1796 ( .A(B[3]), .B(A[598]), .Z(\ab[598][3] ) );
  AND U1797 ( .A(B[2]), .B(A[598]), .Z(\ab[598][2] ) );
  AND U1798 ( .A(B[1]), .B(A[598]), .Z(\ab[598][1] ) );
  AND U1799 ( .A(A[598]), .B(B[0]), .Z(\ab[598][0] ) );
  AND U1800 ( .A(B[3]), .B(A[597]), .Z(\ab[597][3] ) );
  AND U1801 ( .A(B[2]), .B(A[597]), .Z(\ab[597][2] ) );
  AND U1802 ( .A(B[1]), .B(A[597]), .Z(\ab[597][1] ) );
  AND U1803 ( .A(A[597]), .B(B[0]), .Z(\ab[597][0] ) );
  AND U1804 ( .A(B[3]), .B(A[596]), .Z(\ab[596][3] ) );
  AND U1805 ( .A(B[2]), .B(A[596]), .Z(\ab[596][2] ) );
  AND U1806 ( .A(B[1]), .B(A[596]), .Z(\ab[596][1] ) );
  AND U1807 ( .A(A[596]), .B(B[0]), .Z(\ab[596][0] ) );
  AND U1808 ( .A(B[3]), .B(A[595]), .Z(\ab[595][3] ) );
  AND U1809 ( .A(B[2]), .B(A[595]), .Z(\ab[595][2] ) );
  AND U1810 ( .A(B[1]), .B(A[595]), .Z(\ab[595][1] ) );
  AND U1811 ( .A(A[595]), .B(B[0]), .Z(\ab[595][0] ) );
  AND U1812 ( .A(B[3]), .B(A[594]), .Z(\ab[594][3] ) );
  AND U1813 ( .A(B[2]), .B(A[594]), .Z(\ab[594][2] ) );
  AND U1814 ( .A(B[1]), .B(A[594]), .Z(\ab[594][1] ) );
  AND U1815 ( .A(A[594]), .B(B[0]), .Z(\ab[594][0] ) );
  AND U1816 ( .A(B[3]), .B(A[593]), .Z(\ab[593][3] ) );
  AND U1817 ( .A(B[2]), .B(A[593]), .Z(\ab[593][2] ) );
  AND U1818 ( .A(B[1]), .B(A[593]), .Z(\ab[593][1] ) );
  AND U1819 ( .A(A[593]), .B(B[0]), .Z(\ab[593][0] ) );
  AND U1820 ( .A(B[3]), .B(A[592]), .Z(\ab[592][3] ) );
  AND U1821 ( .A(B[2]), .B(A[592]), .Z(\ab[592][2] ) );
  AND U1822 ( .A(B[1]), .B(A[592]), .Z(\ab[592][1] ) );
  AND U1823 ( .A(A[592]), .B(B[0]), .Z(\ab[592][0] ) );
  AND U1824 ( .A(B[3]), .B(A[591]), .Z(\ab[591][3] ) );
  AND U1825 ( .A(B[2]), .B(A[591]), .Z(\ab[591][2] ) );
  AND U1826 ( .A(B[1]), .B(A[591]), .Z(\ab[591][1] ) );
  AND U1827 ( .A(A[591]), .B(B[0]), .Z(\ab[591][0] ) );
  AND U1828 ( .A(B[3]), .B(A[590]), .Z(\ab[590][3] ) );
  AND U1829 ( .A(B[2]), .B(A[590]), .Z(\ab[590][2] ) );
  AND U1830 ( .A(B[1]), .B(A[590]), .Z(\ab[590][1] ) );
  AND U1831 ( .A(A[590]), .B(B[0]), .Z(\ab[590][0] ) );
  AND U1832 ( .A(B[3]), .B(A[58]), .Z(\ab[58][3] ) );
  AND U1833 ( .A(B[2]), .B(A[58]), .Z(\ab[58][2] ) );
  AND U1834 ( .A(B[1]), .B(A[58]), .Z(\ab[58][1] ) );
  AND U1835 ( .A(A[58]), .B(B[0]), .Z(\ab[58][0] ) );
  AND U1836 ( .A(B[3]), .B(A[589]), .Z(\ab[589][3] ) );
  AND U1837 ( .A(B[2]), .B(A[589]), .Z(\ab[589][2] ) );
  AND U1838 ( .A(B[1]), .B(A[589]), .Z(\ab[589][1] ) );
  AND U1839 ( .A(A[589]), .B(B[0]), .Z(\ab[589][0] ) );
  AND U1840 ( .A(B[3]), .B(A[588]), .Z(\ab[588][3] ) );
  AND U1841 ( .A(B[2]), .B(A[588]), .Z(\ab[588][2] ) );
  AND U1842 ( .A(B[1]), .B(A[588]), .Z(\ab[588][1] ) );
  AND U1843 ( .A(A[588]), .B(B[0]), .Z(\ab[588][0] ) );
  AND U1844 ( .A(B[3]), .B(A[587]), .Z(\ab[587][3] ) );
  AND U1845 ( .A(B[2]), .B(A[587]), .Z(\ab[587][2] ) );
  AND U1846 ( .A(B[1]), .B(A[587]), .Z(\ab[587][1] ) );
  AND U1847 ( .A(A[587]), .B(B[0]), .Z(\ab[587][0] ) );
  AND U1848 ( .A(B[3]), .B(A[586]), .Z(\ab[586][3] ) );
  AND U1849 ( .A(B[2]), .B(A[586]), .Z(\ab[586][2] ) );
  AND U1850 ( .A(B[1]), .B(A[586]), .Z(\ab[586][1] ) );
  AND U1851 ( .A(A[586]), .B(B[0]), .Z(\ab[586][0] ) );
  AND U1852 ( .A(B[3]), .B(A[585]), .Z(\ab[585][3] ) );
  AND U1853 ( .A(B[2]), .B(A[585]), .Z(\ab[585][2] ) );
  AND U1854 ( .A(B[1]), .B(A[585]), .Z(\ab[585][1] ) );
  AND U1855 ( .A(A[585]), .B(B[0]), .Z(\ab[585][0] ) );
  AND U1856 ( .A(B[3]), .B(A[584]), .Z(\ab[584][3] ) );
  AND U1857 ( .A(B[2]), .B(A[584]), .Z(\ab[584][2] ) );
  AND U1858 ( .A(B[1]), .B(A[584]), .Z(\ab[584][1] ) );
  AND U1859 ( .A(A[584]), .B(B[0]), .Z(\ab[584][0] ) );
  AND U1860 ( .A(B[3]), .B(A[583]), .Z(\ab[583][3] ) );
  AND U1861 ( .A(B[2]), .B(A[583]), .Z(\ab[583][2] ) );
  AND U1862 ( .A(B[1]), .B(A[583]), .Z(\ab[583][1] ) );
  AND U1863 ( .A(A[583]), .B(B[0]), .Z(\ab[583][0] ) );
  AND U1864 ( .A(B[3]), .B(A[582]), .Z(\ab[582][3] ) );
  AND U1865 ( .A(B[2]), .B(A[582]), .Z(\ab[582][2] ) );
  AND U1866 ( .A(B[1]), .B(A[582]), .Z(\ab[582][1] ) );
  AND U1867 ( .A(A[582]), .B(B[0]), .Z(\ab[582][0] ) );
  AND U1868 ( .A(B[3]), .B(A[581]), .Z(\ab[581][3] ) );
  AND U1869 ( .A(B[2]), .B(A[581]), .Z(\ab[581][2] ) );
  AND U1870 ( .A(B[1]), .B(A[581]), .Z(\ab[581][1] ) );
  AND U1871 ( .A(A[581]), .B(B[0]), .Z(\ab[581][0] ) );
  AND U1872 ( .A(B[3]), .B(A[580]), .Z(\ab[580][3] ) );
  AND U1873 ( .A(B[2]), .B(A[580]), .Z(\ab[580][2] ) );
  AND U1874 ( .A(B[1]), .B(A[580]), .Z(\ab[580][1] ) );
  AND U1875 ( .A(A[580]), .B(B[0]), .Z(\ab[580][0] ) );
  AND U1876 ( .A(B[3]), .B(A[57]), .Z(\ab[57][3] ) );
  AND U1877 ( .A(B[2]), .B(A[57]), .Z(\ab[57][2] ) );
  AND U1878 ( .A(B[1]), .B(A[57]), .Z(\ab[57][1] ) );
  AND U1879 ( .A(A[57]), .B(B[0]), .Z(\ab[57][0] ) );
  AND U1880 ( .A(B[3]), .B(A[579]), .Z(\ab[579][3] ) );
  AND U1881 ( .A(B[2]), .B(A[579]), .Z(\ab[579][2] ) );
  AND U1882 ( .A(B[1]), .B(A[579]), .Z(\ab[579][1] ) );
  AND U1883 ( .A(A[579]), .B(B[0]), .Z(\ab[579][0] ) );
  AND U1884 ( .A(B[3]), .B(A[578]), .Z(\ab[578][3] ) );
  AND U1885 ( .A(B[2]), .B(A[578]), .Z(\ab[578][2] ) );
  AND U1886 ( .A(B[1]), .B(A[578]), .Z(\ab[578][1] ) );
  AND U1887 ( .A(A[578]), .B(B[0]), .Z(\ab[578][0] ) );
  AND U1888 ( .A(B[3]), .B(A[577]), .Z(\ab[577][3] ) );
  AND U1889 ( .A(B[2]), .B(A[577]), .Z(\ab[577][2] ) );
  AND U1890 ( .A(B[1]), .B(A[577]), .Z(\ab[577][1] ) );
  AND U1891 ( .A(A[577]), .B(B[0]), .Z(\ab[577][0] ) );
  AND U1892 ( .A(B[3]), .B(A[576]), .Z(\ab[576][3] ) );
  AND U1893 ( .A(B[2]), .B(A[576]), .Z(\ab[576][2] ) );
  AND U1894 ( .A(B[1]), .B(A[576]), .Z(\ab[576][1] ) );
  AND U1895 ( .A(A[576]), .B(B[0]), .Z(\ab[576][0] ) );
  AND U1896 ( .A(B[3]), .B(A[575]), .Z(\ab[575][3] ) );
  AND U1897 ( .A(B[2]), .B(A[575]), .Z(\ab[575][2] ) );
  AND U1898 ( .A(B[1]), .B(A[575]), .Z(\ab[575][1] ) );
  AND U1899 ( .A(A[575]), .B(B[0]), .Z(\ab[575][0] ) );
  AND U1900 ( .A(B[3]), .B(A[574]), .Z(\ab[574][3] ) );
  AND U1901 ( .A(B[2]), .B(A[574]), .Z(\ab[574][2] ) );
  AND U1902 ( .A(B[1]), .B(A[574]), .Z(\ab[574][1] ) );
  AND U1903 ( .A(A[574]), .B(B[0]), .Z(\ab[574][0] ) );
  AND U1904 ( .A(B[3]), .B(A[573]), .Z(\ab[573][3] ) );
  AND U1905 ( .A(B[2]), .B(A[573]), .Z(\ab[573][2] ) );
  AND U1906 ( .A(B[1]), .B(A[573]), .Z(\ab[573][1] ) );
  AND U1907 ( .A(A[573]), .B(B[0]), .Z(\ab[573][0] ) );
  AND U1908 ( .A(B[3]), .B(A[572]), .Z(\ab[572][3] ) );
  AND U1909 ( .A(B[2]), .B(A[572]), .Z(\ab[572][2] ) );
  AND U1910 ( .A(B[1]), .B(A[572]), .Z(\ab[572][1] ) );
  AND U1911 ( .A(A[572]), .B(B[0]), .Z(\ab[572][0] ) );
  AND U1912 ( .A(B[3]), .B(A[571]), .Z(\ab[571][3] ) );
  AND U1913 ( .A(B[2]), .B(A[571]), .Z(\ab[571][2] ) );
  AND U1914 ( .A(B[1]), .B(A[571]), .Z(\ab[571][1] ) );
  AND U1915 ( .A(A[571]), .B(B[0]), .Z(\ab[571][0] ) );
  AND U1916 ( .A(B[3]), .B(A[570]), .Z(\ab[570][3] ) );
  AND U1917 ( .A(B[2]), .B(A[570]), .Z(\ab[570][2] ) );
  AND U1918 ( .A(B[1]), .B(A[570]), .Z(\ab[570][1] ) );
  AND U1919 ( .A(A[570]), .B(B[0]), .Z(\ab[570][0] ) );
  AND U1920 ( .A(B[3]), .B(A[56]), .Z(\ab[56][3] ) );
  AND U1921 ( .A(B[2]), .B(A[56]), .Z(\ab[56][2] ) );
  AND U1922 ( .A(B[1]), .B(A[56]), .Z(\ab[56][1] ) );
  AND U1923 ( .A(A[56]), .B(B[0]), .Z(\ab[56][0] ) );
  AND U1924 ( .A(B[3]), .B(A[569]), .Z(\ab[569][3] ) );
  AND U1925 ( .A(B[2]), .B(A[569]), .Z(\ab[569][2] ) );
  AND U1926 ( .A(B[1]), .B(A[569]), .Z(\ab[569][1] ) );
  AND U1927 ( .A(A[569]), .B(B[0]), .Z(\ab[569][0] ) );
  AND U1928 ( .A(B[3]), .B(A[568]), .Z(\ab[568][3] ) );
  AND U1929 ( .A(B[2]), .B(A[568]), .Z(\ab[568][2] ) );
  AND U1930 ( .A(B[1]), .B(A[568]), .Z(\ab[568][1] ) );
  AND U1931 ( .A(A[568]), .B(B[0]), .Z(\ab[568][0] ) );
  AND U1932 ( .A(B[3]), .B(A[567]), .Z(\ab[567][3] ) );
  AND U1933 ( .A(B[2]), .B(A[567]), .Z(\ab[567][2] ) );
  AND U1934 ( .A(B[1]), .B(A[567]), .Z(\ab[567][1] ) );
  AND U1935 ( .A(A[567]), .B(B[0]), .Z(\ab[567][0] ) );
  AND U1936 ( .A(B[3]), .B(A[566]), .Z(\ab[566][3] ) );
  AND U1937 ( .A(B[2]), .B(A[566]), .Z(\ab[566][2] ) );
  AND U1938 ( .A(B[1]), .B(A[566]), .Z(\ab[566][1] ) );
  AND U1939 ( .A(A[566]), .B(B[0]), .Z(\ab[566][0] ) );
  AND U1940 ( .A(B[3]), .B(A[565]), .Z(\ab[565][3] ) );
  AND U1941 ( .A(B[2]), .B(A[565]), .Z(\ab[565][2] ) );
  AND U1942 ( .A(B[1]), .B(A[565]), .Z(\ab[565][1] ) );
  AND U1943 ( .A(A[565]), .B(B[0]), .Z(\ab[565][0] ) );
  AND U1944 ( .A(B[3]), .B(A[564]), .Z(\ab[564][3] ) );
  AND U1945 ( .A(B[2]), .B(A[564]), .Z(\ab[564][2] ) );
  AND U1946 ( .A(B[1]), .B(A[564]), .Z(\ab[564][1] ) );
  AND U1947 ( .A(A[564]), .B(B[0]), .Z(\ab[564][0] ) );
  AND U1948 ( .A(B[3]), .B(A[563]), .Z(\ab[563][3] ) );
  AND U1949 ( .A(B[2]), .B(A[563]), .Z(\ab[563][2] ) );
  AND U1950 ( .A(B[1]), .B(A[563]), .Z(\ab[563][1] ) );
  AND U1951 ( .A(A[563]), .B(B[0]), .Z(\ab[563][0] ) );
  AND U1952 ( .A(B[3]), .B(A[562]), .Z(\ab[562][3] ) );
  AND U1953 ( .A(B[2]), .B(A[562]), .Z(\ab[562][2] ) );
  AND U1954 ( .A(B[1]), .B(A[562]), .Z(\ab[562][1] ) );
  AND U1955 ( .A(A[562]), .B(B[0]), .Z(\ab[562][0] ) );
  AND U1956 ( .A(B[3]), .B(A[561]), .Z(\ab[561][3] ) );
  AND U1957 ( .A(B[2]), .B(A[561]), .Z(\ab[561][2] ) );
  AND U1958 ( .A(B[1]), .B(A[561]), .Z(\ab[561][1] ) );
  AND U1959 ( .A(A[561]), .B(B[0]), .Z(\ab[561][0] ) );
  AND U1960 ( .A(B[3]), .B(A[560]), .Z(\ab[560][3] ) );
  AND U1961 ( .A(B[2]), .B(A[560]), .Z(\ab[560][2] ) );
  AND U1962 ( .A(B[1]), .B(A[560]), .Z(\ab[560][1] ) );
  AND U1963 ( .A(A[560]), .B(B[0]), .Z(\ab[560][0] ) );
  AND U1964 ( .A(B[3]), .B(A[55]), .Z(\ab[55][3] ) );
  AND U1965 ( .A(B[2]), .B(A[55]), .Z(\ab[55][2] ) );
  AND U1966 ( .A(B[1]), .B(A[55]), .Z(\ab[55][1] ) );
  AND U1967 ( .A(A[55]), .B(B[0]), .Z(\ab[55][0] ) );
  AND U1968 ( .A(B[3]), .B(A[559]), .Z(\ab[559][3] ) );
  AND U1969 ( .A(B[2]), .B(A[559]), .Z(\ab[559][2] ) );
  AND U1970 ( .A(B[1]), .B(A[559]), .Z(\ab[559][1] ) );
  AND U1971 ( .A(A[559]), .B(B[0]), .Z(\ab[559][0] ) );
  AND U1972 ( .A(B[3]), .B(A[558]), .Z(\ab[558][3] ) );
  AND U1973 ( .A(B[2]), .B(A[558]), .Z(\ab[558][2] ) );
  AND U1974 ( .A(B[1]), .B(A[558]), .Z(\ab[558][1] ) );
  AND U1975 ( .A(A[558]), .B(B[0]), .Z(\ab[558][0] ) );
  AND U1976 ( .A(B[3]), .B(A[557]), .Z(\ab[557][3] ) );
  AND U1977 ( .A(B[2]), .B(A[557]), .Z(\ab[557][2] ) );
  AND U1978 ( .A(B[1]), .B(A[557]), .Z(\ab[557][1] ) );
  AND U1979 ( .A(A[557]), .B(B[0]), .Z(\ab[557][0] ) );
  AND U1980 ( .A(B[3]), .B(A[556]), .Z(\ab[556][3] ) );
  AND U1981 ( .A(B[2]), .B(A[556]), .Z(\ab[556][2] ) );
  AND U1982 ( .A(B[1]), .B(A[556]), .Z(\ab[556][1] ) );
  AND U1983 ( .A(A[556]), .B(B[0]), .Z(\ab[556][0] ) );
  AND U1984 ( .A(B[3]), .B(A[555]), .Z(\ab[555][3] ) );
  AND U1985 ( .A(B[2]), .B(A[555]), .Z(\ab[555][2] ) );
  AND U1986 ( .A(B[1]), .B(A[555]), .Z(\ab[555][1] ) );
  AND U1987 ( .A(A[555]), .B(B[0]), .Z(\ab[555][0] ) );
  AND U1988 ( .A(B[3]), .B(A[554]), .Z(\ab[554][3] ) );
  AND U1989 ( .A(B[2]), .B(A[554]), .Z(\ab[554][2] ) );
  AND U1990 ( .A(B[1]), .B(A[554]), .Z(\ab[554][1] ) );
  AND U1991 ( .A(A[554]), .B(B[0]), .Z(\ab[554][0] ) );
  AND U1992 ( .A(B[3]), .B(A[553]), .Z(\ab[553][3] ) );
  AND U1993 ( .A(B[2]), .B(A[553]), .Z(\ab[553][2] ) );
  AND U1994 ( .A(B[1]), .B(A[553]), .Z(\ab[553][1] ) );
  AND U1995 ( .A(A[553]), .B(B[0]), .Z(\ab[553][0] ) );
  AND U1996 ( .A(B[3]), .B(A[552]), .Z(\ab[552][3] ) );
  AND U1997 ( .A(B[2]), .B(A[552]), .Z(\ab[552][2] ) );
  AND U1998 ( .A(B[1]), .B(A[552]), .Z(\ab[552][1] ) );
  AND U1999 ( .A(A[552]), .B(B[0]), .Z(\ab[552][0] ) );
  AND U2000 ( .A(B[3]), .B(A[551]), .Z(\ab[551][3] ) );
  AND U2001 ( .A(B[2]), .B(A[551]), .Z(\ab[551][2] ) );
  AND U2002 ( .A(B[1]), .B(A[551]), .Z(\ab[551][1] ) );
  AND U2003 ( .A(A[551]), .B(B[0]), .Z(\ab[551][0] ) );
  AND U2004 ( .A(B[3]), .B(A[550]), .Z(\ab[550][3] ) );
  AND U2005 ( .A(B[2]), .B(A[550]), .Z(\ab[550][2] ) );
  AND U2006 ( .A(B[1]), .B(A[550]), .Z(\ab[550][1] ) );
  AND U2007 ( .A(A[550]), .B(B[0]), .Z(\ab[550][0] ) );
  AND U2008 ( .A(B[3]), .B(A[54]), .Z(\ab[54][3] ) );
  AND U2009 ( .A(B[2]), .B(A[54]), .Z(\ab[54][2] ) );
  AND U2010 ( .A(B[1]), .B(A[54]), .Z(\ab[54][1] ) );
  AND U2011 ( .A(A[54]), .B(B[0]), .Z(\ab[54][0] ) );
  AND U2012 ( .A(B[3]), .B(A[549]), .Z(\ab[549][3] ) );
  AND U2013 ( .A(B[2]), .B(A[549]), .Z(\ab[549][2] ) );
  AND U2014 ( .A(B[1]), .B(A[549]), .Z(\ab[549][1] ) );
  AND U2015 ( .A(A[549]), .B(B[0]), .Z(\ab[549][0] ) );
  AND U2016 ( .A(B[3]), .B(A[548]), .Z(\ab[548][3] ) );
  AND U2017 ( .A(B[2]), .B(A[548]), .Z(\ab[548][2] ) );
  AND U2018 ( .A(B[1]), .B(A[548]), .Z(\ab[548][1] ) );
  AND U2019 ( .A(A[548]), .B(B[0]), .Z(\ab[548][0] ) );
  AND U2020 ( .A(B[3]), .B(A[547]), .Z(\ab[547][3] ) );
  AND U2021 ( .A(B[2]), .B(A[547]), .Z(\ab[547][2] ) );
  AND U2022 ( .A(B[1]), .B(A[547]), .Z(\ab[547][1] ) );
  AND U2023 ( .A(A[547]), .B(B[0]), .Z(\ab[547][0] ) );
  AND U2024 ( .A(B[3]), .B(A[546]), .Z(\ab[546][3] ) );
  AND U2025 ( .A(B[2]), .B(A[546]), .Z(\ab[546][2] ) );
  AND U2026 ( .A(B[1]), .B(A[546]), .Z(\ab[546][1] ) );
  AND U2027 ( .A(A[546]), .B(B[0]), .Z(\ab[546][0] ) );
  AND U2028 ( .A(B[3]), .B(A[545]), .Z(\ab[545][3] ) );
  AND U2029 ( .A(B[2]), .B(A[545]), .Z(\ab[545][2] ) );
  AND U2030 ( .A(B[1]), .B(A[545]), .Z(\ab[545][1] ) );
  AND U2031 ( .A(A[545]), .B(B[0]), .Z(\ab[545][0] ) );
  AND U2032 ( .A(B[3]), .B(A[544]), .Z(\ab[544][3] ) );
  AND U2033 ( .A(B[2]), .B(A[544]), .Z(\ab[544][2] ) );
  AND U2034 ( .A(B[1]), .B(A[544]), .Z(\ab[544][1] ) );
  AND U2035 ( .A(A[544]), .B(B[0]), .Z(\ab[544][0] ) );
  AND U2036 ( .A(B[3]), .B(A[543]), .Z(\ab[543][3] ) );
  AND U2037 ( .A(B[2]), .B(A[543]), .Z(\ab[543][2] ) );
  AND U2038 ( .A(B[1]), .B(A[543]), .Z(\ab[543][1] ) );
  AND U2039 ( .A(A[543]), .B(B[0]), .Z(\ab[543][0] ) );
  AND U2040 ( .A(B[3]), .B(A[542]), .Z(\ab[542][3] ) );
  AND U2041 ( .A(B[2]), .B(A[542]), .Z(\ab[542][2] ) );
  AND U2042 ( .A(B[1]), .B(A[542]), .Z(\ab[542][1] ) );
  AND U2043 ( .A(A[542]), .B(B[0]), .Z(\ab[542][0] ) );
  AND U2044 ( .A(B[3]), .B(A[541]), .Z(\ab[541][3] ) );
  AND U2045 ( .A(B[2]), .B(A[541]), .Z(\ab[541][2] ) );
  AND U2046 ( .A(B[1]), .B(A[541]), .Z(\ab[541][1] ) );
  AND U2047 ( .A(A[541]), .B(B[0]), .Z(\ab[541][0] ) );
  AND U2048 ( .A(B[3]), .B(A[540]), .Z(\ab[540][3] ) );
  AND U2049 ( .A(B[2]), .B(A[540]), .Z(\ab[540][2] ) );
  AND U2050 ( .A(B[1]), .B(A[540]), .Z(\ab[540][1] ) );
  AND U2051 ( .A(A[540]), .B(B[0]), .Z(\ab[540][0] ) );
  AND U2052 ( .A(B[3]), .B(A[53]), .Z(\ab[53][3] ) );
  AND U2053 ( .A(B[2]), .B(A[53]), .Z(\ab[53][2] ) );
  AND U2054 ( .A(B[1]), .B(A[53]), .Z(\ab[53][1] ) );
  AND U2055 ( .A(A[53]), .B(B[0]), .Z(\ab[53][0] ) );
  AND U2056 ( .A(B[3]), .B(A[539]), .Z(\ab[539][3] ) );
  AND U2057 ( .A(B[2]), .B(A[539]), .Z(\ab[539][2] ) );
  AND U2058 ( .A(B[1]), .B(A[539]), .Z(\ab[539][1] ) );
  AND U2059 ( .A(A[539]), .B(B[0]), .Z(\ab[539][0] ) );
  AND U2060 ( .A(B[3]), .B(A[538]), .Z(\ab[538][3] ) );
  AND U2061 ( .A(B[2]), .B(A[538]), .Z(\ab[538][2] ) );
  AND U2062 ( .A(B[1]), .B(A[538]), .Z(\ab[538][1] ) );
  AND U2063 ( .A(A[538]), .B(B[0]), .Z(\ab[538][0] ) );
  AND U2064 ( .A(B[3]), .B(A[537]), .Z(\ab[537][3] ) );
  AND U2065 ( .A(B[2]), .B(A[537]), .Z(\ab[537][2] ) );
  AND U2066 ( .A(B[1]), .B(A[537]), .Z(\ab[537][1] ) );
  AND U2067 ( .A(A[537]), .B(B[0]), .Z(\ab[537][0] ) );
  AND U2068 ( .A(B[3]), .B(A[536]), .Z(\ab[536][3] ) );
  AND U2069 ( .A(B[2]), .B(A[536]), .Z(\ab[536][2] ) );
  AND U2070 ( .A(B[1]), .B(A[536]), .Z(\ab[536][1] ) );
  AND U2071 ( .A(A[536]), .B(B[0]), .Z(\ab[536][0] ) );
  AND U2072 ( .A(B[3]), .B(A[535]), .Z(\ab[535][3] ) );
  AND U2073 ( .A(B[2]), .B(A[535]), .Z(\ab[535][2] ) );
  AND U2074 ( .A(B[1]), .B(A[535]), .Z(\ab[535][1] ) );
  AND U2075 ( .A(A[535]), .B(B[0]), .Z(\ab[535][0] ) );
  AND U2076 ( .A(B[3]), .B(A[534]), .Z(\ab[534][3] ) );
  AND U2077 ( .A(B[2]), .B(A[534]), .Z(\ab[534][2] ) );
  AND U2078 ( .A(B[1]), .B(A[534]), .Z(\ab[534][1] ) );
  AND U2079 ( .A(A[534]), .B(B[0]), .Z(\ab[534][0] ) );
  AND U2080 ( .A(B[3]), .B(A[533]), .Z(\ab[533][3] ) );
  AND U2081 ( .A(B[2]), .B(A[533]), .Z(\ab[533][2] ) );
  AND U2082 ( .A(B[1]), .B(A[533]), .Z(\ab[533][1] ) );
  AND U2083 ( .A(A[533]), .B(B[0]), .Z(\ab[533][0] ) );
  AND U2084 ( .A(B[3]), .B(A[532]), .Z(\ab[532][3] ) );
  AND U2085 ( .A(B[2]), .B(A[532]), .Z(\ab[532][2] ) );
  AND U2086 ( .A(B[1]), .B(A[532]), .Z(\ab[532][1] ) );
  AND U2087 ( .A(A[532]), .B(B[0]), .Z(\ab[532][0] ) );
  AND U2088 ( .A(B[3]), .B(A[531]), .Z(\ab[531][3] ) );
  AND U2089 ( .A(B[2]), .B(A[531]), .Z(\ab[531][2] ) );
  AND U2090 ( .A(B[1]), .B(A[531]), .Z(\ab[531][1] ) );
  AND U2091 ( .A(A[531]), .B(B[0]), .Z(\ab[531][0] ) );
  AND U2092 ( .A(B[3]), .B(A[530]), .Z(\ab[530][3] ) );
  AND U2093 ( .A(B[2]), .B(A[530]), .Z(\ab[530][2] ) );
  AND U2094 ( .A(B[1]), .B(A[530]), .Z(\ab[530][1] ) );
  AND U2095 ( .A(A[530]), .B(B[0]), .Z(\ab[530][0] ) );
  AND U2096 ( .A(B[3]), .B(A[52]), .Z(\ab[52][3] ) );
  AND U2097 ( .A(B[2]), .B(A[52]), .Z(\ab[52][2] ) );
  AND U2098 ( .A(B[1]), .B(A[52]), .Z(\ab[52][1] ) );
  AND U2099 ( .A(A[52]), .B(B[0]), .Z(\ab[52][0] ) );
  AND U2100 ( .A(B[3]), .B(A[529]), .Z(\ab[529][3] ) );
  AND U2101 ( .A(B[2]), .B(A[529]), .Z(\ab[529][2] ) );
  AND U2102 ( .A(B[1]), .B(A[529]), .Z(\ab[529][1] ) );
  AND U2103 ( .A(A[529]), .B(B[0]), .Z(\ab[529][0] ) );
  AND U2104 ( .A(B[3]), .B(A[528]), .Z(\ab[528][3] ) );
  AND U2105 ( .A(B[2]), .B(A[528]), .Z(\ab[528][2] ) );
  AND U2106 ( .A(B[1]), .B(A[528]), .Z(\ab[528][1] ) );
  AND U2107 ( .A(A[528]), .B(B[0]), .Z(\ab[528][0] ) );
  AND U2108 ( .A(B[3]), .B(A[527]), .Z(\ab[527][3] ) );
  AND U2109 ( .A(B[2]), .B(A[527]), .Z(\ab[527][2] ) );
  AND U2110 ( .A(B[1]), .B(A[527]), .Z(\ab[527][1] ) );
  AND U2111 ( .A(A[527]), .B(B[0]), .Z(\ab[527][0] ) );
  AND U2112 ( .A(B[3]), .B(A[526]), .Z(\ab[526][3] ) );
  AND U2113 ( .A(B[2]), .B(A[526]), .Z(\ab[526][2] ) );
  AND U2114 ( .A(B[1]), .B(A[526]), .Z(\ab[526][1] ) );
  AND U2115 ( .A(A[526]), .B(B[0]), .Z(\ab[526][0] ) );
  AND U2116 ( .A(B[3]), .B(A[525]), .Z(\ab[525][3] ) );
  AND U2117 ( .A(B[2]), .B(A[525]), .Z(\ab[525][2] ) );
  AND U2118 ( .A(B[1]), .B(A[525]), .Z(\ab[525][1] ) );
  AND U2119 ( .A(A[525]), .B(B[0]), .Z(\ab[525][0] ) );
  AND U2120 ( .A(B[3]), .B(A[524]), .Z(\ab[524][3] ) );
  AND U2121 ( .A(B[2]), .B(A[524]), .Z(\ab[524][2] ) );
  AND U2122 ( .A(B[1]), .B(A[524]), .Z(\ab[524][1] ) );
  AND U2123 ( .A(A[524]), .B(B[0]), .Z(\ab[524][0] ) );
  AND U2124 ( .A(B[3]), .B(A[523]), .Z(\ab[523][3] ) );
  AND U2125 ( .A(B[2]), .B(A[523]), .Z(\ab[523][2] ) );
  AND U2126 ( .A(B[1]), .B(A[523]), .Z(\ab[523][1] ) );
  AND U2127 ( .A(A[523]), .B(B[0]), .Z(\ab[523][0] ) );
  AND U2128 ( .A(B[3]), .B(A[522]), .Z(\ab[522][3] ) );
  AND U2129 ( .A(B[2]), .B(A[522]), .Z(\ab[522][2] ) );
  AND U2130 ( .A(B[1]), .B(A[522]), .Z(\ab[522][1] ) );
  AND U2131 ( .A(A[522]), .B(B[0]), .Z(\ab[522][0] ) );
  AND U2132 ( .A(B[3]), .B(A[521]), .Z(\ab[521][3] ) );
  AND U2133 ( .A(B[2]), .B(A[521]), .Z(\ab[521][2] ) );
  AND U2134 ( .A(B[1]), .B(A[521]), .Z(\ab[521][1] ) );
  AND U2135 ( .A(A[521]), .B(B[0]), .Z(\ab[521][0] ) );
  AND U2136 ( .A(B[3]), .B(A[520]), .Z(\ab[520][3] ) );
  AND U2137 ( .A(B[2]), .B(A[520]), .Z(\ab[520][2] ) );
  AND U2138 ( .A(B[1]), .B(A[520]), .Z(\ab[520][1] ) );
  AND U2139 ( .A(A[520]), .B(B[0]), .Z(\ab[520][0] ) );
  AND U2140 ( .A(B[3]), .B(A[51]), .Z(\ab[51][3] ) );
  AND U2141 ( .A(B[2]), .B(A[51]), .Z(\ab[51][2] ) );
  AND U2142 ( .A(B[1]), .B(A[51]), .Z(\ab[51][1] ) );
  AND U2143 ( .A(A[51]), .B(B[0]), .Z(\ab[51][0] ) );
  AND U2144 ( .A(B[3]), .B(A[519]), .Z(\ab[519][3] ) );
  AND U2145 ( .A(B[2]), .B(A[519]), .Z(\ab[519][2] ) );
  AND U2146 ( .A(B[1]), .B(A[519]), .Z(\ab[519][1] ) );
  AND U2147 ( .A(A[519]), .B(B[0]), .Z(\ab[519][0] ) );
  AND U2148 ( .A(B[3]), .B(A[518]), .Z(\ab[518][3] ) );
  AND U2149 ( .A(B[2]), .B(A[518]), .Z(\ab[518][2] ) );
  AND U2150 ( .A(B[1]), .B(A[518]), .Z(\ab[518][1] ) );
  AND U2151 ( .A(A[518]), .B(B[0]), .Z(\ab[518][0] ) );
  AND U2152 ( .A(B[3]), .B(A[517]), .Z(\ab[517][3] ) );
  AND U2153 ( .A(B[2]), .B(A[517]), .Z(\ab[517][2] ) );
  AND U2154 ( .A(B[1]), .B(A[517]), .Z(\ab[517][1] ) );
  AND U2155 ( .A(A[517]), .B(B[0]), .Z(\ab[517][0] ) );
  AND U2156 ( .A(B[3]), .B(A[516]), .Z(\ab[516][3] ) );
  AND U2157 ( .A(B[2]), .B(A[516]), .Z(\ab[516][2] ) );
  AND U2158 ( .A(B[1]), .B(A[516]), .Z(\ab[516][1] ) );
  AND U2159 ( .A(A[516]), .B(B[0]), .Z(\ab[516][0] ) );
  AND U2160 ( .A(B[3]), .B(A[515]), .Z(\ab[515][3] ) );
  AND U2161 ( .A(B[2]), .B(A[515]), .Z(\ab[515][2] ) );
  AND U2162 ( .A(B[1]), .B(A[515]), .Z(\ab[515][1] ) );
  AND U2163 ( .A(A[515]), .B(B[0]), .Z(\ab[515][0] ) );
  AND U2164 ( .A(B[3]), .B(A[514]), .Z(\ab[514][3] ) );
  AND U2165 ( .A(B[2]), .B(A[514]), .Z(\ab[514][2] ) );
  AND U2166 ( .A(B[1]), .B(A[514]), .Z(\ab[514][1] ) );
  AND U2167 ( .A(A[514]), .B(B[0]), .Z(\ab[514][0] ) );
  AND U2168 ( .A(B[3]), .B(A[513]), .Z(\ab[513][3] ) );
  AND U2169 ( .A(B[2]), .B(A[513]), .Z(\ab[513][2] ) );
  AND U2170 ( .A(B[1]), .B(A[513]), .Z(\ab[513][1] ) );
  AND U2171 ( .A(A[513]), .B(B[0]), .Z(\ab[513][0] ) );
  AND U2172 ( .A(B[3]), .B(A[512]), .Z(\ab[512][3] ) );
  AND U2173 ( .A(B[2]), .B(A[512]), .Z(\ab[512][2] ) );
  AND U2174 ( .A(B[1]), .B(A[512]), .Z(\ab[512][1] ) );
  AND U2175 ( .A(A[512]), .B(B[0]), .Z(\ab[512][0] ) );
  AND U2176 ( .A(B[3]), .B(A[511]), .Z(\ab[511][3] ) );
  AND U2177 ( .A(B[2]), .B(A[511]), .Z(\ab[511][2] ) );
  AND U2178 ( .A(B[1]), .B(A[511]), .Z(\ab[511][1] ) );
  AND U2179 ( .A(A[511]), .B(B[0]), .Z(\ab[511][0] ) );
  AND U2180 ( .A(B[3]), .B(A[510]), .Z(\ab[510][3] ) );
  AND U2181 ( .A(B[2]), .B(A[510]), .Z(\ab[510][2] ) );
  AND U2182 ( .A(B[1]), .B(A[510]), .Z(\ab[510][1] ) );
  AND U2183 ( .A(A[510]), .B(B[0]), .Z(\ab[510][0] ) );
  AND U2184 ( .A(B[3]), .B(A[50]), .Z(\ab[50][3] ) );
  AND U2185 ( .A(B[2]), .B(A[50]), .Z(\ab[50][2] ) );
  AND U2186 ( .A(B[1]), .B(A[50]), .Z(\ab[50][1] ) );
  AND U2187 ( .A(A[50]), .B(B[0]), .Z(\ab[50][0] ) );
  AND U2188 ( .A(B[3]), .B(A[509]), .Z(\ab[509][3] ) );
  AND U2189 ( .A(B[2]), .B(A[509]), .Z(\ab[509][2] ) );
  AND U2190 ( .A(B[1]), .B(A[509]), .Z(\ab[509][1] ) );
  AND U2191 ( .A(A[509]), .B(B[0]), .Z(\ab[509][0] ) );
  AND U2192 ( .A(B[3]), .B(A[508]), .Z(\ab[508][3] ) );
  AND U2193 ( .A(B[2]), .B(A[508]), .Z(\ab[508][2] ) );
  AND U2194 ( .A(B[1]), .B(A[508]), .Z(\ab[508][1] ) );
  AND U2195 ( .A(A[508]), .B(B[0]), .Z(\ab[508][0] ) );
  AND U2196 ( .A(B[3]), .B(A[507]), .Z(\ab[507][3] ) );
  AND U2197 ( .A(B[2]), .B(A[507]), .Z(\ab[507][2] ) );
  AND U2198 ( .A(B[1]), .B(A[507]), .Z(\ab[507][1] ) );
  AND U2199 ( .A(A[507]), .B(B[0]), .Z(\ab[507][0] ) );
  AND U2200 ( .A(B[3]), .B(A[506]), .Z(\ab[506][3] ) );
  AND U2201 ( .A(B[2]), .B(A[506]), .Z(\ab[506][2] ) );
  AND U2202 ( .A(B[1]), .B(A[506]), .Z(\ab[506][1] ) );
  AND U2203 ( .A(A[506]), .B(B[0]), .Z(\ab[506][0] ) );
  AND U2204 ( .A(B[3]), .B(A[505]), .Z(\ab[505][3] ) );
  AND U2205 ( .A(B[2]), .B(A[505]), .Z(\ab[505][2] ) );
  AND U2206 ( .A(B[1]), .B(A[505]), .Z(\ab[505][1] ) );
  AND U2207 ( .A(A[505]), .B(B[0]), .Z(\ab[505][0] ) );
  AND U2208 ( .A(B[3]), .B(A[504]), .Z(\ab[504][3] ) );
  AND U2209 ( .A(B[2]), .B(A[504]), .Z(\ab[504][2] ) );
  AND U2210 ( .A(B[1]), .B(A[504]), .Z(\ab[504][1] ) );
  AND U2211 ( .A(A[504]), .B(B[0]), .Z(\ab[504][0] ) );
  AND U2212 ( .A(B[3]), .B(A[503]), .Z(\ab[503][3] ) );
  AND U2213 ( .A(B[2]), .B(A[503]), .Z(\ab[503][2] ) );
  AND U2214 ( .A(B[1]), .B(A[503]), .Z(\ab[503][1] ) );
  AND U2215 ( .A(A[503]), .B(B[0]), .Z(\ab[503][0] ) );
  AND U2216 ( .A(B[3]), .B(A[502]), .Z(\ab[502][3] ) );
  AND U2217 ( .A(B[2]), .B(A[502]), .Z(\ab[502][2] ) );
  AND U2218 ( .A(B[1]), .B(A[502]), .Z(\ab[502][1] ) );
  AND U2219 ( .A(A[502]), .B(B[0]), .Z(\ab[502][0] ) );
  AND U2220 ( .A(B[3]), .B(A[501]), .Z(\ab[501][3] ) );
  AND U2221 ( .A(B[2]), .B(A[501]), .Z(\ab[501][2] ) );
  AND U2222 ( .A(B[1]), .B(A[501]), .Z(\ab[501][1] ) );
  AND U2223 ( .A(A[501]), .B(B[0]), .Z(\ab[501][0] ) );
  AND U2224 ( .A(B[3]), .B(A[500]), .Z(\ab[500][3] ) );
  AND U2225 ( .A(B[2]), .B(A[500]), .Z(\ab[500][2] ) );
  AND U2226 ( .A(B[1]), .B(A[500]), .Z(\ab[500][1] ) );
  AND U2227 ( .A(A[500]), .B(B[0]), .Z(\ab[500][0] ) );
  AND U2228 ( .A(B[3]), .B(A[4]), .Z(\ab[4][3] ) );
  AND U2229 ( .A(B[2]), .B(A[4]), .Z(\ab[4][2] ) );
  AND U2230 ( .A(B[1]), .B(A[4]), .Z(\ab[4][1] ) );
  AND U2231 ( .A(A[4]), .B(B[0]), .Z(\ab[4][0] ) );
  AND U2232 ( .A(B[3]), .B(A[49]), .Z(\ab[49][3] ) );
  AND U2233 ( .A(B[2]), .B(A[49]), .Z(\ab[49][2] ) );
  AND U2234 ( .A(B[1]), .B(A[49]), .Z(\ab[49][1] ) );
  AND U2235 ( .A(A[49]), .B(B[0]), .Z(\ab[49][0] ) );
  AND U2236 ( .A(B[3]), .B(A[499]), .Z(\ab[499][3] ) );
  AND U2237 ( .A(B[2]), .B(A[499]), .Z(\ab[499][2] ) );
  AND U2238 ( .A(B[1]), .B(A[499]), .Z(\ab[499][1] ) );
  AND U2239 ( .A(A[499]), .B(B[0]), .Z(\ab[499][0] ) );
  AND U2240 ( .A(B[3]), .B(A[498]), .Z(\ab[498][3] ) );
  AND U2241 ( .A(B[2]), .B(A[498]), .Z(\ab[498][2] ) );
  AND U2242 ( .A(B[1]), .B(A[498]), .Z(\ab[498][1] ) );
  AND U2243 ( .A(A[498]), .B(B[0]), .Z(\ab[498][0] ) );
  AND U2244 ( .A(B[3]), .B(A[497]), .Z(\ab[497][3] ) );
  AND U2245 ( .A(B[2]), .B(A[497]), .Z(\ab[497][2] ) );
  AND U2246 ( .A(B[1]), .B(A[497]), .Z(\ab[497][1] ) );
  AND U2247 ( .A(A[497]), .B(B[0]), .Z(\ab[497][0] ) );
  AND U2248 ( .A(B[3]), .B(A[496]), .Z(\ab[496][3] ) );
  AND U2249 ( .A(B[2]), .B(A[496]), .Z(\ab[496][2] ) );
  AND U2250 ( .A(B[1]), .B(A[496]), .Z(\ab[496][1] ) );
  AND U2251 ( .A(A[496]), .B(B[0]), .Z(\ab[496][0] ) );
  AND U2252 ( .A(B[3]), .B(A[495]), .Z(\ab[495][3] ) );
  AND U2253 ( .A(B[2]), .B(A[495]), .Z(\ab[495][2] ) );
  AND U2254 ( .A(B[1]), .B(A[495]), .Z(\ab[495][1] ) );
  AND U2255 ( .A(A[495]), .B(B[0]), .Z(\ab[495][0] ) );
  AND U2256 ( .A(B[3]), .B(A[494]), .Z(\ab[494][3] ) );
  AND U2257 ( .A(B[2]), .B(A[494]), .Z(\ab[494][2] ) );
  AND U2258 ( .A(B[1]), .B(A[494]), .Z(\ab[494][1] ) );
  AND U2259 ( .A(A[494]), .B(B[0]), .Z(\ab[494][0] ) );
  AND U2260 ( .A(B[3]), .B(A[493]), .Z(\ab[493][3] ) );
  AND U2261 ( .A(B[2]), .B(A[493]), .Z(\ab[493][2] ) );
  AND U2262 ( .A(B[1]), .B(A[493]), .Z(\ab[493][1] ) );
  AND U2263 ( .A(A[493]), .B(B[0]), .Z(\ab[493][0] ) );
  AND U2264 ( .A(B[3]), .B(A[492]), .Z(\ab[492][3] ) );
  AND U2265 ( .A(B[2]), .B(A[492]), .Z(\ab[492][2] ) );
  AND U2266 ( .A(B[1]), .B(A[492]), .Z(\ab[492][1] ) );
  AND U2267 ( .A(A[492]), .B(B[0]), .Z(\ab[492][0] ) );
  AND U2268 ( .A(B[3]), .B(A[491]), .Z(\ab[491][3] ) );
  AND U2269 ( .A(B[2]), .B(A[491]), .Z(\ab[491][2] ) );
  AND U2270 ( .A(B[1]), .B(A[491]), .Z(\ab[491][1] ) );
  AND U2271 ( .A(A[491]), .B(B[0]), .Z(\ab[491][0] ) );
  AND U2272 ( .A(B[3]), .B(A[490]), .Z(\ab[490][3] ) );
  AND U2273 ( .A(B[2]), .B(A[490]), .Z(\ab[490][2] ) );
  AND U2274 ( .A(B[1]), .B(A[490]), .Z(\ab[490][1] ) );
  AND U2275 ( .A(A[490]), .B(B[0]), .Z(\ab[490][0] ) );
  AND U2276 ( .A(B[3]), .B(A[48]), .Z(\ab[48][3] ) );
  AND U2277 ( .A(B[2]), .B(A[48]), .Z(\ab[48][2] ) );
  AND U2278 ( .A(B[1]), .B(A[48]), .Z(\ab[48][1] ) );
  AND U2279 ( .A(A[48]), .B(B[0]), .Z(\ab[48][0] ) );
  AND U2280 ( .A(B[3]), .B(A[489]), .Z(\ab[489][3] ) );
  AND U2281 ( .A(B[2]), .B(A[489]), .Z(\ab[489][2] ) );
  AND U2282 ( .A(B[1]), .B(A[489]), .Z(\ab[489][1] ) );
  AND U2283 ( .A(A[489]), .B(B[0]), .Z(\ab[489][0] ) );
  AND U2284 ( .A(B[3]), .B(A[488]), .Z(\ab[488][3] ) );
  AND U2285 ( .A(B[2]), .B(A[488]), .Z(\ab[488][2] ) );
  AND U2286 ( .A(B[1]), .B(A[488]), .Z(\ab[488][1] ) );
  AND U2287 ( .A(A[488]), .B(B[0]), .Z(\ab[488][0] ) );
  AND U2288 ( .A(B[3]), .B(A[487]), .Z(\ab[487][3] ) );
  AND U2289 ( .A(B[2]), .B(A[487]), .Z(\ab[487][2] ) );
  AND U2290 ( .A(B[1]), .B(A[487]), .Z(\ab[487][1] ) );
  AND U2291 ( .A(A[487]), .B(B[0]), .Z(\ab[487][0] ) );
  AND U2292 ( .A(B[3]), .B(A[486]), .Z(\ab[486][3] ) );
  AND U2293 ( .A(B[2]), .B(A[486]), .Z(\ab[486][2] ) );
  AND U2294 ( .A(B[1]), .B(A[486]), .Z(\ab[486][1] ) );
  AND U2295 ( .A(A[486]), .B(B[0]), .Z(\ab[486][0] ) );
  AND U2296 ( .A(B[3]), .B(A[485]), .Z(\ab[485][3] ) );
  AND U2297 ( .A(B[2]), .B(A[485]), .Z(\ab[485][2] ) );
  AND U2298 ( .A(B[1]), .B(A[485]), .Z(\ab[485][1] ) );
  AND U2299 ( .A(A[485]), .B(B[0]), .Z(\ab[485][0] ) );
  AND U2300 ( .A(B[3]), .B(A[484]), .Z(\ab[484][3] ) );
  AND U2301 ( .A(B[2]), .B(A[484]), .Z(\ab[484][2] ) );
  AND U2302 ( .A(B[1]), .B(A[484]), .Z(\ab[484][1] ) );
  AND U2303 ( .A(A[484]), .B(B[0]), .Z(\ab[484][0] ) );
  AND U2304 ( .A(B[3]), .B(A[483]), .Z(\ab[483][3] ) );
  AND U2305 ( .A(B[2]), .B(A[483]), .Z(\ab[483][2] ) );
  AND U2306 ( .A(B[1]), .B(A[483]), .Z(\ab[483][1] ) );
  AND U2307 ( .A(A[483]), .B(B[0]), .Z(\ab[483][0] ) );
  AND U2308 ( .A(B[3]), .B(A[482]), .Z(\ab[482][3] ) );
  AND U2309 ( .A(B[2]), .B(A[482]), .Z(\ab[482][2] ) );
  AND U2310 ( .A(B[1]), .B(A[482]), .Z(\ab[482][1] ) );
  AND U2311 ( .A(A[482]), .B(B[0]), .Z(\ab[482][0] ) );
  AND U2312 ( .A(B[3]), .B(A[481]), .Z(\ab[481][3] ) );
  AND U2313 ( .A(B[2]), .B(A[481]), .Z(\ab[481][2] ) );
  AND U2314 ( .A(B[1]), .B(A[481]), .Z(\ab[481][1] ) );
  AND U2315 ( .A(A[481]), .B(B[0]), .Z(\ab[481][0] ) );
  AND U2316 ( .A(B[3]), .B(A[480]), .Z(\ab[480][3] ) );
  AND U2317 ( .A(B[2]), .B(A[480]), .Z(\ab[480][2] ) );
  AND U2318 ( .A(B[1]), .B(A[480]), .Z(\ab[480][1] ) );
  AND U2319 ( .A(A[480]), .B(B[0]), .Z(\ab[480][0] ) );
  AND U2320 ( .A(B[3]), .B(A[47]), .Z(\ab[47][3] ) );
  AND U2321 ( .A(B[2]), .B(A[47]), .Z(\ab[47][2] ) );
  AND U2322 ( .A(B[1]), .B(A[47]), .Z(\ab[47][1] ) );
  AND U2323 ( .A(A[47]), .B(B[0]), .Z(\ab[47][0] ) );
  AND U2324 ( .A(B[3]), .B(A[479]), .Z(\ab[479][3] ) );
  AND U2325 ( .A(B[2]), .B(A[479]), .Z(\ab[479][2] ) );
  AND U2326 ( .A(B[1]), .B(A[479]), .Z(\ab[479][1] ) );
  AND U2327 ( .A(A[479]), .B(B[0]), .Z(\ab[479][0] ) );
  AND U2328 ( .A(B[3]), .B(A[478]), .Z(\ab[478][3] ) );
  AND U2329 ( .A(B[2]), .B(A[478]), .Z(\ab[478][2] ) );
  AND U2330 ( .A(B[1]), .B(A[478]), .Z(\ab[478][1] ) );
  AND U2331 ( .A(A[478]), .B(B[0]), .Z(\ab[478][0] ) );
  AND U2332 ( .A(B[3]), .B(A[477]), .Z(\ab[477][3] ) );
  AND U2333 ( .A(B[2]), .B(A[477]), .Z(\ab[477][2] ) );
  AND U2334 ( .A(B[1]), .B(A[477]), .Z(\ab[477][1] ) );
  AND U2335 ( .A(A[477]), .B(B[0]), .Z(\ab[477][0] ) );
  AND U2336 ( .A(B[3]), .B(A[476]), .Z(\ab[476][3] ) );
  AND U2337 ( .A(B[2]), .B(A[476]), .Z(\ab[476][2] ) );
  AND U2338 ( .A(B[1]), .B(A[476]), .Z(\ab[476][1] ) );
  AND U2339 ( .A(A[476]), .B(B[0]), .Z(\ab[476][0] ) );
  AND U2340 ( .A(B[3]), .B(A[475]), .Z(\ab[475][3] ) );
  AND U2341 ( .A(B[2]), .B(A[475]), .Z(\ab[475][2] ) );
  AND U2342 ( .A(B[1]), .B(A[475]), .Z(\ab[475][1] ) );
  AND U2343 ( .A(A[475]), .B(B[0]), .Z(\ab[475][0] ) );
  AND U2344 ( .A(B[3]), .B(A[474]), .Z(\ab[474][3] ) );
  AND U2345 ( .A(B[2]), .B(A[474]), .Z(\ab[474][2] ) );
  AND U2346 ( .A(B[1]), .B(A[474]), .Z(\ab[474][1] ) );
  AND U2347 ( .A(A[474]), .B(B[0]), .Z(\ab[474][0] ) );
  AND U2348 ( .A(B[3]), .B(A[473]), .Z(\ab[473][3] ) );
  AND U2349 ( .A(B[2]), .B(A[473]), .Z(\ab[473][2] ) );
  AND U2350 ( .A(B[1]), .B(A[473]), .Z(\ab[473][1] ) );
  AND U2351 ( .A(A[473]), .B(B[0]), .Z(\ab[473][0] ) );
  AND U2352 ( .A(B[3]), .B(A[472]), .Z(\ab[472][3] ) );
  AND U2353 ( .A(B[2]), .B(A[472]), .Z(\ab[472][2] ) );
  AND U2354 ( .A(B[1]), .B(A[472]), .Z(\ab[472][1] ) );
  AND U2355 ( .A(A[472]), .B(B[0]), .Z(\ab[472][0] ) );
  AND U2356 ( .A(B[3]), .B(A[471]), .Z(\ab[471][3] ) );
  AND U2357 ( .A(B[2]), .B(A[471]), .Z(\ab[471][2] ) );
  AND U2358 ( .A(B[1]), .B(A[471]), .Z(\ab[471][1] ) );
  AND U2359 ( .A(A[471]), .B(B[0]), .Z(\ab[471][0] ) );
  AND U2360 ( .A(B[3]), .B(A[470]), .Z(\ab[470][3] ) );
  AND U2361 ( .A(B[2]), .B(A[470]), .Z(\ab[470][2] ) );
  AND U2362 ( .A(B[1]), .B(A[470]), .Z(\ab[470][1] ) );
  AND U2363 ( .A(A[470]), .B(B[0]), .Z(\ab[470][0] ) );
  AND U2364 ( .A(B[3]), .B(A[46]), .Z(\ab[46][3] ) );
  AND U2365 ( .A(B[2]), .B(A[46]), .Z(\ab[46][2] ) );
  AND U2366 ( .A(B[1]), .B(A[46]), .Z(\ab[46][1] ) );
  AND U2367 ( .A(A[46]), .B(B[0]), .Z(\ab[46][0] ) );
  AND U2368 ( .A(B[3]), .B(A[469]), .Z(\ab[469][3] ) );
  AND U2369 ( .A(B[2]), .B(A[469]), .Z(\ab[469][2] ) );
  AND U2370 ( .A(B[1]), .B(A[469]), .Z(\ab[469][1] ) );
  AND U2371 ( .A(A[469]), .B(B[0]), .Z(\ab[469][0] ) );
  AND U2372 ( .A(B[3]), .B(A[468]), .Z(\ab[468][3] ) );
  AND U2373 ( .A(B[2]), .B(A[468]), .Z(\ab[468][2] ) );
  AND U2374 ( .A(B[1]), .B(A[468]), .Z(\ab[468][1] ) );
  AND U2375 ( .A(A[468]), .B(B[0]), .Z(\ab[468][0] ) );
  AND U2376 ( .A(B[3]), .B(A[467]), .Z(\ab[467][3] ) );
  AND U2377 ( .A(B[2]), .B(A[467]), .Z(\ab[467][2] ) );
  AND U2378 ( .A(B[1]), .B(A[467]), .Z(\ab[467][1] ) );
  AND U2379 ( .A(A[467]), .B(B[0]), .Z(\ab[467][0] ) );
  AND U2380 ( .A(B[3]), .B(A[466]), .Z(\ab[466][3] ) );
  AND U2381 ( .A(B[2]), .B(A[466]), .Z(\ab[466][2] ) );
  AND U2382 ( .A(B[1]), .B(A[466]), .Z(\ab[466][1] ) );
  AND U2383 ( .A(A[466]), .B(B[0]), .Z(\ab[466][0] ) );
  AND U2384 ( .A(B[3]), .B(A[465]), .Z(\ab[465][3] ) );
  AND U2385 ( .A(B[2]), .B(A[465]), .Z(\ab[465][2] ) );
  AND U2386 ( .A(B[1]), .B(A[465]), .Z(\ab[465][1] ) );
  AND U2387 ( .A(A[465]), .B(B[0]), .Z(\ab[465][0] ) );
  AND U2388 ( .A(B[3]), .B(A[464]), .Z(\ab[464][3] ) );
  AND U2389 ( .A(B[2]), .B(A[464]), .Z(\ab[464][2] ) );
  AND U2390 ( .A(B[1]), .B(A[464]), .Z(\ab[464][1] ) );
  AND U2391 ( .A(A[464]), .B(B[0]), .Z(\ab[464][0] ) );
  AND U2392 ( .A(B[3]), .B(A[463]), .Z(\ab[463][3] ) );
  AND U2393 ( .A(B[2]), .B(A[463]), .Z(\ab[463][2] ) );
  AND U2394 ( .A(B[1]), .B(A[463]), .Z(\ab[463][1] ) );
  AND U2395 ( .A(A[463]), .B(B[0]), .Z(\ab[463][0] ) );
  AND U2396 ( .A(B[3]), .B(A[462]), .Z(\ab[462][3] ) );
  AND U2397 ( .A(B[2]), .B(A[462]), .Z(\ab[462][2] ) );
  AND U2398 ( .A(B[1]), .B(A[462]), .Z(\ab[462][1] ) );
  AND U2399 ( .A(A[462]), .B(B[0]), .Z(\ab[462][0] ) );
  AND U2400 ( .A(B[3]), .B(A[461]), .Z(\ab[461][3] ) );
  AND U2401 ( .A(B[2]), .B(A[461]), .Z(\ab[461][2] ) );
  AND U2402 ( .A(B[1]), .B(A[461]), .Z(\ab[461][1] ) );
  AND U2403 ( .A(A[461]), .B(B[0]), .Z(\ab[461][0] ) );
  AND U2404 ( .A(B[3]), .B(A[460]), .Z(\ab[460][3] ) );
  AND U2405 ( .A(B[2]), .B(A[460]), .Z(\ab[460][2] ) );
  AND U2406 ( .A(B[1]), .B(A[460]), .Z(\ab[460][1] ) );
  AND U2407 ( .A(A[460]), .B(B[0]), .Z(\ab[460][0] ) );
  AND U2408 ( .A(B[3]), .B(A[45]), .Z(\ab[45][3] ) );
  AND U2409 ( .A(B[2]), .B(A[45]), .Z(\ab[45][2] ) );
  AND U2410 ( .A(B[1]), .B(A[45]), .Z(\ab[45][1] ) );
  AND U2411 ( .A(A[45]), .B(B[0]), .Z(\ab[45][0] ) );
  AND U2412 ( .A(B[3]), .B(A[459]), .Z(\ab[459][3] ) );
  AND U2413 ( .A(B[2]), .B(A[459]), .Z(\ab[459][2] ) );
  AND U2414 ( .A(B[1]), .B(A[459]), .Z(\ab[459][1] ) );
  AND U2415 ( .A(A[459]), .B(B[0]), .Z(\ab[459][0] ) );
  AND U2416 ( .A(B[3]), .B(A[458]), .Z(\ab[458][3] ) );
  AND U2417 ( .A(B[2]), .B(A[458]), .Z(\ab[458][2] ) );
  AND U2418 ( .A(B[1]), .B(A[458]), .Z(\ab[458][1] ) );
  AND U2419 ( .A(A[458]), .B(B[0]), .Z(\ab[458][0] ) );
  AND U2420 ( .A(B[3]), .B(A[457]), .Z(\ab[457][3] ) );
  AND U2421 ( .A(B[2]), .B(A[457]), .Z(\ab[457][2] ) );
  AND U2422 ( .A(B[1]), .B(A[457]), .Z(\ab[457][1] ) );
  AND U2423 ( .A(A[457]), .B(B[0]), .Z(\ab[457][0] ) );
  AND U2424 ( .A(B[3]), .B(A[456]), .Z(\ab[456][3] ) );
  AND U2425 ( .A(B[2]), .B(A[456]), .Z(\ab[456][2] ) );
  AND U2426 ( .A(B[1]), .B(A[456]), .Z(\ab[456][1] ) );
  AND U2427 ( .A(A[456]), .B(B[0]), .Z(\ab[456][0] ) );
  AND U2428 ( .A(B[3]), .B(A[455]), .Z(\ab[455][3] ) );
  AND U2429 ( .A(B[2]), .B(A[455]), .Z(\ab[455][2] ) );
  AND U2430 ( .A(B[1]), .B(A[455]), .Z(\ab[455][1] ) );
  AND U2431 ( .A(A[455]), .B(B[0]), .Z(\ab[455][0] ) );
  AND U2432 ( .A(B[3]), .B(A[454]), .Z(\ab[454][3] ) );
  AND U2433 ( .A(B[2]), .B(A[454]), .Z(\ab[454][2] ) );
  AND U2434 ( .A(B[1]), .B(A[454]), .Z(\ab[454][1] ) );
  AND U2435 ( .A(A[454]), .B(B[0]), .Z(\ab[454][0] ) );
  AND U2436 ( .A(B[3]), .B(A[453]), .Z(\ab[453][3] ) );
  AND U2437 ( .A(B[2]), .B(A[453]), .Z(\ab[453][2] ) );
  AND U2438 ( .A(B[1]), .B(A[453]), .Z(\ab[453][1] ) );
  AND U2439 ( .A(A[453]), .B(B[0]), .Z(\ab[453][0] ) );
  AND U2440 ( .A(B[3]), .B(A[452]), .Z(\ab[452][3] ) );
  AND U2441 ( .A(B[2]), .B(A[452]), .Z(\ab[452][2] ) );
  AND U2442 ( .A(B[1]), .B(A[452]), .Z(\ab[452][1] ) );
  AND U2443 ( .A(A[452]), .B(B[0]), .Z(\ab[452][0] ) );
  AND U2444 ( .A(B[3]), .B(A[451]), .Z(\ab[451][3] ) );
  AND U2445 ( .A(B[2]), .B(A[451]), .Z(\ab[451][2] ) );
  AND U2446 ( .A(B[1]), .B(A[451]), .Z(\ab[451][1] ) );
  AND U2447 ( .A(A[451]), .B(B[0]), .Z(\ab[451][0] ) );
  AND U2448 ( .A(B[3]), .B(A[450]), .Z(\ab[450][3] ) );
  AND U2449 ( .A(B[2]), .B(A[450]), .Z(\ab[450][2] ) );
  AND U2450 ( .A(B[1]), .B(A[450]), .Z(\ab[450][1] ) );
  AND U2451 ( .A(A[450]), .B(B[0]), .Z(\ab[450][0] ) );
  AND U2452 ( .A(B[3]), .B(A[44]), .Z(\ab[44][3] ) );
  AND U2453 ( .A(B[2]), .B(A[44]), .Z(\ab[44][2] ) );
  AND U2454 ( .A(B[1]), .B(A[44]), .Z(\ab[44][1] ) );
  AND U2455 ( .A(A[44]), .B(B[0]), .Z(\ab[44][0] ) );
  AND U2456 ( .A(B[3]), .B(A[449]), .Z(\ab[449][3] ) );
  AND U2457 ( .A(B[2]), .B(A[449]), .Z(\ab[449][2] ) );
  AND U2458 ( .A(B[1]), .B(A[449]), .Z(\ab[449][1] ) );
  AND U2459 ( .A(A[449]), .B(B[0]), .Z(\ab[449][0] ) );
  AND U2460 ( .A(B[3]), .B(A[448]), .Z(\ab[448][3] ) );
  AND U2461 ( .A(B[2]), .B(A[448]), .Z(\ab[448][2] ) );
  AND U2462 ( .A(B[1]), .B(A[448]), .Z(\ab[448][1] ) );
  AND U2463 ( .A(A[448]), .B(B[0]), .Z(\ab[448][0] ) );
  AND U2464 ( .A(B[3]), .B(A[447]), .Z(\ab[447][3] ) );
  AND U2465 ( .A(B[2]), .B(A[447]), .Z(\ab[447][2] ) );
  AND U2466 ( .A(B[1]), .B(A[447]), .Z(\ab[447][1] ) );
  AND U2467 ( .A(A[447]), .B(B[0]), .Z(\ab[447][0] ) );
  AND U2468 ( .A(B[3]), .B(A[446]), .Z(\ab[446][3] ) );
  AND U2469 ( .A(B[2]), .B(A[446]), .Z(\ab[446][2] ) );
  AND U2470 ( .A(B[1]), .B(A[446]), .Z(\ab[446][1] ) );
  AND U2471 ( .A(A[446]), .B(B[0]), .Z(\ab[446][0] ) );
  AND U2472 ( .A(B[3]), .B(A[445]), .Z(\ab[445][3] ) );
  AND U2473 ( .A(B[2]), .B(A[445]), .Z(\ab[445][2] ) );
  AND U2474 ( .A(B[1]), .B(A[445]), .Z(\ab[445][1] ) );
  AND U2475 ( .A(A[445]), .B(B[0]), .Z(\ab[445][0] ) );
  AND U2476 ( .A(B[3]), .B(A[444]), .Z(\ab[444][3] ) );
  AND U2477 ( .A(B[2]), .B(A[444]), .Z(\ab[444][2] ) );
  AND U2478 ( .A(B[1]), .B(A[444]), .Z(\ab[444][1] ) );
  AND U2479 ( .A(A[444]), .B(B[0]), .Z(\ab[444][0] ) );
  AND U2480 ( .A(B[3]), .B(A[443]), .Z(\ab[443][3] ) );
  AND U2481 ( .A(B[2]), .B(A[443]), .Z(\ab[443][2] ) );
  AND U2482 ( .A(B[1]), .B(A[443]), .Z(\ab[443][1] ) );
  AND U2483 ( .A(A[443]), .B(B[0]), .Z(\ab[443][0] ) );
  AND U2484 ( .A(B[3]), .B(A[442]), .Z(\ab[442][3] ) );
  AND U2485 ( .A(B[2]), .B(A[442]), .Z(\ab[442][2] ) );
  AND U2486 ( .A(B[1]), .B(A[442]), .Z(\ab[442][1] ) );
  AND U2487 ( .A(A[442]), .B(B[0]), .Z(\ab[442][0] ) );
  AND U2488 ( .A(B[3]), .B(A[441]), .Z(\ab[441][3] ) );
  AND U2489 ( .A(B[2]), .B(A[441]), .Z(\ab[441][2] ) );
  AND U2490 ( .A(B[1]), .B(A[441]), .Z(\ab[441][1] ) );
  AND U2491 ( .A(A[441]), .B(B[0]), .Z(\ab[441][0] ) );
  AND U2492 ( .A(B[3]), .B(A[440]), .Z(\ab[440][3] ) );
  AND U2493 ( .A(B[2]), .B(A[440]), .Z(\ab[440][2] ) );
  AND U2494 ( .A(B[1]), .B(A[440]), .Z(\ab[440][1] ) );
  AND U2495 ( .A(A[440]), .B(B[0]), .Z(\ab[440][0] ) );
  AND U2496 ( .A(B[3]), .B(A[43]), .Z(\ab[43][3] ) );
  AND U2497 ( .A(B[2]), .B(A[43]), .Z(\ab[43][2] ) );
  AND U2498 ( .A(B[1]), .B(A[43]), .Z(\ab[43][1] ) );
  AND U2499 ( .A(A[43]), .B(B[0]), .Z(\ab[43][0] ) );
  AND U2500 ( .A(B[3]), .B(A[439]), .Z(\ab[439][3] ) );
  AND U2501 ( .A(B[2]), .B(A[439]), .Z(\ab[439][2] ) );
  AND U2502 ( .A(B[1]), .B(A[439]), .Z(\ab[439][1] ) );
  AND U2503 ( .A(A[439]), .B(B[0]), .Z(\ab[439][0] ) );
  AND U2504 ( .A(B[3]), .B(A[438]), .Z(\ab[438][3] ) );
  AND U2505 ( .A(B[2]), .B(A[438]), .Z(\ab[438][2] ) );
  AND U2506 ( .A(B[1]), .B(A[438]), .Z(\ab[438][1] ) );
  AND U2507 ( .A(A[438]), .B(B[0]), .Z(\ab[438][0] ) );
  AND U2508 ( .A(B[3]), .B(A[437]), .Z(\ab[437][3] ) );
  AND U2509 ( .A(B[2]), .B(A[437]), .Z(\ab[437][2] ) );
  AND U2510 ( .A(B[1]), .B(A[437]), .Z(\ab[437][1] ) );
  AND U2511 ( .A(A[437]), .B(B[0]), .Z(\ab[437][0] ) );
  AND U2512 ( .A(B[3]), .B(A[436]), .Z(\ab[436][3] ) );
  AND U2513 ( .A(B[2]), .B(A[436]), .Z(\ab[436][2] ) );
  AND U2514 ( .A(B[1]), .B(A[436]), .Z(\ab[436][1] ) );
  AND U2515 ( .A(A[436]), .B(B[0]), .Z(\ab[436][0] ) );
  AND U2516 ( .A(B[3]), .B(A[435]), .Z(\ab[435][3] ) );
  AND U2517 ( .A(B[2]), .B(A[435]), .Z(\ab[435][2] ) );
  AND U2518 ( .A(B[1]), .B(A[435]), .Z(\ab[435][1] ) );
  AND U2519 ( .A(A[435]), .B(B[0]), .Z(\ab[435][0] ) );
  AND U2520 ( .A(B[3]), .B(A[434]), .Z(\ab[434][3] ) );
  AND U2521 ( .A(B[2]), .B(A[434]), .Z(\ab[434][2] ) );
  AND U2522 ( .A(B[1]), .B(A[434]), .Z(\ab[434][1] ) );
  AND U2523 ( .A(A[434]), .B(B[0]), .Z(\ab[434][0] ) );
  AND U2524 ( .A(B[3]), .B(A[433]), .Z(\ab[433][3] ) );
  AND U2525 ( .A(B[2]), .B(A[433]), .Z(\ab[433][2] ) );
  AND U2526 ( .A(B[1]), .B(A[433]), .Z(\ab[433][1] ) );
  AND U2527 ( .A(A[433]), .B(B[0]), .Z(\ab[433][0] ) );
  AND U2528 ( .A(B[3]), .B(A[432]), .Z(\ab[432][3] ) );
  AND U2529 ( .A(B[2]), .B(A[432]), .Z(\ab[432][2] ) );
  AND U2530 ( .A(B[1]), .B(A[432]), .Z(\ab[432][1] ) );
  AND U2531 ( .A(A[432]), .B(B[0]), .Z(\ab[432][0] ) );
  AND U2532 ( .A(B[3]), .B(A[431]), .Z(\ab[431][3] ) );
  AND U2533 ( .A(B[2]), .B(A[431]), .Z(\ab[431][2] ) );
  AND U2534 ( .A(B[1]), .B(A[431]), .Z(\ab[431][1] ) );
  AND U2535 ( .A(A[431]), .B(B[0]), .Z(\ab[431][0] ) );
  AND U2536 ( .A(B[3]), .B(A[430]), .Z(\ab[430][3] ) );
  AND U2537 ( .A(B[2]), .B(A[430]), .Z(\ab[430][2] ) );
  AND U2538 ( .A(B[1]), .B(A[430]), .Z(\ab[430][1] ) );
  AND U2539 ( .A(A[430]), .B(B[0]), .Z(\ab[430][0] ) );
  AND U2540 ( .A(B[3]), .B(A[42]), .Z(\ab[42][3] ) );
  AND U2541 ( .A(B[2]), .B(A[42]), .Z(\ab[42][2] ) );
  AND U2542 ( .A(B[1]), .B(A[42]), .Z(\ab[42][1] ) );
  AND U2543 ( .A(A[42]), .B(B[0]), .Z(\ab[42][0] ) );
  AND U2544 ( .A(B[3]), .B(A[429]), .Z(\ab[429][3] ) );
  AND U2545 ( .A(B[2]), .B(A[429]), .Z(\ab[429][2] ) );
  AND U2546 ( .A(B[1]), .B(A[429]), .Z(\ab[429][1] ) );
  AND U2547 ( .A(A[429]), .B(B[0]), .Z(\ab[429][0] ) );
  AND U2548 ( .A(B[3]), .B(A[428]), .Z(\ab[428][3] ) );
  AND U2549 ( .A(B[2]), .B(A[428]), .Z(\ab[428][2] ) );
  AND U2550 ( .A(B[1]), .B(A[428]), .Z(\ab[428][1] ) );
  AND U2551 ( .A(A[428]), .B(B[0]), .Z(\ab[428][0] ) );
  AND U2552 ( .A(B[3]), .B(A[427]), .Z(\ab[427][3] ) );
  AND U2553 ( .A(B[2]), .B(A[427]), .Z(\ab[427][2] ) );
  AND U2554 ( .A(B[1]), .B(A[427]), .Z(\ab[427][1] ) );
  AND U2555 ( .A(A[427]), .B(B[0]), .Z(\ab[427][0] ) );
  AND U2556 ( .A(B[3]), .B(A[426]), .Z(\ab[426][3] ) );
  AND U2557 ( .A(B[2]), .B(A[426]), .Z(\ab[426][2] ) );
  AND U2558 ( .A(B[1]), .B(A[426]), .Z(\ab[426][1] ) );
  AND U2559 ( .A(A[426]), .B(B[0]), .Z(\ab[426][0] ) );
  AND U2560 ( .A(B[3]), .B(A[425]), .Z(\ab[425][3] ) );
  AND U2561 ( .A(B[2]), .B(A[425]), .Z(\ab[425][2] ) );
  AND U2562 ( .A(B[1]), .B(A[425]), .Z(\ab[425][1] ) );
  AND U2563 ( .A(A[425]), .B(B[0]), .Z(\ab[425][0] ) );
  AND U2564 ( .A(B[3]), .B(A[424]), .Z(\ab[424][3] ) );
  AND U2565 ( .A(B[2]), .B(A[424]), .Z(\ab[424][2] ) );
  AND U2566 ( .A(B[1]), .B(A[424]), .Z(\ab[424][1] ) );
  AND U2567 ( .A(A[424]), .B(B[0]), .Z(\ab[424][0] ) );
  AND U2568 ( .A(B[3]), .B(A[423]), .Z(\ab[423][3] ) );
  AND U2569 ( .A(B[2]), .B(A[423]), .Z(\ab[423][2] ) );
  AND U2570 ( .A(B[1]), .B(A[423]), .Z(\ab[423][1] ) );
  AND U2571 ( .A(A[423]), .B(B[0]), .Z(\ab[423][0] ) );
  AND U2572 ( .A(B[3]), .B(A[422]), .Z(\ab[422][3] ) );
  AND U2573 ( .A(B[2]), .B(A[422]), .Z(\ab[422][2] ) );
  AND U2574 ( .A(B[1]), .B(A[422]), .Z(\ab[422][1] ) );
  AND U2575 ( .A(A[422]), .B(B[0]), .Z(\ab[422][0] ) );
  AND U2576 ( .A(B[3]), .B(A[421]), .Z(\ab[421][3] ) );
  AND U2577 ( .A(B[2]), .B(A[421]), .Z(\ab[421][2] ) );
  AND U2578 ( .A(B[1]), .B(A[421]), .Z(\ab[421][1] ) );
  AND U2579 ( .A(A[421]), .B(B[0]), .Z(\ab[421][0] ) );
  AND U2580 ( .A(B[3]), .B(A[420]), .Z(\ab[420][3] ) );
  AND U2581 ( .A(B[2]), .B(A[420]), .Z(\ab[420][2] ) );
  AND U2582 ( .A(B[1]), .B(A[420]), .Z(\ab[420][1] ) );
  AND U2583 ( .A(A[420]), .B(B[0]), .Z(\ab[420][0] ) );
  AND U2584 ( .A(B[3]), .B(A[41]), .Z(\ab[41][3] ) );
  AND U2585 ( .A(B[2]), .B(A[41]), .Z(\ab[41][2] ) );
  AND U2586 ( .A(B[1]), .B(A[41]), .Z(\ab[41][1] ) );
  AND U2587 ( .A(A[41]), .B(B[0]), .Z(\ab[41][0] ) );
  AND U2588 ( .A(B[3]), .B(A[419]), .Z(\ab[419][3] ) );
  AND U2589 ( .A(B[2]), .B(A[419]), .Z(\ab[419][2] ) );
  AND U2590 ( .A(B[1]), .B(A[419]), .Z(\ab[419][1] ) );
  AND U2591 ( .A(A[419]), .B(B[0]), .Z(\ab[419][0] ) );
  AND U2592 ( .A(B[3]), .B(A[418]), .Z(\ab[418][3] ) );
  AND U2593 ( .A(B[2]), .B(A[418]), .Z(\ab[418][2] ) );
  AND U2594 ( .A(B[1]), .B(A[418]), .Z(\ab[418][1] ) );
  AND U2595 ( .A(A[418]), .B(B[0]), .Z(\ab[418][0] ) );
  AND U2596 ( .A(B[3]), .B(A[417]), .Z(\ab[417][3] ) );
  AND U2597 ( .A(B[2]), .B(A[417]), .Z(\ab[417][2] ) );
  AND U2598 ( .A(B[1]), .B(A[417]), .Z(\ab[417][1] ) );
  AND U2599 ( .A(A[417]), .B(B[0]), .Z(\ab[417][0] ) );
  AND U2600 ( .A(B[3]), .B(A[416]), .Z(\ab[416][3] ) );
  AND U2601 ( .A(B[2]), .B(A[416]), .Z(\ab[416][2] ) );
  AND U2602 ( .A(B[1]), .B(A[416]), .Z(\ab[416][1] ) );
  AND U2603 ( .A(A[416]), .B(B[0]), .Z(\ab[416][0] ) );
  AND U2604 ( .A(B[3]), .B(A[415]), .Z(\ab[415][3] ) );
  AND U2605 ( .A(B[2]), .B(A[415]), .Z(\ab[415][2] ) );
  AND U2606 ( .A(B[1]), .B(A[415]), .Z(\ab[415][1] ) );
  AND U2607 ( .A(A[415]), .B(B[0]), .Z(\ab[415][0] ) );
  AND U2608 ( .A(B[3]), .B(A[414]), .Z(\ab[414][3] ) );
  AND U2609 ( .A(B[2]), .B(A[414]), .Z(\ab[414][2] ) );
  AND U2610 ( .A(B[1]), .B(A[414]), .Z(\ab[414][1] ) );
  AND U2611 ( .A(A[414]), .B(B[0]), .Z(\ab[414][0] ) );
  AND U2612 ( .A(B[3]), .B(A[413]), .Z(\ab[413][3] ) );
  AND U2613 ( .A(B[2]), .B(A[413]), .Z(\ab[413][2] ) );
  AND U2614 ( .A(B[1]), .B(A[413]), .Z(\ab[413][1] ) );
  AND U2615 ( .A(A[413]), .B(B[0]), .Z(\ab[413][0] ) );
  AND U2616 ( .A(B[3]), .B(A[412]), .Z(\ab[412][3] ) );
  AND U2617 ( .A(B[2]), .B(A[412]), .Z(\ab[412][2] ) );
  AND U2618 ( .A(B[1]), .B(A[412]), .Z(\ab[412][1] ) );
  AND U2619 ( .A(A[412]), .B(B[0]), .Z(\ab[412][0] ) );
  AND U2620 ( .A(B[3]), .B(A[411]), .Z(\ab[411][3] ) );
  AND U2621 ( .A(B[2]), .B(A[411]), .Z(\ab[411][2] ) );
  AND U2622 ( .A(B[1]), .B(A[411]), .Z(\ab[411][1] ) );
  AND U2623 ( .A(A[411]), .B(B[0]), .Z(\ab[411][0] ) );
  AND U2624 ( .A(B[3]), .B(A[410]), .Z(\ab[410][3] ) );
  AND U2625 ( .A(B[2]), .B(A[410]), .Z(\ab[410][2] ) );
  AND U2626 ( .A(B[1]), .B(A[410]), .Z(\ab[410][1] ) );
  AND U2627 ( .A(A[410]), .B(B[0]), .Z(\ab[410][0] ) );
  AND U2628 ( .A(B[3]), .B(A[40]), .Z(\ab[40][3] ) );
  AND U2629 ( .A(B[2]), .B(A[40]), .Z(\ab[40][2] ) );
  AND U2630 ( .A(B[1]), .B(A[40]), .Z(\ab[40][1] ) );
  AND U2631 ( .A(A[40]), .B(B[0]), .Z(\ab[40][0] ) );
  AND U2632 ( .A(B[3]), .B(A[409]), .Z(\ab[409][3] ) );
  AND U2633 ( .A(B[2]), .B(A[409]), .Z(\ab[409][2] ) );
  AND U2634 ( .A(B[1]), .B(A[409]), .Z(\ab[409][1] ) );
  AND U2635 ( .A(A[409]), .B(B[0]), .Z(\ab[409][0] ) );
  AND U2636 ( .A(B[3]), .B(A[408]), .Z(\ab[408][3] ) );
  AND U2637 ( .A(B[2]), .B(A[408]), .Z(\ab[408][2] ) );
  AND U2638 ( .A(B[1]), .B(A[408]), .Z(\ab[408][1] ) );
  AND U2639 ( .A(A[408]), .B(B[0]), .Z(\ab[408][0] ) );
  AND U2640 ( .A(B[3]), .B(A[407]), .Z(\ab[407][3] ) );
  AND U2641 ( .A(B[2]), .B(A[407]), .Z(\ab[407][2] ) );
  AND U2642 ( .A(B[1]), .B(A[407]), .Z(\ab[407][1] ) );
  AND U2643 ( .A(A[407]), .B(B[0]), .Z(\ab[407][0] ) );
  AND U2644 ( .A(B[3]), .B(A[406]), .Z(\ab[406][3] ) );
  AND U2645 ( .A(B[2]), .B(A[406]), .Z(\ab[406][2] ) );
  AND U2646 ( .A(B[1]), .B(A[406]), .Z(\ab[406][1] ) );
  AND U2647 ( .A(A[406]), .B(B[0]), .Z(\ab[406][0] ) );
  AND U2648 ( .A(B[3]), .B(A[405]), .Z(\ab[405][3] ) );
  AND U2649 ( .A(B[2]), .B(A[405]), .Z(\ab[405][2] ) );
  AND U2650 ( .A(B[1]), .B(A[405]), .Z(\ab[405][1] ) );
  AND U2651 ( .A(A[405]), .B(B[0]), .Z(\ab[405][0] ) );
  AND U2652 ( .A(B[3]), .B(A[404]), .Z(\ab[404][3] ) );
  AND U2653 ( .A(B[2]), .B(A[404]), .Z(\ab[404][2] ) );
  AND U2654 ( .A(B[1]), .B(A[404]), .Z(\ab[404][1] ) );
  AND U2655 ( .A(A[404]), .B(B[0]), .Z(\ab[404][0] ) );
  AND U2656 ( .A(B[3]), .B(A[403]), .Z(\ab[403][3] ) );
  AND U2657 ( .A(B[2]), .B(A[403]), .Z(\ab[403][2] ) );
  AND U2658 ( .A(B[1]), .B(A[403]), .Z(\ab[403][1] ) );
  AND U2659 ( .A(A[403]), .B(B[0]), .Z(\ab[403][0] ) );
  AND U2660 ( .A(B[3]), .B(A[402]), .Z(\ab[402][3] ) );
  AND U2661 ( .A(B[2]), .B(A[402]), .Z(\ab[402][2] ) );
  AND U2662 ( .A(B[1]), .B(A[402]), .Z(\ab[402][1] ) );
  AND U2663 ( .A(A[402]), .B(B[0]), .Z(\ab[402][0] ) );
  AND U2664 ( .A(B[3]), .B(A[401]), .Z(\ab[401][3] ) );
  AND U2665 ( .A(B[2]), .B(A[401]), .Z(\ab[401][2] ) );
  AND U2666 ( .A(B[1]), .B(A[401]), .Z(\ab[401][1] ) );
  AND U2667 ( .A(A[401]), .B(B[0]), .Z(\ab[401][0] ) );
  AND U2668 ( .A(B[3]), .B(A[400]), .Z(\ab[400][3] ) );
  AND U2669 ( .A(B[2]), .B(A[400]), .Z(\ab[400][2] ) );
  AND U2670 ( .A(B[1]), .B(A[400]), .Z(\ab[400][1] ) );
  AND U2671 ( .A(A[400]), .B(B[0]), .Z(\ab[400][0] ) );
  AND U2672 ( .A(B[3]), .B(A[3]), .Z(\ab[3][3] ) );
  AND U2673 ( .A(B[2]), .B(A[3]), .Z(\ab[3][2] ) );
  AND U2674 ( .A(B[1]), .B(A[3]), .Z(\ab[3][1] ) );
  AND U2675 ( .A(A[3]), .B(B[0]), .Z(\ab[3][0] ) );
  AND U2676 ( .A(B[3]), .B(A[39]), .Z(\ab[39][3] ) );
  AND U2677 ( .A(B[2]), .B(A[39]), .Z(\ab[39][2] ) );
  AND U2678 ( .A(B[1]), .B(A[39]), .Z(\ab[39][1] ) );
  AND U2679 ( .A(A[39]), .B(B[0]), .Z(\ab[39][0] ) );
  AND U2680 ( .A(B[3]), .B(A[399]), .Z(\ab[399][3] ) );
  AND U2681 ( .A(B[2]), .B(A[399]), .Z(\ab[399][2] ) );
  AND U2682 ( .A(B[1]), .B(A[399]), .Z(\ab[399][1] ) );
  AND U2683 ( .A(A[399]), .B(B[0]), .Z(\ab[399][0] ) );
  AND U2684 ( .A(B[3]), .B(A[398]), .Z(\ab[398][3] ) );
  AND U2685 ( .A(B[2]), .B(A[398]), .Z(\ab[398][2] ) );
  AND U2686 ( .A(B[1]), .B(A[398]), .Z(\ab[398][1] ) );
  AND U2687 ( .A(A[398]), .B(B[0]), .Z(\ab[398][0] ) );
  AND U2688 ( .A(B[3]), .B(A[397]), .Z(\ab[397][3] ) );
  AND U2689 ( .A(B[2]), .B(A[397]), .Z(\ab[397][2] ) );
  AND U2690 ( .A(B[1]), .B(A[397]), .Z(\ab[397][1] ) );
  AND U2691 ( .A(A[397]), .B(B[0]), .Z(\ab[397][0] ) );
  AND U2692 ( .A(B[3]), .B(A[396]), .Z(\ab[396][3] ) );
  AND U2693 ( .A(B[2]), .B(A[396]), .Z(\ab[396][2] ) );
  AND U2694 ( .A(B[1]), .B(A[396]), .Z(\ab[396][1] ) );
  AND U2695 ( .A(A[396]), .B(B[0]), .Z(\ab[396][0] ) );
  AND U2696 ( .A(B[3]), .B(A[395]), .Z(\ab[395][3] ) );
  AND U2697 ( .A(B[2]), .B(A[395]), .Z(\ab[395][2] ) );
  AND U2698 ( .A(B[1]), .B(A[395]), .Z(\ab[395][1] ) );
  AND U2699 ( .A(A[395]), .B(B[0]), .Z(\ab[395][0] ) );
  AND U2700 ( .A(B[3]), .B(A[394]), .Z(\ab[394][3] ) );
  AND U2701 ( .A(B[2]), .B(A[394]), .Z(\ab[394][2] ) );
  AND U2702 ( .A(B[1]), .B(A[394]), .Z(\ab[394][1] ) );
  AND U2703 ( .A(A[394]), .B(B[0]), .Z(\ab[394][0] ) );
  AND U2704 ( .A(B[3]), .B(A[393]), .Z(\ab[393][3] ) );
  AND U2705 ( .A(B[2]), .B(A[393]), .Z(\ab[393][2] ) );
  AND U2706 ( .A(B[1]), .B(A[393]), .Z(\ab[393][1] ) );
  AND U2707 ( .A(A[393]), .B(B[0]), .Z(\ab[393][0] ) );
  AND U2708 ( .A(B[3]), .B(A[392]), .Z(\ab[392][3] ) );
  AND U2709 ( .A(B[2]), .B(A[392]), .Z(\ab[392][2] ) );
  AND U2710 ( .A(B[1]), .B(A[392]), .Z(\ab[392][1] ) );
  AND U2711 ( .A(A[392]), .B(B[0]), .Z(\ab[392][0] ) );
  AND U2712 ( .A(B[3]), .B(A[391]), .Z(\ab[391][3] ) );
  AND U2713 ( .A(B[2]), .B(A[391]), .Z(\ab[391][2] ) );
  AND U2714 ( .A(B[1]), .B(A[391]), .Z(\ab[391][1] ) );
  AND U2715 ( .A(A[391]), .B(B[0]), .Z(\ab[391][0] ) );
  AND U2716 ( .A(B[3]), .B(A[390]), .Z(\ab[390][3] ) );
  AND U2717 ( .A(B[2]), .B(A[390]), .Z(\ab[390][2] ) );
  AND U2718 ( .A(B[1]), .B(A[390]), .Z(\ab[390][1] ) );
  AND U2719 ( .A(A[390]), .B(B[0]), .Z(\ab[390][0] ) );
  AND U2720 ( .A(B[3]), .B(A[38]), .Z(\ab[38][3] ) );
  AND U2721 ( .A(B[2]), .B(A[38]), .Z(\ab[38][2] ) );
  AND U2722 ( .A(B[1]), .B(A[38]), .Z(\ab[38][1] ) );
  AND U2723 ( .A(A[38]), .B(B[0]), .Z(\ab[38][0] ) );
  AND U2724 ( .A(B[3]), .B(A[389]), .Z(\ab[389][3] ) );
  AND U2725 ( .A(B[2]), .B(A[389]), .Z(\ab[389][2] ) );
  AND U2726 ( .A(B[1]), .B(A[389]), .Z(\ab[389][1] ) );
  AND U2727 ( .A(A[389]), .B(B[0]), .Z(\ab[389][0] ) );
  AND U2728 ( .A(B[3]), .B(A[388]), .Z(\ab[388][3] ) );
  AND U2729 ( .A(B[2]), .B(A[388]), .Z(\ab[388][2] ) );
  AND U2730 ( .A(B[1]), .B(A[388]), .Z(\ab[388][1] ) );
  AND U2731 ( .A(A[388]), .B(B[0]), .Z(\ab[388][0] ) );
  AND U2732 ( .A(B[3]), .B(A[387]), .Z(\ab[387][3] ) );
  AND U2733 ( .A(B[2]), .B(A[387]), .Z(\ab[387][2] ) );
  AND U2734 ( .A(B[1]), .B(A[387]), .Z(\ab[387][1] ) );
  AND U2735 ( .A(A[387]), .B(B[0]), .Z(\ab[387][0] ) );
  AND U2736 ( .A(B[3]), .B(A[386]), .Z(\ab[386][3] ) );
  AND U2737 ( .A(B[2]), .B(A[386]), .Z(\ab[386][2] ) );
  AND U2738 ( .A(B[1]), .B(A[386]), .Z(\ab[386][1] ) );
  AND U2739 ( .A(A[386]), .B(B[0]), .Z(\ab[386][0] ) );
  AND U2740 ( .A(B[3]), .B(A[385]), .Z(\ab[385][3] ) );
  AND U2741 ( .A(B[2]), .B(A[385]), .Z(\ab[385][2] ) );
  AND U2742 ( .A(B[1]), .B(A[385]), .Z(\ab[385][1] ) );
  AND U2743 ( .A(A[385]), .B(B[0]), .Z(\ab[385][0] ) );
  AND U2744 ( .A(B[3]), .B(A[384]), .Z(\ab[384][3] ) );
  AND U2745 ( .A(B[2]), .B(A[384]), .Z(\ab[384][2] ) );
  AND U2746 ( .A(B[1]), .B(A[384]), .Z(\ab[384][1] ) );
  AND U2747 ( .A(A[384]), .B(B[0]), .Z(\ab[384][0] ) );
  AND U2748 ( .A(B[3]), .B(A[383]), .Z(\ab[383][3] ) );
  AND U2749 ( .A(B[2]), .B(A[383]), .Z(\ab[383][2] ) );
  AND U2750 ( .A(B[1]), .B(A[383]), .Z(\ab[383][1] ) );
  AND U2751 ( .A(A[383]), .B(B[0]), .Z(\ab[383][0] ) );
  AND U2752 ( .A(B[3]), .B(A[382]), .Z(\ab[382][3] ) );
  AND U2753 ( .A(B[2]), .B(A[382]), .Z(\ab[382][2] ) );
  AND U2754 ( .A(B[1]), .B(A[382]), .Z(\ab[382][1] ) );
  AND U2755 ( .A(A[382]), .B(B[0]), .Z(\ab[382][0] ) );
  AND U2756 ( .A(B[3]), .B(A[381]), .Z(\ab[381][3] ) );
  AND U2757 ( .A(B[2]), .B(A[381]), .Z(\ab[381][2] ) );
  AND U2758 ( .A(B[1]), .B(A[381]), .Z(\ab[381][1] ) );
  AND U2759 ( .A(A[381]), .B(B[0]), .Z(\ab[381][0] ) );
  AND U2760 ( .A(B[3]), .B(A[380]), .Z(\ab[380][3] ) );
  AND U2761 ( .A(B[2]), .B(A[380]), .Z(\ab[380][2] ) );
  AND U2762 ( .A(B[1]), .B(A[380]), .Z(\ab[380][1] ) );
  AND U2763 ( .A(A[380]), .B(B[0]), .Z(\ab[380][0] ) );
  AND U2764 ( .A(B[3]), .B(A[37]), .Z(\ab[37][3] ) );
  AND U2765 ( .A(B[2]), .B(A[37]), .Z(\ab[37][2] ) );
  AND U2766 ( .A(B[1]), .B(A[37]), .Z(\ab[37][1] ) );
  AND U2767 ( .A(A[37]), .B(B[0]), .Z(\ab[37][0] ) );
  AND U2768 ( .A(B[3]), .B(A[379]), .Z(\ab[379][3] ) );
  AND U2769 ( .A(B[2]), .B(A[379]), .Z(\ab[379][2] ) );
  AND U2770 ( .A(B[1]), .B(A[379]), .Z(\ab[379][1] ) );
  AND U2771 ( .A(A[379]), .B(B[0]), .Z(\ab[379][0] ) );
  AND U2772 ( .A(B[3]), .B(A[378]), .Z(\ab[378][3] ) );
  AND U2773 ( .A(B[2]), .B(A[378]), .Z(\ab[378][2] ) );
  AND U2774 ( .A(B[1]), .B(A[378]), .Z(\ab[378][1] ) );
  AND U2775 ( .A(A[378]), .B(B[0]), .Z(\ab[378][0] ) );
  AND U2776 ( .A(B[3]), .B(A[377]), .Z(\ab[377][3] ) );
  AND U2777 ( .A(B[2]), .B(A[377]), .Z(\ab[377][2] ) );
  AND U2778 ( .A(B[1]), .B(A[377]), .Z(\ab[377][1] ) );
  AND U2779 ( .A(A[377]), .B(B[0]), .Z(\ab[377][0] ) );
  AND U2780 ( .A(B[3]), .B(A[376]), .Z(\ab[376][3] ) );
  AND U2781 ( .A(B[2]), .B(A[376]), .Z(\ab[376][2] ) );
  AND U2782 ( .A(B[1]), .B(A[376]), .Z(\ab[376][1] ) );
  AND U2783 ( .A(A[376]), .B(B[0]), .Z(\ab[376][0] ) );
  AND U2784 ( .A(B[3]), .B(A[375]), .Z(\ab[375][3] ) );
  AND U2785 ( .A(B[2]), .B(A[375]), .Z(\ab[375][2] ) );
  AND U2786 ( .A(B[1]), .B(A[375]), .Z(\ab[375][1] ) );
  AND U2787 ( .A(A[375]), .B(B[0]), .Z(\ab[375][0] ) );
  AND U2788 ( .A(B[3]), .B(A[374]), .Z(\ab[374][3] ) );
  AND U2789 ( .A(B[2]), .B(A[374]), .Z(\ab[374][2] ) );
  AND U2790 ( .A(B[1]), .B(A[374]), .Z(\ab[374][1] ) );
  AND U2791 ( .A(A[374]), .B(B[0]), .Z(\ab[374][0] ) );
  AND U2792 ( .A(B[3]), .B(A[373]), .Z(\ab[373][3] ) );
  AND U2793 ( .A(B[2]), .B(A[373]), .Z(\ab[373][2] ) );
  AND U2794 ( .A(B[1]), .B(A[373]), .Z(\ab[373][1] ) );
  AND U2795 ( .A(A[373]), .B(B[0]), .Z(\ab[373][0] ) );
  AND U2796 ( .A(B[3]), .B(A[372]), .Z(\ab[372][3] ) );
  AND U2797 ( .A(B[2]), .B(A[372]), .Z(\ab[372][2] ) );
  AND U2798 ( .A(B[1]), .B(A[372]), .Z(\ab[372][1] ) );
  AND U2799 ( .A(A[372]), .B(B[0]), .Z(\ab[372][0] ) );
  AND U2800 ( .A(B[3]), .B(A[371]), .Z(\ab[371][3] ) );
  AND U2801 ( .A(B[2]), .B(A[371]), .Z(\ab[371][2] ) );
  AND U2802 ( .A(B[1]), .B(A[371]), .Z(\ab[371][1] ) );
  AND U2803 ( .A(A[371]), .B(B[0]), .Z(\ab[371][0] ) );
  AND U2804 ( .A(B[3]), .B(A[370]), .Z(\ab[370][3] ) );
  AND U2805 ( .A(B[2]), .B(A[370]), .Z(\ab[370][2] ) );
  AND U2806 ( .A(B[1]), .B(A[370]), .Z(\ab[370][1] ) );
  AND U2807 ( .A(A[370]), .B(B[0]), .Z(\ab[370][0] ) );
  AND U2808 ( .A(B[3]), .B(A[36]), .Z(\ab[36][3] ) );
  AND U2809 ( .A(B[2]), .B(A[36]), .Z(\ab[36][2] ) );
  AND U2810 ( .A(B[1]), .B(A[36]), .Z(\ab[36][1] ) );
  AND U2811 ( .A(A[36]), .B(B[0]), .Z(\ab[36][0] ) );
  AND U2812 ( .A(B[3]), .B(A[369]), .Z(\ab[369][3] ) );
  AND U2813 ( .A(B[2]), .B(A[369]), .Z(\ab[369][2] ) );
  AND U2814 ( .A(B[1]), .B(A[369]), .Z(\ab[369][1] ) );
  AND U2815 ( .A(A[369]), .B(B[0]), .Z(\ab[369][0] ) );
  AND U2816 ( .A(B[3]), .B(A[368]), .Z(\ab[368][3] ) );
  AND U2817 ( .A(B[2]), .B(A[368]), .Z(\ab[368][2] ) );
  AND U2818 ( .A(B[1]), .B(A[368]), .Z(\ab[368][1] ) );
  AND U2819 ( .A(A[368]), .B(B[0]), .Z(\ab[368][0] ) );
  AND U2820 ( .A(B[3]), .B(A[367]), .Z(\ab[367][3] ) );
  AND U2821 ( .A(B[2]), .B(A[367]), .Z(\ab[367][2] ) );
  AND U2822 ( .A(B[1]), .B(A[367]), .Z(\ab[367][1] ) );
  AND U2823 ( .A(A[367]), .B(B[0]), .Z(\ab[367][0] ) );
  AND U2824 ( .A(B[3]), .B(A[366]), .Z(\ab[366][3] ) );
  AND U2825 ( .A(B[2]), .B(A[366]), .Z(\ab[366][2] ) );
  AND U2826 ( .A(B[1]), .B(A[366]), .Z(\ab[366][1] ) );
  AND U2827 ( .A(A[366]), .B(B[0]), .Z(\ab[366][0] ) );
  AND U2828 ( .A(B[3]), .B(A[365]), .Z(\ab[365][3] ) );
  AND U2829 ( .A(B[2]), .B(A[365]), .Z(\ab[365][2] ) );
  AND U2830 ( .A(B[1]), .B(A[365]), .Z(\ab[365][1] ) );
  AND U2831 ( .A(A[365]), .B(B[0]), .Z(\ab[365][0] ) );
  AND U2832 ( .A(B[3]), .B(A[364]), .Z(\ab[364][3] ) );
  AND U2833 ( .A(B[2]), .B(A[364]), .Z(\ab[364][2] ) );
  AND U2834 ( .A(B[1]), .B(A[364]), .Z(\ab[364][1] ) );
  AND U2835 ( .A(A[364]), .B(B[0]), .Z(\ab[364][0] ) );
  AND U2836 ( .A(B[3]), .B(A[363]), .Z(\ab[363][3] ) );
  AND U2837 ( .A(B[2]), .B(A[363]), .Z(\ab[363][2] ) );
  AND U2838 ( .A(B[1]), .B(A[363]), .Z(\ab[363][1] ) );
  AND U2839 ( .A(A[363]), .B(B[0]), .Z(\ab[363][0] ) );
  AND U2840 ( .A(B[3]), .B(A[362]), .Z(\ab[362][3] ) );
  AND U2841 ( .A(B[2]), .B(A[362]), .Z(\ab[362][2] ) );
  AND U2842 ( .A(B[1]), .B(A[362]), .Z(\ab[362][1] ) );
  AND U2843 ( .A(A[362]), .B(B[0]), .Z(\ab[362][0] ) );
  AND U2844 ( .A(B[3]), .B(A[361]), .Z(\ab[361][3] ) );
  AND U2845 ( .A(B[2]), .B(A[361]), .Z(\ab[361][2] ) );
  AND U2846 ( .A(B[1]), .B(A[361]), .Z(\ab[361][1] ) );
  AND U2847 ( .A(A[361]), .B(B[0]), .Z(\ab[361][0] ) );
  AND U2848 ( .A(B[3]), .B(A[360]), .Z(\ab[360][3] ) );
  AND U2849 ( .A(B[2]), .B(A[360]), .Z(\ab[360][2] ) );
  AND U2850 ( .A(B[1]), .B(A[360]), .Z(\ab[360][1] ) );
  AND U2851 ( .A(A[360]), .B(B[0]), .Z(\ab[360][0] ) );
  AND U2852 ( .A(B[3]), .B(A[35]), .Z(\ab[35][3] ) );
  AND U2853 ( .A(B[2]), .B(A[35]), .Z(\ab[35][2] ) );
  AND U2854 ( .A(B[1]), .B(A[35]), .Z(\ab[35][1] ) );
  AND U2855 ( .A(A[35]), .B(B[0]), .Z(\ab[35][0] ) );
  AND U2856 ( .A(B[3]), .B(A[359]), .Z(\ab[359][3] ) );
  AND U2857 ( .A(B[2]), .B(A[359]), .Z(\ab[359][2] ) );
  AND U2858 ( .A(B[1]), .B(A[359]), .Z(\ab[359][1] ) );
  AND U2859 ( .A(A[359]), .B(B[0]), .Z(\ab[359][0] ) );
  AND U2860 ( .A(B[3]), .B(A[358]), .Z(\ab[358][3] ) );
  AND U2861 ( .A(B[2]), .B(A[358]), .Z(\ab[358][2] ) );
  AND U2862 ( .A(B[1]), .B(A[358]), .Z(\ab[358][1] ) );
  AND U2863 ( .A(A[358]), .B(B[0]), .Z(\ab[358][0] ) );
  AND U2864 ( .A(B[3]), .B(A[357]), .Z(\ab[357][3] ) );
  AND U2865 ( .A(B[2]), .B(A[357]), .Z(\ab[357][2] ) );
  AND U2866 ( .A(B[1]), .B(A[357]), .Z(\ab[357][1] ) );
  AND U2867 ( .A(A[357]), .B(B[0]), .Z(\ab[357][0] ) );
  AND U2868 ( .A(B[3]), .B(A[356]), .Z(\ab[356][3] ) );
  AND U2869 ( .A(B[2]), .B(A[356]), .Z(\ab[356][2] ) );
  AND U2870 ( .A(B[1]), .B(A[356]), .Z(\ab[356][1] ) );
  AND U2871 ( .A(A[356]), .B(B[0]), .Z(\ab[356][0] ) );
  AND U2872 ( .A(B[3]), .B(A[355]), .Z(\ab[355][3] ) );
  AND U2873 ( .A(B[2]), .B(A[355]), .Z(\ab[355][2] ) );
  AND U2874 ( .A(B[1]), .B(A[355]), .Z(\ab[355][1] ) );
  AND U2875 ( .A(A[355]), .B(B[0]), .Z(\ab[355][0] ) );
  AND U2876 ( .A(B[3]), .B(A[354]), .Z(\ab[354][3] ) );
  AND U2877 ( .A(B[2]), .B(A[354]), .Z(\ab[354][2] ) );
  AND U2878 ( .A(B[1]), .B(A[354]), .Z(\ab[354][1] ) );
  AND U2879 ( .A(A[354]), .B(B[0]), .Z(\ab[354][0] ) );
  AND U2880 ( .A(B[3]), .B(A[353]), .Z(\ab[353][3] ) );
  AND U2881 ( .A(B[2]), .B(A[353]), .Z(\ab[353][2] ) );
  AND U2882 ( .A(B[1]), .B(A[353]), .Z(\ab[353][1] ) );
  AND U2883 ( .A(A[353]), .B(B[0]), .Z(\ab[353][0] ) );
  AND U2884 ( .A(B[3]), .B(A[352]), .Z(\ab[352][3] ) );
  AND U2885 ( .A(B[2]), .B(A[352]), .Z(\ab[352][2] ) );
  AND U2886 ( .A(B[1]), .B(A[352]), .Z(\ab[352][1] ) );
  AND U2887 ( .A(A[352]), .B(B[0]), .Z(\ab[352][0] ) );
  AND U2888 ( .A(B[3]), .B(A[351]), .Z(\ab[351][3] ) );
  AND U2889 ( .A(B[2]), .B(A[351]), .Z(\ab[351][2] ) );
  AND U2890 ( .A(B[1]), .B(A[351]), .Z(\ab[351][1] ) );
  AND U2891 ( .A(A[351]), .B(B[0]), .Z(\ab[351][0] ) );
  AND U2892 ( .A(B[3]), .B(A[350]), .Z(\ab[350][3] ) );
  AND U2893 ( .A(B[2]), .B(A[350]), .Z(\ab[350][2] ) );
  AND U2894 ( .A(B[1]), .B(A[350]), .Z(\ab[350][1] ) );
  AND U2895 ( .A(A[350]), .B(B[0]), .Z(\ab[350][0] ) );
  AND U2896 ( .A(B[3]), .B(A[34]), .Z(\ab[34][3] ) );
  AND U2897 ( .A(B[2]), .B(A[34]), .Z(\ab[34][2] ) );
  AND U2898 ( .A(B[1]), .B(A[34]), .Z(\ab[34][1] ) );
  AND U2899 ( .A(A[34]), .B(B[0]), .Z(\ab[34][0] ) );
  AND U2900 ( .A(B[3]), .B(A[349]), .Z(\ab[349][3] ) );
  AND U2901 ( .A(B[2]), .B(A[349]), .Z(\ab[349][2] ) );
  AND U2902 ( .A(B[1]), .B(A[349]), .Z(\ab[349][1] ) );
  AND U2903 ( .A(A[349]), .B(B[0]), .Z(\ab[349][0] ) );
  AND U2904 ( .A(B[3]), .B(A[348]), .Z(\ab[348][3] ) );
  AND U2905 ( .A(B[2]), .B(A[348]), .Z(\ab[348][2] ) );
  AND U2906 ( .A(B[1]), .B(A[348]), .Z(\ab[348][1] ) );
  AND U2907 ( .A(A[348]), .B(B[0]), .Z(\ab[348][0] ) );
  AND U2908 ( .A(B[3]), .B(A[347]), .Z(\ab[347][3] ) );
  AND U2909 ( .A(B[2]), .B(A[347]), .Z(\ab[347][2] ) );
  AND U2910 ( .A(B[1]), .B(A[347]), .Z(\ab[347][1] ) );
  AND U2911 ( .A(A[347]), .B(B[0]), .Z(\ab[347][0] ) );
  AND U2912 ( .A(B[3]), .B(A[346]), .Z(\ab[346][3] ) );
  AND U2913 ( .A(B[2]), .B(A[346]), .Z(\ab[346][2] ) );
  AND U2914 ( .A(B[1]), .B(A[346]), .Z(\ab[346][1] ) );
  AND U2915 ( .A(A[346]), .B(B[0]), .Z(\ab[346][0] ) );
  AND U2916 ( .A(B[3]), .B(A[345]), .Z(\ab[345][3] ) );
  AND U2917 ( .A(B[2]), .B(A[345]), .Z(\ab[345][2] ) );
  AND U2918 ( .A(B[1]), .B(A[345]), .Z(\ab[345][1] ) );
  AND U2919 ( .A(A[345]), .B(B[0]), .Z(\ab[345][0] ) );
  AND U2920 ( .A(B[3]), .B(A[344]), .Z(\ab[344][3] ) );
  AND U2921 ( .A(B[2]), .B(A[344]), .Z(\ab[344][2] ) );
  AND U2922 ( .A(B[1]), .B(A[344]), .Z(\ab[344][1] ) );
  AND U2923 ( .A(A[344]), .B(B[0]), .Z(\ab[344][0] ) );
  AND U2924 ( .A(B[3]), .B(A[343]), .Z(\ab[343][3] ) );
  AND U2925 ( .A(B[2]), .B(A[343]), .Z(\ab[343][2] ) );
  AND U2926 ( .A(B[1]), .B(A[343]), .Z(\ab[343][1] ) );
  AND U2927 ( .A(A[343]), .B(B[0]), .Z(\ab[343][0] ) );
  AND U2928 ( .A(B[3]), .B(A[342]), .Z(\ab[342][3] ) );
  AND U2929 ( .A(B[2]), .B(A[342]), .Z(\ab[342][2] ) );
  AND U2930 ( .A(B[1]), .B(A[342]), .Z(\ab[342][1] ) );
  AND U2931 ( .A(A[342]), .B(B[0]), .Z(\ab[342][0] ) );
  AND U2932 ( .A(B[3]), .B(A[341]), .Z(\ab[341][3] ) );
  AND U2933 ( .A(B[2]), .B(A[341]), .Z(\ab[341][2] ) );
  AND U2934 ( .A(B[1]), .B(A[341]), .Z(\ab[341][1] ) );
  AND U2935 ( .A(A[341]), .B(B[0]), .Z(\ab[341][0] ) );
  AND U2936 ( .A(B[3]), .B(A[340]), .Z(\ab[340][3] ) );
  AND U2937 ( .A(B[2]), .B(A[340]), .Z(\ab[340][2] ) );
  AND U2938 ( .A(B[1]), .B(A[340]), .Z(\ab[340][1] ) );
  AND U2939 ( .A(A[340]), .B(B[0]), .Z(\ab[340][0] ) );
  AND U2940 ( .A(B[3]), .B(A[33]), .Z(\ab[33][3] ) );
  AND U2941 ( .A(B[2]), .B(A[33]), .Z(\ab[33][2] ) );
  AND U2942 ( .A(B[1]), .B(A[33]), .Z(\ab[33][1] ) );
  AND U2943 ( .A(A[33]), .B(B[0]), .Z(\ab[33][0] ) );
  AND U2944 ( .A(B[3]), .B(A[339]), .Z(\ab[339][3] ) );
  AND U2945 ( .A(B[2]), .B(A[339]), .Z(\ab[339][2] ) );
  AND U2946 ( .A(B[1]), .B(A[339]), .Z(\ab[339][1] ) );
  AND U2947 ( .A(A[339]), .B(B[0]), .Z(\ab[339][0] ) );
  AND U2948 ( .A(B[3]), .B(A[338]), .Z(\ab[338][3] ) );
  AND U2949 ( .A(B[2]), .B(A[338]), .Z(\ab[338][2] ) );
  AND U2950 ( .A(B[1]), .B(A[338]), .Z(\ab[338][1] ) );
  AND U2951 ( .A(A[338]), .B(B[0]), .Z(\ab[338][0] ) );
  AND U2952 ( .A(B[3]), .B(A[337]), .Z(\ab[337][3] ) );
  AND U2953 ( .A(B[2]), .B(A[337]), .Z(\ab[337][2] ) );
  AND U2954 ( .A(B[1]), .B(A[337]), .Z(\ab[337][1] ) );
  AND U2955 ( .A(A[337]), .B(B[0]), .Z(\ab[337][0] ) );
  AND U2956 ( .A(B[3]), .B(A[336]), .Z(\ab[336][3] ) );
  AND U2957 ( .A(B[2]), .B(A[336]), .Z(\ab[336][2] ) );
  AND U2958 ( .A(B[1]), .B(A[336]), .Z(\ab[336][1] ) );
  AND U2959 ( .A(A[336]), .B(B[0]), .Z(\ab[336][0] ) );
  AND U2960 ( .A(B[3]), .B(A[335]), .Z(\ab[335][3] ) );
  AND U2961 ( .A(B[2]), .B(A[335]), .Z(\ab[335][2] ) );
  AND U2962 ( .A(B[1]), .B(A[335]), .Z(\ab[335][1] ) );
  AND U2963 ( .A(A[335]), .B(B[0]), .Z(\ab[335][0] ) );
  AND U2964 ( .A(B[3]), .B(A[334]), .Z(\ab[334][3] ) );
  AND U2965 ( .A(B[2]), .B(A[334]), .Z(\ab[334][2] ) );
  AND U2966 ( .A(B[1]), .B(A[334]), .Z(\ab[334][1] ) );
  AND U2967 ( .A(A[334]), .B(B[0]), .Z(\ab[334][0] ) );
  AND U2968 ( .A(B[3]), .B(A[333]), .Z(\ab[333][3] ) );
  AND U2969 ( .A(B[2]), .B(A[333]), .Z(\ab[333][2] ) );
  AND U2970 ( .A(B[1]), .B(A[333]), .Z(\ab[333][1] ) );
  AND U2971 ( .A(A[333]), .B(B[0]), .Z(\ab[333][0] ) );
  AND U2972 ( .A(B[3]), .B(A[332]), .Z(\ab[332][3] ) );
  AND U2973 ( .A(B[2]), .B(A[332]), .Z(\ab[332][2] ) );
  AND U2974 ( .A(B[1]), .B(A[332]), .Z(\ab[332][1] ) );
  AND U2975 ( .A(A[332]), .B(B[0]), .Z(\ab[332][0] ) );
  AND U2976 ( .A(B[3]), .B(A[331]), .Z(\ab[331][3] ) );
  AND U2977 ( .A(B[2]), .B(A[331]), .Z(\ab[331][2] ) );
  AND U2978 ( .A(B[1]), .B(A[331]), .Z(\ab[331][1] ) );
  AND U2979 ( .A(A[331]), .B(B[0]), .Z(\ab[331][0] ) );
  AND U2980 ( .A(B[3]), .B(A[330]), .Z(\ab[330][3] ) );
  AND U2981 ( .A(B[2]), .B(A[330]), .Z(\ab[330][2] ) );
  AND U2982 ( .A(B[1]), .B(A[330]), .Z(\ab[330][1] ) );
  AND U2983 ( .A(A[330]), .B(B[0]), .Z(\ab[330][0] ) );
  AND U2984 ( .A(B[3]), .B(A[32]), .Z(\ab[32][3] ) );
  AND U2985 ( .A(B[2]), .B(A[32]), .Z(\ab[32][2] ) );
  AND U2986 ( .A(B[1]), .B(A[32]), .Z(\ab[32][1] ) );
  AND U2987 ( .A(A[32]), .B(B[0]), .Z(\ab[32][0] ) );
  AND U2988 ( .A(B[3]), .B(A[329]), .Z(\ab[329][3] ) );
  AND U2989 ( .A(B[2]), .B(A[329]), .Z(\ab[329][2] ) );
  AND U2990 ( .A(B[1]), .B(A[329]), .Z(\ab[329][1] ) );
  AND U2991 ( .A(A[329]), .B(B[0]), .Z(\ab[329][0] ) );
  AND U2992 ( .A(B[3]), .B(A[328]), .Z(\ab[328][3] ) );
  AND U2993 ( .A(B[2]), .B(A[328]), .Z(\ab[328][2] ) );
  AND U2994 ( .A(B[1]), .B(A[328]), .Z(\ab[328][1] ) );
  AND U2995 ( .A(A[328]), .B(B[0]), .Z(\ab[328][0] ) );
  AND U2996 ( .A(B[3]), .B(A[327]), .Z(\ab[327][3] ) );
  AND U2997 ( .A(B[2]), .B(A[327]), .Z(\ab[327][2] ) );
  AND U2998 ( .A(B[1]), .B(A[327]), .Z(\ab[327][1] ) );
  AND U2999 ( .A(A[327]), .B(B[0]), .Z(\ab[327][0] ) );
  AND U3000 ( .A(B[3]), .B(A[326]), .Z(\ab[326][3] ) );
  AND U3001 ( .A(B[2]), .B(A[326]), .Z(\ab[326][2] ) );
  AND U3002 ( .A(B[1]), .B(A[326]), .Z(\ab[326][1] ) );
  AND U3003 ( .A(A[326]), .B(B[0]), .Z(\ab[326][0] ) );
  AND U3004 ( .A(B[3]), .B(A[325]), .Z(\ab[325][3] ) );
  AND U3005 ( .A(B[2]), .B(A[325]), .Z(\ab[325][2] ) );
  AND U3006 ( .A(B[1]), .B(A[325]), .Z(\ab[325][1] ) );
  AND U3007 ( .A(A[325]), .B(B[0]), .Z(\ab[325][0] ) );
  AND U3008 ( .A(B[3]), .B(A[324]), .Z(\ab[324][3] ) );
  AND U3009 ( .A(B[2]), .B(A[324]), .Z(\ab[324][2] ) );
  AND U3010 ( .A(B[1]), .B(A[324]), .Z(\ab[324][1] ) );
  AND U3011 ( .A(A[324]), .B(B[0]), .Z(\ab[324][0] ) );
  AND U3012 ( .A(B[3]), .B(A[323]), .Z(\ab[323][3] ) );
  AND U3013 ( .A(B[2]), .B(A[323]), .Z(\ab[323][2] ) );
  AND U3014 ( .A(B[1]), .B(A[323]), .Z(\ab[323][1] ) );
  AND U3015 ( .A(A[323]), .B(B[0]), .Z(\ab[323][0] ) );
  AND U3016 ( .A(B[3]), .B(A[322]), .Z(\ab[322][3] ) );
  AND U3017 ( .A(B[2]), .B(A[322]), .Z(\ab[322][2] ) );
  AND U3018 ( .A(B[1]), .B(A[322]), .Z(\ab[322][1] ) );
  AND U3019 ( .A(A[322]), .B(B[0]), .Z(\ab[322][0] ) );
  AND U3020 ( .A(B[3]), .B(A[321]), .Z(\ab[321][3] ) );
  AND U3021 ( .A(B[2]), .B(A[321]), .Z(\ab[321][2] ) );
  AND U3022 ( .A(B[1]), .B(A[321]), .Z(\ab[321][1] ) );
  AND U3023 ( .A(A[321]), .B(B[0]), .Z(\ab[321][0] ) );
  AND U3024 ( .A(B[3]), .B(A[320]), .Z(\ab[320][3] ) );
  AND U3025 ( .A(B[2]), .B(A[320]), .Z(\ab[320][2] ) );
  AND U3026 ( .A(B[1]), .B(A[320]), .Z(\ab[320][1] ) );
  AND U3027 ( .A(A[320]), .B(B[0]), .Z(\ab[320][0] ) );
  AND U3028 ( .A(B[3]), .B(A[31]), .Z(\ab[31][3] ) );
  AND U3029 ( .A(B[2]), .B(A[31]), .Z(\ab[31][2] ) );
  AND U3030 ( .A(B[1]), .B(A[31]), .Z(\ab[31][1] ) );
  AND U3031 ( .A(A[31]), .B(B[0]), .Z(\ab[31][0] ) );
  AND U3032 ( .A(B[3]), .B(A[319]), .Z(\ab[319][3] ) );
  AND U3033 ( .A(B[2]), .B(A[319]), .Z(\ab[319][2] ) );
  AND U3034 ( .A(B[1]), .B(A[319]), .Z(\ab[319][1] ) );
  AND U3035 ( .A(A[319]), .B(B[0]), .Z(\ab[319][0] ) );
  AND U3036 ( .A(B[3]), .B(A[318]), .Z(\ab[318][3] ) );
  AND U3037 ( .A(B[2]), .B(A[318]), .Z(\ab[318][2] ) );
  AND U3038 ( .A(B[1]), .B(A[318]), .Z(\ab[318][1] ) );
  AND U3039 ( .A(A[318]), .B(B[0]), .Z(\ab[318][0] ) );
  AND U3040 ( .A(B[3]), .B(A[317]), .Z(\ab[317][3] ) );
  AND U3041 ( .A(B[2]), .B(A[317]), .Z(\ab[317][2] ) );
  AND U3042 ( .A(B[1]), .B(A[317]), .Z(\ab[317][1] ) );
  AND U3043 ( .A(A[317]), .B(B[0]), .Z(\ab[317][0] ) );
  AND U3044 ( .A(B[3]), .B(A[316]), .Z(\ab[316][3] ) );
  AND U3045 ( .A(B[2]), .B(A[316]), .Z(\ab[316][2] ) );
  AND U3046 ( .A(B[1]), .B(A[316]), .Z(\ab[316][1] ) );
  AND U3047 ( .A(A[316]), .B(B[0]), .Z(\ab[316][0] ) );
  AND U3048 ( .A(B[3]), .B(A[315]), .Z(\ab[315][3] ) );
  AND U3049 ( .A(B[2]), .B(A[315]), .Z(\ab[315][2] ) );
  AND U3050 ( .A(B[1]), .B(A[315]), .Z(\ab[315][1] ) );
  AND U3051 ( .A(A[315]), .B(B[0]), .Z(\ab[315][0] ) );
  AND U3052 ( .A(B[3]), .B(A[314]), .Z(\ab[314][3] ) );
  AND U3053 ( .A(B[2]), .B(A[314]), .Z(\ab[314][2] ) );
  AND U3054 ( .A(B[1]), .B(A[314]), .Z(\ab[314][1] ) );
  AND U3055 ( .A(A[314]), .B(B[0]), .Z(\ab[314][0] ) );
  AND U3056 ( .A(B[3]), .B(A[313]), .Z(\ab[313][3] ) );
  AND U3057 ( .A(B[2]), .B(A[313]), .Z(\ab[313][2] ) );
  AND U3058 ( .A(B[1]), .B(A[313]), .Z(\ab[313][1] ) );
  AND U3059 ( .A(A[313]), .B(B[0]), .Z(\ab[313][0] ) );
  AND U3060 ( .A(B[3]), .B(A[312]), .Z(\ab[312][3] ) );
  AND U3061 ( .A(B[2]), .B(A[312]), .Z(\ab[312][2] ) );
  AND U3062 ( .A(B[1]), .B(A[312]), .Z(\ab[312][1] ) );
  AND U3063 ( .A(A[312]), .B(B[0]), .Z(\ab[312][0] ) );
  AND U3064 ( .A(B[3]), .B(A[311]), .Z(\ab[311][3] ) );
  AND U3065 ( .A(B[2]), .B(A[311]), .Z(\ab[311][2] ) );
  AND U3066 ( .A(B[1]), .B(A[311]), .Z(\ab[311][1] ) );
  AND U3067 ( .A(A[311]), .B(B[0]), .Z(\ab[311][0] ) );
  AND U3068 ( .A(B[3]), .B(A[310]), .Z(\ab[310][3] ) );
  AND U3069 ( .A(B[2]), .B(A[310]), .Z(\ab[310][2] ) );
  AND U3070 ( .A(B[1]), .B(A[310]), .Z(\ab[310][1] ) );
  AND U3071 ( .A(A[310]), .B(B[0]), .Z(\ab[310][0] ) );
  AND U3072 ( .A(B[3]), .B(A[30]), .Z(\ab[30][3] ) );
  AND U3073 ( .A(B[2]), .B(A[30]), .Z(\ab[30][2] ) );
  AND U3074 ( .A(B[1]), .B(A[30]), .Z(\ab[30][1] ) );
  AND U3075 ( .A(A[30]), .B(B[0]), .Z(\ab[30][0] ) );
  AND U3076 ( .A(B[3]), .B(A[309]), .Z(\ab[309][3] ) );
  AND U3077 ( .A(B[2]), .B(A[309]), .Z(\ab[309][2] ) );
  AND U3078 ( .A(B[1]), .B(A[309]), .Z(\ab[309][1] ) );
  AND U3079 ( .A(A[309]), .B(B[0]), .Z(\ab[309][0] ) );
  AND U3080 ( .A(B[3]), .B(A[308]), .Z(\ab[308][3] ) );
  AND U3081 ( .A(B[2]), .B(A[308]), .Z(\ab[308][2] ) );
  AND U3082 ( .A(B[1]), .B(A[308]), .Z(\ab[308][1] ) );
  AND U3083 ( .A(A[308]), .B(B[0]), .Z(\ab[308][0] ) );
  AND U3084 ( .A(B[3]), .B(A[307]), .Z(\ab[307][3] ) );
  AND U3085 ( .A(B[2]), .B(A[307]), .Z(\ab[307][2] ) );
  AND U3086 ( .A(B[1]), .B(A[307]), .Z(\ab[307][1] ) );
  AND U3087 ( .A(A[307]), .B(B[0]), .Z(\ab[307][0] ) );
  AND U3088 ( .A(B[3]), .B(A[306]), .Z(\ab[306][3] ) );
  AND U3089 ( .A(B[2]), .B(A[306]), .Z(\ab[306][2] ) );
  AND U3090 ( .A(B[1]), .B(A[306]), .Z(\ab[306][1] ) );
  AND U3091 ( .A(A[306]), .B(B[0]), .Z(\ab[306][0] ) );
  AND U3092 ( .A(B[3]), .B(A[305]), .Z(\ab[305][3] ) );
  AND U3093 ( .A(B[2]), .B(A[305]), .Z(\ab[305][2] ) );
  AND U3094 ( .A(B[1]), .B(A[305]), .Z(\ab[305][1] ) );
  AND U3095 ( .A(A[305]), .B(B[0]), .Z(\ab[305][0] ) );
  AND U3096 ( .A(B[3]), .B(A[304]), .Z(\ab[304][3] ) );
  AND U3097 ( .A(B[2]), .B(A[304]), .Z(\ab[304][2] ) );
  AND U3098 ( .A(B[1]), .B(A[304]), .Z(\ab[304][1] ) );
  AND U3099 ( .A(A[304]), .B(B[0]), .Z(\ab[304][0] ) );
  AND U3100 ( .A(B[3]), .B(A[303]), .Z(\ab[303][3] ) );
  AND U3101 ( .A(B[2]), .B(A[303]), .Z(\ab[303][2] ) );
  AND U3102 ( .A(B[1]), .B(A[303]), .Z(\ab[303][1] ) );
  AND U3103 ( .A(A[303]), .B(B[0]), .Z(\ab[303][0] ) );
  AND U3104 ( .A(B[3]), .B(A[302]), .Z(\ab[302][3] ) );
  AND U3105 ( .A(B[2]), .B(A[302]), .Z(\ab[302][2] ) );
  AND U3106 ( .A(B[1]), .B(A[302]), .Z(\ab[302][1] ) );
  AND U3107 ( .A(A[302]), .B(B[0]), .Z(\ab[302][0] ) );
  AND U3108 ( .A(B[3]), .B(A[301]), .Z(\ab[301][3] ) );
  AND U3109 ( .A(B[2]), .B(A[301]), .Z(\ab[301][2] ) );
  AND U3110 ( .A(B[1]), .B(A[301]), .Z(\ab[301][1] ) );
  AND U3111 ( .A(A[301]), .B(B[0]), .Z(\ab[301][0] ) );
  AND U3112 ( .A(B[3]), .B(A[300]), .Z(\ab[300][3] ) );
  AND U3113 ( .A(B[2]), .B(A[300]), .Z(\ab[300][2] ) );
  AND U3114 ( .A(B[1]), .B(A[300]), .Z(\ab[300][1] ) );
  AND U3115 ( .A(A[300]), .B(B[0]), .Z(\ab[300][0] ) );
  AND U3116 ( .A(B[3]), .B(A[2]), .Z(\ab[2][3] ) );
  AND U3117 ( .A(B[2]), .B(A[2]), .Z(\ab[2][2] ) );
  AND U3118 ( .A(B[1]), .B(A[2]), .Z(\ab[2][1] ) );
  AND U3119 ( .A(A[2]), .B(B[0]), .Z(\ab[2][0] ) );
  AND U3120 ( .A(B[3]), .B(A[29]), .Z(\ab[29][3] ) );
  AND U3121 ( .A(B[2]), .B(A[29]), .Z(\ab[29][2] ) );
  AND U3122 ( .A(B[1]), .B(A[29]), .Z(\ab[29][1] ) );
  AND U3123 ( .A(A[29]), .B(B[0]), .Z(\ab[29][0] ) );
  AND U3124 ( .A(B[3]), .B(A[299]), .Z(\ab[299][3] ) );
  AND U3125 ( .A(B[2]), .B(A[299]), .Z(\ab[299][2] ) );
  AND U3126 ( .A(B[1]), .B(A[299]), .Z(\ab[299][1] ) );
  AND U3127 ( .A(A[299]), .B(B[0]), .Z(\ab[299][0] ) );
  AND U3128 ( .A(B[3]), .B(A[298]), .Z(\ab[298][3] ) );
  AND U3129 ( .A(B[2]), .B(A[298]), .Z(\ab[298][2] ) );
  AND U3130 ( .A(B[1]), .B(A[298]), .Z(\ab[298][1] ) );
  AND U3131 ( .A(A[298]), .B(B[0]), .Z(\ab[298][0] ) );
  AND U3132 ( .A(B[3]), .B(A[297]), .Z(\ab[297][3] ) );
  AND U3133 ( .A(B[2]), .B(A[297]), .Z(\ab[297][2] ) );
  AND U3134 ( .A(B[1]), .B(A[297]), .Z(\ab[297][1] ) );
  AND U3135 ( .A(A[297]), .B(B[0]), .Z(\ab[297][0] ) );
  AND U3136 ( .A(B[3]), .B(A[296]), .Z(\ab[296][3] ) );
  AND U3137 ( .A(B[2]), .B(A[296]), .Z(\ab[296][2] ) );
  AND U3138 ( .A(B[1]), .B(A[296]), .Z(\ab[296][1] ) );
  AND U3139 ( .A(A[296]), .B(B[0]), .Z(\ab[296][0] ) );
  AND U3140 ( .A(B[3]), .B(A[295]), .Z(\ab[295][3] ) );
  AND U3141 ( .A(B[2]), .B(A[295]), .Z(\ab[295][2] ) );
  AND U3142 ( .A(B[1]), .B(A[295]), .Z(\ab[295][1] ) );
  AND U3143 ( .A(A[295]), .B(B[0]), .Z(\ab[295][0] ) );
  AND U3144 ( .A(B[3]), .B(A[294]), .Z(\ab[294][3] ) );
  AND U3145 ( .A(B[2]), .B(A[294]), .Z(\ab[294][2] ) );
  AND U3146 ( .A(B[1]), .B(A[294]), .Z(\ab[294][1] ) );
  AND U3147 ( .A(A[294]), .B(B[0]), .Z(\ab[294][0] ) );
  AND U3148 ( .A(B[3]), .B(A[293]), .Z(\ab[293][3] ) );
  AND U3149 ( .A(B[2]), .B(A[293]), .Z(\ab[293][2] ) );
  AND U3150 ( .A(B[1]), .B(A[293]), .Z(\ab[293][1] ) );
  AND U3151 ( .A(A[293]), .B(B[0]), .Z(\ab[293][0] ) );
  AND U3152 ( .A(B[3]), .B(A[292]), .Z(\ab[292][3] ) );
  AND U3153 ( .A(B[2]), .B(A[292]), .Z(\ab[292][2] ) );
  AND U3154 ( .A(B[1]), .B(A[292]), .Z(\ab[292][1] ) );
  AND U3155 ( .A(A[292]), .B(B[0]), .Z(\ab[292][0] ) );
  AND U3156 ( .A(B[3]), .B(A[291]), .Z(\ab[291][3] ) );
  AND U3157 ( .A(B[2]), .B(A[291]), .Z(\ab[291][2] ) );
  AND U3158 ( .A(B[1]), .B(A[291]), .Z(\ab[291][1] ) );
  AND U3159 ( .A(A[291]), .B(B[0]), .Z(\ab[291][0] ) );
  AND U3160 ( .A(B[3]), .B(A[290]), .Z(\ab[290][3] ) );
  AND U3161 ( .A(B[2]), .B(A[290]), .Z(\ab[290][2] ) );
  AND U3162 ( .A(B[1]), .B(A[290]), .Z(\ab[290][1] ) );
  AND U3163 ( .A(A[290]), .B(B[0]), .Z(\ab[290][0] ) );
  AND U3164 ( .A(B[3]), .B(A[28]), .Z(\ab[28][3] ) );
  AND U3165 ( .A(B[2]), .B(A[28]), .Z(\ab[28][2] ) );
  AND U3166 ( .A(B[1]), .B(A[28]), .Z(\ab[28][1] ) );
  AND U3167 ( .A(A[28]), .B(B[0]), .Z(\ab[28][0] ) );
  AND U3168 ( .A(B[3]), .B(A[289]), .Z(\ab[289][3] ) );
  AND U3169 ( .A(B[2]), .B(A[289]), .Z(\ab[289][2] ) );
  AND U3170 ( .A(B[1]), .B(A[289]), .Z(\ab[289][1] ) );
  AND U3171 ( .A(A[289]), .B(B[0]), .Z(\ab[289][0] ) );
  AND U3172 ( .A(B[3]), .B(A[288]), .Z(\ab[288][3] ) );
  AND U3173 ( .A(B[2]), .B(A[288]), .Z(\ab[288][2] ) );
  AND U3174 ( .A(B[1]), .B(A[288]), .Z(\ab[288][1] ) );
  AND U3175 ( .A(A[288]), .B(B[0]), .Z(\ab[288][0] ) );
  AND U3176 ( .A(B[3]), .B(A[287]), .Z(\ab[287][3] ) );
  AND U3177 ( .A(B[2]), .B(A[287]), .Z(\ab[287][2] ) );
  AND U3178 ( .A(B[1]), .B(A[287]), .Z(\ab[287][1] ) );
  AND U3179 ( .A(A[287]), .B(B[0]), .Z(\ab[287][0] ) );
  AND U3180 ( .A(B[3]), .B(A[286]), .Z(\ab[286][3] ) );
  AND U3181 ( .A(B[2]), .B(A[286]), .Z(\ab[286][2] ) );
  AND U3182 ( .A(B[1]), .B(A[286]), .Z(\ab[286][1] ) );
  AND U3183 ( .A(A[286]), .B(B[0]), .Z(\ab[286][0] ) );
  AND U3184 ( .A(B[3]), .B(A[285]), .Z(\ab[285][3] ) );
  AND U3185 ( .A(B[2]), .B(A[285]), .Z(\ab[285][2] ) );
  AND U3186 ( .A(B[1]), .B(A[285]), .Z(\ab[285][1] ) );
  AND U3187 ( .A(A[285]), .B(B[0]), .Z(\ab[285][0] ) );
  AND U3188 ( .A(B[3]), .B(A[284]), .Z(\ab[284][3] ) );
  AND U3189 ( .A(B[2]), .B(A[284]), .Z(\ab[284][2] ) );
  AND U3190 ( .A(B[1]), .B(A[284]), .Z(\ab[284][1] ) );
  AND U3191 ( .A(A[284]), .B(B[0]), .Z(\ab[284][0] ) );
  AND U3192 ( .A(B[3]), .B(A[283]), .Z(\ab[283][3] ) );
  AND U3193 ( .A(B[2]), .B(A[283]), .Z(\ab[283][2] ) );
  AND U3194 ( .A(B[1]), .B(A[283]), .Z(\ab[283][1] ) );
  AND U3195 ( .A(A[283]), .B(B[0]), .Z(\ab[283][0] ) );
  AND U3196 ( .A(B[3]), .B(A[282]), .Z(\ab[282][3] ) );
  AND U3197 ( .A(B[2]), .B(A[282]), .Z(\ab[282][2] ) );
  AND U3198 ( .A(B[1]), .B(A[282]), .Z(\ab[282][1] ) );
  AND U3199 ( .A(A[282]), .B(B[0]), .Z(\ab[282][0] ) );
  AND U3200 ( .A(B[3]), .B(A[281]), .Z(\ab[281][3] ) );
  AND U3201 ( .A(B[2]), .B(A[281]), .Z(\ab[281][2] ) );
  AND U3202 ( .A(B[1]), .B(A[281]), .Z(\ab[281][1] ) );
  AND U3203 ( .A(A[281]), .B(B[0]), .Z(\ab[281][0] ) );
  AND U3204 ( .A(B[3]), .B(A[280]), .Z(\ab[280][3] ) );
  AND U3205 ( .A(B[2]), .B(A[280]), .Z(\ab[280][2] ) );
  AND U3206 ( .A(B[1]), .B(A[280]), .Z(\ab[280][1] ) );
  AND U3207 ( .A(A[280]), .B(B[0]), .Z(\ab[280][0] ) );
  AND U3208 ( .A(B[3]), .B(A[27]), .Z(\ab[27][3] ) );
  AND U3209 ( .A(B[2]), .B(A[27]), .Z(\ab[27][2] ) );
  AND U3210 ( .A(B[1]), .B(A[27]), .Z(\ab[27][1] ) );
  AND U3211 ( .A(A[27]), .B(B[0]), .Z(\ab[27][0] ) );
  AND U3212 ( .A(B[3]), .B(A[279]), .Z(\ab[279][3] ) );
  AND U3213 ( .A(B[2]), .B(A[279]), .Z(\ab[279][2] ) );
  AND U3214 ( .A(B[1]), .B(A[279]), .Z(\ab[279][1] ) );
  AND U3215 ( .A(A[279]), .B(B[0]), .Z(\ab[279][0] ) );
  AND U3216 ( .A(B[3]), .B(A[278]), .Z(\ab[278][3] ) );
  AND U3217 ( .A(B[2]), .B(A[278]), .Z(\ab[278][2] ) );
  AND U3218 ( .A(B[1]), .B(A[278]), .Z(\ab[278][1] ) );
  AND U3219 ( .A(A[278]), .B(B[0]), .Z(\ab[278][0] ) );
  AND U3220 ( .A(B[3]), .B(A[277]), .Z(\ab[277][3] ) );
  AND U3221 ( .A(B[2]), .B(A[277]), .Z(\ab[277][2] ) );
  AND U3222 ( .A(B[1]), .B(A[277]), .Z(\ab[277][1] ) );
  AND U3223 ( .A(A[277]), .B(B[0]), .Z(\ab[277][0] ) );
  AND U3224 ( .A(B[3]), .B(A[276]), .Z(\ab[276][3] ) );
  AND U3225 ( .A(B[2]), .B(A[276]), .Z(\ab[276][2] ) );
  AND U3226 ( .A(B[1]), .B(A[276]), .Z(\ab[276][1] ) );
  AND U3227 ( .A(A[276]), .B(B[0]), .Z(\ab[276][0] ) );
  AND U3228 ( .A(B[3]), .B(A[275]), .Z(\ab[275][3] ) );
  AND U3229 ( .A(B[2]), .B(A[275]), .Z(\ab[275][2] ) );
  AND U3230 ( .A(B[1]), .B(A[275]), .Z(\ab[275][1] ) );
  AND U3231 ( .A(A[275]), .B(B[0]), .Z(\ab[275][0] ) );
  AND U3232 ( .A(B[3]), .B(A[274]), .Z(\ab[274][3] ) );
  AND U3233 ( .A(B[2]), .B(A[274]), .Z(\ab[274][2] ) );
  AND U3234 ( .A(B[1]), .B(A[274]), .Z(\ab[274][1] ) );
  AND U3235 ( .A(A[274]), .B(B[0]), .Z(\ab[274][0] ) );
  AND U3236 ( .A(B[3]), .B(A[273]), .Z(\ab[273][3] ) );
  AND U3237 ( .A(B[2]), .B(A[273]), .Z(\ab[273][2] ) );
  AND U3238 ( .A(B[1]), .B(A[273]), .Z(\ab[273][1] ) );
  AND U3239 ( .A(A[273]), .B(B[0]), .Z(\ab[273][0] ) );
  AND U3240 ( .A(B[3]), .B(A[272]), .Z(\ab[272][3] ) );
  AND U3241 ( .A(B[2]), .B(A[272]), .Z(\ab[272][2] ) );
  AND U3242 ( .A(B[1]), .B(A[272]), .Z(\ab[272][1] ) );
  AND U3243 ( .A(A[272]), .B(B[0]), .Z(\ab[272][0] ) );
  AND U3244 ( .A(B[3]), .B(A[271]), .Z(\ab[271][3] ) );
  AND U3245 ( .A(B[2]), .B(A[271]), .Z(\ab[271][2] ) );
  AND U3246 ( .A(B[1]), .B(A[271]), .Z(\ab[271][1] ) );
  AND U3247 ( .A(A[271]), .B(B[0]), .Z(\ab[271][0] ) );
  AND U3248 ( .A(B[3]), .B(A[270]), .Z(\ab[270][3] ) );
  AND U3249 ( .A(B[2]), .B(A[270]), .Z(\ab[270][2] ) );
  AND U3250 ( .A(B[1]), .B(A[270]), .Z(\ab[270][1] ) );
  AND U3251 ( .A(A[270]), .B(B[0]), .Z(\ab[270][0] ) );
  AND U3252 ( .A(B[3]), .B(A[26]), .Z(\ab[26][3] ) );
  AND U3253 ( .A(B[2]), .B(A[26]), .Z(\ab[26][2] ) );
  AND U3254 ( .A(B[1]), .B(A[26]), .Z(\ab[26][1] ) );
  AND U3255 ( .A(A[26]), .B(B[0]), .Z(\ab[26][0] ) );
  AND U3256 ( .A(B[3]), .B(A[269]), .Z(\ab[269][3] ) );
  AND U3257 ( .A(B[2]), .B(A[269]), .Z(\ab[269][2] ) );
  AND U3258 ( .A(B[1]), .B(A[269]), .Z(\ab[269][1] ) );
  AND U3259 ( .A(A[269]), .B(B[0]), .Z(\ab[269][0] ) );
  AND U3260 ( .A(B[3]), .B(A[268]), .Z(\ab[268][3] ) );
  AND U3261 ( .A(B[2]), .B(A[268]), .Z(\ab[268][2] ) );
  AND U3262 ( .A(B[1]), .B(A[268]), .Z(\ab[268][1] ) );
  AND U3263 ( .A(A[268]), .B(B[0]), .Z(\ab[268][0] ) );
  AND U3264 ( .A(B[3]), .B(A[267]), .Z(\ab[267][3] ) );
  AND U3265 ( .A(B[2]), .B(A[267]), .Z(\ab[267][2] ) );
  AND U3266 ( .A(B[1]), .B(A[267]), .Z(\ab[267][1] ) );
  AND U3267 ( .A(A[267]), .B(B[0]), .Z(\ab[267][0] ) );
  AND U3268 ( .A(B[3]), .B(A[266]), .Z(\ab[266][3] ) );
  AND U3269 ( .A(B[2]), .B(A[266]), .Z(\ab[266][2] ) );
  AND U3270 ( .A(B[1]), .B(A[266]), .Z(\ab[266][1] ) );
  AND U3271 ( .A(A[266]), .B(B[0]), .Z(\ab[266][0] ) );
  AND U3272 ( .A(B[3]), .B(A[265]), .Z(\ab[265][3] ) );
  AND U3273 ( .A(B[2]), .B(A[265]), .Z(\ab[265][2] ) );
  AND U3274 ( .A(B[1]), .B(A[265]), .Z(\ab[265][1] ) );
  AND U3275 ( .A(A[265]), .B(B[0]), .Z(\ab[265][0] ) );
  AND U3276 ( .A(B[3]), .B(A[264]), .Z(\ab[264][3] ) );
  AND U3277 ( .A(B[2]), .B(A[264]), .Z(\ab[264][2] ) );
  AND U3278 ( .A(B[1]), .B(A[264]), .Z(\ab[264][1] ) );
  AND U3279 ( .A(A[264]), .B(B[0]), .Z(\ab[264][0] ) );
  AND U3280 ( .A(B[3]), .B(A[263]), .Z(\ab[263][3] ) );
  AND U3281 ( .A(B[2]), .B(A[263]), .Z(\ab[263][2] ) );
  AND U3282 ( .A(B[1]), .B(A[263]), .Z(\ab[263][1] ) );
  AND U3283 ( .A(A[263]), .B(B[0]), .Z(\ab[263][0] ) );
  AND U3284 ( .A(B[3]), .B(A[262]), .Z(\ab[262][3] ) );
  AND U3285 ( .A(B[2]), .B(A[262]), .Z(\ab[262][2] ) );
  AND U3286 ( .A(B[1]), .B(A[262]), .Z(\ab[262][1] ) );
  AND U3287 ( .A(A[262]), .B(B[0]), .Z(\ab[262][0] ) );
  AND U3288 ( .A(B[3]), .B(A[261]), .Z(\ab[261][3] ) );
  AND U3289 ( .A(B[2]), .B(A[261]), .Z(\ab[261][2] ) );
  AND U3290 ( .A(B[1]), .B(A[261]), .Z(\ab[261][1] ) );
  AND U3291 ( .A(A[261]), .B(B[0]), .Z(\ab[261][0] ) );
  AND U3292 ( .A(B[3]), .B(A[260]), .Z(\ab[260][3] ) );
  AND U3293 ( .A(B[2]), .B(A[260]), .Z(\ab[260][2] ) );
  AND U3294 ( .A(B[1]), .B(A[260]), .Z(\ab[260][1] ) );
  AND U3295 ( .A(A[260]), .B(B[0]), .Z(\ab[260][0] ) );
  AND U3296 ( .A(B[3]), .B(A[25]), .Z(\ab[25][3] ) );
  AND U3297 ( .A(B[2]), .B(A[25]), .Z(\ab[25][2] ) );
  AND U3298 ( .A(B[1]), .B(A[25]), .Z(\ab[25][1] ) );
  AND U3299 ( .A(A[25]), .B(B[0]), .Z(\ab[25][0] ) );
  AND U3300 ( .A(B[3]), .B(A[259]), .Z(\ab[259][3] ) );
  AND U3301 ( .A(B[2]), .B(A[259]), .Z(\ab[259][2] ) );
  AND U3302 ( .A(B[1]), .B(A[259]), .Z(\ab[259][1] ) );
  AND U3303 ( .A(A[259]), .B(B[0]), .Z(\ab[259][0] ) );
  AND U3304 ( .A(B[3]), .B(A[258]), .Z(\ab[258][3] ) );
  AND U3305 ( .A(B[2]), .B(A[258]), .Z(\ab[258][2] ) );
  AND U3306 ( .A(B[1]), .B(A[258]), .Z(\ab[258][1] ) );
  AND U3307 ( .A(A[258]), .B(B[0]), .Z(\ab[258][0] ) );
  AND U3308 ( .A(B[3]), .B(A[257]), .Z(\ab[257][3] ) );
  AND U3309 ( .A(B[2]), .B(A[257]), .Z(\ab[257][2] ) );
  AND U3310 ( .A(B[1]), .B(A[257]), .Z(\ab[257][1] ) );
  AND U3311 ( .A(A[257]), .B(B[0]), .Z(\ab[257][0] ) );
  AND U3312 ( .A(B[3]), .B(A[256]), .Z(\ab[256][3] ) );
  AND U3313 ( .A(B[2]), .B(A[256]), .Z(\ab[256][2] ) );
  AND U3314 ( .A(B[1]), .B(A[256]), .Z(\ab[256][1] ) );
  AND U3315 ( .A(A[256]), .B(B[0]), .Z(\ab[256][0] ) );
  AND U3316 ( .A(B[3]), .B(A[255]), .Z(\ab[255][3] ) );
  AND U3317 ( .A(B[2]), .B(A[255]), .Z(\ab[255][2] ) );
  AND U3318 ( .A(B[1]), .B(A[255]), .Z(\ab[255][1] ) );
  AND U3319 ( .A(A[255]), .B(B[0]), .Z(\ab[255][0] ) );
  AND U3320 ( .A(B[3]), .B(A[254]), .Z(\ab[254][3] ) );
  AND U3321 ( .A(B[2]), .B(A[254]), .Z(\ab[254][2] ) );
  AND U3322 ( .A(B[1]), .B(A[254]), .Z(\ab[254][1] ) );
  AND U3323 ( .A(A[254]), .B(B[0]), .Z(\ab[254][0] ) );
  AND U3324 ( .A(B[3]), .B(A[253]), .Z(\ab[253][3] ) );
  AND U3325 ( .A(B[2]), .B(A[253]), .Z(\ab[253][2] ) );
  AND U3326 ( .A(B[1]), .B(A[253]), .Z(\ab[253][1] ) );
  AND U3327 ( .A(A[253]), .B(B[0]), .Z(\ab[253][0] ) );
  AND U3328 ( .A(B[3]), .B(A[252]), .Z(\ab[252][3] ) );
  AND U3329 ( .A(B[2]), .B(A[252]), .Z(\ab[252][2] ) );
  AND U3330 ( .A(B[1]), .B(A[252]), .Z(\ab[252][1] ) );
  AND U3331 ( .A(A[252]), .B(B[0]), .Z(\ab[252][0] ) );
  AND U3332 ( .A(B[3]), .B(A[251]), .Z(\ab[251][3] ) );
  AND U3333 ( .A(B[2]), .B(A[251]), .Z(\ab[251][2] ) );
  AND U3334 ( .A(B[1]), .B(A[251]), .Z(\ab[251][1] ) );
  AND U3335 ( .A(A[251]), .B(B[0]), .Z(\ab[251][0] ) );
  AND U3336 ( .A(B[3]), .B(A[250]), .Z(\ab[250][3] ) );
  AND U3337 ( .A(B[2]), .B(A[250]), .Z(\ab[250][2] ) );
  AND U3338 ( .A(B[1]), .B(A[250]), .Z(\ab[250][1] ) );
  AND U3339 ( .A(A[250]), .B(B[0]), .Z(\ab[250][0] ) );
  AND U3340 ( .A(B[3]), .B(A[24]), .Z(\ab[24][3] ) );
  AND U3341 ( .A(B[2]), .B(A[24]), .Z(\ab[24][2] ) );
  AND U3342 ( .A(B[1]), .B(A[24]), .Z(\ab[24][1] ) );
  AND U3343 ( .A(A[24]), .B(B[0]), .Z(\ab[24][0] ) );
  AND U3344 ( .A(B[3]), .B(A[249]), .Z(\ab[249][3] ) );
  AND U3345 ( .A(B[2]), .B(A[249]), .Z(\ab[249][2] ) );
  AND U3346 ( .A(B[1]), .B(A[249]), .Z(\ab[249][1] ) );
  AND U3347 ( .A(A[249]), .B(B[0]), .Z(\ab[249][0] ) );
  AND U3348 ( .A(B[3]), .B(A[248]), .Z(\ab[248][3] ) );
  AND U3349 ( .A(B[2]), .B(A[248]), .Z(\ab[248][2] ) );
  AND U3350 ( .A(B[1]), .B(A[248]), .Z(\ab[248][1] ) );
  AND U3351 ( .A(A[248]), .B(B[0]), .Z(\ab[248][0] ) );
  AND U3352 ( .A(B[3]), .B(A[247]), .Z(\ab[247][3] ) );
  AND U3353 ( .A(B[2]), .B(A[247]), .Z(\ab[247][2] ) );
  AND U3354 ( .A(B[1]), .B(A[247]), .Z(\ab[247][1] ) );
  AND U3355 ( .A(A[247]), .B(B[0]), .Z(\ab[247][0] ) );
  AND U3356 ( .A(B[3]), .B(A[246]), .Z(\ab[246][3] ) );
  AND U3357 ( .A(B[2]), .B(A[246]), .Z(\ab[246][2] ) );
  AND U3358 ( .A(B[1]), .B(A[246]), .Z(\ab[246][1] ) );
  AND U3359 ( .A(A[246]), .B(B[0]), .Z(\ab[246][0] ) );
  AND U3360 ( .A(B[3]), .B(A[245]), .Z(\ab[245][3] ) );
  AND U3361 ( .A(B[2]), .B(A[245]), .Z(\ab[245][2] ) );
  AND U3362 ( .A(B[1]), .B(A[245]), .Z(\ab[245][1] ) );
  AND U3363 ( .A(A[245]), .B(B[0]), .Z(\ab[245][0] ) );
  AND U3364 ( .A(B[3]), .B(A[244]), .Z(\ab[244][3] ) );
  AND U3365 ( .A(B[2]), .B(A[244]), .Z(\ab[244][2] ) );
  AND U3366 ( .A(B[1]), .B(A[244]), .Z(\ab[244][1] ) );
  AND U3367 ( .A(A[244]), .B(B[0]), .Z(\ab[244][0] ) );
  AND U3368 ( .A(B[3]), .B(A[243]), .Z(\ab[243][3] ) );
  AND U3369 ( .A(B[2]), .B(A[243]), .Z(\ab[243][2] ) );
  AND U3370 ( .A(B[1]), .B(A[243]), .Z(\ab[243][1] ) );
  AND U3371 ( .A(A[243]), .B(B[0]), .Z(\ab[243][0] ) );
  AND U3372 ( .A(B[3]), .B(A[242]), .Z(\ab[242][3] ) );
  AND U3373 ( .A(B[2]), .B(A[242]), .Z(\ab[242][2] ) );
  AND U3374 ( .A(B[1]), .B(A[242]), .Z(\ab[242][1] ) );
  AND U3375 ( .A(A[242]), .B(B[0]), .Z(\ab[242][0] ) );
  AND U3376 ( .A(B[3]), .B(A[241]), .Z(\ab[241][3] ) );
  AND U3377 ( .A(B[2]), .B(A[241]), .Z(\ab[241][2] ) );
  AND U3378 ( .A(B[1]), .B(A[241]), .Z(\ab[241][1] ) );
  AND U3379 ( .A(A[241]), .B(B[0]), .Z(\ab[241][0] ) );
  AND U3380 ( .A(B[3]), .B(A[240]), .Z(\ab[240][3] ) );
  AND U3381 ( .A(B[2]), .B(A[240]), .Z(\ab[240][2] ) );
  AND U3382 ( .A(B[1]), .B(A[240]), .Z(\ab[240][1] ) );
  AND U3383 ( .A(A[240]), .B(B[0]), .Z(\ab[240][0] ) );
  AND U3384 ( .A(B[3]), .B(A[23]), .Z(\ab[23][3] ) );
  AND U3385 ( .A(B[2]), .B(A[23]), .Z(\ab[23][2] ) );
  AND U3386 ( .A(B[1]), .B(A[23]), .Z(\ab[23][1] ) );
  AND U3387 ( .A(A[23]), .B(B[0]), .Z(\ab[23][0] ) );
  AND U3388 ( .A(B[3]), .B(A[239]), .Z(\ab[239][3] ) );
  AND U3389 ( .A(B[2]), .B(A[239]), .Z(\ab[239][2] ) );
  AND U3390 ( .A(B[1]), .B(A[239]), .Z(\ab[239][1] ) );
  AND U3391 ( .A(A[239]), .B(B[0]), .Z(\ab[239][0] ) );
  AND U3392 ( .A(B[3]), .B(A[238]), .Z(\ab[238][3] ) );
  AND U3393 ( .A(B[2]), .B(A[238]), .Z(\ab[238][2] ) );
  AND U3394 ( .A(B[1]), .B(A[238]), .Z(\ab[238][1] ) );
  AND U3395 ( .A(A[238]), .B(B[0]), .Z(\ab[238][0] ) );
  AND U3396 ( .A(B[3]), .B(A[237]), .Z(\ab[237][3] ) );
  AND U3397 ( .A(B[2]), .B(A[237]), .Z(\ab[237][2] ) );
  AND U3398 ( .A(B[1]), .B(A[237]), .Z(\ab[237][1] ) );
  AND U3399 ( .A(A[237]), .B(B[0]), .Z(\ab[237][0] ) );
  AND U3400 ( .A(B[3]), .B(A[236]), .Z(\ab[236][3] ) );
  AND U3401 ( .A(B[2]), .B(A[236]), .Z(\ab[236][2] ) );
  AND U3402 ( .A(B[1]), .B(A[236]), .Z(\ab[236][1] ) );
  AND U3403 ( .A(A[236]), .B(B[0]), .Z(\ab[236][0] ) );
  AND U3404 ( .A(B[3]), .B(A[235]), .Z(\ab[235][3] ) );
  AND U3405 ( .A(B[2]), .B(A[235]), .Z(\ab[235][2] ) );
  AND U3406 ( .A(B[1]), .B(A[235]), .Z(\ab[235][1] ) );
  AND U3407 ( .A(A[235]), .B(B[0]), .Z(\ab[235][0] ) );
  AND U3408 ( .A(B[3]), .B(A[234]), .Z(\ab[234][3] ) );
  AND U3409 ( .A(B[2]), .B(A[234]), .Z(\ab[234][2] ) );
  AND U3410 ( .A(B[1]), .B(A[234]), .Z(\ab[234][1] ) );
  AND U3411 ( .A(A[234]), .B(B[0]), .Z(\ab[234][0] ) );
  AND U3412 ( .A(B[3]), .B(A[233]), .Z(\ab[233][3] ) );
  AND U3413 ( .A(B[2]), .B(A[233]), .Z(\ab[233][2] ) );
  AND U3414 ( .A(B[1]), .B(A[233]), .Z(\ab[233][1] ) );
  AND U3415 ( .A(A[233]), .B(B[0]), .Z(\ab[233][0] ) );
  AND U3416 ( .A(B[3]), .B(A[232]), .Z(\ab[232][3] ) );
  AND U3417 ( .A(B[2]), .B(A[232]), .Z(\ab[232][2] ) );
  AND U3418 ( .A(B[1]), .B(A[232]), .Z(\ab[232][1] ) );
  AND U3419 ( .A(A[232]), .B(B[0]), .Z(\ab[232][0] ) );
  AND U3420 ( .A(B[3]), .B(A[231]), .Z(\ab[231][3] ) );
  AND U3421 ( .A(B[2]), .B(A[231]), .Z(\ab[231][2] ) );
  AND U3422 ( .A(B[1]), .B(A[231]), .Z(\ab[231][1] ) );
  AND U3423 ( .A(A[231]), .B(B[0]), .Z(\ab[231][0] ) );
  AND U3424 ( .A(B[3]), .B(A[230]), .Z(\ab[230][3] ) );
  AND U3425 ( .A(B[2]), .B(A[230]), .Z(\ab[230][2] ) );
  AND U3426 ( .A(B[1]), .B(A[230]), .Z(\ab[230][1] ) );
  AND U3427 ( .A(A[230]), .B(B[0]), .Z(\ab[230][0] ) );
  AND U3428 ( .A(B[3]), .B(A[22]), .Z(\ab[22][3] ) );
  AND U3429 ( .A(B[2]), .B(A[22]), .Z(\ab[22][2] ) );
  AND U3430 ( .A(B[1]), .B(A[22]), .Z(\ab[22][1] ) );
  AND U3431 ( .A(A[22]), .B(B[0]), .Z(\ab[22][0] ) );
  AND U3432 ( .A(B[3]), .B(A[229]), .Z(\ab[229][3] ) );
  AND U3433 ( .A(B[2]), .B(A[229]), .Z(\ab[229][2] ) );
  AND U3434 ( .A(B[1]), .B(A[229]), .Z(\ab[229][1] ) );
  AND U3435 ( .A(A[229]), .B(B[0]), .Z(\ab[229][0] ) );
  AND U3436 ( .A(B[3]), .B(A[228]), .Z(\ab[228][3] ) );
  AND U3437 ( .A(B[2]), .B(A[228]), .Z(\ab[228][2] ) );
  AND U3438 ( .A(B[1]), .B(A[228]), .Z(\ab[228][1] ) );
  AND U3439 ( .A(A[228]), .B(B[0]), .Z(\ab[228][0] ) );
  AND U3440 ( .A(B[3]), .B(A[227]), .Z(\ab[227][3] ) );
  AND U3441 ( .A(B[2]), .B(A[227]), .Z(\ab[227][2] ) );
  AND U3442 ( .A(B[1]), .B(A[227]), .Z(\ab[227][1] ) );
  AND U3443 ( .A(A[227]), .B(B[0]), .Z(\ab[227][0] ) );
  AND U3444 ( .A(B[3]), .B(A[226]), .Z(\ab[226][3] ) );
  AND U3445 ( .A(B[2]), .B(A[226]), .Z(\ab[226][2] ) );
  AND U3446 ( .A(B[1]), .B(A[226]), .Z(\ab[226][1] ) );
  AND U3447 ( .A(A[226]), .B(B[0]), .Z(\ab[226][0] ) );
  AND U3448 ( .A(B[3]), .B(A[225]), .Z(\ab[225][3] ) );
  AND U3449 ( .A(B[2]), .B(A[225]), .Z(\ab[225][2] ) );
  AND U3450 ( .A(B[1]), .B(A[225]), .Z(\ab[225][1] ) );
  AND U3451 ( .A(A[225]), .B(B[0]), .Z(\ab[225][0] ) );
  AND U3452 ( .A(B[3]), .B(A[224]), .Z(\ab[224][3] ) );
  AND U3453 ( .A(B[2]), .B(A[224]), .Z(\ab[224][2] ) );
  AND U3454 ( .A(B[1]), .B(A[224]), .Z(\ab[224][1] ) );
  AND U3455 ( .A(A[224]), .B(B[0]), .Z(\ab[224][0] ) );
  AND U3456 ( .A(B[3]), .B(A[223]), .Z(\ab[223][3] ) );
  AND U3457 ( .A(B[2]), .B(A[223]), .Z(\ab[223][2] ) );
  AND U3458 ( .A(B[1]), .B(A[223]), .Z(\ab[223][1] ) );
  AND U3459 ( .A(A[223]), .B(B[0]), .Z(\ab[223][0] ) );
  AND U3460 ( .A(B[3]), .B(A[222]), .Z(\ab[222][3] ) );
  AND U3461 ( .A(B[2]), .B(A[222]), .Z(\ab[222][2] ) );
  AND U3462 ( .A(B[1]), .B(A[222]), .Z(\ab[222][1] ) );
  AND U3463 ( .A(A[222]), .B(B[0]), .Z(\ab[222][0] ) );
  AND U3464 ( .A(B[3]), .B(A[221]), .Z(\ab[221][3] ) );
  AND U3465 ( .A(B[2]), .B(A[221]), .Z(\ab[221][2] ) );
  AND U3466 ( .A(B[1]), .B(A[221]), .Z(\ab[221][1] ) );
  AND U3467 ( .A(A[221]), .B(B[0]), .Z(\ab[221][0] ) );
  AND U3468 ( .A(B[3]), .B(A[220]), .Z(\ab[220][3] ) );
  AND U3469 ( .A(B[2]), .B(A[220]), .Z(\ab[220][2] ) );
  AND U3470 ( .A(B[1]), .B(A[220]), .Z(\ab[220][1] ) );
  AND U3471 ( .A(A[220]), .B(B[0]), .Z(\ab[220][0] ) );
  AND U3472 ( .A(B[3]), .B(A[21]), .Z(\ab[21][3] ) );
  AND U3473 ( .A(B[2]), .B(A[21]), .Z(\ab[21][2] ) );
  AND U3474 ( .A(B[1]), .B(A[21]), .Z(\ab[21][1] ) );
  AND U3475 ( .A(A[21]), .B(B[0]), .Z(\ab[21][0] ) );
  AND U3476 ( .A(B[3]), .B(A[219]), .Z(\ab[219][3] ) );
  AND U3477 ( .A(B[2]), .B(A[219]), .Z(\ab[219][2] ) );
  AND U3478 ( .A(B[1]), .B(A[219]), .Z(\ab[219][1] ) );
  AND U3479 ( .A(A[219]), .B(B[0]), .Z(\ab[219][0] ) );
  AND U3480 ( .A(B[3]), .B(A[218]), .Z(\ab[218][3] ) );
  AND U3481 ( .A(B[2]), .B(A[218]), .Z(\ab[218][2] ) );
  AND U3482 ( .A(B[1]), .B(A[218]), .Z(\ab[218][1] ) );
  AND U3483 ( .A(A[218]), .B(B[0]), .Z(\ab[218][0] ) );
  AND U3484 ( .A(B[3]), .B(A[217]), .Z(\ab[217][3] ) );
  AND U3485 ( .A(B[2]), .B(A[217]), .Z(\ab[217][2] ) );
  AND U3486 ( .A(B[1]), .B(A[217]), .Z(\ab[217][1] ) );
  AND U3487 ( .A(A[217]), .B(B[0]), .Z(\ab[217][0] ) );
  AND U3488 ( .A(B[3]), .B(A[216]), .Z(\ab[216][3] ) );
  AND U3489 ( .A(B[2]), .B(A[216]), .Z(\ab[216][2] ) );
  AND U3490 ( .A(B[1]), .B(A[216]), .Z(\ab[216][1] ) );
  AND U3491 ( .A(A[216]), .B(B[0]), .Z(\ab[216][0] ) );
  AND U3492 ( .A(B[3]), .B(A[215]), .Z(\ab[215][3] ) );
  AND U3493 ( .A(B[2]), .B(A[215]), .Z(\ab[215][2] ) );
  AND U3494 ( .A(B[1]), .B(A[215]), .Z(\ab[215][1] ) );
  AND U3495 ( .A(A[215]), .B(B[0]), .Z(\ab[215][0] ) );
  AND U3496 ( .A(B[3]), .B(A[214]), .Z(\ab[214][3] ) );
  AND U3497 ( .A(B[2]), .B(A[214]), .Z(\ab[214][2] ) );
  AND U3498 ( .A(B[1]), .B(A[214]), .Z(\ab[214][1] ) );
  AND U3499 ( .A(A[214]), .B(B[0]), .Z(\ab[214][0] ) );
  AND U3500 ( .A(B[3]), .B(A[213]), .Z(\ab[213][3] ) );
  AND U3501 ( .A(B[2]), .B(A[213]), .Z(\ab[213][2] ) );
  AND U3502 ( .A(B[1]), .B(A[213]), .Z(\ab[213][1] ) );
  AND U3503 ( .A(A[213]), .B(B[0]), .Z(\ab[213][0] ) );
  AND U3504 ( .A(B[3]), .B(A[212]), .Z(\ab[212][3] ) );
  AND U3505 ( .A(B[2]), .B(A[212]), .Z(\ab[212][2] ) );
  AND U3506 ( .A(B[1]), .B(A[212]), .Z(\ab[212][1] ) );
  AND U3507 ( .A(A[212]), .B(B[0]), .Z(\ab[212][0] ) );
  AND U3508 ( .A(B[3]), .B(A[211]), .Z(\ab[211][3] ) );
  AND U3509 ( .A(B[2]), .B(A[211]), .Z(\ab[211][2] ) );
  AND U3510 ( .A(B[1]), .B(A[211]), .Z(\ab[211][1] ) );
  AND U3511 ( .A(A[211]), .B(B[0]), .Z(\ab[211][0] ) );
  AND U3512 ( .A(B[3]), .B(A[210]), .Z(\ab[210][3] ) );
  AND U3513 ( .A(B[2]), .B(A[210]), .Z(\ab[210][2] ) );
  AND U3514 ( .A(B[1]), .B(A[210]), .Z(\ab[210][1] ) );
  AND U3515 ( .A(A[210]), .B(B[0]), .Z(\ab[210][0] ) );
  AND U3516 ( .A(B[3]), .B(A[20]), .Z(\ab[20][3] ) );
  AND U3517 ( .A(B[2]), .B(A[20]), .Z(\ab[20][2] ) );
  AND U3518 ( .A(B[1]), .B(A[20]), .Z(\ab[20][1] ) );
  AND U3519 ( .A(A[20]), .B(B[0]), .Z(\ab[20][0] ) );
  AND U3520 ( .A(B[3]), .B(A[209]), .Z(\ab[209][3] ) );
  AND U3521 ( .A(B[2]), .B(A[209]), .Z(\ab[209][2] ) );
  AND U3522 ( .A(B[1]), .B(A[209]), .Z(\ab[209][1] ) );
  AND U3523 ( .A(A[209]), .B(B[0]), .Z(\ab[209][0] ) );
  AND U3524 ( .A(B[3]), .B(A[208]), .Z(\ab[208][3] ) );
  AND U3525 ( .A(B[2]), .B(A[208]), .Z(\ab[208][2] ) );
  AND U3526 ( .A(B[1]), .B(A[208]), .Z(\ab[208][1] ) );
  AND U3527 ( .A(A[208]), .B(B[0]), .Z(\ab[208][0] ) );
  AND U3528 ( .A(B[3]), .B(A[207]), .Z(\ab[207][3] ) );
  AND U3529 ( .A(B[2]), .B(A[207]), .Z(\ab[207][2] ) );
  AND U3530 ( .A(B[1]), .B(A[207]), .Z(\ab[207][1] ) );
  AND U3531 ( .A(A[207]), .B(B[0]), .Z(\ab[207][0] ) );
  AND U3532 ( .A(B[3]), .B(A[206]), .Z(\ab[206][3] ) );
  AND U3533 ( .A(B[2]), .B(A[206]), .Z(\ab[206][2] ) );
  AND U3534 ( .A(B[1]), .B(A[206]), .Z(\ab[206][1] ) );
  AND U3535 ( .A(A[206]), .B(B[0]), .Z(\ab[206][0] ) );
  AND U3536 ( .A(B[3]), .B(A[205]), .Z(\ab[205][3] ) );
  AND U3537 ( .A(B[2]), .B(A[205]), .Z(\ab[205][2] ) );
  AND U3538 ( .A(B[1]), .B(A[205]), .Z(\ab[205][1] ) );
  AND U3539 ( .A(A[205]), .B(B[0]), .Z(\ab[205][0] ) );
  AND U3540 ( .A(B[3]), .B(A[204]), .Z(\ab[204][3] ) );
  AND U3541 ( .A(B[2]), .B(A[204]), .Z(\ab[204][2] ) );
  AND U3542 ( .A(B[1]), .B(A[204]), .Z(\ab[204][1] ) );
  AND U3543 ( .A(A[204]), .B(B[0]), .Z(\ab[204][0] ) );
  AND U3544 ( .A(B[3]), .B(A[203]), .Z(\ab[203][3] ) );
  AND U3545 ( .A(B[2]), .B(A[203]), .Z(\ab[203][2] ) );
  AND U3546 ( .A(B[1]), .B(A[203]), .Z(\ab[203][1] ) );
  AND U3547 ( .A(A[203]), .B(B[0]), .Z(\ab[203][0] ) );
  AND U3548 ( .A(B[3]), .B(A[202]), .Z(\ab[202][3] ) );
  AND U3549 ( .A(B[2]), .B(A[202]), .Z(\ab[202][2] ) );
  AND U3550 ( .A(B[1]), .B(A[202]), .Z(\ab[202][1] ) );
  AND U3551 ( .A(A[202]), .B(B[0]), .Z(\ab[202][0] ) );
  AND U3552 ( .A(B[3]), .B(A[201]), .Z(\ab[201][3] ) );
  AND U3553 ( .A(B[2]), .B(A[201]), .Z(\ab[201][2] ) );
  AND U3554 ( .A(B[1]), .B(A[201]), .Z(\ab[201][1] ) );
  AND U3555 ( .A(A[201]), .B(B[0]), .Z(\ab[201][0] ) );
  AND U3556 ( .A(B[3]), .B(A[200]), .Z(\ab[200][3] ) );
  AND U3557 ( .A(B[2]), .B(A[200]), .Z(\ab[200][2] ) );
  AND U3558 ( .A(B[1]), .B(A[200]), .Z(\ab[200][1] ) );
  AND U3559 ( .A(A[200]), .B(B[0]), .Z(\ab[200][0] ) );
  AND U3560 ( .A(B[3]), .B(A[1]), .Z(\ab[1][3] ) );
  AND U3561 ( .A(B[2]), .B(A[1]), .Z(\ab[1][2] ) );
  AND U3562 ( .A(B[1]), .B(A[1]), .Z(\ab[1][1] ) );
  AND U3563 ( .A(A[1]), .B(B[0]), .Z(\ab[1][0] ) );
  AND U3564 ( .A(B[3]), .B(A[19]), .Z(\ab[19][3] ) );
  AND U3565 ( .A(B[2]), .B(A[19]), .Z(\ab[19][2] ) );
  AND U3566 ( .A(B[1]), .B(A[19]), .Z(\ab[19][1] ) );
  AND U3567 ( .A(A[19]), .B(B[0]), .Z(\ab[19][0] ) );
  AND U3568 ( .A(B[3]), .B(A[199]), .Z(\ab[199][3] ) );
  AND U3569 ( .A(B[2]), .B(A[199]), .Z(\ab[199][2] ) );
  AND U3570 ( .A(B[1]), .B(A[199]), .Z(\ab[199][1] ) );
  AND U3571 ( .A(A[199]), .B(B[0]), .Z(\ab[199][0] ) );
  AND U3572 ( .A(B[3]), .B(A[198]), .Z(\ab[198][3] ) );
  AND U3573 ( .A(B[2]), .B(A[198]), .Z(\ab[198][2] ) );
  AND U3574 ( .A(B[1]), .B(A[198]), .Z(\ab[198][1] ) );
  AND U3575 ( .A(A[198]), .B(B[0]), .Z(\ab[198][0] ) );
  AND U3576 ( .A(B[3]), .B(A[197]), .Z(\ab[197][3] ) );
  AND U3577 ( .A(B[2]), .B(A[197]), .Z(\ab[197][2] ) );
  AND U3578 ( .A(B[1]), .B(A[197]), .Z(\ab[197][1] ) );
  AND U3579 ( .A(A[197]), .B(B[0]), .Z(\ab[197][0] ) );
  AND U3580 ( .A(B[3]), .B(A[196]), .Z(\ab[196][3] ) );
  AND U3581 ( .A(B[2]), .B(A[196]), .Z(\ab[196][2] ) );
  AND U3582 ( .A(B[1]), .B(A[196]), .Z(\ab[196][1] ) );
  AND U3583 ( .A(A[196]), .B(B[0]), .Z(\ab[196][0] ) );
  AND U3584 ( .A(B[3]), .B(A[195]), .Z(\ab[195][3] ) );
  AND U3585 ( .A(B[2]), .B(A[195]), .Z(\ab[195][2] ) );
  AND U3586 ( .A(B[1]), .B(A[195]), .Z(\ab[195][1] ) );
  AND U3587 ( .A(A[195]), .B(B[0]), .Z(\ab[195][0] ) );
  AND U3588 ( .A(B[3]), .B(A[194]), .Z(\ab[194][3] ) );
  AND U3589 ( .A(B[2]), .B(A[194]), .Z(\ab[194][2] ) );
  AND U3590 ( .A(B[1]), .B(A[194]), .Z(\ab[194][1] ) );
  AND U3591 ( .A(A[194]), .B(B[0]), .Z(\ab[194][0] ) );
  AND U3592 ( .A(B[3]), .B(A[193]), .Z(\ab[193][3] ) );
  AND U3593 ( .A(B[2]), .B(A[193]), .Z(\ab[193][2] ) );
  AND U3594 ( .A(B[1]), .B(A[193]), .Z(\ab[193][1] ) );
  AND U3595 ( .A(A[193]), .B(B[0]), .Z(\ab[193][0] ) );
  AND U3596 ( .A(B[3]), .B(A[192]), .Z(\ab[192][3] ) );
  AND U3597 ( .A(B[2]), .B(A[192]), .Z(\ab[192][2] ) );
  AND U3598 ( .A(B[1]), .B(A[192]), .Z(\ab[192][1] ) );
  AND U3599 ( .A(A[192]), .B(B[0]), .Z(\ab[192][0] ) );
  AND U3600 ( .A(B[3]), .B(A[191]), .Z(\ab[191][3] ) );
  AND U3601 ( .A(B[2]), .B(A[191]), .Z(\ab[191][2] ) );
  AND U3602 ( .A(B[1]), .B(A[191]), .Z(\ab[191][1] ) );
  AND U3603 ( .A(A[191]), .B(B[0]), .Z(\ab[191][0] ) );
  AND U3604 ( .A(B[3]), .B(A[190]), .Z(\ab[190][3] ) );
  AND U3605 ( .A(B[2]), .B(A[190]), .Z(\ab[190][2] ) );
  AND U3606 ( .A(B[1]), .B(A[190]), .Z(\ab[190][1] ) );
  AND U3607 ( .A(A[190]), .B(B[0]), .Z(\ab[190][0] ) );
  AND U3608 ( .A(B[3]), .B(A[18]), .Z(\ab[18][3] ) );
  AND U3609 ( .A(B[2]), .B(A[18]), .Z(\ab[18][2] ) );
  AND U3610 ( .A(B[1]), .B(A[18]), .Z(\ab[18][1] ) );
  AND U3611 ( .A(A[18]), .B(B[0]), .Z(\ab[18][0] ) );
  AND U3612 ( .A(B[3]), .B(A[189]), .Z(\ab[189][3] ) );
  AND U3613 ( .A(B[2]), .B(A[189]), .Z(\ab[189][2] ) );
  AND U3614 ( .A(B[1]), .B(A[189]), .Z(\ab[189][1] ) );
  AND U3615 ( .A(A[189]), .B(B[0]), .Z(\ab[189][0] ) );
  AND U3616 ( .A(B[3]), .B(A[188]), .Z(\ab[188][3] ) );
  AND U3617 ( .A(B[2]), .B(A[188]), .Z(\ab[188][2] ) );
  AND U3618 ( .A(B[1]), .B(A[188]), .Z(\ab[188][1] ) );
  AND U3619 ( .A(A[188]), .B(B[0]), .Z(\ab[188][0] ) );
  AND U3620 ( .A(B[3]), .B(A[187]), .Z(\ab[187][3] ) );
  AND U3621 ( .A(B[2]), .B(A[187]), .Z(\ab[187][2] ) );
  AND U3622 ( .A(B[1]), .B(A[187]), .Z(\ab[187][1] ) );
  AND U3623 ( .A(A[187]), .B(B[0]), .Z(\ab[187][0] ) );
  AND U3624 ( .A(B[3]), .B(A[186]), .Z(\ab[186][3] ) );
  AND U3625 ( .A(B[2]), .B(A[186]), .Z(\ab[186][2] ) );
  AND U3626 ( .A(B[1]), .B(A[186]), .Z(\ab[186][1] ) );
  AND U3627 ( .A(A[186]), .B(B[0]), .Z(\ab[186][0] ) );
  AND U3628 ( .A(B[3]), .B(A[185]), .Z(\ab[185][3] ) );
  AND U3629 ( .A(B[2]), .B(A[185]), .Z(\ab[185][2] ) );
  AND U3630 ( .A(B[1]), .B(A[185]), .Z(\ab[185][1] ) );
  AND U3631 ( .A(A[185]), .B(B[0]), .Z(\ab[185][0] ) );
  AND U3632 ( .A(B[3]), .B(A[184]), .Z(\ab[184][3] ) );
  AND U3633 ( .A(B[2]), .B(A[184]), .Z(\ab[184][2] ) );
  AND U3634 ( .A(B[1]), .B(A[184]), .Z(\ab[184][1] ) );
  AND U3635 ( .A(A[184]), .B(B[0]), .Z(\ab[184][0] ) );
  AND U3636 ( .A(B[3]), .B(A[183]), .Z(\ab[183][3] ) );
  AND U3637 ( .A(B[2]), .B(A[183]), .Z(\ab[183][2] ) );
  AND U3638 ( .A(B[1]), .B(A[183]), .Z(\ab[183][1] ) );
  AND U3639 ( .A(A[183]), .B(B[0]), .Z(\ab[183][0] ) );
  AND U3640 ( .A(B[3]), .B(A[182]), .Z(\ab[182][3] ) );
  AND U3641 ( .A(B[2]), .B(A[182]), .Z(\ab[182][2] ) );
  AND U3642 ( .A(B[1]), .B(A[182]), .Z(\ab[182][1] ) );
  AND U3643 ( .A(A[182]), .B(B[0]), .Z(\ab[182][0] ) );
  AND U3644 ( .A(B[3]), .B(A[181]), .Z(\ab[181][3] ) );
  AND U3645 ( .A(B[2]), .B(A[181]), .Z(\ab[181][2] ) );
  AND U3646 ( .A(B[1]), .B(A[181]), .Z(\ab[181][1] ) );
  AND U3647 ( .A(A[181]), .B(B[0]), .Z(\ab[181][0] ) );
  AND U3648 ( .A(B[3]), .B(A[180]), .Z(\ab[180][3] ) );
  AND U3649 ( .A(B[2]), .B(A[180]), .Z(\ab[180][2] ) );
  AND U3650 ( .A(B[1]), .B(A[180]), .Z(\ab[180][1] ) );
  AND U3651 ( .A(A[180]), .B(B[0]), .Z(\ab[180][0] ) );
  AND U3652 ( .A(B[3]), .B(A[17]), .Z(\ab[17][3] ) );
  AND U3653 ( .A(B[2]), .B(A[17]), .Z(\ab[17][2] ) );
  AND U3654 ( .A(B[1]), .B(A[17]), .Z(\ab[17][1] ) );
  AND U3655 ( .A(A[17]), .B(B[0]), .Z(\ab[17][0] ) );
  AND U3656 ( .A(B[3]), .B(A[179]), .Z(\ab[179][3] ) );
  AND U3657 ( .A(B[2]), .B(A[179]), .Z(\ab[179][2] ) );
  AND U3658 ( .A(B[1]), .B(A[179]), .Z(\ab[179][1] ) );
  AND U3659 ( .A(A[179]), .B(B[0]), .Z(\ab[179][0] ) );
  AND U3660 ( .A(B[3]), .B(A[178]), .Z(\ab[178][3] ) );
  AND U3661 ( .A(B[2]), .B(A[178]), .Z(\ab[178][2] ) );
  AND U3662 ( .A(B[1]), .B(A[178]), .Z(\ab[178][1] ) );
  AND U3663 ( .A(A[178]), .B(B[0]), .Z(\ab[178][0] ) );
  AND U3664 ( .A(B[3]), .B(A[177]), .Z(\ab[177][3] ) );
  AND U3665 ( .A(B[2]), .B(A[177]), .Z(\ab[177][2] ) );
  AND U3666 ( .A(B[1]), .B(A[177]), .Z(\ab[177][1] ) );
  AND U3667 ( .A(A[177]), .B(B[0]), .Z(\ab[177][0] ) );
  AND U3668 ( .A(B[3]), .B(A[176]), .Z(\ab[176][3] ) );
  AND U3669 ( .A(B[2]), .B(A[176]), .Z(\ab[176][2] ) );
  AND U3670 ( .A(B[1]), .B(A[176]), .Z(\ab[176][1] ) );
  AND U3671 ( .A(A[176]), .B(B[0]), .Z(\ab[176][0] ) );
  AND U3672 ( .A(B[3]), .B(A[175]), .Z(\ab[175][3] ) );
  AND U3673 ( .A(B[2]), .B(A[175]), .Z(\ab[175][2] ) );
  AND U3674 ( .A(B[1]), .B(A[175]), .Z(\ab[175][1] ) );
  AND U3675 ( .A(A[175]), .B(B[0]), .Z(\ab[175][0] ) );
  AND U3676 ( .A(B[3]), .B(A[174]), .Z(\ab[174][3] ) );
  AND U3677 ( .A(B[2]), .B(A[174]), .Z(\ab[174][2] ) );
  AND U3678 ( .A(B[1]), .B(A[174]), .Z(\ab[174][1] ) );
  AND U3679 ( .A(A[174]), .B(B[0]), .Z(\ab[174][0] ) );
  AND U3680 ( .A(B[3]), .B(A[173]), .Z(\ab[173][3] ) );
  AND U3681 ( .A(B[2]), .B(A[173]), .Z(\ab[173][2] ) );
  AND U3682 ( .A(B[1]), .B(A[173]), .Z(\ab[173][1] ) );
  AND U3683 ( .A(A[173]), .B(B[0]), .Z(\ab[173][0] ) );
  AND U3684 ( .A(B[3]), .B(A[172]), .Z(\ab[172][3] ) );
  AND U3685 ( .A(B[2]), .B(A[172]), .Z(\ab[172][2] ) );
  AND U3686 ( .A(B[1]), .B(A[172]), .Z(\ab[172][1] ) );
  AND U3687 ( .A(A[172]), .B(B[0]), .Z(\ab[172][0] ) );
  AND U3688 ( .A(B[3]), .B(A[171]), .Z(\ab[171][3] ) );
  AND U3689 ( .A(B[2]), .B(A[171]), .Z(\ab[171][2] ) );
  AND U3690 ( .A(B[1]), .B(A[171]), .Z(\ab[171][1] ) );
  AND U3691 ( .A(A[171]), .B(B[0]), .Z(\ab[171][0] ) );
  AND U3692 ( .A(B[3]), .B(A[170]), .Z(\ab[170][3] ) );
  AND U3693 ( .A(B[2]), .B(A[170]), .Z(\ab[170][2] ) );
  AND U3694 ( .A(B[1]), .B(A[170]), .Z(\ab[170][1] ) );
  AND U3695 ( .A(A[170]), .B(B[0]), .Z(\ab[170][0] ) );
  AND U3696 ( .A(B[3]), .B(A[16]), .Z(\ab[16][3] ) );
  AND U3697 ( .A(B[2]), .B(A[16]), .Z(\ab[16][2] ) );
  AND U3698 ( .A(B[1]), .B(A[16]), .Z(\ab[16][1] ) );
  AND U3699 ( .A(A[16]), .B(B[0]), .Z(\ab[16][0] ) );
  AND U3700 ( .A(B[3]), .B(A[169]), .Z(\ab[169][3] ) );
  AND U3701 ( .A(B[2]), .B(A[169]), .Z(\ab[169][2] ) );
  AND U3702 ( .A(B[1]), .B(A[169]), .Z(\ab[169][1] ) );
  AND U3703 ( .A(A[169]), .B(B[0]), .Z(\ab[169][0] ) );
  AND U3704 ( .A(B[3]), .B(A[168]), .Z(\ab[168][3] ) );
  AND U3705 ( .A(B[2]), .B(A[168]), .Z(\ab[168][2] ) );
  AND U3706 ( .A(B[1]), .B(A[168]), .Z(\ab[168][1] ) );
  AND U3707 ( .A(A[168]), .B(B[0]), .Z(\ab[168][0] ) );
  AND U3708 ( .A(B[3]), .B(A[167]), .Z(\ab[167][3] ) );
  AND U3709 ( .A(B[2]), .B(A[167]), .Z(\ab[167][2] ) );
  AND U3710 ( .A(B[1]), .B(A[167]), .Z(\ab[167][1] ) );
  AND U3711 ( .A(A[167]), .B(B[0]), .Z(\ab[167][0] ) );
  AND U3712 ( .A(B[3]), .B(A[166]), .Z(\ab[166][3] ) );
  AND U3713 ( .A(B[2]), .B(A[166]), .Z(\ab[166][2] ) );
  AND U3714 ( .A(B[1]), .B(A[166]), .Z(\ab[166][1] ) );
  AND U3715 ( .A(A[166]), .B(B[0]), .Z(\ab[166][0] ) );
  AND U3716 ( .A(B[3]), .B(A[165]), .Z(\ab[165][3] ) );
  AND U3717 ( .A(B[2]), .B(A[165]), .Z(\ab[165][2] ) );
  AND U3718 ( .A(B[1]), .B(A[165]), .Z(\ab[165][1] ) );
  AND U3719 ( .A(A[165]), .B(B[0]), .Z(\ab[165][0] ) );
  AND U3720 ( .A(B[3]), .B(A[164]), .Z(\ab[164][3] ) );
  AND U3721 ( .A(B[2]), .B(A[164]), .Z(\ab[164][2] ) );
  AND U3722 ( .A(B[1]), .B(A[164]), .Z(\ab[164][1] ) );
  AND U3723 ( .A(A[164]), .B(B[0]), .Z(\ab[164][0] ) );
  AND U3724 ( .A(B[3]), .B(A[163]), .Z(\ab[163][3] ) );
  AND U3725 ( .A(B[2]), .B(A[163]), .Z(\ab[163][2] ) );
  AND U3726 ( .A(B[1]), .B(A[163]), .Z(\ab[163][1] ) );
  AND U3727 ( .A(A[163]), .B(B[0]), .Z(\ab[163][0] ) );
  AND U3728 ( .A(B[3]), .B(A[162]), .Z(\ab[162][3] ) );
  AND U3729 ( .A(B[2]), .B(A[162]), .Z(\ab[162][2] ) );
  AND U3730 ( .A(B[1]), .B(A[162]), .Z(\ab[162][1] ) );
  AND U3731 ( .A(A[162]), .B(B[0]), .Z(\ab[162][0] ) );
  AND U3732 ( .A(B[3]), .B(A[161]), .Z(\ab[161][3] ) );
  AND U3733 ( .A(B[2]), .B(A[161]), .Z(\ab[161][2] ) );
  AND U3734 ( .A(B[1]), .B(A[161]), .Z(\ab[161][1] ) );
  AND U3735 ( .A(A[161]), .B(B[0]), .Z(\ab[161][0] ) );
  AND U3736 ( .A(B[3]), .B(A[160]), .Z(\ab[160][3] ) );
  AND U3737 ( .A(B[2]), .B(A[160]), .Z(\ab[160][2] ) );
  AND U3738 ( .A(B[1]), .B(A[160]), .Z(\ab[160][1] ) );
  AND U3739 ( .A(A[160]), .B(B[0]), .Z(\ab[160][0] ) );
  AND U3740 ( .A(B[3]), .B(A[15]), .Z(\ab[15][3] ) );
  AND U3741 ( .A(B[2]), .B(A[15]), .Z(\ab[15][2] ) );
  AND U3742 ( .A(B[1]), .B(A[15]), .Z(\ab[15][1] ) );
  AND U3743 ( .A(A[15]), .B(B[0]), .Z(\ab[15][0] ) );
  AND U3744 ( .A(B[3]), .B(A[159]), .Z(\ab[159][3] ) );
  AND U3745 ( .A(B[2]), .B(A[159]), .Z(\ab[159][2] ) );
  AND U3746 ( .A(B[1]), .B(A[159]), .Z(\ab[159][1] ) );
  AND U3747 ( .A(A[159]), .B(B[0]), .Z(\ab[159][0] ) );
  AND U3748 ( .A(B[3]), .B(A[158]), .Z(\ab[158][3] ) );
  AND U3749 ( .A(B[2]), .B(A[158]), .Z(\ab[158][2] ) );
  AND U3750 ( .A(B[1]), .B(A[158]), .Z(\ab[158][1] ) );
  AND U3751 ( .A(A[158]), .B(B[0]), .Z(\ab[158][0] ) );
  AND U3752 ( .A(B[3]), .B(A[157]), .Z(\ab[157][3] ) );
  AND U3753 ( .A(B[2]), .B(A[157]), .Z(\ab[157][2] ) );
  AND U3754 ( .A(B[1]), .B(A[157]), .Z(\ab[157][1] ) );
  AND U3755 ( .A(A[157]), .B(B[0]), .Z(\ab[157][0] ) );
  AND U3756 ( .A(B[3]), .B(A[156]), .Z(\ab[156][3] ) );
  AND U3757 ( .A(B[2]), .B(A[156]), .Z(\ab[156][2] ) );
  AND U3758 ( .A(B[1]), .B(A[156]), .Z(\ab[156][1] ) );
  AND U3759 ( .A(A[156]), .B(B[0]), .Z(\ab[156][0] ) );
  AND U3760 ( .A(B[3]), .B(A[155]), .Z(\ab[155][3] ) );
  AND U3761 ( .A(B[2]), .B(A[155]), .Z(\ab[155][2] ) );
  AND U3762 ( .A(B[1]), .B(A[155]), .Z(\ab[155][1] ) );
  AND U3763 ( .A(A[155]), .B(B[0]), .Z(\ab[155][0] ) );
  AND U3764 ( .A(B[3]), .B(A[154]), .Z(\ab[154][3] ) );
  AND U3765 ( .A(B[2]), .B(A[154]), .Z(\ab[154][2] ) );
  AND U3766 ( .A(B[1]), .B(A[154]), .Z(\ab[154][1] ) );
  AND U3767 ( .A(A[154]), .B(B[0]), .Z(\ab[154][0] ) );
  AND U3768 ( .A(B[3]), .B(A[153]), .Z(\ab[153][3] ) );
  AND U3769 ( .A(B[2]), .B(A[153]), .Z(\ab[153][2] ) );
  AND U3770 ( .A(B[1]), .B(A[153]), .Z(\ab[153][1] ) );
  AND U3771 ( .A(A[153]), .B(B[0]), .Z(\ab[153][0] ) );
  AND U3772 ( .A(B[3]), .B(A[152]), .Z(\ab[152][3] ) );
  AND U3773 ( .A(B[2]), .B(A[152]), .Z(\ab[152][2] ) );
  AND U3774 ( .A(B[1]), .B(A[152]), .Z(\ab[152][1] ) );
  AND U3775 ( .A(A[152]), .B(B[0]), .Z(\ab[152][0] ) );
  AND U3776 ( .A(B[3]), .B(A[151]), .Z(\ab[151][3] ) );
  AND U3777 ( .A(B[2]), .B(A[151]), .Z(\ab[151][2] ) );
  AND U3778 ( .A(B[1]), .B(A[151]), .Z(\ab[151][1] ) );
  AND U3779 ( .A(A[151]), .B(B[0]), .Z(\ab[151][0] ) );
  AND U3780 ( .A(B[3]), .B(A[150]), .Z(\ab[150][3] ) );
  AND U3781 ( .A(B[2]), .B(A[150]), .Z(\ab[150][2] ) );
  AND U3782 ( .A(B[1]), .B(A[150]), .Z(\ab[150][1] ) );
  AND U3783 ( .A(A[150]), .B(B[0]), .Z(\ab[150][0] ) );
  AND U3784 ( .A(B[3]), .B(A[14]), .Z(\ab[14][3] ) );
  AND U3785 ( .A(B[2]), .B(A[14]), .Z(\ab[14][2] ) );
  AND U3786 ( .A(B[1]), .B(A[14]), .Z(\ab[14][1] ) );
  AND U3787 ( .A(A[14]), .B(B[0]), .Z(\ab[14][0] ) );
  AND U3788 ( .A(B[3]), .B(A[149]), .Z(\ab[149][3] ) );
  AND U3789 ( .A(B[2]), .B(A[149]), .Z(\ab[149][2] ) );
  AND U3790 ( .A(B[1]), .B(A[149]), .Z(\ab[149][1] ) );
  AND U3791 ( .A(A[149]), .B(B[0]), .Z(\ab[149][0] ) );
  AND U3792 ( .A(B[3]), .B(A[148]), .Z(\ab[148][3] ) );
  AND U3793 ( .A(B[2]), .B(A[148]), .Z(\ab[148][2] ) );
  AND U3794 ( .A(B[1]), .B(A[148]), .Z(\ab[148][1] ) );
  AND U3795 ( .A(A[148]), .B(B[0]), .Z(\ab[148][0] ) );
  AND U3796 ( .A(B[3]), .B(A[147]), .Z(\ab[147][3] ) );
  AND U3797 ( .A(B[2]), .B(A[147]), .Z(\ab[147][2] ) );
  AND U3798 ( .A(B[1]), .B(A[147]), .Z(\ab[147][1] ) );
  AND U3799 ( .A(A[147]), .B(B[0]), .Z(\ab[147][0] ) );
  AND U3800 ( .A(B[3]), .B(A[146]), .Z(\ab[146][3] ) );
  AND U3801 ( .A(B[2]), .B(A[146]), .Z(\ab[146][2] ) );
  AND U3802 ( .A(B[1]), .B(A[146]), .Z(\ab[146][1] ) );
  AND U3803 ( .A(A[146]), .B(B[0]), .Z(\ab[146][0] ) );
  AND U3804 ( .A(B[3]), .B(A[145]), .Z(\ab[145][3] ) );
  AND U3805 ( .A(B[2]), .B(A[145]), .Z(\ab[145][2] ) );
  AND U3806 ( .A(B[1]), .B(A[145]), .Z(\ab[145][1] ) );
  AND U3807 ( .A(A[145]), .B(B[0]), .Z(\ab[145][0] ) );
  AND U3808 ( .A(B[3]), .B(A[144]), .Z(\ab[144][3] ) );
  AND U3809 ( .A(B[2]), .B(A[144]), .Z(\ab[144][2] ) );
  AND U3810 ( .A(B[1]), .B(A[144]), .Z(\ab[144][1] ) );
  AND U3811 ( .A(A[144]), .B(B[0]), .Z(\ab[144][0] ) );
  AND U3812 ( .A(B[3]), .B(A[143]), .Z(\ab[143][3] ) );
  AND U3813 ( .A(B[2]), .B(A[143]), .Z(\ab[143][2] ) );
  AND U3814 ( .A(B[1]), .B(A[143]), .Z(\ab[143][1] ) );
  AND U3815 ( .A(A[143]), .B(B[0]), .Z(\ab[143][0] ) );
  AND U3816 ( .A(B[3]), .B(A[142]), .Z(\ab[142][3] ) );
  AND U3817 ( .A(B[2]), .B(A[142]), .Z(\ab[142][2] ) );
  AND U3818 ( .A(B[1]), .B(A[142]), .Z(\ab[142][1] ) );
  AND U3819 ( .A(A[142]), .B(B[0]), .Z(\ab[142][0] ) );
  AND U3820 ( .A(B[3]), .B(A[141]), .Z(\ab[141][3] ) );
  AND U3821 ( .A(B[2]), .B(A[141]), .Z(\ab[141][2] ) );
  AND U3822 ( .A(B[1]), .B(A[141]), .Z(\ab[141][1] ) );
  AND U3823 ( .A(A[141]), .B(B[0]), .Z(\ab[141][0] ) );
  AND U3824 ( .A(B[3]), .B(A[140]), .Z(\ab[140][3] ) );
  AND U3825 ( .A(B[2]), .B(A[140]), .Z(\ab[140][2] ) );
  AND U3826 ( .A(B[1]), .B(A[140]), .Z(\ab[140][1] ) );
  AND U3827 ( .A(A[140]), .B(B[0]), .Z(\ab[140][0] ) );
  AND U3828 ( .A(B[3]), .B(A[13]), .Z(\ab[13][3] ) );
  AND U3829 ( .A(B[2]), .B(A[13]), .Z(\ab[13][2] ) );
  AND U3830 ( .A(B[1]), .B(A[13]), .Z(\ab[13][1] ) );
  AND U3831 ( .A(A[13]), .B(B[0]), .Z(\ab[13][0] ) );
  AND U3832 ( .A(B[3]), .B(A[139]), .Z(\ab[139][3] ) );
  AND U3833 ( .A(B[2]), .B(A[139]), .Z(\ab[139][2] ) );
  AND U3834 ( .A(B[1]), .B(A[139]), .Z(\ab[139][1] ) );
  AND U3835 ( .A(A[139]), .B(B[0]), .Z(\ab[139][0] ) );
  AND U3836 ( .A(B[3]), .B(A[138]), .Z(\ab[138][3] ) );
  AND U3837 ( .A(B[2]), .B(A[138]), .Z(\ab[138][2] ) );
  AND U3838 ( .A(B[1]), .B(A[138]), .Z(\ab[138][1] ) );
  AND U3839 ( .A(A[138]), .B(B[0]), .Z(\ab[138][0] ) );
  AND U3840 ( .A(B[3]), .B(A[137]), .Z(\ab[137][3] ) );
  AND U3841 ( .A(B[2]), .B(A[137]), .Z(\ab[137][2] ) );
  AND U3842 ( .A(B[1]), .B(A[137]), .Z(\ab[137][1] ) );
  AND U3843 ( .A(A[137]), .B(B[0]), .Z(\ab[137][0] ) );
  AND U3844 ( .A(B[3]), .B(A[136]), .Z(\ab[136][3] ) );
  AND U3845 ( .A(B[2]), .B(A[136]), .Z(\ab[136][2] ) );
  AND U3846 ( .A(B[1]), .B(A[136]), .Z(\ab[136][1] ) );
  AND U3847 ( .A(A[136]), .B(B[0]), .Z(\ab[136][0] ) );
  AND U3848 ( .A(B[3]), .B(A[135]), .Z(\ab[135][3] ) );
  AND U3849 ( .A(B[2]), .B(A[135]), .Z(\ab[135][2] ) );
  AND U3850 ( .A(B[1]), .B(A[135]), .Z(\ab[135][1] ) );
  AND U3851 ( .A(A[135]), .B(B[0]), .Z(\ab[135][0] ) );
  AND U3852 ( .A(B[3]), .B(A[134]), .Z(\ab[134][3] ) );
  AND U3853 ( .A(B[2]), .B(A[134]), .Z(\ab[134][2] ) );
  AND U3854 ( .A(B[1]), .B(A[134]), .Z(\ab[134][1] ) );
  AND U3855 ( .A(A[134]), .B(B[0]), .Z(\ab[134][0] ) );
  AND U3856 ( .A(B[3]), .B(A[133]), .Z(\ab[133][3] ) );
  AND U3857 ( .A(B[2]), .B(A[133]), .Z(\ab[133][2] ) );
  AND U3858 ( .A(B[1]), .B(A[133]), .Z(\ab[133][1] ) );
  AND U3859 ( .A(A[133]), .B(B[0]), .Z(\ab[133][0] ) );
  AND U3860 ( .A(B[3]), .B(A[132]), .Z(\ab[132][3] ) );
  AND U3861 ( .A(B[2]), .B(A[132]), .Z(\ab[132][2] ) );
  AND U3862 ( .A(B[1]), .B(A[132]), .Z(\ab[132][1] ) );
  AND U3863 ( .A(A[132]), .B(B[0]), .Z(\ab[132][0] ) );
  AND U3864 ( .A(B[3]), .B(A[131]), .Z(\ab[131][3] ) );
  AND U3865 ( .A(B[2]), .B(A[131]), .Z(\ab[131][2] ) );
  AND U3866 ( .A(B[1]), .B(A[131]), .Z(\ab[131][1] ) );
  AND U3867 ( .A(A[131]), .B(B[0]), .Z(\ab[131][0] ) );
  AND U3868 ( .A(B[3]), .B(A[130]), .Z(\ab[130][3] ) );
  AND U3869 ( .A(B[2]), .B(A[130]), .Z(\ab[130][2] ) );
  AND U3870 ( .A(B[1]), .B(A[130]), .Z(\ab[130][1] ) );
  AND U3871 ( .A(A[130]), .B(B[0]), .Z(\ab[130][0] ) );
  AND U3872 ( .A(B[3]), .B(A[12]), .Z(\ab[12][3] ) );
  AND U3873 ( .A(B[2]), .B(A[12]), .Z(\ab[12][2] ) );
  AND U3874 ( .A(B[1]), .B(A[12]), .Z(\ab[12][1] ) );
  AND U3875 ( .A(A[12]), .B(B[0]), .Z(\ab[12][0] ) );
  AND U3876 ( .A(B[3]), .B(A[129]), .Z(\ab[129][3] ) );
  AND U3877 ( .A(B[2]), .B(A[129]), .Z(\ab[129][2] ) );
  AND U3878 ( .A(B[1]), .B(A[129]), .Z(\ab[129][1] ) );
  AND U3879 ( .A(A[129]), .B(B[0]), .Z(\ab[129][0] ) );
  AND U3880 ( .A(B[3]), .B(A[128]), .Z(\ab[128][3] ) );
  AND U3881 ( .A(B[2]), .B(A[128]), .Z(\ab[128][2] ) );
  AND U3882 ( .A(B[1]), .B(A[128]), .Z(\ab[128][1] ) );
  AND U3883 ( .A(A[128]), .B(B[0]), .Z(\ab[128][0] ) );
  AND U3884 ( .A(B[3]), .B(A[127]), .Z(\ab[127][3] ) );
  AND U3885 ( .A(B[2]), .B(A[127]), .Z(\ab[127][2] ) );
  AND U3886 ( .A(B[1]), .B(A[127]), .Z(\ab[127][1] ) );
  AND U3887 ( .A(A[127]), .B(B[0]), .Z(\ab[127][0] ) );
  AND U3888 ( .A(B[3]), .B(A[126]), .Z(\ab[126][3] ) );
  AND U3889 ( .A(B[2]), .B(A[126]), .Z(\ab[126][2] ) );
  AND U3890 ( .A(B[1]), .B(A[126]), .Z(\ab[126][1] ) );
  AND U3891 ( .A(A[126]), .B(B[0]), .Z(\ab[126][0] ) );
  AND U3892 ( .A(B[3]), .B(A[125]), .Z(\ab[125][3] ) );
  AND U3893 ( .A(B[2]), .B(A[125]), .Z(\ab[125][2] ) );
  AND U3894 ( .A(B[1]), .B(A[125]), .Z(\ab[125][1] ) );
  AND U3895 ( .A(A[125]), .B(B[0]), .Z(\ab[125][0] ) );
  AND U3896 ( .A(B[3]), .B(A[124]), .Z(\ab[124][3] ) );
  AND U3897 ( .A(B[2]), .B(A[124]), .Z(\ab[124][2] ) );
  AND U3898 ( .A(B[1]), .B(A[124]), .Z(\ab[124][1] ) );
  AND U3899 ( .A(A[124]), .B(B[0]), .Z(\ab[124][0] ) );
  AND U3900 ( .A(B[3]), .B(A[123]), .Z(\ab[123][3] ) );
  AND U3901 ( .A(B[2]), .B(A[123]), .Z(\ab[123][2] ) );
  AND U3902 ( .A(B[1]), .B(A[123]), .Z(\ab[123][1] ) );
  AND U3903 ( .A(A[123]), .B(B[0]), .Z(\ab[123][0] ) );
  AND U3904 ( .A(B[3]), .B(A[122]), .Z(\ab[122][3] ) );
  AND U3905 ( .A(B[2]), .B(A[122]), .Z(\ab[122][2] ) );
  AND U3906 ( .A(B[1]), .B(A[122]), .Z(\ab[122][1] ) );
  AND U3907 ( .A(A[122]), .B(B[0]), .Z(\ab[122][0] ) );
  AND U3908 ( .A(B[3]), .B(A[121]), .Z(\ab[121][3] ) );
  AND U3909 ( .A(B[2]), .B(A[121]), .Z(\ab[121][2] ) );
  AND U3910 ( .A(B[1]), .B(A[121]), .Z(\ab[121][1] ) );
  AND U3911 ( .A(A[121]), .B(B[0]), .Z(\ab[121][0] ) );
  AND U3912 ( .A(B[3]), .B(A[120]), .Z(\ab[120][3] ) );
  AND U3913 ( .A(B[2]), .B(A[120]), .Z(\ab[120][2] ) );
  AND U3914 ( .A(B[1]), .B(A[120]), .Z(\ab[120][1] ) );
  AND U3915 ( .A(A[120]), .B(B[0]), .Z(\ab[120][0] ) );
  AND U3916 ( .A(B[3]), .B(A[11]), .Z(\ab[11][3] ) );
  AND U3917 ( .A(B[2]), .B(A[11]), .Z(\ab[11][2] ) );
  AND U3918 ( .A(B[1]), .B(A[11]), .Z(\ab[11][1] ) );
  AND U3919 ( .A(A[11]), .B(B[0]), .Z(\ab[11][0] ) );
  AND U3920 ( .A(B[3]), .B(A[119]), .Z(\ab[119][3] ) );
  AND U3921 ( .A(B[2]), .B(A[119]), .Z(\ab[119][2] ) );
  AND U3922 ( .A(B[1]), .B(A[119]), .Z(\ab[119][1] ) );
  AND U3923 ( .A(A[119]), .B(B[0]), .Z(\ab[119][0] ) );
  AND U3924 ( .A(B[3]), .B(A[118]), .Z(\ab[118][3] ) );
  AND U3925 ( .A(B[2]), .B(A[118]), .Z(\ab[118][2] ) );
  AND U3926 ( .A(B[1]), .B(A[118]), .Z(\ab[118][1] ) );
  AND U3927 ( .A(A[118]), .B(B[0]), .Z(\ab[118][0] ) );
  AND U3928 ( .A(B[3]), .B(A[117]), .Z(\ab[117][3] ) );
  AND U3929 ( .A(B[2]), .B(A[117]), .Z(\ab[117][2] ) );
  AND U3930 ( .A(B[1]), .B(A[117]), .Z(\ab[117][1] ) );
  AND U3931 ( .A(A[117]), .B(B[0]), .Z(\ab[117][0] ) );
  AND U3932 ( .A(B[3]), .B(A[116]), .Z(\ab[116][3] ) );
  AND U3933 ( .A(B[2]), .B(A[116]), .Z(\ab[116][2] ) );
  AND U3934 ( .A(B[1]), .B(A[116]), .Z(\ab[116][1] ) );
  AND U3935 ( .A(A[116]), .B(B[0]), .Z(\ab[116][0] ) );
  AND U3936 ( .A(B[3]), .B(A[115]), .Z(\ab[115][3] ) );
  AND U3937 ( .A(B[2]), .B(A[115]), .Z(\ab[115][2] ) );
  AND U3938 ( .A(B[1]), .B(A[115]), .Z(\ab[115][1] ) );
  AND U3939 ( .A(A[115]), .B(B[0]), .Z(\ab[115][0] ) );
  AND U3940 ( .A(B[3]), .B(A[114]), .Z(\ab[114][3] ) );
  AND U3941 ( .A(B[2]), .B(A[114]), .Z(\ab[114][2] ) );
  AND U3942 ( .A(B[1]), .B(A[114]), .Z(\ab[114][1] ) );
  AND U3943 ( .A(A[114]), .B(B[0]), .Z(\ab[114][0] ) );
  AND U3944 ( .A(B[3]), .B(A[113]), .Z(\ab[113][3] ) );
  AND U3945 ( .A(B[2]), .B(A[113]), .Z(\ab[113][2] ) );
  AND U3946 ( .A(B[1]), .B(A[113]), .Z(\ab[113][1] ) );
  AND U3947 ( .A(A[113]), .B(B[0]), .Z(\ab[113][0] ) );
  AND U3948 ( .A(B[3]), .B(A[112]), .Z(\ab[112][3] ) );
  AND U3949 ( .A(B[2]), .B(A[112]), .Z(\ab[112][2] ) );
  AND U3950 ( .A(B[1]), .B(A[112]), .Z(\ab[112][1] ) );
  AND U3951 ( .A(A[112]), .B(B[0]), .Z(\ab[112][0] ) );
  AND U3952 ( .A(B[3]), .B(A[111]), .Z(\ab[111][3] ) );
  AND U3953 ( .A(B[2]), .B(A[111]), .Z(\ab[111][2] ) );
  AND U3954 ( .A(B[1]), .B(A[111]), .Z(\ab[111][1] ) );
  AND U3955 ( .A(A[111]), .B(B[0]), .Z(\ab[111][0] ) );
  AND U3956 ( .A(B[3]), .B(A[110]), .Z(\ab[110][3] ) );
  AND U3957 ( .A(B[2]), .B(A[110]), .Z(\ab[110][2] ) );
  AND U3958 ( .A(B[1]), .B(A[110]), .Z(\ab[110][1] ) );
  AND U3959 ( .A(A[110]), .B(B[0]), .Z(\ab[110][0] ) );
  AND U3960 ( .A(B[3]), .B(A[10]), .Z(\ab[10][3] ) );
  AND U3961 ( .A(B[2]), .B(A[10]), .Z(\ab[10][2] ) );
  AND U3962 ( .A(B[1]), .B(A[10]), .Z(\ab[10][1] ) );
  AND U3963 ( .A(A[10]), .B(B[0]), .Z(\ab[10][0] ) );
  AND U3964 ( .A(B[3]), .B(A[109]), .Z(\ab[109][3] ) );
  AND U3965 ( .A(B[2]), .B(A[109]), .Z(\ab[109][2] ) );
  AND U3966 ( .A(B[1]), .B(A[109]), .Z(\ab[109][1] ) );
  AND U3967 ( .A(A[109]), .B(B[0]), .Z(\ab[109][0] ) );
  AND U3968 ( .A(B[3]), .B(A[108]), .Z(\ab[108][3] ) );
  AND U3969 ( .A(B[2]), .B(A[108]), .Z(\ab[108][2] ) );
  AND U3970 ( .A(B[1]), .B(A[108]), .Z(\ab[108][1] ) );
  AND U3971 ( .A(A[108]), .B(B[0]), .Z(\ab[108][0] ) );
  AND U3972 ( .A(B[3]), .B(A[107]), .Z(\ab[107][3] ) );
  AND U3973 ( .A(B[2]), .B(A[107]), .Z(\ab[107][2] ) );
  AND U3974 ( .A(B[1]), .B(A[107]), .Z(\ab[107][1] ) );
  AND U3975 ( .A(A[107]), .B(B[0]), .Z(\ab[107][0] ) );
  AND U3976 ( .A(B[3]), .B(A[106]), .Z(\ab[106][3] ) );
  AND U3977 ( .A(B[2]), .B(A[106]), .Z(\ab[106][2] ) );
  AND U3978 ( .A(B[1]), .B(A[106]), .Z(\ab[106][1] ) );
  AND U3979 ( .A(A[106]), .B(B[0]), .Z(\ab[106][0] ) );
  AND U3980 ( .A(B[3]), .B(A[105]), .Z(\ab[105][3] ) );
  AND U3981 ( .A(B[2]), .B(A[105]), .Z(\ab[105][2] ) );
  AND U3982 ( .A(B[1]), .B(A[105]), .Z(\ab[105][1] ) );
  AND U3983 ( .A(A[105]), .B(B[0]), .Z(\ab[105][0] ) );
  AND U3984 ( .A(B[3]), .B(A[104]), .Z(\ab[104][3] ) );
  AND U3985 ( .A(B[2]), .B(A[104]), .Z(\ab[104][2] ) );
  AND U3986 ( .A(B[1]), .B(A[104]), .Z(\ab[104][1] ) );
  AND U3987 ( .A(A[104]), .B(B[0]), .Z(\ab[104][0] ) );
  AND U3988 ( .A(B[3]), .B(A[103]), .Z(\ab[103][3] ) );
  AND U3989 ( .A(B[2]), .B(A[103]), .Z(\ab[103][2] ) );
  AND U3990 ( .A(B[1]), .B(A[103]), .Z(\ab[103][1] ) );
  AND U3991 ( .A(A[103]), .B(B[0]), .Z(\ab[103][0] ) );
  AND U3992 ( .A(B[3]), .B(A[102]), .Z(\ab[102][3] ) );
  AND U3993 ( .A(B[2]), .B(A[102]), .Z(\ab[102][2] ) );
  AND U3994 ( .A(B[1]), .B(A[102]), .Z(\ab[102][1] ) );
  AND U3995 ( .A(A[102]), .B(B[0]), .Z(\ab[102][0] ) );
  AND U3996 ( .A(A[1023]), .B(B[0]), .Z(\ab[1023][0] ) );
  AND U3997 ( .A(B[1]), .B(A[1022]), .Z(\ab[1022][1] ) );
  AND U3998 ( .A(A[1022]), .B(B[0]), .Z(\ab[1022][0] ) );
  AND U3999 ( .A(B[2]), .B(A[1021]), .Z(\ab[1021][2] ) );
  AND U4000 ( .A(B[1]), .B(A[1021]), .Z(\ab[1021][1] ) );
  AND U4001 ( .A(A[1021]), .B(B[0]), .Z(\ab[1021][0] ) );
  AND U4002 ( .A(B[3]), .B(A[1020]), .Z(\ab[1020][3] ) );
  AND U4003 ( .A(B[2]), .B(A[1020]), .Z(\ab[1020][2] ) );
  AND U4004 ( .A(B[1]), .B(A[1020]), .Z(\ab[1020][1] ) );
  AND U4005 ( .A(A[1020]), .B(B[0]), .Z(\ab[1020][0] ) );
  AND U4006 ( .A(B[3]), .B(A[101]), .Z(\ab[101][3] ) );
  AND U4007 ( .A(B[2]), .B(A[101]), .Z(\ab[101][2] ) );
  AND U4008 ( .A(B[1]), .B(A[101]), .Z(\ab[101][1] ) );
  AND U4009 ( .A(A[101]), .B(B[0]), .Z(\ab[101][0] ) );
  AND U4010 ( .A(B[3]), .B(A[1019]), .Z(\ab[1019][3] ) );
  AND U4011 ( .A(B[2]), .B(A[1019]), .Z(\ab[1019][2] ) );
  AND U4012 ( .A(B[1]), .B(A[1019]), .Z(\ab[1019][1] ) );
  AND U4013 ( .A(A[1019]), .B(B[0]), .Z(\ab[1019][0] ) );
  AND U4014 ( .A(B[3]), .B(A[1018]), .Z(\ab[1018][3] ) );
  AND U4015 ( .A(B[2]), .B(A[1018]), .Z(\ab[1018][2] ) );
  AND U4016 ( .A(B[1]), .B(A[1018]), .Z(\ab[1018][1] ) );
  AND U4017 ( .A(A[1018]), .B(B[0]), .Z(\ab[1018][0] ) );
  AND U4018 ( .A(B[3]), .B(A[1017]), .Z(\ab[1017][3] ) );
  AND U4019 ( .A(B[2]), .B(A[1017]), .Z(\ab[1017][2] ) );
  AND U4020 ( .A(B[1]), .B(A[1017]), .Z(\ab[1017][1] ) );
  AND U4021 ( .A(A[1017]), .B(B[0]), .Z(\ab[1017][0] ) );
  AND U4022 ( .A(B[3]), .B(A[1016]), .Z(\ab[1016][3] ) );
  AND U4023 ( .A(B[2]), .B(A[1016]), .Z(\ab[1016][2] ) );
  AND U4024 ( .A(B[1]), .B(A[1016]), .Z(\ab[1016][1] ) );
  AND U4025 ( .A(A[1016]), .B(B[0]), .Z(\ab[1016][0] ) );
  AND U4026 ( .A(B[3]), .B(A[1015]), .Z(\ab[1015][3] ) );
  AND U4027 ( .A(B[2]), .B(A[1015]), .Z(\ab[1015][2] ) );
  AND U4028 ( .A(B[1]), .B(A[1015]), .Z(\ab[1015][1] ) );
  AND U4029 ( .A(A[1015]), .B(B[0]), .Z(\ab[1015][0] ) );
  AND U4030 ( .A(B[3]), .B(A[1014]), .Z(\ab[1014][3] ) );
  AND U4031 ( .A(B[2]), .B(A[1014]), .Z(\ab[1014][2] ) );
  AND U4032 ( .A(B[1]), .B(A[1014]), .Z(\ab[1014][1] ) );
  AND U4033 ( .A(A[1014]), .B(B[0]), .Z(\ab[1014][0] ) );
  AND U4034 ( .A(B[3]), .B(A[1013]), .Z(\ab[1013][3] ) );
  AND U4035 ( .A(B[2]), .B(A[1013]), .Z(\ab[1013][2] ) );
  AND U4036 ( .A(B[1]), .B(A[1013]), .Z(\ab[1013][1] ) );
  AND U4037 ( .A(A[1013]), .B(B[0]), .Z(\ab[1013][0] ) );
  AND U4038 ( .A(B[3]), .B(A[1012]), .Z(\ab[1012][3] ) );
  AND U4039 ( .A(B[2]), .B(A[1012]), .Z(\ab[1012][2] ) );
  AND U4040 ( .A(B[1]), .B(A[1012]), .Z(\ab[1012][1] ) );
  AND U4041 ( .A(A[1012]), .B(B[0]), .Z(\ab[1012][0] ) );
  AND U4042 ( .A(B[3]), .B(A[1011]), .Z(\ab[1011][3] ) );
  AND U4043 ( .A(B[2]), .B(A[1011]), .Z(\ab[1011][2] ) );
  AND U4044 ( .A(B[1]), .B(A[1011]), .Z(\ab[1011][1] ) );
  AND U4045 ( .A(A[1011]), .B(B[0]), .Z(\ab[1011][0] ) );
  AND U4046 ( .A(B[3]), .B(A[1010]), .Z(\ab[1010][3] ) );
  AND U4047 ( .A(B[2]), .B(A[1010]), .Z(\ab[1010][2] ) );
  AND U4048 ( .A(B[1]), .B(A[1010]), .Z(\ab[1010][1] ) );
  AND U4049 ( .A(A[1010]), .B(B[0]), .Z(\ab[1010][0] ) );
  AND U4050 ( .A(B[3]), .B(A[100]), .Z(\ab[100][3] ) );
  AND U4051 ( .A(B[2]), .B(A[100]), .Z(\ab[100][2] ) );
  AND U4052 ( .A(B[1]), .B(A[100]), .Z(\ab[100][1] ) );
  AND U4053 ( .A(A[100]), .B(B[0]), .Z(\ab[100][0] ) );
  AND U4054 ( .A(B[3]), .B(A[1009]), .Z(\ab[1009][3] ) );
  AND U4055 ( .A(B[2]), .B(A[1009]), .Z(\ab[1009][2] ) );
  AND U4056 ( .A(B[1]), .B(A[1009]), .Z(\ab[1009][1] ) );
  AND U4057 ( .A(A[1009]), .B(B[0]), .Z(\ab[1009][0] ) );
  AND U4058 ( .A(B[3]), .B(A[1008]), .Z(\ab[1008][3] ) );
  AND U4059 ( .A(B[2]), .B(A[1008]), .Z(\ab[1008][2] ) );
  AND U4060 ( .A(B[1]), .B(A[1008]), .Z(\ab[1008][1] ) );
  AND U4061 ( .A(A[1008]), .B(B[0]), .Z(\ab[1008][0] ) );
  AND U4062 ( .A(B[3]), .B(A[1007]), .Z(\ab[1007][3] ) );
  AND U4063 ( .A(B[2]), .B(A[1007]), .Z(\ab[1007][2] ) );
  AND U4064 ( .A(B[1]), .B(A[1007]), .Z(\ab[1007][1] ) );
  AND U4065 ( .A(A[1007]), .B(B[0]), .Z(\ab[1007][0] ) );
  AND U4066 ( .A(B[3]), .B(A[1006]), .Z(\ab[1006][3] ) );
  AND U4067 ( .A(B[2]), .B(A[1006]), .Z(\ab[1006][2] ) );
  AND U4068 ( .A(B[1]), .B(A[1006]), .Z(\ab[1006][1] ) );
  AND U4069 ( .A(A[1006]), .B(B[0]), .Z(\ab[1006][0] ) );
  AND U4070 ( .A(B[3]), .B(A[1005]), .Z(\ab[1005][3] ) );
  AND U4071 ( .A(B[2]), .B(A[1005]), .Z(\ab[1005][2] ) );
  AND U4072 ( .A(B[1]), .B(A[1005]), .Z(\ab[1005][1] ) );
  AND U4073 ( .A(A[1005]), .B(B[0]), .Z(\ab[1005][0] ) );
  AND U4074 ( .A(B[3]), .B(A[1004]), .Z(\ab[1004][3] ) );
  AND U4075 ( .A(B[2]), .B(A[1004]), .Z(\ab[1004][2] ) );
  AND U4076 ( .A(B[1]), .B(A[1004]), .Z(\ab[1004][1] ) );
  AND U4077 ( .A(A[1004]), .B(B[0]), .Z(\ab[1004][0] ) );
  AND U4078 ( .A(B[3]), .B(A[1003]), .Z(\ab[1003][3] ) );
  AND U4079 ( .A(B[2]), .B(A[1003]), .Z(\ab[1003][2] ) );
  AND U4080 ( .A(B[1]), .B(A[1003]), .Z(\ab[1003][1] ) );
  AND U4081 ( .A(A[1003]), .B(B[0]), .Z(\ab[1003][0] ) );
  AND U4082 ( .A(B[3]), .B(A[1002]), .Z(\ab[1002][3] ) );
  AND U4083 ( .A(B[2]), .B(A[1002]), .Z(\ab[1002][2] ) );
  AND U4084 ( .A(B[1]), .B(A[1002]), .Z(\ab[1002][1] ) );
  AND U4085 ( .A(A[1002]), .B(B[0]), .Z(\ab[1002][0] ) );
  AND U4086 ( .A(B[3]), .B(A[1001]), .Z(\ab[1001][3] ) );
  AND U4087 ( .A(B[2]), .B(A[1001]), .Z(\ab[1001][2] ) );
  AND U4088 ( .A(B[1]), .B(A[1001]), .Z(\ab[1001][1] ) );
  AND U4089 ( .A(A[1001]), .B(B[0]), .Z(\ab[1001][0] ) );
  AND U4090 ( .A(B[3]), .B(A[1000]), .Z(\ab[1000][3] ) );
  AND U4091 ( .A(B[2]), .B(A[1000]), .Z(\ab[1000][2] ) );
  AND U4092 ( .A(B[1]), .B(A[1000]), .Z(\ab[1000][1] ) );
  AND U4093 ( .A(A[1000]), .B(B[0]), .Z(\ab[1000][0] ) );
  AND U4094 ( .A(B[3]), .B(A[0]), .Z(\ab[0][3] ) );
  AND U4095 ( .A(B[2]), .B(A[0]), .Z(\ab[0][2] ) );
  AND U4096 ( .A(B[1]), .B(A[0]), .Z(\ab[0][1] ) );
  AND U4097 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module mult_N1024_CC256 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [3:0] b;
  output [1023:0] c;
  input clk, rst;

  wire   [1023:4] swire;
  wire   [1023:0] clocal;
  wire   [2047:1024] sreg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  DFF \sreg_reg[1024]  ( .D(swire[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1024]) );
  DFF \sreg_reg[1025]  ( .D(swire[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1025]) );
  DFF \sreg_reg[1026]  ( .D(swire[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1026]) );
  DFF \sreg_reg[1027]  ( .D(swire[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1027]) );
  DFF \sreg_reg[1028]  ( .D(swire[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1028]) );
  DFF \sreg_reg[1029]  ( .D(swire[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1029]) );
  DFF \sreg_reg[1030]  ( .D(swire[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1030]) );
  DFF \sreg_reg[1031]  ( .D(swire[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1031]) );
  DFF \sreg_reg[1032]  ( .D(swire[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1032]) );
  DFF \sreg_reg[1033]  ( .D(swire[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1033]) );
  DFF \sreg_reg[1034]  ( .D(swire[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1034]) );
  DFF \sreg_reg[1035]  ( .D(swire[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1035]) );
  DFF \sreg_reg[1036]  ( .D(swire[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1036]) );
  DFF \sreg_reg[1037]  ( .D(swire[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1037]) );
  DFF \sreg_reg[1038]  ( .D(swire[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1038]) );
  DFF \sreg_reg[1039]  ( .D(swire[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1039]) );
  DFF \sreg_reg[1040]  ( .D(swire[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1040]) );
  DFF \sreg_reg[1041]  ( .D(swire[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1041]) );
  DFF \sreg_reg[1042]  ( .D(swire[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1042]) );
  DFF \sreg_reg[1043]  ( .D(swire[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1043]) );
  DFF \sreg_reg[1044]  ( .D(swire[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1044]) );
  DFF \sreg_reg[1045]  ( .D(swire[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1045]) );
  DFF \sreg_reg[1046]  ( .D(swire[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1046]) );
  DFF \sreg_reg[1047]  ( .D(swire[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1047]) );
  DFF \sreg_reg[1048]  ( .D(swire[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1048]) );
  DFF \sreg_reg[1049]  ( .D(swire[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1049]) );
  DFF \sreg_reg[1050]  ( .D(swire[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1050]) );
  DFF \sreg_reg[1051]  ( .D(swire[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1051]) );
  DFF \sreg_reg[1052]  ( .D(swire[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1052]) );
  DFF \sreg_reg[1053]  ( .D(swire[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1053]) );
  DFF \sreg_reg[1054]  ( .D(swire[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1054]) );
  DFF \sreg_reg[1055]  ( .D(swire[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1055]) );
  DFF \sreg_reg[1056]  ( .D(swire[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1056]) );
  DFF \sreg_reg[1057]  ( .D(swire[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1057]) );
  DFF \sreg_reg[1058]  ( .D(swire[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1058]) );
  DFF \sreg_reg[1059]  ( .D(swire[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1059]) );
  DFF \sreg_reg[1060]  ( .D(swire[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1060]) );
  DFF \sreg_reg[1061]  ( .D(swire[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1061]) );
  DFF \sreg_reg[1062]  ( .D(swire[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1062]) );
  DFF \sreg_reg[1063]  ( .D(swire[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1063]) );
  DFF \sreg_reg[1064]  ( .D(swire[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1064]) );
  DFF \sreg_reg[1065]  ( .D(swire[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1065]) );
  DFF \sreg_reg[1066]  ( .D(swire[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1066]) );
  DFF \sreg_reg[1067]  ( .D(swire[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1067]) );
  DFF \sreg_reg[1068]  ( .D(swire[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1068]) );
  DFF \sreg_reg[1069]  ( .D(swire[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1069]) );
  DFF \sreg_reg[1070]  ( .D(swire[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1070]) );
  DFF \sreg_reg[1071]  ( .D(swire[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1071]) );
  DFF \sreg_reg[1072]  ( .D(swire[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1072]) );
  DFF \sreg_reg[1073]  ( .D(swire[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1073]) );
  DFF \sreg_reg[1074]  ( .D(swire[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1074]) );
  DFF \sreg_reg[1075]  ( .D(swire[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1075]) );
  DFF \sreg_reg[1076]  ( .D(swire[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1076]) );
  DFF \sreg_reg[1077]  ( .D(swire[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1077]) );
  DFF \sreg_reg[1078]  ( .D(swire[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1078]) );
  DFF \sreg_reg[1079]  ( .D(swire[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1079]) );
  DFF \sreg_reg[1080]  ( .D(swire[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1080]) );
  DFF \sreg_reg[1081]  ( .D(swire[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1081]) );
  DFF \sreg_reg[1082]  ( .D(swire[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1082]) );
  DFF \sreg_reg[1083]  ( .D(swire[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1083]) );
  DFF \sreg_reg[1084]  ( .D(swire[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1084]) );
  DFF \sreg_reg[1085]  ( .D(swire[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1085]) );
  DFF \sreg_reg[1086]  ( .D(swire[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1086]) );
  DFF \sreg_reg[1087]  ( .D(swire[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1087]) );
  DFF \sreg_reg[1088]  ( .D(swire[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1088]) );
  DFF \sreg_reg[1089]  ( .D(swire[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1089]) );
  DFF \sreg_reg[1090]  ( .D(swire[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1090]) );
  DFF \sreg_reg[1091]  ( .D(swire[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1091]) );
  DFF \sreg_reg[1092]  ( .D(swire[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1092]) );
  DFF \sreg_reg[1093]  ( .D(swire[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1093]) );
  DFF \sreg_reg[1094]  ( .D(swire[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1094]) );
  DFF \sreg_reg[1095]  ( .D(swire[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1095]) );
  DFF \sreg_reg[1096]  ( .D(swire[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1096]) );
  DFF \sreg_reg[1097]  ( .D(swire[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1097]) );
  DFF \sreg_reg[1098]  ( .D(swire[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1098]) );
  DFF \sreg_reg[1099]  ( .D(swire[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1099]) );
  DFF \sreg_reg[1100]  ( .D(swire[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1100]) );
  DFF \sreg_reg[1101]  ( .D(swire[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1101]) );
  DFF \sreg_reg[1102]  ( .D(swire[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1102]) );
  DFF \sreg_reg[1103]  ( .D(swire[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1103]) );
  DFF \sreg_reg[1104]  ( .D(swire[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1104]) );
  DFF \sreg_reg[1105]  ( .D(swire[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1105]) );
  DFF \sreg_reg[1106]  ( .D(swire[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1106]) );
  DFF \sreg_reg[1107]  ( .D(swire[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1107]) );
  DFF \sreg_reg[1108]  ( .D(swire[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1108]) );
  DFF \sreg_reg[1109]  ( .D(swire[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1109]) );
  DFF \sreg_reg[1110]  ( .D(swire[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1110]) );
  DFF \sreg_reg[1111]  ( .D(swire[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1111]) );
  DFF \sreg_reg[1112]  ( .D(swire[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1112]) );
  DFF \sreg_reg[1113]  ( .D(swire[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1113]) );
  DFF \sreg_reg[1114]  ( .D(swire[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1114]) );
  DFF \sreg_reg[1115]  ( .D(swire[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1115]) );
  DFF \sreg_reg[1116]  ( .D(swire[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1116]) );
  DFF \sreg_reg[1117]  ( .D(swire[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1117]) );
  DFF \sreg_reg[1118]  ( .D(swire[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1118]) );
  DFF \sreg_reg[1119]  ( .D(swire[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1119]) );
  DFF \sreg_reg[1120]  ( .D(swire[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1120]) );
  DFF \sreg_reg[1121]  ( .D(swire[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1121]) );
  DFF \sreg_reg[1122]  ( .D(swire[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1122]) );
  DFF \sreg_reg[1123]  ( .D(swire[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1123]) );
  DFF \sreg_reg[1124]  ( .D(swire[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1124]) );
  DFF \sreg_reg[1125]  ( .D(swire[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1125]) );
  DFF \sreg_reg[1126]  ( .D(swire[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1126]) );
  DFF \sreg_reg[1127]  ( .D(swire[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1127]) );
  DFF \sreg_reg[1128]  ( .D(swire[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1128]) );
  DFF \sreg_reg[1129]  ( .D(swire[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1129]) );
  DFF \sreg_reg[1130]  ( .D(swire[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1130]) );
  DFF \sreg_reg[1131]  ( .D(swire[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1131]) );
  DFF \sreg_reg[1132]  ( .D(swire[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1132]) );
  DFF \sreg_reg[1133]  ( .D(swire[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1133]) );
  DFF \sreg_reg[1134]  ( .D(swire[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1134]) );
  DFF \sreg_reg[1135]  ( .D(swire[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1135]) );
  DFF \sreg_reg[1136]  ( .D(swire[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1136]) );
  DFF \sreg_reg[1137]  ( .D(swire[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1137]) );
  DFF \sreg_reg[1138]  ( .D(swire[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1138]) );
  DFF \sreg_reg[1139]  ( .D(swire[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1139]) );
  DFF \sreg_reg[1140]  ( .D(swire[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1140]) );
  DFF \sreg_reg[1141]  ( .D(swire[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1141]) );
  DFF \sreg_reg[1142]  ( .D(swire[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1142]) );
  DFF \sreg_reg[1143]  ( .D(swire[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1143]) );
  DFF \sreg_reg[1144]  ( .D(swire[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1144]) );
  DFF \sreg_reg[1145]  ( .D(swire[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1145]) );
  DFF \sreg_reg[1146]  ( .D(swire[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1146]) );
  DFF \sreg_reg[1147]  ( .D(swire[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1147]) );
  DFF \sreg_reg[1148]  ( .D(swire[128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1148]) );
  DFF \sreg_reg[1149]  ( .D(swire[129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1149]) );
  DFF \sreg_reg[1150]  ( .D(swire[130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1150]) );
  DFF \sreg_reg[1151]  ( .D(swire[131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1151]) );
  DFF \sreg_reg[1152]  ( .D(swire[132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1152]) );
  DFF \sreg_reg[1153]  ( .D(swire[133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1153]) );
  DFF \sreg_reg[1154]  ( .D(swire[134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1154]) );
  DFF \sreg_reg[1155]  ( .D(swire[135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1155]) );
  DFF \sreg_reg[1156]  ( .D(swire[136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1156]) );
  DFF \sreg_reg[1157]  ( .D(swire[137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1157]) );
  DFF \sreg_reg[1158]  ( .D(swire[138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1158]) );
  DFF \sreg_reg[1159]  ( .D(swire[139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1159]) );
  DFF \sreg_reg[1160]  ( .D(swire[140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1160]) );
  DFF \sreg_reg[1161]  ( .D(swire[141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1161]) );
  DFF \sreg_reg[1162]  ( .D(swire[142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1162]) );
  DFF \sreg_reg[1163]  ( .D(swire[143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1163]) );
  DFF \sreg_reg[1164]  ( .D(swire[144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1164]) );
  DFF \sreg_reg[1165]  ( .D(swire[145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1165]) );
  DFF \sreg_reg[1166]  ( .D(swire[146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1166]) );
  DFF \sreg_reg[1167]  ( .D(swire[147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1167]) );
  DFF \sreg_reg[1168]  ( .D(swire[148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1168]) );
  DFF \sreg_reg[1169]  ( .D(swire[149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1169]) );
  DFF \sreg_reg[1170]  ( .D(swire[150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1170]) );
  DFF \sreg_reg[1171]  ( .D(swire[151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1171]) );
  DFF \sreg_reg[1172]  ( .D(swire[152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1172]) );
  DFF \sreg_reg[1173]  ( .D(swire[153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1173]) );
  DFF \sreg_reg[1174]  ( .D(swire[154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1174]) );
  DFF \sreg_reg[1175]  ( .D(swire[155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1175]) );
  DFF \sreg_reg[1176]  ( .D(swire[156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1176]) );
  DFF \sreg_reg[1177]  ( .D(swire[157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1177]) );
  DFF \sreg_reg[1178]  ( .D(swire[158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1178]) );
  DFF \sreg_reg[1179]  ( .D(swire[159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1179]) );
  DFF \sreg_reg[1180]  ( .D(swire[160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1180]) );
  DFF \sreg_reg[1181]  ( .D(swire[161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1181]) );
  DFF \sreg_reg[1182]  ( .D(swire[162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1182]) );
  DFF \sreg_reg[1183]  ( .D(swire[163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1183]) );
  DFF \sreg_reg[1184]  ( .D(swire[164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1184]) );
  DFF \sreg_reg[1185]  ( .D(swire[165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1185]) );
  DFF \sreg_reg[1186]  ( .D(swire[166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1186]) );
  DFF \sreg_reg[1187]  ( .D(swire[167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1187]) );
  DFF \sreg_reg[1188]  ( .D(swire[168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1188]) );
  DFF \sreg_reg[1189]  ( .D(swire[169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1189]) );
  DFF \sreg_reg[1190]  ( .D(swire[170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1190]) );
  DFF \sreg_reg[1191]  ( .D(swire[171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1191]) );
  DFF \sreg_reg[1192]  ( .D(swire[172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1192]) );
  DFF \sreg_reg[1193]  ( .D(swire[173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1193]) );
  DFF \sreg_reg[1194]  ( .D(swire[174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1194]) );
  DFF \sreg_reg[1195]  ( .D(swire[175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1195]) );
  DFF \sreg_reg[1196]  ( .D(swire[176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1196]) );
  DFF \sreg_reg[1197]  ( .D(swire[177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1197]) );
  DFF \sreg_reg[1198]  ( .D(swire[178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1198]) );
  DFF \sreg_reg[1199]  ( .D(swire[179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1199]) );
  DFF \sreg_reg[1200]  ( .D(swire[180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1200]) );
  DFF \sreg_reg[1201]  ( .D(swire[181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1201]) );
  DFF \sreg_reg[1202]  ( .D(swire[182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1202]) );
  DFF \sreg_reg[1203]  ( .D(swire[183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1203]) );
  DFF \sreg_reg[1204]  ( .D(swire[184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1204]) );
  DFF \sreg_reg[1205]  ( .D(swire[185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1205]) );
  DFF \sreg_reg[1206]  ( .D(swire[186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1206]) );
  DFF \sreg_reg[1207]  ( .D(swire[187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1207]) );
  DFF \sreg_reg[1208]  ( .D(swire[188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1208]) );
  DFF \sreg_reg[1209]  ( .D(swire[189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1209]) );
  DFF \sreg_reg[1210]  ( .D(swire[190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1210]) );
  DFF \sreg_reg[1211]  ( .D(swire[191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1211]) );
  DFF \sreg_reg[1212]  ( .D(swire[192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1212]) );
  DFF \sreg_reg[1213]  ( .D(swire[193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1213]) );
  DFF \sreg_reg[1214]  ( .D(swire[194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1214]) );
  DFF \sreg_reg[1215]  ( .D(swire[195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1215]) );
  DFF \sreg_reg[1216]  ( .D(swire[196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1216]) );
  DFF \sreg_reg[1217]  ( .D(swire[197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1217]) );
  DFF \sreg_reg[1218]  ( .D(swire[198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1218]) );
  DFF \sreg_reg[1219]  ( .D(swire[199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1219]) );
  DFF \sreg_reg[1220]  ( .D(swire[200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1220]) );
  DFF \sreg_reg[1221]  ( .D(swire[201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1221]) );
  DFF \sreg_reg[1222]  ( .D(swire[202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1222]) );
  DFF \sreg_reg[1223]  ( .D(swire[203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1223]) );
  DFF \sreg_reg[1224]  ( .D(swire[204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1224]) );
  DFF \sreg_reg[1225]  ( .D(swire[205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1225]) );
  DFF \sreg_reg[1226]  ( .D(swire[206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1226]) );
  DFF \sreg_reg[1227]  ( .D(swire[207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1227]) );
  DFF \sreg_reg[1228]  ( .D(swire[208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1228]) );
  DFF \sreg_reg[1229]  ( .D(swire[209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1229]) );
  DFF \sreg_reg[1230]  ( .D(swire[210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1230]) );
  DFF \sreg_reg[1231]  ( .D(swire[211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1231]) );
  DFF \sreg_reg[1232]  ( .D(swire[212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1232]) );
  DFF \sreg_reg[1233]  ( .D(swire[213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1233]) );
  DFF \sreg_reg[1234]  ( .D(swire[214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1234]) );
  DFF \sreg_reg[1235]  ( .D(swire[215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1235]) );
  DFF \sreg_reg[1236]  ( .D(swire[216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1236]) );
  DFF \sreg_reg[1237]  ( .D(swire[217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1237]) );
  DFF \sreg_reg[1238]  ( .D(swire[218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1238]) );
  DFF \sreg_reg[1239]  ( .D(swire[219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1239]) );
  DFF \sreg_reg[1240]  ( .D(swire[220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1240]) );
  DFF \sreg_reg[1241]  ( .D(swire[221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1241]) );
  DFF \sreg_reg[1242]  ( .D(swire[222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1242]) );
  DFF \sreg_reg[1243]  ( .D(swire[223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1243]) );
  DFF \sreg_reg[1244]  ( .D(swire[224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1244]) );
  DFF \sreg_reg[1245]  ( .D(swire[225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1245]) );
  DFF \sreg_reg[1246]  ( .D(swire[226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1246]) );
  DFF \sreg_reg[1247]  ( .D(swire[227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1247]) );
  DFF \sreg_reg[1248]  ( .D(swire[228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1248]) );
  DFF \sreg_reg[1249]  ( .D(swire[229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1249]) );
  DFF \sreg_reg[1250]  ( .D(swire[230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1250]) );
  DFF \sreg_reg[1251]  ( .D(swire[231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1251]) );
  DFF \sreg_reg[1252]  ( .D(swire[232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1252]) );
  DFF \sreg_reg[1253]  ( .D(swire[233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1253]) );
  DFF \sreg_reg[1254]  ( .D(swire[234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1254]) );
  DFF \sreg_reg[1255]  ( .D(swire[235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1255]) );
  DFF \sreg_reg[1256]  ( .D(swire[236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1256]) );
  DFF \sreg_reg[1257]  ( .D(swire[237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1257]) );
  DFF \sreg_reg[1258]  ( .D(swire[238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1258]) );
  DFF \sreg_reg[1259]  ( .D(swire[239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1259]) );
  DFF \sreg_reg[1260]  ( .D(swire[240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1260]) );
  DFF \sreg_reg[1261]  ( .D(swire[241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1261]) );
  DFF \sreg_reg[1262]  ( .D(swire[242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1262]) );
  DFF \sreg_reg[1263]  ( .D(swire[243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1263]) );
  DFF \sreg_reg[1264]  ( .D(swire[244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1264]) );
  DFF \sreg_reg[1265]  ( .D(swire[245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1265]) );
  DFF \sreg_reg[1266]  ( .D(swire[246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1266]) );
  DFF \sreg_reg[1267]  ( .D(swire[247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1267]) );
  DFF \sreg_reg[1268]  ( .D(swire[248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1268]) );
  DFF \sreg_reg[1269]  ( .D(swire[249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1269]) );
  DFF \sreg_reg[1270]  ( .D(swire[250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1270]) );
  DFF \sreg_reg[1271]  ( .D(swire[251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1271]) );
  DFF \sreg_reg[1272]  ( .D(swire[252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1272]) );
  DFF \sreg_reg[1273]  ( .D(swire[253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1273]) );
  DFF \sreg_reg[1274]  ( .D(swire[254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1274]) );
  DFF \sreg_reg[1275]  ( .D(swire[255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1275]) );
  DFF \sreg_reg[1276]  ( .D(swire[256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1276]) );
  DFF \sreg_reg[1277]  ( .D(swire[257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1277]) );
  DFF \sreg_reg[1278]  ( .D(swire[258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1278]) );
  DFF \sreg_reg[1279]  ( .D(swire[259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1279]) );
  DFF \sreg_reg[1280]  ( .D(swire[260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1280]) );
  DFF \sreg_reg[1281]  ( .D(swire[261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1281]) );
  DFF \sreg_reg[1282]  ( .D(swire[262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1282]) );
  DFF \sreg_reg[1283]  ( .D(swire[263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1283]) );
  DFF \sreg_reg[1284]  ( .D(swire[264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1284]) );
  DFF \sreg_reg[1285]  ( .D(swire[265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1285]) );
  DFF \sreg_reg[1286]  ( .D(swire[266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1286]) );
  DFF \sreg_reg[1287]  ( .D(swire[267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1287]) );
  DFF \sreg_reg[1288]  ( .D(swire[268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1288]) );
  DFF \sreg_reg[1289]  ( .D(swire[269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1289]) );
  DFF \sreg_reg[1290]  ( .D(swire[270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1290]) );
  DFF \sreg_reg[1291]  ( .D(swire[271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1291]) );
  DFF \sreg_reg[1292]  ( .D(swire[272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1292]) );
  DFF \sreg_reg[1293]  ( .D(swire[273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1293]) );
  DFF \sreg_reg[1294]  ( .D(swire[274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1294]) );
  DFF \sreg_reg[1295]  ( .D(swire[275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1295]) );
  DFF \sreg_reg[1296]  ( .D(swire[276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1296]) );
  DFF \sreg_reg[1297]  ( .D(swire[277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1297]) );
  DFF \sreg_reg[1298]  ( .D(swire[278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1298]) );
  DFF \sreg_reg[1299]  ( .D(swire[279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1299]) );
  DFF \sreg_reg[1300]  ( .D(swire[280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1300]) );
  DFF \sreg_reg[1301]  ( .D(swire[281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1301]) );
  DFF \sreg_reg[1302]  ( .D(swire[282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1302]) );
  DFF \sreg_reg[1303]  ( .D(swire[283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1303]) );
  DFF \sreg_reg[1304]  ( .D(swire[284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1304]) );
  DFF \sreg_reg[1305]  ( .D(swire[285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1305]) );
  DFF \sreg_reg[1306]  ( .D(swire[286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1306]) );
  DFF \sreg_reg[1307]  ( .D(swire[287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1307]) );
  DFF \sreg_reg[1308]  ( .D(swire[288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1308]) );
  DFF \sreg_reg[1309]  ( .D(swire[289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1309]) );
  DFF \sreg_reg[1310]  ( .D(swire[290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1310]) );
  DFF \sreg_reg[1311]  ( .D(swire[291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1311]) );
  DFF \sreg_reg[1312]  ( .D(swire[292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1312]) );
  DFF \sreg_reg[1313]  ( .D(swire[293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1313]) );
  DFF \sreg_reg[1314]  ( .D(swire[294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1314]) );
  DFF \sreg_reg[1315]  ( .D(swire[295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1315]) );
  DFF \sreg_reg[1316]  ( .D(swire[296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1316]) );
  DFF \sreg_reg[1317]  ( .D(swire[297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1317]) );
  DFF \sreg_reg[1318]  ( .D(swire[298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1318]) );
  DFF \sreg_reg[1319]  ( .D(swire[299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1319]) );
  DFF \sreg_reg[1320]  ( .D(swire[300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1320]) );
  DFF \sreg_reg[1321]  ( .D(swire[301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1321]) );
  DFF \sreg_reg[1322]  ( .D(swire[302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1322]) );
  DFF \sreg_reg[1323]  ( .D(swire[303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1323]) );
  DFF \sreg_reg[1324]  ( .D(swire[304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1324]) );
  DFF \sreg_reg[1325]  ( .D(swire[305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1325]) );
  DFF \sreg_reg[1326]  ( .D(swire[306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1326]) );
  DFF \sreg_reg[1327]  ( .D(swire[307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1327]) );
  DFF \sreg_reg[1328]  ( .D(swire[308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1328]) );
  DFF \sreg_reg[1329]  ( .D(swire[309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1329]) );
  DFF \sreg_reg[1330]  ( .D(swire[310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1330]) );
  DFF \sreg_reg[1331]  ( .D(swire[311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1331]) );
  DFF \sreg_reg[1332]  ( .D(swire[312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1332]) );
  DFF \sreg_reg[1333]  ( .D(swire[313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1333]) );
  DFF \sreg_reg[1334]  ( .D(swire[314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1334]) );
  DFF \sreg_reg[1335]  ( .D(swire[315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1335]) );
  DFF \sreg_reg[1336]  ( .D(swire[316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1336]) );
  DFF \sreg_reg[1337]  ( .D(swire[317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1337]) );
  DFF \sreg_reg[1338]  ( .D(swire[318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1338]) );
  DFF \sreg_reg[1339]  ( .D(swire[319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1339]) );
  DFF \sreg_reg[1340]  ( .D(swire[320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1340]) );
  DFF \sreg_reg[1341]  ( .D(swire[321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1341]) );
  DFF \sreg_reg[1342]  ( .D(swire[322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1342]) );
  DFF \sreg_reg[1343]  ( .D(swire[323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1343]) );
  DFF \sreg_reg[1344]  ( .D(swire[324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1344]) );
  DFF \sreg_reg[1345]  ( .D(swire[325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1345]) );
  DFF \sreg_reg[1346]  ( .D(swire[326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1346]) );
  DFF \sreg_reg[1347]  ( .D(swire[327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1347]) );
  DFF \sreg_reg[1348]  ( .D(swire[328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1348]) );
  DFF \sreg_reg[1349]  ( .D(swire[329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1349]) );
  DFF \sreg_reg[1350]  ( .D(swire[330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1350]) );
  DFF \sreg_reg[1351]  ( .D(swire[331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1351]) );
  DFF \sreg_reg[1352]  ( .D(swire[332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1352]) );
  DFF \sreg_reg[1353]  ( .D(swire[333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1353]) );
  DFF \sreg_reg[1354]  ( .D(swire[334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1354]) );
  DFF \sreg_reg[1355]  ( .D(swire[335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1355]) );
  DFF \sreg_reg[1356]  ( .D(swire[336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1356]) );
  DFF \sreg_reg[1357]  ( .D(swire[337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1357]) );
  DFF \sreg_reg[1358]  ( .D(swire[338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1358]) );
  DFF \sreg_reg[1359]  ( .D(swire[339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1359]) );
  DFF \sreg_reg[1360]  ( .D(swire[340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1360]) );
  DFF \sreg_reg[1361]  ( .D(swire[341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1361]) );
  DFF \sreg_reg[1362]  ( .D(swire[342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1362]) );
  DFF \sreg_reg[1363]  ( .D(swire[343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1363]) );
  DFF \sreg_reg[1364]  ( .D(swire[344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1364]) );
  DFF \sreg_reg[1365]  ( .D(swire[345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1365]) );
  DFF \sreg_reg[1366]  ( .D(swire[346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1366]) );
  DFF \sreg_reg[1367]  ( .D(swire[347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1367]) );
  DFF \sreg_reg[1368]  ( .D(swire[348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1368]) );
  DFF \sreg_reg[1369]  ( .D(swire[349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1369]) );
  DFF \sreg_reg[1370]  ( .D(swire[350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1370]) );
  DFF \sreg_reg[1371]  ( .D(swire[351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1371]) );
  DFF \sreg_reg[1372]  ( .D(swire[352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1372]) );
  DFF \sreg_reg[1373]  ( .D(swire[353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1373]) );
  DFF \sreg_reg[1374]  ( .D(swire[354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1374]) );
  DFF \sreg_reg[1375]  ( .D(swire[355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1375]) );
  DFF \sreg_reg[1376]  ( .D(swire[356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1376]) );
  DFF \sreg_reg[1377]  ( .D(swire[357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1377]) );
  DFF \sreg_reg[1378]  ( .D(swire[358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1378]) );
  DFF \sreg_reg[1379]  ( .D(swire[359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1379]) );
  DFF \sreg_reg[1380]  ( .D(swire[360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1380]) );
  DFF \sreg_reg[1381]  ( .D(swire[361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1381]) );
  DFF \sreg_reg[1382]  ( .D(swire[362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1382]) );
  DFF \sreg_reg[1383]  ( .D(swire[363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1383]) );
  DFF \sreg_reg[1384]  ( .D(swire[364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1384]) );
  DFF \sreg_reg[1385]  ( .D(swire[365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1385]) );
  DFF \sreg_reg[1386]  ( .D(swire[366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1386]) );
  DFF \sreg_reg[1387]  ( .D(swire[367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1387]) );
  DFF \sreg_reg[1388]  ( .D(swire[368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1388]) );
  DFF \sreg_reg[1389]  ( .D(swire[369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1389]) );
  DFF \sreg_reg[1390]  ( .D(swire[370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1390]) );
  DFF \sreg_reg[1391]  ( .D(swire[371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1391]) );
  DFF \sreg_reg[1392]  ( .D(swire[372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1392]) );
  DFF \sreg_reg[1393]  ( .D(swire[373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1393]) );
  DFF \sreg_reg[1394]  ( .D(swire[374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1394]) );
  DFF \sreg_reg[1395]  ( .D(swire[375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1395]) );
  DFF \sreg_reg[1396]  ( .D(swire[376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1396]) );
  DFF \sreg_reg[1397]  ( .D(swire[377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1397]) );
  DFF \sreg_reg[1398]  ( .D(swire[378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1398]) );
  DFF \sreg_reg[1399]  ( .D(swire[379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1399]) );
  DFF \sreg_reg[1400]  ( .D(swire[380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1400]) );
  DFF \sreg_reg[1401]  ( .D(swire[381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1401]) );
  DFF \sreg_reg[1402]  ( .D(swire[382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1402]) );
  DFF \sreg_reg[1403]  ( .D(swire[383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1403]) );
  DFF \sreg_reg[1404]  ( .D(swire[384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1404]) );
  DFF \sreg_reg[1405]  ( .D(swire[385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1405]) );
  DFF \sreg_reg[1406]  ( .D(swire[386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1406]) );
  DFF \sreg_reg[1407]  ( .D(swire[387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1407]) );
  DFF \sreg_reg[1408]  ( .D(swire[388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1408]) );
  DFF \sreg_reg[1409]  ( .D(swire[389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1409]) );
  DFF \sreg_reg[1410]  ( .D(swire[390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1410]) );
  DFF \sreg_reg[1411]  ( .D(swire[391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1411]) );
  DFF \sreg_reg[1412]  ( .D(swire[392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1412]) );
  DFF \sreg_reg[1413]  ( .D(swire[393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1413]) );
  DFF \sreg_reg[1414]  ( .D(swire[394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1414]) );
  DFF \sreg_reg[1415]  ( .D(swire[395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1415]) );
  DFF \sreg_reg[1416]  ( .D(swire[396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1416]) );
  DFF \sreg_reg[1417]  ( .D(swire[397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1417]) );
  DFF \sreg_reg[1418]  ( .D(swire[398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1418]) );
  DFF \sreg_reg[1419]  ( .D(swire[399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1419]) );
  DFF \sreg_reg[1420]  ( .D(swire[400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1420]) );
  DFF \sreg_reg[1421]  ( .D(swire[401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1421]) );
  DFF \sreg_reg[1422]  ( .D(swire[402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1422]) );
  DFF \sreg_reg[1423]  ( .D(swire[403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1423]) );
  DFF \sreg_reg[1424]  ( .D(swire[404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1424]) );
  DFF \sreg_reg[1425]  ( .D(swire[405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1425]) );
  DFF \sreg_reg[1426]  ( .D(swire[406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1426]) );
  DFF \sreg_reg[1427]  ( .D(swire[407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1427]) );
  DFF \sreg_reg[1428]  ( .D(swire[408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1428]) );
  DFF \sreg_reg[1429]  ( .D(swire[409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1429]) );
  DFF \sreg_reg[1430]  ( .D(swire[410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1430]) );
  DFF \sreg_reg[1431]  ( .D(swire[411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1431]) );
  DFF \sreg_reg[1432]  ( .D(swire[412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1432]) );
  DFF \sreg_reg[1433]  ( .D(swire[413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1433]) );
  DFF \sreg_reg[1434]  ( .D(swire[414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1434]) );
  DFF \sreg_reg[1435]  ( .D(swire[415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1435]) );
  DFF \sreg_reg[1436]  ( .D(swire[416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1436]) );
  DFF \sreg_reg[1437]  ( .D(swire[417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1437]) );
  DFF \sreg_reg[1438]  ( .D(swire[418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1438]) );
  DFF \sreg_reg[1439]  ( .D(swire[419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1439]) );
  DFF \sreg_reg[1440]  ( .D(swire[420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1440]) );
  DFF \sreg_reg[1441]  ( .D(swire[421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1441]) );
  DFF \sreg_reg[1442]  ( .D(swire[422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1442]) );
  DFF \sreg_reg[1443]  ( .D(swire[423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1443]) );
  DFF \sreg_reg[1444]  ( .D(swire[424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1444]) );
  DFF \sreg_reg[1445]  ( .D(swire[425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1445]) );
  DFF \sreg_reg[1446]  ( .D(swire[426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1446]) );
  DFF \sreg_reg[1447]  ( .D(swire[427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1447]) );
  DFF \sreg_reg[1448]  ( .D(swire[428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1448]) );
  DFF \sreg_reg[1449]  ( .D(swire[429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1449]) );
  DFF \sreg_reg[1450]  ( .D(swire[430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1450]) );
  DFF \sreg_reg[1451]  ( .D(swire[431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1451]) );
  DFF \sreg_reg[1452]  ( .D(swire[432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1452]) );
  DFF \sreg_reg[1453]  ( .D(swire[433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1453]) );
  DFF \sreg_reg[1454]  ( .D(swire[434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1454]) );
  DFF \sreg_reg[1455]  ( .D(swire[435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1455]) );
  DFF \sreg_reg[1456]  ( .D(swire[436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1456]) );
  DFF \sreg_reg[1457]  ( .D(swire[437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1457]) );
  DFF \sreg_reg[1458]  ( .D(swire[438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1458]) );
  DFF \sreg_reg[1459]  ( .D(swire[439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1459]) );
  DFF \sreg_reg[1460]  ( .D(swire[440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1460]) );
  DFF \sreg_reg[1461]  ( .D(swire[441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1461]) );
  DFF \sreg_reg[1462]  ( .D(swire[442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1462]) );
  DFF \sreg_reg[1463]  ( .D(swire[443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1463]) );
  DFF \sreg_reg[1464]  ( .D(swire[444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1464]) );
  DFF \sreg_reg[1465]  ( .D(swire[445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1465]) );
  DFF \sreg_reg[1466]  ( .D(swire[446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1466]) );
  DFF \sreg_reg[1467]  ( .D(swire[447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1467]) );
  DFF \sreg_reg[1468]  ( .D(swire[448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1468]) );
  DFF \sreg_reg[1469]  ( .D(swire[449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1469]) );
  DFF \sreg_reg[1470]  ( .D(swire[450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1470]) );
  DFF \sreg_reg[1471]  ( .D(swire[451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1471]) );
  DFF \sreg_reg[1472]  ( .D(swire[452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1472]) );
  DFF \sreg_reg[1473]  ( .D(swire[453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1473]) );
  DFF \sreg_reg[1474]  ( .D(swire[454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1474]) );
  DFF \sreg_reg[1475]  ( .D(swire[455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1475]) );
  DFF \sreg_reg[1476]  ( .D(swire[456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1476]) );
  DFF \sreg_reg[1477]  ( .D(swire[457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1477]) );
  DFF \sreg_reg[1478]  ( .D(swire[458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1478]) );
  DFF \sreg_reg[1479]  ( .D(swire[459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1479]) );
  DFF \sreg_reg[1480]  ( .D(swire[460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1480]) );
  DFF \sreg_reg[1481]  ( .D(swire[461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1481]) );
  DFF \sreg_reg[1482]  ( .D(swire[462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1482]) );
  DFF \sreg_reg[1483]  ( .D(swire[463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1483]) );
  DFF \sreg_reg[1484]  ( .D(swire[464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1484]) );
  DFF \sreg_reg[1485]  ( .D(swire[465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1485]) );
  DFF \sreg_reg[1486]  ( .D(swire[466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1486]) );
  DFF \sreg_reg[1487]  ( .D(swire[467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1487]) );
  DFF \sreg_reg[1488]  ( .D(swire[468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1488]) );
  DFF \sreg_reg[1489]  ( .D(swire[469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1489]) );
  DFF \sreg_reg[1490]  ( .D(swire[470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1490]) );
  DFF \sreg_reg[1491]  ( .D(swire[471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1491]) );
  DFF \sreg_reg[1492]  ( .D(swire[472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1492]) );
  DFF \sreg_reg[1493]  ( .D(swire[473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1493]) );
  DFF \sreg_reg[1494]  ( .D(swire[474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1494]) );
  DFF \sreg_reg[1495]  ( .D(swire[475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1495]) );
  DFF \sreg_reg[1496]  ( .D(swire[476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1496]) );
  DFF \sreg_reg[1497]  ( .D(swire[477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1497]) );
  DFF \sreg_reg[1498]  ( .D(swire[478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1498]) );
  DFF \sreg_reg[1499]  ( .D(swire[479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1499]) );
  DFF \sreg_reg[1500]  ( .D(swire[480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1500]) );
  DFF \sreg_reg[1501]  ( .D(swire[481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1501]) );
  DFF \sreg_reg[1502]  ( .D(swire[482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1502]) );
  DFF \sreg_reg[1503]  ( .D(swire[483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1503]) );
  DFF \sreg_reg[1504]  ( .D(swire[484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1504]) );
  DFF \sreg_reg[1505]  ( .D(swire[485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1505]) );
  DFF \sreg_reg[1506]  ( .D(swire[486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1506]) );
  DFF \sreg_reg[1507]  ( .D(swire[487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1507]) );
  DFF \sreg_reg[1508]  ( .D(swire[488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1508]) );
  DFF \sreg_reg[1509]  ( .D(swire[489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1509]) );
  DFF \sreg_reg[1510]  ( .D(swire[490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1510]) );
  DFF \sreg_reg[1511]  ( .D(swire[491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1511]) );
  DFF \sreg_reg[1512]  ( .D(swire[492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1512]) );
  DFF \sreg_reg[1513]  ( .D(swire[493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1513]) );
  DFF \sreg_reg[1514]  ( .D(swire[494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1514]) );
  DFF \sreg_reg[1515]  ( .D(swire[495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1515]) );
  DFF \sreg_reg[1516]  ( .D(swire[496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1516]) );
  DFF \sreg_reg[1517]  ( .D(swire[497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1517]) );
  DFF \sreg_reg[1518]  ( .D(swire[498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1518]) );
  DFF \sreg_reg[1519]  ( .D(swire[499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1519]) );
  DFF \sreg_reg[1520]  ( .D(swire[500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1520]) );
  DFF \sreg_reg[1521]  ( .D(swire[501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1521]) );
  DFF \sreg_reg[1522]  ( .D(swire[502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1522]) );
  DFF \sreg_reg[1523]  ( .D(swire[503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1523]) );
  DFF \sreg_reg[1524]  ( .D(swire[504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1524]) );
  DFF \sreg_reg[1525]  ( .D(swire[505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1525]) );
  DFF \sreg_reg[1526]  ( .D(swire[506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1526]) );
  DFF \sreg_reg[1527]  ( .D(swire[507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1527]) );
  DFF \sreg_reg[1528]  ( .D(swire[508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1528]) );
  DFF \sreg_reg[1529]  ( .D(swire[509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1529]) );
  DFF \sreg_reg[1530]  ( .D(swire[510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1530]) );
  DFF \sreg_reg[1531]  ( .D(swire[511]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1531]) );
  DFF \sreg_reg[1532]  ( .D(swire[512]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1532]) );
  DFF \sreg_reg[1533]  ( .D(swire[513]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1533]) );
  DFF \sreg_reg[1534]  ( .D(swire[514]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1534]) );
  DFF \sreg_reg[1535]  ( .D(swire[515]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1535]) );
  DFF \sreg_reg[1536]  ( .D(swire[516]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1536]) );
  DFF \sreg_reg[1537]  ( .D(swire[517]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1537]) );
  DFF \sreg_reg[1538]  ( .D(swire[518]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1538]) );
  DFF \sreg_reg[1539]  ( .D(swire[519]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1539]) );
  DFF \sreg_reg[1540]  ( .D(swire[520]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1540]) );
  DFF \sreg_reg[1541]  ( .D(swire[521]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1541]) );
  DFF \sreg_reg[1542]  ( .D(swire[522]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1542]) );
  DFF \sreg_reg[1543]  ( .D(swire[523]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1543]) );
  DFF \sreg_reg[1544]  ( .D(swire[524]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1544]) );
  DFF \sreg_reg[1545]  ( .D(swire[525]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1545]) );
  DFF \sreg_reg[1546]  ( .D(swire[526]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1546]) );
  DFF \sreg_reg[1547]  ( .D(swire[527]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1547]) );
  DFF \sreg_reg[1548]  ( .D(swire[528]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1548]) );
  DFF \sreg_reg[1549]  ( .D(swire[529]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1549]) );
  DFF \sreg_reg[1550]  ( .D(swire[530]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1550]) );
  DFF \sreg_reg[1551]  ( .D(swire[531]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1551]) );
  DFF \sreg_reg[1552]  ( .D(swire[532]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1552]) );
  DFF \sreg_reg[1553]  ( .D(swire[533]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1553]) );
  DFF \sreg_reg[1554]  ( .D(swire[534]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1554]) );
  DFF \sreg_reg[1555]  ( .D(swire[535]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1555]) );
  DFF \sreg_reg[1556]  ( .D(swire[536]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1556]) );
  DFF \sreg_reg[1557]  ( .D(swire[537]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1557]) );
  DFF \sreg_reg[1558]  ( .D(swire[538]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1558]) );
  DFF \sreg_reg[1559]  ( .D(swire[539]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1559]) );
  DFF \sreg_reg[1560]  ( .D(swire[540]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1560]) );
  DFF \sreg_reg[1561]  ( .D(swire[541]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1561]) );
  DFF \sreg_reg[1562]  ( .D(swire[542]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1562]) );
  DFF \sreg_reg[1563]  ( .D(swire[543]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1563]) );
  DFF \sreg_reg[1564]  ( .D(swire[544]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1564]) );
  DFF \sreg_reg[1565]  ( .D(swire[545]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1565]) );
  DFF \sreg_reg[1566]  ( .D(swire[546]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1566]) );
  DFF \sreg_reg[1567]  ( .D(swire[547]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1567]) );
  DFF \sreg_reg[1568]  ( .D(swire[548]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1568]) );
  DFF \sreg_reg[1569]  ( .D(swire[549]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1569]) );
  DFF \sreg_reg[1570]  ( .D(swire[550]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1570]) );
  DFF \sreg_reg[1571]  ( .D(swire[551]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1571]) );
  DFF \sreg_reg[1572]  ( .D(swire[552]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1572]) );
  DFF \sreg_reg[1573]  ( .D(swire[553]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1573]) );
  DFF \sreg_reg[1574]  ( .D(swire[554]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1574]) );
  DFF \sreg_reg[1575]  ( .D(swire[555]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1575]) );
  DFF \sreg_reg[1576]  ( .D(swire[556]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1576]) );
  DFF \sreg_reg[1577]  ( .D(swire[557]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1577]) );
  DFF \sreg_reg[1578]  ( .D(swire[558]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1578]) );
  DFF \sreg_reg[1579]  ( .D(swire[559]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1579]) );
  DFF \sreg_reg[1580]  ( .D(swire[560]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1580]) );
  DFF \sreg_reg[1581]  ( .D(swire[561]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1581]) );
  DFF \sreg_reg[1582]  ( .D(swire[562]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1582]) );
  DFF \sreg_reg[1583]  ( .D(swire[563]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1583]) );
  DFF \sreg_reg[1584]  ( .D(swire[564]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1584]) );
  DFF \sreg_reg[1585]  ( .D(swire[565]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1585]) );
  DFF \sreg_reg[1586]  ( .D(swire[566]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1586]) );
  DFF \sreg_reg[1587]  ( .D(swire[567]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1587]) );
  DFF \sreg_reg[1588]  ( .D(swire[568]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1588]) );
  DFF \sreg_reg[1589]  ( .D(swire[569]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1589]) );
  DFF \sreg_reg[1590]  ( .D(swire[570]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1590]) );
  DFF \sreg_reg[1591]  ( .D(swire[571]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1591]) );
  DFF \sreg_reg[1592]  ( .D(swire[572]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1592]) );
  DFF \sreg_reg[1593]  ( .D(swire[573]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1593]) );
  DFF \sreg_reg[1594]  ( .D(swire[574]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1594]) );
  DFF \sreg_reg[1595]  ( .D(swire[575]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1595]) );
  DFF \sreg_reg[1596]  ( .D(swire[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1596]) );
  DFF \sreg_reg[1597]  ( .D(swire[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1597]) );
  DFF \sreg_reg[1598]  ( .D(swire[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1598]) );
  DFF \sreg_reg[1599]  ( .D(swire[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1599]) );
  DFF \sreg_reg[1600]  ( .D(swire[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1600]) );
  DFF \sreg_reg[1601]  ( .D(swire[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1601]) );
  DFF \sreg_reg[1602]  ( .D(swire[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1602]) );
  DFF \sreg_reg[1603]  ( .D(swire[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1603]) );
  DFF \sreg_reg[1604]  ( .D(swire[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1604]) );
  DFF \sreg_reg[1605]  ( .D(swire[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1605]) );
  DFF \sreg_reg[1606]  ( .D(swire[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1606]) );
  DFF \sreg_reg[1607]  ( .D(swire[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1607]) );
  DFF \sreg_reg[1608]  ( .D(swire[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1608]) );
  DFF \sreg_reg[1609]  ( .D(swire[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1609]) );
  DFF \sreg_reg[1610]  ( .D(swire[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1610]) );
  DFF \sreg_reg[1611]  ( .D(swire[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1611]) );
  DFF \sreg_reg[1612]  ( .D(swire[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1612]) );
  DFF \sreg_reg[1613]  ( .D(swire[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1613]) );
  DFF \sreg_reg[1614]  ( .D(swire[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1614]) );
  DFF \sreg_reg[1615]  ( .D(swire[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1615]) );
  DFF \sreg_reg[1616]  ( .D(swire[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1616]) );
  DFF \sreg_reg[1617]  ( .D(swire[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1617]) );
  DFF \sreg_reg[1618]  ( .D(swire[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1618]) );
  DFF \sreg_reg[1619]  ( .D(swire[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1619]) );
  DFF \sreg_reg[1620]  ( .D(swire[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1620]) );
  DFF \sreg_reg[1621]  ( .D(swire[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1621]) );
  DFF \sreg_reg[1622]  ( .D(swire[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1622]) );
  DFF \sreg_reg[1623]  ( .D(swire[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1623]) );
  DFF \sreg_reg[1624]  ( .D(swire[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1624]) );
  DFF \sreg_reg[1625]  ( .D(swire[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1625]) );
  DFF \sreg_reg[1626]  ( .D(swire[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1626]) );
  DFF \sreg_reg[1627]  ( .D(swire[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1627]) );
  DFF \sreg_reg[1628]  ( .D(swire[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1628]) );
  DFF \sreg_reg[1629]  ( .D(swire[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1629]) );
  DFF \sreg_reg[1630]  ( .D(swire[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1630]) );
  DFF \sreg_reg[1631]  ( .D(swire[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1631]) );
  DFF \sreg_reg[1632]  ( .D(swire[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1632]) );
  DFF \sreg_reg[1633]  ( .D(swire[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1633]) );
  DFF \sreg_reg[1634]  ( .D(swire[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1634]) );
  DFF \sreg_reg[1635]  ( .D(swire[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1635]) );
  DFF \sreg_reg[1636]  ( .D(swire[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1636]) );
  DFF \sreg_reg[1637]  ( .D(swire[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1637]) );
  DFF \sreg_reg[1638]  ( .D(swire[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1638]) );
  DFF \sreg_reg[1639]  ( .D(swire[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1639]) );
  DFF \sreg_reg[1640]  ( .D(swire[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1640]) );
  DFF \sreg_reg[1641]  ( .D(swire[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1641]) );
  DFF \sreg_reg[1642]  ( .D(swire[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1642]) );
  DFF \sreg_reg[1643]  ( .D(swire[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1643]) );
  DFF \sreg_reg[1644]  ( .D(swire[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1644]) );
  DFF \sreg_reg[1645]  ( .D(swire[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1645]) );
  DFF \sreg_reg[1646]  ( .D(swire[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1646]) );
  DFF \sreg_reg[1647]  ( .D(swire[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1647]) );
  DFF \sreg_reg[1648]  ( .D(swire[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1648]) );
  DFF \sreg_reg[1649]  ( .D(swire[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1649]) );
  DFF \sreg_reg[1650]  ( .D(swire[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1650]) );
  DFF \sreg_reg[1651]  ( .D(swire[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1651]) );
  DFF \sreg_reg[1652]  ( .D(swire[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1652]) );
  DFF \sreg_reg[1653]  ( .D(swire[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1653]) );
  DFF \sreg_reg[1654]  ( .D(swire[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1654]) );
  DFF \sreg_reg[1655]  ( .D(swire[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1655]) );
  DFF \sreg_reg[1656]  ( .D(swire[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1656]) );
  DFF \sreg_reg[1657]  ( .D(swire[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1657]) );
  DFF \sreg_reg[1658]  ( .D(swire[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1658]) );
  DFF \sreg_reg[1659]  ( .D(swire[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1659]) );
  DFF \sreg_reg[1660]  ( .D(swire[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1660]) );
  DFF \sreg_reg[1661]  ( .D(swire[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1661]) );
  DFF \sreg_reg[1662]  ( .D(swire[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1662]) );
  DFF \sreg_reg[1663]  ( .D(swire[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1663]) );
  DFF \sreg_reg[1664]  ( .D(swire[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1664]) );
  DFF \sreg_reg[1665]  ( .D(swire[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1665]) );
  DFF \sreg_reg[1666]  ( .D(swire[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1666]) );
  DFF \sreg_reg[1667]  ( .D(swire[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1667]) );
  DFF \sreg_reg[1668]  ( .D(swire[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1668]) );
  DFF \sreg_reg[1669]  ( .D(swire[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1669]) );
  DFF \sreg_reg[1670]  ( .D(swire[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1670]) );
  DFF \sreg_reg[1671]  ( .D(swire[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1671]) );
  DFF \sreg_reg[1672]  ( .D(swire[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1672]) );
  DFF \sreg_reg[1673]  ( .D(swire[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1673]) );
  DFF \sreg_reg[1674]  ( .D(swire[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1674]) );
  DFF \sreg_reg[1675]  ( .D(swire[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1675]) );
  DFF \sreg_reg[1676]  ( .D(swire[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1676]) );
  DFF \sreg_reg[1677]  ( .D(swire[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1677]) );
  DFF \sreg_reg[1678]  ( .D(swire[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1678]) );
  DFF \sreg_reg[1679]  ( .D(swire[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1679]) );
  DFF \sreg_reg[1680]  ( .D(swire[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1680]) );
  DFF \sreg_reg[1681]  ( .D(swire[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1681]) );
  DFF \sreg_reg[1682]  ( .D(swire[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1682]) );
  DFF \sreg_reg[1683]  ( .D(swire[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1683]) );
  DFF \sreg_reg[1684]  ( .D(swire[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1684]) );
  DFF \sreg_reg[1685]  ( .D(swire[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1685]) );
  DFF \sreg_reg[1686]  ( .D(swire[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1686]) );
  DFF \sreg_reg[1687]  ( .D(swire[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1687]) );
  DFF \sreg_reg[1688]  ( .D(swire[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1688]) );
  DFF \sreg_reg[1689]  ( .D(swire[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1689]) );
  DFF \sreg_reg[1690]  ( .D(swire[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1690]) );
  DFF \sreg_reg[1691]  ( .D(swire[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1691]) );
  DFF \sreg_reg[1692]  ( .D(swire[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1692]) );
  DFF \sreg_reg[1693]  ( .D(swire[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1693]) );
  DFF \sreg_reg[1694]  ( .D(swire[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1694]) );
  DFF \sreg_reg[1695]  ( .D(swire[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1695]) );
  DFF \sreg_reg[1696]  ( .D(swire[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1696]) );
  DFF \sreg_reg[1697]  ( .D(swire[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1697]) );
  DFF \sreg_reg[1698]  ( .D(swire[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1698]) );
  DFF \sreg_reg[1699]  ( .D(swire[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1699]) );
  DFF \sreg_reg[1700]  ( .D(swire[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1700]) );
  DFF \sreg_reg[1701]  ( .D(swire[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1701]) );
  DFF \sreg_reg[1702]  ( .D(swire[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1702]) );
  DFF \sreg_reg[1703]  ( .D(swire[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1703]) );
  DFF \sreg_reg[1704]  ( .D(swire[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1704]) );
  DFF \sreg_reg[1705]  ( .D(swire[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1705]) );
  DFF \sreg_reg[1706]  ( .D(swire[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1706]) );
  DFF \sreg_reg[1707]  ( .D(swire[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1707]) );
  DFF \sreg_reg[1708]  ( .D(swire[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1708]) );
  DFF \sreg_reg[1709]  ( .D(swire[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1709]) );
  DFF \sreg_reg[1710]  ( .D(swire[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1710]) );
  DFF \sreg_reg[1711]  ( .D(swire[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1711]) );
  DFF \sreg_reg[1712]  ( .D(swire[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1712]) );
  DFF \sreg_reg[1713]  ( .D(swire[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1713]) );
  DFF \sreg_reg[1714]  ( .D(swire[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1714]) );
  DFF \sreg_reg[1715]  ( .D(swire[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1715]) );
  DFF \sreg_reg[1716]  ( .D(swire[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1716]) );
  DFF \sreg_reg[1717]  ( .D(swire[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1717]) );
  DFF \sreg_reg[1718]  ( .D(swire[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1718]) );
  DFF \sreg_reg[1719]  ( .D(swire[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1719]) );
  DFF \sreg_reg[1720]  ( .D(swire[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1720]) );
  DFF \sreg_reg[1721]  ( .D(swire[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1721]) );
  DFF \sreg_reg[1722]  ( .D(swire[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1722]) );
  DFF \sreg_reg[1723]  ( .D(swire[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1723]) );
  DFF \sreg_reg[1724]  ( .D(swire[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1724]) );
  DFF \sreg_reg[1725]  ( .D(swire[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1725]) );
  DFF \sreg_reg[1726]  ( .D(swire[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1726]) );
  DFF \sreg_reg[1727]  ( .D(swire[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1727]) );
  DFF \sreg_reg[1728]  ( .D(swire[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1728]) );
  DFF \sreg_reg[1729]  ( .D(swire[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1729]) );
  DFF \sreg_reg[1730]  ( .D(swire[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1730]) );
  DFF \sreg_reg[1731]  ( .D(swire[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1731]) );
  DFF \sreg_reg[1732]  ( .D(swire[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1732]) );
  DFF \sreg_reg[1733]  ( .D(swire[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1733]) );
  DFF \sreg_reg[1734]  ( .D(swire[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1734]) );
  DFF \sreg_reg[1735]  ( .D(swire[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1735]) );
  DFF \sreg_reg[1736]  ( .D(swire[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1736]) );
  DFF \sreg_reg[1737]  ( .D(swire[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1737]) );
  DFF \sreg_reg[1738]  ( .D(swire[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1738]) );
  DFF \sreg_reg[1739]  ( .D(swire[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1739]) );
  DFF \sreg_reg[1740]  ( .D(swire[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1740]) );
  DFF \sreg_reg[1741]  ( .D(swire[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1741]) );
  DFF \sreg_reg[1742]  ( .D(swire[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1742]) );
  DFF \sreg_reg[1743]  ( .D(swire[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1743]) );
  DFF \sreg_reg[1744]  ( .D(swire[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1744]) );
  DFF \sreg_reg[1745]  ( .D(swire[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1745]) );
  DFF \sreg_reg[1746]  ( .D(swire[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1746]) );
  DFF \sreg_reg[1747]  ( .D(swire[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1747]) );
  DFF \sreg_reg[1748]  ( .D(swire[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1748]) );
  DFF \sreg_reg[1749]  ( .D(swire[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1749]) );
  DFF \sreg_reg[1750]  ( .D(swire[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1750]) );
  DFF \sreg_reg[1751]  ( .D(swire[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1751]) );
  DFF \sreg_reg[1752]  ( .D(swire[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1752]) );
  DFF \sreg_reg[1753]  ( .D(swire[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1753]) );
  DFF \sreg_reg[1754]  ( .D(swire[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1754]) );
  DFF \sreg_reg[1755]  ( .D(swire[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1755]) );
  DFF \sreg_reg[1756]  ( .D(swire[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1756]) );
  DFF \sreg_reg[1757]  ( .D(swire[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1757]) );
  DFF \sreg_reg[1758]  ( .D(swire[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1758]) );
  DFF \sreg_reg[1759]  ( .D(swire[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1759]) );
  DFF \sreg_reg[1760]  ( .D(swire[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1760]) );
  DFF \sreg_reg[1761]  ( .D(swire[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1761]) );
  DFF \sreg_reg[1762]  ( .D(swire[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1762]) );
  DFF \sreg_reg[1763]  ( .D(swire[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1763]) );
  DFF \sreg_reg[1764]  ( .D(swire[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1764]) );
  DFF \sreg_reg[1765]  ( .D(swire[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1765]) );
  DFF \sreg_reg[1766]  ( .D(swire[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1766]) );
  DFF \sreg_reg[1767]  ( .D(swire[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1767]) );
  DFF \sreg_reg[1768]  ( .D(swire[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1768]) );
  DFF \sreg_reg[1769]  ( .D(swire[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1769]) );
  DFF \sreg_reg[1770]  ( .D(swire[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1770]) );
  DFF \sreg_reg[1771]  ( .D(swire[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1771]) );
  DFF \sreg_reg[1772]  ( .D(swire[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1772]) );
  DFF \sreg_reg[1773]  ( .D(swire[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1773]) );
  DFF \sreg_reg[1774]  ( .D(swire[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1774]) );
  DFF \sreg_reg[1775]  ( .D(swire[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1775]) );
  DFF \sreg_reg[1776]  ( .D(swire[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1776]) );
  DFF \sreg_reg[1777]  ( .D(swire[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1777]) );
  DFF \sreg_reg[1778]  ( .D(swire[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1778]) );
  DFF \sreg_reg[1779]  ( .D(swire[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1779]) );
  DFF \sreg_reg[1780]  ( .D(swire[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1780]) );
  DFF \sreg_reg[1781]  ( .D(swire[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1781]) );
  DFF \sreg_reg[1782]  ( .D(swire[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1782]) );
  DFF \sreg_reg[1783]  ( .D(swire[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1783]) );
  DFF \sreg_reg[1784]  ( .D(swire[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1784]) );
  DFF \sreg_reg[1785]  ( .D(swire[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1785]) );
  DFF \sreg_reg[1786]  ( .D(swire[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1786]) );
  DFF \sreg_reg[1787]  ( .D(swire[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1787]) );
  DFF \sreg_reg[1788]  ( .D(swire[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1788]) );
  DFF \sreg_reg[1789]  ( .D(swire[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1789]) );
  DFF \sreg_reg[1790]  ( .D(swire[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1790]) );
  DFF \sreg_reg[1791]  ( .D(swire[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1791]) );
  DFF \sreg_reg[1792]  ( .D(swire[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1792]) );
  DFF \sreg_reg[1793]  ( .D(swire[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1793]) );
  DFF \sreg_reg[1794]  ( .D(swire[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1794]) );
  DFF \sreg_reg[1795]  ( .D(swire[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1795]) );
  DFF \sreg_reg[1796]  ( .D(swire[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1796]) );
  DFF \sreg_reg[1797]  ( .D(swire[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1797]) );
  DFF \sreg_reg[1798]  ( .D(swire[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1798]) );
  DFF \sreg_reg[1799]  ( .D(swire[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1799]) );
  DFF \sreg_reg[1800]  ( .D(swire[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1800]) );
  DFF \sreg_reg[1801]  ( .D(swire[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1801]) );
  DFF \sreg_reg[1802]  ( .D(swire[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1802]) );
  DFF \sreg_reg[1803]  ( .D(swire[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1803]) );
  DFF \sreg_reg[1804]  ( .D(swire[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1804]) );
  DFF \sreg_reg[1805]  ( .D(swire[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1805]) );
  DFF \sreg_reg[1806]  ( .D(swire[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1806]) );
  DFF \sreg_reg[1807]  ( .D(swire[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1807]) );
  DFF \sreg_reg[1808]  ( .D(swire[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1808]) );
  DFF \sreg_reg[1809]  ( .D(swire[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1809]) );
  DFF \sreg_reg[1810]  ( .D(swire[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1810]) );
  DFF \sreg_reg[1811]  ( .D(swire[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1811]) );
  DFF \sreg_reg[1812]  ( .D(swire[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1812]) );
  DFF \sreg_reg[1813]  ( .D(swire[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1813]) );
  DFF \sreg_reg[1814]  ( .D(swire[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1814]) );
  DFF \sreg_reg[1815]  ( .D(swire[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1815]) );
  DFF \sreg_reg[1816]  ( .D(swire[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1816]) );
  DFF \sreg_reg[1817]  ( .D(swire[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1817]) );
  DFF \sreg_reg[1818]  ( .D(swire[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1818]) );
  DFF \sreg_reg[1819]  ( .D(swire[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1819]) );
  DFF \sreg_reg[1820]  ( .D(swire[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1820]) );
  DFF \sreg_reg[1821]  ( .D(swire[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1821]) );
  DFF \sreg_reg[1822]  ( .D(swire[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1822]) );
  DFF \sreg_reg[1823]  ( .D(swire[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1823]) );
  DFF \sreg_reg[1824]  ( .D(swire[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1824]) );
  DFF \sreg_reg[1825]  ( .D(swire[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1825]) );
  DFF \sreg_reg[1826]  ( .D(swire[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1826]) );
  DFF \sreg_reg[1827]  ( .D(swire[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1827]) );
  DFF \sreg_reg[1828]  ( .D(swire[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1828]) );
  DFF \sreg_reg[1829]  ( .D(swire[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1829]) );
  DFF \sreg_reg[1830]  ( .D(swire[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1830]) );
  DFF \sreg_reg[1831]  ( .D(swire[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1831]) );
  DFF \sreg_reg[1832]  ( .D(swire[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1832]) );
  DFF \sreg_reg[1833]  ( .D(swire[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1833]) );
  DFF \sreg_reg[1834]  ( .D(swire[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1834]) );
  DFF \sreg_reg[1835]  ( .D(swire[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1835]) );
  DFF \sreg_reg[1836]  ( .D(swire[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1836]) );
  DFF \sreg_reg[1837]  ( .D(swire[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1837]) );
  DFF \sreg_reg[1838]  ( .D(swire[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1838]) );
  DFF \sreg_reg[1839]  ( .D(swire[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1839]) );
  DFF \sreg_reg[1840]  ( .D(swire[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1840]) );
  DFF \sreg_reg[1841]  ( .D(swire[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1841]) );
  DFF \sreg_reg[1842]  ( .D(swire[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1842]) );
  DFF \sreg_reg[1843]  ( .D(swire[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1843]) );
  DFF \sreg_reg[1844]  ( .D(swire[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1844]) );
  DFF \sreg_reg[1845]  ( .D(swire[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1845]) );
  DFF \sreg_reg[1846]  ( .D(swire[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1846]) );
  DFF \sreg_reg[1847]  ( .D(swire[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1847]) );
  DFF \sreg_reg[1848]  ( .D(swire[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1848]) );
  DFF \sreg_reg[1849]  ( .D(swire[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1849]) );
  DFF \sreg_reg[1850]  ( .D(swire[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1850]) );
  DFF \sreg_reg[1851]  ( .D(swire[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1851]) );
  DFF \sreg_reg[1852]  ( .D(swire[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1852]) );
  DFF \sreg_reg[1853]  ( .D(swire[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1853]) );
  DFF \sreg_reg[1854]  ( .D(swire[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1854]) );
  DFF \sreg_reg[1855]  ( .D(swire[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1855]) );
  DFF \sreg_reg[1856]  ( .D(swire[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1856]) );
  DFF \sreg_reg[1857]  ( .D(swire[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1857]) );
  DFF \sreg_reg[1858]  ( .D(swire[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1858]) );
  DFF \sreg_reg[1859]  ( .D(swire[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1859]) );
  DFF \sreg_reg[1860]  ( .D(swire[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1860]) );
  DFF \sreg_reg[1861]  ( .D(swire[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1861]) );
  DFF \sreg_reg[1862]  ( .D(swire[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1862]) );
  DFF \sreg_reg[1863]  ( .D(swire[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1863]) );
  DFF \sreg_reg[1864]  ( .D(swire[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1864]) );
  DFF \sreg_reg[1865]  ( .D(swire[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1865]) );
  DFF \sreg_reg[1866]  ( .D(swire[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1866]) );
  DFF \sreg_reg[1867]  ( .D(swire[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1867]) );
  DFF \sreg_reg[1868]  ( .D(swire[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1868]) );
  DFF \sreg_reg[1869]  ( .D(swire[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1869]) );
  DFF \sreg_reg[1870]  ( .D(swire[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1870]) );
  DFF \sreg_reg[1871]  ( .D(swire[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1871]) );
  DFF \sreg_reg[1872]  ( .D(swire[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1872]) );
  DFF \sreg_reg[1873]  ( .D(swire[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1873]) );
  DFF \sreg_reg[1874]  ( .D(swire[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1874]) );
  DFF \sreg_reg[1875]  ( .D(swire[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1875]) );
  DFF \sreg_reg[1876]  ( .D(swire[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1876]) );
  DFF \sreg_reg[1877]  ( .D(swire[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1877]) );
  DFF \sreg_reg[1878]  ( .D(swire[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1878]) );
  DFF \sreg_reg[1879]  ( .D(swire[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1879]) );
  DFF \sreg_reg[1880]  ( .D(swire[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1880]) );
  DFF \sreg_reg[1881]  ( .D(swire[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1881]) );
  DFF \sreg_reg[1882]  ( .D(swire[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1882]) );
  DFF \sreg_reg[1883]  ( .D(swire[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1883]) );
  DFF \sreg_reg[1884]  ( .D(swire[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1884]) );
  DFF \sreg_reg[1885]  ( .D(swire[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1885]) );
  DFF \sreg_reg[1886]  ( .D(swire[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1886]) );
  DFF \sreg_reg[1887]  ( .D(swire[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1887]) );
  DFF \sreg_reg[1888]  ( .D(swire[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1888]) );
  DFF \sreg_reg[1889]  ( .D(swire[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1889]) );
  DFF \sreg_reg[1890]  ( .D(swire[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1890]) );
  DFF \sreg_reg[1891]  ( .D(swire[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1891]) );
  DFF \sreg_reg[1892]  ( .D(swire[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1892]) );
  DFF \sreg_reg[1893]  ( .D(swire[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1893]) );
  DFF \sreg_reg[1894]  ( .D(swire[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1894]) );
  DFF \sreg_reg[1895]  ( .D(swire[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1895]) );
  DFF \sreg_reg[1896]  ( .D(swire[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1896]) );
  DFF \sreg_reg[1897]  ( .D(swire[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1897]) );
  DFF \sreg_reg[1898]  ( .D(swire[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1898]) );
  DFF \sreg_reg[1899]  ( .D(swire[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1899]) );
  DFF \sreg_reg[1900]  ( .D(swire[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1900]) );
  DFF \sreg_reg[1901]  ( .D(swire[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1901]) );
  DFF \sreg_reg[1902]  ( .D(swire[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1902]) );
  DFF \sreg_reg[1903]  ( .D(swire[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1903]) );
  DFF \sreg_reg[1904]  ( .D(swire[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1904]) );
  DFF \sreg_reg[1905]  ( .D(swire[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1905]) );
  DFF \sreg_reg[1906]  ( .D(swire[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1906]) );
  DFF \sreg_reg[1907]  ( .D(swire[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1907]) );
  DFF \sreg_reg[1908]  ( .D(swire[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1908]) );
  DFF \sreg_reg[1909]  ( .D(swire[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1909]) );
  DFF \sreg_reg[1910]  ( .D(swire[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1910]) );
  DFF \sreg_reg[1911]  ( .D(swire[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1911]) );
  DFF \sreg_reg[1912]  ( .D(swire[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1912]) );
  DFF \sreg_reg[1913]  ( .D(swire[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1913]) );
  DFF \sreg_reg[1914]  ( .D(swire[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1914]) );
  DFF \sreg_reg[1915]  ( .D(swire[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1915]) );
  DFF \sreg_reg[1916]  ( .D(swire[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1916]) );
  DFF \sreg_reg[1917]  ( .D(swire[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1917]) );
  DFF \sreg_reg[1918]  ( .D(swire[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1918]) );
  DFF \sreg_reg[1919]  ( .D(swire[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1919]) );
  DFF \sreg_reg[1920]  ( .D(swire[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1920]) );
  DFF \sreg_reg[1921]  ( .D(swire[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1921]) );
  DFF \sreg_reg[1922]  ( .D(swire[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1922]) );
  DFF \sreg_reg[1923]  ( .D(swire[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1923]) );
  DFF \sreg_reg[1924]  ( .D(swire[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1924]) );
  DFF \sreg_reg[1925]  ( .D(swire[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1925]) );
  DFF \sreg_reg[1926]  ( .D(swire[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1926]) );
  DFF \sreg_reg[1927]  ( .D(swire[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1927]) );
  DFF \sreg_reg[1928]  ( .D(swire[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1928]) );
  DFF \sreg_reg[1929]  ( .D(swire[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1929]) );
  DFF \sreg_reg[1930]  ( .D(swire[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1930]) );
  DFF \sreg_reg[1931]  ( .D(swire[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1931]) );
  DFF \sreg_reg[1932]  ( .D(swire[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1932]) );
  DFF \sreg_reg[1933]  ( .D(swire[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1933]) );
  DFF \sreg_reg[1934]  ( .D(swire[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1934]) );
  DFF \sreg_reg[1935]  ( .D(swire[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1935]) );
  DFF \sreg_reg[1936]  ( .D(swire[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1936]) );
  DFF \sreg_reg[1937]  ( .D(swire[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1937]) );
  DFF \sreg_reg[1938]  ( .D(swire[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1938]) );
  DFF \sreg_reg[1939]  ( .D(swire[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1939]) );
  DFF \sreg_reg[1940]  ( .D(swire[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1940]) );
  DFF \sreg_reg[1941]  ( .D(swire[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1941]) );
  DFF \sreg_reg[1942]  ( .D(swire[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1942]) );
  DFF \sreg_reg[1943]  ( .D(swire[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1943]) );
  DFF \sreg_reg[1944]  ( .D(swire[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1944]) );
  DFF \sreg_reg[1945]  ( .D(swire[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1945]) );
  DFF \sreg_reg[1946]  ( .D(swire[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1946]) );
  DFF \sreg_reg[1947]  ( .D(swire[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1947]) );
  DFF \sreg_reg[1948]  ( .D(swire[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1948]) );
  DFF \sreg_reg[1949]  ( .D(swire[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1949]) );
  DFF \sreg_reg[1950]  ( .D(swire[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1950]) );
  DFF \sreg_reg[1951]  ( .D(swire[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1951]) );
  DFF \sreg_reg[1952]  ( .D(swire[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1952]) );
  DFF \sreg_reg[1953]  ( .D(swire[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1953]) );
  DFF \sreg_reg[1954]  ( .D(swire[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1954]) );
  DFF \sreg_reg[1955]  ( .D(swire[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1955]) );
  DFF \sreg_reg[1956]  ( .D(swire[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1956]) );
  DFF \sreg_reg[1957]  ( .D(swire[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1957]) );
  DFF \sreg_reg[1958]  ( .D(swire[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1958]) );
  DFF \sreg_reg[1959]  ( .D(swire[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1959]) );
  DFF \sreg_reg[1960]  ( .D(swire[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1960]) );
  DFF \sreg_reg[1961]  ( .D(swire[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1961]) );
  DFF \sreg_reg[1962]  ( .D(swire[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1962]) );
  DFF \sreg_reg[1963]  ( .D(swire[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1963]) );
  DFF \sreg_reg[1964]  ( .D(swire[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1964]) );
  DFF \sreg_reg[1965]  ( .D(swire[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1965]) );
  DFF \sreg_reg[1966]  ( .D(swire[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1966]) );
  DFF \sreg_reg[1967]  ( .D(swire[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1967]) );
  DFF \sreg_reg[1968]  ( .D(swire[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1968]) );
  DFF \sreg_reg[1969]  ( .D(swire[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1969]) );
  DFF \sreg_reg[1970]  ( .D(swire[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1970]) );
  DFF \sreg_reg[1971]  ( .D(swire[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1971]) );
  DFF \sreg_reg[1972]  ( .D(swire[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1972]) );
  DFF \sreg_reg[1973]  ( .D(swire[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1973]) );
  DFF \sreg_reg[1974]  ( .D(swire[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1974]) );
  DFF \sreg_reg[1975]  ( .D(swire[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1975]) );
  DFF \sreg_reg[1976]  ( .D(swire[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1976]) );
  DFF \sreg_reg[1977]  ( .D(swire[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1977]) );
  DFF \sreg_reg[1978]  ( .D(swire[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1978]) );
  DFF \sreg_reg[1979]  ( .D(swire[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1979]) );
  DFF \sreg_reg[1980]  ( .D(swire[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1980]) );
  DFF \sreg_reg[1981]  ( .D(swire[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1981]) );
  DFF \sreg_reg[1982]  ( .D(swire[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1982]) );
  DFF \sreg_reg[1983]  ( .D(swire[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1983]) );
  DFF \sreg_reg[1984]  ( .D(swire[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1984]) );
  DFF \sreg_reg[1985]  ( .D(swire[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1985]) );
  DFF \sreg_reg[1986]  ( .D(swire[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1986]) );
  DFF \sreg_reg[1987]  ( .D(swire[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1987]) );
  DFF \sreg_reg[1988]  ( .D(swire[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1988]) );
  DFF \sreg_reg[1989]  ( .D(swire[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1989]) );
  DFF \sreg_reg[1990]  ( .D(swire[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1990]) );
  DFF \sreg_reg[1991]  ( .D(swire[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1991]) );
  DFF \sreg_reg[1992]  ( .D(swire[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1992]) );
  DFF \sreg_reg[1993]  ( .D(swire[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1993]) );
  DFF \sreg_reg[1994]  ( .D(swire[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1994]) );
  DFF \sreg_reg[1995]  ( .D(swire[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1995]) );
  DFF \sreg_reg[1996]  ( .D(swire[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1996]) );
  DFF \sreg_reg[1997]  ( .D(swire[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1997]) );
  DFF \sreg_reg[1998]  ( .D(swire[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1998]) );
  DFF \sreg_reg[1999]  ( .D(swire[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[1999]) );
  DFF \sreg_reg[2000]  ( .D(swire[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2000]) );
  DFF \sreg_reg[2001]  ( .D(swire[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2001]) );
  DFF \sreg_reg[2002]  ( .D(swire[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2002]) );
  DFF \sreg_reg[2003]  ( .D(swire[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2003]) );
  DFF \sreg_reg[2004]  ( .D(swire[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2004]) );
  DFF \sreg_reg[2005]  ( .D(swire[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2005]) );
  DFF \sreg_reg[2006]  ( .D(swire[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2006]) );
  DFF \sreg_reg[2007]  ( .D(swire[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2007]) );
  DFF \sreg_reg[2008]  ( .D(swire[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2008]) );
  DFF \sreg_reg[2009]  ( .D(swire[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2009]) );
  DFF \sreg_reg[2010]  ( .D(swire[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2010]) );
  DFF \sreg_reg[2011]  ( .D(swire[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2011]) );
  DFF \sreg_reg[2012]  ( .D(swire[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2012]) );
  DFF \sreg_reg[2013]  ( .D(swire[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2013]) );
  DFF \sreg_reg[2014]  ( .D(swire[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2014]) );
  DFF \sreg_reg[2015]  ( .D(swire[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2015]) );
  DFF \sreg_reg[2016]  ( .D(swire[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2016]) );
  DFF \sreg_reg[2017]  ( .D(swire[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2017]) );
  DFF \sreg_reg[2018]  ( .D(swire[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2018]) );
  DFF \sreg_reg[2019]  ( .D(swire[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2019]) );
  DFF \sreg_reg[2020]  ( .D(swire[1000]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2020]) );
  DFF \sreg_reg[2021]  ( .D(swire[1001]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2021]) );
  DFF \sreg_reg[2022]  ( .D(swire[1002]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2022]) );
  DFF \sreg_reg[2023]  ( .D(swire[1003]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2023]) );
  DFF \sreg_reg[2024]  ( .D(swire[1004]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2024]) );
  DFF \sreg_reg[2025]  ( .D(swire[1005]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2025]) );
  DFF \sreg_reg[2026]  ( .D(swire[1006]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2026]) );
  DFF \sreg_reg[2027]  ( .D(swire[1007]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2027]) );
  DFF \sreg_reg[2028]  ( .D(swire[1008]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2028]) );
  DFF \sreg_reg[2029]  ( .D(swire[1009]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2029]) );
  DFF \sreg_reg[2030]  ( .D(swire[1010]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2030]) );
  DFF \sreg_reg[2031]  ( .D(swire[1011]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2031]) );
  DFF \sreg_reg[2032]  ( .D(swire[1012]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2032]) );
  DFF \sreg_reg[2033]  ( .D(swire[1013]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2033]) );
  DFF \sreg_reg[2034]  ( .D(swire[1014]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2034]) );
  DFF \sreg_reg[2035]  ( .D(swire[1015]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2035]) );
  DFF \sreg_reg[2036]  ( .D(swire[1016]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2036]) );
  DFF \sreg_reg[2037]  ( .D(swire[1017]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2037]) );
  DFF \sreg_reg[2038]  ( .D(swire[1018]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2038]) );
  DFF \sreg_reg[2039]  ( .D(swire[1019]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2039]) );
  DFF \sreg_reg[2040]  ( .D(swire[1020]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2040]) );
  DFF \sreg_reg[2041]  ( .D(swire[1021]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2041]) );
  DFF \sreg_reg[2042]  ( .D(swire[1022]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2042]) );
  DFF \sreg_reg[2043]  ( .D(swire[1023]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        sreg[2043]) );
  DFF \sreg_reg[1023]  ( .D(c[1023]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1019]) );
  DFF \sreg_reg[1022]  ( .D(c[1022]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1018]) );
  DFF \sreg_reg[1021]  ( .D(c[1021]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1017]) );
  DFF \sreg_reg[1020]  ( .D(c[1020]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1016]) );
  DFF \sreg_reg[1019]  ( .D(c[1019]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1015]) );
  DFF \sreg_reg[1018]  ( .D(c[1018]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1014]) );
  DFF \sreg_reg[1017]  ( .D(c[1017]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1013]) );
  DFF \sreg_reg[1016]  ( .D(c[1016]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1012]) );
  DFF \sreg_reg[1015]  ( .D(c[1015]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1011]) );
  DFF \sreg_reg[1014]  ( .D(c[1014]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1010]) );
  DFF \sreg_reg[1013]  ( .D(c[1013]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1009]) );
  DFF \sreg_reg[1012]  ( .D(c[1012]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1008]) );
  DFF \sreg_reg[1011]  ( .D(c[1011]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1007]) );
  DFF \sreg_reg[1010]  ( .D(c[1010]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1006]) );
  DFF \sreg_reg[1009]  ( .D(c[1009]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1005]) );
  DFF \sreg_reg[1008]  ( .D(c[1008]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1004]) );
  DFF \sreg_reg[1007]  ( .D(c[1007]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1003]) );
  DFF \sreg_reg[1006]  ( .D(c[1006]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1002]) );
  DFF \sreg_reg[1005]  ( .D(c[1005]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1001]) );
  DFF \sreg_reg[1004]  ( .D(c[1004]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[1000]) );
  DFF \sreg_reg[1003]  ( .D(c[1003]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[999]) );
  DFF \sreg_reg[1002]  ( .D(c[1002]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[998]) );
  DFF \sreg_reg[1001]  ( .D(c[1001]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[997]) );
  DFF \sreg_reg[1000]  ( .D(c[1000]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        c[996]) );
  DFF \sreg_reg[999]  ( .D(c[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[995])
         );
  DFF \sreg_reg[998]  ( .D(c[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[994])
         );
  DFF \sreg_reg[997]  ( .D(c[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[993])
         );
  DFF \sreg_reg[996]  ( .D(c[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[992])
         );
  DFF \sreg_reg[995]  ( .D(c[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[991])
         );
  DFF \sreg_reg[994]  ( .D(c[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[990])
         );
  DFF \sreg_reg[993]  ( .D(c[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[989])
         );
  DFF \sreg_reg[992]  ( .D(c[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[988])
         );
  DFF \sreg_reg[991]  ( .D(c[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[987])
         );
  DFF \sreg_reg[990]  ( .D(c[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[986])
         );
  DFF \sreg_reg[989]  ( .D(c[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[985])
         );
  DFF \sreg_reg[988]  ( .D(c[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[984])
         );
  DFF \sreg_reg[987]  ( .D(c[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[983])
         );
  DFF \sreg_reg[986]  ( .D(c[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[982])
         );
  DFF \sreg_reg[985]  ( .D(c[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[981])
         );
  DFF \sreg_reg[984]  ( .D(c[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[980])
         );
  DFF \sreg_reg[983]  ( .D(c[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[979])
         );
  DFF \sreg_reg[982]  ( .D(c[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[978])
         );
  DFF \sreg_reg[981]  ( .D(c[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[977])
         );
  DFF \sreg_reg[980]  ( .D(c[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[976])
         );
  DFF \sreg_reg[979]  ( .D(c[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[975])
         );
  DFF \sreg_reg[978]  ( .D(c[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[974])
         );
  DFF \sreg_reg[977]  ( .D(c[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[973])
         );
  DFF \sreg_reg[976]  ( .D(c[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[972])
         );
  DFF \sreg_reg[975]  ( .D(c[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[971])
         );
  DFF \sreg_reg[974]  ( .D(c[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[970])
         );
  DFF \sreg_reg[973]  ( .D(c[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[969])
         );
  DFF \sreg_reg[972]  ( .D(c[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[968])
         );
  DFF \sreg_reg[971]  ( .D(c[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[967])
         );
  DFF \sreg_reg[970]  ( .D(c[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[966])
         );
  DFF \sreg_reg[969]  ( .D(c[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[965])
         );
  DFF \sreg_reg[968]  ( .D(c[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[964])
         );
  DFF \sreg_reg[967]  ( .D(c[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[963])
         );
  DFF \sreg_reg[966]  ( .D(c[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[962])
         );
  DFF \sreg_reg[965]  ( .D(c[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[961])
         );
  DFF \sreg_reg[964]  ( .D(c[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[960])
         );
  DFF \sreg_reg[963]  ( .D(c[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[959])
         );
  DFF \sreg_reg[962]  ( .D(c[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[958])
         );
  DFF \sreg_reg[961]  ( .D(c[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[957])
         );
  DFF \sreg_reg[960]  ( .D(c[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[956])
         );
  DFF \sreg_reg[959]  ( .D(c[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[955])
         );
  DFF \sreg_reg[958]  ( .D(c[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[954])
         );
  DFF \sreg_reg[957]  ( .D(c[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[953])
         );
  DFF \sreg_reg[956]  ( .D(c[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[952])
         );
  DFF \sreg_reg[955]  ( .D(c[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[951])
         );
  DFF \sreg_reg[954]  ( .D(c[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[950])
         );
  DFF \sreg_reg[953]  ( .D(c[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[949])
         );
  DFF \sreg_reg[952]  ( .D(c[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[948])
         );
  DFF \sreg_reg[951]  ( .D(c[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[947])
         );
  DFF \sreg_reg[950]  ( .D(c[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[946])
         );
  DFF \sreg_reg[949]  ( .D(c[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[945])
         );
  DFF \sreg_reg[948]  ( .D(c[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[944])
         );
  DFF \sreg_reg[947]  ( .D(c[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[943])
         );
  DFF \sreg_reg[946]  ( .D(c[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[942])
         );
  DFF \sreg_reg[945]  ( .D(c[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[941])
         );
  DFF \sreg_reg[944]  ( .D(c[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[940])
         );
  DFF \sreg_reg[943]  ( .D(c[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[939])
         );
  DFF \sreg_reg[942]  ( .D(c[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[938])
         );
  DFF \sreg_reg[941]  ( .D(c[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[937])
         );
  DFF \sreg_reg[940]  ( .D(c[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[936])
         );
  DFF \sreg_reg[939]  ( .D(c[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[935])
         );
  DFF \sreg_reg[938]  ( .D(c[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[934])
         );
  DFF \sreg_reg[937]  ( .D(c[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[933])
         );
  DFF \sreg_reg[936]  ( .D(c[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[932])
         );
  DFF \sreg_reg[935]  ( .D(c[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[931])
         );
  DFF \sreg_reg[934]  ( .D(c[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[930])
         );
  DFF \sreg_reg[933]  ( .D(c[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[929])
         );
  DFF \sreg_reg[932]  ( .D(c[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[928])
         );
  DFF \sreg_reg[931]  ( .D(c[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[927])
         );
  DFF \sreg_reg[930]  ( .D(c[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[926])
         );
  DFF \sreg_reg[929]  ( .D(c[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[925])
         );
  DFF \sreg_reg[928]  ( .D(c[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[924])
         );
  DFF \sreg_reg[927]  ( .D(c[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[923])
         );
  DFF \sreg_reg[926]  ( .D(c[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[922])
         );
  DFF \sreg_reg[925]  ( .D(c[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[921])
         );
  DFF \sreg_reg[924]  ( .D(c[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[920])
         );
  DFF \sreg_reg[923]  ( .D(c[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[919])
         );
  DFF \sreg_reg[922]  ( .D(c[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[918])
         );
  DFF \sreg_reg[921]  ( .D(c[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[917])
         );
  DFF \sreg_reg[920]  ( .D(c[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[916])
         );
  DFF \sreg_reg[919]  ( .D(c[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[915])
         );
  DFF \sreg_reg[918]  ( .D(c[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[914])
         );
  DFF \sreg_reg[917]  ( .D(c[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[913])
         );
  DFF \sreg_reg[916]  ( .D(c[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[912])
         );
  DFF \sreg_reg[915]  ( .D(c[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[911])
         );
  DFF \sreg_reg[914]  ( .D(c[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[910])
         );
  DFF \sreg_reg[913]  ( .D(c[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[909])
         );
  DFF \sreg_reg[912]  ( .D(c[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[908])
         );
  DFF \sreg_reg[911]  ( .D(c[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[907])
         );
  DFF \sreg_reg[910]  ( .D(c[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[906])
         );
  DFF \sreg_reg[909]  ( .D(c[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[905])
         );
  DFF \sreg_reg[908]  ( .D(c[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[904])
         );
  DFF \sreg_reg[907]  ( .D(c[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[903])
         );
  DFF \sreg_reg[906]  ( .D(c[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[902])
         );
  DFF \sreg_reg[905]  ( .D(c[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[901])
         );
  DFF \sreg_reg[904]  ( .D(c[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[900])
         );
  DFF \sreg_reg[903]  ( .D(c[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[899])
         );
  DFF \sreg_reg[902]  ( .D(c[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[898])
         );
  DFF \sreg_reg[901]  ( .D(c[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[897])
         );
  DFF \sreg_reg[900]  ( .D(c[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[896])
         );
  DFF \sreg_reg[899]  ( .D(c[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[895])
         );
  DFF \sreg_reg[898]  ( .D(c[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[894])
         );
  DFF \sreg_reg[897]  ( .D(c[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[893])
         );
  DFF \sreg_reg[896]  ( .D(c[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[892])
         );
  DFF \sreg_reg[895]  ( .D(c[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[891])
         );
  DFF \sreg_reg[894]  ( .D(c[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[890])
         );
  DFF \sreg_reg[893]  ( .D(c[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[889])
         );
  DFF \sreg_reg[892]  ( .D(c[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[888])
         );
  DFF \sreg_reg[891]  ( .D(c[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[887])
         );
  DFF \sreg_reg[890]  ( .D(c[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[886])
         );
  DFF \sreg_reg[889]  ( .D(c[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[885])
         );
  DFF \sreg_reg[888]  ( .D(c[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[884])
         );
  DFF \sreg_reg[887]  ( .D(c[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[883])
         );
  DFF \sreg_reg[886]  ( .D(c[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[882])
         );
  DFF \sreg_reg[885]  ( .D(c[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[881])
         );
  DFF \sreg_reg[884]  ( .D(c[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[880])
         );
  DFF \sreg_reg[883]  ( .D(c[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[879])
         );
  DFF \sreg_reg[882]  ( .D(c[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[878])
         );
  DFF \sreg_reg[881]  ( .D(c[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[877])
         );
  DFF \sreg_reg[880]  ( .D(c[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[876])
         );
  DFF \sreg_reg[879]  ( .D(c[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[875])
         );
  DFF \sreg_reg[878]  ( .D(c[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[874])
         );
  DFF \sreg_reg[877]  ( .D(c[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[873])
         );
  DFF \sreg_reg[876]  ( .D(c[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[872])
         );
  DFF \sreg_reg[875]  ( .D(c[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[871])
         );
  DFF \sreg_reg[874]  ( .D(c[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[870])
         );
  DFF \sreg_reg[873]  ( .D(c[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[869])
         );
  DFF \sreg_reg[872]  ( .D(c[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[868])
         );
  DFF \sreg_reg[871]  ( .D(c[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[867])
         );
  DFF \sreg_reg[870]  ( .D(c[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[866])
         );
  DFF \sreg_reg[869]  ( .D(c[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[865])
         );
  DFF \sreg_reg[868]  ( .D(c[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[864])
         );
  DFF \sreg_reg[867]  ( .D(c[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[863])
         );
  DFF \sreg_reg[866]  ( .D(c[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[862])
         );
  DFF \sreg_reg[865]  ( .D(c[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[861])
         );
  DFF \sreg_reg[864]  ( .D(c[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[860])
         );
  DFF \sreg_reg[863]  ( .D(c[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[859])
         );
  DFF \sreg_reg[862]  ( .D(c[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[858])
         );
  DFF \sreg_reg[861]  ( .D(c[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[857])
         );
  DFF \sreg_reg[860]  ( .D(c[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[856])
         );
  DFF \sreg_reg[859]  ( .D(c[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[855])
         );
  DFF \sreg_reg[858]  ( .D(c[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[854])
         );
  DFF \sreg_reg[857]  ( .D(c[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[853])
         );
  DFF \sreg_reg[856]  ( .D(c[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[852])
         );
  DFF \sreg_reg[855]  ( .D(c[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[851])
         );
  DFF \sreg_reg[854]  ( .D(c[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[850])
         );
  DFF \sreg_reg[853]  ( .D(c[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[849])
         );
  DFF \sreg_reg[852]  ( .D(c[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[848])
         );
  DFF \sreg_reg[851]  ( .D(c[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[847])
         );
  DFF \sreg_reg[850]  ( .D(c[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[846])
         );
  DFF \sreg_reg[849]  ( .D(c[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[845])
         );
  DFF \sreg_reg[848]  ( .D(c[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[844])
         );
  DFF \sreg_reg[847]  ( .D(c[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[843])
         );
  DFF \sreg_reg[846]  ( .D(c[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[842])
         );
  DFF \sreg_reg[845]  ( .D(c[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[841])
         );
  DFF \sreg_reg[844]  ( .D(c[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[840])
         );
  DFF \sreg_reg[843]  ( .D(c[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[839])
         );
  DFF \sreg_reg[842]  ( .D(c[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[838])
         );
  DFF \sreg_reg[841]  ( .D(c[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[837])
         );
  DFF \sreg_reg[840]  ( .D(c[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[836])
         );
  DFF \sreg_reg[839]  ( .D(c[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[835])
         );
  DFF \sreg_reg[838]  ( .D(c[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[834])
         );
  DFF \sreg_reg[837]  ( .D(c[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[833])
         );
  DFF \sreg_reg[836]  ( .D(c[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[832])
         );
  DFF \sreg_reg[835]  ( .D(c[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[831])
         );
  DFF \sreg_reg[834]  ( .D(c[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[830])
         );
  DFF \sreg_reg[833]  ( .D(c[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[829])
         );
  DFF \sreg_reg[832]  ( .D(c[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[828])
         );
  DFF \sreg_reg[831]  ( .D(c[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[827])
         );
  DFF \sreg_reg[830]  ( .D(c[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[826])
         );
  DFF \sreg_reg[829]  ( .D(c[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[825])
         );
  DFF \sreg_reg[828]  ( .D(c[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[824])
         );
  DFF \sreg_reg[827]  ( .D(c[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[823])
         );
  DFF \sreg_reg[826]  ( .D(c[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[822])
         );
  DFF \sreg_reg[825]  ( .D(c[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[821])
         );
  DFF \sreg_reg[824]  ( .D(c[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[820])
         );
  DFF \sreg_reg[823]  ( .D(c[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[819])
         );
  DFF \sreg_reg[822]  ( .D(c[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[818])
         );
  DFF \sreg_reg[821]  ( .D(c[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[817])
         );
  DFF \sreg_reg[820]  ( .D(c[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[816])
         );
  DFF \sreg_reg[819]  ( .D(c[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[815])
         );
  DFF \sreg_reg[818]  ( .D(c[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[814])
         );
  DFF \sreg_reg[817]  ( .D(c[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[813])
         );
  DFF \sreg_reg[816]  ( .D(c[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[812])
         );
  DFF \sreg_reg[815]  ( .D(c[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[811])
         );
  DFF \sreg_reg[814]  ( .D(c[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[810])
         );
  DFF \sreg_reg[813]  ( .D(c[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[809])
         );
  DFF \sreg_reg[812]  ( .D(c[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[808])
         );
  DFF \sreg_reg[811]  ( .D(c[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[807])
         );
  DFF \sreg_reg[810]  ( .D(c[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[806])
         );
  DFF \sreg_reg[809]  ( .D(c[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[805])
         );
  DFF \sreg_reg[808]  ( .D(c[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[804])
         );
  DFF \sreg_reg[807]  ( .D(c[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[803])
         );
  DFF \sreg_reg[806]  ( .D(c[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[802])
         );
  DFF \sreg_reg[805]  ( .D(c[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[801])
         );
  DFF \sreg_reg[804]  ( .D(c[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[800])
         );
  DFF \sreg_reg[803]  ( .D(c[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[799])
         );
  DFF \sreg_reg[802]  ( .D(c[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[798])
         );
  DFF \sreg_reg[801]  ( .D(c[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[797])
         );
  DFF \sreg_reg[800]  ( .D(c[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[796])
         );
  DFF \sreg_reg[799]  ( .D(c[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[795])
         );
  DFF \sreg_reg[798]  ( .D(c[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[794])
         );
  DFF \sreg_reg[797]  ( .D(c[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[793])
         );
  DFF \sreg_reg[796]  ( .D(c[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[792])
         );
  DFF \sreg_reg[795]  ( .D(c[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[791])
         );
  DFF \sreg_reg[794]  ( .D(c[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[790])
         );
  DFF \sreg_reg[793]  ( .D(c[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[789])
         );
  DFF \sreg_reg[792]  ( .D(c[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[788])
         );
  DFF \sreg_reg[791]  ( .D(c[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[787])
         );
  DFF \sreg_reg[790]  ( .D(c[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[786])
         );
  DFF \sreg_reg[789]  ( .D(c[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[785])
         );
  DFF \sreg_reg[788]  ( .D(c[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[784])
         );
  DFF \sreg_reg[787]  ( .D(c[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[783])
         );
  DFF \sreg_reg[786]  ( .D(c[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[782])
         );
  DFF \sreg_reg[785]  ( .D(c[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[781])
         );
  DFF \sreg_reg[784]  ( .D(c[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[780])
         );
  DFF \sreg_reg[783]  ( .D(c[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[779])
         );
  DFF \sreg_reg[782]  ( .D(c[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[778])
         );
  DFF \sreg_reg[781]  ( .D(c[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[777])
         );
  DFF \sreg_reg[780]  ( .D(c[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[776])
         );
  DFF \sreg_reg[779]  ( .D(c[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[775])
         );
  DFF \sreg_reg[778]  ( .D(c[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[774])
         );
  DFF \sreg_reg[777]  ( .D(c[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[773])
         );
  DFF \sreg_reg[776]  ( .D(c[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[772])
         );
  DFF \sreg_reg[775]  ( .D(c[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[771])
         );
  DFF \sreg_reg[774]  ( .D(c[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[770])
         );
  DFF \sreg_reg[773]  ( .D(c[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[769])
         );
  DFF \sreg_reg[772]  ( .D(c[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[768])
         );
  DFF \sreg_reg[771]  ( .D(c[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[767])
         );
  DFF \sreg_reg[770]  ( .D(c[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[766])
         );
  DFF \sreg_reg[769]  ( .D(c[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[765])
         );
  DFF \sreg_reg[768]  ( .D(c[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[764])
         );
  DFF \sreg_reg[767]  ( .D(c[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[763])
         );
  DFF \sreg_reg[766]  ( .D(c[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[762])
         );
  DFF \sreg_reg[765]  ( .D(c[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[761])
         );
  DFF \sreg_reg[764]  ( .D(c[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[760])
         );
  DFF \sreg_reg[763]  ( .D(c[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[759])
         );
  DFF \sreg_reg[762]  ( .D(c[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[758])
         );
  DFF \sreg_reg[761]  ( .D(c[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[757])
         );
  DFF \sreg_reg[760]  ( .D(c[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[756])
         );
  DFF \sreg_reg[759]  ( .D(c[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[755])
         );
  DFF \sreg_reg[758]  ( .D(c[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[754])
         );
  DFF \sreg_reg[757]  ( .D(c[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[753])
         );
  DFF \sreg_reg[756]  ( .D(c[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[752])
         );
  DFF \sreg_reg[755]  ( .D(c[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[751])
         );
  DFF \sreg_reg[754]  ( .D(c[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[750])
         );
  DFF \sreg_reg[753]  ( .D(c[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[749])
         );
  DFF \sreg_reg[752]  ( .D(c[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[748])
         );
  DFF \sreg_reg[751]  ( .D(c[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[747])
         );
  DFF \sreg_reg[750]  ( .D(c[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[746])
         );
  DFF \sreg_reg[749]  ( .D(c[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[745])
         );
  DFF \sreg_reg[748]  ( .D(c[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[744])
         );
  DFF \sreg_reg[747]  ( .D(c[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[743])
         );
  DFF \sreg_reg[746]  ( .D(c[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[742])
         );
  DFF \sreg_reg[745]  ( .D(c[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[741])
         );
  DFF \sreg_reg[744]  ( .D(c[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[740])
         );
  DFF \sreg_reg[743]  ( .D(c[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[739])
         );
  DFF \sreg_reg[742]  ( .D(c[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[738])
         );
  DFF \sreg_reg[741]  ( .D(c[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[737])
         );
  DFF \sreg_reg[740]  ( .D(c[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[736])
         );
  DFF \sreg_reg[739]  ( .D(c[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[735])
         );
  DFF \sreg_reg[738]  ( .D(c[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[734])
         );
  DFF \sreg_reg[737]  ( .D(c[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[733])
         );
  DFF \sreg_reg[736]  ( .D(c[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[732])
         );
  DFF \sreg_reg[735]  ( .D(c[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[731])
         );
  DFF \sreg_reg[734]  ( .D(c[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[730])
         );
  DFF \sreg_reg[733]  ( .D(c[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[729])
         );
  DFF \sreg_reg[732]  ( .D(c[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[728])
         );
  DFF \sreg_reg[731]  ( .D(c[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[727])
         );
  DFF \sreg_reg[730]  ( .D(c[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[726])
         );
  DFF \sreg_reg[729]  ( .D(c[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[725])
         );
  DFF \sreg_reg[728]  ( .D(c[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[724])
         );
  DFF \sreg_reg[727]  ( .D(c[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[723])
         );
  DFF \sreg_reg[726]  ( .D(c[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[722])
         );
  DFF \sreg_reg[725]  ( .D(c[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[721])
         );
  DFF \sreg_reg[724]  ( .D(c[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[720])
         );
  DFF \sreg_reg[723]  ( .D(c[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[719])
         );
  DFF \sreg_reg[722]  ( .D(c[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[718])
         );
  DFF \sreg_reg[721]  ( .D(c[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[717])
         );
  DFF \sreg_reg[720]  ( .D(c[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[716])
         );
  DFF \sreg_reg[719]  ( .D(c[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[715])
         );
  DFF \sreg_reg[718]  ( .D(c[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[714])
         );
  DFF \sreg_reg[717]  ( .D(c[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[713])
         );
  DFF \sreg_reg[716]  ( .D(c[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[712])
         );
  DFF \sreg_reg[715]  ( .D(c[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[711])
         );
  DFF \sreg_reg[714]  ( .D(c[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[710])
         );
  DFF \sreg_reg[713]  ( .D(c[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[709])
         );
  DFF \sreg_reg[712]  ( .D(c[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[708])
         );
  DFF \sreg_reg[711]  ( .D(c[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[707])
         );
  DFF \sreg_reg[710]  ( .D(c[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[706])
         );
  DFF \sreg_reg[709]  ( .D(c[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[705])
         );
  DFF \sreg_reg[708]  ( .D(c[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[704])
         );
  DFF \sreg_reg[707]  ( .D(c[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[703])
         );
  DFF \sreg_reg[706]  ( .D(c[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[702])
         );
  DFF \sreg_reg[705]  ( .D(c[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[701])
         );
  DFF \sreg_reg[704]  ( .D(c[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[700])
         );
  DFF \sreg_reg[703]  ( .D(c[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[699])
         );
  DFF \sreg_reg[702]  ( .D(c[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[698])
         );
  DFF \sreg_reg[701]  ( .D(c[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[697])
         );
  DFF \sreg_reg[700]  ( .D(c[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[696])
         );
  DFF \sreg_reg[699]  ( .D(c[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[695])
         );
  DFF \sreg_reg[698]  ( .D(c[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[694])
         );
  DFF \sreg_reg[697]  ( .D(c[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[693])
         );
  DFF \sreg_reg[696]  ( .D(c[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[692])
         );
  DFF \sreg_reg[695]  ( .D(c[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[691])
         );
  DFF \sreg_reg[694]  ( .D(c[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[690])
         );
  DFF \sreg_reg[693]  ( .D(c[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[689])
         );
  DFF \sreg_reg[692]  ( .D(c[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[688])
         );
  DFF \sreg_reg[691]  ( .D(c[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[687])
         );
  DFF \sreg_reg[690]  ( .D(c[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[686])
         );
  DFF \sreg_reg[689]  ( .D(c[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[685])
         );
  DFF \sreg_reg[688]  ( .D(c[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[684])
         );
  DFF \sreg_reg[687]  ( .D(c[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[683])
         );
  DFF \sreg_reg[686]  ( .D(c[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[682])
         );
  DFF \sreg_reg[685]  ( .D(c[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[681])
         );
  DFF \sreg_reg[684]  ( .D(c[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[680])
         );
  DFF \sreg_reg[683]  ( .D(c[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[679])
         );
  DFF \sreg_reg[682]  ( .D(c[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[678])
         );
  DFF \sreg_reg[681]  ( .D(c[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[677])
         );
  DFF \sreg_reg[680]  ( .D(c[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[676])
         );
  DFF \sreg_reg[679]  ( .D(c[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[675])
         );
  DFF \sreg_reg[678]  ( .D(c[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[674])
         );
  DFF \sreg_reg[677]  ( .D(c[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[673])
         );
  DFF \sreg_reg[676]  ( .D(c[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[672])
         );
  DFF \sreg_reg[675]  ( .D(c[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[671])
         );
  DFF \sreg_reg[674]  ( .D(c[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[670])
         );
  DFF \sreg_reg[673]  ( .D(c[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[669])
         );
  DFF \sreg_reg[672]  ( .D(c[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[668])
         );
  DFF \sreg_reg[671]  ( .D(c[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[667])
         );
  DFF \sreg_reg[670]  ( .D(c[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[666])
         );
  DFF \sreg_reg[669]  ( .D(c[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[665])
         );
  DFF \sreg_reg[668]  ( .D(c[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[664])
         );
  DFF \sreg_reg[667]  ( .D(c[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[663])
         );
  DFF \sreg_reg[666]  ( .D(c[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[662])
         );
  DFF \sreg_reg[665]  ( .D(c[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[661])
         );
  DFF \sreg_reg[664]  ( .D(c[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[660])
         );
  DFF \sreg_reg[663]  ( .D(c[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[659])
         );
  DFF \sreg_reg[662]  ( .D(c[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[658])
         );
  DFF \sreg_reg[661]  ( .D(c[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[657])
         );
  DFF \sreg_reg[660]  ( .D(c[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[656])
         );
  DFF \sreg_reg[659]  ( .D(c[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[655])
         );
  DFF \sreg_reg[658]  ( .D(c[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[654])
         );
  DFF \sreg_reg[657]  ( .D(c[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[653])
         );
  DFF \sreg_reg[656]  ( .D(c[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[652])
         );
  DFF \sreg_reg[655]  ( .D(c[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[651])
         );
  DFF \sreg_reg[654]  ( .D(c[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[650])
         );
  DFF \sreg_reg[653]  ( .D(c[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[649])
         );
  DFF \sreg_reg[652]  ( .D(c[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[648])
         );
  DFF \sreg_reg[651]  ( .D(c[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[647])
         );
  DFF \sreg_reg[650]  ( .D(c[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[646])
         );
  DFF \sreg_reg[649]  ( .D(c[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[645])
         );
  DFF \sreg_reg[648]  ( .D(c[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[644])
         );
  DFF \sreg_reg[647]  ( .D(c[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[643])
         );
  DFF \sreg_reg[646]  ( .D(c[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[642])
         );
  DFF \sreg_reg[645]  ( .D(c[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[641])
         );
  DFF \sreg_reg[644]  ( .D(c[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[640])
         );
  DFF \sreg_reg[643]  ( .D(c[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[639])
         );
  DFF \sreg_reg[642]  ( .D(c[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[638])
         );
  DFF \sreg_reg[641]  ( .D(c[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[637])
         );
  DFF \sreg_reg[640]  ( .D(c[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[636])
         );
  DFF \sreg_reg[639]  ( .D(c[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[635])
         );
  DFF \sreg_reg[638]  ( .D(c[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[634])
         );
  DFF \sreg_reg[637]  ( .D(c[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[633])
         );
  DFF \sreg_reg[636]  ( .D(c[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[632])
         );
  DFF \sreg_reg[635]  ( .D(c[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[631])
         );
  DFF \sreg_reg[634]  ( .D(c[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[630])
         );
  DFF \sreg_reg[633]  ( .D(c[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[629])
         );
  DFF \sreg_reg[632]  ( .D(c[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[628])
         );
  DFF \sreg_reg[631]  ( .D(c[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[627])
         );
  DFF \sreg_reg[630]  ( .D(c[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[626])
         );
  DFF \sreg_reg[629]  ( .D(c[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[625])
         );
  DFF \sreg_reg[628]  ( .D(c[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[624])
         );
  DFF \sreg_reg[627]  ( .D(c[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[623])
         );
  DFF \sreg_reg[626]  ( .D(c[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[622])
         );
  DFF \sreg_reg[625]  ( .D(c[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[621])
         );
  DFF \sreg_reg[624]  ( .D(c[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[620])
         );
  DFF \sreg_reg[623]  ( .D(c[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[619])
         );
  DFF \sreg_reg[622]  ( .D(c[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[618])
         );
  DFF \sreg_reg[621]  ( .D(c[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[617])
         );
  DFF \sreg_reg[620]  ( .D(c[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[616])
         );
  DFF \sreg_reg[619]  ( .D(c[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[615])
         );
  DFF \sreg_reg[618]  ( .D(c[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[614])
         );
  DFF \sreg_reg[617]  ( .D(c[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[613])
         );
  DFF \sreg_reg[616]  ( .D(c[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[612])
         );
  DFF \sreg_reg[615]  ( .D(c[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[611])
         );
  DFF \sreg_reg[614]  ( .D(c[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[610])
         );
  DFF \sreg_reg[613]  ( .D(c[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[609])
         );
  DFF \sreg_reg[612]  ( .D(c[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[608])
         );
  DFF \sreg_reg[611]  ( .D(c[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[607])
         );
  DFF \sreg_reg[610]  ( .D(c[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[606])
         );
  DFF \sreg_reg[609]  ( .D(c[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[605])
         );
  DFF \sreg_reg[608]  ( .D(c[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[604])
         );
  DFF \sreg_reg[607]  ( .D(c[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[603])
         );
  DFF \sreg_reg[606]  ( .D(c[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[602])
         );
  DFF \sreg_reg[605]  ( .D(c[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[601])
         );
  DFF \sreg_reg[604]  ( .D(c[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[600])
         );
  DFF \sreg_reg[603]  ( .D(c[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[599])
         );
  DFF \sreg_reg[602]  ( .D(c[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[598])
         );
  DFF \sreg_reg[601]  ( .D(c[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[597])
         );
  DFF \sreg_reg[600]  ( .D(c[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[596])
         );
  DFF \sreg_reg[599]  ( .D(c[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[595])
         );
  DFF \sreg_reg[598]  ( .D(c[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[594])
         );
  DFF \sreg_reg[597]  ( .D(c[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[593])
         );
  DFF \sreg_reg[596]  ( .D(c[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[592])
         );
  DFF \sreg_reg[595]  ( .D(c[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[591])
         );
  DFF \sreg_reg[594]  ( .D(c[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[590])
         );
  DFF \sreg_reg[593]  ( .D(c[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[589])
         );
  DFF \sreg_reg[592]  ( .D(c[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[588])
         );
  DFF \sreg_reg[591]  ( .D(c[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[587])
         );
  DFF \sreg_reg[590]  ( .D(c[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[586])
         );
  DFF \sreg_reg[589]  ( .D(c[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[585])
         );
  DFF \sreg_reg[588]  ( .D(c[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[584])
         );
  DFF \sreg_reg[587]  ( .D(c[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[583])
         );
  DFF \sreg_reg[586]  ( .D(c[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[582])
         );
  DFF \sreg_reg[585]  ( .D(c[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[581])
         );
  DFF \sreg_reg[584]  ( .D(c[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[580])
         );
  DFF \sreg_reg[583]  ( .D(c[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[579])
         );
  DFF \sreg_reg[582]  ( .D(c[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[578])
         );
  DFF \sreg_reg[581]  ( .D(c[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[577])
         );
  DFF \sreg_reg[580]  ( .D(c[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[576])
         );
  DFF \sreg_reg[579]  ( .D(c[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[575])
         );
  DFF \sreg_reg[578]  ( .D(c[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[574])
         );
  DFF \sreg_reg[577]  ( .D(c[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[573])
         );
  DFF \sreg_reg[576]  ( .D(c[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[572])
         );
  DFF \sreg_reg[575]  ( .D(c[575]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[571])
         );
  DFF \sreg_reg[574]  ( .D(c[574]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[570])
         );
  DFF \sreg_reg[573]  ( .D(c[573]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[569])
         );
  DFF \sreg_reg[572]  ( .D(c[572]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[568])
         );
  DFF \sreg_reg[571]  ( .D(c[571]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[567])
         );
  DFF \sreg_reg[570]  ( .D(c[570]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[566])
         );
  DFF \sreg_reg[569]  ( .D(c[569]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[565])
         );
  DFF \sreg_reg[568]  ( .D(c[568]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[564])
         );
  DFF \sreg_reg[567]  ( .D(c[567]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[563])
         );
  DFF \sreg_reg[566]  ( .D(c[566]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[562])
         );
  DFF \sreg_reg[565]  ( .D(c[565]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[561])
         );
  DFF \sreg_reg[564]  ( .D(c[564]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[560])
         );
  DFF \sreg_reg[563]  ( .D(c[563]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[559])
         );
  DFF \sreg_reg[562]  ( .D(c[562]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[558])
         );
  DFF \sreg_reg[561]  ( .D(c[561]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[557])
         );
  DFF \sreg_reg[560]  ( .D(c[560]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[556])
         );
  DFF \sreg_reg[559]  ( .D(c[559]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[555])
         );
  DFF \sreg_reg[558]  ( .D(c[558]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[554])
         );
  DFF \sreg_reg[557]  ( .D(c[557]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[553])
         );
  DFF \sreg_reg[556]  ( .D(c[556]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[552])
         );
  DFF \sreg_reg[555]  ( .D(c[555]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[551])
         );
  DFF \sreg_reg[554]  ( .D(c[554]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[550])
         );
  DFF \sreg_reg[553]  ( .D(c[553]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[549])
         );
  DFF \sreg_reg[552]  ( .D(c[552]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[548])
         );
  DFF \sreg_reg[551]  ( .D(c[551]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[547])
         );
  DFF \sreg_reg[550]  ( .D(c[550]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[546])
         );
  DFF \sreg_reg[549]  ( .D(c[549]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[545])
         );
  DFF \sreg_reg[548]  ( .D(c[548]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[544])
         );
  DFF \sreg_reg[547]  ( .D(c[547]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[543])
         );
  DFF \sreg_reg[546]  ( .D(c[546]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[542])
         );
  DFF \sreg_reg[545]  ( .D(c[545]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[541])
         );
  DFF \sreg_reg[544]  ( .D(c[544]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[540])
         );
  DFF \sreg_reg[543]  ( .D(c[543]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[539])
         );
  DFF \sreg_reg[542]  ( .D(c[542]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[538])
         );
  DFF \sreg_reg[541]  ( .D(c[541]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[537])
         );
  DFF \sreg_reg[540]  ( .D(c[540]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[536])
         );
  DFF \sreg_reg[539]  ( .D(c[539]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[535])
         );
  DFF \sreg_reg[538]  ( .D(c[538]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[534])
         );
  DFF \sreg_reg[537]  ( .D(c[537]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[533])
         );
  DFF \sreg_reg[536]  ( .D(c[536]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[532])
         );
  DFF \sreg_reg[535]  ( .D(c[535]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[531])
         );
  DFF \sreg_reg[534]  ( .D(c[534]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[530])
         );
  DFF \sreg_reg[533]  ( .D(c[533]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[529])
         );
  DFF \sreg_reg[532]  ( .D(c[532]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[528])
         );
  DFF \sreg_reg[531]  ( .D(c[531]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[527])
         );
  DFF \sreg_reg[530]  ( .D(c[530]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[526])
         );
  DFF \sreg_reg[529]  ( .D(c[529]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[525])
         );
  DFF \sreg_reg[528]  ( .D(c[528]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[524])
         );
  DFF \sreg_reg[527]  ( .D(c[527]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[523])
         );
  DFF \sreg_reg[526]  ( .D(c[526]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[522])
         );
  DFF \sreg_reg[525]  ( .D(c[525]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[521])
         );
  DFF \sreg_reg[524]  ( .D(c[524]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[520])
         );
  DFF \sreg_reg[523]  ( .D(c[523]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[519])
         );
  DFF \sreg_reg[522]  ( .D(c[522]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[518])
         );
  DFF \sreg_reg[521]  ( .D(c[521]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[517])
         );
  DFF \sreg_reg[520]  ( .D(c[520]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[516])
         );
  DFF \sreg_reg[519]  ( .D(c[519]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[515])
         );
  DFF \sreg_reg[518]  ( .D(c[518]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[514])
         );
  DFF \sreg_reg[517]  ( .D(c[517]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[513])
         );
  DFF \sreg_reg[516]  ( .D(c[516]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[512])
         );
  DFF \sreg_reg[515]  ( .D(c[515]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[511])
         );
  DFF \sreg_reg[514]  ( .D(c[514]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[510])
         );
  DFF \sreg_reg[513]  ( .D(c[513]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[509])
         );
  DFF \sreg_reg[512]  ( .D(c[512]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[508])
         );
  DFF \sreg_reg[511]  ( .D(c[511]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[507])
         );
  DFF \sreg_reg[510]  ( .D(c[510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[506])
         );
  DFF \sreg_reg[509]  ( .D(c[509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[505])
         );
  DFF \sreg_reg[508]  ( .D(c[508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[504])
         );
  DFF \sreg_reg[507]  ( .D(c[507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[503])
         );
  DFF \sreg_reg[506]  ( .D(c[506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[502])
         );
  DFF \sreg_reg[505]  ( .D(c[505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[501])
         );
  DFF \sreg_reg[504]  ( .D(c[504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[500])
         );
  DFF \sreg_reg[503]  ( .D(c[503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[499])
         );
  DFF \sreg_reg[502]  ( .D(c[502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[498])
         );
  DFF \sreg_reg[501]  ( .D(c[501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[497])
         );
  DFF \sreg_reg[500]  ( .D(c[500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[496])
         );
  DFF \sreg_reg[499]  ( .D(c[499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[495])
         );
  DFF \sreg_reg[498]  ( .D(c[498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[494])
         );
  DFF \sreg_reg[497]  ( .D(c[497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[493])
         );
  DFF \sreg_reg[496]  ( .D(c[496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[492])
         );
  DFF \sreg_reg[495]  ( .D(c[495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[491])
         );
  DFF \sreg_reg[494]  ( .D(c[494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[490])
         );
  DFF \sreg_reg[493]  ( .D(c[493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[489])
         );
  DFF \sreg_reg[492]  ( .D(c[492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[488])
         );
  DFF \sreg_reg[491]  ( .D(c[491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[487])
         );
  DFF \sreg_reg[490]  ( .D(c[490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[486])
         );
  DFF \sreg_reg[489]  ( .D(c[489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[485])
         );
  DFF \sreg_reg[488]  ( .D(c[488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[484])
         );
  DFF \sreg_reg[487]  ( .D(c[487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[483])
         );
  DFF \sreg_reg[486]  ( .D(c[486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[482])
         );
  DFF \sreg_reg[485]  ( .D(c[485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[481])
         );
  DFF \sreg_reg[484]  ( .D(c[484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[480])
         );
  DFF \sreg_reg[483]  ( .D(c[483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[479])
         );
  DFF \sreg_reg[482]  ( .D(c[482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[478])
         );
  DFF \sreg_reg[481]  ( .D(c[481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[477])
         );
  DFF \sreg_reg[480]  ( .D(c[480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[476])
         );
  DFF \sreg_reg[479]  ( .D(c[479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[475])
         );
  DFF \sreg_reg[478]  ( .D(c[478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[474])
         );
  DFF \sreg_reg[477]  ( .D(c[477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[473])
         );
  DFF \sreg_reg[476]  ( .D(c[476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[472])
         );
  DFF \sreg_reg[475]  ( .D(c[475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[471])
         );
  DFF \sreg_reg[474]  ( .D(c[474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[470])
         );
  DFF \sreg_reg[473]  ( .D(c[473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[469])
         );
  DFF \sreg_reg[472]  ( .D(c[472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[468])
         );
  DFF \sreg_reg[471]  ( .D(c[471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[467])
         );
  DFF \sreg_reg[470]  ( .D(c[470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[466])
         );
  DFF \sreg_reg[469]  ( .D(c[469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[465])
         );
  DFF \sreg_reg[468]  ( .D(c[468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[464])
         );
  DFF \sreg_reg[467]  ( .D(c[467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[463])
         );
  DFF \sreg_reg[466]  ( .D(c[466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[462])
         );
  DFF \sreg_reg[465]  ( .D(c[465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[461])
         );
  DFF \sreg_reg[464]  ( .D(c[464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[460])
         );
  DFF \sreg_reg[463]  ( .D(c[463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[459])
         );
  DFF \sreg_reg[462]  ( .D(c[462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[458])
         );
  DFF \sreg_reg[461]  ( .D(c[461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[457])
         );
  DFF \sreg_reg[460]  ( .D(c[460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[456])
         );
  DFF \sreg_reg[459]  ( .D(c[459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[455])
         );
  DFF \sreg_reg[458]  ( .D(c[458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[454])
         );
  DFF \sreg_reg[457]  ( .D(c[457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[453])
         );
  DFF \sreg_reg[456]  ( .D(c[456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[452])
         );
  DFF \sreg_reg[455]  ( .D(c[455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[451])
         );
  DFF \sreg_reg[454]  ( .D(c[454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[450])
         );
  DFF \sreg_reg[453]  ( .D(c[453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[449])
         );
  DFF \sreg_reg[452]  ( .D(c[452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[448])
         );
  DFF \sreg_reg[451]  ( .D(c[451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[447])
         );
  DFF \sreg_reg[450]  ( .D(c[450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[446])
         );
  DFF \sreg_reg[449]  ( .D(c[449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[445])
         );
  DFF \sreg_reg[448]  ( .D(c[448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[444])
         );
  DFF \sreg_reg[447]  ( .D(c[447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[443])
         );
  DFF \sreg_reg[446]  ( .D(c[446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[442])
         );
  DFF \sreg_reg[445]  ( .D(c[445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[441])
         );
  DFF \sreg_reg[444]  ( .D(c[444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[440])
         );
  DFF \sreg_reg[443]  ( .D(c[443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[439])
         );
  DFF \sreg_reg[442]  ( .D(c[442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[438])
         );
  DFF \sreg_reg[441]  ( .D(c[441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[437])
         );
  DFF \sreg_reg[440]  ( .D(c[440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[436])
         );
  DFF \sreg_reg[439]  ( .D(c[439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[435])
         );
  DFF \sreg_reg[438]  ( .D(c[438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[434])
         );
  DFF \sreg_reg[437]  ( .D(c[437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[433])
         );
  DFF \sreg_reg[436]  ( .D(c[436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[432])
         );
  DFF \sreg_reg[435]  ( .D(c[435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[431])
         );
  DFF \sreg_reg[434]  ( .D(c[434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[430])
         );
  DFF \sreg_reg[433]  ( .D(c[433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[429])
         );
  DFF \sreg_reg[432]  ( .D(c[432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[428])
         );
  DFF \sreg_reg[431]  ( .D(c[431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[427])
         );
  DFF \sreg_reg[430]  ( .D(c[430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[426])
         );
  DFF \sreg_reg[429]  ( .D(c[429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[425])
         );
  DFF \sreg_reg[428]  ( .D(c[428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[424])
         );
  DFF \sreg_reg[427]  ( .D(c[427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[423])
         );
  DFF \sreg_reg[426]  ( .D(c[426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[422])
         );
  DFF \sreg_reg[425]  ( .D(c[425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[421])
         );
  DFF \sreg_reg[424]  ( .D(c[424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[420])
         );
  DFF \sreg_reg[423]  ( .D(c[423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[419])
         );
  DFF \sreg_reg[422]  ( .D(c[422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[418])
         );
  DFF \sreg_reg[421]  ( .D(c[421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[417])
         );
  DFF \sreg_reg[420]  ( .D(c[420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[416])
         );
  DFF \sreg_reg[419]  ( .D(c[419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[415])
         );
  DFF \sreg_reg[418]  ( .D(c[418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[414])
         );
  DFF \sreg_reg[417]  ( .D(c[417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[413])
         );
  DFF \sreg_reg[416]  ( .D(c[416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[412])
         );
  DFF \sreg_reg[415]  ( .D(c[415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[411])
         );
  DFF \sreg_reg[414]  ( .D(c[414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[410])
         );
  DFF \sreg_reg[413]  ( .D(c[413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[409])
         );
  DFF \sreg_reg[412]  ( .D(c[412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[408])
         );
  DFF \sreg_reg[411]  ( .D(c[411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[407])
         );
  DFF \sreg_reg[410]  ( .D(c[410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[406])
         );
  DFF \sreg_reg[409]  ( .D(c[409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[405])
         );
  DFF \sreg_reg[408]  ( .D(c[408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[404])
         );
  DFF \sreg_reg[407]  ( .D(c[407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[403])
         );
  DFF \sreg_reg[406]  ( .D(c[406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[402])
         );
  DFF \sreg_reg[405]  ( .D(c[405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[401])
         );
  DFF \sreg_reg[404]  ( .D(c[404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[400])
         );
  DFF \sreg_reg[403]  ( .D(c[403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[399])
         );
  DFF \sreg_reg[402]  ( .D(c[402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[398])
         );
  DFF \sreg_reg[401]  ( .D(c[401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[397])
         );
  DFF \sreg_reg[400]  ( .D(c[400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[396])
         );
  DFF \sreg_reg[399]  ( .D(c[399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[395])
         );
  DFF \sreg_reg[398]  ( .D(c[398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[394])
         );
  DFF \sreg_reg[397]  ( .D(c[397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[393])
         );
  DFF \sreg_reg[396]  ( .D(c[396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[392])
         );
  DFF \sreg_reg[395]  ( .D(c[395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[391])
         );
  DFF \sreg_reg[394]  ( .D(c[394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[390])
         );
  DFF \sreg_reg[393]  ( .D(c[393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[389])
         );
  DFF \sreg_reg[392]  ( .D(c[392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[388])
         );
  DFF \sreg_reg[391]  ( .D(c[391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[387])
         );
  DFF \sreg_reg[390]  ( .D(c[390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[386])
         );
  DFF \sreg_reg[389]  ( .D(c[389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[385])
         );
  DFF \sreg_reg[388]  ( .D(c[388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[384])
         );
  DFF \sreg_reg[387]  ( .D(c[387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[383])
         );
  DFF \sreg_reg[386]  ( .D(c[386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[382])
         );
  DFF \sreg_reg[385]  ( .D(c[385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[381])
         );
  DFF \sreg_reg[384]  ( .D(c[384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[380])
         );
  DFF \sreg_reg[383]  ( .D(c[383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[379])
         );
  DFF \sreg_reg[382]  ( .D(c[382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[378])
         );
  DFF \sreg_reg[381]  ( .D(c[381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[377])
         );
  DFF \sreg_reg[380]  ( .D(c[380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[376])
         );
  DFF \sreg_reg[379]  ( .D(c[379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[375])
         );
  DFF \sreg_reg[378]  ( .D(c[378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[374])
         );
  DFF \sreg_reg[377]  ( .D(c[377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[373])
         );
  DFF \sreg_reg[376]  ( .D(c[376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[372])
         );
  DFF \sreg_reg[375]  ( .D(c[375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[371])
         );
  DFF \sreg_reg[374]  ( .D(c[374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[370])
         );
  DFF \sreg_reg[373]  ( .D(c[373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[369])
         );
  DFF \sreg_reg[372]  ( .D(c[372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[368])
         );
  DFF \sreg_reg[371]  ( .D(c[371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[367])
         );
  DFF \sreg_reg[370]  ( .D(c[370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[366])
         );
  DFF \sreg_reg[369]  ( .D(c[369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[365])
         );
  DFF \sreg_reg[368]  ( .D(c[368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[364])
         );
  DFF \sreg_reg[367]  ( .D(c[367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[363])
         );
  DFF \sreg_reg[366]  ( .D(c[366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[362])
         );
  DFF \sreg_reg[365]  ( .D(c[365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[361])
         );
  DFF \sreg_reg[364]  ( .D(c[364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[360])
         );
  DFF \sreg_reg[363]  ( .D(c[363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[359])
         );
  DFF \sreg_reg[362]  ( .D(c[362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[358])
         );
  DFF \sreg_reg[361]  ( .D(c[361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[357])
         );
  DFF \sreg_reg[360]  ( .D(c[360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[356])
         );
  DFF \sreg_reg[359]  ( .D(c[359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[355])
         );
  DFF \sreg_reg[358]  ( .D(c[358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[354])
         );
  DFF \sreg_reg[357]  ( .D(c[357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[353])
         );
  DFF \sreg_reg[356]  ( .D(c[356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[352])
         );
  DFF \sreg_reg[355]  ( .D(c[355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[351])
         );
  DFF \sreg_reg[354]  ( .D(c[354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[350])
         );
  DFF \sreg_reg[353]  ( .D(c[353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[349])
         );
  DFF \sreg_reg[352]  ( .D(c[352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[348])
         );
  DFF \sreg_reg[351]  ( .D(c[351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[347])
         );
  DFF \sreg_reg[350]  ( .D(c[350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[346])
         );
  DFF \sreg_reg[349]  ( .D(c[349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[345])
         );
  DFF \sreg_reg[348]  ( .D(c[348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[344])
         );
  DFF \sreg_reg[347]  ( .D(c[347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[343])
         );
  DFF \sreg_reg[346]  ( .D(c[346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[342])
         );
  DFF \sreg_reg[345]  ( .D(c[345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[341])
         );
  DFF \sreg_reg[344]  ( .D(c[344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[340])
         );
  DFF \sreg_reg[343]  ( .D(c[343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[339])
         );
  DFF \sreg_reg[342]  ( .D(c[342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[338])
         );
  DFF \sreg_reg[341]  ( .D(c[341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[337])
         );
  DFF \sreg_reg[340]  ( .D(c[340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[336])
         );
  DFF \sreg_reg[339]  ( .D(c[339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[335])
         );
  DFF \sreg_reg[338]  ( .D(c[338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[334])
         );
  DFF \sreg_reg[337]  ( .D(c[337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[333])
         );
  DFF \sreg_reg[336]  ( .D(c[336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[332])
         );
  DFF \sreg_reg[335]  ( .D(c[335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[331])
         );
  DFF \sreg_reg[334]  ( .D(c[334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[330])
         );
  DFF \sreg_reg[333]  ( .D(c[333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[329])
         );
  DFF \sreg_reg[332]  ( .D(c[332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[328])
         );
  DFF \sreg_reg[331]  ( .D(c[331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[327])
         );
  DFF \sreg_reg[330]  ( .D(c[330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[326])
         );
  DFF \sreg_reg[329]  ( .D(c[329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[325])
         );
  DFF \sreg_reg[328]  ( .D(c[328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[324])
         );
  DFF \sreg_reg[327]  ( .D(c[327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[323])
         );
  DFF \sreg_reg[326]  ( .D(c[326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[322])
         );
  DFF \sreg_reg[325]  ( .D(c[325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[321])
         );
  DFF \sreg_reg[324]  ( .D(c[324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[320])
         );
  DFF \sreg_reg[323]  ( .D(c[323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[319])
         );
  DFF \sreg_reg[322]  ( .D(c[322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[318])
         );
  DFF \sreg_reg[321]  ( .D(c[321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[317])
         );
  DFF \sreg_reg[320]  ( .D(c[320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[316])
         );
  DFF \sreg_reg[319]  ( .D(c[319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[315])
         );
  DFF \sreg_reg[318]  ( .D(c[318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[314])
         );
  DFF \sreg_reg[317]  ( .D(c[317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[313])
         );
  DFF \sreg_reg[316]  ( .D(c[316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[312])
         );
  DFF \sreg_reg[315]  ( .D(c[315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[311])
         );
  DFF \sreg_reg[314]  ( .D(c[314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[310])
         );
  DFF \sreg_reg[313]  ( .D(c[313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[309])
         );
  DFF \sreg_reg[312]  ( .D(c[312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[308])
         );
  DFF \sreg_reg[311]  ( .D(c[311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[307])
         );
  DFF \sreg_reg[310]  ( .D(c[310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[306])
         );
  DFF \sreg_reg[309]  ( .D(c[309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[305])
         );
  DFF \sreg_reg[308]  ( .D(c[308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[304])
         );
  DFF \sreg_reg[307]  ( .D(c[307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[303])
         );
  DFF \sreg_reg[306]  ( .D(c[306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[302])
         );
  DFF \sreg_reg[305]  ( .D(c[305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[301])
         );
  DFF \sreg_reg[304]  ( .D(c[304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[300])
         );
  DFF \sreg_reg[303]  ( .D(c[303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[299])
         );
  DFF \sreg_reg[302]  ( .D(c[302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[298])
         );
  DFF \sreg_reg[301]  ( .D(c[301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[297])
         );
  DFF \sreg_reg[300]  ( .D(c[300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[296])
         );
  DFF \sreg_reg[299]  ( .D(c[299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[295])
         );
  DFF \sreg_reg[298]  ( .D(c[298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[294])
         );
  DFF \sreg_reg[297]  ( .D(c[297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[293])
         );
  DFF \sreg_reg[296]  ( .D(c[296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[292])
         );
  DFF \sreg_reg[295]  ( .D(c[295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[291])
         );
  DFF \sreg_reg[294]  ( .D(c[294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[290])
         );
  DFF \sreg_reg[293]  ( .D(c[293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[289])
         );
  DFF \sreg_reg[292]  ( .D(c[292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[288])
         );
  DFF \sreg_reg[291]  ( .D(c[291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[287])
         );
  DFF \sreg_reg[290]  ( .D(c[290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[286])
         );
  DFF \sreg_reg[289]  ( .D(c[289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[285])
         );
  DFF \sreg_reg[288]  ( .D(c[288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[284])
         );
  DFF \sreg_reg[287]  ( .D(c[287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[283])
         );
  DFF \sreg_reg[286]  ( .D(c[286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[282])
         );
  DFF \sreg_reg[285]  ( .D(c[285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[281])
         );
  DFF \sreg_reg[284]  ( .D(c[284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[280])
         );
  DFF \sreg_reg[283]  ( .D(c[283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[279])
         );
  DFF \sreg_reg[282]  ( .D(c[282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[278])
         );
  DFF \sreg_reg[281]  ( .D(c[281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[277])
         );
  DFF \sreg_reg[280]  ( .D(c[280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[276])
         );
  DFF \sreg_reg[279]  ( .D(c[279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[275])
         );
  DFF \sreg_reg[278]  ( .D(c[278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[274])
         );
  DFF \sreg_reg[277]  ( .D(c[277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[273])
         );
  DFF \sreg_reg[276]  ( .D(c[276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[272])
         );
  DFF \sreg_reg[275]  ( .D(c[275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[271])
         );
  DFF \sreg_reg[274]  ( .D(c[274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[270])
         );
  DFF \sreg_reg[273]  ( .D(c[273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[269])
         );
  DFF \sreg_reg[272]  ( .D(c[272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[268])
         );
  DFF \sreg_reg[271]  ( .D(c[271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[267])
         );
  DFF \sreg_reg[270]  ( .D(c[270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[266])
         );
  DFF \sreg_reg[269]  ( .D(c[269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[265])
         );
  DFF \sreg_reg[268]  ( .D(c[268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[264])
         );
  DFF \sreg_reg[267]  ( .D(c[267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[263])
         );
  DFF \sreg_reg[266]  ( .D(c[266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[262])
         );
  DFF \sreg_reg[265]  ( .D(c[265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[261])
         );
  DFF \sreg_reg[264]  ( .D(c[264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[260])
         );
  DFF \sreg_reg[263]  ( .D(c[263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[259])
         );
  DFF \sreg_reg[262]  ( .D(c[262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[258])
         );
  DFF \sreg_reg[261]  ( .D(c[261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[257])
         );
  DFF \sreg_reg[260]  ( .D(c[260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[256])
         );
  DFF \sreg_reg[259]  ( .D(c[259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[255])
         );
  DFF \sreg_reg[258]  ( .D(c[258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[254])
         );
  DFF \sreg_reg[257]  ( .D(c[257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[253])
         );
  DFF \sreg_reg[256]  ( .D(c[256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[252])
         );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[251])
         );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[250])
         );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[249])
         );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[248])
         );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[247])
         );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[246])
         );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[245])
         );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[244])
         );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[243])
         );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[242])
         );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[241])
         );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[240])
         );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[239])
         );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[238])
         );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[237])
         );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[236])
         );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[235])
         );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[234])
         );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[233])
         );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[232])
         );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[231])
         );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[230])
         );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[229])
         );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[228])
         );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[227])
         );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[226])
         );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[225])
         );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[224])
         );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[223])
         );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[222])
         );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[221])
         );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[220])
         );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[219])
         );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[218])
         );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[217])
         );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[216])
         );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[215])
         );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[214])
         );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[213])
         );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[212])
         );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[211])
         );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[210])
         );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[209])
         );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[208])
         );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[207])
         );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[206])
         );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[205])
         );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[204])
         );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[203])
         );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[202])
         );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[201])
         );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[200])
         );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[199])
         );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[198])
         );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[197])
         );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[196])
         );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[195])
         );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[194])
         );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[193])
         );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[192])
         );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[191])
         );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[190])
         );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[189])
         );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[188])
         );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[187])
         );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[186])
         );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[185])
         );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[184])
         );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[183])
         );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[182])
         );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[181])
         );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[180])
         );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[179])
         );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[178])
         );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[177])
         );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[176])
         );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[175])
         );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[174])
         );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[173])
         );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[172])
         );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[171])
         );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[170])
         );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[169])
         );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[168])
         );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[167])
         );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[166])
         );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[165])
         );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[164])
         );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[163])
         );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[162])
         );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[161])
         );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[160])
         );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[159])
         );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[158])
         );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[157])
         );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[156])
         );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[155])
         );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[154])
         );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[153])
         );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[152])
         );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[151])
         );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[150])
         );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[149])
         );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[148])
         );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[147])
         );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[146])
         );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[145])
         );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[144])
         );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[143])
         );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[142])
         );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[141])
         );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[140])
         );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[139])
         );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[138])
         );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[137])
         );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[136])
         );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[135])
         );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[134])
         );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[133])
         );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[132])
         );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[131])
         );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[130])
         );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[129])
         );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[128])
         );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[127])
         );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[126])
         );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[125])
         );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[124])
         );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[123])
         );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[122])
         );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[121])
         );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[120])
         );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[119])
         );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[118])
         );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[117])
         );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[116])
         );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[115])
         );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[114])
         );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[113])
         );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[112])
         );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[111])
         );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[110])
         );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[109])
         );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[108])
         );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[107])
         );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[106])
         );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[105])
         );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[104])
         );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[103])
         );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[102])
         );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[101])
         );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[100])
         );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[99])
         );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[98])
         );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[97])
         );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[96])
         );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[95]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[94]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[93]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[92]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[91]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[90]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[89]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[88]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[87]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[86]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[85]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[84]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[83]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[82]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[81]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[80]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[79]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[78]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[77]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[76]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[75]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[74]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[73]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[72]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[71]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[70]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[69]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[68]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[67]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[66]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[65]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[64]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[63]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[62]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[61]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[60]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(c[0]) );
  ADD_N1024 ADD_ ( .A({1'b0, 1'b0, 1'b0, 1'b0, sreg[2043:1024]}), .B(clocal), 
        .CI(1'b0), .S({swire, c[1023:1020]}) );
  mult_N1024_CC256_DW02_mult_0 mult_44 ( .A(a), .B(b), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, clocal}) );
endmodule

