
module round_2 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XOR U1 ( .A(n1390), .B(n1431), .Z(n4463) );
  AND U2 ( .A(n4755), .B(n4362), .Z(n1) );
  XNOR U3 ( .A(n4583), .B(n1), .Z(out[713]) );
  ANDN U4 ( .B(n5051), .A(n1646), .Z(n2) );
  XNOR U5 ( .A(n1841), .B(n2), .Z(out[1100]) );
  XNOR U6 ( .A(n1455), .B(n1036), .Z(n2780) );
  XNOR U7 ( .A(n1461), .B(n1062), .Z(n2817) );
  XOR U8 ( .A(n1448), .B(n766), .Z(n4491) );
  XNOR U9 ( .A(n1701), .B(n1702), .Z(n3083) );
  XOR U10 ( .A(n781), .B(n1450), .Z(n4494) );
  XOR U11 ( .A(n796), .B(n1452), .Z(n4497) );
  XNOR U12 ( .A(n1714), .B(n1715), .Z(n3088) );
  XOR U13 ( .A(n822), .B(n1454), .Z(n4500) );
  XOR U14 ( .A(n1456), .B(n837), .Z(n4503) );
  XOR U15 ( .A(n1460), .B(n852), .Z(n4506) );
  AND U16 ( .A(n2599), .B(n2399), .Z(n3) );
  XNOR U17 ( .A(n2600), .B(n3), .Z(out[1513]) );
  AND U18 ( .A(n4759), .B(n4365), .Z(n4) );
  XNOR U19 ( .A(n4585), .B(n4), .Z(out[714]) );
  NANDN U20 ( .A(n4464), .B(n4883), .Z(n5) );
  XNOR U21 ( .A(n4663), .B(n5), .Z(out[742]) );
  ANDN U22 ( .B(n3505), .A(n3692), .Z(n6) );
  XNOR U23 ( .A(n3693), .B(n6), .Z(out[530]) );
  ANDN U24 ( .B(n3500), .A(n3688), .Z(n7) );
  XNOR U25 ( .A(n3689), .B(n7), .Z(out[529]) );
  ANDN U26 ( .B(n3507), .A(n3700), .Z(n8) );
  XNOR U27 ( .A(n3701), .B(n8), .Z(out[532]) );
  ANDN U28 ( .B(n3512), .A(n3726), .Z(n9) );
  XNOR U29 ( .A(n3727), .B(n9), .Z(out[537]) );
  NAND U30 ( .A(n3837), .B(n3417), .Z(n10) );
  XNOR U31 ( .A(n3416), .B(n10), .Z(out[434]) );
  NAND U32 ( .A(n3841), .B(n3420), .Z(n11) );
  XNOR U33 ( .A(n3419), .B(n11), .Z(out[435]) );
  ANDN U34 ( .B(n3845), .A(n3428), .Z(n12) );
  XNOR U35 ( .A(n3586), .B(n12), .Z(out[436]) );
  NANDN U36 ( .A(n3449), .B(n3877), .Z(n13) );
  XNOR U37 ( .A(n3603), .B(n13), .Z(out[443]) );
  AND U38 ( .A(n3889), .B(n3462), .Z(n14) );
  XNOR U39 ( .A(n3608), .B(n14), .Z(out[446]) );
  ANDN U40 ( .B(n3615), .A(n3261), .Z(n15) );
  XNOR U41 ( .A(n3467), .B(n15), .Z(out[384]) );
  NANDN U42 ( .A(n3277), .B(n3635), .Z(n16) );
  XNOR U43 ( .A(n3475), .B(n16), .Z(out[388]) );
  NANDN U44 ( .A(n3280), .B(n3639), .Z(n17) );
  XNOR U45 ( .A(n3476), .B(n17), .Z(out[389]) );
  NANDN U46 ( .A(n3283), .B(n3643), .Z(n18) );
  XNOR U47 ( .A(n3477), .B(n18), .Z(out[390]) );
  NANDN U48 ( .A(n3286), .B(n3647), .Z(n19) );
  XNOR U49 ( .A(n3478), .B(n19), .Z(out[391]) );
  NANDN U50 ( .A(n3289), .B(n3651), .Z(n20) );
  XNOR U51 ( .A(n3483), .B(n20), .Z(out[392]) );
  ANDN U52 ( .B(n2435), .A(n2434), .Z(n21) );
  XNOR U53 ( .A(n2436), .B(round_const[0]), .Z(n22) );
  XOR U54 ( .A(n21), .B(n22), .Z(out[1536]) );
  ANDN U55 ( .B(n2478), .A(n2477), .Z(n23) );
  XNOR U56 ( .A(n2476), .B(n23), .Z(out[1547]) );
  XNOR U57 ( .A(n1449), .B(n1756), .Z(n3217) );
  XNOR U58 ( .A(n1459), .B(n1049), .Z(n2794) );
  XNOR U59 ( .A(n1463), .B(n1075), .Z(n2840) );
  XNOR U60 ( .A(n1685), .B(n1686), .Z(n3073) );
  XOR U61 ( .A(n1437), .B(n1402), .Z(n4472) );
  XNOR U62 ( .A(n1473), .B(n1103), .Z(n2888) );
  XOR U63 ( .A(n1439), .B(n1406), .Z(n4479) );
  XNOR U64 ( .A(n1477), .B(n1123), .Z(n2921) );
  XOR U65 ( .A(n736), .B(n1442), .Z(n4485) );
  XNOR U66 ( .A(n1718), .B(n1719), .Z(n3090) );
  XNOR U67 ( .A(n1710), .B(n1352), .Z(n3931) );
  XNOR U68 ( .A(n1436), .B(n1731), .Z(n3199) );
  XNOR U69 ( .A(n1751), .B(n1752), .Z(n3104) );
  XNOR U70 ( .A(n1451), .B(n1010), .Z(n2756) );
  XOR U71 ( .A(n1398), .B(n1435), .Z(n4469) );
  XOR U72 ( .A(n1394), .B(n1433), .Z(n4466) );
  XOR U73 ( .A(n1386), .B(n1429), .Z(n4460) );
  XNOR U74 ( .A(n3962), .B(in[1486]), .Z(n4783) );
  XNOR U75 ( .A(n3946), .B(in[1482]), .Z(n4763) );
  AND U76 ( .A(n4739), .B(n4351), .Z(n24) );
  XNOR U77 ( .A(n4570), .B(n24), .Z(out[709]) );
  NANDN U78 ( .A(n4458), .B(n4875), .Z(n25) );
  XNOR U79 ( .A(n4655), .B(n25), .Z(out[740]) );
  ANDN U80 ( .B(n3506), .A(n3696), .Z(n26) );
  XNOR U81 ( .A(n3697), .B(n26), .Z(out[531]) );
  ANDN U82 ( .B(n3509), .A(n3708), .Z(n27) );
  XNOR U83 ( .A(n3709), .B(n27), .Z(out[534]) );
  NANDN U84 ( .A(n3446), .B(n3873), .Z(n28) );
  XNOR U85 ( .A(n3602), .B(n28), .Z(out[442]) );
  ANDN U86 ( .B(n3881), .A(n3452), .Z(n29) );
  XNOR U87 ( .A(n3604), .B(n29), .Z(out[444]) );
  ANDN U88 ( .B(n3885), .A(n3455), .Z(n30) );
  XNOR U89 ( .A(n3606), .B(n30), .Z(out[445]) );
  ANDN U90 ( .B(n3893), .A(n3465), .Z(n31) );
  XNOR U91 ( .A(n3610), .B(n31), .Z(out[447]) );
  ANDN U92 ( .B(n1948), .A(n1541), .Z(n32) );
  XNOR U93 ( .A(n1780), .B(n32), .Z(out[1074]) );
  ANDN U94 ( .B(n1952), .A(n1545), .Z(n33) );
  XNOR U95 ( .A(n1782), .B(n33), .Z(out[1075]) );
  NAND U96 ( .A(n3483), .B(n3649), .Z(n34) );
  XNOR U97 ( .A(n3648), .B(n34), .Z(out[520]) );
  ANDN U98 ( .B(n1960), .A(n1555), .Z(n35) );
  XNOR U99 ( .A(n1786), .B(n35), .Z(out[1077]) );
  NAND U100 ( .A(n4642), .B(n4849), .Z(n36) );
  XNOR U101 ( .A(n4848), .B(n36), .Z(out[863]) );
  NAND U102 ( .A(n2895), .B(n4440), .Z(n37) );
  XNOR U103 ( .A(n2894), .B(n37), .Z(out[207]) );
  NAND U104 ( .A(n2901), .B(n4512), .Z(n38) );
  XNOR U105 ( .A(n2900), .B(n38), .Z(out[209]) );
  ANDN U106 ( .B(n2952), .A(n5158), .Z(n39) );
  XNOR U107 ( .A(n3096), .B(n39), .Z(out[227]) );
  AND U108 ( .A(n4631), .B(n4630), .Z(n40) );
  XNOR U109 ( .A(n4632), .B(n40), .Z(out[85]) );
  ANDN U110 ( .B(n5055), .A(n1650), .Z(n41) );
  XNOR U111 ( .A(n1843), .B(n41), .Z(out[1101]) );
  AND U112 ( .A(n5066), .B(n1662), .Z(n42) );
  XNOR U113 ( .A(n1851), .B(n42), .Z(out[1104]) );
  NANDN U114 ( .A(n4881), .B(n4663), .Z(n43) );
  XNOR U115 ( .A(n4880), .B(n43), .Z(out[870]) );
  AND U116 ( .A(n4743), .B(n4354), .Z(n44) );
  XNOR U117 ( .A(n4572), .B(n44), .Z(out[710]) );
  ANDN U118 ( .B(n4671), .A(n4912), .Z(n45) );
  XNOR U119 ( .A(n4913), .B(n45), .Z(out[877]) );
  ANDN U120 ( .B(n4672), .A(n4916), .Z(n46) );
  XNOR U121 ( .A(n4917), .B(n46), .Z(out[878]) );
  NAND U122 ( .A(n2856), .B(n2855), .Z(n47) );
  XNOR U123 ( .A(n3939), .B(n47), .Z(out[256]) );
  NANDN U124 ( .A(n3641), .B(n3477), .Z(n48) );
  XNOR U125 ( .A(n3640), .B(n48), .Z(out[518]) );
  XNOR U126 ( .A(n1660), .B(n1661), .Z(n3059) );
  XNOR U127 ( .A(n1407), .B(n1682), .Z(n3171) );
  XNOR U128 ( .A(n1689), .B(n1690), .Z(n3077) );
  XNOR U129 ( .A(n1705), .B(n1706), .Z(n3085) );
  XOR U130 ( .A(n1440), .B(n721), .Z(n4482) );
  XNOR U131 ( .A(n1486), .B(n1162), .Z(n4062) );
  XNOR U132 ( .A(n1411), .B(n1686), .Z(n3173) );
  XNOR U133 ( .A(n1462), .B(n867), .Z(n4513) );
  XNOR U134 ( .A(n1464), .B(n882), .Z(n4516) );
  XNOR U135 ( .A(n1438), .B(n1735), .Z(n3202) );
  XOR U136 ( .A(n1484), .B(n687), .Z(n4534) );
  XOR U137 ( .A(n1482), .B(n942), .Z(n4530) );
  XNOR U138 ( .A(n1426), .B(n1711), .Z(n3185) );
  XNOR U139 ( .A(n1445), .B(n1747), .Z(n3211) );
  XNOR U140 ( .A(n1428), .B(n1715), .Z(n3187) );
  XNOR U141 ( .A(n1447), .B(n1752), .Z(n3214) );
  XNOR U142 ( .A(n1430), .B(n1719), .Z(n2294) );
  XNOR U143 ( .A(n1417), .B(n1698), .Z(n3179) );
  XOR U144 ( .A(n1474), .B(n912), .Z(n4522) );
  XNOR U145 ( .A(n1419), .B(n1702), .Z(n3181) );
  XNOR U146 ( .A(n1432), .B(n1723), .Z(n3194) );
  XNOR U147 ( .A(n1755), .B(n1756), .Z(n3106) );
  XOR U148 ( .A(n1489), .B(n815), .Z(n4542) );
  XNOR U149 ( .A(n1434), .B(n1727), .Z(n3196) );
  XNOR U150 ( .A(n3950), .B(in[1483]), .Z(n4767) );
  XNOR U151 ( .A(n3954), .B(in[1484]), .Z(n4771) );
  XNOR U152 ( .A(n3970), .B(in[1488]), .Z(n4791) );
  AND U153 ( .A(n3422), .B(n2984), .Z(n49) );
  XNOR U154 ( .A(n3423), .B(n49), .Z(out[305]) );
  AND U155 ( .A(n4751), .B(n4359), .Z(n50) );
  XNOR U156 ( .A(n4581), .B(n50), .Z(out[712]) );
  ANDN U157 ( .B(n3510), .A(n3712), .Z(n51) );
  XNOR U158 ( .A(n3713), .B(n51), .Z(out[535]) );
  ANDN U159 ( .B(n1998), .A(n1591), .Z(n52) );
  XNOR U160 ( .A(n1806), .B(n52), .Z(out[1086]) );
  ANDN U161 ( .B(n3861), .A(n3437), .Z(n53) );
  XNOR U162 ( .A(n3592), .B(n53), .Z(out[439]) );
  ANDN U163 ( .B(n3869), .A(n3443), .Z(n54) );
  XNOR U164 ( .A(n3596), .B(n54), .Z(out[441]) );
  ANDN U165 ( .B(n1940), .A(n1533), .Z(n55) );
  XNOR U166 ( .A(n1776), .B(n55), .Z(out[1072]) );
  ANDN U167 ( .B(n1966), .A(n1559), .Z(n56) );
  XNOR U168 ( .A(n1788), .B(n56), .Z(out[1078]) );
  NAND U169 ( .A(n2892), .B(n4406), .Z(n57) );
  XNOR U170 ( .A(n2891), .B(n57), .Z(out[206]) );
  NANDN U171 ( .A(n2934), .B(n4819), .Z(n58) );
  XNOR U172 ( .A(n2933), .B(n58), .Z(out[219]) );
  ANDN U173 ( .B(n2454), .A(n2453), .Z(n59) );
  XNOR U174 ( .A(n2452), .B(n59), .Z(out[1540]) );
  ANDN U175 ( .B(n2457), .A(n2456), .Z(n60) );
  XNOR U176 ( .A(n2455), .B(n60), .Z(out[1541]) );
  AND U177 ( .A(n4675), .B(n4674), .Z(n61) );
  XNOR U178 ( .A(n4676), .B(n61), .Z(out[87]) );
  AND U179 ( .A(n4691), .B(n4690), .Z(n62) );
  XNOR U180 ( .A(n4692), .B(n62), .Z(out[88]) );
  AND U181 ( .A(n5072), .B(n1671), .Z(n63) );
  XNOR U182 ( .A(n1855), .B(n63), .Z(out[1106]) );
  NANDN U183 ( .A(n4877), .B(n4658), .Z(n64) );
  XNOR U184 ( .A(n4876), .B(n64), .Z(out[869]) );
  ANDN U185 ( .B(n2469), .A(n2468), .Z(n65) );
  XNOR U186 ( .A(n2467), .B(n65), .Z(out[1544]) );
  ANDN U187 ( .B(n5083), .A(n1679), .Z(n66) );
  XNOR U188 ( .A(n1859), .B(n66), .Z(out[1108]) );
  ANDN U189 ( .B(n2472), .A(n2471), .Z(n67) );
  XNOR U190 ( .A(n2470), .B(n67), .Z(out[1545]) );
  ANDN U191 ( .B(n2475), .A(n2474), .Z(n68) );
  XNOR U192 ( .A(n2473), .B(n68), .Z(out[1546]) );
  NANDN U193 ( .A(n4889), .B(n4665), .Z(n69) );
  XNOR U194 ( .A(n4888), .B(n69), .Z(out[872]) );
  NANDN U195 ( .A(n4897), .B(n4667), .Z(n70) );
  XNOR U196 ( .A(n4896), .B(n70), .Z(out[874]) );
  ANDN U197 ( .B(n5098), .A(n1699), .Z(n71) );
  XNOR U198 ( .A(n1871), .B(n71), .Z(out[1113]) );
  ANDN U199 ( .B(n4670), .A(n4908), .Z(n72) );
  XNOR U200 ( .A(n4909), .B(n72), .Z(out[876]) );
  ANDN U201 ( .B(n2648), .A(n2290), .Z(n73) );
  XNOR U202 ( .A(n2412), .B(n73), .Z(out[1396]) );
  ANDN U203 ( .B(n4673), .A(n4920), .Z(n74) );
  XNOR U204 ( .A(n4921), .B(n74), .Z(out[879]) );
  NAND U205 ( .A(n2575), .B(n2392), .Z(n75) );
  XNOR U206 ( .A(n2576), .B(n75), .Z(out[1507]) );
  AND U207 ( .A(n3015), .B(n3806), .Z(n76) );
  XNOR U208 ( .A(n3807), .B(n76), .Z(out[317]) );
  ANDN U209 ( .B(n4678), .A(n4928), .Z(n77) );
  XNOR U210 ( .A(n4929), .B(n77), .Z(out[881]) );
  ANDN U211 ( .B(n4679), .A(n4932), .Z(n78) );
  XNOR U212 ( .A(n4933), .B(n78), .Z(out[882]) );
  ANDN U213 ( .B(n2674), .A(n2303), .Z(n79) );
  XNOR U214 ( .A(n2422), .B(n79), .Z(out[1402]) );
  NANDN U215 ( .A(n1916), .B(n1765), .Z(n80) );
  XNOR U216 ( .A(n1915), .B(n80), .Z(out[1195]) );
  ANDN U217 ( .B(n5134), .A(n1736), .Z(n81) );
  XNOR U218 ( .A(n1891), .B(n81), .Z(out[1122]) );
  ANDN U219 ( .B(n4683), .A(n4952), .Z(n82) );
  XNOR U220 ( .A(n4953), .B(n82), .Z(out[886]) );
  NANDN U221 ( .A(n3637), .B(n3476), .Z(n83) );
  XNOR U222 ( .A(n3636), .B(n83), .Z(out[517]) );
  ANDN U223 ( .B(n1924), .A(n1517), .Z(n84) );
  XNOR U224 ( .A(n1766), .B(n84), .Z(out[1068]) );
  NANDN U225 ( .A(n2885), .B(n2884), .Z(n85) );
  XNOR U226 ( .A(n4340), .B(n85), .Z(out[268]) );
  NAND U227 ( .A(n2571), .B(n2391), .Z(n86) );
  XNOR U228 ( .A(n2572), .B(n86), .Z(out[1506]) );
  NANDN U229 ( .A(n4452), .B(n4867), .Z(n87) );
  XNOR U230 ( .A(n4649), .B(n87), .Z(out[738]) );
  OR U231 ( .A(n5093), .B(n5094), .Z(n88) );
  XNOR U232 ( .A(n5095), .B(n88), .Z(out[984]) );
  ANDN U233 ( .B(n2510), .A(n2220), .Z(n89) );
  XNOR U234 ( .A(n2361), .B(n89), .Z(out[1363]) );
  ANDN U235 ( .B(n2535), .A(n2233), .Z(n90) );
  XNOR U236 ( .A(n2373), .B(n90), .Z(out[1369]) );
  ANDN U237 ( .B(n2539), .A(n2235), .Z(n91) );
  XNOR U238 ( .A(n2375), .B(n91), .Z(out[1370]) );
  ANDN U239 ( .B(n2555), .A(n2243), .Z(n92) );
  XNOR U240 ( .A(n2384), .B(n92), .Z(out[1374]) );
  ANDN U241 ( .B(n2558), .A(n2245), .Z(n93) );
  XNOR U242 ( .A(n2386), .B(n93), .Z(out[1375]) );
  ANDN U243 ( .B(n2564), .A(n2248), .Z(n94) );
  XNOR U244 ( .A(n2388), .B(n94), .Z(out[1376]) );
  XNOR U245 ( .A(n1481), .B(n1136), .Z(n4054) );
  XNOR U246 ( .A(n1664), .B(n1665), .Z(n3061) );
  XNOR U247 ( .A(n1669), .B(n1670), .Z(n3063) );
  XNOR U248 ( .A(n1677), .B(n1678), .Z(n3068) );
  XNOR U249 ( .A(n570), .B(n687), .Z(n4049) );
  XNOR U250 ( .A(n1467), .B(n1090), .Z(n2864) );
  XNOR U251 ( .A(n1413), .B(n1690), .Z(n3175) );
  XNOR U252 ( .A(n1501), .B(n1237), .Z(n2213) );
  XNOR U253 ( .A(n1491), .B(n1192), .Z(n4074) );
  XNOR U254 ( .A(n1415), .B(n1694), .Z(n3177) );
  XNOR U255 ( .A(n1494), .B(n1207), .Z(n4078) );
  XNOR U256 ( .A(n1222), .B(n1497), .Z(n4082) );
  XOR U257 ( .A(n704), .B(n1487), .Z(n4538) );
  XNOR U258 ( .A(n1468), .B(n897), .Z(n4519) );
  XOR U259 ( .A(n1478), .B(n927), .Z(n4526) );
  XNOR U260 ( .A(n1424), .B(n1706), .Z(n3183) );
  XNOR U261 ( .A(n1453), .B(n1023), .Z(n2773) );
  XNOR U262 ( .A(n3966), .B(in[1487]), .Z(n4787) );
  AND U263 ( .A(n4763), .B(n4368), .Z(n95) );
  XNOR U264 ( .A(n4587), .B(n95), .Z(out[715]) );
  NANDN U265 ( .A(n4461), .B(n4879), .Z(n96) );
  XNOR U266 ( .A(n4658), .B(n96), .Z(out[741]) );
  ANDN U267 ( .B(n3511), .A(n3722), .Z(n97) );
  XNOR U268 ( .A(n3723), .B(n97), .Z(out[536]) );
  ANDN U269 ( .B(n1982), .A(n1575), .Z(n98) );
  XNOR U270 ( .A(n1798), .B(n98), .Z(out[1082]) );
  AND U271 ( .A(n2002), .B(n1593), .Z(n99) );
  XNOR U272 ( .A(n1808), .B(n99), .Z(out[1087]) );
  ANDN U273 ( .B(n3508), .A(n3704), .Z(n100) );
  XNOR U274 ( .A(n3705), .B(n100), .Z(out[533]) );
  ANDN U275 ( .B(n3857), .A(n3434), .Z(n101) );
  XNOR U276 ( .A(n3590), .B(n101), .Z(out[438]) );
  NOR U277 ( .A(n4699), .B(n4547), .Z(n102) );
  XNOR U278 ( .A(n4980), .B(n102), .Z(out[829]) );
  ANDN U279 ( .B(n1932), .A(n1525), .Z(n103) );
  XNOR U280 ( .A(n1770), .B(n103), .Z(out[1070]) );
  NOR U281 ( .A(n4702), .B(n4553), .Z(n104) );
  XNOR U282 ( .A(n4984), .B(n104), .Z(out[830]) );
  ANDN U283 ( .B(n1936), .A(n1529), .Z(n105) );
  XNOR U284 ( .A(n1772), .B(n105), .Z(out[1071]) );
  NOR U285 ( .A(n4556), .B(n4336), .Z(n106) );
  XNOR U286 ( .A(n4708), .B(n106), .Z(out[768]) );
  NOR U287 ( .A(n4559), .B(n4338), .Z(n107) );
  XNOR U288 ( .A(n4712), .B(n107), .Z(out[769]) );
  ANDN U289 ( .B(n1944), .A(n1537), .Z(n108) );
  XNOR U290 ( .A(n1778), .B(n108), .Z(out[1073]) );
  NOR U291 ( .A(n4562), .B(n4344), .Z(n109) );
  XNOR U292 ( .A(n4716), .B(n109), .Z(out[770]) );
  NOR U293 ( .A(n4565), .B(n4346), .Z(n110) );
  XNOR U294 ( .A(n4720), .B(n110), .Z(out[771]) );
  ANDN U295 ( .B(n1956), .A(n1551), .Z(n111) );
  XNOR U296 ( .A(n1784), .B(n111), .Z(out[1076]) );
  NANDN U297 ( .A(n2237), .B(n2543), .Z(n112) );
  XNOR U298 ( .A(n2377), .B(n112), .Z(out[1371]) );
  NOR U299 ( .A(n4574), .B(n4357), .Z(n113) );
  XNOR U300 ( .A(n4744), .B(n113), .Z(out[775]) );
  NAND U301 ( .A(n2898), .B(n4478), .Z(n114) );
  XNOR U302 ( .A(n2897), .B(n114), .Z(out[208]) );
  ANDN U303 ( .B(n5059), .A(n1654), .Z(n115) );
  XNOR U304 ( .A(n1847), .B(n115), .Z(out[1102]) );
  AND U305 ( .A(n5069), .B(n1666), .Z(n116) );
  XNOR U306 ( .A(n1853), .B(n116), .Z(out[1105]) );
  NANDN U307 ( .A(n4885), .B(n4664), .Z(n117) );
  XNOR U308 ( .A(n4884), .B(n117), .Z(out[871]) );
  ANDN U309 ( .B(n5089), .A(n1687), .Z(n118) );
  XNOR U310 ( .A(n1863), .B(n118), .Z(out[1110]) );
  ANDN U311 ( .B(n2481), .A(n2480), .Z(n119) );
  XNOR U312 ( .A(n2479), .B(n119), .Z(out[1548]) );
  ANDN U313 ( .B(n5092), .A(n1691), .Z(n120) );
  XNOR U314 ( .A(n1865), .B(n120), .Z(out[1111]) );
  ANDN U315 ( .B(n5101), .A(n1703), .Z(n121) );
  XNOR U316 ( .A(n1873), .B(n121), .Z(out[1114]) );
  ANDN U317 ( .B(n5108), .A(n1712), .Z(n122) );
  XNOR U318 ( .A(n1877), .B(n122), .Z(out[1116]) );
  ANDN U319 ( .B(n2652), .A(n2292), .Z(n123) );
  XNOR U320 ( .A(n2414), .B(n123), .Z(out[1397]) );
  ANDN U321 ( .B(n4677), .A(n4924), .Z(n124) );
  XNOR U322 ( .A(n4925), .B(n124), .Z(out[880]) );
  AND U323 ( .A(n4767), .B(n4375), .Z(n125) );
  XNOR U324 ( .A(n4589), .B(n125), .Z(out[716]) );
  NAND U325 ( .A(n2583), .B(n2394), .Z(n126) );
  XNOR U326 ( .A(n2584), .B(n126), .Z(out[1509]) );
  ANDN U327 ( .B(n4680), .A(n4936), .Z(n127) );
  XNOR U328 ( .A(n4937), .B(n127), .Z(out[883]) );
  ANDN U329 ( .B(n4681), .A(n4940), .Z(n128) );
  XNOR U330 ( .A(n4941), .B(n128), .Z(out[884]) );
  ANDN U331 ( .B(n4682), .A(n4944), .Z(n129) );
  XNOR U332 ( .A(n4945), .B(n129), .Z(out[885]) );
  ANDN U333 ( .B(n1906), .A(n1499), .Z(n130) );
  XNOR U334 ( .A(n1759), .B(n130), .Z(out[1064]) );
  NAND U335 ( .A(n3475), .B(n3633), .Z(n131) );
  XNOR U336 ( .A(n3632), .B(n131), .Z(out[516]) );
  OR U337 ( .A(n5021), .B(n1830), .Z(n132) );
  XNOR U338 ( .A(n5020), .B(n132), .Z(out[1222]) );
  ANDN U339 ( .B(n1910), .A(n1503), .Z(n133) );
  XNOR U340 ( .A(n1761), .B(n133), .Z(out[1065]) );
  NANDN U341 ( .A(n1513), .B(n1918), .Z(n134) );
  XNOR U342 ( .A(n1765), .B(n134), .Z(out[1067]) );
  NANDN U343 ( .A(n4414), .B(n4823), .Z(n135) );
  XNOR U344 ( .A(n4620), .B(n135), .Z(out[728]) );
  NANDN U345 ( .A(n4417), .B(n4827), .Z(n136) );
  XNOR U346 ( .A(n4623), .B(n136), .Z(out[729]) );
  NANDN U347 ( .A(n2883), .B(n2882), .Z(n137) );
  XNOR U348 ( .A(n4308), .B(n137), .Z(out[267]) );
  ANDN U349 ( .B(n1928), .A(n1521), .Z(n138) );
  XNOR U350 ( .A(n1768), .B(n138), .Z(out[1069]) );
  ANDN U351 ( .B(n4831), .A(n4420), .Z(n139) );
  XNOR U352 ( .A(n4626), .B(n139), .Z(out[730]) );
  NANDN U353 ( .A(n2887), .B(n2886), .Z(n140) );
  XNOR U354 ( .A(n4371), .B(n140), .Z(out[269]) );
  NANDN U355 ( .A(n4429), .B(n4843), .Z(n141) );
  XNOR U356 ( .A(n4636), .B(n141), .Z(out[733]) );
  AND U357 ( .A(n2655), .B(n2416), .Z(n142) );
  XNOR U358 ( .A(n2656), .B(n142), .Z(out[1526]) );
  NANDN U359 ( .A(n4432), .B(n4847), .Z(n143) );
  XNOR U360 ( .A(n4639), .B(n143), .Z(out[734]) );
  NANDN U361 ( .A(n4435), .B(n4851), .Z(n144) );
  XNOR U362 ( .A(n4642), .B(n144), .Z(out[735]) );
  OR U363 ( .A(n5084), .B(n5085), .Z(n145) );
  XNOR U364 ( .A(n5086), .B(n145), .Z(out[981]) );
  NANDN U365 ( .A(n2211), .B(n2492), .Z(n146) );
  XNOR U366 ( .A(n2353), .B(n146), .Z(out[1359]) );
  NAND U367 ( .A(n3939), .B(n3938), .Z(n147) );
  XNOR U368 ( .A(n3940), .B(n147), .Z(out[64]) );
  NANDN U369 ( .A(n2214), .B(n2498), .Z(n148) );
  XNOR U370 ( .A(n2355), .B(n148), .Z(out[1360]) );
  NANDN U371 ( .A(n3982), .B(n3981), .Z(n149) );
  XNOR U372 ( .A(n3983), .B(n149), .Z(out[65]) );
  ANDN U373 ( .B(n2502), .A(n2216), .Z(n150) );
  XNOR U374 ( .A(n2356), .B(n150), .Z(out[1361]) );
  OR U375 ( .A(n5096), .B(n5097), .Z(n151) );
  XNOR U376 ( .A(n5098), .B(n151), .Z(out[985]) );
  ANDN U377 ( .B(n2514), .A(n2222), .Z(n152) );
  XNOR U378 ( .A(n2363), .B(n152), .Z(out[1364]) );
  OR U379 ( .A(n5109), .B(n5110), .Z(n153) );
  XNOR U380 ( .A(n5111), .B(n153), .Z(out[989]) );
  OR U381 ( .A(n5116), .B(n5117), .Z(n154) );
  XNOR U382 ( .A(n5118), .B(n154), .Z(out[990]) );
  ANDN U383 ( .B(n3515), .A(n3734), .Z(n155) );
  XNOR U384 ( .A(n3735), .B(n155), .Z(out[539]) );
  NANDN U385 ( .A(n2853), .B(n3897), .Z(n156) );
  XNOR U386 ( .A(n3019), .B(n156), .Z(out[191]) );
  XNOR U387 ( .A(n1681), .B(n1682), .Z(n3071) );
  XNOR U388 ( .A(n1693), .B(n1694), .Z(n3079) );
  XNOR U389 ( .A(n1697), .B(n1698), .Z(n3081) );
  XNOR U390 ( .A(n1483), .B(n1149), .Z(n4058) );
  XNOR U391 ( .A(n1722), .B(n1723), .Z(n3092) );
  XNOR U392 ( .A(n1726), .B(n1727), .Z(n3094) );
  XNOR U393 ( .A(n1730), .B(n1731), .Z(n3098) );
  XNOR U394 ( .A(n1441), .B(n1743), .Z(n3208) );
  XOR U395 ( .A(n1446), .B(n751), .Z(n4488) );
  XNOR U396 ( .A(n3958), .B(in[1485]), .Z(n4779) );
  XNOR U397 ( .A(n3974), .B(in[1489]), .Z(n4795) );
  XNOR U398 ( .A(n3978), .B(in[1490]), .Z(n4799) );
  XNOR U399 ( .A(n3935), .B(in[1480]), .Z(n4755) );
  XNOR U400 ( .A(n3942), .B(in[1481]), .Z(n4759) );
  NAND U401 ( .A(n4747), .B(n4357), .Z(n157) );
  XNOR U402 ( .A(n4574), .B(n157), .Z(out[711]) );
  NAND U403 ( .A(n2587), .B(n2396), .Z(n158) );
  XNOR U404 ( .A(n2588), .B(n158), .Z(out[1510]) );
  AND U405 ( .A(n2591), .B(n2397), .Z(n159) );
  XNOR U406 ( .A(n2592), .B(n159), .Z(out[1511]) );
  AND U407 ( .A(n2595), .B(n2398), .Z(n160) );
  XNOR U408 ( .A(n2596), .B(n160), .Z(out[1512]) );
  ANDN U409 ( .B(n1986), .A(n1579), .Z(n161) );
  XNOR U410 ( .A(n1800), .B(n161), .Z(out[1083]) );
  NOR U411 ( .A(n4597), .B(n4387), .Z(n162) );
  XNOR U412 ( .A(n4785), .B(n162), .Z(out[784]) );
  ANDN U413 ( .B(n3849), .A(n3431), .Z(n163) );
  XNOR U414 ( .A(n3588), .B(n163), .Z(out[437]) );
  ANDN U415 ( .B(n3865), .A(n3440), .Z(n164) );
  XNOR U416 ( .A(n3594), .B(n164), .Z(out[440]) );
  NAND U417 ( .A(n3602), .B(n3871), .Z(n165) );
  XNOR U418 ( .A(n3870), .B(n165), .Z(out[570]) );
  NOR U419 ( .A(n4705), .B(n4555), .Z(n166) );
  XNOR U420 ( .A(n4988), .B(n166), .Z(out[831]) );
  ANDN U421 ( .B(n2547), .A(n2239), .Z(n167) );
  XNOR U422 ( .A(n2380), .B(n167), .Z(out[1372]) );
  ANDN U423 ( .B(n2551), .A(n2241), .Z(n168) );
  XNOR U424 ( .A(n2382), .B(n168), .Z(out[1373]) );
  NAND U425 ( .A(n2904), .B(n4551), .Z(n169) );
  XNOR U426 ( .A(n2903), .B(n169), .Z(out[210]) );
  NAND U427 ( .A(n2907), .B(n4580), .Z(n170) );
  XNOR U428 ( .A(n2906), .B(n170), .Z(out[211]) );
  NAND U429 ( .A(n2910), .B(n4605), .Z(n171) );
  XNOR U430 ( .A(n2909), .B(n171), .Z(out[212]) );
  NANDN U431 ( .A(n2916), .B(n4662), .Z(n172) );
  XNOR U432 ( .A(n2915), .B(n172), .Z(out[214]) );
  NANDN U433 ( .A(n2928), .B(n4727), .Z(n173) );
  XNOR U434 ( .A(n2927), .B(n173), .Z(out[217]) );
  NANDN U435 ( .A(n2931), .B(n4775), .Z(n174) );
  XNOR U436 ( .A(n2930), .B(n174), .Z(out[218]) );
  ANDN U437 ( .B(n5047), .A(n1642), .Z(n175) );
  XNOR U438 ( .A(n1839), .B(n175), .Z(out[1099]) );
  AND U439 ( .A(n5063), .B(n1658), .Z(n176) );
  XNOR U440 ( .A(n1849), .B(n176), .Z(out[1103]) );
  ANDN U441 ( .B(n5076), .A(n1675), .Z(n177) );
  XNOR U442 ( .A(n1857), .B(n177), .Z(out[1107]) );
  ANDN U443 ( .B(n5086), .A(n1683), .Z(n178) );
  XNOR U444 ( .A(n1861), .B(n178), .Z(out[1109]) );
  NANDN U445 ( .A(n4893), .B(n4666), .Z(n179) );
  XNOR U446 ( .A(n4892), .B(n179), .Z(out[873]) );
  ANDN U447 ( .B(n5095), .A(n1695), .Z(n180) );
  XNOR U448 ( .A(n1869), .B(n180), .Z(out[1112]) );
  ANDN U449 ( .B(n2484), .A(n2483), .Z(n181) );
  XNOR U450 ( .A(n2482), .B(n181), .Z(out[1549]) );
  ANDN U451 ( .B(n2644), .A(n2287), .Z(n182) );
  XNOR U452 ( .A(n2410), .B(n182), .Z(out[1395]) );
  ANDN U453 ( .B(n5111), .A(n1716), .Z(n183) );
  XNOR U454 ( .A(n1879), .B(n183), .Z(out[1117]) );
  NAND U455 ( .A(n3603), .B(n3875), .Z(n184) );
  XNOR U456 ( .A(n3874), .B(n184), .Z(out[571]) );
  NAND U457 ( .A(n2579), .B(n2393), .Z(n185) );
  XNOR U458 ( .A(n2580), .B(n185), .Z(out[1508]) );
  ANDN U459 ( .B(n2670), .A(n2301), .Z(n186) );
  XNOR U460 ( .A(n2419), .B(n186), .Z(out[1401]) );
  AND U461 ( .A(n2495), .B(n2355), .Z(n187) );
  XNOR U462 ( .A(n2496), .B(n187), .Z(out[1488]) );
  ANDN U463 ( .B(n2403), .A(n2617), .Z(n188) );
  XNOR U464 ( .A(n2618), .B(n188), .Z(out[1517]) );
  ANDN U465 ( .B(n1914), .A(n1509), .Z(n189) );
  XNOR U466 ( .A(n1763), .B(n189), .Z(out[1066]) );
  NANDN U467 ( .A(n3645), .B(n3478), .Z(n190) );
  XNOR U468 ( .A(n3644), .B(n190), .Z(out[519]) );
  NAND U469 ( .A(n2540), .B(n2377), .Z(n191) );
  XNOR U470 ( .A(n2541), .B(n191), .Z(out[1499]) );
  OR U471 ( .A(n5064), .B(n5065), .Z(n192) );
  XNOR U472 ( .A(n5066), .B(n192), .Z(out[976]) );
  OR U473 ( .A(n5067), .B(n5068), .Z(n193) );
  XNOR U474 ( .A(n5069), .B(n193), .Z(out[977]) );
  OR U475 ( .A(n5070), .B(n5071), .Z(n194) );
  XNOR U476 ( .A(n5072), .B(n194), .Z(out[978]) );
  NAND U477 ( .A(n2565), .B(n2390), .Z(n195) );
  XNOR U478 ( .A(n2566), .B(n195), .Z(out[1505]) );
  AND U479 ( .A(n2663), .B(n2418), .Z(n196) );
  XNOR U480 ( .A(n2664), .B(n196), .Z(out[1528]) );
  NANDN U481 ( .A(n4446), .B(n4855), .Z(n197) );
  XNOR U482 ( .A(n4643), .B(n197), .Z(out[736]) );
  OR U483 ( .A(n5081), .B(n5082), .Z(n198) );
  XNOR U484 ( .A(n5083), .B(n198), .Z(out[980]) );
  NANDN U485 ( .A(n4449), .B(n4859), .Z(n199) );
  XNOR U486 ( .A(n4646), .B(n199), .Z(out[737]) );
  OR U487 ( .A(n5087), .B(n5088), .Z(n200) );
  XNOR U488 ( .A(n5089), .B(n200), .Z(out[982]) );
  NANDN U489 ( .A(n4455), .B(n4871), .Z(n201) );
  XNOR U490 ( .A(n4652), .B(n201), .Z(out[739]) );
  OR U491 ( .A(n5090), .B(n5091), .Z(n202) );
  XNOR U492 ( .A(n5092), .B(n202), .Z(out[983]) );
  OR U493 ( .A(n5099), .B(n5100), .Z(n203) );
  XNOR U494 ( .A(n5101), .B(n203), .Z(out[986]) );
  OR U495 ( .A(n5102), .B(n5103), .Z(n204) );
  XNOR U496 ( .A(n5104), .B(n204), .Z(out[987]) );
  NAND U497 ( .A(n2603), .B(n2400), .Z(n205) );
  XNOR U498 ( .A(n2604), .B(n205), .Z(out[1514]) );
  AND U499 ( .A(n2607), .B(n2401), .Z(n206) );
  XNOR U500 ( .A(n2608), .B(n206), .Z(out[1515]) );
  ANDN U501 ( .B(n1990), .A(n1583), .Z(n207) );
  XNOR U502 ( .A(n1802), .B(n207), .Z(out[1084]) );
  AND U503 ( .A(n2613), .B(n2402), .Z(n208) );
  XNOR U504 ( .A(n2614), .B(n208), .Z(out[1516]) );
  ANDN U505 ( .B(n1994), .A(n1587), .Z(n209) );
  XNOR U506 ( .A(n1804), .B(n209), .Z(out[1085]) );
  AND U507 ( .A(n2621), .B(n2404), .Z(n210) );
  XNOR U508 ( .A(n2622), .B(n210), .Z(out[1518]) );
  ANDN U509 ( .B(n2531), .A(n2231), .Z(n211) );
  XNOR U510 ( .A(n2371), .B(n211), .Z(out[1368]) );
  AND U511 ( .A(n2625), .B(n2405), .Z(n212) );
  XNOR U512 ( .A(n2626), .B(n212), .Z(out[1519]) );
  ANDN U513 ( .B(n4999), .A(n1597), .Z(n213) );
  XNOR U514 ( .A(n1811), .B(n213), .Z(out[1088]) );
  AND U515 ( .A(n2629), .B(n2407), .Z(n214) );
  XNOR U516 ( .A(n2630), .B(n214), .Z(out[1520]) );
  ANDN U517 ( .B(n5003), .A(n1601), .Z(n215) );
  XNOR U518 ( .A(n1814), .B(n215), .Z(out[1089]) );
  AND U519 ( .A(n2633), .B(n2408), .Z(n216) );
  XNOR U520 ( .A(n2634), .B(n216), .Z(out[1521]) );
  ANDN U521 ( .B(n5007), .A(n1605), .Z(n217) );
  XNOR U522 ( .A(n1817), .B(n217), .Z(out[1090]) );
  AND U523 ( .A(n2637), .B(n2409), .Z(n218) );
  XNOR U524 ( .A(n2638), .B(n218), .Z(out[1522]) );
  ANDN U525 ( .B(n5011), .A(n1609), .Z(n219) );
  XNOR U526 ( .A(n1820), .B(n219), .Z(out[1091]) );
  ANDN U527 ( .B(n5015), .A(n1613), .Z(n220) );
  XNOR U528 ( .A(n1825), .B(n220), .Z(out[1092]) );
  ANDN U529 ( .B(n5019), .A(n1617), .Z(n221) );
  XNOR U530 ( .A(n1828), .B(n221), .Z(out[1093]) );
  NANDN U531 ( .A(n2849), .B(n3809), .Z(n222) );
  XNOR U532 ( .A(n3015), .B(n222), .Z(out[189]) );
  ANDN U533 ( .B(n5023), .A(n1621), .Z(n223) );
  XNOR U534 ( .A(n1830), .B(n223), .Z(out[1094]) );
  NANDN U535 ( .A(n2851), .B(n3853), .Z(n224) );
  XNOR U536 ( .A(n3016), .B(n224), .Z(out[190]) );
  ANDN U537 ( .B(n5027), .A(n1625), .Z(n225) );
  XNOR U538 ( .A(n1831), .B(n225), .Z(out[1095]) );
  AND U539 ( .A(n2659), .B(n2417), .Z(n226) );
  XNOR U540 ( .A(n2660), .B(n226), .Z(out[1527]) );
  ANDN U541 ( .B(n5031), .A(n1630), .Z(n227) );
  XNOR U542 ( .A(n1833), .B(n227), .Z(out[1096]) );
  ANDN U543 ( .B(n5035), .A(n1634), .Z(n228) );
  XNOR U544 ( .A(n1835), .B(n228), .Z(out[1097]) );
  NANDN U545 ( .A(n2252), .B(n2574), .Z(n229) );
  XNOR U546 ( .A(n2391), .B(n229), .Z(out[1378]) );
  ANDN U547 ( .B(n5043), .A(n1638), .Z(n230) );
  XNOR U548 ( .A(n1837), .B(n230), .Z(out[1098]) );
  NAND U549 ( .A(n2491), .B(n2353), .Z(n231) );
  XNOR U550 ( .A(n2490), .B(n231), .Z(out[1487]) );
  XNOR U551 ( .A(in[1168]), .B(n934), .Z(n232) );
  XNOR U552 ( .A(in[545]), .B(n1176), .Z(n233) );
  XOR U553 ( .A(in[1469]), .B(in[509]), .Z(n235) );
  XNOR U554 ( .A(in[829]), .B(in[189]), .Z(n234) );
  XNOR U555 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U556 ( .A(in[1149]), .B(n236), .Z(n1105) );
  XOR U557 ( .A(in[1598]), .B(in[638]), .Z(n238) );
  XNOR U558 ( .A(in[958]), .B(in[318]), .Z(n237) );
  XNOR U559 ( .A(n238), .B(n237), .Z(n239) );
  XNOR U560 ( .A(in[1278]), .B(n239), .Z(n1674) );
  XNOR U561 ( .A(n1105), .B(n1674), .Z(n3288) );
  XOR U562 ( .A(in[254]), .B(n3288), .Z(n3938) );
  XOR U563 ( .A(in[1345]), .B(in[65]), .Z(n241) );
  XNOR U564 ( .A(in[1025]), .B(in[385]), .Z(n240) );
  XNOR U565 ( .A(n241), .B(n240), .Z(n242) );
  XNOR U566 ( .A(in[705]), .B(n242), .Z(n1682) );
  XOR U567 ( .A(in[1474]), .B(in[514]), .Z(n244) );
  XNOR U568 ( .A(in[834]), .B(in[194]), .Z(n243) );
  XNOR U569 ( .A(n244), .B(n243), .Z(n245) );
  XOR U570 ( .A(in[1154]), .B(n245), .Z(n1407) );
  XOR U571 ( .A(in[1410]), .B(n3171), .Z(n3939) );
  XOR U572 ( .A(in[137]), .B(in[457]), .Z(n247) );
  XNOR U573 ( .A(in[777]), .B(in[1417]), .Z(n246) );
  XNOR U574 ( .A(n247), .B(n246), .Z(n248) );
  XNOR U575 ( .A(in[1097]), .B(n248), .Z(n1364) );
  XOR U576 ( .A(in[328]), .B(in[8]), .Z(n250) );
  XNOR U577 ( .A(in[968]), .B(in[648]), .Z(n249) );
  XNOR U578 ( .A(n250), .B(n249), .Z(n251) );
  XNOR U579 ( .A(in[1288]), .B(n251), .Z(n1420) );
  XOR U580 ( .A(n1364), .B(n1420), .Z(n4451) );
  XNOR U581 ( .A(in[1033]), .B(n4451), .Z(n2856) );
  OR U582 ( .A(n3939), .B(n2856), .Z(n252) );
  XOR U583 ( .A(n3938), .B(n252), .Z(out[0]) );
  XOR U584 ( .A(in[1386]), .B(in[106]), .Z(n254) );
  XNOR U585 ( .A(in[1066]), .B(in[746]), .Z(n253) );
  XNOR U586 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U587 ( .A(in[426]), .B(n255), .Z(n708) );
  XOR U588 ( .A(in[1515]), .B(in[555]), .Z(n257) );
  XNOR U589 ( .A(in[875]), .B(in[235]), .Z(n256) );
  XNOR U590 ( .A(n257), .B(n256), .Z(n258) );
  XNOR U591 ( .A(in[1195]), .B(n258), .Z(n1528) );
  XOR U592 ( .A(n708), .B(n1528), .Z(n4109) );
  XOR U593 ( .A(in[171]), .B(n4109), .Z(n1499) );
  XOR U594 ( .A(in[971]), .B(in[1291]), .Z(n260) );
  XNOR U595 ( .A(in[11]), .B(in[331]), .Z(n259) );
  XNOR U596 ( .A(n260), .B(n259), .Z(n261) );
  XNOR U597 ( .A(in[651]), .B(n261), .Z(n1429) );
  XOR U598 ( .A(in[140]), .B(in[460]), .Z(n263) );
  XNOR U599 ( .A(in[1100]), .B(in[1420]), .Z(n262) );
  XNOR U600 ( .A(n263), .B(n262), .Z(n264) );
  XOR U601 ( .A(in[780]), .B(n264), .Z(n1386) );
  XNOR U602 ( .A(in[1356]), .B(n4460), .Z(n1906) );
  XOR U603 ( .A(in[1364]), .B(in[724]), .Z(n266) );
  XNOR U604 ( .A(in[84]), .B(in[404]), .Z(n265) );
  XNOR U605 ( .A(n266), .B(n265), .Z(n267) );
  XNOR U606 ( .A(in[1044]), .B(n267), .Z(n1010) );
  XOR U607 ( .A(in[1555]), .B(in[595]), .Z(n269) );
  XNOR U608 ( .A(in[915]), .B(in[275]), .Z(n268) );
  XNOR U609 ( .A(n269), .B(n268), .Z(n270) );
  XNOR U610 ( .A(in[1235]), .B(n270), .Z(n722) );
  XOR U611 ( .A(n1010), .B(n722), .Z(n4248) );
  XOR U612 ( .A(in[980]), .B(n4248), .Z(n1903) );
  NANDN U613 ( .A(n1906), .B(n1903), .Z(n271) );
  XNOR U614 ( .A(n1499), .B(n271), .Z(out[1000]) );
  XOR U615 ( .A(in[1387]), .B(in[107]), .Z(n273) );
  XNOR U616 ( .A(in[1067]), .B(in[747]), .Z(n272) );
  XNOR U617 ( .A(n273), .B(n272), .Z(n274) );
  XNOR U618 ( .A(in[427]), .B(n274), .Z(n719) );
  XOR U619 ( .A(in[1516]), .B(in[556]), .Z(n276) );
  XNOR U620 ( .A(in[876]), .B(in[236]), .Z(n275) );
  XNOR U621 ( .A(n276), .B(n275), .Z(n277) );
  XNOR U622 ( .A(in[1196]), .B(n277), .Z(n1532) );
  XOR U623 ( .A(n719), .B(n1532), .Z(n4117) );
  XOR U624 ( .A(in[172]), .B(n4117), .Z(n1503) );
  XOR U625 ( .A(in[972]), .B(in[12]), .Z(n279) );
  XNOR U626 ( .A(in[1292]), .B(in[332]), .Z(n278) );
  XNOR U627 ( .A(n279), .B(n278), .Z(n280) );
  XNOR U628 ( .A(in[652]), .B(n280), .Z(n1431) );
  XOR U629 ( .A(in[141]), .B(in[461]), .Z(n282) );
  XNOR U630 ( .A(in[1101]), .B(in[1421]), .Z(n281) );
  XNOR U631 ( .A(n282), .B(n281), .Z(n283) );
  XOR U632 ( .A(in[781]), .B(n283), .Z(n1390) );
  XNOR U633 ( .A(in[1357]), .B(n4463), .Z(n1910) );
  XOR U634 ( .A(in[1365]), .B(in[725]), .Z(n285) );
  XNOR U635 ( .A(in[85]), .B(in[405]), .Z(n284) );
  XNOR U636 ( .A(n285), .B(n284), .Z(n286) );
  XNOR U637 ( .A(in[1045]), .B(n286), .Z(n1023) );
  XOR U638 ( .A(in[1556]), .B(in[596]), .Z(n288) );
  XNOR U639 ( .A(in[916]), .B(in[276]), .Z(n287) );
  XNOR U640 ( .A(n288), .B(n287), .Z(n289) );
  XNOR U641 ( .A(in[1236]), .B(n289), .Z(n737) );
  XOR U642 ( .A(n1023), .B(n737), .Z(n4251) );
  XOR U643 ( .A(in[981]), .B(n4251), .Z(n1907) );
  NANDN U644 ( .A(n1910), .B(n1907), .Z(n290) );
  XNOR U645 ( .A(n1503), .B(n290), .Z(out[1001]) );
  XOR U646 ( .A(in[1388]), .B(in[108]), .Z(n292) );
  XNOR U647 ( .A(in[1068]), .B(in[748]), .Z(n291) );
  XNOR U648 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U649 ( .A(in[428]), .B(n293), .Z(n1596) );
  XOR U650 ( .A(in[1517]), .B(in[557]), .Z(n295) );
  XNOR U651 ( .A(in[877]), .B(in[237]), .Z(n294) );
  XNOR U652 ( .A(n295), .B(n294), .Z(n296) );
  XNOR U653 ( .A(in[1197]), .B(n296), .Z(n1536) );
  XOR U654 ( .A(n1596), .B(n1536), .Z(n1369) );
  XOR U655 ( .A(in[173]), .B(n1369), .Z(n1509) );
  XOR U656 ( .A(in[973]), .B(in[13]), .Z(n298) );
  XNOR U657 ( .A(in[1293]), .B(in[333]), .Z(n297) );
  XNOR U658 ( .A(n298), .B(n297), .Z(n299) );
  XNOR U659 ( .A(in[653]), .B(n299), .Z(n1433) );
  XOR U660 ( .A(in[142]), .B(in[1422]), .Z(n301) );
  XNOR U661 ( .A(in[1102]), .B(in[782]), .Z(n300) );
  XNOR U662 ( .A(n301), .B(n300), .Z(n302) );
  XOR U663 ( .A(in[462]), .B(n302), .Z(n1394) );
  XNOR U664 ( .A(in[1358]), .B(n4466), .Z(n1914) );
  XOR U665 ( .A(in[1366]), .B(in[726]), .Z(n304) );
  XNOR U666 ( .A(in[86]), .B(in[406]), .Z(n303) );
  XNOR U667 ( .A(n304), .B(n303), .Z(n305) );
  XNOR U668 ( .A(in[1046]), .B(n305), .Z(n1036) );
  XOR U669 ( .A(in[1557]), .B(in[597]), .Z(n307) );
  XNOR U670 ( .A(in[917]), .B(in[277]), .Z(n306) );
  XNOR U671 ( .A(n307), .B(n306), .Z(n308) );
  XNOR U672 ( .A(in[1237]), .B(n308), .Z(n752) );
  XOR U673 ( .A(n1036), .B(n752), .Z(n4252) );
  XOR U674 ( .A(in[982]), .B(n4252), .Z(n1911) );
  NANDN U675 ( .A(n1914), .B(n1911), .Z(n309) );
  XNOR U676 ( .A(n1509), .B(n309), .Z(out[1002]) );
  XOR U677 ( .A(in[1389]), .B(in[109]), .Z(n311) );
  XNOR U678 ( .A(in[1069]), .B(in[749]), .Z(n310) );
  XNOR U679 ( .A(n311), .B(n310), .Z(n312) );
  XNOR U680 ( .A(in[429]), .B(n312), .Z(n1600) );
  XOR U681 ( .A(in[1518]), .B(in[558]), .Z(n314) );
  XNOR U682 ( .A(in[878]), .B(in[238]), .Z(n313) );
  XNOR U683 ( .A(n314), .B(n313), .Z(n315) );
  XNOR U684 ( .A(in[1198]), .B(n315), .Z(n1540) );
  XOR U685 ( .A(n1600), .B(n1540), .Z(n1409) );
  XOR U686 ( .A(in[174]), .B(n1409), .Z(n1513) );
  XOR U687 ( .A(in[974]), .B(in[14]), .Z(n317) );
  XNOR U688 ( .A(in[1294]), .B(in[334]), .Z(n316) );
  XNOR U689 ( .A(n317), .B(n316), .Z(n318) );
  XNOR U690 ( .A(in[654]), .B(n318), .Z(n1435) );
  XOR U691 ( .A(in[143]), .B(in[1423]), .Z(n320) );
  XNOR U692 ( .A(in[1103]), .B(in[783]), .Z(n319) );
  XNOR U693 ( .A(n320), .B(n319), .Z(n321) );
  XOR U694 ( .A(in[463]), .B(n321), .Z(n1398) );
  XNOR U695 ( .A(in[1359]), .B(n4469), .Z(n1918) );
  XOR U696 ( .A(in[1367]), .B(in[727]), .Z(n323) );
  XNOR U697 ( .A(in[87]), .B(in[407]), .Z(n322) );
  XNOR U698 ( .A(n323), .B(n322), .Z(n324) );
  XNOR U699 ( .A(in[1047]), .B(n324), .Z(n1049) );
  XOR U700 ( .A(in[1558]), .B(in[598]), .Z(n326) );
  XNOR U701 ( .A(in[918]), .B(in[278]), .Z(n325) );
  XNOR U702 ( .A(n326), .B(n325), .Z(n327) );
  XNOR U703 ( .A(in[1238]), .B(n327), .Z(n767) );
  XOR U704 ( .A(n1049), .B(n767), .Z(n4253) );
  XOR U705 ( .A(in[983]), .B(n4253), .Z(n1915) );
  NANDN U706 ( .A(n1918), .B(n1915), .Z(n328) );
  XNOR U707 ( .A(n1513), .B(n328), .Z(out[1003]) );
  XOR U708 ( .A(in[1390]), .B(in[110]), .Z(n330) );
  XNOR U709 ( .A(in[1070]), .B(in[750]), .Z(n329) );
  XNOR U710 ( .A(n330), .B(n329), .Z(n331) );
  XNOR U711 ( .A(in[430]), .B(n331), .Z(n1604) );
  XOR U712 ( .A(in[1519]), .B(in[559]), .Z(n333) );
  XNOR U713 ( .A(in[879]), .B(in[239]), .Z(n332) );
  XNOR U714 ( .A(n333), .B(n332), .Z(n334) );
  XNOR U715 ( .A(in[1199]), .B(n334), .Z(n1544) );
  XOR U716 ( .A(n1604), .B(n1544), .Z(n1421) );
  XOR U717 ( .A(in[175]), .B(n1421), .Z(n1517) );
  XOR U718 ( .A(in[144]), .B(in[1424]), .Z(n336) );
  XNOR U719 ( .A(in[1104]), .B(in[784]), .Z(n335) );
  XNOR U720 ( .A(n336), .B(n335), .Z(n337) );
  XNOR U721 ( .A(in[464]), .B(n337), .Z(n1402) );
  XOR U722 ( .A(in[975]), .B(in[15]), .Z(n339) );
  XNOR U723 ( .A(in[1295]), .B(in[335]), .Z(n338) );
  XNOR U724 ( .A(n339), .B(n338), .Z(n340) );
  XOR U725 ( .A(in[655]), .B(n340), .Z(n1437) );
  XNOR U726 ( .A(in[1360]), .B(n4472), .Z(n1924) );
  XOR U727 ( .A(in[1368]), .B(in[728]), .Z(n342) );
  XNOR U728 ( .A(in[88]), .B(in[408]), .Z(n341) );
  XNOR U729 ( .A(n342), .B(n341), .Z(n343) );
  XNOR U730 ( .A(in[1048]), .B(n343), .Z(n1062) );
  XOR U731 ( .A(in[1559]), .B(in[599]), .Z(n345) );
  XNOR U732 ( .A(in[919]), .B(in[279]), .Z(n344) );
  XNOR U733 ( .A(n345), .B(n344), .Z(n346) );
  XNOR U734 ( .A(in[1239]), .B(n346), .Z(n782) );
  XOR U735 ( .A(n1062), .B(n782), .Z(n4254) );
  XOR U736 ( .A(in[984]), .B(n4254), .Z(n1921) );
  NANDN U737 ( .A(n1924), .B(n1921), .Z(n347) );
  XNOR U738 ( .A(n1517), .B(n347), .Z(out[1004]) );
  XOR U739 ( .A(in[1391]), .B(in[111]), .Z(n349) );
  XNOR U740 ( .A(in[1071]), .B(in[751]), .Z(n348) );
  XNOR U741 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U742 ( .A(in[431]), .B(n350), .Z(n1608) );
  XOR U743 ( .A(in[1520]), .B(in[560]), .Z(n352) );
  XNOR U744 ( .A(in[880]), .B(in[240]), .Z(n351) );
  XNOR U745 ( .A(n352), .B(n351), .Z(n353) );
  XNOR U746 ( .A(in[1200]), .B(n353), .Z(n1550) );
  XOR U747 ( .A(n1608), .B(n1550), .Z(n1443) );
  XOR U748 ( .A(in[176]), .B(n1443), .Z(n1521) );
  XOR U749 ( .A(in[145]), .B(in[1425]), .Z(n355) );
  XNOR U750 ( .A(in[1105]), .B(in[785]), .Z(n354) );
  XNOR U751 ( .A(n355), .B(n354), .Z(n356) );
  XNOR U752 ( .A(in[465]), .B(n356), .Z(n1406) );
  XOR U753 ( .A(in[976]), .B(in[16]), .Z(n358) );
  XNOR U754 ( .A(in[1296]), .B(in[336]), .Z(n357) );
  XNOR U755 ( .A(n358), .B(n357), .Z(n359) );
  XOR U756 ( .A(in[656]), .B(n359), .Z(n1439) );
  XNOR U757 ( .A(in[1361]), .B(n4479), .Z(n1928) );
  XOR U758 ( .A(in[1369]), .B(in[729]), .Z(n361) );
  XNOR U759 ( .A(in[89]), .B(in[409]), .Z(n360) );
  XNOR U760 ( .A(n361), .B(n360), .Z(n362) );
  XNOR U761 ( .A(in[1049]), .B(n362), .Z(n1075) );
  XOR U762 ( .A(in[1560]), .B(in[600]), .Z(n364) );
  XNOR U763 ( .A(in[920]), .B(in[280]), .Z(n363) );
  XNOR U764 ( .A(n364), .B(n363), .Z(n365) );
  XNOR U765 ( .A(in[1240]), .B(n365), .Z(n797) );
  XOR U766 ( .A(n1075), .B(n797), .Z(n4255) );
  XOR U767 ( .A(in[985]), .B(n4255), .Z(n1925) );
  NANDN U768 ( .A(n1928), .B(n1925), .Z(n366) );
  XNOR U769 ( .A(n1521), .B(n366), .Z(out[1005]) );
  XOR U770 ( .A(in[1392]), .B(in[112]), .Z(n368) );
  XNOR U771 ( .A(in[1072]), .B(in[752]), .Z(n367) );
  XNOR U772 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U773 ( .A(in[432]), .B(n369), .Z(n1612) );
  XOR U774 ( .A(in[1521]), .B(in[561]), .Z(n371) );
  XNOR U775 ( .A(in[881]), .B(in[241]), .Z(n370) );
  XNOR U776 ( .A(n371), .B(n370), .Z(n372) );
  XNOR U777 ( .A(in[1201]), .B(n372), .Z(n1554) );
  XOR U778 ( .A(n1612), .B(n1554), .Z(n1471) );
  XOR U779 ( .A(in[177]), .B(n1471), .Z(n1525) );
  XOR U780 ( .A(in[1426]), .B(in[466]), .Z(n374) );
  XNOR U781 ( .A(in[786]), .B(in[146]), .Z(n373) );
  XNOR U782 ( .A(n374), .B(n373), .Z(n375) );
  XNOR U783 ( .A(in[1106]), .B(n375), .Z(n721) );
  XOR U784 ( .A(in[17]), .B(in[657]), .Z(n377) );
  XNOR U785 ( .A(in[977]), .B(in[337]), .Z(n376) );
  XNOR U786 ( .A(n377), .B(n376), .Z(n378) );
  XOR U787 ( .A(in[1297]), .B(n378), .Z(n1440) );
  XNOR U788 ( .A(n4482), .B(in[1362]), .Z(n1932) );
  XOR U789 ( .A(in[1370]), .B(in[730]), .Z(n380) );
  XNOR U790 ( .A(in[90]), .B(in[410]), .Z(n379) );
  XNOR U791 ( .A(n380), .B(n379), .Z(n381) );
  XNOR U792 ( .A(in[1050]), .B(n381), .Z(n1090) );
  XOR U793 ( .A(in[1561]), .B(in[601]), .Z(n383) );
  XNOR U794 ( .A(in[921]), .B(in[281]), .Z(n382) );
  XNOR U795 ( .A(n383), .B(n382), .Z(n384) );
  XNOR U796 ( .A(in[1241]), .B(n384), .Z(n823) );
  XOR U797 ( .A(n1090), .B(n823), .Z(n4256) );
  XOR U798 ( .A(in[986]), .B(n4256), .Z(n1929) );
  NANDN U799 ( .A(n1932), .B(n1929), .Z(n385) );
  XNOR U800 ( .A(n1525), .B(n385), .Z(out[1006]) );
  XOR U801 ( .A(in[1393]), .B(in[113]), .Z(n387) );
  XNOR U802 ( .A(in[1073]), .B(in[753]), .Z(n386) );
  XNOR U803 ( .A(n387), .B(n386), .Z(n388) );
  XNOR U804 ( .A(in[433]), .B(n388), .Z(n1616) );
  XOR U805 ( .A(in[1522]), .B(in[562]), .Z(n390) );
  XNOR U806 ( .A(in[882]), .B(in[242]), .Z(n389) );
  XNOR U807 ( .A(n390), .B(n389), .Z(n391) );
  XNOR U808 ( .A(in[1202]), .B(n391), .Z(n1558) );
  XOR U809 ( .A(n1616), .B(n1558), .Z(n1505) );
  XOR U810 ( .A(in[178]), .B(n1505), .Z(n1529) );
  XOR U811 ( .A(in[978]), .B(in[18]), .Z(n393) );
  XNOR U812 ( .A(in[1298]), .B(in[338]), .Z(n392) );
  XNOR U813 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U814 ( .A(in[658]), .B(n394), .Z(n1442) );
  XOR U815 ( .A(in[147]), .B(in[1427]), .Z(n396) );
  XNOR U816 ( .A(in[1107]), .B(in[787]), .Z(n395) );
  XNOR U817 ( .A(n396), .B(n395), .Z(n397) );
  XOR U818 ( .A(in[467]), .B(n397), .Z(n736) );
  XNOR U819 ( .A(in[1363]), .B(n4485), .Z(n1936) );
  XOR U820 ( .A(in[1371]), .B(in[731]), .Z(n399) );
  XNOR U821 ( .A(in[91]), .B(in[411]), .Z(n398) );
  XNOR U822 ( .A(n399), .B(n398), .Z(n400) );
  XNOR U823 ( .A(in[1051]), .B(n400), .Z(n1103) );
  XOR U824 ( .A(in[1562]), .B(in[602]), .Z(n402) );
  XNOR U825 ( .A(in[922]), .B(in[282]), .Z(n401) );
  XNOR U826 ( .A(n402), .B(n401), .Z(n403) );
  XNOR U827 ( .A(in[1242]), .B(n403), .Z(n838) );
  XOR U828 ( .A(n1103), .B(n838), .Z(n4257) );
  XOR U829 ( .A(in[987]), .B(n4257), .Z(n1933) );
  NANDN U830 ( .A(n1936), .B(n1933), .Z(n404) );
  XNOR U831 ( .A(n1529), .B(n404), .Z(out[1007]) );
  XOR U832 ( .A(in[1394]), .B(in[114]), .Z(n406) );
  XNOR U833 ( .A(in[1074]), .B(in[754]), .Z(n405) );
  XNOR U834 ( .A(n406), .B(n405), .Z(n407) );
  XNOR U835 ( .A(in[434]), .B(n407), .Z(n1620) );
  XOR U836 ( .A(in[1523]), .B(in[563]), .Z(n409) );
  XNOR U837 ( .A(in[883]), .B(in[243]), .Z(n408) );
  XNOR U838 ( .A(n409), .B(n408), .Z(n410) );
  XNOR U839 ( .A(in[1203]), .B(n410), .Z(n1562) );
  XOR U840 ( .A(n1620), .B(n1562), .Z(n1547) );
  XOR U841 ( .A(in[179]), .B(n1547), .Z(n1533) );
  XOR U842 ( .A(in[148]), .B(in[1428]), .Z(n412) );
  XNOR U843 ( .A(in[1108]), .B(in[788]), .Z(n411) );
  XNOR U844 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U845 ( .A(in[468]), .B(n413), .Z(n751) );
  XOR U846 ( .A(in[979]), .B(in[19]), .Z(n415) );
  XNOR U847 ( .A(in[1299]), .B(in[339]), .Z(n414) );
  XNOR U848 ( .A(n415), .B(n414), .Z(n416) );
  XOR U849 ( .A(in[659]), .B(n416), .Z(n1446) );
  XNOR U850 ( .A(in[1364]), .B(n4488), .Z(n1940) );
  XOR U851 ( .A(in[1372]), .B(in[732]), .Z(n418) );
  XNOR U852 ( .A(in[92]), .B(in[412]), .Z(n417) );
  XNOR U853 ( .A(n418), .B(n417), .Z(n419) );
  XNOR U854 ( .A(in[1052]), .B(n419), .Z(n1123) );
  XOR U855 ( .A(in[1563]), .B(in[603]), .Z(n421) );
  XNOR U856 ( .A(in[923]), .B(in[283]), .Z(n420) );
  XNOR U857 ( .A(n421), .B(n420), .Z(n422) );
  XNOR U858 ( .A(in[1243]), .B(n422), .Z(n853) );
  XOR U859 ( .A(n1123), .B(n853), .Z(n4260) );
  XOR U860 ( .A(in[988]), .B(n4260), .Z(n1937) );
  NANDN U861 ( .A(n1940), .B(n1937), .Z(n423) );
  XNOR U862 ( .A(n1533), .B(n423), .Z(out[1008]) );
  XOR U863 ( .A(in[1395]), .B(in[115]), .Z(n425) );
  XNOR U864 ( .A(in[1075]), .B(in[755]), .Z(n424) );
  XNOR U865 ( .A(n425), .B(n424), .Z(n426) );
  XNOR U866 ( .A(in[435]), .B(n426), .Z(n1624) );
  XOR U867 ( .A(in[1524]), .B(in[564]), .Z(n428) );
  XNOR U868 ( .A(in[884]), .B(in[244]), .Z(n427) );
  XNOR U869 ( .A(n428), .B(n427), .Z(n429) );
  XNOR U870 ( .A(in[1204]), .B(n429), .Z(n1566) );
  XOR U871 ( .A(n1624), .B(n1566), .Z(n1589) );
  XOR U872 ( .A(in[180]), .B(n1589), .Z(n1537) );
  XOR U873 ( .A(in[149]), .B(in[1429]), .Z(n431) );
  XNOR U874 ( .A(in[1109]), .B(in[789]), .Z(n430) );
  XNOR U875 ( .A(n431), .B(n430), .Z(n432) );
  XNOR U876 ( .A(in[469]), .B(n432), .Z(n766) );
  XOR U877 ( .A(in[340]), .B(in[660]), .Z(n434) );
  XNOR U878 ( .A(in[20]), .B(in[1300]), .Z(n433) );
  XNOR U879 ( .A(n434), .B(n433), .Z(n435) );
  XOR U880 ( .A(in[980]), .B(n435), .Z(n1448) );
  XNOR U881 ( .A(in[1365]), .B(n4491), .Z(n1944) );
  XOR U882 ( .A(in[1373]), .B(in[733]), .Z(n437) );
  XNOR U883 ( .A(in[93]), .B(in[413]), .Z(n436) );
  XNOR U884 ( .A(n437), .B(n436), .Z(n438) );
  XNOR U885 ( .A(in[1053]), .B(n438), .Z(n1136) );
  XOR U886 ( .A(in[1564]), .B(in[604]), .Z(n440) );
  XNOR U887 ( .A(in[924]), .B(in[284]), .Z(n439) );
  XNOR U888 ( .A(n440), .B(n439), .Z(n441) );
  XNOR U889 ( .A(in[1244]), .B(n441), .Z(n868) );
  XOR U890 ( .A(n1136), .B(n868), .Z(n4261) );
  XOR U891 ( .A(in[989]), .B(n4261), .Z(n1941) );
  NANDN U892 ( .A(n1944), .B(n1941), .Z(n442) );
  XNOR U893 ( .A(n1537), .B(n442), .Z(out[1009]) );
  XOR U894 ( .A(in[1339]), .B(in[59]), .Z(n444) );
  XNOR U895 ( .A(in[699]), .B(in[379]), .Z(n443) );
  XNOR U896 ( .A(n444), .B(n443), .Z(n445) );
  XNOR U897 ( .A(in[1019]), .B(n445), .Z(n1094) );
  XOR U898 ( .A(in[1530]), .B(in[570]), .Z(n447) );
  XNOR U899 ( .A(in[1210]), .B(in[250]), .Z(n446) );
  XNOR U900 ( .A(n447), .B(n446), .Z(n448) );
  XNOR U901 ( .A(in[890]), .B(n448), .Z(n560) );
  XOR U902 ( .A(n1094), .B(n560), .Z(n3953) );
  XOR U903 ( .A(in[635]), .B(n3953), .Z(n2704) );
  IV U904 ( .A(n2704), .Z(n2790) );
  XOR U905 ( .A(in[161]), .B(in[1441]), .Z(n450) );
  XNOR U906 ( .A(in[801]), .B(in[1121]), .Z(n449) );
  XNOR U907 ( .A(n450), .B(n449), .Z(n451) );
  XNOR U908 ( .A(in[481]), .B(n451), .Z(n687) );
  XOR U909 ( .A(in[1570]), .B(in[610]), .Z(n453) );
  XNOR U910 ( .A(in[930]), .B(in[290]), .Z(n452) );
  XNOR U911 ( .A(n453), .B(n452), .Z(n454) );
  XOR U912 ( .A(in[1250]), .B(n454), .Z(n570) );
  XOR U913 ( .A(in[226]), .B(n4049), .Z(n3115) );
  XOR U914 ( .A(in[1510]), .B(in[550]), .Z(n456) );
  XNOR U915 ( .A(in[870]), .B(in[230]), .Z(n455) );
  XNOR U916 ( .A(n456), .B(n455), .Z(n457) );
  XNOR U917 ( .A(in[1190]), .B(n457), .Z(n1508) );
  XOR U918 ( .A(in[1061]), .B(in[421]), .Z(n459) );
  XNOR U919 ( .A(in[741]), .B(in[1381]), .Z(n458) );
  XNOR U920 ( .A(n459), .B(n458), .Z(n460) );
  XNOR U921 ( .A(in[101]), .B(n460), .Z(n606) );
  XNOR U922 ( .A(n1508), .B(n606), .Z(n4089) );
  IV U923 ( .A(n4089), .Z(n1249) );
  XOR U924 ( .A(in[1446]), .B(n1249), .Z(n3112) );
  NANDN U925 ( .A(n3115), .B(n3112), .Z(n461) );
  XOR U926 ( .A(n2790), .B(n461), .Z(out[100]) );
  XOR U927 ( .A(in[1396]), .B(in[116]), .Z(n463) );
  XNOR U928 ( .A(in[1076]), .B(in[756]), .Z(n462) );
  XNOR U929 ( .A(n463), .B(n462), .Z(n464) );
  XNOR U930 ( .A(in[436]), .B(n464), .Z(n1629) );
  XOR U931 ( .A(in[1525]), .B(in[565]), .Z(n466) );
  XNOR U932 ( .A(in[885]), .B(in[245]), .Z(n465) );
  XNOR U933 ( .A(n466), .B(n465), .Z(n467) );
  XNOR U934 ( .A(in[1205]), .B(n467), .Z(n1570) );
  XOR U935 ( .A(n1629), .B(n1570), .Z(n4153) );
  XOR U936 ( .A(in[181]), .B(n4153), .Z(n1541) );
  XOR U937 ( .A(in[341]), .B(in[661]), .Z(n469) );
  XNOR U938 ( .A(in[21]), .B(in[1301]), .Z(n468) );
  XNOR U939 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U940 ( .A(in[981]), .B(n470), .Z(n1450) );
  XOR U941 ( .A(in[150]), .B(in[1430]), .Z(n472) );
  XNOR U942 ( .A(in[1110]), .B(in[790]), .Z(n471) );
  XNOR U943 ( .A(n472), .B(n471), .Z(n473) );
  XOR U944 ( .A(in[470]), .B(n473), .Z(n781) );
  XNOR U945 ( .A(in[1366]), .B(n4494), .Z(n1948) );
  XOR U946 ( .A(in[1374]), .B(in[734]), .Z(n475) );
  XNOR U947 ( .A(in[94]), .B(in[414]), .Z(n474) );
  XNOR U948 ( .A(n475), .B(n474), .Z(n476) );
  XNOR U949 ( .A(in[1054]), .B(n476), .Z(n1149) );
  XOR U950 ( .A(in[1565]), .B(in[605]), .Z(n478) );
  XNOR U951 ( .A(in[925]), .B(in[285]), .Z(n477) );
  XNOR U952 ( .A(n478), .B(n477), .Z(n479) );
  XNOR U953 ( .A(in[1245]), .B(n479), .Z(n883) );
  XOR U954 ( .A(n1149), .B(n883), .Z(n4262) );
  XOR U955 ( .A(in[990]), .B(n4262), .Z(n1945) );
  NANDN U956 ( .A(n1948), .B(n1945), .Z(n480) );
  XNOR U957 ( .A(n1541), .B(n480), .Z(out[1010]) );
  XOR U958 ( .A(in[1526]), .B(in[566]), .Z(n482) );
  XNOR U959 ( .A(in[886]), .B(in[246]), .Z(n481) );
  XNOR U960 ( .A(n482), .B(n481), .Z(n483) );
  XNOR U961 ( .A(in[1206]), .B(n483), .Z(n1574) );
  XOR U962 ( .A(in[1397]), .B(in[117]), .Z(n485) );
  XNOR U963 ( .A(in[1077]), .B(in[757]), .Z(n484) );
  XNOR U964 ( .A(n485), .B(n484), .Z(n486) );
  XNOR U965 ( .A(in[437]), .B(n486), .Z(n1633) );
  XOR U966 ( .A(n1574), .B(n1633), .Z(n4163) );
  XOR U967 ( .A(in[182]), .B(n4163), .Z(n1545) );
  XOR U968 ( .A(in[342]), .B(in[662]), .Z(n488) );
  XNOR U969 ( .A(in[22]), .B(in[1302]), .Z(n487) );
  XNOR U970 ( .A(n488), .B(n487), .Z(n489) );
  XNOR U971 ( .A(in[982]), .B(n489), .Z(n1452) );
  XOR U972 ( .A(in[151]), .B(in[1431]), .Z(n491) );
  XNOR U973 ( .A(in[1111]), .B(in[791]), .Z(n490) );
  XNOR U974 ( .A(n491), .B(n490), .Z(n492) );
  XOR U975 ( .A(in[471]), .B(n492), .Z(n796) );
  XNOR U976 ( .A(in[1367]), .B(n4497), .Z(n1952) );
  XOR U977 ( .A(in[1375]), .B(in[735]), .Z(n494) );
  XNOR U978 ( .A(in[95]), .B(in[415]), .Z(n493) );
  XNOR U979 ( .A(n494), .B(n493), .Z(n495) );
  XNOR U980 ( .A(in[1055]), .B(n495), .Z(n1162) );
  XOR U981 ( .A(in[1566]), .B(in[606]), .Z(n497) );
  XNOR U982 ( .A(in[926]), .B(in[286]), .Z(n496) );
  XNOR U983 ( .A(n497), .B(n496), .Z(n498) );
  XNOR U984 ( .A(in[1246]), .B(n498), .Z(n898) );
  XOR U985 ( .A(n1162), .B(n898), .Z(n4263) );
  XOR U986 ( .A(in[991]), .B(n4263), .Z(n1949) );
  NANDN U987 ( .A(n1952), .B(n1949), .Z(n499) );
  XNOR U988 ( .A(n1545), .B(n499), .Z(out[1011]) );
  XOR U989 ( .A(in[1527]), .B(in[567]), .Z(n501) );
  XNOR U990 ( .A(in[887]), .B(in[247]), .Z(n500) );
  XNOR U991 ( .A(n501), .B(n500), .Z(n502) );
  XNOR U992 ( .A(in[1207]), .B(n502), .Z(n1578) );
  XOR U993 ( .A(in[1398]), .B(in[118]), .Z(n504) );
  XNOR U994 ( .A(in[1078]), .B(in[758]), .Z(n503) );
  XNOR U995 ( .A(n504), .B(n503), .Z(n505) );
  XNOR U996 ( .A(in[438]), .B(n505), .Z(n1637) );
  XOR U997 ( .A(n1578), .B(n1637), .Z(n4167) );
  XOR U998 ( .A(in[183]), .B(n4167), .Z(n1551) );
  XOR U999 ( .A(in[343]), .B(in[663]), .Z(n507) );
  XNOR U1000 ( .A(in[23]), .B(in[1303]), .Z(n506) );
  XNOR U1001 ( .A(n507), .B(n506), .Z(n508) );
  XNOR U1002 ( .A(in[983]), .B(n508), .Z(n1454) );
  XOR U1003 ( .A(in[152]), .B(in[1432]), .Z(n510) );
  XNOR U1004 ( .A(in[1112]), .B(in[792]), .Z(n509) );
  XNOR U1005 ( .A(n510), .B(n509), .Z(n511) );
  XOR U1006 ( .A(in[472]), .B(n511), .Z(n822) );
  XNOR U1007 ( .A(in[1368]), .B(n4500), .Z(n1956) );
  XOR U1008 ( .A(in[1376]), .B(in[736]), .Z(n513) );
  XNOR U1009 ( .A(in[96]), .B(in[416]), .Z(n512) );
  XNOR U1010 ( .A(n513), .B(n512), .Z(n514) );
  XNOR U1011 ( .A(in[1056]), .B(n514), .Z(n1177) );
  XOR U1012 ( .A(in[1567]), .B(in[607]), .Z(n516) );
  XNOR U1013 ( .A(in[927]), .B(in[287]), .Z(n515) );
  XNOR U1014 ( .A(n516), .B(n515), .Z(n517) );
  XNOR U1015 ( .A(in[1247]), .B(n517), .Z(n913) );
  XOR U1016 ( .A(n1177), .B(n913), .Z(n4266) );
  XOR U1017 ( .A(in[992]), .B(n4266), .Z(n1953) );
  NANDN U1018 ( .A(n1956), .B(n1953), .Z(n518) );
  XNOR U1019 ( .A(n1551), .B(n518), .Z(out[1012]) );
  XOR U1020 ( .A(in[1528]), .B(in[568]), .Z(n520) );
  XNOR U1021 ( .A(in[888]), .B(in[248]), .Z(n519) );
  XNOR U1022 ( .A(n520), .B(n519), .Z(n521) );
  XNOR U1023 ( .A(in[1208]), .B(n521), .Z(n1582) );
  XOR U1024 ( .A(in[1399]), .B(in[119]), .Z(n523) );
  XNOR U1025 ( .A(in[1079]), .B(in[759]), .Z(n522) );
  XNOR U1026 ( .A(n523), .B(n522), .Z(n524) );
  XNOR U1027 ( .A(in[439]), .B(n524), .Z(n1641) );
  XOR U1028 ( .A(n1582), .B(n1641), .Z(n4171) );
  XOR U1029 ( .A(in[184]), .B(n4171), .Z(n1555) );
  XOR U1030 ( .A(in[153]), .B(in[1433]), .Z(n526) );
  XNOR U1031 ( .A(in[1113]), .B(in[793]), .Z(n525) );
  XNOR U1032 ( .A(n526), .B(n525), .Z(n527) );
  XNOR U1033 ( .A(in[473]), .B(n527), .Z(n837) );
  XOR U1034 ( .A(in[344]), .B(in[664]), .Z(n529) );
  XNOR U1035 ( .A(in[24]), .B(in[1304]), .Z(n528) );
  XNOR U1036 ( .A(n529), .B(n528), .Z(n530) );
  XOR U1037 ( .A(in[984]), .B(n530), .Z(n1456) );
  XNOR U1038 ( .A(in[1369]), .B(n4503), .Z(n1960) );
  XOR U1039 ( .A(in[1377]), .B(in[737]), .Z(n532) );
  XNOR U1040 ( .A(in[97]), .B(in[417]), .Z(n531) );
  XNOR U1041 ( .A(n532), .B(n531), .Z(n533) );
  XNOR U1042 ( .A(in[1057]), .B(n533), .Z(n1192) );
  XOR U1043 ( .A(in[1568]), .B(in[608]), .Z(n535) );
  XNOR U1044 ( .A(in[928]), .B(in[288]), .Z(n534) );
  XNOR U1045 ( .A(n535), .B(n534), .Z(n536) );
  XNOR U1046 ( .A(in[1248]), .B(n536), .Z(n928) );
  XOR U1047 ( .A(n1192), .B(n928), .Z(n4269) );
  XOR U1048 ( .A(in[993]), .B(n4269), .Z(n1957) );
  NANDN U1049 ( .A(n1960), .B(n1957), .Z(n537) );
  XNOR U1050 ( .A(n1555), .B(n537), .Z(out[1013]) );
  XOR U1051 ( .A(in[1529]), .B(in[569]), .Z(n539) );
  XNOR U1052 ( .A(in[889]), .B(in[249]), .Z(n538) );
  XNOR U1053 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U1054 ( .A(in[1209]), .B(n540), .Z(n1586) );
  XOR U1055 ( .A(in[1400]), .B(in[120]), .Z(n542) );
  XNOR U1056 ( .A(in[1080]), .B(in[760]), .Z(n541) );
  XNOR U1057 ( .A(n542), .B(n541), .Z(n543) );
  XNOR U1058 ( .A(in[440]), .B(n543), .Z(n1645) );
  XOR U1059 ( .A(n1586), .B(n1645), .Z(n4175) );
  XOR U1060 ( .A(in[185]), .B(n4175), .Z(n1559) );
  XOR U1061 ( .A(in[154]), .B(in[1434]), .Z(n545) );
  XNOR U1062 ( .A(in[1114]), .B(in[794]), .Z(n544) );
  XNOR U1063 ( .A(n545), .B(n544), .Z(n546) );
  XNOR U1064 ( .A(in[474]), .B(n546), .Z(n852) );
  XOR U1065 ( .A(in[345]), .B(in[665]), .Z(n548) );
  XNOR U1066 ( .A(in[25]), .B(in[1305]), .Z(n547) );
  XNOR U1067 ( .A(n548), .B(n547), .Z(n549) );
  XOR U1068 ( .A(in[985]), .B(n549), .Z(n1460) );
  XNOR U1069 ( .A(in[1370]), .B(n4506), .Z(n1966) );
  XOR U1070 ( .A(in[1569]), .B(in[609]), .Z(n551) );
  XNOR U1071 ( .A(in[929]), .B(in[289]), .Z(n550) );
  XNOR U1072 ( .A(n551), .B(n550), .Z(n552) );
  XNOR U1073 ( .A(in[1249]), .B(n552), .Z(n943) );
  XOR U1074 ( .A(in[1378]), .B(in[738]), .Z(n554) );
  XNOR U1075 ( .A(in[98]), .B(in[418]), .Z(n553) );
  XNOR U1076 ( .A(n554), .B(n553), .Z(n555) );
  XNOR U1077 ( .A(in[1058]), .B(n555), .Z(n1207) );
  XOR U1078 ( .A(n943), .B(n1207), .Z(n4272) );
  XOR U1079 ( .A(in[994]), .B(n4272), .Z(n1963) );
  NANDN U1080 ( .A(n1966), .B(n1963), .Z(n556) );
  XNOR U1081 ( .A(n1559), .B(n556), .Z(out[1014]) );
  XOR U1082 ( .A(in[1401]), .B(in[121]), .Z(n558) );
  XNOR U1083 ( .A(in[1081]), .B(in[761]), .Z(n557) );
  XNOR U1084 ( .A(n558), .B(n557), .Z(n559) );
  XNOR U1085 ( .A(in[441]), .B(n559), .Z(n1649) );
  XOR U1086 ( .A(n560), .B(n1649), .Z(n1796) );
  XOR U1087 ( .A(in[186]), .B(n1796), .Z(n1563) );
  XOR U1088 ( .A(in[155]), .B(in[1435]), .Z(n562) );
  XNOR U1089 ( .A(in[1115]), .B(in[795]), .Z(n561) );
  XNOR U1090 ( .A(n562), .B(n561), .Z(n563) );
  XNOR U1091 ( .A(in[475]), .B(n563), .Z(n867) );
  XOR U1092 ( .A(in[346]), .B(in[666]), .Z(n565) );
  XNOR U1093 ( .A(in[26]), .B(in[1306]), .Z(n564) );
  XNOR U1094 ( .A(n565), .B(n564), .Z(n566) );
  XOR U1095 ( .A(in[986]), .B(n566), .Z(n1462) );
  IV U1096 ( .A(n4513), .Z(n2740) );
  XOR U1097 ( .A(in[1371]), .B(n2740), .Z(n1365) );
  IV U1098 ( .A(n1365), .Z(n1970) );
  XOR U1099 ( .A(in[1379]), .B(in[739]), .Z(n568) );
  XNOR U1100 ( .A(in[99]), .B(in[419]), .Z(n567) );
  XNOR U1101 ( .A(n568), .B(n567), .Z(n569) );
  XOR U1102 ( .A(in[1059]), .B(n569), .Z(n1222) );
  XNOR U1103 ( .A(n570), .B(n1222), .Z(n4275) );
  XNOR U1104 ( .A(in[995]), .B(n4275), .Z(n1967) );
  NANDN U1105 ( .A(n1970), .B(n1967), .Z(n571) );
  XNOR U1106 ( .A(n1563), .B(n571), .Z(out[1015]) );
  XOR U1107 ( .A(in[1402]), .B(in[122]), .Z(n573) );
  XNOR U1108 ( .A(in[1082]), .B(in[762]), .Z(n572) );
  XNOR U1109 ( .A(n573), .B(n572), .Z(n574) );
  XNOR U1110 ( .A(in[442]), .B(n574), .Z(n1653) );
  XOR U1111 ( .A(in[1531]), .B(in[571]), .Z(n576) );
  XNOR U1112 ( .A(in[1211]), .B(in[251]), .Z(n575) );
  XNOR U1113 ( .A(n576), .B(n575), .Z(n577) );
  XNOR U1114 ( .A(in[891]), .B(n577), .Z(n649) );
  XOR U1115 ( .A(n1653), .B(n649), .Z(n1822) );
  XOR U1116 ( .A(in[187]), .B(n1822), .Z(n1567) );
  XOR U1117 ( .A(in[156]), .B(in[1436]), .Z(n579) );
  XNOR U1118 ( .A(in[1116]), .B(in[796]), .Z(n578) );
  XNOR U1119 ( .A(n579), .B(n578), .Z(n580) );
  XNOR U1120 ( .A(in[476]), .B(n580), .Z(n882) );
  XOR U1121 ( .A(in[347]), .B(in[667]), .Z(n582) );
  XNOR U1122 ( .A(in[27]), .B(in[1307]), .Z(n581) );
  XNOR U1123 ( .A(n582), .B(n581), .Z(n583) );
  XOR U1124 ( .A(in[987]), .B(n583), .Z(n1464) );
  IV U1125 ( .A(n4516), .Z(n2757) );
  XOR U1126 ( .A(in[1372]), .B(n2757), .Z(n1375) );
  IV U1127 ( .A(n1375), .Z(n1974) );
  XOR U1128 ( .A(in[1060]), .B(in[420]), .Z(n585) );
  XNOR U1129 ( .A(in[740]), .B(in[1380]), .Z(n584) );
  XNOR U1130 ( .A(n585), .B(n584), .Z(n586) );
  XNOR U1131 ( .A(in[100]), .B(n586), .Z(n1237) );
  XOR U1132 ( .A(in[1571]), .B(in[611]), .Z(n588) );
  XNOR U1133 ( .A(in[931]), .B(in[291]), .Z(n587) );
  XNOR U1134 ( .A(n588), .B(n587), .Z(n589) );
  XNOR U1135 ( .A(in[1251]), .B(n589), .Z(n653) );
  XOR U1136 ( .A(n1237), .B(n653), .Z(n4278) );
  XOR U1137 ( .A(in[996]), .B(n4278), .Z(n1971) );
  NANDN U1138 ( .A(n1974), .B(n1971), .Z(n590) );
  XNOR U1139 ( .A(n1567), .B(n590), .Z(out[1016]) );
  XOR U1140 ( .A(in[1403]), .B(in[123]), .Z(n592) );
  XNOR U1141 ( .A(in[1083]), .B(in[763]), .Z(n591) );
  XNOR U1142 ( .A(n592), .B(n591), .Z(n593) );
  XNOR U1143 ( .A(in[443]), .B(n593), .Z(n1657) );
  XOR U1144 ( .A(in[1532]), .B(in[572]), .Z(n595) );
  XNOR U1145 ( .A(in[1212]), .B(in[252]), .Z(n594) );
  XNOR U1146 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U1147 ( .A(in[892]), .B(n596), .Z(n814) );
  XOR U1148 ( .A(n1657), .B(n814), .Z(n1845) );
  XOR U1149 ( .A(in[188]), .B(n1845), .Z(n1571) );
  XOR U1150 ( .A(in[157]), .B(in[1437]), .Z(n598) );
  XNOR U1151 ( .A(in[1117]), .B(in[797]), .Z(n597) );
  XNOR U1152 ( .A(n598), .B(n597), .Z(n599) );
  XNOR U1153 ( .A(in[477]), .B(n599), .Z(n897) );
  XOR U1154 ( .A(in[348]), .B(in[668]), .Z(n601) );
  XNOR U1155 ( .A(in[28]), .B(in[1308]), .Z(n600) );
  XNOR U1156 ( .A(n601), .B(n600), .Z(n602) );
  XOR U1157 ( .A(in[988]), .B(n602), .Z(n1468) );
  IV U1158 ( .A(n4519), .Z(n2774) );
  XOR U1159 ( .A(in[1373]), .B(n2774), .Z(n1381) );
  IV U1160 ( .A(n1381), .Z(n1978) );
  XOR U1161 ( .A(in[1572]), .B(in[612]), .Z(n604) );
  XNOR U1162 ( .A(in[932]), .B(in[292]), .Z(n603) );
  XNOR U1163 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U1164 ( .A(in[1252]), .B(n605), .Z(n816) );
  XOR U1165 ( .A(n606), .B(n816), .Z(n4280) );
  XOR U1166 ( .A(in[997]), .B(n4280), .Z(n1975) );
  NANDN U1167 ( .A(n1978), .B(n1975), .Z(n607) );
  XNOR U1168 ( .A(n1571), .B(n607), .Z(out[1017]) );
  XOR U1169 ( .A(in[1404]), .B(in[124]), .Z(n609) );
  XNOR U1170 ( .A(in[1084]), .B(in[764]), .Z(n608) );
  XNOR U1171 ( .A(n609), .B(n608), .Z(n610) );
  XNOR U1172 ( .A(in[444]), .B(n610), .Z(n1661) );
  XOR U1173 ( .A(in[1533]), .B(in[573]), .Z(n612) );
  XNOR U1174 ( .A(in[1213]), .B(in[253]), .Z(n611) );
  XNOR U1175 ( .A(n612), .B(n611), .Z(n613) );
  XNOR U1176 ( .A(in[893]), .B(n613), .Z(n973) );
  XOR U1177 ( .A(n1661), .B(n973), .Z(n1867) );
  XOR U1178 ( .A(in[189]), .B(n1867), .Z(n1575) );
  XOR U1179 ( .A(in[158]), .B(in[1438]), .Z(n615) );
  XNOR U1180 ( .A(in[1118]), .B(in[798]), .Z(n614) );
  XNOR U1181 ( .A(n615), .B(n614), .Z(n616) );
  XNOR U1182 ( .A(in[478]), .B(n616), .Z(n912) );
  XOR U1183 ( .A(in[349]), .B(in[669]), .Z(n618) );
  XNOR U1184 ( .A(in[29]), .B(in[1309]), .Z(n617) );
  XNOR U1185 ( .A(n618), .B(n617), .Z(n619) );
  XOR U1186 ( .A(in[989]), .B(n619), .Z(n1474) );
  XNOR U1187 ( .A(in[1374]), .B(n4522), .Z(n1982) );
  XOR U1188 ( .A(in[1062]), .B(in[422]), .Z(n621) );
  XNOR U1189 ( .A(in[742]), .B(in[1382]), .Z(n620) );
  XNOR U1190 ( .A(n621), .B(n620), .Z(n622) );
  XNOR U1191 ( .A(in[102]), .B(n622), .Z(n657) );
  XOR U1192 ( .A(in[1573]), .B(in[613]), .Z(n624) );
  XNOR U1193 ( .A(in[933]), .B(in[293]), .Z(n623) );
  XNOR U1194 ( .A(n624), .B(n623), .Z(n625) );
  XNOR U1195 ( .A(in[1253]), .B(n625), .Z(n975) );
  XOR U1196 ( .A(n657), .B(n975), .Z(n4286) );
  XOR U1197 ( .A(in[998]), .B(n4286), .Z(n1979) );
  NANDN U1198 ( .A(n1982), .B(n1979), .Z(n626) );
  XNOR U1199 ( .A(n1575), .B(n626), .Z(out[1018]) );
  XOR U1200 ( .A(in[1405]), .B(in[125]), .Z(n628) );
  XNOR U1201 ( .A(in[1085]), .B(in[765]), .Z(n627) );
  XNOR U1202 ( .A(n628), .B(n627), .Z(n629) );
  XNOR U1203 ( .A(in[445]), .B(n629), .Z(n1665) );
  XOR U1204 ( .A(in[1534]), .B(in[894]), .Z(n631) );
  XNOR U1205 ( .A(in[574]), .B(in[1214]), .Z(n630) );
  XNOR U1206 ( .A(n631), .B(n630), .Z(n632) );
  XNOR U1207 ( .A(in[254]), .B(n632), .Z(n1110) );
  XOR U1208 ( .A(n1665), .B(n1110), .Z(n1889) );
  XOR U1209 ( .A(in[190]), .B(n1889), .Z(n1579) );
  XOR U1210 ( .A(in[1439]), .B(in[479]), .Z(n634) );
  XNOR U1211 ( .A(in[799]), .B(in[159]), .Z(n633) );
  XNOR U1212 ( .A(n634), .B(n633), .Z(n635) );
  XNOR U1213 ( .A(in[1119]), .B(n635), .Z(n927) );
  XOR U1214 ( .A(in[350]), .B(in[670]), .Z(n637) );
  XNOR U1215 ( .A(in[30]), .B(in[1310]), .Z(n636) );
  XNOR U1216 ( .A(n637), .B(n636), .Z(n638) );
  XOR U1217 ( .A(in[990]), .B(n638), .Z(n1478) );
  XNOR U1218 ( .A(in[1375]), .B(n4526), .Z(n1986) );
  XOR U1219 ( .A(in[1063]), .B(in[423]), .Z(n640) );
  XNOR U1220 ( .A(in[743]), .B(in[1383]), .Z(n639) );
  XNOR U1221 ( .A(n640), .B(n639), .Z(n641) );
  XNOR U1222 ( .A(in[103]), .B(n641), .Z(n820) );
  XOR U1223 ( .A(in[1574]), .B(in[614]), .Z(n643) );
  XNOR U1224 ( .A(in[934]), .B(in[294]), .Z(n642) );
  XNOR U1225 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U1226 ( .A(in[1254]), .B(n644), .Z(n1019) );
  XOR U1227 ( .A(n820), .B(n1019), .Z(n4288) );
  XOR U1228 ( .A(in[999]), .B(n4288), .Z(n1983) );
  NANDN U1229 ( .A(n1986), .B(n1983), .Z(n645) );
  XNOR U1230 ( .A(n1579), .B(n645), .Z(out[1019]) );
  XOR U1231 ( .A(in[1340]), .B(in[60]), .Z(n647) );
  XNOR U1232 ( .A(in[700]), .B(in[380]), .Z(n646) );
  XNOR U1233 ( .A(n647), .B(n646), .Z(n648) );
  XNOR U1234 ( .A(in[1020]), .B(n648), .Z(n1104) );
  XOR U1235 ( .A(n649), .B(n1104), .Z(n3957) );
  XOR U1236 ( .A(in[636]), .B(n3957), .Z(n2706) );
  IV U1237 ( .A(n2706), .Z(n2792) );
  XOR U1238 ( .A(in[162]), .B(in[1442]), .Z(n651) );
  XNOR U1239 ( .A(in[802]), .B(in[1122]), .Z(n650) );
  XNOR U1240 ( .A(n651), .B(n650), .Z(n652) );
  XOR U1241 ( .A(in[482]), .B(n652), .Z(n704) );
  XOR U1242 ( .A(n653), .B(n704), .Z(n3398) );
  IV U1243 ( .A(n3398), .Z(n4053) );
  XOR U1244 ( .A(in[227]), .B(n4053), .Z(n3137) );
  XOR U1245 ( .A(in[1511]), .B(in[551]), .Z(n655) );
  XNOR U1246 ( .A(in[871]), .B(in[231]), .Z(n654) );
  XNOR U1247 ( .A(n655), .B(n654), .Z(n656) );
  XNOR U1248 ( .A(in[1191]), .B(n656), .Z(n1512) );
  XNOR U1249 ( .A(n657), .B(n1512), .Z(n4093) );
  IV U1250 ( .A(n4093), .Z(n1264) );
  XOR U1251 ( .A(in[1447]), .B(n1264), .Z(n3134) );
  NANDN U1252 ( .A(n3137), .B(n3134), .Z(n658) );
  XOR U1253 ( .A(n2792), .B(n658), .Z(out[101]) );
  XOR U1254 ( .A(in[1406]), .B(in[126]), .Z(n660) );
  XNOR U1255 ( .A(in[1086]), .B(in[766]), .Z(n659) );
  XNOR U1256 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U1257 ( .A(in[446]), .B(n661), .Z(n1670) );
  XOR U1258 ( .A(in[1535]), .B(in[575]), .Z(n663) );
  XNOR U1259 ( .A(in[895]), .B(in[255]), .Z(n662) );
  XNOR U1260 ( .A(n663), .B(n662), .Z(n664) );
  XNOR U1261 ( .A(in[1215]), .B(n664), .Z(n1258) );
  XOR U1262 ( .A(n1670), .B(n1258), .Z(n1919) );
  XOR U1263 ( .A(in[191]), .B(n1919), .Z(n1583) );
  XOR U1264 ( .A(in[1440]), .B(in[480]), .Z(n666) );
  XNOR U1265 ( .A(in[800]), .B(in[160]), .Z(n665) );
  XNOR U1266 ( .A(n666), .B(n665), .Z(n667) );
  XNOR U1267 ( .A(in[1120]), .B(n667), .Z(n942) );
  XOR U1268 ( .A(in[351]), .B(in[671]), .Z(n669) );
  XNOR U1269 ( .A(in[31]), .B(in[1311]), .Z(n668) );
  XNOR U1270 ( .A(n669), .B(n668), .Z(n670) );
  XOR U1271 ( .A(in[991]), .B(n670), .Z(n1482) );
  XNOR U1272 ( .A(in[1376]), .B(n4530), .Z(n1990) );
  XOR U1273 ( .A(in[1064]), .B(in[424]), .Z(n672) );
  XNOR U1274 ( .A(in[744]), .B(in[1384]), .Z(n671) );
  XNOR U1275 ( .A(n672), .B(n671), .Z(n673) );
  XNOR U1276 ( .A(in[104]), .B(n673), .Z(n979) );
  XOR U1277 ( .A(in[1575]), .B(in[615]), .Z(n675) );
  XNOR U1278 ( .A(in[935]), .B(in[295]), .Z(n674) );
  XNOR U1279 ( .A(n675), .B(n674), .Z(n676) );
  XNOR U1280 ( .A(in[1255]), .B(n676), .Z(n1032) );
  XOR U1281 ( .A(n979), .B(n1032), .Z(n4290) );
  XOR U1282 ( .A(in[1000]), .B(n4290), .Z(n1987) );
  NANDN U1283 ( .A(n1990), .B(n1987), .Z(n677) );
  XNOR U1284 ( .A(n1583), .B(n677), .Z(out[1020]) );
  XOR U1285 ( .A(in[1407]), .B(in[127]), .Z(n679) );
  XNOR U1286 ( .A(in[1087]), .B(in[767]), .Z(n678) );
  XNOR U1287 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U1288 ( .A(in[447]), .B(n680), .Z(n1673) );
  XOR U1289 ( .A(in[1472]), .B(in[512]), .Z(n682) );
  XNOR U1290 ( .A(in[832]), .B(in[192]), .Z(n681) );
  XNOR U1291 ( .A(n682), .B(n681), .Z(n683) );
  XNOR U1292 ( .A(in[1152]), .B(n683), .Z(n1323) );
  XOR U1293 ( .A(n1673), .B(n1323), .Z(n1961) );
  XOR U1294 ( .A(in[128]), .B(n1961), .Z(n1587) );
  XOR U1295 ( .A(in[352]), .B(in[672]), .Z(n685) );
  XNOR U1296 ( .A(in[32]), .B(in[1312]), .Z(n684) );
  XNOR U1297 ( .A(n685), .B(n684), .Z(n686) );
  XOR U1298 ( .A(in[992]), .B(n686), .Z(n1484) );
  XNOR U1299 ( .A(in[1377]), .B(n4534), .Z(n1994) );
  XOR U1300 ( .A(in[1065]), .B(in[425]), .Z(n689) );
  XNOR U1301 ( .A(in[745]), .B(in[1385]), .Z(n688) );
  XNOR U1302 ( .A(n689), .B(n688), .Z(n690) );
  XNOR U1303 ( .A(in[105]), .B(n690), .Z(n1114) );
  XOR U1304 ( .A(in[1576]), .B(in[616]), .Z(n692) );
  XNOR U1305 ( .A(in[936]), .B(in[296]), .Z(n691) );
  XNOR U1306 ( .A(n692), .B(n691), .Z(n693) );
  XNOR U1307 ( .A(in[1256]), .B(n693), .Z(n1045) );
  XOR U1308 ( .A(n1114), .B(n1045), .Z(n4292) );
  XOR U1309 ( .A(in[1001]), .B(n4292), .Z(n1991) );
  NANDN U1310 ( .A(n1994), .B(n1991), .Z(n694) );
  XNOR U1311 ( .A(n1587), .B(n694), .Z(out[1021]) );
  XOR U1312 ( .A(in[1344]), .B(in[64]), .Z(n696) );
  XNOR U1313 ( .A(in[1024]), .B(in[384]), .Z(n695) );
  XNOR U1314 ( .A(n696), .B(n695), .Z(n697) );
  XNOR U1315 ( .A(in[704]), .B(n697), .Z(n1678) );
  XOR U1316 ( .A(in[1473]), .B(in[513]), .Z(n699) );
  XNOR U1317 ( .A(in[833]), .B(in[193]), .Z(n698) );
  XNOR U1318 ( .A(n699), .B(n698), .Z(n700) );
  XNOR U1319 ( .A(in[1153]), .B(n700), .Z(n1368) );
  XOR U1320 ( .A(n1678), .B(n1368), .Z(n2003) );
  XOR U1321 ( .A(in[129]), .B(n2003), .Z(n1591) );
  XOR U1322 ( .A(in[353]), .B(in[673]), .Z(n702) );
  XNOR U1323 ( .A(in[33]), .B(in[1313]), .Z(n701) );
  XNOR U1324 ( .A(n702), .B(n701), .Z(n703) );
  XNOR U1325 ( .A(in[993]), .B(n703), .Z(n1487) );
  XNOR U1326 ( .A(in[1378]), .B(n4538), .Z(n1998) );
  XOR U1327 ( .A(in[1577]), .B(in[617]), .Z(n706) );
  XNOR U1328 ( .A(in[937]), .B(in[297]), .Z(n705) );
  XNOR U1329 ( .A(n706), .B(n705), .Z(n707) );
  XNOR U1330 ( .A(in[1257]), .B(n707), .Z(n1058) );
  XOR U1331 ( .A(n708), .B(n1058), .Z(n4294) );
  XOR U1332 ( .A(in[1002]), .B(n4294), .Z(n1995) );
  NANDN U1333 ( .A(n1998), .B(n1995), .Z(n709) );
  XNOR U1334 ( .A(n1591), .B(n709), .Z(out[1022]) );
  IV U1335 ( .A(n3171), .Z(n3932) );
  XOR U1336 ( .A(n3932), .B(in[130]), .Z(n1593) );
  XOR U1337 ( .A(in[163]), .B(in[1443]), .Z(n711) );
  XNOR U1338 ( .A(in[803]), .B(in[1123]), .Z(n710) );
  XNOR U1339 ( .A(n711), .B(n710), .Z(n712) );
  XNOR U1340 ( .A(in[483]), .B(n712), .Z(n815) );
  XOR U1341 ( .A(in[354]), .B(in[674]), .Z(n714) );
  XNOR U1342 ( .A(in[34]), .B(in[1314]), .Z(n713) );
  XNOR U1343 ( .A(n714), .B(n713), .Z(n715) );
  XOR U1344 ( .A(in[994]), .B(n715), .Z(n1489) );
  XNOR U1345 ( .A(in[1379]), .B(n4542), .Z(n2002) );
  XOR U1346 ( .A(in[1578]), .B(in[618]), .Z(n717) );
  XNOR U1347 ( .A(in[938]), .B(in[298]), .Z(n716) );
  XNOR U1348 ( .A(n717), .B(n716), .Z(n718) );
  XNOR U1349 ( .A(in[1258]), .B(n718), .Z(n1071) );
  XOR U1350 ( .A(n719), .B(n1071), .Z(n4296) );
  XOR U1351 ( .A(in[1003]), .B(n4296), .Z(n1999) );
  NANDN U1352 ( .A(n2002), .B(n1999), .Z(n720) );
  XOR U1353 ( .A(n1593), .B(n720), .Z(out[1023]) );
  XOR U1354 ( .A(n722), .B(n721), .Z(n3985) );
  XOR U1355 ( .A(in[531]), .B(n3985), .Z(n1597) );
  XOR U1356 ( .A(in[35]), .B(in[675]), .Z(n724) );
  XNOR U1357 ( .A(in[355]), .B(in[1315]), .Z(n723) );
  XNOR U1358 ( .A(n724), .B(n723), .Z(n725) );
  XNOR U1359 ( .A(in[995]), .B(n725), .Z(n1492) );
  XOR U1360 ( .A(in[164]), .B(in[1444]), .Z(n727) );
  XNOR U1361 ( .A(in[804]), .B(in[1124]), .Z(n726) );
  XNOR U1362 ( .A(n727), .B(n726), .Z(n728) );
  XNOR U1363 ( .A(in[484]), .B(n728), .Z(n974) );
  XOR U1364 ( .A(n1492), .B(n974), .Z(n4546) );
  XNOR U1365 ( .A(in[1380]), .B(n4546), .Z(n4997) );
  XOR U1366 ( .A(in[1346]), .B(in[66]), .Z(n730) );
  XNOR U1367 ( .A(in[1026]), .B(in[386]), .Z(n729) );
  XNOR U1368 ( .A(n730), .B(n729), .Z(n731) );
  XNOR U1369 ( .A(in[706]), .B(n731), .Z(n1686) );
  XOR U1370 ( .A(in[1475]), .B(in[515]), .Z(n733) );
  XNOR U1371 ( .A(in[835]), .B(in[195]), .Z(n732) );
  XNOR U1372 ( .A(n733), .B(n732), .Z(n734) );
  XOR U1373 ( .A(in[1155]), .B(n734), .Z(n1411) );
  XOR U1374 ( .A(in[131]), .B(n3173), .Z(n4999) );
  OR U1375 ( .A(n4997), .B(n4999), .Z(n735) );
  XNOR U1376 ( .A(n1597), .B(n735), .Z(out[1024]) );
  XNOR U1377 ( .A(n737), .B(n736), .Z(n3989) );
  XOR U1378 ( .A(in[532]), .B(n3989), .Z(n1601) );
  XOR U1379 ( .A(in[36]), .B(in[676]), .Z(n739) );
  XNOR U1380 ( .A(in[356]), .B(in[1316]), .Z(n738) );
  XNOR U1381 ( .A(n739), .B(n738), .Z(n740) );
  XNOR U1382 ( .A(in[996]), .B(n740), .Z(n1495) );
  XOR U1383 ( .A(in[1445]), .B(in[165]), .Z(n742) );
  XNOR U1384 ( .A(in[805]), .B(in[1125]), .Z(n741) );
  XNOR U1385 ( .A(n742), .B(n741), .Z(n743) );
  XNOR U1386 ( .A(in[485]), .B(n743), .Z(n1018) );
  XOR U1387 ( .A(n1495), .B(n1018), .Z(n4552) );
  XNOR U1388 ( .A(in[1381]), .B(n4552), .Z(n5001) );
  XOR U1389 ( .A(in[1347]), .B(in[67]), .Z(n745) );
  XNOR U1390 ( .A(in[1027]), .B(in[387]), .Z(n744) );
  XNOR U1391 ( .A(n745), .B(n744), .Z(n746) );
  XNOR U1392 ( .A(in[707]), .B(n746), .Z(n1690) );
  XOR U1393 ( .A(in[1476]), .B(in[516]), .Z(n748) );
  XNOR U1394 ( .A(in[836]), .B(in[196]), .Z(n747) );
  XNOR U1395 ( .A(n748), .B(n747), .Z(n749) );
  XOR U1396 ( .A(in[1156]), .B(n749), .Z(n1413) );
  XOR U1397 ( .A(in[132]), .B(n3175), .Z(n5003) );
  OR U1398 ( .A(n5001), .B(n5003), .Z(n750) );
  XNOR U1399 ( .A(n1601), .B(n750), .Z(out[1025]) );
  XOR U1400 ( .A(n752), .B(n751), .Z(n2006) );
  XOR U1401 ( .A(in[533]), .B(n2006), .Z(n1605) );
  XOR U1402 ( .A(in[166]), .B(in[806]), .Z(n754) );
  XNOR U1403 ( .A(in[1126]), .B(in[486]), .Z(n753) );
  XNOR U1404 ( .A(n754), .B(n753), .Z(n755) );
  XNOR U1405 ( .A(in[1446]), .B(n755), .Z(n1031) );
  XOR U1406 ( .A(in[37]), .B(in[677]), .Z(n757) );
  XNOR U1407 ( .A(in[357]), .B(in[1317]), .Z(n756) );
  XNOR U1408 ( .A(n757), .B(n756), .Z(n758) );
  XNOR U1409 ( .A(in[997]), .B(n758), .Z(n1498) );
  XOR U1410 ( .A(n1031), .B(n1498), .Z(n4554) );
  XNOR U1411 ( .A(in[1382]), .B(n4554), .Z(n5005) );
  XOR U1412 ( .A(in[1348]), .B(in[68]), .Z(n760) );
  XNOR U1413 ( .A(in[1028]), .B(in[388]), .Z(n759) );
  XNOR U1414 ( .A(n760), .B(n759), .Z(n761) );
  XNOR U1415 ( .A(in[708]), .B(n761), .Z(n1694) );
  XOR U1416 ( .A(in[1477]), .B(in[517]), .Z(n763) );
  XNOR U1417 ( .A(in[837]), .B(in[197]), .Z(n762) );
  XNOR U1418 ( .A(n763), .B(n762), .Z(n764) );
  XOR U1419 ( .A(in[1157]), .B(n764), .Z(n1415) );
  XOR U1420 ( .A(in[133]), .B(n3177), .Z(n5007) );
  OR U1421 ( .A(n5005), .B(n5007), .Z(n765) );
  XNOR U1422 ( .A(n1605), .B(n765), .Z(out[1026]) );
  XOR U1423 ( .A(n767), .B(n766), .Z(n2008) );
  XOR U1424 ( .A(in[534]), .B(n2008), .Z(n1609) );
  XOR U1425 ( .A(in[38]), .B(in[678]), .Z(n769) );
  XNOR U1426 ( .A(in[358]), .B(in[1318]), .Z(n768) );
  XNOR U1427 ( .A(n769), .B(n768), .Z(n770) );
  XNOR U1428 ( .A(in[998]), .B(n770), .Z(n1502) );
  XOR U1429 ( .A(in[167]), .B(in[807]), .Z(n772) );
  XNOR U1430 ( .A(in[1127]), .B(in[487]), .Z(n771) );
  XNOR U1431 ( .A(n772), .B(n771), .Z(n773) );
  XNOR U1432 ( .A(in[1447]), .B(n773), .Z(n1044) );
  XOR U1433 ( .A(n1502), .B(n1044), .Z(n4335) );
  XNOR U1434 ( .A(in[1383]), .B(n4335), .Z(n5009) );
  XOR U1435 ( .A(in[1349]), .B(in[69]), .Z(n775) );
  XNOR U1436 ( .A(in[1029]), .B(in[389]), .Z(n774) );
  XNOR U1437 ( .A(n775), .B(n774), .Z(n776) );
  XNOR U1438 ( .A(in[709]), .B(n776), .Z(n1698) );
  XOR U1439 ( .A(in[1478]), .B(in[518]), .Z(n778) );
  XNOR U1440 ( .A(in[838]), .B(in[198]), .Z(n777) );
  XNOR U1441 ( .A(n778), .B(n777), .Z(n779) );
  XOR U1442 ( .A(in[1158]), .B(n779), .Z(n1417) );
  XOR U1443 ( .A(in[134]), .B(n3179), .Z(n5011) );
  OR U1444 ( .A(n5009), .B(n5011), .Z(n780) );
  XNOR U1445 ( .A(n1609), .B(n780), .Z(out[1027]) );
  XNOR U1446 ( .A(n782), .B(n781), .Z(n4001) );
  XOR U1447 ( .A(in[535]), .B(n4001), .Z(n1613) );
  XOR U1448 ( .A(in[168]), .B(in[1448]), .Z(n784) );
  XNOR U1449 ( .A(in[1128]), .B(in[808]), .Z(n783) );
  XNOR U1450 ( .A(n784), .B(n783), .Z(n785) );
  XNOR U1451 ( .A(in[488]), .B(n785), .Z(n1057) );
  XOR U1452 ( .A(in[39]), .B(in[679]), .Z(n787) );
  XNOR U1453 ( .A(in[359]), .B(in[1319]), .Z(n786) );
  XNOR U1454 ( .A(n787), .B(n786), .Z(n788) );
  XNOR U1455 ( .A(in[999]), .B(n788), .Z(n1507) );
  XOR U1456 ( .A(n1057), .B(n1507), .Z(n4337) );
  XNOR U1457 ( .A(in[1384]), .B(n4337), .Z(n5013) );
  XOR U1458 ( .A(in[1350]), .B(in[70]), .Z(n790) );
  XNOR U1459 ( .A(in[1030]), .B(in[390]), .Z(n789) );
  XNOR U1460 ( .A(n790), .B(n789), .Z(n791) );
  XNOR U1461 ( .A(in[710]), .B(n791), .Z(n1702) );
  XOR U1462 ( .A(in[199]), .B(in[1479]), .Z(n793) );
  XNOR U1463 ( .A(in[1159]), .B(in[839]), .Z(n792) );
  XNOR U1464 ( .A(n793), .B(n792), .Z(n794) );
  XOR U1465 ( .A(in[519]), .B(n794), .Z(n1419) );
  XOR U1466 ( .A(in[135]), .B(n3181), .Z(n5015) );
  OR U1467 ( .A(n5013), .B(n5015), .Z(n795) );
  XNOR U1468 ( .A(n1613), .B(n795), .Z(out[1028]) );
  XNOR U1469 ( .A(n797), .B(n796), .Z(n4005) );
  XOR U1470 ( .A(in[536]), .B(n4005), .Z(n1617) );
  XOR U1471 ( .A(in[169]), .B(in[1449]), .Z(n799) );
  XNOR U1472 ( .A(in[1129]), .B(in[809]), .Z(n798) );
  XNOR U1473 ( .A(n799), .B(n798), .Z(n800) );
  XNOR U1474 ( .A(in[489]), .B(n800), .Z(n1070) );
  XOR U1475 ( .A(in[680]), .B(in[1320]), .Z(n802) );
  XNOR U1476 ( .A(in[40]), .B(in[360]), .Z(n801) );
  XNOR U1477 ( .A(n802), .B(n801), .Z(n803) );
  XNOR U1478 ( .A(in[1000]), .B(n803), .Z(n1511) );
  XOR U1479 ( .A(n1070), .B(n1511), .Z(n4343) );
  XNOR U1480 ( .A(in[1385]), .B(n4343), .Z(n5017) );
  XOR U1481 ( .A(in[1351]), .B(in[711]), .Z(n805) );
  XNOR U1482 ( .A(in[1031]), .B(in[391]), .Z(n804) );
  XNOR U1483 ( .A(n805), .B(n804), .Z(n806) );
  XNOR U1484 ( .A(in[71]), .B(n806), .Z(n1706) );
  XOR U1485 ( .A(in[1480]), .B(in[520]), .Z(n808) );
  XNOR U1486 ( .A(in[840]), .B(in[200]), .Z(n807) );
  XNOR U1487 ( .A(n808), .B(n807), .Z(n809) );
  XOR U1488 ( .A(in[1160]), .B(n809), .Z(n1424) );
  XOR U1489 ( .A(in[136]), .B(n3183), .Z(n5019) );
  OR U1490 ( .A(n5017), .B(n5019), .Z(n810) );
  XNOR U1491 ( .A(n1617), .B(n810), .Z(out[1029]) );
  XOR U1492 ( .A(in[1341]), .B(in[61]), .Z(n812) );
  XNOR U1493 ( .A(in[701]), .B(in[381]), .Z(n811) );
  XNOR U1494 ( .A(n812), .B(n811), .Z(n813) );
  XNOR U1495 ( .A(in[1021]), .B(n813), .Z(n1127) );
  XOR U1496 ( .A(n814), .B(n1127), .Z(n3961) );
  XOR U1497 ( .A(in[637]), .B(n3961), .Z(n2708) );
  IV U1498 ( .A(n2708), .Z(n2797) );
  XOR U1499 ( .A(n816), .B(n815), .Z(n4057) );
  XOR U1500 ( .A(in[228]), .B(n4057), .Z(n3156) );
  XOR U1501 ( .A(in[1512]), .B(in[552]), .Z(n818) );
  XNOR U1502 ( .A(in[872]), .B(in[232]), .Z(n817) );
  XNOR U1503 ( .A(n818), .B(n817), .Z(n819) );
  XNOR U1504 ( .A(in[1192]), .B(n819), .Z(n1516) );
  XNOR U1505 ( .A(n820), .B(n1516), .Z(n4097) );
  IV U1506 ( .A(n4097), .Z(n1276) );
  XOR U1507 ( .A(in[1448]), .B(n1276), .Z(n3154) );
  NANDN U1508 ( .A(n3156), .B(n3154), .Z(n821) );
  XOR U1509 ( .A(n2797), .B(n821), .Z(out[102]) );
  XNOR U1510 ( .A(n823), .B(n822), .Z(n4009) );
  XOR U1511 ( .A(in[537]), .B(n4009), .Z(n1621) );
  XOR U1512 ( .A(in[1352]), .B(in[712]), .Z(n825) );
  XNOR U1513 ( .A(in[1032]), .B(in[392]), .Z(n824) );
  XNOR U1514 ( .A(n825), .B(n824), .Z(n826) );
  XNOR U1515 ( .A(in[72]), .B(n826), .Z(n1711) );
  XOR U1516 ( .A(in[1481]), .B(in[521]), .Z(n828) );
  XNOR U1517 ( .A(in[841]), .B(in[201]), .Z(n827) );
  XNOR U1518 ( .A(n828), .B(n827), .Z(n829) );
  XOR U1519 ( .A(in[1161]), .B(n829), .Z(n1426) );
  XOR U1520 ( .A(in[137]), .B(n3185), .Z(n5023) );
  XOR U1521 ( .A(in[681]), .B(in[1321]), .Z(n831) );
  XNOR U1522 ( .A(in[41]), .B(in[361]), .Z(n830) );
  XNOR U1523 ( .A(n831), .B(n830), .Z(n832) );
  XNOR U1524 ( .A(in[1001]), .B(n832), .Z(n1515) );
  XOR U1525 ( .A(in[170]), .B(in[1450]), .Z(n834) );
  XNOR U1526 ( .A(in[1130]), .B(in[810]), .Z(n833) );
  XNOR U1527 ( .A(n834), .B(n833), .Z(n835) );
  XNOR U1528 ( .A(in[490]), .B(n835), .Z(n1086) );
  XOR U1529 ( .A(n1515), .B(n1086), .Z(n4345) );
  XOR U1530 ( .A(in[1386]), .B(n4345), .Z(n5020) );
  NANDN U1531 ( .A(n5023), .B(n5020), .Z(n836) );
  XNOR U1532 ( .A(n1621), .B(n836), .Z(out[1030]) );
  XOR U1533 ( .A(n838), .B(n837), .Z(n2015) );
  XOR U1534 ( .A(in[538]), .B(n2015), .Z(n1625) );
  XOR U1535 ( .A(in[1353]), .B(in[393]), .Z(n840) );
  XNOR U1536 ( .A(in[713]), .B(in[73]), .Z(n839) );
  XNOR U1537 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1538 ( .A(in[1033]), .B(n841), .Z(n1715) );
  XOR U1539 ( .A(in[1482]), .B(in[522]), .Z(n843) );
  XNOR U1540 ( .A(in[842]), .B(in[202]), .Z(n842) );
  XNOR U1541 ( .A(n843), .B(n842), .Z(n844) );
  XOR U1542 ( .A(in[1162]), .B(n844), .Z(n1428) );
  XOR U1543 ( .A(in[138]), .B(n3187), .Z(n5027) );
  XOR U1544 ( .A(in[811]), .B(in[491]), .Z(n846) );
  XNOR U1545 ( .A(in[1451]), .B(in[1131]), .Z(n845) );
  XNOR U1546 ( .A(n846), .B(n845), .Z(n847) );
  XNOR U1547 ( .A(in[171]), .B(n847), .Z(n1099) );
  XOR U1548 ( .A(in[682]), .B(in[1322]), .Z(n849) );
  XNOR U1549 ( .A(in[42]), .B(in[362]), .Z(n848) );
  XNOR U1550 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U1551 ( .A(in[1002]), .B(n850), .Z(n1520) );
  XOR U1552 ( .A(n1099), .B(n1520), .Z(n4347) );
  XOR U1553 ( .A(in[1387]), .B(n4347), .Z(n5024) );
  NANDN U1554 ( .A(n5027), .B(n5024), .Z(n851) );
  XNOR U1555 ( .A(n1625), .B(n851), .Z(out[1031]) );
  XOR U1556 ( .A(n853), .B(n852), .Z(n2018) );
  XOR U1557 ( .A(in[539]), .B(n2018), .Z(n1630) );
  XOR U1558 ( .A(in[1354]), .B(in[714]), .Z(n855) );
  XNOR U1559 ( .A(in[74]), .B(in[394]), .Z(n854) );
  XNOR U1560 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1561 ( .A(in[1034]), .B(n856), .Z(n1719) );
  XOR U1562 ( .A(in[1483]), .B(in[523]), .Z(n858) );
  XNOR U1563 ( .A(in[843]), .B(in[203]), .Z(n857) );
  XNOR U1564 ( .A(n858), .B(n857), .Z(n859) );
  XOR U1565 ( .A(in[1163]), .B(n859), .Z(n1430) );
  XOR U1566 ( .A(n2294), .B(in[139]), .Z(n5031) );
  XOR U1567 ( .A(in[812]), .B(in[492]), .Z(n861) );
  XNOR U1568 ( .A(in[1452]), .B(in[1132]), .Z(n860) );
  XNOR U1569 ( .A(n861), .B(n860), .Z(n862) );
  XNOR U1570 ( .A(in[172]), .B(n862), .Z(n1119) );
  XOR U1571 ( .A(in[683]), .B(in[1323]), .Z(n864) );
  XNOR U1572 ( .A(in[43]), .B(in[363]), .Z(n863) );
  XNOR U1573 ( .A(n864), .B(n863), .Z(n865) );
  XNOR U1574 ( .A(in[1003]), .B(n865), .Z(n1524) );
  XOR U1575 ( .A(n1119), .B(n1524), .Z(n4350) );
  XOR U1576 ( .A(in[1388]), .B(n4350), .Z(n5028) );
  NANDN U1577 ( .A(n5031), .B(n5028), .Z(n866) );
  XNOR U1578 ( .A(n1630), .B(n866), .Z(out[1032]) );
  XOR U1579 ( .A(n868), .B(n867), .Z(n4021) );
  XOR U1580 ( .A(in[540]), .B(n4021), .Z(n1634) );
  XOR U1581 ( .A(in[1355]), .B(in[715]), .Z(n870) );
  XNOR U1582 ( .A(in[1035]), .B(in[395]), .Z(n869) );
  XNOR U1583 ( .A(n870), .B(n869), .Z(n871) );
  XNOR U1584 ( .A(in[75]), .B(n871), .Z(n1723) );
  XOR U1585 ( .A(in[1484]), .B(in[524]), .Z(n873) );
  XNOR U1586 ( .A(in[844]), .B(in[204]), .Z(n872) );
  XNOR U1587 ( .A(n873), .B(n872), .Z(n874) );
  XOR U1588 ( .A(in[1164]), .B(n874), .Z(n1432) );
  XOR U1589 ( .A(in[140]), .B(n3194), .Z(n5035) );
  XOR U1590 ( .A(in[1324]), .B(in[44]), .Z(n876) );
  XNOR U1591 ( .A(in[684]), .B(in[364]), .Z(n875) );
  XNOR U1592 ( .A(n876), .B(n875), .Z(n877) );
  XNOR U1593 ( .A(in[1004]), .B(n877), .Z(n1527) );
  XOR U1594 ( .A(in[813]), .B(in[493]), .Z(n879) );
  XNOR U1595 ( .A(in[1453]), .B(in[1133]), .Z(n878) );
  XNOR U1596 ( .A(n879), .B(n878), .Z(n880) );
  XNOR U1597 ( .A(in[173]), .B(n880), .Z(n1132) );
  XOR U1598 ( .A(n1527), .B(n1132), .Z(n4353) );
  XOR U1599 ( .A(in[1389]), .B(n4353), .Z(n5032) );
  NANDN U1600 ( .A(n5035), .B(n5032), .Z(n881) );
  XNOR U1601 ( .A(n1634), .B(n881), .Z(out[1033]) );
  XOR U1602 ( .A(n883), .B(n882), .Z(n4029) );
  XOR U1603 ( .A(in[541]), .B(n4029), .Z(n1638) );
  XOR U1604 ( .A(in[76]), .B(in[1036]), .Z(n885) );
  XNOR U1605 ( .A(in[716]), .B(in[396]), .Z(n884) );
  XNOR U1606 ( .A(n885), .B(n884), .Z(n886) );
  XNOR U1607 ( .A(in[1356]), .B(n886), .Z(n1727) );
  XOR U1608 ( .A(in[1485]), .B(in[525]), .Z(n888) );
  XNOR U1609 ( .A(in[845]), .B(in[205]), .Z(n887) );
  XNOR U1610 ( .A(n888), .B(n887), .Z(n889) );
  XOR U1611 ( .A(in[1165]), .B(n889), .Z(n1434) );
  XOR U1612 ( .A(in[141]), .B(n3196), .Z(n5043) );
  XOR U1613 ( .A(in[1325]), .B(in[45]), .Z(n891) );
  XNOR U1614 ( .A(in[685]), .B(in[365]), .Z(n890) );
  XNOR U1615 ( .A(n891), .B(n890), .Z(n892) );
  XNOR U1616 ( .A(in[1005]), .B(n892), .Z(n1531) );
  XOR U1617 ( .A(in[814]), .B(in[494]), .Z(n894) );
  XNOR U1618 ( .A(in[1454]), .B(in[1134]), .Z(n893) );
  XNOR U1619 ( .A(n894), .B(n893), .Z(n895) );
  XNOR U1620 ( .A(in[174]), .B(n895), .Z(n1145) );
  XOR U1621 ( .A(n1531), .B(n1145), .Z(n4356) );
  XOR U1622 ( .A(in[1390]), .B(n4356), .Z(n5040) );
  NANDN U1623 ( .A(n5043), .B(n5040), .Z(n896) );
  XNOR U1624 ( .A(n1638), .B(n896), .Z(out[1034]) );
  XOR U1625 ( .A(n898), .B(n897), .Z(n4033) );
  XOR U1626 ( .A(in[542]), .B(n4033), .Z(n1642) );
  XOR U1627 ( .A(in[77]), .B(in[1037]), .Z(n900) );
  XNOR U1628 ( .A(in[717]), .B(in[397]), .Z(n899) );
  XNOR U1629 ( .A(n900), .B(n899), .Z(n901) );
  XNOR U1630 ( .A(in[1357]), .B(n901), .Z(n1731) );
  XOR U1631 ( .A(in[1486]), .B(in[526]), .Z(n903) );
  XNOR U1632 ( .A(in[846]), .B(in[206]), .Z(n902) );
  XNOR U1633 ( .A(n903), .B(n902), .Z(n904) );
  XOR U1634 ( .A(in[1166]), .B(n904), .Z(n1436) );
  XOR U1635 ( .A(in[142]), .B(n3199), .Z(n5047) );
  XOR U1636 ( .A(in[1326]), .B(in[46]), .Z(n906) );
  XNOR U1637 ( .A(in[686]), .B(in[366]), .Z(n905) );
  XNOR U1638 ( .A(n906), .B(n905), .Z(n907) );
  XNOR U1639 ( .A(in[1006]), .B(n907), .Z(n1535) );
  XOR U1640 ( .A(in[815]), .B(in[495]), .Z(n909) );
  XNOR U1641 ( .A(in[1455]), .B(in[1135]), .Z(n908) );
  XNOR U1642 ( .A(n909), .B(n908), .Z(n910) );
  XNOR U1643 ( .A(in[175]), .B(n910), .Z(n1158) );
  XOR U1644 ( .A(n1535), .B(n1158), .Z(n4358) );
  XOR U1645 ( .A(in[1391]), .B(n4358), .Z(n5044) );
  NANDN U1646 ( .A(n5047), .B(n5044), .Z(n911) );
  XNOR U1647 ( .A(n1642), .B(n911), .Z(out[1035]) );
  XOR U1648 ( .A(n913), .B(n912), .Z(n4037) );
  XOR U1649 ( .A(in[543]), .B(n4037), .Z(n1646) );
  XOR U1650 ( .A(in[78]), .B(in[1038]), .Z(n915) );
  XNOR U1651 ( .A(in[718]), .B(in[398]), .Z(n914) );
  XNOR U1652 ( .A(n915), .B(n914), .Z(n916) );
  XNOR U1653 ( .A(in[1358]), .B(n916), .Z(n1735) );
  XOR U1654 ( .A(in[1487]), .B(in[527]), .Z(n918) );
  XNOR U1655 ( .A(in[847]), .B(in[207]), .Z(n917) );
  XNOR U1656 ( .A(n918), .B(n917), .Z(n919) );
  XOR U1657 ( .A(in[1167]), .B(n919), .Z(n1438) );
  XOR U1658 ( .A(in[143]), .B(n3202), .Z(n5051) );
  XOR U1659 ( .A(in[816]), .B(in[496]), .Z(n921) );
  XNOR U1660 ( .A(in[1456]), .B(in[1136]), .Z(n920) );
  XNOR U1661 ( .A(n921), .B(n920), .Z(n922) );
  XNOR U1662 ( .A(in[176]), .B(n922), .Z(n1173) );
  XOR U1663 ( .A(in[1327]), .B(in[47]), .Z(n924) );
  XNOR U1664 ( .A(in[687]), .B(in[367]), .Z(n923) );
  XNOR U1665 ( .A(n924), .B(n923), .Z(n925) );
  XNOR U1666 ( .A(in[1007]), .B(n925), .Z(n1539) );
  XOR U1667 ( .A(n1173), .B(n1539), .Z(n4361) );
  XOR U1668 ( .A(in[1392]), .B(n4361), .Z(n5048) );
  NANDN U1669 ( .A(n5051), .B(n5048), .Z(n926) );
  XNOR U1670 ( .A(n1646), .B(n926), .Z(out[1036]) );
  XOR U1671 ( .A(n928), .B(n927), .Z(n4041) );
  XOR U1672 ( .A(in[544]), .B(n4041), .Z(n1650) );
  XOR U1673 ( .A(in[79]), .B(in[1039]), .Z(n930) );
  XNOR U1674 ( .A(in[719]), .B(in[399]), .Z(n929) );
  XNOR U1675 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U1676 ( .A(in[1359]), .B(n931), .Z(n1739) );
  XOR U1677 ( .A(in[1488]), .B(in[528]), .Z(n933) );
  XNOR U1678 ( .A(in[848]), .B(in[208]), .Z(n932) );
  XNOR U1679 ( .A(n933), .B(n932), .Z(n934) );
  XOR U1680 ( .A(n1739), .B(n232), .Z(n3205) );
  XOR U1681 ( .A(in[144]), .B(n3205), .Z(n5055) );
  XOR U1682 ( .A(in[817]), .B(in[497]), .Z(n936) );
  XNOR U1683 ( .A(in[1457]), .B(in[1137]), .Z(n935) );
  XNOR U1684 ( .A(n936), .B(n935), .Z(n937) );
  XNOR U1685 ( .A(in[177]), .B(n937), .Z(n1188) );
  XOR U1686 ( .A(in[1328]), .B(in[48]), .Z(n939) );
  XNOR U1687 ( .A(in[688]), .B(in[368]), .Z(n938) );
  XNOR U1688 ( .A(n939), .B(n938), .Z(n940) );
  XNOR U1689 ( .A(in[1008]), .B(n940), .Z(n1543) );
  XOR U1690 ( .A(n1188), .B(n1543), .Z(n4364) );
  XOR U1691 ( .A(in[1393]), .B(n4364), .Z(n5052) );
  NANDN U1692 ( .A(n5055), .B(n5052), .Z(n941) );
  XNOR U1693 ( .A(n1650), .B(n941), .Z(out[1037]) );
  XOR U1694 ( .A(n943), .B(n942), .Z(n4045) );
  XOR U1695 ( .A(in[545]), .B(n4045), .Z(n1654) );
  XOR U1696 ( .A(in[80]), .B(in[1040]), .Z(n945) );
  XNOR U1697 ( .A(in[720]), .B(in[400]), .Z(n944) );
  XNOR U1698 ( .A(n945), .B(n944), .Z(n946) );
  XNOR U1699 ( .A(in[1360]), .B(n946), .Z(n1743) );
  XOR U1700 ( .A(in[1489]), .B(in[529]), .Z(n948) );
  XNOR U1701 ( .A(in[849]), .B(in[209]), .Z(n947) );
  XNOR U1702 ( .A(n948), .B(n947), .Z(n949) );
  XOR U1703 ( .A(in[1169]), .B(n949), .Z(n1441) );
  XOR U1704 ( .A(in[145]), .B(n3208), .Z(n5059) );
  XOR U1705 ( .A(in[818]), .B(in[498]), .Z(n951) );
  XNOR U1706 ( .A(in[1458]), .B(in[1138]), .Z(n950) );
  XNOR U1707 ( .A(n951), .B(n950), .Z(n952) );
  XNOR U1708 ( .A(in[178]), .B(n952), .Z(n1203) );
  XOR U1709 ( .A(in[1329]), .B(in[49]), .Z(n954) );
  XNOR U1710 ( .A(in[689]), .B(in[369]), .Z(n953) );
  XNOR U1711 ( .A(n954), .B(n953), .Z(n955) );
  XNOR U1712 ( .A(in[1009]), .B(n955), .Z(n1549) );
  XOR U1713 ( .A(n1203), .B(n1549), .Z(n4367) );
  XOR U1714 ( .A(in[1394]), .B(n4367), .Z(n5056) );
  NANDN U1715 ( .A(n5059), .B(n5056), .Z(n956) );
  XNOR U1716 ( .A(n1654), .B(n956), .Z(out[1038]) );
  IV U1717 ( .A(n4049), .Z(n3395) );
  XOR U1718 ( .A(n3395), .B(in[546]), .Z(n1658) );
  XOR U1719 ( .A(in[81]), .B(in[1041]), .Z(n958) );
  XNOR U1720 ( .A(in[721]), .B(in[401]), .Z(n957) );
  XNOR U1721 ( .A(n958), .B(n957), .Z(n959) );
  XNOR U1722 ( .A(in[1361]), .B(n959), .Z(n1747) );
  XOR U1723 ( .A(in[1490]), .B(in[530]), .Z(n961) );
  XNOR U1724 ( .A(in[850]), .B(in[210]), .Z(n960) );
  XNOR U1725 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1726 ( .A(in[1170]), .B(n962), .Z(n1445) );
  XOR U1727 ( .A(in[146]), .B(n3211), .Z(n5063) );
  XOR U1728 ( .A(in[1330]), .B(in[50]), .Z(n964) );
  XNOR U1729 ( .A(in[690]), .B(in[370]), .Z(n963) );
  XNOR U1730 ( .A(n964), .B(n963), .Z(n965) );
  XNOR U1731 ( .A(in[1010]), .B(n965), .Z(n1553) );
  XOR U1732 ( .A(in[819]), .B(in[499]), .Z(n967) );
  XNOR U1733 ( .A(in[1459]), .B(in[1139]), .Z(n966) );
  XNOR U1734 ( .A(n967), .B(n966), .Z(n968) );
  XNOR U1735 ( .A(in[179]), .B(n968), .Z(n1218) );
  XOR U1736 ( .A(n1553), .B(n1218), .Z(n4374) );
  XOR U1737 ( .A(in[1395]), .B(n4374), .Z(n5060) );
  NANDN U1738 ( .A(n5063), .B(n5060), .Z(n969) );
  XOR U1739 ( .A(n1658), .B(n969), .Z(out[1039]) );
  XOR U1740 ( .A(in[1342]), .B(in[62]), .Z(n971) );
  XNOR U1741 ( .A(in[702]), .B(in[382]), .Z(n970) );
  XNOR U1742 ( .A(n971), .B(n970), .Z(n972) );
  XNOR U1743 ( .A(in[1022]), .B(n972), .Z(n1140) );
  XOR U1744 ( .A(n973), .B(n1140), .Z(n3965) );
  XOR U1745 ( .A(in[638]), .B(n3965), .Z(n2710) );
  IV U1746 ( .A(n2710), .Z(n2799) );
  XOR U1747 ( .A(n975), .B(n974), .Z(n4061) );
  XOR U1748 ( .A(in[229]), .B(n4061), .Z(n3167) );
  XOR U1749 ( .A(in[1513]), .B(in[553]), .Z(n977) );
  XNOR U1750 ( .A(in[873]), .B(in[233]), .Z(n976) );
  XNOR U1751 ( .A(n977), .B(n976), .Z(n978) );
  XNOR U1752 ( .A(in[1193]), .B(n978), .Z(n1519) );
  XNOR U1753 ( .A(n979), .B(n1519), .Z(n4101) );
  IV U1754 ( .A(n4101), .Z(n1288) );
  XOR U1755 ( .A(in[1449]), .B(n1288), .Z(n3164) );
  NANDN U1756 ( .A(n3167), .B(n3164), .Z(n980) );
  XOR U1757 ( .A(n2799), .B(n980), .Z(out[103]) );
  XOR U1758 ( .A(n3398), .B(in[547]), .Z(n1662) );
  XOR U1759 ( .A(in[1042]), .B(in[402]), .Z(n982) );
  XNOR U1760 ( .A(in[722]), .B(in[82]), .Z(n981) );
  XNOR U1761 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1762 ( .A(in[1362]), .B(n983), .Z(n1752) );
  XOR U1763 ( .A(in[851]), .B(in[1171]), .Z(n985) );
  XNOR U1764 ( .A(in[1491]), .B(in[211]), .Z(n984) );
  XNOR U1765 ( .A(n985), .B(n984), .Z(n986) );
  XOR U1766 ( .A(in[531]), .B(n986), .Z(n1447) );
  IV U1767 ( .A(n3214), .Z(n4006) );
  XNOR U1768 ( .A(in[147]), .B(n4006), .Z(n5066) );
  XOR U1769 ( .A(in[820]), .B(in[500]), .Z(n988) );
  XNOR U1770 ( .A(in[1460]), .B(in[1140]), .Z(n987) );
  XNOR U1771 ( .A(n988), .B(n987), .Z(n989) );
  XNOR U1772 ( .A(in[180]), .B(n989), .Z(n1233) );
  XOR U1773 ( .A(in[1331]), .B(in[51]), .Z(n991) );
  XNOR U1774 ( .A(in[691]), .B(in[371]), .Z(n990) );
  XNOR U1775 ( .A(n991), .B(n990), .Z(n992) );
  XNOR U1776 ( .A(in[1011]), .B(n992), .Z(n1557) );
  XOR U1777 ( .A(n1233), .B(n1557), .Z(n4377) );
  XOR U1778 ( .A(in[1396]), .B(n4377), .Z(n5065) );
  NANDN U1779 ( .A(n5066), .B(n5065), .Z(n993) );
  XOR U1780 ( .A(n1662), .B(n993), .Z(out[1040]) );
  IV U1781 ( .A(n4057), .Z(n3402) );
  XOR U1782 ( .A(n3402), .B(in[548]), .Z(n1666) );
  XOR U1783 ( .A(in[83]), .B(in[1043]), .Z(n995) );
  XNOR U1784 ( .A(in[723]), .B(in[403]), .Z(n994) );
  XNOR U1785 ( .A(n995), .B(n994), .Z(n996) );
  XNOR U1786 ( .A(in[1363]), .B(n996), .Z(n1756) );
  XOR U1787 ( .A(in[852]), .B(in[1172]), .Z(n998) );
  XNOR U1788 ( .A(in[1492]), .B(in[212]), .Z(n997) );
  XNOR U1789 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1790 ( .A(in[532]), .B(n999), .Z(n1449) );
  IV U1791 ( .A(n3217), .Z(n4010) );
  XNOR U1792 ( .A(in[148]), .B(n4010), .Z(n5069) );
  XOR U1793 ( .A(in[821]), .B(in[501]), .Z(n1001) );
  XNOR U1794 ( .A(in[1461]), .B(in[1141]), .Z(n1000) );
  XNOR U1795 ( .A(n1001), .B(n1000), .Z(n1002) );
  XNOR U1796 ( .A(in[181]), .B(n1002), .Z(n1248) );
  XOR U1797 ( .A(in[1332]), .B(in[52]), .Z(n1004) );
  XNOR U1798 ( .A(in[692]), .B(in[372]), .Z(n1003) );
  XNOR U1799 ( .A(n1004), .B(n1003), .Z(n1005) );
  XNOR U1800 ( .A(in[1012]), .B(n1005), .Z(n1561) );
  XOR U1801 ( .A(n1248), .B(n1561), .Z(n4380) );
  XOR U1802 ( .A(in[1397]), .B(n4380), .Z(n5068) );
  NANDN U1803 ( .A(n5069), .B(n5068), .Z(n1006) );
  XOR U1804 ( .A(n1666), .B(n1006), .Z(out[1041]) );
  IV U1805 ( .A(n4061), .Z(n3406) );
  XOR U1806 ( .A(n3406), .B(in[549]), .Z(n1671) );
  XOR U1807 ( .A(in[853]), .B(in[1173]), .Z(n1008) );
  XNOR U1808 ( .A(in[1493]), .B(in[213]), .Z(n1007) );
  XNOR U1809 ( .A(n1008), .B(n1007), .Z(n1009) );
  XOR U1810 ( .A(in[533]), .B(n1009), .Z(n1451) );
  IV U1811 ( .A(n2756), .Z(n4014) );
  XNOR U1812 ( .A(in[149]), .B(n4014), .Z(n5072) );
  XOR U1813 ( .A(in[822]), .B(in[502]), .Z(n1012) );
  XNOR U1814 ( .A(in[1462]), .B(in[1142]), .Z(n1011) );
  XNOR U1815 ( .A(n1012), .B(n1011), .Z(n1013) );
  XNOR U1816 ( .A(in[182]), .B(n1013), .Z(n1263) );
  XOR U1817 ( .A(in[1333]), .B(in[53]), .Z(n1015) );
  XNOR U1818 ( .A(in[693]), .B(in[373]), .Z(n1014) );
  XNOR U1819 ( .A(n1015), .B(n1014), .Z(n1016) );
  XNOR U1820 ( .A(in[1013]), .B(n1016), .Z(n1565) );
  XOR U1821 ( .A(n1263), .B(n1565), .Z(n4383) );
  XOR U1822 ( .A(in[1398]), .B(n4383), .Z(n5071) );
  NANDN U1823 ( .A(n5072), .B(n5071), .Z(n1017) );
  XOR U1824 ( .A(n1671), .B(n1017), .Z(out[1042]) );
  XOR U1825 ( .A(n1019), .B(n1018), .Z(n2037) );
  XOR U1826 ( .A(in[550]), .B(n2037), .Z(n1675) );
  XOR U1827 ( .A(in[854]), .B(in[1174]), .Z(n1021) );
  XNOR U1828 ( .A(in[1494]), .B(in[214]), .Z(n1020) );
  XNOR U1829 ( .A(n1021), .B(n1020), .Z(n1022) );
  XOR U1830 ( .A(in[534]), .B(n1022), .Z(n1453) );
  XOR U1831 ( .A(in[150]), .B(n2773), .Z(n5076) );
  XOR U1832 ( .A(in[823]), .B(in[503]), .Z(n1025) );
  XNOR U1833 ( .A(in[1463]), .B(in[1143]), .Z(n1024) );
  XNOR U1834 ( .A(n1025), .B(n1024), .Z(n1026) );
  XNOR U1835 ( .A(in[183]), .B(n1026), .Z(n1275) );
  XOR U1836 ( .A(in[1334]), .B(in[54]), .Z(n1028) );
  XNOR U1837 ( .A(in[694]), .B(in[374]), .Z(n1027) );
  XNOR U1838 ( .A(n1028), .B(n1027), .Z(n1029) );
  XNOR U1839 ( .A(in[1014]), .B(n1029), .Z(n1569) );
  XOR U1840 ( .A(n1275), .B(n1569), .Z(n4386) );
  XOR U1841 ( .A(in[1399]), .B(n4386), .Z(n5073) );
  NANDN U1842 ( .A(n5076), .B(n5073), .Z(n1030) );
  XNOR U1843 ( .A(n1675), .B(n1030), .Z(out[1043]) );
  XOR U1844 ( .A(n1032), .B(n1031), .Z(n2040) );
  XOR U1845 ( .A(in[551]), .B(n2040), .Z(n1679) );
  XOR U1846 ( .A(in[855]), .B(in[1175]), .Z(n1034) );
  XNOR U1847 ( .A(in[1495]), .B(in[215]), .Z(n1033) );
  XNOR U1848 ( .A(n1034), .B(n1033), .Z(n1035) );
  XOR U1849 ( .A(in[535]), .B(n1035), .Z(n1455) );
  XOR U1850 ( .A(in[151]), .B(n2780), .Z(n5083) );
  XOR U1851 ( .A(in[824]), .B(in[504]), .Z(n1038) );
  XNOR U1852 ( .A(in[1464]), .B(in[1144]), .Z(n1037) );
  XNOR U1853 ( .A(n1038), .B(n1037), .Z(n1039) );
  XNOR U1854 ( .A(in[184]), .B(n1039), .Z(n1281) );
  XOR U1855 ( .A(in[1335]), .B(in[55]), .Z(n1041) );
  XNOR U1856 ( .A(in[695]), .B(in[375]), .Z(n1040) );
  XNOR U1857 ( .A(n1041), .B(n1040), .Z(n1042) );
  XNOR U1858 ( .A(in[1015]), .B(n1042), .Z(n1573) );
  XOR U1859 ( .A(n1281), .B(n1573), .Z(n4388) );
  XOR U1860 ( .A(in[1400]), .B(n4388), .Z(n5082) );
  NANDN U1861 ( .A(n5083), .B(n5082), .Z(n1043) );
  XNOR U1862 ( .A(n1679), .B(n1043), .Z(out[1044]) );
  XOR U1863 ( .A(n1045), .B(n1044), .Z(n2044) );
  XOR U1864 ( .A(in[552]), .B(n2044), .Z(n1683) );
  XOR U1865 ( .A(in[856]), .B(in[1176]), .Z(n1047) );
  XNOR U1866 ( .A(in[1496]), .B(in[216]), .Z(n1046) );
  XNOR U1867 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1868 ( .A(in[536]), .B(n1048), .Z(n1459) );
  XOR U1869 ( .A(in[152]), .B(n2794), .Z(n5086) );
  XOR U1870 ( .A(in[825]), .B(in[505]), .Z(n1051) );
  XNOR U1871 ( .A(in[1465]), .B(in[1145]), .Z(n1050) );
  XNOR U1872 ( .A(n1051), .B(n1050), .Z(n1052) );
  XNOR U1873 ( .A(in[185]), .B(n1052), .Z(n1293) );
  XOR U1874 ( .A(in[1336]), .B(in[56]), .Z(n1054) );
  XNOR U1875 ( .A(in[696]), .B(in[376]), .Z(n1053) );
  XNOR U1876 ( .A(n1054), .B(n1053), .Z(n1055) );
  XNOR U1877 ( .A(in[1016]), .B(n1055), .Z(n1577) );
  XOR U1878 ( .A(n1293), .B(n1577), .Z(n4391) );
  XOR U1879 ( .A(in[1401]), .B(n4391), .Z(n5085) );
  NANDN U1880 ( .A(n5086), .B(n5085), .Z(n1056) );
  XNOR U1881 ( .A(n1683), .B(n1056), .Z(out[1045]) );
  XOR U1882 ( .A(n1058), .B(n1057), .Z(n2046) );
  XOR U1883 ( .A(in[553]), .B(n2046), .Z(n1687) );
  XOR U1884 ( .A(in[857]), .B(in[1177]), .Z(n1060) );
  XNOR U1885 ( .A(in[1497]), .B(in[217]), .Z(n1059) );
  XNOR U1886 ( .A(n1060), .B(n1059), .Z(n1061) );
  XOR U1887 ( .A(in[537]), .B(n1061), .Z(n1461) );
  XOR U1888 ( .A(in[153]), .B(n2817), .Z(n5089) );
  XOR U1889 ( .A(in[1337]), .B(in[57]), .Z(n1064) );
  XNOR U1890 ( .A(in[697]), .B(in[377]), .Z(n1063) );
  XNOR U1891 ( .A(n1064), .B(n1063), .Z(n1065) );
  XNOR U1892 ( .A(in[1017]), .B(n1065), .Z(n1581) );
  XOR U1893 ( .A(in[826]), .B(in[506]), .Z(n1067) );
  XNOR U1894 ( .A(in[1466]), .B(in[1146]), .Z(n1066) );
  XNOR U1895 ( .A(n1067), .B(n1066), .Z(n1068) );
  XNOR U1896 ( .A(in[186]), .B(n1068), .Z(n1305) );
  XOR U1897 ( .A(n1581), .B(n1305), .Z(n2116) );
  IV U1898 ( .A(n2116), .Z(n4394) );
  XNOR U1899 ( .A(in[1402]), .B(n4394), .Z(n5088) );
  NANDN U1900 ( .A(n5089), .B(n5088), .Z(n1069) );
  XNOR U1901 ( .A(n1687), .B(n1069), .Z(out[1046]) );
  XOR U1902 ( .A(n1071), .B(n1070), .Z(n2048) );
  XOR U1903 ( .A(in[554]), .B(n2048), .Z(n1691) );
  XOR U1904 ( .A(in[858]), .B(in[1178]), .Z(n1073) );
  XNOR U1905 ( .A(in[1498]), .B(in[218]), .Z(n1072) );
  XNOR U1906 ( .A(n1073), .B(n1072), .Z(n1074) );
  XOR U1907 ( .A(in[538]), .B(n1074), .Z(n1463) );
  XOR U1908 ( .A(in[154]), .B(n2840), .Z(n5092) );
  XOR U1909 ( .A(in[1338]), .B(in[58]), .Z(n1077) );
  XNOR U1910 ( .A(in[698]), .B(in[378]), .Z(n1076) );
  XNOR U1911 ( .A(n1077), .B(n1076), .Z(n1078) );
  XNOR U1912 ( .A(in[1018]), .B(n1078), .Z(n1585) );
  XOR U1913 ( .A(in[827]), .B(in[507]), .Z(n1080) );
  XNOR U1914 ( .A(in[1467]), .B(in[1147]), .Z(n1079) );
  XNOR U1915 ( .A(n1080), .B(n1079), .Z(n1081) );
  XNOR U1916 ( .A(in[187]), .B(n1081), .Z(n1309) );
  XOR U1917 ( .A(n1585), .B(n1309), .Z(n2118) );
  IV U1918 ( .A(n2118), .Z(n4397) );
  XNOR U1919 ( .A(in[1403]), .B(n4397), .Z(n5091) );
  NANDN U1920 ( .A(n5092), .B(n5091), .Z(n1082) );
  XNOR U1921 ( .A(n1691), .B(n1082), .Z(out[1047]) );
  XOR U1922 ( .A(in[1579]), .B(in[619]), .Z(n1084) );
  XNOR U1923 ( .A(in[939]), .B(in[299]), .Z(n1083) );
  XNOR U1924 ( .A(n1084), .B(n1083), .Z(n1085) );
  XNOR U1925 ( .A(in[1259]), .B(n1085), .Z(n1595) );
  XNOR U1926 ( .A(n1086), .B(n1595), .Z(n3430) );
  IV U1927 ( .A(n3430), .Z(n4090) );
  XOR U1928 ( .A(in[555]), .B(n4090), .Z(n1695) );
  XOR U1929 ( .A(in[859]), .B(in[1179]), .Z(n1088) );
  XNOR U1930 ( .A(in[1499]), .B(in[219]), .Z(n1087) );
  XNOR U1931 ( .A(n1088), .B(n1087), .Z(n1089) );
  XOR U1932 ( .A(in[539]), .B(n1089), .Z(n1467) );
  XOR U1933 ( .A(in[155]), .B(n2864), .Z(n5095) );
  XOR U1934 ( .A(in[828]), .B(in[508]), .Z(n1092) );
  XNOR U1935 ( .A(in[1468]), .B(in[1148]), .Z(n1091) );
  XNOR U1936 ( .A(n1092), .B(n1091), .Z(n1093) );
  XNOR U1937 ( .A(in[188]), .B(n1093), .Z(n1313) );
  XOR U1938 ( .A(n1094), .B(n1313), .Z(n4400) );
  XOR U1939 ( .A(in[1404]), .B(n4400), .Z(n5094) );
  NANDN U1940 ( .A(n5095), .B(n5094), .Z(n1095) );
  XNOR U1941 ( .A(n1695), .B(n1095), .Z(out[1048]) );
  XOR U1942 ( .A(in[1580]), .B(in[620]), .Z(n1097) );
  XNOR U1943 ( .A(in[940]), .B(in[300]), .Z(n1096) );
  XNOR U1944 ( .A(n1097), .B(n1096), .Z(n1098) );
  XNOR U1945 ( .A(in[1260]), .B(n1098), .Z(n1599) );
  XNOR U1946 ( .A(n1099), .B(n1599), .Z(n3433) );
  IV U1947 ( .A(n3433), .Z(n4094) );
  XOR U1948 ( .A(in[556]), .B(n4094), .Z(n1699) );
  XOR U1949 ( .A(in[860]), .B(in[1180]), .Z(n1101) );
  XNOR U1950 ( .A(in[1500]), .B(in[220]), .Z(n1100) );
  XNOR U1951 ( .A(n1101), .B(n1100), .Z(n1102) );
  XOR U1952 ( .A(in[540]), .B(n1102), .Z(n1473) );
  XOR U1953 ( .A(in[156]), .B(n2888), .Z(n5098) );
  XOR U1954 ( .A(n1105), .B(n1104), .Z(n4407) );
  XOR U1955 ( .A(in[1405]), .B(n4407), .Z(n5097) );
  NANDN U1956 ( .A(n5098), .B(n5097), .Z(n1106) );
  XNOR U1957 ( .A(n1699), .B(n1106), .Z(out[1049]) );
  XOR U1958 ( .A(in[1343]), .B(in[63]), .Z(n1108) );
  XNOR U1959 ( .A(in[703]), .B(in[383]), .Z(n1107) );
  XNOR U1960 ( .A(n1108), .B(n1107), .Z(n1109) );
  XNOR U1961 ( .A(in[1023]), .B(n1109), .Z(n1153) );
  XOR U1962 ( .A(n1110), .B(n1153), .Z(n3969) );
  XOR U1963 ( .A(in[639]), .B(n3969), .Z(n2712) );
  IV U1964 ( .A(n2712), .Z(n2801) );
  XNOR U1965 ( .A(in[230]), .B(n2037), .Z(n3192) );
  XOR U1966 ( .A(in[874]), .B(in[1194]), .Z(n1112) );
  XNOR U1967 ( .A(in[1514]), .B(in[234]), .Z(n1111) );
  XNOR U1968 ( .A(n1112), .B(n1111), .Z(n1113) );
  XNOR U1969 ( .A(in[554]), .B(n1113), .Z(n1523) );
  XNOR U1970 ( .A(n1114), .B(n1523), .Z(n4105) );
  IV U1971 ( .A(n4105), .Z(n1294) );
  XOR U1972 ( .A(in[1450]), .B(n1294), .Z(n3189) );
  NAND U1973 ( .A(n3192), .B(n3189), .Z(n1115) );
  XOR U1974 ( .A(n2801), .B(n1115), .Z(out[104]) );
  XOR U1975 ( .A(in[1581]), .B(in[621]), .Z(n1117) );
  XNOR U1976 ( .A(in[941]), .B(in[301]), .Z(n1116) );
  XNOR U1977 ( .A(n1117), .B(n1116), .Z(n1118) );
  XNOR U1978 ( .A(in[1261]), .B(n1118), .Z(n1603) );
  XNOR U1979 ( .A(n1119), .B(n1603), .Z(n3436) );
  IV U1980 ( .A(n3436), .Z(n4098) );
  XOR U1981 ( .A(in[557]), .B(n4098), .Z(n1703) );
  XOR U1982 ( .A(in[861]), .B(in[1181]), .Z(n1121) );
  XNOR U1983 ( .A(in[1501]), .B(in[221]), .Z(n1120) );
  XNOR U1984 ( .A(n1121), .B(n1120), .Z(n1122) );
  XOR U1985 ( .A(in[541]), .B(n1122), .Z(n1477) );
  XOR U1986 ( .A(in[157]), .B(n2921), .Z(n5101) );
  XOR U1987 ( .A(in[830]), .B(in[510]), .Z(n1125) );
  XNOR U1988 ( .A(in[1470]), .B(in[1150]), .Z(n1124) );
  XNOR U1989 ( .A(n1125), .B(n1124), .Z(n1126) );
  XNOR U1990 ( .A(in[190]), .B(n1126), .Z(n1317) );
  XOR U1991 ( .A(n1127), .B(n1317), .Z(n4410) );
  XOR U1992 ( .A(in[1406]), .B(n4410), .Z(n5100) );
  NANDN U1993 ( .A(n5101), .B(n5100), .Z(n1128) );
  XNOR U1994 ( .A(n1703), .B(n1128), .Z(out[1050]) );
  XOR U1995 ( .A(in[1582]), .B(in[622]), .Z(n1130) );
  XNOR U1996 ( .A(in[942]), .B(in[302]), .Z(n1129) );
  XNOR U1997 ( .A(n1130), .B(n1129), .Z(n1131) );
  XNOR U1998 ( .A(in[1262]), .B(n1131), .Z(n1607) );
  XNOR U1999 ( .A(n1132), .B(n1607), .Z(n3439) );
  IV U2000 ( .A(n3439), .Z(n4102) );
  XOR U2001 ( .A(in[558]), .B(n4102), .Z(n1707) );
  XOR U2002 ( .A(in[862]), .B(in[1182]), .Z(n1134) );
  XNOR U2003 ( .A(in[1502]), .B(in[222]), .Z(n1133) );
  XNOR U2004 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U2005 ( .A(in[542]), .B(n1135), .Z(n1481) );
  XNOR U2006 ( .A(in[158]), .B(n4054), .Z(n1457) );
  IV U2007 ( .A(n1457), .Z(n5104) );
  XOR U2008 ( .A(in[831]), .B(in[511]), .Z(n1138) );
  XNOR U2009 ( .A(in[1471]), .B(in[1151]), .Z(n1137) );
  XNOR U2010 ( .A(n1138), .B(n1137), .Z(n1139) );
  XNOR U2011 ( .A(in[191]), .B(n1139), .Z(n1321) );
  XOR U2012 ( .A(n1140), .B(n1321), .Z(n4413) );
  XOR U2013 ( .A(in[1407]), .B(n4413), .Z(n5103) );
  NANDN U2014 ( .A(n5104), .B(n5103), .Z(n1141) );
  XNOR U2015 ( .A(n1707), .B(n1141), .Z(out[1051]) );
  XOR U2016 ( .A(in[1583]), .B(in[623]), .Z(n1143) );
  XNOR U2017 ( .A(in[943]), .B(in[303]), .Z(n1142) );
  XNOR U2018 ( .A(n1143), .B(n1142), .Z(n1144) );
  XNOR U2019 ( .A(in[1263]), .B(n1144), .Z(n1611) );
  XNOR U2020 ( .A(n1145), .B(n1611), .Z(n3442) );
  IV U2021 ( .A(n3442), .Z(n4106) );
  XOR U2022 ( .A(in[559]), .B(n4106), .Z(n1712) );
  XOR U2023 ( .A(in[863]), .B(in[1183]), .Z(n1147) );
  XNOR U2024 ( .A(in[1503]), .B(in[223]), .Z(n1146) );
  XNOR U2025 ( .A(n1147), .B(n1146), .Z(n1148) );
  XOR U2026 ( .A(in[543]), .B(n1148), .Z(n1483) );
  XOR U2027 ( .A(in[159]), .B(n4058), .Z(n5108) );
  XOR U2028 ( .A(in[768]), .B(in[1088]), .Z(n1151) );
  XNOR U2029 ( .A(in[448]), .B(in[1408]), .Z(n1150) );
  XNOR U2030 ( .A(n1151), .B(n1150), .Z(n1152) );
  XNOR U2031 ( .A(in[128]), .B(n1152), .Z(n1328) );
  XOR U2032 ( .A(n1153), .B(n1328), .Z(n4416) );
  XOR U2033 ( .A(in[1344]), .B(n4416), .Z(n5105) );
  NANDN U2034 ( .A(n5108), .B(n5105), .Z(n1154) );
  XNOR U2035 ( .A(n1712), .B(n1154), .Z(out[1052]) );
  XOR U2036 ( .A(in[1584]), .B(in[624]), .Z(n1156) );
  XNOR U2037 ( .A(in[944]), .B(in[304]), .Z(n1155) );
  XNOR U2038 ( .A(n1156), .B(n1155), .Z(n1157) );
  XNOR U2039 ( .A(in[1264]), .B(n1157), .Z(n1615) );
  XNOR U2040 ( .A(n1158), .B(n1615), .Z(n3445) );
  IV U2041 ( .A(n3445), .Z(n4110) );
  XOR U2042 ( .A(in[560]), .B(n4110), .Z(n1716) );
  XOR U2043 ( .A(in[224]), .B(in[864]), .Z(n1160) );
  XNOR U2044 ( .A(in[1184]), .B(in[1504]), .Z(n1159) );
  XNOR U2045 ( .A(n1160), .B(n1159), .Z(n1161) );
  XOR U2046 ( .A(in[544]), .B(n1161), .Z(n1486) );
  XOR U2047 ( .A(in[160]), .B(n4062), .Z(n5111) );
  XOR U2048 ( .A(in[769]), .B(in[1089]), .Z(n1164) );
  XNOR U2049 ( .A(in[449]), .B(in[1409]), .Z(n1163) );
  XNOR U2050 ( .A(n1164), .B(n1163), .Z(n1165) );
  XNOR U2051 ( .A(in[129]), .B(n1165), .Z(n1332) );
  XOR U2052 ( .A(in[1280]), .B(in[640]), .Z(n1167) );
  XNOR U2053 ( .A(in[960]), .B(in[320]), .Z(n1166) );
  XNOR U2054 ( .A(n1167), .B(n1166), .Z(n1168) );
  XNOR U2055 ( .A(in[0]), .B(n1168), .Z(n1257) );
  XOR U2056 ( .A(n1332), .B(n1257), .Z(n4419) );
  XOR U2057 ( .A(in[1345]), .B(n4419), .Z(n5110) );
  NANDN U2058 ( .A(n5111), .B(n5110), .Z(n1169) );
  XNOR U2059 ( .A(n1716), .B(n1169), .Z(out[1053]) );
  XOR U2060 ( .A(in[1585]), .B(in[625]), .Z(n1171) );
  XNOR U2061 ( .A(in[945]), .B(in[305]), .Z(n1170) );
  XNOR U2062 ( .A(n1171), .B(n1170), .Z(n1172) );
  XNOR U2063 ( .A(in[1265]), .B(n1172), .Z(n1619) );
  XNOR U2064 ( .A(n1173), .B(n1619), .Z(n3448) );
  IV U2065 ( .A(n3448), .Z(n4118) );
  XOR U2066 ( .A(in[561]), .B(n4118), .Z(n1720) );
  XOR U2067 ( .A(in[225]), .B(in[865]), .Z(n1175) );
  XNOR U2068 ( .A(in[1185]), .B(in[1505]), .Z(n1174) );
  XNOR U2069 ( .A(n1175), .B(n1174), .Z(n1176) );
  XOR U2070 ( .A(n1177), .B(n233), .Z(n4066) );
  XNOR U2071 ( .A(in[161]), .B(n4066), .Z(n1465) );
  IV U2072 ( .A(n1465), .Z(n5118) );
  XOR U2073 ( .A(in[1]), .B(in[641]), .Z(n1179) );
  XNOR U2074 ( .A(in[961]), .B(in[321]), .Z(n1178) );
  XNOR U2075 ( .A(n1179), .B(n1178), .Z(n1180) );
  XNOR U2076 ( .A(in[1281]), .B(n1180), .Z(n1322) );
  XOR U2077 ( .A(in[1090]), .B(in[450]), .Z(n1182) );
  XNOR U2078 ( .A(in[130]), .B(in[770]), .Z(n1181) );
  XNOR U2079 ( .A(n1182), .B(n1181), .Z(n1183) );
  XNOR U2080 ( .A(in[1410]), .B(n1183), .Z(n1336) );
  XOR U2081 ( .A(n1322), .B(n1336), .Z(n4422) );
  XOR U2082 ( .A(in[1346]), .B(n4422), .Z(n5117) );
  NANDN U2083 ( .A(n5118), .B(n5117), .Z(n1184) );
  XNOR U2084 ( .A(n1720), .B(n1184), .Z(out[1054]) );
  XOR U2085 ( .A(in[1586]), .B(in[626]), .Z(n1186) );
  XNOR U2086 ( .A(in[946]), .B(in[306]), .Z(n1185) );
  XNOR U2087 ( .A(n1186), .B(n1185), .Z(n1187) );
  XNOR U2088 ( .A(in[1266]), .B(n1187), .Z(n1623) );
  XNOR U2089 ( .A(n1188), .B(n1623), .Z(n3451) );
  IV U2090 ( .A(n3451), .Z(n4122) );
  XOR U2091 ( .A(in[562]), .B(n4122), .Z(n1724) );
  XOR U2092 ( .A(in[1186]), .B(in[1506]), .Z(n1190) );
  XNOR U2093 ( .A(in[546]), .B(in[866]), .Z(n1189) );
  XNOR U2094 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U2095 ( .A(in[226]), .B(n1191), .Z(n1491) );
  XNOR U2096 ( .A(in[162]), .B(n4074), .Z(n1469) );
  IV U2097 ( .A(n1469), .Z(n5122) );
  XOR U2098 ( .A(in[2]), .B(in[642]), .Z(n1194) );
  XNOR U2099 ( .A(in[962]), .B(in[322]), .Z(n1193) );
  XNOR U2100 ( .A(n1194), .B(n1193), .Z(n1195) );
  XNOR U2101 ( .A(in[1282]), .B(n1195), .Z(n1367) );
  XOR U2102 ( .A(in[771]), .B(in[1091]), .Z(n1197) );
  XNOR U2103 ( .A(in[451]), .B(in[1411]), .Z(n1196) );
  XNOR U2104 ( .A(n1197), .B(n1196), .Z(n1198) );
  XNOR U2105 ( .A(in[131]), .B(n1198), .Z(n1340) );
  XOR U2106 ( .A(n1367), .B(n1340), .Z(n4425) );
  XOR U2107 ( .A(in[1347]), .B(n4425), .Z(n5119) );
  NANDN U2108 ( .A(n5122), .B(n5119), .Z(n1199) );
  XNOR U2109 ( .A(n1724), .B(n1199), .Z(out[1055]) );
  XOR U2110 ( .A(in[1587]), .B(in[627]), .Z(n1201) );
  XNOR U2111 ( .A(in[947]), .B(in[307]), .Z(n1200) );
  XNOR U2112 ( .A(n1201), .B(n1200), .Z(n1202) );
  XNOR U2113 ( .A(in[1267]), .B(n1202), .Z(n1628) );
  XNOR U2114 ( .A(n1203), .B(n1628), .Z(n3454) );
  IV U2115 ( .A(n3454), .Z(n4126) );
  XOR U2116 ( .A(in[563]), .B(n4126), .Z(n1728) );
  XOR U2117 ( .A(in[1187]), .B(in[1507]), .Z(n1205) );
  XNOR U2118 ( .A(in[547]), .B(in[867]), .Z(n1204) );
  XNOR U2119 ( .A(n1205), .B(n1204), .Z(n1206) );
  XOR U2120 ( .A(in[227]), .B(n1206), .Z(n1494) );
  XNOR U2121 ( .A(in[163]), .B(n4078), .Z(n1475) );
  IV U2122 ( .A(n1475), .Z(n5126) );
  XOR U2123 ( .A(in[772]), .B(in[1092]), .Z(n1209) );
  XNOR U2124 ( .A(in[452]), .B(in[1412]), .Z(n1208) );
  XNOR U2125 ( .A(n1209), .B(n1208), .Z(n1210) );
  XNOR U2126 ( .A(in[132]), .B(n1210), .Z(n1344) );
  XOR U2127 ( .A(in[323]), .B(in[643]), .Z(n1212) );
  XNOR U2128 ( .A(in[963]), .B(in[3]), .Z(n1211) );
  XNOR U2129 ( .A(n1212), .B(n1211), .Z(n1213) );
  XNOR U2130 ( .A(in[1283]), .B(n1213), .Z(n1408) );
  XOR U2131 ( .A(n1344), .B(n1408), .Z(n4428) );
  XOR U2132 ( .A(in[1348]), .B(n4428), .Z(n5123) );
  NANDN U2133 ( .A(n5126), .B(n5123), .Z(n1214) );
  XNOR U2134 ( .A(n1728), .B(n1214), .Z(out[1056]) );
  XOR U2135 ( .A(in[1588]), .B(in[628]), .Z(n1216) );
  XNOR U2136 ( .A(in[948]), .B(in[308]), .Z(n1215) );
  XNOR U2137 ( .A(n1216), .B(n1215), .Z(n1217) );
  XNOR U2138 ( .A(in[1268]), .B(n1217), .Z(n1632) );
  XNOR U2139 ( .A(n1218), .B(n1632), .Z(n3461) );
  IV U2140 ( .A(n3461), .Z(n4130) );
  XOR U2141 ( .A(in[564]), .B(n4130), .Z(n1732) );
  XOR U2142 ( .A(in[1188]), .B(in[1508]), .Z(n1220) );
  XNOR U2143 ( .A(in[548]), .B(in[868]), .Z(n1219) );
  XNOR U2144 ( .A(n1220), .B(n1219), .Z(n1221) );
  XNOR U2145 ( .A(in[228]), .B(n1221), .Z(n1497) );
  XNOR U2146 ( .A(in[164]), .B(n4082), .Z(n1479) );
  IV U2147 ( .A(n1479), .Z(n5130) );
  XOR U2148 ( .A(in[324]), .B(in[644]), .Z(n1224) );
  XNOR U2149 ( .A(in[964]), .B(in[4]), .Z(n1223) );
  XNOR U2150 ( .A(n1224), .B(n1223), .Z(n1225) );
  XNOR U2151 ( .A(in[1284]), .B(n1225), .Z(n1412) );
  XOR U2152 ( .A(in[773]), .B(in[1093]), .Z(n1227) );
  XNOR U2153 ( .A(in[453]), .B(in[1413]), .Z(n1226) );
  XNOR U2154 ( .A(n1227), .B(n1226), .Z(n1228) );
  XNOR U2155 ( .A(in[133]), .B(n1228), .Z(n1348) );
  XOR U2156 ( .A(n1412), .B(n1348), .Z(n4431) );
  XOR U2157 ( .A(in[1349]), .B(n4431), .Z(n5127) );
  NANDN U2158 ( .A(n5130), .B(n5127), .Z(n1229) );
  XNOR U2159 ( .A(n1732), .B(n1229), .Z(out[1057]) );
  XOR U2160 ( .A(in[1589]), .B(in[629]), .Z(n1231) );
  XNOR U2161 ( .A(in[949]), .B(in[309]), .Z(n1230) );
  XNOR U2162 ( .A(n1231), .B(n1230), .Z(n1232) );
  XNOR U2163 ( .A(in[1269]), .B(n1232), .Z(n1636) );
  XNOR U2164 ( .A(n1233), .B(n1636), .Z(n3464) );
  IV U2165 ( .A(n3464), .Z(n4134) );
  XOR U2166 ( .A(in[565]), .B(n4134), .Z(n1736) );
  XOR U2167 ( .A(in[1189]), .B(in[1509]), .Z(n1235) );
  XNOR U2168 ( .A(in[549]), .B(in[869]), .Z(n1234) );
  XNOR U2169 ( .A(n1235), .B(n1234), .Z(n1236) );
  XOR U2170 ( .A(in[229]), .B(n1236), .Z(n1501) );
  XOR U2171 ( .A(in[165]), .B(n2213), .Z(n5134) );
  XOR U2172 ( .A(in[774]), .B(in[1094]), .Z(n1239) );
  XNOR U2173 ( .A(in[454]), .B(in[1414]), .Z(n1238) );
  XNOR U2174 ( .A(n1239), .B(n1238), .Z(n1240) );
  XNOR U2175 ( .A(in[134]), .B(n1240), .Z(n1352) );
  XOR U2176 ( .A(in[325]), .B(in[645]), .Z(n1242) );
  XNOR U2177 ( .A(in[965]), .B(in[5]), .Z(n1241) );
  XNOR U2178 ( .A(n1242), .B(n1241), .Z(n1243) );
  XNOR U2179 ( .A(in[1285]), .B(n1243), .Z(n1414) );
  XOR U2180 ( .A(n1352), .B(n1414), .Z(n2128) );
  IV U2181 ( .A(n2128), .Z(n4434) );
  XNOR U2182 ( .A(in[1350]), .B(n4434), .Z(n5131) );
  NANDN U2183 ( .A(n5134), .B(n5131), .Z(n1244) );
  XNOR U2184 ( .A(n1736), .B(n1244), .Z(out[1058]) );
  XOR U2185 ( .A(in[1590]), .B(in[630]), .Z(n1246) );
  XNOR U2186 ( .A(in[950]), .B(in[310]), .Z(n1245) );
  XNOR U2187 ( .A(n1246), .B(n1245), .Z(n1247) );
  XNOR U2188 ( .A(in[1270]), .B(n1247), .Z(n1640) );
  XNOR U2189 ( .A(n1248), .B(n1640), .Z(n3260) );
  IV U2190 ( .A(n3260), .Z(n4138) );
  XOR U2191 ( .A(in[566]), .B(n4138), .Z(n1740) );
  XNOR U2192 ( .A(in[166]), .B(n1249), .Z(n5138) );
  XOR U2193 ( .A(in[775]), .B(in[1095]), .Z(n1251) );
  XNOR U2194 ( .A(in[455]), .B(in[1415]), .Z(n1250) );
  XNOR U2195 ( .A(n1251), .B(n1250), .Z(n1252) );
  XNOR U2196 ( .A(in[135]), .B(n1252), .Z(n1356) );
  XOR U2197 ( .A(in[326]), .B(in[6]), .Z(n1254) );
  XNOR U2198 ( .A(in[966]), .B(in[646]), .Z(n1253) );
  XNOR U2199 ( .A(n1254), .B(n1253), .Z(n1255) );
  XNOR U2200 ( .A(in[1286]), .B(n1255), .Z(n1416) );
  XOR U2201 ( .A(n1356), .B(n1416), .Z(n4445) );
  XOR U2202 ( .A(in[1351]), .B(n4445), .Z(n5135) );
  NAND U2203 ( .A(n5138), .B(n5135), .Z(n1256) );
  XNOR U2204 ( .A(n1740), .B(n1256), .Z(out[1059]) );
  XOR U2205 ( .A(n1258), .B(n1257), .Z(n3973) );
  XOR U2206 ( .A(in[576]), .B(n3973), .Z(n2714) );
  IV U2207 ( .A(n2714), .Z(n2803) );
  XNOR U2208 ( .A(in[1451]), .B(n4109), .Z(n3221) );
  XNOR U2209 ( .A(in[231]), .B(n2040), .Z(n3223) );
  NANDN U2210 ( .A(n3221), .B(n3223), .Z(n1259) );
  XOR U2211 ( .A(n2803), .B(n1259), .Z(out[105]) );
  XOR U2212 ( .A(in[1591]), .B(in[631]), .Z(n1261) );
  XNOR U2213 ( .A(in[951]), .B(in[311]), .Z(n1260) );
  XNOR U2214 ( .A(n1261), .B(n1260), .Z(n1262) );
  XNOR U2215 ( .A(in[1271]), .B(n1262), .Z(n1644) );
  XNOR U2216 ( .A(n1263), .B(n1644), .Z(n3263) );
  IV U2217 ( .A(n3263), .Z(n4142) );
  XOR U2218 ( .A(in[567]), .B(n4142), .Z(n1744) );
  XNOR U2219 ( .A(in[167]), .B(n1264), .Z(n5142) );
  XOR U2220 ( .A(in[776]), .B(in[1096]), .Z(n1266) );
  XNOR U2221 ( .A(in[456]), .B(in[1416]), .Z(n1265) );
  XNOR U2222 ( .A(n1266), .B(n1265), .Z(n1267) );
  XNOR U2223 ( .A(in[136]), .B(n1267), .Z(n1360) );
  XOR U2224 ( .A(in[327]), .B(in[7]), .Z(n1269) );
  XNOR U2225 ( .A(in[967]), .B(in[647]), .Z(n1268) );
  XNOR U2226 ( .A(n1269), .B(n1268), .Z(n1270) );
  XNOR U2227 ( .A(in[1287]), .B(n1270), .Z(n1418) );
  XOR U2228 ( .A(n1360), .B(n1418), .Z(n4448) );
  XOR U2229 ( .A(in[1352]), .B(n4448), .Z(n5139) );
  NAND U2230 ( .A(n5142), .B(n5139), .Z(n1271) );
  XNOR U2231 ( .A(n1744), .B(n1271), .Z(out[1060]) );
  XOR U2232 ( .A(in[632]), .B(in[1592]), .Z(n1273) );
  XNOR U2233 ( .A(in[1272]), .B(in[312]), .Z(n1272) );
  XNOR U2234 ( .A(n1273), .B(n1272), .Z(n1274) );
  XNOR U2235 ( .A(in[952]), .B(n1274), .Z(n1648) );
  XNOR U2236 ( .A(n1275), .B(n1648), .Z(n3270) );
  IV U2237 ( .A(n3270), .Z(n4146) );
  XOR U2238 ( .A(in[568]), .B(n4146), .Z(n1748) );
  XNOR U2239 ( .A(in[168]), .B(n1276), .Z(n5146) );
  XOR U2240 ( .A(in[1353]), .B(n4451), .Z(n5143) );
  NAND U2241 ( .A(n5146), .B(n5143), .Z(n1277) );
  XNOR U2242 ( .A(n1748), .B(n1277), .Z(out[1061]) );
  XOR U2243 ( .A(in[633]), .B(in[1593]), .Z(n1279) );
  XNOR U2244 ( .A(in[1273]), .B(in[313]), .Z(n1278) );
  XNOR U2245 ( .A(n1279), .B(n1278), .Z(n1280) );
  XNOR U2246 ( .A(in[953]), .B(n1280), .Z(n1652) );
  XNOR U2247 ( .A(n1281), .B(n1652), .Z(n3273) );
  IV U2248 ( .A(n3273), .Z(n4150) );
  XOR U2249 ( .A(in[569]), .B(n4150), .Z(n1753) );
  XOR U2250 ( .A(in[329]), .B(in[969]), .Z(n1283) );
  XNOR U2251 ( .A(in[9]), .B(in[649]), .Z(n1282) );
  XNOR U2252 ( .A(n1283), .B(n1282), .Z(n1284) );
  XNOR U2253 ( .A(in[1289]), .B(n1284), .Z(n1425) );
  XOR U2254 ( .A(in[778]), .B(in[1098]), .Z(n1286) );
  XNOR U2255 ( .A(in[458]), .B(in[1418]), .Z(n1285) );
  XNOR U2256 ( .A(n1286), .B(n1285), .Z(n1287) );
  XNOR U2257 ( .A(in[138]), .B(n1287), .Z(n1374) );
  XOR U2258 ( .A(n1425), .B(n1374), .Z(n4454) );
  XNOR U2259 ( .A(in[1354]), .B(n4454), .Z(n5148) );
  XNOR U2260 ( .A(in[169]), .B(n1288), .Z(n5150) );
  NANDN U2261 ( .A(n5148), .B(n5150), .Z(n1289) );
  XNOR U2262 ( .A(n1753), .B(n1289), .Z(out[1062]) );
  XOR U2263 ( .A(in[634]), .B(in[1594]), .Z(n1291) );
  XNOR U2264 ( .A(in[1274]), .B(in[314]), .Z(n1290) );
  XNOR U2265 ( .A(n1291), .B(n1290), .Z(n1292) );
  XNOR U2266 ( .A(in[954]), .B(n1292), .Z(n1656) );
  XNOR U2267 ( .A(n1293), .B(n1656), .Z(n3276) );
  IV U2268 ( .A(n3276), .Z(n4154) );
  XOR U2269 ( .A(in[570]), .B(n4154), .Z(n1757) );
  XNOR U2270 ( .A(in[170]), .B(n1294), .Z(n5154) );
  XOR U2271 ( .A(in[1419]), .B(in[779]), .Z(n1296) );
  XNOR U2272 ( .A(in[1099]), .B(in[459]), .Z(n1295) );
  XNOR U2273 ( .A(n1296), .B(n1295), .Z(n1297) );
  XNOR U2274 ( .A(in[139]), .B(n1297), .Z(n1380) );
  XOR U2275 ( .A(in[1290]), .B(in[650]), .Z(n1299) );
  XNOR U2276 ( .A(in[970]), .B(in[330]), .Z(n1298) );
  XNOR U2277 ( .A(n1299), .B(n1298), .Z(n1300) );
  XNOR U2278 ( .A(in[10]), .B(n1300), .Z(n1427) );
  XOR U2279 ( .A(n1380), .B(n1427), .Z(n4457) );
  XOR U2280 ( .A(in[1355]), .B(n4457), .Z(n5151) );
  NAND U2281 ( .A(n5154), .B(n5151), .Z(n1301) );
  XNOR U2282 ( .A(n1757), .B(n1301), .Z(out[1063]) );
  XOR U2283 ( .A(in[955]), .B(in[1275]), .Z(n1303) );
  XNOR U2284 ( .A(in[1595]), .B(in[315]), .Z(n1302) );
  XNOR U2285 ( .A(n1303), .B(n1302), .Z(n1304) );
  XOR U2286 ( .A(in[635]), .B(n1304), .Z(n1660) );
  XOR U2287 ( .A(n1305), .B(n1660), .Z(n4164) );
  XOR U2288 ( .A(in[571]), .B(n4164), .Z(n1759) );
  XOR U2289 ( .A(in[956]), .B(in[1276]), .Z(n1307) );
  XNOR U2290 ( .A(in[1596]), .B(in[316]), .Z(n1306) );
  XNOR U2291 ( .A(n1307), .B(n1306), .Z(n1308) );
  XOR U2292 ( .A(in[636]), .B(n1308), .Z(n1664) );
  XOR U2293 ( .A(n1309), .B(n1664), .Z(n4168) );
  XOR U2294 ( .A(in[572]), .B(n4168), .Z(n1761) );
  XOR U2295 ( .A(in[957]), .B(in[1277]), .Z(n1311) );
  XNOR U2296 ( .A(in[1597]), .B(in[317]), .Z(n1310) );
  XNOR U2297 ( .A(n1311), .B(n1310), .Z(n1312) );
  XOR U2298 ( .A(in[637]), .B(n1312), .Z(n1669) );
  XOR U2299 ( .A(n1313), .B(n1669), .Z(n4172) );
  XOR U2300 ( .A(in[573]), .B(n4172), .Z(n1763) );
  IV U2301 ( .A(n3288), .Z(n4176) );
  XOR U2302 ( .A(in[574]), .B(n4176), .Z(n1765) );
  XOR U2303 ( .A(in[959]), .B(in[1279]), .Z(n1315) );
  XNOR U2304 ( .A(in[1599]), .B(in[319]), .Z(n1314) );
  XNOR U2305 ( .A(n1315), .B(n1314), .Z(n1316) );
  XOR U2306 ( .A(in[639]), .B(n1316), .Z(n1677) );
  XOR U2307 ( .A(n1317), .B(n1677), .Z(n3291) );
  XOR U2308 ( .A(in[575]), .B(n3291), .Z(n1766) );
  XOR U2309 ( .A(in[896]), .B(in[1216]), .Z(n1319) );
  XNOR U2310 ( .A(in[1536]), .B(in[256]), .Z(n1318) );
  XNOR U2311 ( .A(n1319), .B(n1318), .Z(n1320) );
  XOR U2312 ( .A(in[576]), .B(n1320), .Z(n1681) );
  XOR U2313 ( .A(n1321), .B(n1681), .Z(n3294) );
  XOR U2314 ( .A(in[512]), .B(n3294), .Z(n1768) );
  XOR U2315 ( .A(n1323), .B(n1322), .Z(n3977) );
  XOR U2316 ( .A(in[577]), .B(n3977), .Z(n2717) );
  IV U2317 ( .A(n2717), .Z(n2805) );
  XNOR U2318 ( .A(in[1452]), .B(n4117), .Z(n3245) );
  XNOR U2319 ( .A(in[232]), .B(n2044), .Z(n3247) );
  NANDN U2320 ( .A(n3245), .B(n3247), .Z(n1324) );
  XOR U2321 ( .A(n2805), .B(n1324), .Z(out[106]) );
  XOR U2322 ( .A(in[897]), .B(in[1217]), .Z(n1326) );
  XNOR U2323 ( .A(in[1537]), .B(in[257]), .Z(n1325) );
  XNOR U2324 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U2325 ( .A(in[577]), .B(n1327), .Z(n1685) );
  XOR U2326 ( .A(n1328), .B(n1685), .Z(n3297) );
  XOR U2327 ( .A(in[513]), .B(n3297), .Z(n1770) );
  XOR U2328 ( .A(in[1538]), .B(in[578]), .Z(n1330) );
  XNOR U2329 ( .A(in[898]), .B(in[258]), .Z(n1329) );
  XNOR U2330 ( .A(n1330), .B(n1329), .Z(n1331) );
  XOR U2331 ( .A(in[1218]), .B(n1331), .Z(n1689) );
  XOR U2332 ( .A(n1332), .B(n1689), .Z(n3304) );
  XOR U2333 ( .A(in[514]), .B(n3304), .Z(n1772) );
  XOR U2334 ( .A(in[1539]), .B(in[579]), .Z(n1334) );
  XNOR U2335 ( .A(in[899]), .B(in[259]), .Z(n1333) );
  XNOR U2336 ( .A(n1334), .B(n1333), .Z(n1335) );
  XOR U2337 ( .A(in[1219]), .B(n1335), .Z(n1693) );
  XOR U2338 ( .A(n1336), .B(n1693), .Z(n3307) );
  XOR U2339 ( .A(in[515]), .B(n3307), .Z(n1776) );
  XOR U2340 ( .A(in[1540]), .B(in[580]), .Z(n1338) );
  XNOR U2341 ( .A(in[900]), .B(in[260]), .Z(n1337) );
  XNOR U2342 ( .A(n1338), .B(n1337), .Z(n1339) );
  XOR U2343 ( .A(in[1220]), .B(n1339), .Z(n1697) );
  XOR U2344 ( .A(n1340), .B(n1697), .Z(n3310) );
  XOR U2345 ( .A(in[516]), .B(n3310), .Z(n1778) );
  XOR U2346 ( .A(in[1541]), .B(in[581]), .Z(n1342) );
  XNOR U2347 ( .A(in[901]), .B(in[261]), .Z(n1341) );
  XNOR U2348 ( .A(n1342), .B(n1341), .Z(n1343) );
  XOR U2349 ( .A(in[1221]), .B(n1343), .Z(n1701) );
  XOR U2350 ( .A(n1344), .B(n1701), .Z(n3313) );
  XOR U2351 ( .A(in[517]), .B(n3313), .Z(n1780) );
  XOR U2352 ( .A(in[1542]), .B(in[582]), .Z(n1346) );
  XNOR U2353 ( .A(in[902]), .B(in[262]), .Z(n1345) );
  XNOR U2354 ( .A(n1346), .B(n1345), .Z(n1347) );
  XOR U2355 ( .A(in[1222]), .B(n1347), .Z(n1705) );
  XOR U2356 ( .A(n1348), .B(n1705), .Z(n3316) );
  XOR U2357 ( .A(in[518]), .B(n3316), .Z(n1782) );
  XOR U2358 ( .A(in[1543]), .B(in[583]), .Z(n1350) );
  XNOR U2359 ( .A(in[903]), .B(in[263]), .Z(n1349) );
  XNOR U2360 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U2361 ( .A(in[1223]), .B(n1351), .Z(n1710) );
  IV U2362 ( .A(n3931), .Z(n3319) );
  XOR U2363 ( .A(in[519]), .B(n3319), .Z(n1784) );
  XOR U2364 ( .A(in[1544]), .B(in[584]), .Z(n1354) );
  XNOR U2365 ( .A(in[904]), .B(in[264]), .Z(n1353) );
  XNOR U2366 ( .A(n1354), .B(n1353), .Z(n1355) );
  XOR U2367 ( .A(in[1224]), .B(n1355), .Z(n1714) );
  XOR U2368 ( .A(n1356), .B(n1714), .Z(n3935) );
  XOR U2369 ( .A(in[520]), .B(n3935), .Z(n1786) );
  XOR U2370 ( .A(in[1545]), .B(in[585]), .Z(n1358) );
  XNOR U2371 ( .A(in[905]), .B(in[265]), .Z(n1357) );
  XNOR U2372 ( .A(n1358), .B(n1357), .Z(n1359) );
  XOR U2373 ( .A(in[1225]), .B(n1359), .Z(n1718) );
  XOR U2374 ( .A(n1360), .B(n1718), .Z(n3942) );
  XOR U2375 ( .A(in[521]), .B(n3942), .Z(n1788) );
  XOR U2376 ( .A(in[1546]), .B(in[586]), .Z(n1362) );
  XNOR U2377 ( .A(in[906]), .B(in[266]), .Z(n1361) );
  XNOR U2378 ( .A(n1362), .B(n1361), .Z(n1363) );
  XOR U2379 ( .A(in[1226]), .B(n1363), .Z(n1722) );
  XOR U2380 ( .A(n1364), .B(n1722), .Z(n3946) );
  XOR U2381 ( .A(in[522]), .B(n3946), .Z(n1790) );
  NOR U2382 ( .A(n1365), .B(n1563), .Z(n1366) );
  XNOR U2383 ( .A(n1790), .B(n1366), .Z(out[1079]) );
  XOR U2384 ( .A(n1368), .B(n1367), .Z(n3984) );
  XOR U2385 ( .A(in[578]), .B(n3984), .Z(n2719) );
  IV U2386 ( .A(n2719), .Z(n2807) );
  IV U2387 ( .A(n1369), .Z(n4121) );
  XOR U2388 ( .A(in[1453]), .B(n4121), .Z(n3257) );
  XNOR U2389 ( .A(in[233]), .B(n2046), .Z(n3259) );
  NANDN U2390 ( .A(n3257), .B(n3259), .Z(n1370) );
  XOR U2391 ( .A(n2807), .B(n1370), .Z(out[107]) );
  XOR U2392 ( .A(in[1547]), .B(in[587]), .Z(n1372) );
  XNOR U2393 ( .A(in[907]), .B(in[267]), .Z(n1371) );
  XNOR U2394 ( .A(n1372), .B(n1371), .Z(n1373) );
  XOR U2395 ( .A(in[1227]), .B(n1373), .Z(n1726) );
  XOR U2396 ( .A(n1374), .B(n1726), .Z(n3950) );
  XOR U2397 ( .A(in[523]), .B(n3950), .Z(n1792) );
  NOR U2398 ( .A(n1375), .B(n1567), .Z(n1376) );
  XNOR U2399 ( .A(n1792), .B(n1376), .Z(out[1080]) );
  XOR U2400 ( .A(in[1548]), .B(in[588]), .Z(n1378) );
  XNOR U2401 ( .A(in[908]), .B(in[268]), .Z(n1377) );
  XNOR U2402 ( .A(n1378), .B(n1377), .Z(n1379) );
  XOR U2403 ( .A(in[1228]), .B(n1379), .Z(n1730) );
  XOR U2404 ( .A(n1380), .B(n1730), .Z(n3954) );
  XOR U2405 ( .A(in[524]), .B(n3954), .Z(n1794) );
  NOR U2406 ( .A(n1381), .B(n1571), .Z(n1382) );
  XNOR U2407 ( .A(n1794), .B(n1382), .Z(out[1081]) );
  XOR U2408 ( .A(in[1549]), .B(in[589]), .Z(n1384) );
  XNOR U2409 ( .A(in[909]), .B(in[269]), .Z(n1383) );
  XNOR U2410 ( .A(n1384), .B(n1383), .Z(n1385) );
  XNOR U2411 ( .A(in[1229]), .B(n1385), .Z(n1734) );
  XOR U2412 ( .A(n1734), .B(n1386), .Z(n3958) );
  XOR U2413 ( .A(in[525]), .B(n3958), .Z(n1798) );
  XOR U2414 ( .A(in[1550]), .B(in[590]), .Z(n1388) );
  XNOR U2415 ( .A(in[910]), .B(in[270]), .Z(n1387) );
  XNOR U2416 ( .A(n1388), .B(n1387), .Z(n1389) );
  XNOR U2417 ( .A(in[1230]), .B(n1389), .Z(n1738) );
  XOR U2418 ( .A(n1738), .B(n1390), .Z(n3962) );
  XOR U2419 ( .A(in[526]), .B(n3962), .Z(n1800) );
  XOR U2420 ( .A(in[1551]), .B(in[591]), .Z(n1392) );
  XNOR U2421 ( .A(in[911]), .B(in[271]), .Z(n1391) );
  XNOR U2422 ( .A(n1392), .B(n1391), .Z(n1393) );
  XNOR U2423 ( .A(in[1231]), .B(n1393), .Z(n1742) );
  XOR U2424 ( .A(n1742), .B(n1394), .Z(n3966) );
  XOR U2425 ( .A(in[527]), .B(n3966), .Z(n1802) );
  XOR U2426 ( .A(in[1552]), .B(in[592]), .Z(n1396) );
  XNOR U2427 ( .A(in[912]), .B(in[272]), .Z(n1395) );
  XNOR U2428 ( .A(n1396), .B(n1395), .Z(n1397) );
  XNOR U2429 ( .A(in[1232]), .B(n1397), .Z(n1746) );
  XOR U2430 ( .A(n1746), .B(n1398), .Z(n3970) );
  XOR U2431 ( .A(in[528]), .B(n3970), .Z(n1804) );
  XOR U2432 ( .A(in[1553]), .B(in[593]), .Z(n1400) );
  XNOR U2433 ( .A(in[913]), .B(in[273]), .Z(n1399) );
  XNOR U2434 ( .A(n1400), .B(n1399), .Z(n1401) );
  XOR U2435 ( .A(in[1233]), .B(n1401), .Z(n1751) );
  XOR U2436 ( .A(n1402), .B(n1751), .Z(n3974) );
  XOR U2437 ( .A(in[529]), .B(n3974), .Z(n1806) );
  XOR U2438 ( .A(in[1554]), .B(in[594]), .Z(n1404) );
  XNOR U2439 ( .A(in[914]), .B(in[274]), .Z(n1403) );
  XNOR U2440 ( .A(n1404), .B(n1403), .Z(n1405) );
  XOR U2441 ( .A(in[1234]), .B(n1405), .Z(n1755) );
  XOR U2442 ( .A(n1406), .B(n1755), .Z(n3978) );
  XOR U2443 ( .A(in[530]), .B(n3978), .Z(n1808) );
  XNOR U2444 ( .A(in[957]), .B(n3961), .Z(n1811) );
  XNOR U2445 ( .A(in[958]), .B(n3965), .Z(n1814) );
  XNOR U2446 ( .A(n1408), .B(n1407), .Z(n3988) );
  XOR U2447 ( .A(in[579]), .B(n3988), .Z(n2721) );
  IV U2448 ( .A(n2721), .Z(n2809) );
  IV U2449 ( .A(n1409), .Z(n4125) );
  XOR U2450 ( .A(in[1454]), .B(n4125), .Z(n3267) );
  XNOR U2451 ( .A(in[234]), .B(n2048), .Z(n3269) );
  NANDN U2452 ( .A(n3267), .B(n3269), .Z(n1410) );
  XOR U2453 ( .A(n2809), .B(n1410), .Z(out[108]) );
  XNOR U2454 ( .A(in[959]), .B(n3969), .Z(n1817) );
  XNOR U2455 ( .A(in[896]), .B(n3973), .Z(n1820) );
  XNOR U2456 ( .A(in[897]), .B(n3977), .Z(n1825) );
  XNOR U2457 ( .A(in[898]), .B(n3984), .Z(n1828) );
  XNOR U2458 ( .A(in[899]), .B(n3988), .Z(n1830) );
  XOR U2459 ( .A(n1412), .B(n1411), .Z(n2011) );
  XOR U2460 ( .A(in[900]), .B(n2011), .Z(n1831) );
  XOR U2461 ( .A(n1414), .B(n1413), .Z(n2013) );
  XOR U2462 ( .A(in[901]), .B(n2013), .Z(n1833) );
  XOR U2463 ( .A(n1416), .B(n1415), .Z(n2016) );
  XOR U2464 ( .A(in[902]), .B(n2016), .Z(n1835) );
  XOR U2465 ( .A(n1418), .B(n1417), .Z(n2019) );
  XOR U2466 ( .A(in[903]), .B(n2019), .Z(n1837) );
  XOR U2467 ( .A(n1420), .B(n1419), .Z(n2021) );
  XOR U2468 ( .A(in[904]), .B(n2021), .Z(n1839) );
  IV U2469 ( .A(n2011), .Z(n3992) );
  XOR U2470 ( .A(in[580]), .B(n3992), .Z(n2811) );
  IV U2471 ( .A(n1421), .Z(n4129) );
  XOR U2472 ( .A(in[1455]), .B(n4129), .Z(n3301) );
  XNOR U2473 ( .A(in[235]), .B(n4090), .Z(n3303) );
  NANDN U2474 ( .A(n3301), .B(n3303), .Z(n1422) );
  XNOR U2475 ( .A(n2811), .B(n1422), .Z(out[109]) );
  XNOR U2476 ( .A(in[200]), .B(n3935), .Z(n4282) );
  XOR U2477 ( .A(in[1420]), .B(n3194), .Z(n4283) );
  XNOR U2478 ( .A(n4485), .B(in[1043]), .Z(n2879) );
  NANDN U2479 ( .A(n4283), .B(n2879), .Z(n1423) );
  XNOR U2480 ( .A(n4282), .B(n1423), .Z(out[10]) );
  XOR U2481 ( .A(n1425), .B(n1424), .Z(n2023) );
  XOR U2482 ( .A(in[905]), .B(n2023), .Z(n1841) );
  XOR U2483 ( .A(n1427), .B(n1426), .Z(n2026) );
  XOR U2484 ( .A(in[906]), .B(n2026), .Z(n1843) );
  XOR U2485 ( .A(n1429), .B(n1428), .Z(n2028) );
  XOR U2486 ( .A(in[907]), .B(n2028), .Z(n1847) );
  XOR U2487 ( .A(n1431), .B(n1430), .Z(n2030) );
  XOR U2488 ( .A(in[908]), .B(n2030), .Z(n1849) );
  XOR U2489 ( .A(n1433), .B(n1432), .Z(n3110) );
  XOR U2490 ( .A(in[909]), .B(n3110), .Z(n1851) );
  XOR U2491 ( .A(n1435), .B(n1434), .Z(n3116) );
  XOR U2492 ( .A(in[910]), .B(n3116), .Z(n1853) );
  XNOR U2493 ( .A(n1437), .B(n1436), .Z(n3118) );
  XOR U2494 ( .A(in[911]), .B(n3118), .Z(n1855) );
  XNOR U2495 ( .A(n1439), .B(n1438), .Z(n3120) );
  XOR U2496 ( .A(in[912]), .B(n3120), .Z(n1857) );
  XOR U2497 ( .A(n1440), .B(n232), .Z(n4048) );
  XOR U2498 ( .A(in[913]), .B(n4048), .Z(n1859) );
  XOR U2499 ( .A(n1442), .B(n1441), .Z(n2038) );
  XOR U2500 ( .A(in[914]), .B(n2038), .Z(n1861) );
  IV U2501 ( .A(n2013), .Z(n3996) );
  XOR U2502 ( .A(in[581]), .B(n3996), .Z(n2813) );
  IV U2503 ( .A(n1443), .Z(n4133) );
  XOR U2504 ( .A(in[1456]), .B(n4133), .Z(n3331) );
  XNOR U2505 ( .A(in[236]), .B(n4094), .Z(n3333) );
  NANDN U2506 ( .A(n3331), .B(n3333), .Z(n1444) );
  XNOR U2507 ( .A(n2813), .B(n1444), .Z(out[110]) );
  XNOR U2508 ( .A(n1446), .B(n1445), .Z(n3124) );
  XOR U2509 ( .A(in[915]), .B(n3124), .Z(n1863) );
  XNOR U2510 ( .A(n1448), .B(n1447), .Z(n3126) );
  XOR U2511 ( .A(in[916]), .B(n3126), .Z(n1865) );
  XOR U2512 ( .A(n1450), .B(n1449), .Z(n3128) );
  XOR U2513 ( .A(in[917]), .B(n3128), .Z(n1869) );
  XOR U2514 ( .A(n1452), .B(n1451), .Z(n3130) );
  XOR U2515 ( .A(in[918]), .B(n3130), .Z(n1871) );
  XOR U2516 ( .A(n1454), .B(n1453), .Z(n3132) );
  XOR U2517 ( .A(in[919]), .B(n3132), .Z(n1873) );
  XNOR U2518 ( .A(n1456), .B(n1455), .Z(n3138) );
  XOR U2519 ( .A(in[920]), .B(n3138), .Z(n1875) );
  NOR U2520 ( .A(n1457), .B(n1707), .Z(n1458) );
  XNOR U2521 ( .A(n1875), .B(n1458), .Z(out[1115]) );
  XNOR U2522 ( .A(n1460), .B(n1459), .Z(n3140) );
  XOR U2523 ( .A(in[921]), .B(n3140), .Z(n1877) );
  XNOR U2524 ( .A(n1462), .B(n1461), .Z(n3143) );
  XOR U2525 ( .A(in[922]), .B(n3143), .Z(n1879) );
  XNOR U2526 ( .A(n1464), .B(n1463), .Z(n3145) );
  XOR U2527 ( .A(in[923]), .B(n3145), .Z(n1881) );
  NOR U2528 ( .A(n1465), .B(n1720), .Z(n1466) );
  XNOR U2529 ( .A(n1881), .B(n1466), .Z(out[1118]) );
  XNOR U2530 ( .A(n1468), .B(n1467), .Z(n3024) );
  XOR U2531 ( .A(in[924]), .B(n3024), .Z(n1883) );
  NOR U2532 ( .A(n1469), .B(n1724), .Z(n1470) );
  XNOR U2533 ( .A(n1883), .B(n1470), .Z(out[1119]) );
  IV U2534 ( .A(n2016), .Z(n4000) );
  XOR U2535 ( .A(in[582]), .B(n4000), .Z(n2815) );
  IV U2536 ( .A(n1471), .Z(n4137) );
  XOR U2537 ( .A(in[1457]), .B(n4137), .Z(n3360) );
  XNOR U2538 ( .A(in[237]), .B(n4098), .Z(n3362) );
  NANDN U2539 ( .A(n3360), .B(n3362), .Z(n1472) );
  XNOR U2540 ( .A(n2815), .B(n1472), .Z(out[111]) );
  XNOR U2541 ( .A(n1474), .B(n1473), .Z(n3026) );
  XOR U2542 ( .A(in[925]), .B(n3026), .Z(n1885) );
  NOR U2543 ( .A(n1475), .B(n1728), .Z(n1476) );
  XNOR U2544 ( .A(n1885), .B(n1476), .Z(out[1120]) );
  XNOR U2545 ( .A(n1478), .B(n1477), .Z(n3028) );
  XOR U2546 ( .A(in[926]), .B(n3028), .Z(n1887) );
  NOR U2547 ( .A(n1479), .B(n1732), .Z(n1480) );
  XNOR U2548 ( .A(n1887), .B(n1480), .Z(out[1121]) );
  XNOR U2549 ( .A(n1482), .B(n1481), .Z(n3030) );
  XOR U2550 ( .A(in[927]), .B(n3030), .Z(n1891) );
  XNOR U2551 ( .A(n1484), .B(n1483), .Z(n3032) );
  XOR U2552 ( .A(in[928]), .B(n3032), .Z(n1893) );
  NOR U2553 ( .A(n5138), .B(n1740), .Z(n1485) );
  XNOR U2554 ( .A(n1893), .B(n1485), .Z(out[1123]) );
  XOR U2555 ( .A(n1487), .B(n1486), .Z(n3034) );
  XOR U2556 ( .A(in[929]), .B(n3034), .Z(n1895) );
  NOR U2557 ( .A(n5142), .B(n1744), .Z(n1488) );
  XNOR U2558 ( .A(n1895), .B(n1488), .Z(out[1124]) );
  XOR U2559 ( .A(n1489), .B(n233), .Z(n4124) );
  XOR U2560 ( .A(in[930]), .B(n4124), .Z(n1897) );
  NOR U2561 ( .A(n5146), .B(n1748), .Z(n1490) );
  XNOR U2562 ( .A(n1897), .B(n1490), .Z(out[1125]) );
  XOR U2563 ( .A(n1492), .B(n1491), .Z(n3037) );
  XOR U2564 ( .A(in[931]), .B(n3037), .Z(n1899) );
  NOR U2565 ( .A(n5150), .B(n1753), .Z(n1493) );
  XNOR U2566 ( .A(n1899), .B(n1493), .Z(out[1126]) );
  XOR U2567 ( .A(n1495), .B(n1494), .Z(n3039) );
  XOR U2568 ( .A(in[932]), .B(n3039), .Z(n1901) );
  NOR U2569 ( .A(n5154), .B(n1757), .Z(n1496) );
  XNOR U2570 ( .A(n1901), .B(n1496), .Z(out[1127]) );
  XOR U2571 ( .A(n1498), .B(n1497), .Z(n4136) );
  XOR U2572 ( .A(in[933]), .B(n4136), .Z(n1904) );
  NAND U2573 ( .A(n1499), .B(n1759), .Z(n1500) );
  XNOR U2574 ( .A(n1904), .B(n1500), .Z(out[1128]) );
  XNOR U2575 ( .A(n1502), .B(n1501), .Z(n4140) );
  XOR U2576 ( .A(in[934]), .B(n4140), .Z(n1908) );
  NAND U2577 ( .A(n1503), .B(n1761), .Z(n1504) );
  XNOR U2578 ( .A(n1908), .B(n1504), .Z(out[1129]) );
  IV U2579 ( .A(n2019), .Z(n4004) );
  XOR U2580 ( .A(in[583]), .B(n4004), .Z(n2820) );
  IV U2581 ( .A(n1505), .Z(n4141) );
  XOR U2582 ( .A(in[1458]), .B(n4141), .Z(n3388) );
  XNOR U2583 ( .A(in[238]), .B(n4102), .Z(n3390) );
  NANDN U2584 ( .A(n3388), .B(n3390), .Z(n1506) );
  XNOR U2585 ( .A(n2820), .B(n1506), .Z(out[112]) );
  XOR U2586 ( .A(n1508), .B(n1507), .Z(n4144) );
  XOR U2587 ( .A(in[935]), .B(n4144), .Z(n1912) );
  NAND U2588 ( .A(n1509), .B(n1763), .Z(n1510) );
  XNOR U2589 ( .A(n1912), .B(n1510), .Z(out[1130]) );
  XOR U2590 ( .A(n1512), .B(n1511), .Z(n4148) );
  XOR U2591 ( .A(in[936]), .B(n4148), .Z(n1916) );
  NANDN U2592 ( .A(n1765), .B(n1513), .Z(n1514) );
  XNOR U2593 ( .A(n1916), .B(n1514), .Z(out[1131]) );
  XOR U2594 ( .A(n1516), .B(n1515), .Z(n4152) );
  XOR U2595 ( .A(in[937]), .B(n4152), .Z(n1922) );
  NAND U2596 ( .A(n1517), .B(n1766), .Z(n1518) );
  XNOR U2597 ( .A(n1922), .B(n1518), .Z(out[1132]) );
  XOR U2598 ( .A(n1520), .B(n1519), .Z(n4162) );
  XOR U2599 ( .A(in[938]), .B(n4162), .Z(n1926) );
  NAND U2600 ( .A(n1521), .B(n1768), .Z(n1522) );
  XNOR U2601 ( .A(n1926), .B(n1522), .Z(out[1133]) );
  XOR U2602 ( .A(n1524), .B(n1523), .Z(n4166) );
  XOR U2603 ( .A(in[939]), .B(n4166), .Z(n1930) );
  NAND U2604 ( .A(n1525), .B(n1770), .Z(n1526) );
  XNOR U2605 ( .A(n1930), .B(n1526), .Z(out[1134]) );
  XOR U2606 ( .A(n1528), .B(n1527), .Z(n4170) );
  XOR U2607 ( .A(in[940]), .B(n4170), .Z(n1934) );
  NAND U2608 ( .A(n1529), .B(n1772), .Z(n1530) );
  XNOR U2609 ( .A(n1934), .B(n1530), .Z(out[1135]) );
  XOR U2610 ( .A(n1532), .B(n1531), .Z(n4174) );
  XOR U2611 ( .A(in[941]), .B(n4174), .Z(n1938) );
  NAND U2612 ( .A(n1533), .B(n1776), .Z(n1534) );
  XNOR U2613 ( .A(n1938), .B(n1534), .Z(out[1136]) );
  XOR U2614 ( .A(n1536), .B(n1535), .Z(n3898) );
  XOR U2615 ( .A(in[942]), .B(n3898), .Z(n1942) );
  NAND U2616 ( .A(n1537), .B(n1778), .Z(n1538) );
  XNOR U2617 ( .A(n1942), .B(n1538), .Z(out[1137]) );
  XOR U2618 ( .A(n1540), .B(n1539), .Z(n3902) );
  XOR U2619 ( .A(in[943]), .B(n3902), .Z(n1946) );
  NAND U2620 ( .A(n1541), .B(n1780), .Z(n1542) );
  XNOR U2621 ( .A(n1946), .B(n1542), .Z(out[1138]) );
  XOR U2622 ( .A(n1544), .B(n1543), .Z(n3906) );
  XOR U2623 ( .A(in[944]), .B(n3906), .Z(n1950) );
  NAND U2624 ( .A(n1545), .B(n1782), .Z(n1546) );
  XNOR U2625 ( .A(n1950), .B(n1546), .Z(out[1139]) );
  IV U2626 ( .A(n2021), .Z(n4008) );
  XOR U2627 ( .A(in[584]), .B(n4008), .Z(n2822) );
  IV U2628 ( .A(n1547), .Z(n4145) );
  XOR U2629 ( .A(in[1459]), .B(n4145), .Z(n3423) );
  XNOR U2630 ( .A(in[239]), .B(n4106), .Z(n3425) );
  NANDN U2631 ( .A(n3423), .B(n3425), .Z(n1548) );
  XNOR U2632 ( .A(n2822), .B(n1548), .Z(out[113]) );
  XOR U2633 ( .A(n1550), .B(n1549), .Z(n3910) );
  XOR U2634 ( .A(in[945]), .B(n3910), .Z(n1954) );
  NAND U2635 ( .A(n1551), .B(n1784), .Z(n1552) );
  XNOR U2636 ( .A(n1954), .B(n1552), .Z(out[1140]) );
  XOR U2637 ( .A(n1554), .B(n1553), .Z(n3914) );
  XOR U2638 ( .A(in[946]), .B(n3914), .Z(n1958) );
  NAND U2639 ( .A(n1555), .B(n1786), .Z(n1556) );
  XNOR U2640 ( .A(n1958), .B(n1556), .Z(out[1141]) );
  XNOR U2641 ( .A(n1558), .B(n1557), .Z(n3918) );
  IV U2642 ( .A(n3918), .Z(n2569) );
  XOR U2643 ( .A(in[947]), .B(n2569), .Z(n1964) );
  NAND U2644 ( .A(n1559), .B(n1788), .Z(n1560) );
  XNOR U2645 ( .A(n1964), .B(n1560), .Z(out[1142]) );
  XNOR U2646 ( .A(n1562), .B(n1561), .Z(n3922) );
  IV U2647 ( .A(n3922), .Z(n2611) );
  XOR U2648 ( .A(in[948]), .B(n2611), .Z(n1968) );
  NAND U2649 ( .A(n1563), .B(n1790), .Z(n1564) );
  XNOR U2650 ( .A(n1968), .B(n1564), .Z(out[1143]) );
  XNOR U2651 ( .A(n1566), .B(n1565), .Z(n3926) );
  IV U2652 ( .A(n3926), .Z(n2653) );
  XOR U2653 ( .A(in[949]), .B(n2653), .Z(n1972) );
  NAND U2654 ( .A(n1567), .B(n1792), .Z(n1568) );
  XNOR U2655 ( .A(n1972), .B(n1568), .Z(out[1144]) );
  XOR U2656 ( .A(n1570), .B(n1569), .Z(n3065) );
  XOR U2657 ( .A(in[950]), .B(n3065), .Z(n1976) );
  NAND U2658 ( .A(n1571), .B(n1794), .Z(n1572) );
  XNOR U2659 ( .A(n1976), .B(n1572), .Z(out[1145]) );
  XOR U2660 ( .A(n1574), .B(n1573), .Z(n3067) );
  XOR U2661 ( .A(in[951]), .B(n3067), .Z(n1980) );
  NAND U2662 ( .A(n1575), .B(n1798), .Z(n1576) );
  XNOR U2663 ( .A(n1980), .B(n1576), .Z(out[1146]) );
  XOR U2664 ( .A(n1578), .B(n1577), .Z(n3070) );
  XOR U2665 ( .A(in[952]), .B(n3070), .Z(n1984) );
  NAND U2666 ( .A(n1579), .B(n1800), .Z(n1580) );
  XNOR U2667 ( .A(n1984), .B(n1580), .Z(out[1147]) );
  XNOR U2668 ( .A(n1582), .B(n1581), .Z(n3945) );
  IV U2669 ( .A(n3945), .Z(n2700) );
  XOR U2670 ( .A(in[953]), .B(n2700), .Z(n1988) );
  NAND U2671 ( .A(n1583), .B(n1802), .Z(n1584) );
  XNOR U2672 ( .A(n1988), .B(n1584), .Z(out[1148]) );
  XNOR U2673 ( .A(n1586), .B(n1585), .Z(n3949) );
  IV U2674 ( .A(n3949), .Z(n2702) );
  XOR U2675 ( .A(in[954]), .B(n2702), .Z(n1992) );
  NAND U2676 ( .A(n1587), .B(n1804), .Z(n1588) );
  XNOR U2677 ( .A(n1992), .B(n1588), .Z(out[1149]) );
  IV U2678 ( .A(n2023), .Z(n4012) );
  XOR U2679 ( .A(in[585]), .B(n4012), .Z(n2824) );
  IV U2680 ( .A(n1589), .Z(n4149) );
  XOR U2681 ( .A(in[1460]), .B(n4149), .Z(n3458) );
  XNOR U2682 ( .A(in[240]), .B(n4110), .Z(n3460) );
  NANDN U2683 ( .A(n3458), .B(n3460), .Z(n1590) );
  XNOR U2684 ( .A(n2824), .B(n1590), .Z(out[114]) );
  XOR U2685 ( .A(in[955]), .B(n3953), .Z(n1996) );
  NAND U2686 ( .A(n1591), .B(n1806), .Z(n1592) );
  XNOR U2687 ( .A(n1996), .B(n1592), .Z(out[1150]) );
  XOR U2688 ( .A(in[956]), .B(n3957), .Z(n2000) );
  NANDN U2689 ( .A(n1593), .B(n1808), .Z(n1594) );
  XNOR U2690 ( .A(n2000), .B(n1594), .Z(out[1151]) );
  XOR U2691 ( .A(n1596), .B(n1595), .Z(n4298) );
  XOR U2692 ( .A(in[1004]), .B(n4298), .Z(n1810) );
  NAND U2693 ( .A(n1597), .B(n1811), .Z(n1598) );
  XNOR U2694 ( .A(n1810), .B(n1598), .Z(out[1152]) );
  XOR U2695 ( .A(n1600), .B(n1599), .Z(n4300) );
  XOR U2696 ( .A(in[1005]), .B(n4300), .Z(n1813) );
  NAND U2697 ( .A(n1601), .B(n1814), .Z(n1602) );
  XNOR U2698 ( .A(n1813), .B(n1602), .Z(out[1153]) );
  XOR U2699 ( .A(n1604), .B(n1603), .Z(n4302) );
  XOR U2700 ( .A(in[1006]), .B(n4302), .Z(n1816) );
  NAND U2701 ( .A(n1605), .B(n1817), .Z(n1606) );
  XNOR U2702 ( .A(n1816), .B(n1606), .Z(out[1154]) );
  XOR U2703 ( .A(n1608), .B(n1607), .Z(n4304) );
  XOR U2704 ( .A(in[1007]), .B(n4304), .Z(n1819) );
  NAND U2705 ( .A(n1609), .B(n1820), .Z(n1610) );
  XNOR U2706 ( .A(n1819), .B(n1610), .Z(out[1155]) );
  XOR U2707 ( .A(n1612), .B(n1611), .Z(n4311) );
  XOR U2708 ( .A(in[1008]), .B(n4311), .Z(n1824) );
  NAND U2709 ( .A(n1613), .B(n1825), .Z(n1614) );
  XNOR U2710 ( .A(n1824), .B(n1614), .Z(out[1156]) );
  XOR U2711 ( .A(n1616), .B(n1615), .Z(n4314) );
  XOR U2712 ( .A(in[1009]), .B(n4314), .Z(n1827) );
  NAND U2713 ( .A(n1617), .B(n1828), .Z(n1618) );
  XNOR U2714 ( .A(n1827), .B(n1618), .Z(out[1157]) );
  XOR U2715 ( .A(n1620), .B(n1619), .Z(n4317) );
  XOR U2716 ( .A(in[1010]), .B(n4317), .Z(n5021) );
  NAND U2717 ( .A(n1621), .B(n1830), .Z(n1622) );
  XNOR U2718 ( .A(n5021), .B(n1622), .Z(out[1158]) );
  XOR U2719 ( .A(n1624), .B(n1623), .Z(n4320) );
  XOR U2720 ( .A(in[1011]), .B(n4320), .Z(n5025) );
  NAND U2721 ( .A(n1625), .B(n1831), .Z(n1626) );
  XNOR U2722 ( .A(n5025), .B(n1626), .Z(out[1159]) );
  IV U2723 ( .A(n2026), .Z(n4016) );
  XOR U2724 ( .A(in[586]), .B(n4016), .Z(n2826) );
  XNOR U2725 ( .A(in[1461]), .B(n4153), .Z(n3480) );
  XNOR U2726 ( .A(in[241]), .B(n4118), .Z(n3482) );
  NANDN U2727 ( .A(n3480), .B(n3482), .Z(n1627) );
  XNOR U2728 ( .A(n2826), .B(n1627), .Z(out[115]) );
  XOR U2729 ( .A(n1629), .B(n1628), .Z(n4323) );
  XOR U2730 ( .A(in[1012]), .B(n4323), .Z(n5029) );
  NAND U2731 ( .A(n1630), .B(n1833), .Z(n1631) );
  XNOR U2732 ( .A(n5029), .B(n1631), .Z(out[1160]) );
  XOR U2733 ( .A(n1633), .B(n1632), .Z(n4326) );
  XOR U2734 ( .A(in[1013]), .B(n4326), .Z(n5033) );
  NAND U2735 ( .A(n1634), .B(n1835), .Z(n1635) );
  XNOR U2736 ( .A(n5033), .B(n1635), .Z(out[1161]) );
  XOR U2737 ( .A(n1637), .B(n1636), .Z(n4329) );
  XOR U2738 ( .A(in[1014]), .B(n4329), .Z(n5041) );
  NAND U2739 ( .A(n1638), .B(n1837), .Z(n1639) );
  XNOR U2740 ( .A(n5041), .B(n1639), .Z(out[1162]) );
  XOR U2741 ( .A(n1641), .B(n1640), .Z(n4332) );
  XOR U2742 ( .A(in[1015]), .B(n4332), .Z(n5045) );
  NAND U2743 ( .A(n1642), .B(n1839), .Z(n1643) );
  XNOR U2744 ( .A(n5045), .B(n1643), .Z(out[1163]) );
  XOR U2745 ( .A(n1645), .B(n1644), .Z(n4178) );
  XOR U2746 ( .A(in[1016]), .B(n4178), .Z(n5049) );
  NAND U2747 ( .A(n1646), .B(n1841), .Z(n1647) );
  XNOR U2748 ( .A(n5049), .B(n1647), .Z(out[1164]) );
  XOR U2749 ( .A(n1649), .B(n1648), .Z(n4181) );
  XOR U2750 ( .A(in[1017]), .B(n4181), .Z(n5053) );
  NAND U2751 ( .A(n1650), .B(n1843), .Z(n1651) );
  XNOR U2752 ( .A(n5053), .B(n1651), .Z(out[1165]) );
  XOR U2753 ( .A(n1653), .B(n1652), .Z(n4184) );
  XOR U2754 ( .A(in[1018]), .B(n4184), .Z(n5057) );
  NAND U2755 ( .A(n1654), .B(n1847), .Z(n1655) );
  XNOR U2756 ( .A(n5057), .B(n1655), .Z(out[1166]) );
  XOR U2757 ( .A(n1657), .B(n1656), .Z(n4187) );
  XOR U2758 ( .A(in[1019]), .B(n4187), .Z(n5061) );
  NANDN U2759 ( .A(n1658), .B(n1849), .Z(n1659) );
  XNOR U2760 ( .A(n5061), .B(n1659), .Z(out[1167]) );
  IV U2761 ( .A(n3059), .Z(n4190) );
  XOR U2762 ( .A(in[1020]), .B(n4190), .Z(n5064) );
  NANDN U2763 ( .A(n1662), .B(n1851), .Z(n1663) );
  XOR U2764 ( .A(n5064), .B(n1663), .Z(out[1168]) );
  IV U2765 ( .A(n3061), .Z(n4193) );
  XOR U2766 ( .A(in[1021]), .B(n4193), .Z(n5067) );
  NANDN U2767 ( .A(n1666), .B(n1853), .Z(n1667) );
  XOR U2768 ( .A(n5067), .B(n1667), .Z(out[1169]) );
  IV U2769 ( .A(n2028), .Z(n4020) );
  XOR U2770 ( .A(in[587]), .B(n4020), .Z(n2828) );
  XNOR U2771 ( .A(in[1462]), .B(n4163), .Z(n3502) );
  XNOR U2772 ( .A(in[242]), .B(n4122), .Z(n3504) );
  NANDN U2773 ( .A(n3502), .B(n3504), .Z(n1668) );
  XNOR U2774 ( .A(n2828), .B(n1668), .Z(out[116]) );
  IV U2775 ( .A(n3063), .Z(n4198) );
  XOR U2776 ( .A(in[1022]), .B(n4198), .Z(n5070) );
  NANDN U2777 ( .A(n1671), .B(n1855), .Z(n1672) );
  XOR U2778 ( .A(n5070), .B(n1672), .Z(out[1170]) );
  XOR U2779 ( .A(n1674), .B(n1673), .Z(n4199) );
  XOR U2780 ( .A(in[1023]), .B(n4199), .Z(n5074) );
  NAND U2781 ( .A(n1675), .B(n1857), .Z(n1676) );
  XNOR U2782 ( .A(n5074), .B(n1676), .Z(out[1171]) );
  IV U2783 ( .A(n3068), .Z(n4200) );
  XOR U2784 ( .A(in[960]), .B(n4200), .Z(n5081) );
  NAND U2785 ( .A(n1679), .B(n1859), .Z(n1680) );
  XOR U2786 ( .A(n5081), .B(n1680), .Z(out[1172]) );
  IV U2787 ( .A(n3071), .Z(n4201) );
  XOR U2788 ( .A(in[961]), .B(n4201), .Z(n5084) );
  NAND U2789 ( .A(n1683), .B(n1861), .Z(n1684) );
  XOR U2790 ( .A(n5084), .B(n1684), .Z(out[1173]) );
  IV U2791 ( .A(n3073), .Z(n4202) );
  XOR U2792 ( .A(in[962]), .B(n4202), .Z(n5087) );
  NAND U2793 ( .A(n1687), .B(n1863), .Z(n1688) );
  XOR U2794 ( .A(n5087), .B(n1688), .Z(out[1174]) );
  IV U2795 ( .A(n3077), .Z(n4203) );
  XOR U2796 ( .A(in[963]), .B(n4203), .Z(n5090) );
  NAND U2797 ( .A(n1691), .B(n1865), .Z(n1692) );
  XOR U2798 ( .A(n5090), .B(n1692), .Z(out[1175]) );
  IV U2799 ( .A(n3079), .Z(n4204) );
  XOR U2800 ( .A(in[964]), .B(n4204), .Z(n5093) );
  NAND U2801 ( .A(n1695), .B(n1869), .Z(n1696) );
  XOR U2802 ( .A(n5093), .B(n1696), .Z(out[1176]) );
  IV U2803 ( .A(n3081), .Z(n4205) );
  XOR U2804 ( .A(in[965]), .B(n4205), .Z(n5096) );
  NAND U2805 ( .A(n1699), .B(n1871), .Z(n1700) );
  XOR U2806 ( .A(n5096), .B(n1700), .Z(out[1177]) );
  IV U2807 ( .A(n3083), .Z(n4208) );
  XOR U2808 ( .A(in[966]), .B(n4208), .Z(n5099) );
  NAND U2809 ( .A(n1703), .B(n1873), .Z(n1704) );
  XOR U2810 ( .A(n5099), .B(n1704), .Z(out[1178]) );
  IV U2811 ( .A(n3085), .Z(n4211) );
  XOR U2812 ( .A(in[967]), .B(n4211), .Z(n5102) );
  NAND U2813 ( .A(n1707), .B(n1875), .Z(n1708) );
  XOR U2814 ( .A(n5102), .B(n1708), .Z(out[1179]) );
  IV U2815 ( .A(n2030), .Z(n4028) );
  XOR U2816 ( .A(in[588]), .B(n4028), .Z(n2830) );
  XNOR U2817 ( .A(in[1463]), .B(n4167), .Z(n3517) );
  XNOR U2818 ( .A(in[243]), .B(n4126), .Z(n3519) );
  NANDN U2819 ( .A(n3517), .B(n3519), .Z(n1709) );
  XNOR U2820 ( .A(n2830), .B(n1709), .Z(out[117]) );
  XNOR U2821 ( .A(n1711), .B(n1710), .Z(n4216) );
  XOR U2822 ( .A(in[968]), .B(n4216), .Z(n5106) );
  NAND U2823 ( .A(n1712), .B(n1877), .Z(n1713) );
  XNOR U2824 ( .A(n5106), .B(n1713), .Z(out[1180]) );
  IV U2825 ( .A(n3088), .Z(n4219) );
  XOR U2826 ( .A(in[969]), .B(n4219), .Z(n5109) );
  NAND U2827 ( .A(n1716), .B(n1879), .Z(n1717) );
  XOR U2828 ( .A(n5109), .B(n1717), .Z(out[1181]) );
  IV U2829 ( .A(n3090), .Z(n4222) );
  XOR U2830 ( .A(in[970]), .B(n4222), .Z(n5116) );
  NAND U2831 ( .A(n1720), .B(n1881), .Z(n1721) );
  XOR U2832 ( .A(n5116), .B(n1721), .Z(out[1182]) );
  XOR U2833 ( .A(in[971]), .B(n3092), .Z(n5120) );
  NAND U2834 ( .A(n1724), .B(n1883), .Z(n1725) );
  XNOR U2835 ( .A(n5120), .B(n1725), .Z(out[1183]) );
  XOR U2836 ( .A(in[972]), .B(n3094), .Z(n5124) );
  NAND U2837 ( .A(n1728), .B(n1885), .Z(n1729) );
  XNOR U2838 ( .A(n5124), .B(n1729), .Z(out[1184]) );
  XOR U2839 ( .A(in[973]), .B(n3098), .Z(n5128) );
  NAND U2840 ( .A(n1732), .B(n1887), .Z(n1733) );
  XNOR U2841 ( .A(n5128), .B(n1733), .Z(out[1185]) );
  XOR U2842 ( .A(n1735), .B(n1734), .Z(n4234) );
  XOR U2843 ( .A(in[974]), .B(n4234), .Z(n5132) );
  NAND U2844 ( .A(n1736), .B(n1891), .Z(n1737) );
  XNOR U2845 ( .A(n5132), .B(n1737), .Z(out[1186]) );
  XOR U2846 ( .A(n1739), .B(n1738), .Z(n4237) );
  XOR U2847 ( .A(in[975]), .B(n4237), .Z(n5136) );
  NAND U2848 ( .A(n1740), .B(n1893), .Z(n1741) );
  XNOR U2849 ( .A(n5136), .B(n1741), .Z(out[1187]) );
  XOR U2850 ( .A(n1743), .B(n1742), .Z(n4240) );
  XOR U2851 ( .A(in[976]), .B(n4240), .Z(n5140) );
  NAND U2852 ( .A(n1744), .B(n1895), .Z(n1745) );
  XNOR U2853 ( .A(n5140), .B(n1745), .Z(out[1188]) );
  XOR U2854 ( .A(n1747), .B(n1746), .Z(n4241) );
  XOR U2855 ( .A(in[977]), .B(n4241), .Z(n5144) );
  NAND U2856 ( .A(n1748), .B(n1897), .Z(n1749) );
  XNOR U2857 ( .A(n5144), .B(n1749), .Z(out[1189]) );
  IV U2858 ( .A(n3110), .Z(n4032) );
  XOR U2859 ( .A(in[589]), .B(n4032), .Z(n2832) );
  XNOR U2860 ( .A(in[1464]), .B(n4171), .Z(n3545) );
  XNOR U2861 ( .A(in[244]), .B(n4130), .Z(n3547) );
  NANDN U2862 ( .A(n3545), .B(n3547), .Z(n1750) );
  XNOR U2863 ( .A(n2832), .B(n1750), .Z(out[118]) );
  XOR U2864 ( .A(in[978]), .B(n3104), .Z(n5147) );
  NAND U2865 ( .A(n1753), .B(n1899), .Z(n1754) );
  XNOR U2866 ( .A(n5147), .B(n1754), .Z(out[1190]) );
  XOR U2867 ( .A(in[979]), .B(n3106), .Z(n5152) );
  NAND U2868 ( .A(n1757), .B(n1901), .Z(n1758) );
  XNOR U2869 ( .A(n5152), .B(n1758), .Z(out[1191]) );
  OR U2870 ( .A(n1904), .B(n1759), .Z(n1760) );
  XNOR U2871 ( .A(n1903), .B(n1760), .Z(out[1192]) );
  OR U2872 ( .A(n1908), .B(n1761), .Z(n1762) );
  XNOR U2873 ( .A(n1907), .B(n1762), .Z(out[1193]) );
  OR U2874 ( .A(n1912), .B(n1763), .Z(n1764) );
  XNOR U2875 ( .A(n1911), .B(n1764), .Z(out[1194]) );
  OR U2876 ( .A(n1922), .B(n1766), .Z(n1767) );
  XNOR U2877 ( .A(n1921), .B(n1767), .Z(out[1196]) );
  OR U2878 ( .A(n1926), .B(n1768), .Z(n1769) );
  XNOR U2879 ( .A(n1925), .B(n1769), .Z(out[1197]) );
  OR U2880 ( .A(n1930), .B(n1770), .Z(n1771) );
  XNOR U2881 ( .A(n1929), .B(n1771), .Z(out[1198]) );
  OR U2882 ( .A(n1934), .B(n1772), .Z(n1773) );
  XNOR U2883 ( .A(n1933), .B(n1773), .Z(out[1199]) );
  IV U2884 ( .A(n3116), .Z(n4036) );
  XOR U2885 ( .A(in[590]), .B(n4036), .Z(n2834) );
  XNOR U2886 ( .A(in[1465]), .B(n4175), .Z(n3575) );
  XNOR U2887 ( .A(in[245]), .B(n4134), .Z(n3577) );
  NANDN U2888 ( .A(n3575), .B(n3577), .Z(n1774) );
  XNOR U2889 ( .A(n2834), .B(n1774), .Z(out[119]) );
  XNOR U2890 ( .A(in[201]), .B(n3942), .Z(n4307) );
  XOR U2891 ( .A(in[1421]), .B(n3196), .Z(n4308) );
  XNOR U2892 ( .A(in[1044]), .B(n4488), .Z(n2883) );
  NANDN U2893 ( .A(n4308), .B(n2883), .Z(n1775) );
  XNOR U2894 ( .A(n4307), .B(n1775), .Z(out[11]) );
  OR U2895 ( .A(n1938), .B(n1776), .Z(n1777) );
  XNOR U2896 ( .A(n1937), .B(n1777), .Z(out[1200]) );
  OR U2897 ( .A(n1942), .B(n1778), .Z(n1779) );
  XNOR U2898 ( .A(n1941), .B(n1779), .Z(out[1201]) );
  OR U2899 ( .A(n1946), .B(n1780), .Z(n1781) );
  XNOR U2900 ( .A(n1945), .B(n1781), .Z(out[1202]) );
  OR U2901 ( .A(n1950), .B(n1782), .Z(n1783) );
  XNOR U2902 ( .A(n1949), .B(n1783), .Z(out[1203]) );
  OR U2903 ( .A(n1954), .B(n1784), .Z(n1785) );
  XNOR U2904 ( .A(n1953), .B(n1785), .Z(out[1204]) );
  OR U2905 ( .A(n1958), .B(n1786), .Z(n1787) );
  XNOR U2906 ( .A(n1957), .B(n1787), .Z(out[1205]) );
  OR U2907 ( .A(n1964), .B(n1788), .Z(n1789) );
  XNOR U2908 ( .A(n1963), .B(n1789), .Z(out[1206]) );
  OR U2909 ( .A(n1968), .B(n1790), .Z(n1791) );
  XNOR U2910 ( .A(n1967), .B(n1791), .Z(out[1207]) );
  OR U2911 ( .A(n1972), .B(n1792), .Z(n1793) );
  XNOR U2912 ( .A(n1971), .B(n1793), .Z(out[1208]) );
  OR U2913 ( .A(n1976), .B(n1794), .Z(n1795) );
  XNOR U2914 ( .A(n1975), .B(n1795), .Z(out[1209]) );
  IV U2915 ( .A(n3118), .Z(n4040) );
  XOR U2916 ( .A(in[591]), .B(n4040), .Z(n2836) );
  IV U2917 ( .A(n1796), .Z(n3899) );
  XOR U2918 ( .A(in[1466]), .B(n3899), .Z(n3599) );
  XNOR U2919 ( .A(in[246]), .B(n4138), .Z(n3601) );
  NANDN U2920 ( .A(n3599), .B(n3601), .Z(n1797) );
  XNOR U2921 ( .A(n2836), .B(n1797), .Z(out[120]) );
  OR U2922 ( .A(n1980), .B(n1798), .Z(n1799) );
  XNOR U2923 ( .A(n1979), .B(n1799), .Z(out[1210]) );
  OR U2924 ( .A(n1984), .B(n1800), .Z(n1801) );
  XNOR U2925 ( .A(n1983), .B(n1801), .Z(out[1211]) );
  OR U2926 ( .A(n1988), .B(n1802), .Z(n1803) );
  XNOR U2927 ( .A(n1987), .B(n1803), .Z(out[1212]) );
  OR U2928 ( .A(n1992), .B(n1804), .Z(n1805) );
  XNOR U2929 ( .A(n1991), .B(n1805), .Z(out[1213]) );
  OR U2930 ( .A(n1996), .B(n1806), .Z(n1807) );
  XNOR U2931 ( .A(n1995), .B(n1807), .Z(out[1214]) );
  OR U2932 ( .A(n2000), .B(n1808), .Z(n1809) );
  XNOR U2933 ( .A(n1999), .B(n1809), .Z(out[1215]) );
  IV U2934 ( .A(n1810), .Z(n4996) );
  NANDN U2935 ( .A(n1811), .B(n4996), .Z(n1812) );
  XOR U2936 ( .A(n4997), .B(n1812), .Z(out[1216]) );
  IV U2937 ( .A(n1813), .Z(n5000) );
  NANDN U2938 ( .A(n1814), .B(n5000), .Z(n1815) );
  XOR U2939 ( .A(n5001), .B(n1815), .Z(out[1217]) );
  IV U2940 ( .A(n1816), .Z(n5004) );
  NANDN U2941 ( .A(n1817), .B(n5004), .Z(n1818) );
  XOR U2942 ( .A(n5005), .B(n1818), .Z(out[1218]) );
  IV U2943 ( .A(n1819), .Z(n5008) );
  NANDN U2944 ( .A(n1820), .B(n5008), .Z(n1821) );
  XOR U2945 ( .A(n5009), .B(n1821), .Z(out[1219]) );
  IV U2946 ( .A(n3120), .Z(n4044) );
  XOR U2947 ( .A(in[592]), .B(n4044), .Z(n2838) );
  IV U2948 ( .A(n1822), .Z(n3903) );
  XOR U2949 ( .A(in[1467]), .B(n3903), .Z(n3629) );
  XNOR U2950 ( .A(in[247]), .B(n4142), .Z(n3631) );
  NANDN U2951 ( .A(n3629), .B(n3631), .Z(n1823) );
  XNOR U2952 ( .A(n2838), .B(n1823), .Z(out[121]) );
  IV U2953 ( .A(n1824), .Z(n5012) );
  NANDN U2954 ( .A(n1825), .B(n5012), .Z(n1826) );
  XOR U2955 ( .A(n5013), .B(n1826), .Z(out[1220]) );
  IV U2956 ( .A(n1827), .Z(n5016) );
  NANDN U2957 ( .A(n1828), .B(n5016), .Z(n1829) );
  XOR U2958 ( .A(n5017), .B(n1829), .Z(out[1221]) );
  OR U2959 ( .A(n5025), .B(n1831), .Z(n1832) );
  XNOR U2960 ( .A(n5024), .B(n1832), .Z(out[1223]) );
  OR U2961 ( .A(n5029), .B(n1833), .Z(n1834) );
  XNOR U2962 ( .A(n5028), .B(n1834), .Z(out[1224]) );
  OR U2963 ( .A(n5033), .B(n1835), .Z(n1836) );
  XNOR U2964 ( .A(n5032), .B(n1836), .Z(out[1225]) );
  OR U2965 ( .A(n5041), .B(n1837), .Z(n1838) );
  XNOR U2966 ( .A(n5040), .B(n1838), .Z(out[1226]) );
  OR U2967 ( .A(n5045), .B(n1839), .Z(n1840) );
  XNOR U2968 ( .A(n5044), .B(n1840), .Z(out[1227]) );
  OR U2969 ( .A(n5049), .B(n1841), .Z(n1842) );
  XNOR U2970 ( .A(n5048), .B(n1842), .Z(out[1228]) );
  OR U2971 ( .A(n5053), .B(n1843), .Z(n1844) );
  XNOR U2972 ( .A(n5052), .B(n1844), .Z(out[1229]) );
  XNOR U2973 ( .A(in[593]), .B(n4048), .Z(n2843) );
  IV U2974 ( .A(n1845), .Z(n3907) );
  XOR U2975 ( .A(in[1468]), .B(n3907), .Z(n3673) );
  XNOR U2976 ( .A(in[248]), .B(n4146), .Z(n3675) );
  NANDN U2977 ( .A(n3673), .B(n3675), .Z(n1846) );
  XNOR U2978 ( .A(n2843), .B(n1846), .Z(out[122]) );
  OR U2979 ( .A(n5057), .B(n1847), .Z(n1848) );
  XNOR U2980 ( .A(n5056), .B(n1848), .Z(out[1230]) );
  OR U2981 ( .A(n5061), .B(n1849), .Z(n1850) );
  XNOR U2982 ( .A(n5060), .B(n1850), .Z(out[1231]) );
  NANDN U2983 ( .A(n1851), .B(n5064), .Z(n1852) );
  XNOR U2984 ( .A(n5065), .B(n1852), .Z(out[1232]) );
  NANDN U2985 ( .A(n1853), .B(n5067), .Z(n1854) );
  XNOR U2986 ( .A(n5068), .B(n1854), .Z(out[1233]) );
  NANDN U2987 ( .A(n1855), .B(n5070), .Z(n1856) );
  XNOR U2988 ( .A(n5071), .B(n1856), .Z(out[1234]) );
  OR U2989 ( .A(n5074), .B(n1857), .Z(n1858) );
  XNOR U2990 ( .A(n5073), .B(n1858), .Z(out[1235]) );
  NANDN U2991 ( .A(n1859), .B(n5081), .Z(n1860) );
  XNOR U2992 ( .A(n5082), .B(n1860), .Z(out[1236]) );
  NANDN U2993 ( .A(n1861), .B(n5084), .Z(n1862) );
  XNOR U2994 ( .A(n5085), .B(n1862), .Z(out[1237]) );
  NANDN U2995 ( .A(n1863), .B(n5087), .Z(n1864) );
  XNOR U2996 ( .A(n5088), .B(n1864), .Z(out[1238]) );
  NANDN U2997 ( .A(n1865), .B(n5090), .Z(n1866) );
  XNOR U2998 ( .A(n5091), .B(n1866), .Z(out[1239]) );
  IV U2999 ( .A(n2038), .Z(n4052) );
  XOR U3000 ( .A(in[594]), .B(n4052), .Z(n2845) );
  IV U3001 ( .A(n1867), .Z(n3911) );
  XOR U3002 ( .A(in[1469]), .B(n3911), .Z(n3717) );
  XNOR U3003 ( .A(in[249]), .B(n4150), .Z(n3719) );
  NANDN U3004 ( .A(n3717), .B(n3719), .Z(n1868) );
  XNOR U3005 ( .A(n2845), .B(n1868), .Z(out[123]) );
  NANDN U3006 ( .A(n1869), .B(n5093), .Z(n1870) );
  XNOR U3007 ( .A(n5094), .B(n1870), .Z(out[1240]) );
  NANDN U3008 ( .A(n1871), .B(n5096), .Z(n1872) );
  XNOR U3009 ( .A(n5097), .B(n1872), .Z(out[1241]) );
  NANDN U3010 ( .A(n1873), .B(n5099), .Z(n1874) );
  XNOR U3011 ( .A(n5100), .B(n1874), .Z(out[1242]) );
  NANDN U3012 ( .A(n1875), .B(n5102), .Z(n1876) );
  XNOR U3013 ( .A(n5103), .B(n1876), .Z(out[1243]) );
  OR U3014 ( .A(n5106), .B(n1877), .Z(n1878) );
  XNOR U3015 ( .A(n5105), .B(n1878), .Z(out[1244]) );
  NANDN U3016 ( .A(n1879), .B(n5109), .Z(n1880) );
  XNOR U3017 ( .A(n5110), .B(n1880), .Z(out[1245]) );
  NANDN U3018 ( .A(n1881), .B(n5116), .Z(n1882) );
  XNOR U3019 ( .A(n5117), .B(n1882), .Z(out[1246]) );
  OR U3020 ( .A(n5120), .B(n1883), .Z(n1884) );
  XNOR U3021 ( .A(n5119), .B(n1884), .Z(out[1247]) );
  OR U3022 ( .A(n5124), .B(n1885), .Z(n1886) );
  XNOR U3023 ( .A(n5123), .B(n1886), .Z(out[1248]) );
  OR U3024 ( .A(n5128), .B(n1887), .Z(n1888) );
  XNOR U3025 ( .A(n5127), .B(n1888), .Z(out[1249]) );
  IV U3026 ( .A(n3124), .Z(n4056) );
  XOR U3027 ( .A(in[595]), .B(n4056), .Z(n2847) );
  IV U3028 ( .A(n1889), .Z(n3915) );
  XOR U3029 ( .A(in[1470]), .B(n3915), .Z(n3763) );
  XNOR U3030 ( .A(in[250]), .B(n4154), .Z(n3765) );
  NANDN U3031 ( .A(n3763), .B(n3765), .Z(n1890) );
  XNOR U3032 ( .A(n2847), .B(n1890), .Z(out[124]) );
  OR U3033 ( .A(n5132), .B(n1891), .Z(n1892) );
  XNOR U3034 ( .A(n5131), .B(n1892), .Z(out[1250]) );
  OR U3035 ( .A(n5136), .B(n1893), .Z(n1894) );
  XNOR U3036 ( .A(n5135), .B(n1894), .Z(out[1251]) );
  OR U3037 ( .A(n5140), .B(n1895), .Z(n1896) );
  XNOR U3038 ( .A(n5139), .B(n1896), .Z(out[1252]) );
  OR U3039 ( .A(n5144), .B(n1897), .Z(n1898) );
  XNOR U3040 ( .A(n5143), .B(n1898), .Z(out[1253]) );
  OR U3041 ( .A(n5147), .B(n1899), .Z(n1900) );
  XOR U3042 ( .A(n5148), .B(n1900), .Z(out[1254]) );
  OR U3043 ( .A(n5152), .B(n1901), .Z(n1902) );
  XNOR U3044 ( .A(n5151), .B(n1902), .Z(out[1255]) );
  ANDN U3045 ( .B(n1904), .A(n1903), .Z(n1905) );
  XOR U3046 ( .A(n1906), .B(n1905), .Z(out[1256]) );
  ANDN U3047 ( .B(n1908), .A(n1907), .Z(n1909) );
  XOR U3048 ( .A(n1910), .B(n1909), .Z(out[1257]) );
  ANDN U3049 ( .B(n1912), .A(n1911), .Z(n1913) );
  XOR U3050 ( .A(n1914), .B(n1913), .Z(out[1258]) );
  ANDN U3051 ( .B(n1916), .A(n1915), .Z(n1917) );
  XOR U3052 ( .A(n1918), .B(n1917), .Z(out[1259]) );
  IV U3053 ( .A(n3126), .Z(n4060) );
  XOR U3054 ( .A(in[596]), .B(n4060), .Z(n2849) );
  IV U3055 ( .A(n1919), .Z(n3919) );
  XOR U3056 ( .A(in[1471]), .B(n3919), .Z(n3807) );
  IV U3057 ( .A(n4164), .Z(n3279) );
  XOR U3058 ( .A(in[251]), .B(n3279), .Z(n3809) );
  OR U3059 ( .A(n3807), .B(n3809), .Z(n1920) );
  XNOR U3060 ( .A(n2849), .B(n1920), .Z(out[125]) );
  ANDN U3061 ( .B(n1922), .A(n1921), .Z(n1923) );
  XOR U3062 ( .A(n1924), .B(n1923), .Z(out[1260]) );
  ANDN U3063 ( .B(n1926), .A(n1925), .Z(n1927) );
  XOR U3064 ( .A(n1928), .B(n1927), .Z(out[1261]) );
  ANDN U3065 ( .B(n1930), .A(n1929), .Z(n1931) );
  XOR U3066 ( .A(n1932), .B(n1931), .Z(out[1262]) );
  ANDN U3067 ( .B(n1934), .A(n1933), .Z(n1935) );
  XOR U3068 ( .A(n1936), .B(n1935), .Z(out[1263]) );
  ANDN U3069 ( .B(n1938), .A(n1937), .Z(n1939) );
  XOR U3070 ( .A(n1940), .B(n1939), .Z(out[1264]) );
  ANDN U3071 ( .B(n1942), .A(n1941), .Z(n1943) );
  XOR U3072 ( .A(n1944), .B(n1943), .Z(out[1265]) );
  ANDN U3073 ( .B(n1946), .A(n1945), .Z(n1947) );
  XOR U3074 ( .A(n1948), .B(n1947), .Z(out[1266]) );
  ANDN U3075 ( .B(n1950), .A(n1949), .Z(n1951) );
  XOR U3076 ( .A(n1952), .B(n1951), .Z(out[1267]) );
  ANDN U3077 ( .B(n1954), .A(n1953), .Z(n1955) );
  XOR U3078 ( .A(n1956), .B(n1955), .Z(out[1268]) );
  ANDN U3079 ( .B(n1958), .A(n1957), .Z(n1959) );
  XOR U3080 ( .A(n1960), .B(n1959), .Z(out[1269]) );
  IV U3081 ( .A(n3128), .Z(n4064) );
  XOR U3082 ( .A(in[597]), .B(n4064), .Z(n2851) );
  IV U3083 ( .A(n1961), .Z(n3923) );
  XOR U3084 ( .A(in[1408]), .B(n3923), .Z(n3851) );
  IV U3085 ( .A(n4168), .Z(n3282) );
  XOR U3086 ( .A(in[252]), .B(n3282), .Z(n3853) );
  OR U3087 ( .A(n3851), .B(n3853), .Z(n1962) );
  XNOR U3088 ( .A(n2851), .B(n1962), .Z(out[126]) );
  ANDN U3089 ( .B(n1964), .A(n1963), .Z(n1965) );
  XOR U3090 ( .A(n1966), .B(n1965), .Z(out[1270]) );
  ANDN U3091 ( .B(n1968), .A(n1967), .Z(n1969) );
  XOR U3092 ( .A(n1970), .B(n1969), .Z(out[1271]) );
  ANDN U3093 ( .B(n1972), .A(n1971), .Z(n1973) );
  XOR U3094 ( .A(n1974), .B(n1973), .Z(out[1272]) );
  ANDN U3095 ( .B(n1976), .A(n1975), .Z(n1977) );
  XOR U3096 ( .A(n1978), .B(n1977), .Z(out[1273]) );
  ANDN U3097 ( .B(n1980), .A(n1979), .Z(n1981) );
  XOR U3098 ( .A(n1982), .B(n1981), .Z(out[1274]) );
  ANDN U3099 ( .B(n1984), .A(n1983), .Z(n1985) );
  XOR U3100 ( .A(n1986), .B(n1985), .Z(out[1275]) );
  ANDN U3101 ( .B(n1988), .A(n1987), .Z(n1989) );
  XOR U3102 ( .A(n1990), .B(n1989), .Z(out[1276]) );
  ANDN U3103 ( .B(n1992), .A(n1991), .Z(n1993) );
  XOR U3104 ( .A(n1994), .B(n1993), .Z(out[1277]) );
  ANDN U3105 ( .B(n1996), .A(n1995), .Z(n1997) );
  XOR U3106 ( .A(n1998), .B(n1997), .Z(out[1278]) );
  ANDN U3107 ( .B(n2000), .A(n1999), .Z(n2001) );
  XOR U3108 ( .A(n2002), .B(n2001), .Z(out[1279]) );
  IV U3109 ( .A(n3130), .Z(n4072) );
  XOR U3110 ( .A(in[598]), .B(n4072), .Z(n2853) );
  IV U3111 ( .A(n2003), .Z(n3927) );
  XOR U3112 ( .A(in[1409]), .B(n3927), .Z(n3895) );
  IV U3113 ( .A(n4172), .Z(n3285) );
  XOR U3114 ( .A(in[253]), .B(n3285), .Z(n3897) );
  OR U3115 ( .A(n3895), .B(n3897), .Z(n2004) );
  XNOR U3116 ( .A(n2853), .B(n2004), .Z(out[127]) );
  XOR U3117 ( .A(in[50]), .B(n4317), .Z(n2179) );
  XNOR U3118 ( .A(in[1172]), .B(n3989), .Z(n2435) );
  XNOR U3119 ( .A(in[1536]), .B(n3973), .Z(n2436) );
  NANDN U3120 ( .A(n2435), .B(n2436), .Z(n2005) );
  XNOR U3121 ( .A(n2179), .B(n2005), .Z(out[1280]) );
  XOR U3122 ( .A(in[51]), .B(n4320), .Z(n2181) );
  IV U3123 ( .A(n2006), .Z(n3993) );
  XOR U3124 ( .A(in[1173]), .B(n3993), .Z(n2438) );
  XNOR U3125 ( .A(in[1537]), .B(n3977), .Z(n2096) );
  IV U3126 ( .A(n2096), .Z(n2439) );
  OR U3127 ( .A(n2438), .B(n2439), .Z(n2007) );
  XNOR U3128 ( .A(n2181), .B(n2007), .Z(out[1281]) );
  XOR U3129 ( .A(in[52]), .B(n4323), .Z(n2184) );
  IV U3130 ( .A(n2008), .Z(n3997) );
  XOR U3131 ( .A(in[1174]), .B(n3997), .Z(n2443) );
  XNOR U3132 ( .A(in[1538]), .B(n3984), .Z(n2098) );
  IV U3133 ( .A(n2098), .Z(n2445) );
  OR U3134 ( .A(n2443), .B(n2445), .Z(n2009) );
  XNOR U3135 ( .A(n2184), .B(n2009), .Z(out[1282]) );
  XOR U3136 ( .A(in[53]), .B(n4326), .Z(n2186) );
  XNOR U3137 ( .A(in[1175]), .B(n4001), .Z(n2447) );
  XNOR U3138 ( .A(in[1539]), .B(n3988), .Z(n2448) );
  NANDN U3139 ( .A(n2447), .B(n2448), .Z(n2010) );
  XNOR U3140 ( .A(n2186), .B(n2010), .Z(out[1283]) );
  XOR U3141 ( .A(in[54]), .B(n4329), .Z(n2188) );
  XNOR U3142 ( .A(in[1176]), .B(n4005), .Z(n2454) );
  XOR U3143 ( .A(in[1540]), .B(n2011), .Z(n2452) );
  NANDN U3144 ( .A(n2454), .B(n2452), .Z(n2012) );
  XNOR U3145 ( .A(n2188), .B(n2012), .Z(out[1284]) );
  XOR U3146 ( .A(in[55]), .B(n4332), .Z(n2190) );
  XNOR U3147 ( .A(in[1177]), .B(n4009), .Z(n2457) );
  XOR U3148 ( .A(in[1541]), .B(n2013), .Z(n2455) );
  NANDN U3149 ( .A(n2457), .B(n2455), .Z(n2014) );
  XNOR U3150 ( .A(n2190), .B(n2014), .Z(out[1285]) );
  XOR U3151 ( .A(in[56]), .B(n4178), .Z(n2192) );
  IV U3152 ( .A(n2015), .Z(n4013) );
  XOR U3153 ( .A(in[1178]), .B(n4013), .Z(n2459) );
  XOR U3154 ( .A(in[1542]), .B(n2016), .Z(n2104) );
  IV U3155 ( .A(n2104), .Z(n2461) );
  OR U3156 ( .A(n2459), .B(n2461), .Z(n2017) );
  XNOR U3157 ( .A(n2192), .B(n2017), .Z(out[1286]) );
  XOR U3158 ( .A(in[57]), .B(n4181), .Z(n2194) );
  IV U3159 ( .A(n2018), .Z(n4017) );
  XOR U3160 ( .A(in[1179]), .B(n4017), .Z(n2463) );
  XOR U3161 ( .A(in[1543]), .B(n2019), .Z(n2106) );
  IV U3162 ( .A(n2106), .Z(n2464) );
  OR U3163 ( .A(n2463), .B(n2464), .Z(n2020) );
  XNOR U3164 ( .A(n2194), .B(n2020), .Z(out[1287]) );
  XOR U3165 ( .A(in[58]), .B(n4184), .Z(n2196) );
  XNOR U3166 ( .A(in[1180]), .B(n4021), .Z(n2469) );
  XOR U3167 ( .A(in[1544]), .B(n2021), .Z(n2467) );
  NANDN U3168 ( .A(n2469), .B(n2467), .Z(n2022) );
  XNOR U3169 ( .A(n2196), .B(n2022), .Z(out[1288]) );
  XOR U3170 ( .A(in[59]), .B(n4187), .Z(n2198) );
  XNOR U3171 ( .A(in[1181]), .B(n4029), .Z(n2472) );
  XOR U3172 ( .A(in[1545]), .B(n2023), .Z(n2470) );
  NANDN U3173 ( .A(n2472), .B(n2470), .Z(n2024) );
  XNOR U3174 ( .A(n2198), .B(n2024), .Z(out[1289]) );
  XOR U3175 ( .A(in[665]), .B(n4255), .Z(n2855) );
  IV U3176 ( .A(n3132), .Z(n4076) );
  XOR U3177 ( .A(in[599]), .B(n4076), .Z(n3940) );
  OR U3178 ( .A(n3940), .B(n3938), .Z(n2025) );
  XNOR U3179 ( .A(n2855), .B(n2025), .Z(out[128]) );
  XOR U3180 ( .A(in[60]), .B(n3059), .Z(n2200) );
  XNOR U3181 ( .A(in[1182]), .B(n4033), .Z(n2475) );
  XOR U3182 ( .A(in[1546]), .B(n2026), .Z(n2473) );
  NANDN U3183 ( .A(n2475), .B(n2473), .Z(n2027) );
  XNOR U3184 ( .A(n2200), .B(n2027), .Z(out[1290]) );
  XOR U3185 ( .A(in[61]), .B(n3061), .Z(n2202) );
  XNOR U3186 ( .A(in[1183]), .B(n4037), .Z(n2478) );
  XOR U3187 ( .A(in[1547]), .B(n2028), .Z(n2476) );
  NANDN U3188 ( .A(n2478), .B(n2476), .Z(n2029) );
  XNOR U3189 ( .A(n2202), .B(n2029), .Z(out[1291]) );
  XOR U3190 ( .A(in[62]), .B(n3063), .Z(n2205) );
  XNOR U3191 ( .A(in[1184]), .B(n4041), .Z(n2481) );
  XOR U3192 ( .A(in[1548]), .B(n2030), .Z(n2479) );
  NANDN U3193 ( .A(n2481), .B(n2479), .Z(n2031) );
  XNOR U3194 ( .A(n2205), .B(n2031), .Z(out[1292]) );
  XOR U3195 ( .A(in[63]), .B(n4199), .Z(n2207) );
  XNOR U3196 ( .A(in[1185]), .B(n4045), .Z(n2484) );
  XOR U3197 ( .A(in[1549]), .B(n3110), .Z(n2482) );
  NANDN U3198 ( .A(n2484), .B(n2482), .Z(n2032) );
  XNOR U3199 ( .A(n2207), .B(n2032), .Z(out[1293]) );
  XOR U3200 ( .A(in[0]), .B(n3068), .Z(n2209) );
  XOR U3201 ( .A(in[1550]), .B(n3116), .Z(n2114) );
  IV U3202 ( .A(n2114), .Z(n2489) );
  XNOR U3203 ( .A(n3395), .B(in[1186]), .Z(n2486) );
  NANDN U3204 ( .A(n2489), .B(n2486), .Z(n2033) );
  XNOR U3205 ( .A(n2209), .B(n2033), .Z(out[1294]) );
  XOR U3206 ( .A(in[1]), .B(n3071), .Z(n2211) );
  XOR U3207 ( .A(in[1551]), .B(n4040), .Z(n2492) );
  XNOR U3208 ( .A(n3398), .B(in[1187]), .Z(n2490) );
  NANDN U3209 ( .A(n2492), .B(n2490), .Z(n2034) );
  XNOR U3210 ( .A(n2211), .B(n2034), .Z(out[1295]) );
  XOR U3211 ( .A(in[2]), .B(n3073), .Z(n2214) );
  XOR U3212 ( .A(n3402), .B(in[1188]), .Z(n2496) );
  XOR U3213 ( .A(in[1552]), .B(n4044), .Z(n2498) );
  OR U3214 ( .A(n2496), .B(n2498), .Z(n2035) );
  XNOR U3215 ( .A(n2214), .B(n2035), .Z(out[1296]) );
  XOR U3216 ( .A(in[3]), .B(n3077), .Z(n2216) );
  XOR U3217 ( .A(n3406), .B(in[1189]), .Z(n2500) );
  XNOR U3218 ( .A(in[1553]), .B(n4048), .Z(n2502) );
  OR U3219 ( .A(n2500), .B(n2502), .Z(n2036) );
  XNOR U3220 ( .A(n2216), .B(n2036), .Z(out[1297]) );
  XOR U3221 ( .A(in[4]), .B(n3079), .Z(n2218) );
  IV U3222 ( .A(n2037), .Z(n4065) );
  XOR U3223 ( .A(in[1190]), .B(n4065), .Z(n2504) );
  XOR U3224 ( .A(in[1554]), .B(n2038), .Z(n2119) );
  IV U3225 ( .A(n2119), .Z(n2506) );
  OR U3226 ( .A(n2504), .B(n2506), .Z(n2039) );
  XNOR U3227 ( .A(n2218), .B(n2039), .Z(out[1298]) );
  XOR U3228 ( .A(in[5]), .B(n3081), .Z(n2220) );
  IV U3229 ( .A(n2040), .Z(n4073) );
  XOR U3230 ( .A(in[1191]), .B(n4073), .Z(n2508) );
  XOR U3231 ( .A(in[1555]), .B(n4056), .Z(n2510) );
  OR U3232 ( .A(n2508), .B(n2510), .Z(n2041) );
  XNOR U3233 ( .A(n2220), .B(n2041), .Z(out[1299]) );
  XOR U3234 ( .A(in[666]), .B(n4256), .Z(n2858) );
  IV U3235 ( .A(n3138), .Z(n4080) );
  XOR U3236 ( .A(in[600]), .B(n4080), .Z(n3983) );
  XNOR U3237 ( .A(in[255]), .B(n3291), .Z(n3982) );
  NANDN U3238 ( .A(n3983), .B(n3982), .Z(n2042) );
  XNOR U3239 ( .A(n2858), .B(n2042), .Z(out[129]) );
  XNOR U3240 ( .A(in[202]), .B(n3946), .Z(n4339) );
  XOR U3241 ( .A(in[1422]), .B(n3199), .Z(n4340) );
  XNOR U3242 ( .A(in[1045]), .B(n4491), .Z(n2885) );
  NANDN U3243 ( .A(n4340), .B(n2885), .Z(n2043) );
  XNOR U3244 ( .A(n4339), .B(n2043), .Z(out[12]) );
  XOR U3245 ( .A(in[6]), .B(n3083), .Z(n2222) );
  IV U3246 ( .A(n2044), .Z(n4077) );
  XOR U3247 ( .A(in[1192]), .B(n4077), .Z(n2512) );
  XOR U3248 ( .A(in[1556]), .B(n4060), .Z(n2514) );
  OR U3249 ( .A(n2512), .B(n2514), .Z(n2045) );
  XNOR U3250 ( .A(n2222), .B(n2045), .Z(out[1300]) );
  XOR U3251 ( .A(in[7]), .B(n3085), .Z(n2224) );
  IV U3252 ( .A(n2046), .Z(n4081) );
  XOR U3253 ( .A(in[1193]), .B(n4081), .Z(n2516) );
  XOR U3254 ( .A(in[1557]), .B(n3128), .Z(n2121) );
  IV U3255 ( .A(n2121), .Z(n2518) );
  OR U3256 ( .A(n2516), .B(n2518), .Z(n2047) );
  XNOR U3257 ( .A(n2224), .B(n2047), .Z(out[1301]) );
  XOR U3258 ( .A(in[8]), .B(n4216), .Z(n2227) );
  IV U3259 ( .A(n2048), .Z(n4085) );
  XOR U3260 ( .A(in[1194]), .B(n4085), .Z(n2520) );
  XOR U3261 ( .A(in[1558]), .B(n3130), .Z(n2123) );
  IV U3262 ( .A(n2123), .Z(n2522) );
  OR U3263 ( .A(n2520), .B(n2522), .Z(n2049) );
  XNOR U3264 ( .A(n2227), .B(n2049), .Z(out[1302]) );
  XOR U3265 ( .A(in[9]), .B(n3088), .Z(n2229) );
  XOR U3266 ( .A(in[1559]), .B(n3132), .Z(n2125) );
  IV U3267 ( .A(n2125), .Z(n2526) );
  XOR U3268 ( .A(in[1195]), .B(n4090), .Z(n2524) );
  NANDN U3269 ( .A(n2526), .B(n2524), .Z(n2050) );
  XNOR U3270 ( .A(n2229), .B(n2050), .Z(out[1303]) );
  XOR U3271 ( .A(in[10]), .B(n3090), .Z(n2231) );
  XOR U3272 ( .A(in[1560]), .B(n4080), .Z(n2531) );
  XOR U3273 ( .A(in[1196]), .B(n4094), .Z(n2529) );
  NANDN U3274 ( .A(n2531), .B(n2529), .Z(n2051) );
  XNOR U3275 ( .A(n2231), .B(n2051), .Z(out[1304]) );
  XOR U3276 ( .A(in[11]), .B(n3092), .Z(n2233) );
  IV U3277 ( .A(n3140), .Z(n4084) );
  XOR U3278 ( .A(in[1561]), .B(n4084), .Z(n2535) );
  XOR U3279 ( .A(in[1197]), .B(n4098), .Z(n2533) );
  NANDN U3280 ( .A(n2535), .B(n2533), .Z(n2052) );
  XNOR U3281 ( .A(n2233), .B(n2052), .Z(out[1305]) );
  XOR U3282 ( .A(in[12]), .B(n3094), .Z(n2235) );
  IV U3283 ( .A(n3143), .Z(n4088) );
  XOR U3284 ( .A(in[1562]), .B(n4088), .Z(n2539) );
  XOR U3285 ( .A(in[1198]), .B(n4102), .Z(n2537) );
  NANDN U3286 ( .A(n2539), .B(n2537), .Z(n2053) );
  XNOR U3287 ( .A(n2235), .B(n2053), .Z(out[1306]) );
  XOR U3288 ( .A(in[13]), .B(n3098), .Z(n2237) );
  IV U3289 ( .A(n3145), .Z(n4092) );
  XOR U3290 ( .A(in[1563]), .B(n4092), .Z(n2543) );
  XOR U3291 ( .A(in[1199]), .B(n4106), .Z(n2541) );
  NANDN U3292 ( .A(n2543), .B(n2541), .Z(n2054) );
  XNOR U3293 ( .A(n2237), .B(n2054), .Z(out[1307]) );
  XOR U3294 ( .A(in[14]), .B(n4234), .Z(n2239) );
  IV U3295 ( .A(n3024), .Z(n4096) );
  XOR U3296 ( .A(in[1564]), .B(n4096), .Z(n2547) );
  XOR U3297 ( .A(in[1200]), .B(n4110), .Z(n2545) );
  NANDN U3298 ( .A(n2547), .B(n2545), .Z(n2055) );
  XNOR U3299 ( .A(n2239), .B(n2055), .Z(out[1308]) );
  XOR U3300 ( .A(in[15]), .B(n4237), .Z(n2241) );
  IV U3301 ( .A(n3026), .Z(n4100) );
  XOR U3302 ( .A(in[1565]), .B(n4100), .Z(n2551) );
  XOR U3303 ( .A(in[1201]), .B(n4118), .Z(n2549) );
  NANDN U3304 ( .A(n2551), .B(n2549), .Z(n2056) );
  XNOR U3305 ( .A(n2241), .B(n2056), .Z(out[1309]) );
  XOR U3306 ( .A(in[667]), .B(n4257), .Z(n2744) );
  IV U3307 ( .A(n2744), .Z(n2860) );
  XOR U3308 ( .A(in[601]), .B(n4084), .Z(n4027) );
  XNOR U3309 ( .A(in[192]), .B(n3294), .Z(n4024) );
  NANDN U3310 ( .A(n4027), .B(n4024), .Z(n2057) );
  XOR U3311 ( .A(n2860), .B(n2057), .Z(out[130]) );
  XOR U3312 ( .A(in[16]), .B(n4240), .Z(n2243) );
  IV U3313 ( .A(n3028), .Z(n4104) );
  XOR U3314 ( .A(in[1566]), .B(n4104), .Z(n2555) );
  XOR U3315 ( .A(in[1202]), .B(n4122), .Z(n2553) );
  NANDN U3316 ( .A(n2555), .B(n2553), .Z(n2058) );
  XNOR U3317 ( .A(n2243), .B(n2058), .Z(out[1310]) );
  XOR U3318 ( .A(in[17]), .B(n4241), .Z(n2245) );
  IV U3319 ( .A(n3030), .Z(n4108) );
  XOR U3320 ( .A(in[1567]), .B(n4108), .Z(n2558) );
  XOR U3321 ( .A(in[1203]), .B(n4126), .Z(n2557) );
  NANDN U3322 ( .A(n2558), .B(n2557), .Z(n2059) );
  XNOR U3323 ( .A(n2245), .B(n2059), .Z(out[1311]) );
  XOR U3324 ( .A(in[18]), .B(n3104), .Z(n2248) );
  IV U3325 ( .A(n3032), .Z(n4116) );
  XOR U3326 ( .A(in[1568]), .B(n4116), .Z(n2564) );
  XOR U3327 ( .A(in[1204]), .B(n4130), .Z(n2562) );
  NANDN U3328 ( .A(n2564), .B(n2562), .Z(n2060) );
  XNOR U3329 ( .A(n2248), .B(n2060), .Z(out[1312]) );
  XOR U3330 ( .A(in[19]), .B(n3106), .Z(n2250) );
  XOR U3331 ( .A(in[1569]), .B(n3034), .Z(n2129) );
  IV U3332 ( .A(n2129), .Z(n2568) );
  XOR U3333 ( .A(in[1205]), .B(n4134), .Z(n2566) );
  NANDN U3334 ( .A(n2568), .B(n2566), .Z(n2061) );
  XNOR U3335 ( .A(n2250), .B(n2061), .Z(out[1313]) );
  XOR U3336 ( .A(in[20]), .B(n4248), .Z(n2252) );
  XNOR U3337 ( .A(in[1570]), .B(n4124), .Z(n2574) );
  XOR U3338 ( .A(in[1206]), .B(n4138), .Z(n2572) );
  NANDN U3339 ( .A(n2574), .B(n2572), .Z(n2062) );
  XNOR U3340 ( .A(n2252), .B(n2062), .Z(out[1314]) );
  XOR U3341 ( .A(in[21]), .B(n4251), .Z(n2254) );
  XOR U3342 ( .A(in[1571]), .B(n3037), .Z(n2131) );
  IV U3343 ( .A(n2131), .Z(n2578) );
  XOR U3344 ( .A(in[1207]), .B(n4142), .Z(n2576) );
  NANDN U3345 ( .A(n2578), .B(n2576), .Z(n2063) );
  XNOR U3346 ( .A(n2254), .B(n2063), .Z(out[1315]) );
  XOR U3347 ( .A(in[22]), .B(n4252), .Z(n2256) );
  XOR U3348 ( .A(in[1572]), .B(n3039), .Z(n2134) );
  IV U3349 ( .A(n2134), .Z(n2582) );
  XOR U3350 ( .A(in[1208]), .B(n4146), .Z(n2580) );
  NANDN U3351 ( .A(n2582), .B(n2580), .Z(n2064) );
  XNOR U3352 ( .A(n2256), .B(n2064), .Z(out[1316]) );
  XOR U3353 ( .A(in[23]), .B(n4253), .Z(n2258) );
  XNOR U3354 ( .A(in[1573]), .B(n4136), .Z(n2136) );
  IV U3355 ( .A(n2136), .Z(n2586) );
  XOR U3356 ( .A(in[1209]), .B(n4150), .Z(n2584) );
  NANDN U3357 ( .A(n2586), .B(n2584), .Z(n2065) );
  XNOR U3358 ( .A(n2258), .B(n2065), .Z(out[1317]) );
  XOR U3359 ( .A(in[24]), .B(n4254), .Z(n2260) );
  XNOR U3360 ( .A(in[1574]), .B(n4140), .Z(n2590) );
  XOR U3361 ( .A(in[1210]), .B(n4154), .Z(n2588) );
  NAND U3362 ( .A(n2590), .B(n2588), .Z(n2066) );
  XNOR U3363 ( .A(n2260), .B(n2066), .Z(out[1318]) );
  XOR U3364 ( .A(in[25]), .B(n4255), .Z(n2262) );
  XOR U3365 ( .A(in[1211]), .B(n4164), .Z(n2592) );
  XNOR U3366 ( .A(in[1575]), .B(n4144), .Z(n2139) );
  IV U3367 ( .A(n2139), .Z(n2594) );
  OR U3368 ( .A(n2592), .B(n2594), .Z(n2067) );
  XNOR U3369 ( .A(n2262), .B(n2067), .Z(out[1319]) );
  XOR U3370 ( .A(in[668]), .B(n4260), .Z(n2746) );
  IV U3371 ( .A(n2746), .Z(n2862) );
  XOR U3372 ( .A(in[602]), .B(n4088), .Z(n4071) );
  XNOR U3373 ( .A(in[193]), .B(n3297), .Z(n4068) );
  NANDN U3374 ( .A(n4071), .B(n4068), .Z(n2068) );
  XOR U3375 ( .A(n2862), .B(n2068), .Z(out[131]) );
  XOR U3376 ( .A(in[26]), .B(n4256), .Z(n2264) );
  XOR U3377 ( .A(in[1212]), .B(n4168), .Z(n2596) );
  XNOR U3378 ( .A(in[1576]), .B(n4148), .Z(n2141) );
  IV U3379 ( .A(n2141), .Z(n2598) );
  OR U3380 ( .A(n2596), .B(n2598), .Z(n2069) );
  XNOR U3381 ( .A(n2264), .B(n2069), .Z(out[1320]) );
  XOR U3382 ( .A(in[27]), .B(n4257), .Z(n2266) );
  XOR U3383 ( .A(in[1213]), .B(n4172), .Z(n2600) );
  XNOR U3384 ( .A(in[1577]), .B(n4152), .Z(n2143) );
  IV U3385 ( .A(n2143), .Z(n2602) );
  OR U3386 ( .A(n2600), .B(n2602), .Z(n2070) );
  XNOR U3387 ( .A(n2266), .B(n2070), .Z(out[1321]) );
  XOR U3388 ( .A(in[28]), .B(n4260), .Z(n2269) );
  XNOR U3389 ( .A(in[1578]), .B(n4162), .Z(n2145) );
  IV U3390 ( .A(n2145), .Z(n2606) );
  XOR U3391 ( .A(in[1214]), .B(n4176), .Z(n2604) );
  NANDN U3392 ( .A(n2606), .B(n2604), .Z(n2071) );
  XNOR U3393 ( .A(n2269), .B(n2071), .Z(out[1322]) );
  XOR U3394 ( .A(in[29]), .B(n4261), .Z(n2271) );
  XOR U3395 ( .A(in[1215]), .B(n3291), .Z(n2608) );
  XNOR U3396 ( .A(in[1579]), .B(n4166), .Z(n2147) );
  IV U3397 ( .A(n2147), .Z(n2610) );
  OR U3398 ( .A(n2608), .B(n2610), .Z(n2072) );
  XNOR U3399 ( .A(n2271), .B(n2072), .Z(out[1323]) );
  XOR U3400 ( .A(in[30]), .B(n4262), .Z(n2273) );
  XOR U3401 ( .A(in[1152]), .B(n3294), .Z(n2614) );
  XNOR U3402 ( .A(in[1580]), .B(n4170), .Z(n2149) );
  IV U3403 ( .A(n2149), .Z(n2616) );
  OR U3404 ( .A(n2614), .B(n2616), .Z(n2073) );
  XNOR U3405 ( .A(n2273), .B(n2073), .Z(out[1324]) );
  XOR U3406 ( .A(in[31]), .B(n4263), .Z(n2275) );
  XOR U3407 ( .A(in[1153]), .B(n3297), .Z(n2618) );
  XNOR U3408 ( .A(in[1581]), .B(n4174), .Z(n2151) );
  IV U3409 ( .A(n2151), .Z(n2620) );
  OR U3410 ( .A(n2618), .B(n2620), .Z(n2074) );
  XNOR U3411 ( .A(n2275), .B(n2074), .Z(out[1325]) );
  XOR U3412 ( .A(in[32]), .B(n4266), .Z(n2277) );
  XOR U3413 ( .A(in[1154]), .B(n3304), .Z(n2622) );
  XNOR U3414 ( .A(in[1582]), .B(n3898), .Z(n2154) );
  IV U3415 ( .A(n2154), .Z(n2624) );
  OR U3416 ( .A(n2622), .B(n2624), .Z(n2075) );
  XNOR U3417 ( .A(n2277), .B(n2075), .Z(out[1326]) );
  XOR U3418 ( .A(in[33]), .B(n4269), .Z(n2279) );
  XOR U3419 ( .A(in[1155]), .B(n3307), .Z(n2626) );
  XNOR U3420 ( .A(in[1583]), .B(n3902), .Z(n2156) );
  IV U3421 ( .A(n2156), .Z(n2628) );
  OR U3422 ( .A(n2626), .B(n2628), .Z(n2076) );
  XNOR U3423 ( .A(n2279), .B(n2076), .Z(out[1327]) );
  XOR U3424 ( .A(in[34]), .B(n4272), .Z(n2281) );
  XOR U3425 ( .A(in[1156]), .B(n3310), .Z(n2630) );
  XNOR U3426 ( .A(in[1584]), .B(n3906), .Z(n2158) );
  IV U3427 ( .A(n2158), .Z(n2632) );
  OR U3428 ( .A(n2630), .B(n2632), .Z(n2077) );
  XNOR U3429 ( .A(n2281), .B(n2077), .Z(out[1328]) );
  IV U3430 ( .A(n4275), .Z(n3142) );
  XOR U3431 ( .A(in[35]), .B(n3142), .Z(n2283) );
  XOR U3432 ( .A(in[1157]), .B(n3313), .Z(n2634) );
  XNOR U3433 ( .A(in[1585]), .B(n3910), .Z(n2160) );
  IV U3434 ( .A(n2160), .Z(n2636) );
  OR U3435 ( .A(n2634), .B(n2636), .Z(n2078) );
  XNOR U3436 ( .A(n2283), .B(n2078), .Z(out[1329]) );
  XOR U3437 ( .A(in[669]), .B(n4261), .Z(n2748) );
  IV U3438 ( .A(n2748), .Z(n2867) );
  XOR U3439 ( .A(in[603]), .B(n4092), .Z(n4115) );
  XNOR U3440 ( .A(in[194]), .B(n3304), .Z(n4112) );
  NANDN U3441 ( .A(n4115), .B(n4112), .Z(n2079) );
  XOR U3442 ( .A(n2867), .B(n2079), .Z(out[132]) );
  XOR U3443 ( .A(in[36]), .B(n4278), .Z(n2285) );
  XOR U3444 ( .A(in[1158]), .B(n3316), .Z(n2638) );
  XNOR U3445 ( .A(in[1586]), .B(n3914), .Z(n2162) );
  IV U3446 ( .A(n2162), .Z(n2640) );
  OR U3447 ( .A(n2638), .B(n2640), .Z(n2080) );
  XNOR U3448 ( .A(n2285), .B(n2080), .Z(out[1330]) );
  XOR U3449 ( .A(in[37]), .B(n4280), .Z(n2287) );
  XOR U3450 ( .A(in[1159]), .B(n3319), .Z(n2642) );
  XOR U3451 ( .A(in[1587]), .B(n2569), .Z(n2644) );
  OR U3452 ( .A(n2642), .B(n2644), .Z(n2081) );
  XNOR U3453 ( .A(n2287), .B(n2081), .Z(out[1331]) );
  XOR U3454 ( .A(in[38]), .B(n4286), .Z(n2290) );
  XOR U3455 ( .A(in[1160]), .B(n3935), .Z(n2646) );
  XOR U3456 ( .A(in[1588]), .B(n2611), .Z(n2648) );
  OR U3457 ( .A(n2646), .B(n2648), .Z(n2082) );
  XNOR U3458 ( .A(n2290), .B(n2082), .Z(out[1332]) );
  XOR U3459 ( .A(in[39]), .B(n4288), .Z(n2292) );
  XOR U3460 ( .A(in[1161]), .B(n3942), .Z(n2650) );
  XOR U3461 ( .A(in[1589]), .B(n2653), .Z(n2652) );
  OR U3462 ( .A(n2650), .B(n2652), .Z(n2083) );
  XNOR U3463 ( .A(n2292), .B(n2083), .Z(out[1333]) );
  XOR U3464 ( .A(in[40]), .B(n4290), .Z(n2295) );
  XOR U3465 ( .A(in[1162]), .B(n3946), .Z(n2656) );
  XNOR U3466 ( .A(in[1590]), .B(n3065), .Z(n2658) );
  NANDN U3467 ( .A(n2656), .B(n2658), .Z(n2084) );
  XNOR U3468 ( .A(n2295), .B(n2084), .Z(out[1334]) );
  XOR U3469 ( .A(in[41]), .B(n4292), .Z(n2297) );
  XOR U3470 ( .A(in[1163]), .B(n3950), .Z(n2660) );
  XNOR U3471 ( .A(in[1591]), .B(n3067), .Z(n2662) );
  NANDN U3472 ( .A(n2660), .B(n2662), .Z(n2085) );
  XNOR U3473 ( .A(n2297), .B(n2085), .Z(out[1335]) );
  XOR U3474 ( .A(in[42]), .B(n4294), .Z(n2299) );
  XOR U3475 ( .A(in[1164]), .B(n3954), .Z(n2664) );
  XNOR U3476 ( .A(in[1592]), .B(n3070), .Z(n2666) );
  NANDN U3477 ( .A(n2664), .B(n2666), .Z(n2086) );
  XNOR U3478 ( .A(n2299), .B(n2086), .Z(out[1336]) );
  XOR U3479 ( .A(in[43]), .B(n4296), .Z(n2301) );
  XOR U3480 ( .A(in[1165]), .B(n3958), .Z(n2668) );
  XOR U3481 ( .A(in[1593]), .B(n2700), .Z(n2670) );
  OR U3482 ( .A(n2668), .B(n2670), .Z(n2087) );
  XNOR U3483 ( .A(n2301), .B(n2087), .Z(out[1337]) );
  XOR U3484 ( .A(in[44]), .B(n4298), .Z(n2303) );
  XOR U3485 ( .A(in[1166]), .B(n3962), .Z(n2672) );
  XOR U3486 ( .A(in[1594]), .B(n2702), .Z(n2674) );
  OR U3487 ( .A(n2672), .B(n2674), .Z(n2088) );
  XNOR U3488 ( .A(n2303), .B(n2088), .Z(out[1338]) );
  XOR U3489 ( .A(in[45]), .B(n4300), .Z(n2305) );
  XOR U3490 ( .A(in[1167]), .B(n3966), .Z(n2676) );
  XNOR U3491 ( .A(in[1595]), .B(n3953), .Z(n2169) );
  IV U3492 ( .A(n2169), .Z(n2678) );
  OR U3493 ( .A(n2676), .B(n2678), .Z(n2089) );
  XNOR U3494 ( .A(n2305), .B(n2089), .Z(out[1339]) );
  XOR U3495 ( .A(in[670]), .B(n4262), .Z(n2750) );
  IV U3496 ( .A(n2750), .Z(n2869) );
  XOR U3497 ( .A(in[604]), .B(n4096), .Z(n4159) );
  XNOR U3498 ( .A(in[195]), .B(n3307), .Z(n4156) );
  NANDN U3499 ( .A(n4159), .B(n4156), .Z(n2090) );
  XOR U3500 ( .A(n2869), .B(n2090), .Z(out[133]) );
  XOR U3501 ( .A(in[46]), .B(n4302), .Z(n2307) );
  XOR U3502 ( .A(in[1168]), .B(n3970), .Z(n2680) );
  XNOR U3503 ( .A(in[1596]), .B(n3957), .Z(n2171) );
  IV U3504 ( .A(n2171), .Z(n2682) );
  OR U3505 ( .A(n2680), .B(n2682), .Z(n2091) );
  XNOR U3506 ( .A(n2307), .B(n2091), .Z(out[1340]) );
  XOR U3507 ( .A(in[47]), .B(n4304), .Z(n2309) );
  XOR U3508 ( .A(in[1169]), .B(n3974), .Z(n2684) );
  XNOR U3509 ( .A(in[1597]), .B(n3961), .Z(n2173) );
  IV U3510 ( .A(n2173), .Z(n2686) );
  OR U3511 ( .A(n2684), .B(n2686), .Z(n2092) );
  XNOR U3512 ( .A(n2309), .B(n2092), .Z(out[1341]) );
  XOR U3513 ( .A(in[48]), .B(n4311), .Z(n2312) );
  XOR U3514 ( .A(in[1170]), .B(n3978), .Z(n2688) );
  XNOR U3515 ( .A(in[1598]), .B(n3965), .Z(n2175) );
  IV U3516 ( .A(n2175), .Z(n2690) );
  OR U3517 ( .A(n2688), .B(n2690), .Z(n2093) );
  XNOR U3518 ( .A(n2312), .B(n2093), .Z(out[1342]) );
  XOR U3519 ( .A(in[49]), .B(n4314), .Z(n2314) );
  IV U3520 ( .A(n3985), .Z(n3349) );
  XOR U3521 ( .A(in[1171]), .B(n3349), .Z(n2692) );
  XNOR U3522 ( .A(in[1599]), .B(n3969), .Z(n2177) );
  IV U3523 ( .A(n2177), .Z(n2693) );
  OR U3524 ( .A(n2692), .B(n2693), .Z(n2094) );
  XNOR U3525 ( .A(n2314), .B(n2094), .Z(out[1343]) );
  XNOR U3526 ( .A(in[427]), .B(n4347), .Z(n2316) );
  NOR U3527 ( .A(n2436), .B(n2179), .Z(n2095) );
  XNOR U3528 ( .A(n2316), .B(n2095), .Z(out[1344]) );
  XNOR U3529 ( .A(in[428]), .B(n4350), .Z(n2318) );
  NOR U3530 ( .A(n2096), .B(n2181), .Z(n2097) );
  XNOR U3531 ( .A(n2318), .B(n2097), .Z(out[1345]) );
  XNOR U3532 ( .A(in[429]), .B(n4353), .Z(n2320) );
  NOR U3533 ( .A(n2098), .B(n2184), .Z(n2099) );
  XNOR U3534 ( .A(n2320), .B(n2099), .Z(out[1346]) );
  XNOR U3535 ( .A(in[430]), .B(n4356), .Z(n2322) );
  NOR U3536 ( .A(n2448), .B(n2186), .Z(n2100) );
  XNOR U3537 ( .A(n2322), .B(n2100), .Z(out[1347]) );
  XNOR U3538 ( .A(in[431]), .B(n4358), .Z(n2324) );
  NOR U3539 ( .A(n2452), .B(n2188), .Z(n2101) );
  XNOR U3540 ( .A(n2324), .B(n2101), .Z(out[1348]) );
  XNOR U3541 ( .A(in[432]), .B(n4361), .Z(n2326) );
  NOR U3542 ( .A(n2455), .B(n2190), .Z(n2102) );
  XNOR U3543 ( .A(n2326), .B(n2102), .Z(out[1349]) );
  XOR U3544 ( .A(in[671]), .B(n4263), .Z(n2752) );
  IV U3545 ( .A(n2752), .Z(n2871) );
  XOR U3546 ( .A(in[605]), .B(n4100), .Z(n4197) );
  XNOR U3547 ( .A(in[196]), .B(n3310), .Z(n4194) );
  NANDN U3548 ( .A(n4197), .B(n4194), .Z(n2103) );
  XOR U3549 ( .A(n2871), .B(n2103), .Z(out[134]) );
  XNOR U3550 ( .A(in[433]), .B(n4364), .Z(n2328) );
  NOR U3551 ( .A(n2104), .B(n2192), .Z(n2105) );
  XNOR U3552 ( .A(n2328), .B(n2105), .Z(out[1350]) );
  XNOR U3553 ( .A(in[434]), .B(n4367), .Z(n2330) );
  NOR U3554 ( .A(n2106), .B(n2194), .Z(n2107) );
  XNOR U3555 ( .A(n2330), .B(n2107), .Z(out[1351]) );
  XNOR U3556 ( .A(in[435]), .B(n4374), .Z(n2333) );
  NOR U3557 ( .A(n2467), .B(n2196), .Z(n2108) );
  XNOR U3558 ( .A(n2333), .B(n2108), .Z(out[1352]) );
  XNOR U3559 ( .A(in[436]), .B(n4377), .Z(n2336) );
  NOR U3560 ( .A(n2470), .B(n2198), .Z(n2109) );
  XNOR U3561 ( .A(n2336), .B(n2109), .Z(out[1353]) );
  XNOR U3562 ( .A(in[437]), .B(n4380), .Z(n2339) );
  NOR U3563 ( .A(n2473), .B(n2200), .Z(n2110) );
  XNOR U3564 ( .A(n2339), .B(n2110), .Z(out[1354]) );
  XNOR U3565 ( .A(in[438]), .B(n4383), .Z(n2342) );
  NOR U3566 ( .A(n2476), .B(n2202), .Z(n2111) );
  XNOR U3567 ( .A(n2342), .B(n2111), .Z(out[1355]) );
  XNOR U3568 ( .A(in[439]), .B(n4386), .Z(n2345) );
  NOR U3569 ( .A(n2479), .B(n2205), .Z(n2112) );
  XNOR U3570 ( .A(n2345), .B(n2112), .Z(out[1356]) );
  XNOR U3571 ( .A(in[440]), .B(n4388), .Z(n2348) );
  NOR U3572 ( .A(n2482), .B(n2207), .Z(n2113) );
  XNOR U3573 ( .A(n2348), .B(n2113), .Z(out[1357]) );
  XNOR U3574 ( .A(in[441]), .B(n4391), .Z(n2351) );
  NOR U3575 ( .A(n2114), .B(n2209), .Z(n2115) );
  XNOR U3576 ( .A(n2351), .B(n2115), .Z(out[1358]) );
  XOR U3577 ( .A(in[442]), .B(n2116), .Z(n2353) );
  XOR U3578 ( .A(in[672]), .B(n4266), .Z(n2754) );
  IV U3579 ( .A(n2754), .Z(n2873) );
  XOR U3580 ( .A(in[606]), .B(n4104), .Z(n4215) );
  XNOR U3581 ( .A(in[197]), .B(n3313), .Z(n4444) );
  NANDN U3582 ( .A(n4215), .B(n4444), .Z(n2117) );
  XOR U3583 ( .A(n2873), .B(n2117), .Z(out[135]) );
  XOR U3584 ( .A(in[443]), .B(n2118), .Z(n2355) );
  XNOR U3585 ( .A(in[444]), .B(n4400), .Z(n2356) );
  XNOR U3586 ( .A(in[445]), .B(n4407), .Z(n2359) );
  NOR U3587 ( .A(n2119), .B(n2218), .Z(n2120) );
  XNOR U3588 ( .A(n2359), .B(n2120), .Z(out[1362]) );
  XNOR U3589 ( .A(in[446]), .B(n4410), .Z(n2361) );
  XNOR U3590 ( .A(in[447]), .B(n4413), .Z(n2363) );
  XNOR U3591 ( .A(in[384]), .B(n4416), .Z(n2365) );
  NOR U3592 ( .A(n2121), .B(n2224), .Z(n2122) );
  XNOR U3593 ( .A(n2365), .B(n2122), .Z(out[1365]) );
  XNOR U3594 ( .A(in[385]), .B(n4419), .Z(n2367) );
  NOR U3595 ( .A(n2123), .B(n2227), .Z(n2124) );
  XNOR U3596 ( .A(n2367), .B(n2124), .Z(out[1366]) );
  XNOR U3597 ( .A(in[386]), .B(n4422), .Z(n2369) );
  NOR U3598 ( .A(n2125), .B(n2229), .Z(n2126) );
  XNOR U3599 ( .A(n2369), .B(n2126), .Z(out[1367]) );
  XNOR U3600 ( .A(in[387]), .B(n4425), .Z(n2371) );
  XNOR U3601 ( .A(in[388]), .B(n4428), .Z(n2373) );
  XOR U3602 ( .A(in[673]), .B(n4269), .Z(n2761) );
  IV U3603 ( .A(n2761), .Z(n2875) );
  XOR U3604 ( .A(in[607]), .B(n4108), .Z(n4243) );
  XNOR U3605 ( .A(in[198]), .B(n3316), .Z(n4731) );
  NANDN U3606 ( .A(n4243), .B(n4731), .Z(n2127) );
  XOR U3607 ( .A(n2875), .B(n2127), .Z(out[136]) );
  XNOR U3608 ( .A(in[389]), .B(n4431), .Z(n2375) );
  XOR U3609 ( .A(in[390]), .B(n2128), .Z(n2377) );
  XNOR U3610 ( .A(in[391]), .B(n4445), .Z(n2380) );
  XNOR U3611 ( .A(in[392]), .B(n4448), .Z(n2382) );
  XNOR U3612 ( .A(in[393]), .B(n4451), .Z(n2384) );
  XNOR U3613 ( .A(in[394]), .B(n4454), .Z(n2386) );
  XNOR U3614 ( .A(in[395]), .B(n4457), .Z(n2388) );
  XNOR U3615 ( .A(n4460), .B(in[396]), .Z(n2390) );
  NOR U3616 ( .A(n2129), .B(n2250), .Z(n2130) );
  XOR U3617 ( .A(n2390), .B(n2130), .Z(out[1377]) );
  XNOR U3618 ( .A(n4463), .B(in[397]), .Z(n2391) );
  XNOR U3619 ( .A(n4466), .B(in[398]), .Z(n2392) );
  NOR U3620 ( .A(n2131), .B(n2254), .Z(n2132) );
  XOR U3621 ( .A(n2392), .B(n2132), .Z(out[1379]) );
  XOR U3622 ( .A(in[674]), .B(n4272), .Z(n2763) );
  IV U3623 ( .A(n2763), .Z(n2877) );
  XOR U3624 ( .A(in[608]), .B(n4116), .Z(n4259) );
  XNOR U3625 ( .A(in[199]), .B(n3319), .Z(n5162) );
  NANDN U3626 ( .A(n4259), .B(n5162), .Z(n2133) );
  XOR U3627 ( .A(n2877), .B(n2133), .Z(out[137]) );
  XNOR U3628 ( .A(n4469), .B(in[399]), .Z(n2393) );
  NOR U3629 ( .A(n2134), .B(n2256), .Z(n2135) );
  XOR U3630 ( .A(n2393), .B(n2135), .Z(out[1380]) );
  XNOR U3631 ( .A(n4472), .B(in[400]), .Z(n2394) );
  NOR U3632 ( .A(n2136), .B(n2258), .Z(n2137) );
  XOR U3633 ( .A(n2394), .B(n2137), .Z(out[1381]) );
  XNOR U3634 ( .A(n4479), .B(in[401]), .Z(n2396) );
  NOR U3635 ( .A(n2590), .B(n2260), .Z(n2138) );
  XOR U3636 ( .A(n2396), .B(n2138), .Z(out[1382]) );
  XNOR U3637 ( .A(n4482), .B(in[402]), .Z(n2397) );
  NOR U3638 ( .A(n2139), .B(n2262), .Z(n2140) );
  XOR U3639 ( .A(n2397), .B(n2140), .Z(out[1383]) );
  XNOR U3640 ( .A(n4485), .B(in[403]), .Z(n2398) );
  NOR U3641 ( .A(n2141), .B(n2264), .Z(n2142) );
  XOR U3642 ( .A(n2398), .B(n2142), .Z(out[1384]) );
  XNOR U3643 ( .A(in[404]), .B(n4488), .Z(n2399) );
  NOR U3644 ( .A(n2143), .B(n2266), .Z(n2144) );
  XOR U3645 ( .A(n2399), .B(n2144), .Z(out[1385]) );
  XNOR U3646 ( .A(in[405]), .B(n4491), .Z(n2400) );
  NOR U3647 ( .A(n2145), .B(n2269), .Z(n2146) );
  XOR U3648 ( .A(n2400), .B(n2146), .Z(out[1386]) );
  XNOR U3649 ( .A(in[406]), .B(n4494), .Z(n2401) );
  NOR U3650 ( .A(n2147), .B(n2271), .Z(n2148) );
  XOR U3651 ( .A(n2401), .B(n2148), .Z(out[1387]) );
  XNOR U3652 ( .A(in[407]), .B(n4497), .Z(n2402) );
  NOR U3653 ( .A(n2149), .B(n2273), .Z(n2150) );
  XOR U3654 ( .A(n2402), .B(n2150), .Z(out[1388]) );
  XNOR U3655 ( .A(in[408]), .B(n4500), .Z(n2403) );
  NOR U3656 ( .A(n2151), .B(n2275), .Z(n2152) );
  XOR U3657 ( .A(n2403), .B(n2152), .Z(out[1389]) );
  XOR U3658 ( .A(in[675]), .B(n4275), .Z(n2880) );
  IV U3659 ( .A(n3034), .Z(n4120) );
  XOR U3660 ( .A(in[609]), .B(n4120), .Z(n4285) );
  NANDN U3661 ( .A(n4285), .B(n4282), .Z(n2153) );
  XOR U3662 ( .A(n2880), .B(n2153), .Z(out[138]) );
  XNOR U3663 ( .A(in[409]), .B(n4503), .Z(n2404) );
  NOR U3664 ( .A(n2154), .B(n2277), .Z(n2155) );
  XOR U3665 ( .A(n2404), .B(n2155), .Z(out[1390]) );
  XNOR U3666 ( .A(in[410]), .B(n4506), .Z(n2405) );
  NOR U3667 ( .A(n2156), .B(n2279), .Z(n2157) );
  XOR U3668 ( .A(n2405), .B(n2157), .Z(out[1391]) );
  XOR U3669 ( .A(in[411]), .B(n4513), .Z(n2407) );
  NOR U3670 ( .A(n2158), .B(n2281), .Z(n2159) );
  XOR U3671 ( .A(n2407), .B(n2159), .Z(out[1392]) );
  XOR U3672 ( .A(in[412]), .B(n4516), .Z(n2408) );
  NOR U3673 ( .A(n2160), .B(n2283), .Z(n2161) );
  XOR U3674 ( .A(n2408), .B(n2161), .Z(out[1393]) );
  XOR U3675 ( .A(in[413]), .B(n4519), .Z(n2409) );
  NOR U3676 ( .A(n2162), .B(n2285), .Z(n2163) );
  XOR U3677 ( .A(n2409), .B(n2163), .Z(out[1394]) );
  XOR U3678 ( .A(in[414]), .B(n4522), .Z(n2410) );
  XOR U3679 ( .A(in[415]), .B(n4526), .Z(n2412) );
  XOR U3680 ( .A(in[416]), .B(n4530), .Z(n2414) );
  XNOR U3681 ( .A(in[417]), .B(n4534), .Z(n2416) );
  NOR U3682 ( .A(n2658), .B(n2295), .Z(n2164) );
  XOR U3683 ( .A(n2416), .B(n2164), .Z(out[1398]) );
  XNOR U3684 ( .A(in[418]), .B(n4538), .Z(n2417) );
  NOR U3685 ( .A(n2662), .B(n2297), .Z(n2165) );
  XOR U3686 ( .A(n2417), .B(n2165), .Z(out[1399]) );
  XOR U3687 ( .A(in[676]), .B(n4278), .Z(n2882) );
  XNOR U3688 ( .A(in[610]), .B(n4124), .Z(n4310) );
  NANDN U3689 ( .A(n4310), .B(n4307), .Z(n2166) );
  XNOR U3690 ( .A(n2882), .B(n2166), .Z(out[139]) );
  XNOR U3691 ( .A(in[203]), .B(n3950), .Z(n4370) );
  XOR U3692 ( .A(in[1423]), .B(n3202), .Z(n4371) );
  XNOR U3693 ( .A(in[1046]), .B(n4494), .Z(n2887) );
  NANDN U3694 ( .A(n4371), .B(n2887), .Z(n2167) );
  XNOR U3695 ( .A(n4370), .B(n2167), .Z(out[13]) );
  XNOR U3696 ( .A(in[419]), .B(n4542), .Z(n2418) );
  NOR U3697 ( .A(n2666), .B(n2299), .Z(n2168) );
  XOR U3698 ( .A(n2418), .B(n2168), .Z(out[1400]) );
  XNOR U3699 ( .A(in[420]), .B(n4546), .Z(n2419) );
  XNOR U3700 ( .A(in[421]), .B(n4552), .Z(n2422) );
  XNOR U3701 ( .A(in[422]), .B(n4554), .Z(n2424) );
  NOR U3702 ( .A(n2169), .B(n2305), .Z(n2170) );
  XNOR U3703 ( .A(n2424), .B(n2170), .Z(out[1403]) );
  XNOR U3704 ( .A(in[423]), .B(n4335), .Z(n2426) );
  NOR U3705 ( .A(n2171), .B(n2307), .Z(n2172) );
  XNOR U3706 ( .A(n2426), .B(n2172), .Z(out[1404]) );
  XNOR U3707 ( .A(in[424]), .B(n4337), .Z(n2428) );
  NOR U3708 ( .A(n2173), .B(n2309), .Z(n2174) );
  XNOR U3709 ( .A(n2428), .B(n2174), .Z(out[1405]) );
  XNOR U3710 ( .A(in[425]), .B(n4343), .Z(n2430) );
  NOR U3711 ( .A(n2175), .B(n2312), .Z(n2176) );
  XNOR U3712 ( .A(n2430), .B(n2176), .Z(out[1406]) );
  XNOR U3713 ( .A(in[426]), .B(n4345), .Z(n2432) );
  NOR U3714 ( .A(n2177), .B(n2314), .Z(n2178) );
  XNOR U3715 ( .A(n2432), .B(n2178), .Z(out[1407]) );
  XOR U3716 ( .A(in[789]), .B(n4014), .Z(n2434) );
  NAND U3717 ( .A(n2179), .B(n2316), .Z(n2180) );
  XOR U3718 ( .A(n2434), .B(n2180), .Z(out[1408]) );
  IV U3719 ( .A(n2773), .Z(n4018) );
  XOR U3720 ( .A(in[790]), .B(n4018), .Z(n2437) );
  NAND U3721 ( .A(n2181), .B(n2318), .Z(n2182) );
  XOR U3722 ( .A(n2437), .B(n2182), .Z(out[1409]) );
  XOR U3723 ( .A(in[677]), .B(n4280), .Z(n2884) );
  IV U3724 ( .A(n3037), .Z(n4128) );
  XOR U3725 ( .A(in[611]), .B(n4128), .Z(n4342) );
  NANDN U3726 ( .A(n4342), .B(n4339), .Z(n2183) );
  XNOR U3727 ( .A(n2884), .B(n2183), .Z(out[140]) );
  IV U3728 ( .A(n2780), .Z(n4022) );
  XOR U3729 ( .A(in[791]), .B(n4022), .Z(n2442) );
  NAND U3730 ( .A(n2184), .B(n2320), .Z(n2185) );
  XOR U3731 ( .A(n2442), .B(n2185), .Z(out[1410]) );
  IV U3732 ( .A(n2794), .Z(n4030) );
  XOR U3733 ( .A(in[792]), .B(n4030), .Z(n2446) );
  NAND U3734 ( .A(n2186), .B(n2322), .Z(n2187) );
  XOR U3735 ( .A(n2446), .B(n2187), .Z(out[1411]) );
  IV U3736 ( .A(n2817), .Z(n4034) );
  XOR U3737 ( .A(in[793]), .B(n4034), .Z(n2453) );
  NAND U3738 ( .A(n2188), .B(n2324), .Z(n2189) );
  XOR U3739 ( .A(n2453), .B(n2189), .Z(out[1412]) );
  IV U3740 ( .A(n2840), .Z(n4038) );
  XOR U3741 ( .A(in[794]), .B(n4038), .Z(n2456) );
  NAND U3742 ( .A(n2190), .B(n2326), .Z(n2191) );
  XOR U3743 ( .A(n2456), .B(n2191), .Z(out[1413]) );
  IV U3744 ( .A(n2864), .Z(n4042) );
  XOR U3745 ( .A(in[795]), .B(n4042), .Z(n2458) );
  NAND U3746 ( .A(n2192), .B(n2328), .Z(n2193) );
  XOR U3747 ( .A(n2458), .B(n2193), .Z(out[1414]) );
  IV U3748 ( .A(n2888), .Z(n4046) );
  XOR U3749 ( .A(in[796]), .B(n4046), .Z(n2462) );
  NAND U3750 ( .A(n2194), .B(n2330), .Z(n2195) );
  XOR U3751 ( .A(n2462), .B(n2195), .Z(out[1415]) );
  IV U3752 ( .A(n2921), .Z(n4050) );
  XOR U3753 ( .A(in[797]), .B(n4050), .Z(n2468) );
  NAND U3754 ( .A(n2196), .B(n2333), .Z(n2197) );
  XOR U3755 ( .A(n2468), .B(n2197), .Z(out[1416]) );
  XOR U3756 ( .A(in[798]), .B(n4054), .Z(n2335) );
  NAND U3757 ( .A(n2198), .B(n2336), .Z(n2199) );
  XNOR U3758 ( .A(n2335), .B(n2199), .Z(out[1417]) );
  XOR U3759 ( .A(in[799]), .B(n4058), .Z(n2338) );
  NAND U3760 ( .A(n2200), .B(n2339), .Z(n2201) );
  XNOR U3761 ( .A(n2338), .B(n2201), .Z(out[1418]) );
  XOR U3762 ( .A(in[800]), .B(n4062), .Z(n2341) );
  NAND U3763 ( .A(n2202), .B(n2342), .Z(n2203) );
  XNOR U3764 ( .A(n2341), .B(n2203), .Z(out[1419]) );
  XOR U3765 ( .A(in[678]), .B(n4286), .Z(n2886) );
  IV U3766 ( .A(n3039), .Z(n4132) );
  XOR U3767 ( .A(in[612]), .B(n4132), .Z(n4373) );
  NANDN U3768 ( .A(n4373), .B(n4370), .Z(n2204) );
  XNOR U3769 ( .A(n2886), .B(n2204), .Z(out[141]) );
  XOR U3770 ( .A(in[801]), .B(n4066), .Z(n2344) );
  NAND U3771 ( .A(n2205), .B(n2345), .Z(n2206) );
  XNOR U3772 ( .A(n2344), .B(n2206), .Z(out[1420]) );
  XOR U3773 ( .A(in[802]), .B(n4074), .Z(n2347) );
  NAND U3774 ( .A(n2207), .B(n2348), .Z(n2208) );
  XNOR U3775 ( .A(n2347), .B(n2208), .Z(out[1421]) );
  XOR U3776 ( .A(in[803]), .B(n4078), .Z(n2350) );
  NAND U3777 ( .A(n2209), .B(n2351), .Z(n2210) );
  XNOR U3778 ( .A(n2350), .B(n2210), .Z(out[1422]) );
  XOR U3779 ( .A(in[804]), .B(n4082), .Z(n2354) );
  NANDN U3780 ( .A(n2353), .B(n2211), .Z(n2212) );
  XNOR U3781 ( .A(n2354), .B(n2212), .Z(out[1423]) );
  IV U3782 ( .A(n2213), .Z(n4086) );
  XOR U3783 ( .A(in[805]), .B(n4086), .Z(n2495) );
  NANDN U3784 ( .A(n2355), .B(n2214), .Z(n2215) );
  XOR U3785 ( .A(n2495), .B(n2215), .Z(out[1424]) );
  XNOR U3786 ( .A(in[806]), .B(n4089), .Z(n2499) );
  NAND U3787 ( .A(n2216), .B(n2356), .Z(n2217) );
  XNOR U3788 ( .A(n2499), .B(n2217), .Z(out[1425]) );
  XNOR U3789 ( .A(in[807]), .B(n4093), .Z(n2503) );
  NAND U3790 ( .A(n2218), .B(n2359), .Z(n2219) );
  XNOR U3791 ( .A(n2503), .B(n2219), .Z(out[1426]) );
  XNOR U3792 ( .A(in[808]), .B(n4097), .Z(n2507) );
  NAND U3793 ( .A(n2220), .B(n2361), .Z(n2221) );
  XNOR U3794 ( .A(n2507), .B(n2221), .Z(out[1427]) );
  XNOR U3795 ( .A(in[809]), .B(n4101), .Z(n2511) );
  NAND U3796 ( .A(n2222), .B(n2363), .Z(n2223) );
  XNOR U3797 ( .A(n2511), .B(n2223), .Z(out[1428]) );
  XNOR U3798 ( .A(in[810]), .B(n4105), .Z(n2515) );
  NAND U3799 ( .A(n2224), .B(n2365), .Z(n2225) );
  XNOR U3800 ( .A(n2515), .B(n2225), .Z(out[1429]) );
  XOR U3801 ( .A(in[679]), .B(n4288), .Z(n2769) );
  XOR U3802 ( .A(in[613]), .B(n4136), .Z(n4406) );
  XNOR U3803 ( .A(in[204]), .B(n3954), .Z(n4403) );
  NANDN U3804 ( .A(n4406), .B(n4403), .Z(n2226) );
  XNOR U3805 ( .A(n2769), .B(n2226), .Z(out[142]) );
  XNOR U3806 ( .A(in[811]), .B(n4109), .Z(n2519) );
  NAND U3807 ( .A(n2227), .B(n2367), .Z(n2228) );
  XOR U3808 ( .A(n2519), .B(n2228), .Z(out[1430]) );
  XNOR U3809 ( .A(in[812]), .B(n4117), .Z(n2523) );
  NAND U3810 ( .A(n2229), .B(n2369), .Z(n2230) );
  XOR U3811 ( .A(n2523), .B(n2230), .Z(out[1431]) );
  XOR U3812 ( .A(in[813]), .B(n4121), .Z(n2528) );
  NAND U3813 ( .A(n2231), .B(n2371), .Z(n2232) );
  XOR U3814 ( .A(n2528), .B(n2232), .Z(out[1432]) );
  XOR U3815 ( .A(in[814]), .B(n4125), .Z(n2532) );
  NAND U3816 ( .A(n2233), .B(n2373), .Z(n2234) );
  XOR U3817 ( .A(n2532), .B(n2234), .Z(out[1433]) );
  XOR U3818 ( .A(in[815]), .B(n4129), .Z(n2536) );
  NAND U3819 ( .A(n2235), .B(n2375), .Z(n2236) );
  XOR U3820 ( .A(n2536), .B(n2236), .Z(out[1434]) );
  XOR U3821 ( .A(in[816]), .B(n4133), .Z(n2540) );
  NANDN U3822 ( .A(n2377), .B(n2237), .Z(n2238) );
  XOR U3823 ( .A(n2540), .B(n2238), .Z(out[1435]) );
  XOR U3824 ( .A(in[817]), .B(n4137), .Z(n2544) );
  NAND U3825 ( .A(n2239), .B(n2380), .Z(n2240) );
  XOR U3826 ( .A(n2544), .B(n2240), .Z(out[1436]) );
  XOR U3827 ( .A(in[818]), .B(n4141), .Z(n2548) );
  NAND U3828 ( .A(n2241), .B(n2382), .Z(n2242) );
  XOR U3829 ( .A(n2548), .B(n2242), .Z(out[1437]) );
  XOR U3830 ( .A(in[819]), .B(n4145), .Z(n2552) );
  NAND U3831 ( .A(n2243), .B(n2384), .Z(n2244) );
  XOR U3832 ( .A(n2552), .B(n2244), .Z(out[1438]) );
  XOR U3833 ( .A(in[820]), .B(n4149), .Z(n2556) );
  NAND U3834 ( .A(n2245), .B(n2386), .Z(n2246) );
  XOR U3835 ( .A(n2556), .B(n2246), .Z(out[1439]) );
  XOR U3836 ( .A(in[680]), .B(n4290), .Z(n2770) );
  XOR U3837 ( .A(in[614]), .B(n4140), .Z(n4440) );
  XNOR U3838 ( .A(in[205]), .B(n3958), .Z(n4437) );
  NANDN U3839 ( .A(n4440), .B(n4437), .Z(n2247) );
  XNOR U3840 ( .A(n2770), .B(n2247), .Z(out[143]) );
  XNOR U3841 ( .A(in[821]), .B(n4153), .Z(n2561) );
  NAND U3842 ( .A(n2248), .B(n2388), .Z(n2249) );
  XOR U3843 ( .A(n2561), .B(n2249), .Z(out[1440]) );
  XNOR U3844 ( .A(in[822]), .B(n4163), .Z(n2565) );
  NANDN U3845 ( .A(n2390), .B(n2250), .Z(n2251) );
  XOR U3846 ( .A(n2565), .B(n2251), .Z(out[1441]) );
  XNOR U3847 ( .A(in[823]), .B(n4167), .Z(n2571) );
  NANDN U3848 ( .A(n2391), .B(n2252), .Z(n2253) );
  XOR U3849 ( .A(n2571), .B(n2253), .Z(out[1442]) );
  XNOR U3850 ( .A(in[824]), .B(n4171), .Z(n2575) );
  NANDN U3851 ( .A(n2392), .B(n2254), .Z(n2255) );
  XOR U3852 ( .A(n2575), .B(n2255), .Z(out[1443]) );
  XNOR U3853 ( .A(in[825]), .B(n4175), .Z(n2579) );
  NANDN U3854 ( .A(n2393), .B(n2256), .Z(n2257) );
  XOR U3855 ( .A(n2579), .B(n2257), .Z(out[1444]) );
  XOR U3856 ( .A(in[826]), .B(n3899), .Z(n2583) );
  NANDN U3857 ( .A(n2394), .B(n2258), .Z(n2259) );
  XOR U3858 ( .A(n2583), .B(n2259), .Z(out[1445]) );
  XOR U3859 ( .A(in[827]), .B(n3903), .Z(n2587) );
  NANDN U3860 ( .A(n2396), .B(n2260), .Z(n2261) );
  XOR U3861 ( .A(n2587), .B(n2261), .Z(out[1446]) );
  XOR U3862 ( .A(in[828]), .B(n3907), .Z(n2591) );
  NANDN U3863 ( .A(n2397), .B(n2262), .Z(n2263) );
  XOR U3864 ( .A(n2591), .B(n2263), .Z(out[1447]) );
  XOR U3865 ( .A(in[829]), .B(n3911), .Z(n2595) );
  NANDN U3866 ( .A(n2398), .B(n2264), .Z(n2265) );
  XOR U3867 ( .A(n2595), .B(n2265), .Z(out[1448]) );
  XOR U3868 ( .A(in[830]), .B(n3915), .Z(n2599) );
  NANDN U3869 ( .A(n2399), .B(n2266), .Z(n2267) );
  XOR U3870 ( .A(n2599), .B(n2267), .Z(out[1449]) );
  XOR U3871 ( .A(in[681]), .B(n4292), .Z(n2771) );
  XOR U3872 ( .A(in[615]), .B(n4144), .Z(n4478) );
  XNOR U3873 ( .A(in[206]), .B(n3962), .Z(n4475) );
  NANDN U3874 ( .A(n4478), .B(n4475), .Z(n2268) );
  XNOR U3875 ( .A(n2771), .B(n2268), .Z(out[144]) );
  XOR U3876 ( .A(in[831]), .B(n3919), .Z(n2603) );
  NANDN U3877 ( .A(n2400), .B(n2269), .Z(n2270) );
  XOR U3878 ( .A(n2603), .B(n2270), .Z(out[1450]) );
  XOR U3879 ( .A(in[768]), .B(n3923), .Z(n2607) );
  NANDN U3880 ( .A(n2401), .B(n2271), .Z(n2272) );
  XOR U3881 ( .A(n2607), .B(n2272), .Z(out[1451]) );
  XOR U3882 ( .A(in[769]), .B(n3927), .Z(n2613) );
  NANDN U3883 ( .A(n2402), .B(n2273), .Z(n2274) );
  XOR U3884 ( .A(n2613), .B(n2274), .Z(out[1452]) );
  XNOR U3885 ( .A(n3932), .B(in[770]), .Z(n2617) );
  NANDN U3886 ( .A(n2403), .B(n2275), .Z(n2276) );
  XNOR U3887 ( .A(n2617), .B(n2276), .Z(out[1453]) );
  IV U3888 ( .A(n3173), .Z(n3936) );
  XOR U3889 ( .A(n3936), .B(in[771]), .Z(n2621) );
  NANDN U3890 ( .A(n2404), .B(n2277), .Z(n2278) );
  XOR U3891 ( .A(n2621), .B(n2278), .Z(out[1454]) );
  IV U3892 ( .A(n3175), .Z(n3943) );
  XOR U3893 ( .A(n3943), .B(in[772]), .Z(n2625) );
  NANDN U3894 ( .A(n2405), .B(n2279), .Z(n2280) );
  XOR U3895 ( .A(n2625), .B(n2280), .Z(out[1455]) );
  IV U3896 ( .A(n3177), .Z(n3947) );
  XOR U3897 ( .A(n3947), .B(in[773]), .Z(n2629) );
  NANDN U3898 ( .A(n2407), .B(n2281), .Z(n2282) );
  XOR U3899 ( .A(n2629), .B(n2282), .Z(out[1456]) );
  IV U3900 ( .A(n3179), .Z(n3951) );
  XOR U3901 ( .A(n3951), .B(in[774]), .Z(n2633) );
  NANDN U3902 ( .A(n2408), .B(n2283), .Z(n2284) );
  XOR U3903 ( .A(n2633), .B(n2284), .Z(out[1457]) );
  IV U3904 ( .A(n3181), .Z(n3955) );
  XOR U3905 ( .A(n3955), .B(in[775]), .Z(n2637) );
  NANDN U3906 ( .A(n2409), .B(n2285), .Z(n2286) );
  XOR U3907 ( .A(n2637), .B(n2286), .Z(out[1458]) );
  IV U3908 ( .A(n3183), .Z(n3959) );
  XOR U3909 ( .A(n3959), .B(in[776]), .Z(n2641) );
  NAND U3910 ( .A(n2287), .B(n2410), .Z(n2288) );
  XOR U3911 ( .A(n2641), .B(n2288), .Z(out[1459]) );
  XOR U3912 ( .A(in[682]), .B(n4294), .Z(n2772) );
  XOR U3913 ( .A(in[616]), .B(n4148), .Z(n4512) );
  XNOR U3914 ( .A(in[207]), .B(n3966), .Z(n4509) );
  NANDN U3915 ( .A(n4512), .B(n4509), .Z(n2289) );
  XNOR U3916 ( .A(n2772), .B(n2289), .Z(out[145]) );
  IV U3917 ( .A(n3185), .Z(n3963) );
  XOR U3918 ( .A(in[777]), .B(n3963), .Z(n2645) );
  NAND U3919 ( .A(n2290), .B(n2412), .Z(n2291) );
  XOR U3920 ( .A(n2645), .B(n2291), .Z(out[1460]) );
  IV U3921 ( .A(n3187), .Z(n3967) );
  XOR U3922 ( .A(n3967), .B(in[778]), .Z(n2649) );
  NAND U3923 ( .A(n2292), .B(n2414), .Z(n2293) );
  XOR U3924 ( .A(n2649), .B(n2293), .Z(out[1461]) );
  IV U3925 ( .A(n2294), .Z(n3971) );
  XOR U3926 ( .A(n3971), .B(in[779]), .Z(n2655) );
  NANDN U3927 ( .A(n2416), .B(n2295), .Z(n2296) );
  XOR U3928 ( .A(n2655), .B(n2296), .Z(out[1462]) );
  IV U3929 ( .A(n3194), .Z(n3975) );
  XOR U3930 ( .A(in[780]), .B(n3975), .Z(n2659) );
  NANDN U3931 ( .A(n2417), .B(n2297), .Z(n2298) );
  XOR U3932 ( .A(n2659), .B(n2298), .Z(out[1463]) );
  IV U3933 ( .A(n3196), .Z(n3979) );
  XOR U3934 ( .A(in[781]), .B(n3979), .Z(n2663) );
  NANDN U3935 ( .A(n2418), .B(n2299), .Z(n2300) );
  XOR U3936 ( .A(n2663), .B(n2300), .Z(out[1464]) );
  IV U3937 ( .A(n3199), .Z(n3986) );
  XOR U3938 ( .A(in[782]), .B(n3986), .Z(n2667) );
  NAND U3939 ( .A(n2301), .B(n2419), .Z(n2302) );
  XOR U3940 ( .A(n2667), .B(n2302), .Z(out[1465]) );
  IV U3941 ( .A(n3202), .Z(n3990) );
  XOR U3942 ( .A(in[783]), .B(n3990), .Z(n2671) );
  NAND U3943 ( .A(n2303), .B(n2422), .Z(n2304) );
  XOR U3944 ( .A(n2671), .B(n2304), .Z(out[1466]) );
  IV U3945 ( .A(n3205), .Z(n3994) );
  XOR U3946 ( .A(in[784]), .B(n3994), .Z(n2675) );
  NAND U3947 ( .A(n2305), .B(n2424), .Z(n2306) );
  XOR U3948 ( .A(n2675), .B(n2306), .Z(out[1467]) );
  IV U3949 ( .A(n3208), .Z(n3998) );
  XOR U3950 ( .A(in[785]), .B(n3998), .Z(n2679) );
  NAND U3951 ( .A(n2307), .B(n2426), .Z(n2308) );
  XOR U3952 ( .A(n2679), .B(n2308), .Z(out[1468]) );
  IV U3953 ( .A(n3211), .Z(n4002) );
  XOR U3954 ( .A(in[786]), .B(n4002), .Z(n2683) );
  NAND U3955 ( .A(n2309), .B(n2428), .Z(n2310) );
  XOR U3956 ( .A(n2683), .B(n2310), .Z(out[1469]) );
  XOR U3957 ( .A(in[683]), .B(n4296), .Z(n2776) );
  XOR U3958 ( .A(in[617]), .B(n4152), .Z(n4551) );
  XNOR U3959 ( .A(in[208]), .B(n3970), .Z(n4548) );
  NANDN U3960 ( .A(n4551), .B(n4548), .Z(n2311) );
  XNOR U3961 ( .A(n2776), .B(n2311), .Z(out[146]) );
  XOR U3962 ( .A(in[787]), .B(n4006), .Z(n2687) );
  NAND U3963 ( .A(n2312), .B(n2430), .Z(n2313) );
  XOR U3964 ( .A(n2687), .B(n2313), .Z(out[1470]) );
  XOR U3965 ( .A(in[788]), .B(n4010), .Z(n2691) );
  NAND U3966 ( .A(n2314), .B(n2432), .Z(n2315) );
  XOR U3967 ( .A(n2691), .B(n2315), .Z(out[1471]) );
  NANDN U3968 ( .A(n2316), .B(n2434), .Z(n2317) );
  XOR U3969 ( .A(n2435), .B(n2317), .Z(out[1472]) );
  NANDN U3970 ( .A(n2318), .B(n2437), .Z(n2319) );
  XOR U3971 ( .A(n2438), .B(n2319), .Z(out[1473]) );
  NANDN U3972 ( .A(n2320), .B(n2442), .Z(n2321) );
  XOR U3973 ( .A(n2443), .B(n2321), .Z(out[1474]) );
  NANDN U3974 ( .A(n2322), .B(n2446), .Z(n2323) );
  XOR U3975 ( .A(n2447), .B(n2323), .Z(out[1475]) );
  NANDN U3976 ( .A(n2324), .B(n2453), .Z(n2325) );
  XOR U3977 ( .A(n2454), .B(n2325), .Z(out[1476]) );
  NANDN U3978 ( .A(n2326), .B(n2456), .Z(n2327) );
  XOR U3979 ( .A(n2457), .B(n2327), .Z(out[1477]) );
  NANDN U3980 ( .A(n2328), .B(n2458), .Z(n2329) );
  XOR U3981 ( .A(n2459), .B(n2329), .Z(out[1478]) );
  NANDN U3982 ( .A(n2330), .B(n2462), .Z(n2331) );
  XOR U3983 ( .A(n2463), .B(n2331), .Z(out[1479]) );
  XNOR U3984 ( .A(in[684]), .B(n4298), .Z(n2907) );
  XOR U3985 ( .A(in[618]), .B(n4162), .Z(n4580) );
  XNOR U3986 ( .A(in[209]), .B(n3974), .Z(n4577) );
  NANDN U3987 ( .A(n4580), .B(n4577), .Z(n2332) );
  XOR U3988 ( .A(n2907), .B(n2332), .Z(out[147]) );
  NANDN U3989 ( .A(n2333), .B(n2468), .Z(n2334) );
  XOR U3990 ( .A(n2469), .B(n2334), .Z(out[1480]) );
  IV U3991 ( .A(n2335), .Z(n2471) );
  NANDN U3992 ( .A(n2336), .B(n2471), .Z(n2337) );
  XOR U3993 ( .A(n2472), .B(n2337), .Z(out[1481]) );
  IV U3994 ( .A(n2338), .Z(n2474) );
  NANDN U3995 ( .A(n2339), .B(n2474), .Z(n2340) );
  XOR U3996 ( .A(n2475), .B(n2340), .Z(out[1482]) );
  IV U3997 ( .A(n2341), .Z(n2477) );
  NANDN U3998 ( .A(n2342), .B(n2477), .Z(n2343) );
  XOR U3999 ( .A(n2478), .B(n2343), .Z(out[1483]) );
  IV U4000 ( .A(n2344), .Z(n2480) );
  NANDN U4001 ( .A(n2345), .B(n2480), .Z(n2346) );
  XOR U4002 ( .A(n2481), .B(n2346), .Z(out[1484]) );
  IV U4003 ( .A(n2347), .Z(n2483) );
  NANDN U4004 ( .A(n2348), .B(n2483), .Z(n2349) );
  XOR U4005 ( .A(n2484), .B(n2349), .Z(out[1485]) );
  IV U4006 ( .A(n2350), .Z(n2487) );
  NANDN U4007 ( .A(n2351), .B(n2487), .Z(n2352) );
  XNOR U4008 ( .A(n2486), .B(n2352), .Z(out[1486]) );
  IV U4009 ( .A(n2354), .Z(n2491) );
  OR U4010 ( .A(n2499), .B(n2356), .Z(n2357) );
  XOR U4011 ( .A(n2500), .B(n2357), .Z(out[1489]) );
  XNOR U4012 ( .A(in[685]), .B(n4300), .Z(n2910) );
  XOR U4013 ( .A(in[619]), .B(n4166), .Z(n4605) );
  XNOR U4014 ( .A(in[210]), .B(n3978), .Z(n4602) );
  NANDN U4015 ( .A(n4605), .B(n4602), .Z(n2358) );
  XOR U4016 ( .A(n2910), .B(n2358), .Z(out[148]) );
  OR U4017 ( .A(n2503), .B(n2359), .Z(n2360) );
  XOR U4018 ( .A(n2504), .B(n2360), .Z(out[1490]) );
  OR U4019 ( .A(n2507), .B(n2361), .Z(n2362) );
  XOR U4020 ( .A(n2508), .B(n2362), .Z(out[1491]) );
  OR U4021 ( .A(n2511), .B(n2363), .Z(n2364) );
  XOR U4022 ( .A(n2512), .B(n2364), .Z(out[1492]) );
  OR U4023 ( .A(n2515), .B(n2365), .Z(n2366) );
  XOR U4024 ( .A(n2516), .B(n2366), .Z(out[1493]) );
  NANDN U4025 ( .A(n2367), .B(n2519), .Z(n2368) );
  XOR U4026 ( .A(n2520), .B(n2368), .Z(out[1494]) );
  NANDN U4027 ( .A(n2369), .B(n2523), .Z(n2370) );
  XNOR U4028 ( .A(n2524), .B(n2370), .Z(out[1495]) );
  NANDN U4029 ( .A(n2371), .B(n2528), .Z(n2372) );
  XNOR U4030 ( .A(n2529), .B(n2372), .Z(out[1496]) );
  NANDN U4031 ( .A(n2373), .B(n2532), .Z(n2374) );
  XNOR U4032 ( .A(n2533), .B(n2374), .Z(out[1497]) );
  NANDN U4033 ( .A(n2375), .B(n2536), .Z(n2376) );
  XNOR U4034 ( .A(n2537), .B(n2376), .Z(out[1498]) );
  XOR U4035 ( .A(in[686]), .B(n4302), .Z(n2913) );
  XOR U4036 ( .A(in[211]), .B(n3349), .Z(n4630) );
  XNOR U4037 ( .A(in[620]), .B(n4170), .Z(n4632) );
  NANDN U4038 ( .A(n4630), .B(n4632), .Z(n2378) );
  XNOR U4039 ( .A(n2913), .B(n2378), .Z(out[149]) );
  XOR U4040 ( .A(in[1424]), .B(n3205), .Z(n4404) );
  XNOR U4041 ( .A(in[1047]), .B(n4497), .Z(n2891) );
  NANDN U4042 ( .A(n4404), .B(n2891), .Z(n2379) );
  XNOR U4043 ( .A(n4403), .B(n2379), .Z(out[14]) );
  NANDN U4044 ( .A(n2380), .B(n2544), .Z(n2381) );
  XNOR U4045 ( .A(n2545), .B(n2381), .Z(out[1500]) );
  NANDN U4046 ( .A(n2382), .B(n2548), .Z(n2383) );
  XNOR U4047 ( .A(n2549), .B(n2383), .Z(out[1501]) );
  NANDN U4048 ( .A(n2384), .B(n2552), .Z(n2385) );
  XNOR U4049 ( .A(n2553), .B(n2385), .Z(out[1502]) );
  NANDN U4050 ( .A(n2386), .B(n2556), .Z(n2387) );
  XNOR U4051 ( .A(n2557), .B(n2387), .Z(out[1503]) );
  NANDN U4052 ( .A(n2388), .B(n2561), .Z(n2389) );
  XNOR U4053 ( .A(n2562), .B(n2389), .Z(out[1504]) );
  XOR U4054 ( .A(in[687]), .B(n4304), .Z(n2916) );
  XOR U4055 ( .A(in[621]), .B(n4174), .Z(n4662) );
  XOR U4056 ( .A(in[212]), .B(n3989), .Z(n4659) );
  NANDN U4057 ( .A(n4662), .B(n4659), .Z(n2395) );
  XNOR U4058 ( .A(n2916), .B(n2395), .Z(out[150]) );
  XOR U4059 ( .A(in[688]), .B(n4311), .Z(n2919) );
  XOR U4060 ( .A(in[213]), .B(n3993), .Z(n4674) );
  XNOR U4061 ( .A(in[622]), .B(n3898), .Z(n4676) );
  NANDN U4062 ( .A(n4674), .B(n4676), .Z(n2406) );
  XNOR U4063 ( .A(n2919), .B(n2406), .Z(out[151]) );
  NANDN U4064 ( .A(n2410), .B(n2641), .Z(n2411) );
  XOR U4065 ( .A(n2642), .B(n2411), .Z(out[1523]) );
  NANDN U4066 ( .A(n2412), .B(n2645), .Z(n2413) );
  XOR U4067 ( .A(n2646), .B(n2413), .Z(out[1524]) );
  NANDN U4068 ( .A(n2414), .B(n2649), .Z(n2415) );
  XOR U4069 ( .A(n2650), .B(n2415), .Z(out[1525]) );
  NANDN U4070 ( .A(n2419), .B(n2667), .Z(n2420) );
  XOR U4071 ( .A(n2668), .B(n2420), .Z(out[1529]) );
  XOR U4072 ( .A(in[689]), .B(n4314), .Z(n2925) );
  XOR U4073 ( .A(in[214]), .B(n3997), .Z(n4690) );
  XNOR U4074 ( .A(in[623]), .B(n3902), .Z(n4692) );
  NANDN U4075 ( .A(n4690), .B(n4692), .Z(n2421) );
  XNOR U4076 ( .A(n2925), .B(n2421), .Z(out[152]) );
  NANDN U4077 ( .A(n2422), .B(n2671), .Z(n2423) );
  XOR U4078 ( .A(n2672), .B(n2423), .Z(out[1530]) );
  NANDN U4079 ( .A(n2424), .B(n2675), .Z(n2425) );
  XOR U4080 ( .A(n2676), .B(n2425), .Z(out[1531]) );
  NANDN U4081 ( .A(n2426), .B(n2679), .Z(n2427) );
  XOR U4082 ( .A(n2680), .B(n2427), .Z(out[1532]) );
  NANDN U4083 ( .A(n2428), .B(n2683), .Z(n2429) );
  XOR U4084 ( .A(n2684), .B(n2429), .Z(out[1533]) );
  NANDN U4085 ( .A(n2430), .B(n2687), .Z(n2431) );
  XOR U4086 ( .A(n2688), .B(n2431), .Z(out[1534]) );
  NANDN U4087 ( .A(n2432), .B(n2691), .Z(n2433) );
  XOR U4088 ( .A(n2692), .B(n2433), .Z(out[1535]) );
  ANDN U4089 ( .B(n2438), .A(n2437), .Z(n2441) );
  XNOR U4090 ( .A(n2439), .B(round_const[1]), .Z(n2440) );
  XNOR U4091 ( .A(n2441), .B(n2440), .Z(out[1537]) );
  ANDN U4092 ( .B(n2443), .A(n2442), .Z(n2444) );
  XOR U4093 ( .A(n2445), .B(n2444), .Z(out[1538]) );
  ANDN U4094 ( .B(n2447), .A(n2446), .Z(n2450) );
  XOR U4095 ( .A(n2448), .B(round_const_3), .Z(n2449) );
  XNOR U4096 ( .A(n2450), .B(n2449), .Z(out[1539]) );
  XOR U4097 ( .A(in[690]), .B(n4317), .Z(n2928) );
  XOR U4098 ( .A(in[624]), .B(n3906), .Z(n4727) );
  XOR U4099 ( .A(in[215]), .B(n4001), .Z(n4724) );
  NANDN U4100 ( .A(n4727), .B(n4724), .Z(n2451) );
  XNOR U4101 ( .A(n2928), .B(n2451), .Z(out[153]) );
  ANDN U4102 ( .B(n2459), .A(n2458), .Z(n2460) );
  XOR U4103 ( .A(n2461), .B(n2460), .Z(out[1542]) );
  ANDN U4104 ( .B(n2463), .A(n2462), .Z(n2466) );
  XNOR U4105 ( .A(n2464), .B(round_const_7), .Z(n2465) );
  XNOR U4106 ( .A(n2466), .B(n2465), .Z(out[1543]) );
  XOR U4107 ( .A(in[691]), .B(n4320), .Z(n2931) );
  XOR U4108 ( .A(in[625]), .B(n3910), .Z(n4775) );
  XOR U4109 ( .A(in[216]), .B(n4005), .Z(n4772) );
  NANDN U4110 ( .A(n4775), .B(n4772), .Z(n2485) );
  XNOR U4111 ( .A(n2931), .B(n2485), .Z(out[154]) );
  NOR U4112 ( .A(n2487), .B(n2486), .Z(n2488) );
  XOR U4113 ( .A(n2489), .B(n2488), .Z(out[1550]) );
  NOR U4114 ( .A(n2491), .B(n2490), .Z(n2494) );
  XNOR U4115 ( .A(n2492), .B(round_const_15), .Z(n2493) );
  XNOR U4116 ( .A(n2494), .B(n2493), .Z(out[1551]) );
  ANDN U4117 ( .B(n2496), .A(n2495), .Z(n2497) );
  XOR U4118 ( .A(n2498), .B(n2497), .Z(out[1552]) );
  AND U4119 ( .A(n2500), .B(n2499), .Z(n2501) );
  XOR U4120 ( .A(n2502), .B(n2501), .Z(out[1553]) );
  AND U4121 ( .A(n2504), .B(n2503), .Z(n2505) );
  XOR U4122 ( .A(n2506), .B(n2505), .Z(out[1554]) );
  AND U4123 ( .A(n2508), .B(n2507), .Z(n2509) );
  XOR U4124 ( .A(n2510), .B(n2509), .Z(out[1555]) );
  AND U4125 ( .A(n2512), .B(n2511), .Z(n2513) );
  XOR U4126 ( .A(n2514), .B(n2513), .Z(out[1556]) );
  AND U4127 ( .A(n2516), .B(n2515), .Z(n2517) );
  XOR U4128 ( .A(n2518), .B(n2517), .Z(out[1557]) );
  ANDN U4129 ( .B(n2520), .A(n2519), .Z(n2521) );
  XOR U4130 ( .A(n2522), .B(n2521), .Z(out[1558]) );
  NOR U4131 ( .A(n2524), .B(n2523), .Z(n2525) );
  XOR U4132 ( .A(n2526), .B(n2525), .Z(out[1559]) );
  XOR U4133 ( .A(in[692]), .B(n4323), .Z(n2934) );
  XOR U4134 ( .A(in[626]), .B(n3914), .Z(n4819) );
  XOR U4135 ( .A(in[217]), .B(n4009), .Z(n4816) );
  NANDN U4136 ( .A(n4819), .B(n4816), .Z(n2527) );
  XNOR U4137 ( .A(n2934), .B(n2527), .Z(out[155]) );
  NOR U4138 ( .A(n2529), .B(n2528), .Z(n2530) );
  XOR U4139 ( .A(n2531), .B(n2530), .Z(out[1560]) );
  NOR U4140 ( .A(n2533), .B(n2532), .Z(n2534) );
  XOR U4141 ( .A(n2535), .B(n2534), .Z(out[1561]) );
  NOR U4142 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U4143 ( .A(n2539), .B(n2538), .Z(out[1562]) );
  NOR U4144 ( .A(n2541), .B(n2540), .Z(n2542) );
  XOR U4145 ( .A(n2543), .B(n2542), .Z(out[1563]) );
  NOR U4146 ( .A(n2545), .B(n2544), .Z(n2546) );
  XOR U4147 ( .A(n2547), .B(n2546), .Z(out[1564]) );
  NOR U4148 ( .A(n2549), .B(n2548), .Z(n2550) );
  XOR U4149 ( .A(n2551), .B(n2550), .Z(out[1565]) );
  NOR U4150 ( .A(n2553), .B(n2552), .Z(n2554) );
  XOR U4151 ( .A(n2555), .B(n2554), .Z(out[1566]) );
  NOR U4152 ( .A(n2557), .B(n2556), .Z(n2560) );
  XNOR U4153 ( .A(n2558), .B(round_const_31), .Z(n2559) );
  XNOR U4154 ( .A(n2560), .B(n2559), .Z(out[1567]) );
  NOR U4155 ( .A(n2562), .B(n2561), .Z(n2563) );
  XOR U4156 ( .A(n2564), .B(n2563), .Z(out[1568]) );
  NOR U4157 ( .A(n2566), .B(n2565), .Z(n2567) );
  XOR U4158 ( .A(n2568), .B(n2567), .Z(out[1569]) );
  XOR U4159 ( .A(in[693]), .B(n4326), .Z(n2936) );
  XOR U4160 ( .A(in[218]), .B(n4013), .Z(n4861) );
  XNOR U4161 ( .A(in[627]), .B(n2569), .Z(n4863) );
  NANDN U4162 ( .A(n4861), .B(n4863), .Z(n2570) );
  XNOR U4163 ( .A(n2936), .B(n2570), .Z(out[156]) );
  NOR U4164 ( .A(n2572), .B(n2571), .Z(n2573) );
  XOR U4165 ( .A(n2574), .B(n2573), .Z(out[1570]) );
  NOR U4166 ( .A(n2576), .B(n2575), .Z(n2577) );
  XOR U4167 ( .A(n2578), .B(n2577), .Z(out[1571]) );
  NOR U4168 ( .A(n2580), .B(n2579), .Z(n2581) );
  XOR U4169 ( .A(n2582), .B(n2581), .Z(out[1572]) );
  NOR U4170 ( .A(n2584), .B(n2583), .Z(n2585) );
  XOR U4171 ( .A(n2586), .B(n2585), .Z(out[1573]) );
  NOR U4172 ( .A(n2588), .B(n2587), .Z(n2589) );
  XNOR U4173 ( .A(n2590), .B(n2589), .Z(out[1574]) );
  ANDN U4174 ( .B(n2592), .A(n2591), .Z(n2593) );
  XOR U4175 ( .A(n2594), .B(n2593), .Z(out[1575]) );
  ANDN U4176 ( .B(n2596), .A(n2595), .Z(n2597) );
  XOR U4177 ( .A(n2598), .B(n2597), .Z(out[1576]) );
  ANDN U4178 ( .B(n2600), .A(n2599), .Z(n2601) );
  XOR U4179 ( .A(n2602), .B(n2601), .Z(out[1577]) );
  NOR U4180 ( .A(n2604), .B(n2603), .Z(n2605) );
  XOR U4181 ( .A(n2606), .B(n2605), .Z(out[1578]) );
  ANDN U4182 ( .B(n2608), .A(n2607), .Z(n2609) );
  XOR U4183 ( .A(n2610), .B(n2609), .Z(out[1579]) );
  XOR U4184 ( .A(in[694]), .B(n4329), .Z(n2938) );
  XOR U4185 ( .A(in[219]), .B(n4017), .Z(n4905) );
  XNOR U4186 ( .A(in[628]), .B(n2611), .Z(n4907) );
  NANDN U4187 ( .A(n4905), .B(n4907), .Z(n2612) );
  XNOR U4188 ( .A(n2938), .B(n2612), .Z(out[157]) );
  ANDN U4189 ( .B(n2614), .A(n2613), .Z(n2615) );
  XOR U4190 ( .A(n2616), .B(n2615), .Z(out[1580]) );
  AND U4191 ( .A(n2618), .B(n2617), .Z(n2619) );
  XOR U4192 ( .A(n2620), .B(n2619), .Z(out[1581]) );
  ANDN U4193 ( .B(n2622), .A(n2621), .Z(n2623) );
  XOR U4194 ( .A(n2624), .B(n2623), .Z(out[1582]) );
  ANDN U4195 ( .B(n2626), .A(n2625), .Z(n2627) );
  XOR U4196 ( .A(n2628), .B(n2627), .Z(out[1583]) );
  ANDN U4197 ( .B(n2630), .A(n2629), .Z(n2631) );
  XOR U4198 ( .A(n2632), .B(n2631), .Z(out[1584]) );
  ANDN U4199 ( .B(n2634), .A(n2633), .Z(n2635) );
  XOR U4200 ( .A(n2636), .B(n2635), .Z(out[1585]) );
  ANDN U4201 ( .B(n2638), .A(n2637), .Z(n2639) );
  XOR U4202 ( .A(n2640), .B(n2639), .Z(out[1586]) );
  ANDN U4203 ( .B(n2642), .A(n2641), .Z(n2643) );
  XOR U4204 ( .A(n2644), .B(n2643), .Z(out[1587]) );
  ANDN U4205 ( .B(n2646), .A(n2645), .Z(n2647) );
  XOR U4206 ( .A(n2648), .B(n2647), .Z(out[1588]) );
  ANDN U4207 ( .B(n2650), .A(n2649), .Z(n2651) );
  XOR U4208 ( .A(n2652), .B(n2651), .Z(out[1589]) );
  XOR U4209 ( .A(in[695]), .B(n4332), .Z(n2940) );
  XNOR U4210 ( .A(in[220]), .B(n4021), .Z(n4949) );
  XNOR U4211 ( .A(in[629]), .B(n2653), .Z(n4951) );
  NANDN U4212 ( .A(n4949), .B(n4951), .Z(n2654) );
  XNOR U4213 ( .A(n2940), .B(n2654), .Z(out[158]) );
  ANDN U4214 ( .B(n2656), .A(n2655), .Z(n2657) );
  XNOR U4215 ( .A(n2658), .B(n2657), .Z(out[1590]) );
  ANDN U4216 ( .B(n2660), .A(n2659), .Z(n2661) );
  XNOR U4217 ( .A(n2662), .B(n2661), .Z(out[1591]) );
  ANDN U4218 ( .B(n2664), .A(n2663), .Z(n2665) );
  XNOR U4219 ( .A(n2666), .B(n2665), .Z(out[1592]) );
  ANDN U4220 ( .B(n2668), .A(n2667), .Z(n2669) );
  XOR U4221 ( .A(n2670), .B(n2669), .Z(out[1593]) );
  ANDN U4222 ( .B(n2672), .A(n2671), .Z(n2673) );
  XOR U4223 ( .A(n2674), .B(n2673), .Z(out[1594]) );
  ANDN U4224 ( .B(n2676), .A(n2675), .Z(n2677) );
  XOR U4225 ( .A(n2678), .B(n2677), .Z(out[1595]) );
  ANDN U4226 ( .B(n2680), .A(n2679), .Z(n2681) );
  XOR U4227 ( .A(n2682), .B(n2681), .Z(out[1596]) );
  ANDN U4228 ( .B(n2684), .A(n2683), .Z(n2685) );
  XOR U4229 ( .A(n2686), .B(n2685), .Z(out[1597]) );
  ANDN U4230 ( .B(n2688), .A(n2687), .Z(n2689) );
  XOR U4231 ( .A(n2690), .B(n2689), .Z(out[1598]) );
  ANDN U4232 ( .B(n2692), .A(n2691), .Z(n2695) );
  XNOR U4233 ( .A(n2693), .B(round_const_63), .Z(n2694) );
  XNOR U4234 ( .A(n2695), .B(n2694), .Z(out[1599]) );
  XOR U4235 ( .A(in[696]), .B(n4178), .Z(n2942) );
  XNOR U4236 ( .A(in[221]), .B(n4029), .Z(n4993) );
  XNOR U4237 ( .A(in[630]), .B(n3065), .Z(n4995) );
  NANDN U4238 ( .A(n4993), .B(n4995), .Z(n2696) );
  XNOR U4239 ( .A(n2942), .B(n2696), .Z(out[159]) );
  XOR U4240 ( .A(in[1425]), .B(n3208), .Z(n4438) );
  XNOR U4241 ( .A(in[1048]), .B(n4500), .Z(n2894) );
  NANDN U4242 ( .A(n4438), .B(n2894), .Z(n2697) );
  XNOR U4243 ( .A(n4437), .B(n2697), .Z(out[15]) );
  XOR U4244 ( .A(in[697]), .B(n4181), .Z(n2944) );
  XNOR U4245 ( .A(in[222]), .B(n4033), .Z(n5037) );
  XNOR U4246 ( .A(in[631]), .B(n3067), .Z(n5039) );
  NANDN U4247 ( .A(n5037), .B(n5039), .Z(n2698) );
  XNOR U4248 ( .A(n2944), .B(n2698), .Z(out[160]) );
  XOR U4249 ( .A(in[698]), .B(n4184), .Z(n2946) );
  XNOR U4250 ( .A(in[223]), .B(n4037), .Z(n5078) );
  XNOR U4251 ( .A(in[632]), .B(n3070), .Z(n5080) );
  NANDN U4252 ( .A(n5078), .B(n5080), .Z(n2699) );
  XNOR U4253 ( .A(n2946), .B(n2699), .Z(out[161]) );
  XOR U4254 ( .A(in[699]), .B(n4187), .Z(n2950) );
  XNOR U4255 ( .A(in[633]), .B(n2700), .Z(n5115) );
  XOR U4256 ( .A(in[224]), .B(n4041), .Z(n5112) );
  NAND U4257 ( .A(n5115), .B(n5112), .Z(n2701) );
  XNOR U4258 ( .A(n2950), .B(n2701), .Z(out[162]) );
  XOR U4259 ( .A(in[700]), .B(n4190), .Z(n2952) );
  XNOR U4260 ( .A(in[634]), .B(n2702), .Z(n5158) );
  XOR U4261 ( .A(in[225]), .B(n4045), .Z(n5155) );
  NAND U4262 ( .A(n5158), .B(n5155), .Z(n2703) );
  XOR U4263 ( .A(n2952), .B(n2703), .Z(out[163]) );
  XOR U4264 ( .A(in[701]), .B(n4193), .Z(n2954) );
  ANDN U4265 ( .B(n3115), .A(n2704), .Z(n2705) );
  XNOR U4266 ( .A(n2954), .B(n2705), .Z(out[164]) );
  XOR U4267 ( .A(in[702]), .B(n4198), .Z(n2956) );
  ANDN U4268 ( .B(n3137), .A(n2706), .Z(n2707) );
  XNOR U4269 ( .A(n2956), .B(n2707), .Z(out[165]) );
  XNOR U4270 ( .A(in[703]), .B(n4199), .Z(n2958) );
  ANDN U4271 ( .B(n3156), .A(n2708), .Z(n2709) );
  XNOR U4272 ( .A(n2958), .B(n2709), .Z(out[166]) );
  XOR U4273 ( .A(in[640]), .B(n4200), .Z(n2960) );
  ANDN U4274 ( .B(n3167), .A(n2710), .Z(n2711) );
  XNOR U4275 ( .A(n2960), .B(n2711), .Z(out[167]) );
  XOR U4276 ( .A(in[641]), .B(n4201), .Z(n2962) );
  NOR U4277 ( .A(n2712), .B(n3192), .Z(n2713) );
  XNOR U4278 ( .A(n2962), .B(n2713), .Z(out[168]) );
  XOR U4279 ( .A(in[642]), .B(n4202), .Z(n2964) );
  NOR U4280 ( .A(n2714), .B(n3223), .Z(n2715) );
  XNOR U4281 ( .A(n2964), .B(n2715), .Z(out[169]) );
  XOR U4282 ( .A(in[1426]), .B(n3211), .Z(n4476) );
  XNOR U4283 ( .A(in[1049]), .B(n4503), .Z(n2897) );
  NANDN U4284 ( .A(n4476), .B(n2897), .Z(n2716) );
  XNOR U4285 ( .A(n4475), .B(n2716), .Z(out[16]) );
  XOR U4286 ( .A(in[643]), .B(n4203), .Z(n2966) );
  NOR U4287 ( .A(n2717), .B(n3247), .Z(n2718) );
  XNOR U4288 ( .A(n2966), .B(n2718), .Z(out[170]) );
  XOR U4289 ( .A(in[644]), .B(n4204), .Z(n2968) );
  NOR U4290 ( .A(n2719), .B(n3259), .Z(n2720) );
  XNOR U4291 ( .A(n2968), .B(n2720), .Z(out[171]) );
  XOR U4292 ( .A(in[645]), .B(n4205), .Z(n2974) );
  NOR U4293 ( .A(n2721), .B(n3269), .Z(n2722) );
  XNOR U4294 ( .A(n2974), .B(n2722), .Z(out[172]) );
  XOR U4295 ( .A(in[646]), .B(n4208), .Z(n2976) );
  NOR U4296 ( .A(n3303), .B(n2811), .Z(n2723) );
  XNOR U4297 ( .A(n2976), .B(n2723), .Z(out[173]) );
  XOR U4298 ( .A(in[647]), .B(n4211), .Z(n2978) );
  NOR U4299 ( .A(n3333), .B(n2813), .Z(n2724) );
  XNOR U4300 ( .A(n2978), .B(n2724), .Z(out[174]) );
  XNOR U4301 ( .A(in[648]), .B(n4216), .Z(n2980) );
  NOR U4302 ( .A(n3362), .B(n2815), .Z(n2725) );
  XNOR U4303 ( .A(n2980), .B(n2725), .Z(out[175]) );
  XOR U4304 ( .A(in[649]), .B(n4219), .Z(n2982) );
  NOR U4305 ( .A(n3390), .B(n2820), .Z(n2726) );
  XNOR U4306 ( .A(n2982), .B(n2726), .Z(out[176]) );
  XOR U4307 ( .A(in[650]), .B(n3090), .Z(n2984) );
  NOR U4308 ( .A(n3425), .B(n2822), .Z(n2727) );
  XOR U4309 ( .A(n2984), .B(n2727), .Z(out[177]) );
  IV U4310 ( .A(n3092), .Z(n4225) );
  XOR U4311 ( .A(in[651]), .B(n4225), .Z(n2985) );
  NOR U4312 ( .A(n3460), .B(n2824), .Z(n2728) );
  XNOR U4313 ( .A(n2985), .B(n2728), .Z(out[178]) );
  IV U4314 ( .A(n3094), .Z(n4228) );
  XOR U4315 ( .A(in[652]), .B(n4228), .Z(n2987) );
  NOR U4316 ( .A(n3482), .B(n2826), .Z(n2729) );
  XNOR U4317 ( .A(n2987), .B(n2729), .Z(out[179]) );
  XOR U4318 ( .A(in[1427]), .B(n3214), .Z(n4510) );
  XNOR U4319 ( .A(in[1050]), .B(n4506), .Z(n2900) );
  NANDN U4320 ( .A(n4510), .B(n2900), .Z(n2730) );
  XNOR U4321 ( .A(n4509), .B(n2730), .Z(out[17]) );
  IV U4322 ( .A(n3098), .Z(n4231) );
  XOR U4323 ( .A(in[653]), .B(n4231), .Z(n2989) );
  NOR U4324 ( .A(n3504), .B(n2828), .Z(n2731) );
  XNOR U4325 ( .A(n2989), .B(n2731), .Z(out[180]) );
  XNOR U4326 ( .A(in[654]), .B(n4234), .Z(n2992) );
  NOR U4327 ( .A(n3519), .B(n2830), .Z(n2732) );
  XNOR U4328 ( .A(n2992), .B(n2732), .Z(out[181]) );
  XNOR U4329 ( .A(in[655]), .B(n4237), .Z(n2997) );
  NOR U4330 ( .A(n3547), .B(n2832), .Z(n2733) );
  XNOR U4331 ( .A(n2997), .B(n2733), .Z(out[182]) );
  XNOR U4332 ( .A(in[656]), .B(n4240), .Z(n3000) );
  NOR U4333 ( .A(n3577), .B(n2834), .Z(n2734) );
  XNOR U4334 ( .A(n3000), .B(n2734), .Z(out[183]) );
  XNOR U4335 ( .A(in[657]), .B(n4241), .Z(n3003) );
  NOR U4336 ( .A(n3601), .B(n2836), .Z(n2735) );
  XNOR U4337 ( .A(n3003), .B(n2735), .Z(out[184]) );
  IV U4338 ( .A(n3104), .Z(n4244) );
  XOR U4339 ( .A(in[658]), .B(n4244), .Z(n3005) );
  NOR U4340 ( .A(n3631), .B(n2838), .Z(n2736) );
  XNOR U4341 ( .A(n3005), .B(n2736), .Z(out[185]) );
  IV U4342 ( .A(n3106), .Z(n4245) );
  XOR U4343 ( .A(in[659]), .B(n4245), .Z(n3007) );
  NOR U4344 ( .A(n3675), .B(n2843), .Z(n2737) );
  XNOR U4345 ( .A(n3007), .B(n2737), .Z(out[186]) );
  XOR U4346 ( .A(in[660]), .B(n4248), .Z(n3009) );
  NOR U4347 ( .A(n3719), .B(n2845), .Z(n2738) );
  XOR U4348 ( .A(n3009), .B(n2738), .Z(out[187]) );
  XOR U4349 ( .A(in[661]), .B(n4251), .Z(n3012) );
  NOR U4350 ( .A(n3765), .B(n2847), .Z(n2739) );
  XOR U4351 ( .A(n3012), .B(n2739), .Z(out[188]) );
  XOR U4352 ( .A(in[662]), .B(n4252), .Z(n3015) );
  XOR U4353 ( .A(in[1428]), .B(n3217), .Z(n4549) );
  XNOR U4354 ( .A(in[1051]), .B(n2740), .Z(n2903) );
  NANDN U4355 ( .A(n4549), .B(n2903), .Z(n2741) );
  XNOR U4356 ( .A(n4548), .B(n2741), .Z(out[18]) );
  XOR U4357 ( .A(in[663]), .B(n4253), .Z(n3016) );
  XOR U4358 ( .A(in[664]), .B(n4254), .Z(n3019) );
  NANDN U4359 ( .A(n2855), .B(n3940), .Z(n2742) );
  XOR U4360 ( .A(n2856), .B(n2742), .Z(out[192]) );
  XNOR U4361 ( .A(in[1034]), .B(n4454), .Z(n2759) );
  ANDN U4362 ( .B(n3983), .A(n2858), .Z(n2743) );
  XNOR U4363 ( .A(n2759), .B(n2743), .Z(out[193]) );
  XNOR U4364 ( .A(in[1035]), .B(n4457), .Z(n2972) );
  ANDN U4365 ( .B(n4027), .A(n2744), .Z(n2745) );
  XNOR U4366 ( .A(n2972), .B(n2745), .Z(out[194]) );
  XOR U4367 ( .A(n4460), .B(in[1036]), .Z(n3168) );
  ANDN U4368 ( .B(n4071), .A(n2746), .Z(n2747) );
  XNOR U4369 ( .A(n3168), .B(n2747), .Z(out[195]) );
  XOR U4370 ( .A(n4463), .B(in[1037]), .Z(n3426) );
  ANDN U4371 ( .B(n4115), .A(n2748), .Z(n2749) );
  XNOR U4372 ( .A(n3426), .B(n2749), .Z(out[196]) );
  XOR U4373 ( .A(n4466), .B(in[1038]), .Z(n3720) );
  ANDN U4374 ( .B(n4159), .A(n2750), .Z(n2751) );
  XNOR U4375 ( .A(n3720), .B(n2751), .Z(out[197]) );
  XOR U4376 ( .A(n4469), .B(in[1039]), .Z(n4160) );
  ANDN U4377 ( .B(n4197), .A(n2752), .Z(n2753) );
  XNOR U4378 ( .A(n4160), .B(n2753), .Z(out[198]) );
  XOR U4379 ( .A(n4472), .B(in[1040]), .Z(n4441) );
  ANDN U4380 ( .B(n4215), .A(n2754), .Z(n2755) );
  XNOR U4381 ( .A(n4441), .B(n2755), .Z(out[199]) );
  XOR U4382 ( .A(in[1429]), .B(n2756), .Z(n4578) );
  XNOR U4383 ( .A(in[1052]), .B(n2757), .Z(n2906) );
  NANDN U4384 ( .A(n4578), .B(n2906), .Z(n2758) );
  XNOR U4385 ( .A(n4577), .B(n2758), .Z(out[19]) );
  XOR U4386 ( .A(n3173), .B(in[1411]), .Z(n3981) );
  IV U4387 ( .A(n2759), .Z(n2857) );
  NANDN U4388 ( .A(n3981), .B(n2857), .Z(n2760) );
  XNOR U4389 ( .A(n3982), .B(n2760), .Z(out[1]) );
  XOR U4390 ( .A(n4479), .B(in[1041]), .Z(n4728) );
  ANDN U4391 ( .B(n4243), .A(n2761), .Z(n2762) );
  XNOR U4392 ( .A(n4728), .B(n2762), .Z(out[200]) );
  XOR U4393 ( .A(n4482), .B(in[1042]), .Z(n5159) );
  ANDN U4394 ( .B(n4259), .A(n2763), .Z(n2764) );
  XNOR U4395 ( .A(n5159), .B(n2764), .Z(out[201]) );
  NAND U4396 ( .A(n4285), .B(n2880), .Z(n2765) );
  XNOR U4397 ( .A(n2879), .B(n2765), .Z(out[202]) );
  NANDN U4398 ( .A(n2882), .B(n4310), .Z(n2766) );
  XNOR U4399 ( .A(n2883), .B(n2766), .Z(out[203]) );
  NANDN U4400 ( .A(n2884), .B(n4342), .Z(n2767) );
  XNOR U4401 ( .A(n2885), .B(n2767), .Z(out[204]) );
  NANDN U4402 ( .A(n2886), .B(n4373), .Z(n2768) );
  XNOR U4403 ( .A(n2887), .B(n2768), .Z(out[205]) );
  IV U4404 ( .A(n2769), .Z(n2892) );
  IV U4405 ( .A(n2770), .Z(n2895) );
  IV U4406 ( .A(n2771), .Z(n2898) );
  IV U4407 ( .A(n2772), .Z(n2901) );
  XOR U4408 ( .A(in[1430]), .B(n2773), .Z(n4603) );
  XNOR U4409 ( .A(in[1053]), .B(n2774), .Z(n2909) );
  NANDN U4410 ( .A(n4603), .B(n2909), .Z(n2775) );
  XNOR U4411 ( .A(n4602), .B(n2775), .Z(out[20]) );
  IV U4412 ( .A(n2776), .Z(n2904) );
  XOR U4413 ( .A(in[1054]), .B(n4522), .Z(n2781) );
  IV U4414 ( .A(n2781), .Z(n2912) );
  NOR U4415 ( .A(n4632), .B(n2913), .Z(n2777) );
  XOR U4416 ( .A(n2912), .B(n2777), .Z(out[213]) );
  XOR U4417 ( .A(in[1055]), .B(n4526), .Z(n2795) );
  IV U4418 ( .A(n2795), .Z(n2915) );
  XOR U4419 ( .A(in[1056]), .B(n4530), .Z(n2818) );
  IV U4420 ( .A(n2818), .Z(n2918) );
  NOR U4421 ( .A(n4676), .B(n2919), .Z(n2778) );
  XOR U4422 ( .A(n2918), .B(n2778), .Z(out[215]) );
  XOR U4423 ( .A(in[1057]), .B(n4534), .Z(n2841) );
  IV U4424 ( .A(n2841), .Z(n2924) );
  NOR U4425 ( .A(n4692), .B(n2925), .Z(n2779) );
  XOR U4426 ( .A(n2924), .B(n2779), .Z(out[216]) );
  XOR U4427 ( .A(in[1058]), .B(n4538), .Z(n2865) );
  IV U4428 ( .A(n2865), .Z(n2927) );
  XOR U4429 ( .A(in[1059]), .B(n4542), .Z(n2889) );
  IV U4430 ( .A(n2889), .Z(n2930) );
  XNOR U4431 ( .A(in[1060]), .B(n4546), .Z(n2922) );
  IV U4432 ( .A(n2922), .Z(n2933) );
  XOR U4433 ( .A(in[1431]), .B(n2780), .Z(n4631) );
  OR U4434 ( .A(n4631), .B(n2781), .Z(n2782) );
  XOR U4435 ( .A(n4630), .B(n2782), .Z(out[21]) );
  XNOR U4436 ( .A(in[1061]), .B(n4552), .Z(n2948) );
  NOR U4437 ( .A(n4863), .B(n2936), .Z(n2783) );
  XNOR U4438 ( .A(n2948), .B(n2783), .Z(out[220]) );
  XNOR U4439 ( .A(in[1062]), .B(n4554), .Z(n2970) );
  NOR U4440 ( .A(n4907), .B(n2938), .Z(n2784) );
  XNOR U4441 ( .A(n2970), .B(n2784), .Z(out[221]) );
  XNOR U4442 ( .A(in[1063]), .B(n4335), .Z(n2994) );
  NOR U4443 ( .A(n4951), .B(n2940), .Z(n2785) );
  XNOR U4444 ( .A(n2994), .B(n2785), .Z(out[222]) );
  XNOR U4445 ( .A(in[1064]), .B(n4337), .Z(n3022) );
  NOR U4446 ( .A(n4995), .B(n2942), .Z(n2786) );
  XNOR U4447 ( .A(n3022), .B(n2786), .Z(out[223]) );
  XNOR U4448 ( .A(in[1065]), .B(n4343), .Z(n3042) );
  NOR U4449 ( .A(n5039), .B(n2944), .Z(n2787) );
  XNOR U4450 ( .A(n3042), .B(n2787), .Z(out[224]) );
  XNOR U4451 ( .A(in[1066]), .B(n4345), .Z(n3054) );
  NOR U4452 ( .A(n5080), .B(n2946), .Z(n2788) );
  XNOR U4453 ( .A(n3054), .B(n2788), .Z(out[225]) );
  XNOR U4454 ( .A(in[1067]), .B(n4347), .Z(n3075) );
  NOR U4455 ( .A(n5115), .B(n2950), .Z(n2789) );
  XNOR U4456 ( .A(n3075), .B(n2789), .Z(out[226]) );
  XNOR U4457 ( .A(in[1068]), .B(n4350), .Z(n3096) );
  XOR U4458 ( .A(in[1069]), .B(n4353), .Z(n3113) );
  NANDN U4459 ( .A(n2790), .B(n2954), .Z(n2791) );
  XNOR U4460 ( .A(n3113), .B(n2791), .Z(out[228]) );
  XOR U4461 ( .A(in[1070]), .B(n4356), .Z(n3135) );
  NANDN U4462 ( .A(n2792), .B(n2956), .Z(n2793) );
  XNOR U4463 ( .A(n3135), .B(n2793), .Z(out[229]) );
  XOR U4464 ( .A(in[1432]), .B(n2794), .Z(n4660) );
  OR U4465 ( .A(n4660), .B(n2795), .Z(n2796) );
  XNOR U4466 ( .A(n4659), .B(n2796), .Z(out[22]) );
  XNOR U4467 ( .A(in[1071]), .B(n4358), .Z(n3153) );
  NANDN U4468 ( .A(n2797), .B(n2958), .Z(n2798) );
  XOR U4469 ( .A(n3153), .B(n2798), .Z(out[230]) );
  XOR U4470 ( .A(in[1072]), .B(n4361), .Z(n3165) );
  NANDN U4471 ( .A(n2799), .B(n2960), .Z(n2800) );
  XNOR U4472 ( .A(n3165), .B(n2800), .Z(out[231]) );
  XOR U4473 ( .A(in[1073]), .B(n4364), .Z(n3190) );
  NANDN U4474 ( .A(n2801), .B(n2962), .Z(n2802) );
  XNOR U4475 ( .A(n3190), .B(n2802), .Z(out[232]) );
  XOR U4476 ( .A(in[1074]), .B(n4367), .Z(n3220) );
  NANDN U4477 ( .A(n2803), .B(n2964), .Z(n2804) );
  XNOR U4478 ( .A(n3220), .B(n2804), .Z(out[233]) );
  XOR U4479 ( .A(in[1075]), .B(n4374), .Z(n3244) );
  NANDN U4480 ( .A(n2805), .B(n2966), .Z(n2806) );
  XNOR U4481 ( .A(n3244), .B(n2806), .Z(out[234]) );
  XOR U4482 ( .A(in[1076]), .B(n4377), .Z(n3256) );
  NANDN U4483 ( .A(n2807), .B(n2968), .Z(n2808) );
  XNOR U4484 ( .A(n3256), .B(n2808), .Z(out[235]) );
  XOR U4485 ( .A(in[1077]), .B(n4380), .Z(n3266) );
  NANDN U4486 ( .A(n2809), .B(n2974), .Z(n2810) );
  XNOR U4487 ( .A(n3266), .B(n2810), .Z(out[236]) );
  XOR U4488 ( .A(in[1078]), .B(n4383), .Z(n3300) );
  NAND U4489 ( .A(n2811), .B(n2976), .Z(n2812) );
  XNOR U4490 ( .A(n3300), .B(n2812), .Z(out[237]) );
  XOR U4491 ( .A(in[1079]), .B(n4386), .Z(n3330) );
  NAND U4492 ( .A(n2813), .B(n2978), .Z(n2814) );
  XNOR U4493 ( .A(n3330), .B(n2814), .Z(out[238]) );
  XNOR U4494 ( .A(in[1080]), .B(n4388), .Z(n3359) );
  NAND U4495 ( .A(n2815), .B(n2980), .Z(n2816) );
  XOR U4496 ( .A(n3359), .B(n2816), .Z(out[239]) );
  XOR U4497 ( .A(in[1433]), .B(n2817), .Z(n4675) );
  OR U4498 ( .A(n4675), .B(n2818), .Z(n2819) );
  XOR U4499 ( .A(n4674), .B(n2819), .Z(out[23]) );
  XOR U4500 ( .A(in[1081]), .B(n4391), .Z(n3387) );
  NAND U4501 ( .A(n2820), .B(n2982), .Z(n2821) );
  XNOR U4502 ( .A(n3387), .B(n2821), .Z(out[240]) );
  XOR U4503 ( .A(in[1082]), .B(n4394), .Z(n3422) );
  NANDN U4504 ( .A(n2984), .B(n2822), .Z(n2823) );
  XOR U4505 ( .A(n3422), .B(n2823), .Z(out[241]) );
  XOR U4506 ( .A(in[1083]), .B(n4397), .Z(n3457) );
  NAND U4507 ( .A(n2824), .B(n2985), .Z(n2825) );
  XOR U4508 ( .A(n3457), .B(n2825), .Z(out[242]) );
  XNOR U4509 ( .A(in[1084]), .B(n4400), .Z(n3479) );
  NAND U4510 ( .A(n2826), .B(n2987), .Z(n2827) );
  XOR U4511 ( .A(n3479), .B(n2827), .Z(out[243]) );
  XNOR U4512 ( .A(in[1085]), .B(n4407), .Z(n3501) );
  NAND U4513 ( .A(n2828), .B(n2989), .Z(n2829) );
  XOR U4514 ( .A(n3501), .B(n2829), .Z(out[244]) );
  XOR U4515 ( .A(in[1086]), .B(n4410), .Z(n2991) );
  NAND U4516 ( .A(n2830), .B(n2992), .Z(n2831) );
  XNOR U4517 ( .A(n2991), .B(n2831), .Z(out[245]) );
  XOR U4518 ( .A(in[1087]), .B(n4413), .Z(n2996) );
  NAND U4519 ( .A(n2832), .B(n2997), .Z(n2833) );
  XNOR U4520 ( .A(n2996), .B(n2833), .Z(out[246]) );
  XOR U4521 ( .A(in[1024]), .B(n4416), .Z(n2999) );
  NAND U4522 ( .A(n2834), .B(n3000), .Z(n2835) );
  XNOR U4523 ( .A(n2999), .B(n2835), .Z(out[247]) );
  XOR U4524 ( .A(in[1025]), .B(n4419), .Z(n3002) );
  NAND U4525 ( .A(n2836), .B(n3003), .Z(n2837) );
  XNOR U4526 ( .A(n3002), .B(n2837), .Z(out[248]) );
  XNOR U4527 ( .A(in[1026]), .B(n4422), .Z(n3628) );
  NAND U4528 ( .A(n2838), .B(n3005), .Z(n2839) );
  XOR U4529 ( .A(n3628), .B(n2839), .Z(out[249]) );
  XOR U4530 ( .A(in[1434]), .B(n2840), .Z(n4691) );
  OR U4531 ( .A(n4691), .B(n2841), .Z(n2842) );
  XOR U4532 ( .A(n4690), .B(n2842), .Z(out[24]) );
  XNOR U4533 ( .A(in[1027]), .B(n4425), .Z(n3672) );
  NAND U4534 ( .A(n2843), .B(n3007), .Z(n2844) );
  XOR U4535 ( .A(n3672), .B(n2844), .Z(out[250]) );
  XOR U4536 ( .A(in[1028]), .B(n4428), .Z(n3010) );
  IV U4537 ( .A(n3010), .Z(n3716) );
  NANDN U4538 ( .A(n3009), .B(n2845), .Z(n2846) );
  XOR U4539 ( .A(n3716), .B(n2846), .Z(out[251]) );
  XOR U4540 ( .A(in[1029]), .B(n4431), .Z(n3013) );
  IV U4541 ( .A(n3013), .Z(n3762) );
  NANDN U4542 ( .A(n3012), .B(n2847), .Z(n2848) );
  XOR U4543 ( .A(n3762), .B(n2848), .Z(out[252]) );
  XOR U4544 ( .A(in[1030]), .B(n4434), .Z(n3806) );
  NANDN U4545 ( .A(n3015), .B(n2849), .Z(n2850) );
  XOR U4546 ( .A(n3806), .B(n2850), .Z(out[253]) );
  XOR U4547 ( .A(in[1031]), .B(n4445), .Z(n3017) );
  IV U4548 ( .A(n3017), .Z(n3850) );
  NANDN U4549 ( .A(n3016), .B(n2851), .Z(n2852) );
  XOR U4550 ( .A(n3850), .B(n2852), .Z(out[254]) );
  XOR U4551 ( .A(in[1032]), .B(n4448), .Z(n3020) );
  IV U4552 ( .A(n3020), .Z(n3894) );
  NANDN U4553 ( .A(n3019), .B(n2853), .Z(n2854) );
  XOR U4554 ( .A(n3894), .B(n2854), .Z(out[255]) );
  ANDN U4555 ( .B(n2858), .A(n2857), .Z(n2859) );
  XOR U4556 ( .A(n3981), .B(n2859), .Z(out[257]) );
  XNOR U4557 ( .A(n3943), .B(in[1412]), .Z(n4025) );
  NANDN U4558 ( .A(n2860), .B(n2972), .Z(n2861) );
  XNOR U4559 ( .A(n4025), .B(n2861), .Z(out[258]) );
  XNOR U4560 ( .A(n3947), .B(in[1413]), .Z(n4069) );
  NANDN U4561 ( .A(n2862), .B(n3168), .Z(n2863) );
  XNOR U4562 ( .A(n4069), .B(n2863), .Z(out[259]) );
  XOR U4563 ( .A(in[1435]), .B(n2864), .Z(n4725) );
  OR U4564 ( .A(n4725), .B(n2865), .Z(n2866) );
  XNOR U4565 ( .A(n4724), .B(n2866), .Z(out[25]) );
  XNOR U4566 ( .A(n3951), .B(in[1414]), .Z(n4113) );
  NANDN U4567 ( .A(n2867), .B(n3426), .Z(n2868) );
  XNOR U4568 ( .A(n4113), .B(n2868), .Z(out[260]) );
  XNOR U4569 ( .A(n3955), .B(in[1415]), .Z(n4157) );
  NANDN U4570 ( .A(n2869), .B(n3720), .Z(n2870) );
  XNOR U4571 ( .A(n4157), .B(n2870), .Z(out[261]) );
  XNOR U4572 ( .A(n3959), .B(in[1416]), .Z(n4195) );
  NANDN U4573 ( .A(n2871), .B(n4160), .Z(n2872) );
  XNOR U4574 ( .A(n4195), .B(n2872), .Z(out[262]) );
  XNOR U4575 ( .A(in[1417]), .B(n3963), .Z(n4442) );
  NANDN U4576 ( .A(n2873), .B(n4441), .Z(n2874) );
  XNOR U4577 ( .A(n4442), .B(n2874), .Z(out[263]) );
  XNOR U4578 ( .A(n3967), .B(in[1418]), .Z(n4729) );
  NANDN U4579 ( .A(n2875), .B(n4728), .Z(n2876) );
  XNOR U4580 ( .A(n4729), .B(n2876), .Z(out[264]) );
  XNOR U4581 ( .A(n3971), .B(in[1419]), .Z(n5160) );
  NANDN U4582 ( .A(n2877), .B(n5159), .Z(n2878) );
  XNOR U4583 ( .A(n5160), .B(n2878), .Z(out[265]) );
  NOR U4584 ( .A(n2880), .B(n2879), .Z(n2881) );
  XOR U4585 ( .A(n4283), .B(n2881), .Z(out[266]) );
  XOR U4586 ( .A(in[1436]), .B(n2888), .Z(n4773) );
  OR U4587 ( .A(n4773), .B(n2889), .Z(n2890) );
  XNOR U4588 ( .A(n4772), .B(n2890), .Z(out[26]) );
  NOR U4589 ( .A(n2892), .B(n2891), .Z(n2893) );
  XOR U4590 ( .A(n4404), .B(n2893), .Z(out[270]) );
  NOR U4591 ( .A(n2895), .B(n2894), .Z(n2896) );
  XOR U4592 ( .A(n4438), .B(n2896), .Z(out[271]) );
  NOR U4593 ( .A(n2898), .B(n2897), .Z(n2899) );
  XOR U4594 ( .A(n4476), .B(n2899), .Z(out[272]) );
  NOR U4595 ( .A(n2901), .B(n2900), .Z(n2902) );
  XOR U4596 ( .A(n4510), .B(n2902), .Z(out[273]) );
  NOR U4597 ( .A(n2904), .B(n2903), .Z(n2905) );
  XOR U4598 ( .A(n4549), .B(n2905), .Z(out[274]) );
  NOR U4599 ( .A(n2907), .B(n2906), .Z(n2908) );
  XOR U4600 ( .A(n4578), .B(n2908), .Z(out[275]) );
  NOR U4601 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U4602 ( .A(n4603), .B(n2911), .Z(out[276]) );
  ANDN U4603 ( .B(n2913), .A(n2912), .Z(n2914) );
  XOR U4604 ( .A(n4631), .B(n2914), .Z(out[277]) );
  ANDN U4605 ( .B(n2916), .A(n2915), .Z(n2917) );
  XOR U4606 ( .A(n4660), .B(n2917), .Z(out[278]) );
  ANDN U4607 ( .B(n2919), .A(n2918), .Z(n2920) );
  XOR U4608 ( .A(n4675), .B(n2920), .Z(out[279]) );
  XOR U4609 ( .A(in[1437]), .B(n2921), .Z(n4817) );
  OR U4610 ( .A(n4817), .B(n2922), .Z(n2923) );
  XNOR U4611 ( .A(n4816), .B(n2923), .Z(out[27]) );
  ANDN U4612 ( .B(n2925), .A(n2924), .Z(n2926) );
  XOR U4613 ( .A(n4691), .B(n2926), .Z(out[280]) );
  ANDN U4614 ( .B(n2928), .A(n2927), .Z(n2929) );
  XOR U4615 ( .A(n4725), .B(n2929), .Z(out[281]) );
  ANDN U4616 ( .B(n2931), .A(n2930), .Z(n2932) );
  XOR U4617 ( .A(n4773), .B(n2932), .Z(out[282]) );
  ANDN U4618 ( .B(n2934), .A(n2933), .Z(n2935) );
  XOR U4619 ( .A(n4817), .B(n2935), .Z(out[283]) );
  XOR U4620 ( .A(in[1438]), .B(n4054), .Z(n4860) );
  NAND U4621 ( .A(n2936), .B(n2948), .Z(n2937) );
  XNOR U4622 ( .A(n4860), .B(n2937), .Z(out[284]) );
  XOR U4623 ( .A(in[1439]), .B(n4058), .Z(n4904) );
  NAND U4624 ( .A(n2938), .B(n2970), .Z(n2939) );
  XNOR U4625 ( .A(n4904), .B(n2939), .Z(out[285]) );
  XOR U4626 ( .A(in[1440]), .B(n4062), .Z(n4948) );
  NAND U4627 ( .A(n2940), .B(n2994), .Z(n2941) );
  XNOR U4628 ( .A(n4948), .B(n2941), .Z(out[286]) );
  XOR U4629 ( .A(in[1441]), .B(n4066), .Z(n4992) );
  NAND U4630 ( .A(n2942), .B(n3022), .Z(n2943) );
  XNOR U4631 ( .A(n4992), .B(n2943), .Z(out[287]) );
  XOR U4632 ( .A(in[1442]), .B(n4074), .Z(n5036) );
  NAND U4633 ( .A(n2944), .B(n3042), .Z(n2945) );
  XNOR U4634 ( .A(n5036), .B(n2945), .Z(out[288]) );
  XOR U4635 ( .A(in[1443]), .B(n4078), .Z(n5077) );
  NAND U4636 ( .A(n2946), .B(n3054), .Z(n2947) );
  XNOR U4637 ( .A(n5077), .B(n2947), .Z(out[289]) );
  OR U4638 ( .A(n4860), .B(n2948), .Z(n2949) );
  XOR U4639 ( .A(n4861), .B(n2949), .Z(out[28]) );
  XOR U4640 ( .A(in[1444]), .B(n4082), .Z(n5113) );
  NAND U4641 ( .A(n2950), .B(n3075), .Z(n2951) );
  XNOR U4642 ( .A(n5113), .B(n2951), .Z(out[290]) );
  XNOR U4643 ( .A(in[1445]), .B(n4086), .Z(n5156) );
  NANDN U4644 ( .A(n2952), .B(n3096), .Z(n2953) );
  XNOR U4645 ( .A(n5156), .B(n2953), .Z(out[291]) );
  OR U4646 ( .A(n3113), .B(n2954), .Z(n2955) );
  XNOR U4647 ( .A(n3112), .B(n2955), .Z(out[292]) );
  OR U4648 ( .A(n3135), .B(n2956), .Z(n2957) );
  XNOR U4649 ( .A(n3134), .B(n2957), .Z(out[293]) );
  NANDN U4650 ( .A(n2958), .B(n3153), .Z(n2959) );
  XNOR U4651 ( .A(n3154), .B(n2959), .Z(out[294]) );
  OR U4652 ( .A(n3165), .B(n2960), .Z(n2961) );
  XNOR U4653 ( .A(n3164), .B(n2961), .Z(out[295]) );
  OR U4654 ( .A(n3190), .B(n2962), .Z(n2963) );
  XNOR U4655 ( .A(n3189), .B(n2963), .Z(out[296]) );
  OR U4656 ( .A(n3220), .B(n2964), .Z(n2965) );
  XOR U4657 ( .A(n3221), .B(n2965), .Z(out[297]) );
  OR U4658 ( .A(n3244), .B(n2966), .Z(n2967) );
  XOR U4659 ( .A(n3245), .B(n2967), .Z(out[298]) );
  OR U4660 ( .A(n3256), .B(n2968), .Z(n2969) );
  XOR U4661 ( .A(n3257), .B(n2969), .Z(out[299]) );
  OR U4662 ( .A(n4904), .B(n2970), .Z(n2971) );
  XOR U4663 ( .A(n4905), .B(n2971), .Z(out[29]) );
  OR U4664 ( .A(n4025), .B(n2972), .Z(n2973) );
  XNOR U4665 ( .A(n4024), .B(n2973), .Z(out[2]) );
  OR U4666 ( .A(n3266), .B(n2974), .Z(n2975) );
  XOR U4667 ( .A(n3267), .B(n2975), .Z(out[300]) );
  OR U4668 ( .A(n3300), .B(n2976), .Z(n2977) );
  XOR U4669 ( .A(n3301), .B(n2977), .Z(out[301]) );
  OR U4670 ( .A(n3330), .B(n2978), .Z(n2979) );
  XOR U4671 ( .A(n3331), .B(n2979), .Z(out[302]) );
  NANDN U4672 ( .A(n2980), .B(n3359), .Z(n2981) );
  XOR U4673 ( .A(n3360), .B(n2981), .Z(out[303]) );
  OR U4674 ( .A(n3387), .B(n2982), .Z(n2983) );
  XOR U4675 ( .A(n3388), .B(n2983), .Z(out[304]) );
  NANDN U4676 ( .A(n2985), .B(n3457), .Z(n2986) );
  XOR U4677 ( .A(n3458), .B(n2986), .Z(out[306]) );
  NANDN U4678 ( .A(n2987), .B(n3479), .Z(n2988) );
  XOR U4679 ( .A(n3480), .B(n2988), .Z(out[307]) );
  NANDN U4680 ( .A(n2989), .B(n3501), .Z(n2990) );
  XOR U4681 ( .A(n3502), .B(n2990), .Z(out[308]) );
  IV U4682 ( .A(n2991), .Z(n3516) );
  NANDN U4683 ( .A(n2992), .B(n3516), .Z(n2993) );
  XOR U4684 ( .A(n3517), .B(n2993), .Z(out[309]) );
  OR U4685 ( .A(n4948), .B(n2994), .Z(n2995) );
  XOR U4686 ( .A(n4949), .B(n2995), .Z(out[30]) );
  IV U4687 ( .A(n2996), .Z(n3544) );
  NANDN U4688 ( .A(n2997), .B(n3544), .Z(n2998) );
  XOR U4689 ( .A(n3545), .B(n2998), .Z(out[310]) );
  IV U4690 ( .A(n2999), .Z(n3574) );
  NANDN U4691 ( .A(n3000), .B(n3574), .Z(n3001) );
  XOR U4692 ( .A(n3575), .B(n3001), .Z(out[311]) );
  IV U4693 ( .A(n3002), .Z(n3598) );
  NANDN U4694 ( .A(n3003), .B(n3598), .Z(n3004) );
  XOR U4695 ( .A(n3599), .B(n3004), .Z(out[312]) );
  NANDN U4696 ( .A(n3005), .B(n3628), .Z(n3006) );
  XOR U4697 ( .A(n3629), .B(n3006), .Z(out[313]) );
  NANDN U4698 ( .A(n3007), .B(n3672), .Z(n3008) );
  XOR U4699 ( .A(n3673), .B(n3008), .Z(out[314]) );
  NANDN U4700 ( .A(n3010), .B(n3009), .Z(n3011) );
  XOR U4701 ( .A(n3717), .B(n3011), .Z(out[315]) );
  NANDN U4702 ( .A(n3013), .B(n3012), .Z(n3014) );
  XOR U4703 ( .A(n3763), .B(n3014), .Z(out[316]) );
  NANDN U4704 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U4705 ( .A(n3851), .B(n3018), .Z(out[318]) );
  NANDN U4706 ( .A(n3020), .B(n3019), .Z(n3021) );
  XOR U4707 ( .A(n3895), .B(n3021), .Z(out[319]) );
  OR U4708 ( .A(n4992), .B(n3022), .Z(n3023) );
  XOR U4709 ( .A(n4993), .B(n3023), .Z(out[31]) );
  XOR U4710 ( .A(in[72]), .B(n4448), .Z(n3261) );
  XOR U4711 ( .A(in[1317]), .B(n4280), .Z(n3615) );
  XNOR U4712 ( .A(in[1244]), .B(n3024), .Z(n3612) );
  NANDN U4713 ( .A(n3615), .B(n3612), .Z(n3025) );
  XNOR U4714 ( .A(n3261), .B(n3025), .Z(out[320]) );
  XOR U4715 ( .A(in[73]), .B(n4451), .Z(n3147) );
  IV U4716 ( .A(n3147), .Z(n3264) );
  XOR U4717 ( .A(in[1318]), .B(n4286), .Z(n3619) );
  XNOR U4718 ( .A(in[1245]), .B(n3026), .Z(n3616) );
  NANDN U4719 ( .A(n3619), .B(n3616), .Z(n3027) );
  XOR U4720 ( .A(n3264), .B(n3027), .Z(out[321]) );
  XOR U4721 ( .A(in[74]), .B(n4454), .Z(n3149) );
  IV U4722 ( .A(n3149), .Z(n3271) );
  XOR U4723 ( .A(in[1319]), .B(n4288), .Z(n3623) );
  XNOR U4724 ( .A(in[1246]), .B(n3028), .Z(n3620) );
  NANDN U4725 ( .A(n3623), .B(n3620), .Z(n3029) );
  XOR U4726 ( .A(n3271), .B(n3029), .Z(out[322]) );
  XOR U4727 ( .A(in[75]), .B(n4457), .Z(n3151) );
  IV U4728 ( .A(n3151), .Z(n3274) );
  XOR U4729 ( .A(in[1320]), .B(n4290), .Z(n3627) );
  XNOR U4730 ( .A(in[1247]), .B(n3030), .Z(n3624) );
  NANDN U4731 ( .A(n3627), .B(n3624), .Z(n3031) );
  XOR U4732 ( .A(n3274), .B(n3031), .Z(out[323]) );
  XNOR U4733 ( .A(n4460), .B(in[76]), .Z(n3277) );
  XOR U4734 ( .A(in[1321]), .B(n4292), .Z(n3635) );
  XNOR U4735 ( .A(in[1248]), .B(n3032), .Z(n3632) );
  NANDN U4736 ( .A(n3635), .B(n3632), .Z(n3033) );
  XNOR U4737 ( .A(n3277), .B(n3033), .Z(out[324]) );
  XNOR U4738 ( .A(n4463), .B(in[77]), .Z(n3280) );
  XOR U4739 ( .A(in[1322]), .B(n4294), .Z(n3639) );
  XNOR U4740 ( .A(in[1249]), .B(n3034), .Z(n3636) );
  NANDN U4741 ( .A(n3639), .B(n3636), .Z(n3035) );
  XNOR U4742 ( .A(n3280), .B(n3035), .Z(out[325]) );
  XNOR U4743 ( .A(n4466), .B(in[78]), .Z(n3283) );
  XOR U4744 ( .A(in[1323]), .B(n4296), .Z(n3643) );
  XNOR U4745 ( .A(in[1250]), .B(n4124), .Z(n3640) );
  NANDN U4746 ( .A(n3643), .B(n3640), .Z(n3036) );
  XNOR U4747 ( .A(n3283), .B(n3036), .Z(out[326]) );
  XNOR U4748 ( .A(n4469), .B(in[79]), .Z(n3286) );
  XOR U4749 ( .A(in[1324]), .B(n4298), .Z(n3647) );
  XNOR U4750 ( .A(in[1251]), .B(n3037), .Z(n3644) );
  NANDN U4751 ( .A(n3647), .B(n3644), .Z(n3038) );
  XNOR U4752 ( .A(n3286), .B(n3038), .Z(out[327]) );
  XNOR U4753 ( .A(n4472), .B(in[80]), .Z(n3289) );
  XOR U4754 ( .A(in[1325]), .B(n4300), .Z(n3651) );
  XNOR U4755 ( .A(in[1252]), .B(n3039), .Z(n3648) );
  NANDN U4756 ( .A(n3651), .B(n3648), .Z(n3040) );
  XNOR U4757 ( .A(n3289), .B(n3040), .Z(out[328]) );
  XNOR U4758 ( .A(n4479), .B(in[81]), .Z(n3292) );
  XNOR U4759 ( .A(in[1253]), .B(n4136), .Z(n3653) );
  XNOR U4760 ( .A(in[1326]), .B(n4302), .Z(n3655) );
  NANDN U4761 ( .A(n3653), .B(n3655), .Z(n3041) );
  XNOR U4762 ( .A(n3292), .B(n3041), .Z(out[329]) );
  OR U4763 ( .A(n5036), .B(n3042), .Z(n3043) );
  XOR U4764 ( .A(n5037), .B(n3043), .Z(out[32]) );
  XNOR U4765 ( .A(n4482), .B(in[82]), .Z(n3295) );
  XNOR U4766 ( .A(in[1254]), .B(n4140), .Z(n3657) );
  XNOR U4767 ( .A(in[1327]), .B(n4304), .Z(n3659) );
  NANDN U4768 ( .A(n3657), .B(n3659), .Z(n3044) );
  XNOR U4769 ( .A(n3295), .B(n3044), .Z(out[330]) );
  XNOR U4770 ( .A(n4485), .B(in[83]), .Z(n3298) );
  XNOR U4771 ( .A(in[1255]), .B(n4144), .Z(n3661) );
  XNOR U4772 ( .A(in[1328]), .B(n4311), .Z(n3663) );
  NANDN U4773 ( .A(n3661), .B(n3663), .Z(n3045) );
  XNOR U4774 ( .A(n3298), .B(n3045), .Z(out[331]) );
  XNOR U4775 ( .A(in[84]), .B(n4488), .Z(n3305) );
  XNOR U4776 ( .A(in[1256]), .B(n4148), .Z(n3665) );
  XNOR U4777 ( .A(in[1329]), .B(n4314), .Z(n3667) );
  NANDN U4778 ( .A(n3665), .B(n3667), .Z(n3046) );
  XNOR U4779 ( .A(n3305), .B(n3046), .Z(out[332]) );
  XNOR U4780 ( .A(in[85]), .B(n4491), .Z(n3308) );
  XNOR U4781 ( .A(in[1257]), .B(n4152), .Z(n3669) );
  XNOR U4782 ( .A(in[1330]), .B(n4317), .Z(n3671) );
  NANDN U4783 ( .A(n3669), .B(n3671), .Z(n3047) );
  XNOR U4784 ( .A(n3308), .B(n3047), .Z(out[333]) );
  XNOR U4785 ( .A(in[86]), .B(n4494), .Z(n3311) );
  XNOR U4786 ( .A(in[1258]), .B(n4162), .Z(n3677) );
  XNOR U4787 ( .A(in[1331]), .B(n4320), .Z(n3679) );
  NANDN U4788 ( .A(n3677), .B(n3679), .Z(n3048) );
  XNOR U4789 ( .A(n3311), .B(n3048), .Z(out[334]) );
  XNOR U4790 ( .A(in[87]), .B(n4497), .Z(n3314) );
  XNOR U4791 ( .A(in[1259]), .B(n4166), .Z(n3681) );
  XNOR U4792 ( .A(in[1332]), .B(n4323), .Z(n3683) );
  NANDN U4793 ( .A(n3681), .B(n3683), .Z(n3049) );
  XNOR U4794 ( .A(n3314), .B(n3049), .Z(out[335]) );
  XNOR U4795 ( .A(in[88]), .B(n4500), .Z(n3317) );
  XNOR U4796 ( .A(in[1260]), .B(n4170), .Z(n3685) );
  XNOR U4797 ( .A(in[1333]), .B(n4326), .Z(n3687) );
  NANDN U4798 ( .A(n3685), .B(n3687), .Z(n3050) );
  XNOR U4799 ( .A(n3317), .B(n3050), .Z(out[336]) );
  XNOR U4800 ( .A(in[89]), .B(n4503), .Z(n3320) );
  XNOR U4801 ( .A(in[1261]), .B(n4174), .Z(n3689) );
  XNOR U4802 ( .A(in[1334]), .B(n4329), .Z(n3691) );
  NANDN U4803 ( .A(n3689), .B(n3691), .Z(n3051) );
  XNOR U4804 ( .A(n3320), .B(n3051), .Z(out[337]) );
  XNOR U4805 ( .A(in[90]), .B(n4506), .Z(n3322) );
  XNOR U4806 ( .A(in[1262]), .B(n3898), .Z(n3693) );
  XNOR U4807 ( .A(in[1335]), .B(n4332), .Z(n3695) );
  NANDN U4808 ( .A(n3693), .B(n3695), .Z(n3052) );
  XNOR U4809 ( .A(n3322), .B(n3052), .Z(out[338]) );
  XOR U4810 ( .A(in[91]), .B(n4513), .Z(n3324) );
  XNOR U4811 ( .A(in[1263]), .B(n3902), .Z(n3697) );
  XNOR U4812 ( .A(in[1336]), .B(n4178), .Z(n3699) );
  NANDN U4813 ( .A(n3697), .B(n3699), .Z(n3053) );
  XNOR U4814 ( .A(n3324), .B(n3053), .Z(out[339]) );
  OR U4815 ( .A(n5077), .B(n3054), .Z(n3055) );
  XOR U4816 ( .A(n5078), .B(n3055), .Z(out[33]) );
  XOR U4817 ( .A(in[92]), .B(n4516), .Z(n3326) );
  XNOR U4818 ( .A(in[1264]), .B(n3906), .Z(n3701) );
  XNOR U4819 ( .A(in[1337]), .B(n4181), .Z(n3703) );
  NANDN U4820 ( .A(n3701), .B(n3703), .Z(n3056) );
  XNOR U4821 ( .A(n3326), .B(n3056), .Z(out[340]) );
  XOR U4822 ( .A(in[93]), .B(n4519), .Z(n3328) );
  XNOR U4823 ( .A(in[1265]), .B(n3910), .Z(n3705) );
  XNOR U4824 ( .A(in[1338]), .B(n4184), .Z(n3707) );
  NANDN U4825 ( .A(n3705), .B(n3707), .Z(n3057) );
  XNOR U4826 ( .A(n3328), .B(n3057), .Z(out[341]) );
  XNOR U4827 ( .A(in[94]), .B(n4522), .Z(n3334) );
  XNOR U4828 ( .A(in[1266]), .B(n3914), .Z(n3709) );
  XNOR U4829 ( .A(in[1339]), .B(n4187), .Z(n3711) );
  NANDN U4830 ( .A(n3709), .B(n3711), .Z(n3058) );
  XNOR U4831 ( .A(n3334), .B(n3058), .Z(out[342]) );
  XNOR U4832 ( .A(in[95]), .B(n4526), .Z(n3336) );
  XOR U4833 ( .A(in[1267]), .B(n3918), .Z(n3713) );
  XNOR U4834 ( .A(in[1340]), .B(n3059), .Z(n3715) );
  NANDN U4835 ( .A(n3713), .B(n3715), .Z(n3060) );
  XNOR U4836 ( .A(n3336), .B(n3060), .Z(out[343]) );
  XNOR U4837 ( .A(in[96]), .B(n4530), .Z(n3338) );
  XOR U4838 ( .A(in[1268]), .B(n3922), .Z(n3723) );
  XNOR U4839 ( .A(in[1341]), .B(n3061), .Z(n3725) );
  NANDN U4840 ( .A(n3723), .B(n3725), .Z(n3062) );
  XNOR U4841 ( .A(n3338), .B(n3062), .Z(out[344]) );
  XNOR U4842 ( .A(in[97]), .B(n4534), .Z(n3340) );
  XOR U4843 ( .A(in[1269]), .B(n3926), .Z(n3727) );
  XNOR U4844 ( .A(in[1342]), .B(n3063), .Z(n3729) );
  NANDN U4845 ( .A(n3727), .B(n3729), .Z(n3064) );
  XNOR U4846 ( .A(n3340), .B(n3064), .Z(out[345]) );
  XNOR U4847 ( .A(in[98]), .B(n4538), .Z(n3342) );
  IV U4848 ( .A(n3065), .Z(n3930) );
  XOR U4849 ( .A(in[1270]), .B(n3930), .Z(n3731) );
  XNOR U4850 ( .A(in[1343]), .B(n4199), .Z(n3733) );
  NANDN U4851 ( .A(n3731), .B(n3733), .Z(n3066) );
  XNOR U4852 ( .A(n3342), .B(n3066), .Z(out[346]) );
  XNOR U4853 ( .A(in[99]), .B(n4542), .Z(n3344) );
  IV U4854 ( .A(n3067), .Z(n3934) );
  XOR U4855 ( .A(in[1271]), .B(n3934), .Z(n3735) );
  XNOR U4856 ( .A(in[1280]), .B(n3068), .Z(n3737) );
  NANDN U4857 ( .A(n3735), .B(n3737), .Z(n3069) );
  XNOR U4858 ( .A(n3344), .B(n3069), .Z(out[347]) );
  XOR U4859 ( .A(in[100]), .B(n4546), .Z(n3197) );
  IV U4860 ( .A(n3197), .Z(n3347) );
  IV U4861 ( .A(n3070), .Z(n3941) );
  XOR U4862 ( .A(in[1272]), .B(n3941), .Z(n3739) );
  XNOR U4863 ( .A(in[1281]), .B(n3071), .Z(n3741) );
  NANDN U4864 ( .A(n3739), .B(n3741), .Z(n3072) );
  XOR U4865 ( .A(n3347), .B(n3072), .Z(out[348]) );
  XOR U4866 ( .A(in[101]), .B(n4552), .Z(n3200) );
  IV U4867 ( .A(n3200), .Z(n3351) );
  XOR U4868 ( .A(in[1273]), .B(n3945), .Z(n3743) );
  XNOR U4869 ( .A(in[1282]), .B(n3073), .Z(n3745) );
  NANDN U4870 ( .A(n3743), .B(n3745), .Z(n3074) );
  XOR U4871 ( .A(n3351), .B(n3074), .Z(out[349]) );
  OR U4872 ( .A(n5113), .B(n3075), .Z(n3076) );
  XNOR U4873 ( .A(n5112), .B(n3076), .Z(out[34]) );
  XOR U4874 ( .A(in[102]), .B(n4554), .Z(n3203) );
  IV U4875 ( .A(n3203), .Z(n3354) );
  XOR U4876 ( .A(in[1274]), .B(n3949), .Z(n3747) );
  XNOR U4877 ( .A(in[1283]), .B(n3077), .Z(n3749) );
  NANDN U4878 ( .A(n3747), .B(n3749), .Z(n3078) );
  XOR U4879 ( .A(n3354), .B(n3078), .Z(out[350]) );
  XOR U4880 ( .A(in[103]), .B(n4335), .Z(n3206) );
  IV U4881 ( .A(n3206), .Z(n3357) );
  XNOR U4882 ( .A(in[1275]), .B(n3953), .Z(n3751) );
  XNOR U4883 ( .A(in[1284]), .B(n3079), .Z(n3753) );
  NANDN U4884 ( .A(n3751), .B(n3753), .Z(n3080) );
  XOR U4885 ( .A(n3357), .B(n3080), .Z(out[351]) );
  XOR U4886 ( .A(in[104]), .B(n4337), .Z(n3209) );
  IV U4887 ( .A(n3209), .Z(n3364) );
  XNOR U4888 ( .A(in[1276]), .B(n3957), .Z(n3755) );
  XNOR U4889 ( .A(in[1285]), .B(n3081), .Z(n3757) );
  NANDN U4890 ( .A(n3755), .B(n3757), .Z(n3082) );
  XOR U4891 ( .A(n3364), .B(n3082), .Z(out[352]) );
  XOR U4892 ( .A(in[105]), .B(n4343), .Z(n3212) );
  IV U4893 ( .A(n3212), .Z(n3367) );
  XNOR U4894 ( .A(in[1277]), .B(n3961), .Z(n3759) );
  XNOR U4895 ( .A(in[1286]), .B(n3083), .Z(n3761) );
  NANDN U4896 ( .A(n3759), .B(n3761), .Z(n3084) );
  XOR U4897 ( .A(n3367), .B(n3084), .Z(out[353]) );
  XOR U4898 ( .A(in[106]), .B(n4345), .Z(n3215) );
  IV U4899 ( .A(n3215), .Z(n3370) );
  XNOR U4900 ( .A(in[1278]), .B(n3965), .Z(n3767) );
  XNOR U4901 ( .A(in[1287]), .B(n3085), .Z(n3769) );
  NANDN U4902 ( .A(n3767), .B(n3769), .Z(n3086) );
  XOR U4903 ( .A(n3370), .B(n3086), .Z(out[354]) );
  XOR U4904 ( .A(in[107]), .B(n4347), .Z(n3218) );
  IV U4905 ( .A(n3218), .Z(n3373) );
  XNOR U4906 ( .A(in[1279]), .B(n3969), .Z(n3771) );
  XNOR U4907 ( .A(in[1288]), .B(n4216), .Z(n3773) );
  NANDN U4908 ( .A(n3771), .B(n3773), .Z(n3087) );
  XOR U4909 ( .A(n3373), .B(n3087), .Z(out[355]) );
  XOR U4910 ( .A(in[108]), .B(n4350), .Z(n3224) );
  IV U4911 ( .A(n3224), .Z(n3375) );
  XNOR U4912 ( .A(in[1216]), .B(n3973), .Z(n3775) );
  XNOR U4913 ( .A(in[1289]), .B(n3088), .Z(n3777) );
  NANDN U4914 ( .A(n3775), .B(n3777), .Z(n3089) );
  XOR U4915 ( .A(n3375), .B(n3089), .Z(out[356]) );
  XOR U4916 ( .A(in[109]), .B(n4353), .Z(n3226) );
  IV U4917 ( .A(n3226), .Z(n3377) );
  XNOR U4918 ( .A(in[1217]), .B(n3977), .Z(n3779) );
  XNOR U4919 ( .A(in[1290]), .B(n3090), .Z(n3781) );
  NANDN U4920 ( .A(n3779), .B(n3781), .Z(n3091) );
  XOR U4921 ( .A(n3377), .B(n3091), .Z(out[357]) );
  XOR U4922 ( .A(in[110]), .B(n4356), .Z(n3228) );
  IV U4923 ( .A(n3228), .Z(n3379) );
  XNOR U4924 ( .A(in[1218]), .B(n3984), .Z(n3783) );
  XNOR U4925 ( .A(in[1291]), .B(n3092), .Z(n3785) );
  NANDN U4926 ( .A(n3783), .B(n3785), .Z(n3093) );
  XOR U4927 ( .A(n3379), .B(n3093), .Z(out[358]) );
  XOR U4928 ( .A(in[111]), .B(n4358), .Z(n3230) );
  IV U4929 ( .A(n3230), .Z(n3381) );
  XNOR U4930 ( .A(in[1219]), .B(n3988), .Z(n3787) );
  XNOR U4931 ( .A(in[1292]), .B(n3094), .Z(n3789) );
  NANDN U4932 ( .A(n3787), .B(n3789), .Z(n3095) );
  XOR U4933 ( .A(n3381), .B(n3095), .Z(out[359]) );
  OR U4934 ( .A(n5156), .B(n3096), .Z(n3097) );
  XNOR U4935 ( .A(n5155), .B(n3097), .Z(out[35]) );
  XOR U4936 ( .A(in[112]), .B(n4361), .Z(n3232) );
  IV U4937 ( .A(n3232), .Z(n3383) );
  XOR U4938 ( .A(in[1293]), .B(n3098), .Z(n3793) );
  XOR U4939 ( .A(in[1220]), .B(n3992), .Z(n3790) );
  NANDN U4940 ( .A(n3793), .B(n3790), .Z(n3099) );
  XOR U4941 ( .A(n3383), .B(n3099), .Z(out[360]) );
  XOR U4942 ( .A(in[113]), .B(n4364), .Z(n3234) );
  IV U4943 ( .A(n3234), .Z(n3385) );
  XOR U4944 ( .A(in[1294]), .B(n4234), .Z(n3797) );
  XOR U4945 ( .A(in[1221]), .B(n3996), .Z(n3794) );
  NANDN U4946 ( .A(n3797), .B(n3794), .Z(n3100) );
  XOR U4947 ( .A(n3385), .B(n3100), .Z(out[361]) );
  XOR U4948 ( .A(in[114]), .B(n4367), .Z(n3236) );
  IV U4949 ( .A(n3236), .Z(n3391) );
  XOR U4950 ( .A(in[1295]), .B(n4237), .Z(n3801) );
  XOR U4951 ( .A(in[1222]), .B(n4000), .Z(n3798) );
  NANDN U4952 ( .A(n3801), .B(n3798), .Z(n3101) );
  XOR U4953 ( .A(n3391), .B(n3101), .Z(out[362]) );
  XOR U4954 ( .A(in[115]), .B(n4374), .Z(n3238) );
  IV U4955 ( .A(n3238), .Z(n3393) );
  XOR U4956 ( .A(in[1296]), .B(n4240), .Z(n3805) );
  XOR U4957 ( .A(in[1223]), .B(n4004), .Z(n3802) );
  NANDN U4958 ( .A(n3805), .B(n3802), .Z(n3102) );
  XOR U4959 ( .A(n3393), .B(n3102), .Z(out[363]) );
  XOR U4960 ( .A(in[116]), .B(n4377), .Z(n3240) );
  IV U4961 ( .A(n3240), .Z(n3396) );
  XOR U4962 ( .A(in[1297]), .B(n4241), .Z(n3813) );
  XOR U4963 ( .A(in[1224]), .B(n4008), .Z(n3810) );
  NANDN U4964 ( .A(n3813), .B(n3810), .Z(n3103) );
  XOR U4965 ( .A(n3396), .B(n3103), .Z(out[364]) );
  XOR U4966 ( .A(in[117]), .B(n4380), .Z(n3242) );
  IV U4967 ( .A(n3242), .Z(n3400) );
  XOR U4968 ( .A(in[1298]), .B(n3104), .Z(n3817) );
  XOR U4969 ( .A(in[1225]), .B(n4012), .Z(n3814) );
  NANDN U4970 ( .A(n3817), .B(n3814), .Z(n3105) );
  XOR U4971 ( .A(n3400), .B(n3105), .Z(out[365]) );
  XOR U4972 ( .A(in[118]), .B(n4383), .Z(n3248) );
  IV U4973 ( .A(n3248), .Z(n3404) );
  XOR U4974 ( .A(in[1299]), .B(n3106), .Z(n3821) );
  XOR U4975 ( .A(in[1226]), .B(n4016), .Z(n3818) );
  NANDN U4976 ( .A(n3821), .B(n3818), .Z(n3107) );
  XOR U4977 ( .A(n3404), .B(n3107), .Z(out[366]) );
  XOR U4978 ( .A(in[119]), .B(n4386), .Z(n3250) );
  IV U4979 ( .A(n3250), .Z(n3408) );
  XOR U4980 ( .A(in[1300]), .B(n4248), .Z(n3825) );
  XOR U4981 ( .A(in[1227]), .B(n4020), .Z(n3822) );
  NANDN U4982 ( .A(n3825), .B(n3822), .Z(n3108) );
  XOR U4983 ( .A(n3408), .B(n3108), .Z(out[367]) );
  XOR U4984 ( .A(in[120]), .B(n4388), .Z(n3252) );
  IV U4985 ( .A(n3252), .Z(n3411) );
  XOR U4986 ( .A(in[1301]), .B(n4251), .Z(n3829) );
  XOR U4987 ( .A(in[1228]), .B(n4028), .Z(n3826) );
  NANDN U4988 ( .A(n3829), .B(n3826), .Z(n3109) );
  XOR U4989 ( .A(n3411), .B(n3109), .Z(out[368]) );
  XOR U4990 ( .A(in[121]), .B(n4391), .Z(n3254) );
  IV U4991 ( .A(n3254), .Z(n3414) );
  XOR U4992 ( .A(in[1302]), .B(n4252), .Z(n3833) );
  XNOR U4993 ( .A(in[1229]), .B(n3110), .Z(n3830) );
  NANDN U4994 ( .A(n3833), .B(n3830), .Z(n3111) );
  XOR U4995 ( .A(n3414), .B(n3111), .Z(out[369]) );
  ANDN U4996 ( .B(n3113), .A(n3112), .Z(n3114) );
  XOR U4997 ( .A(n3115), .B(n3114), .Z(out[36]) );
  XOR U4998 ( .A(in[122]), .B(n4394), .Z(n3417) );
  XOR U4999 ( .A(in[1303]), .B(n4253), .Z(n3837) );
  XNOR U5000 ( .A(in[1230]), .B(n3116), .Z(n3834) );
  NANDN U5001 ( .A(n3837), .B(n3834), .Z(n3117) );
  XOR U5002 ( .A(n3417), .B(n3117), .Z(out[370]) );
  XOR U5003 ( .A(in[123]), .B(n4397), .Z(n3420) );
  XOR U5004 ( .A(in[1304]), .B(n4254), .Z(n3841) );
  XNOR U5005 ( .A(in[1231]), .B(n3118), .Z(n3838) );
  NANDN U5006 ( .A(n3841), .B(n3838), .Z(n3119) );
  XOR U5007 ( .A(n3420), .B(n3119), .Z(out[371]) );
  XOR U5008 ( .A(in[124]), .B(n4400), .Z(n3428) );
  XOR U5009 ( .A(in[1305]), .B(n4255), .Z(n3845) );
  XNOR U5010 ( .A(in[1232]), .B(n3120), .Z(n3842) );
  NANDN U5011 ( .A(n3845), .B(n3842), .Z(n3121) );
  XNOR U5012 ( .A(n3428), .B(n3121), .Z(out[372]) );
  XOR U5013 ( .A(in[125]), .B(n4407), .Z(n3431) );
  XOR U5014 ( .A(in[1306]), .B(n4256), .Z(n3849) );
  XNOR U5015 ( .A(in[1233]), .B(n4048), .Z(n3846) );
  NANDN U5016 ( .A(n3849), .B(n3846), .Z(n3122) );
  XNOR U5017 ( .A(n3431), .B(n3122), .Z(out[373]) );
  XOR U5018 ( .A(in[126]), .B(n4410), .Z(n3434) );
  XOR U5019 ( .A(in[1307]), .B(n4257), .Z(n3857) );
  XOR U5020 ( .A(in[1234]), .B(n4052), .Z(n3854) );
  NANDN U5021 ( .A(n3857), .B(n3854), .Z(n3123) );
  XNOR U5022 ( .A(n3434), .B(n3123), .Z(out[374]) );
  XOR U5023 ( .A(in[127]), .B(n4413), .Z(n3437) );
  XOR U5024 ( .A(in[1308]), .B(n4260), .Z(n3861) );
  XNOR U5025 ( .A(in[1235]), .B(n3124), .Z(n3858) );
  NANDN U5026 ( .A(n3861), .B(n3858), .Z(n3125) );
  XNOR U5027 ( .A(n3437), .B(n3125), .Z(out[375]) );
  XOR U5028 ( .A(in[64]), .B(n4416), .Z(n3440) );
  XOR U5029 ( .A(in[1309]), .B(n4261), .Z(n3865) );
  XNOR U5030 ( .A(in[1236]), .B(n3126), .Z(n3862) );
  NANDN U5031 ( .A(n3865), .B(n3862), .Z(n3127) );
  XNOR U5032 ( .A(n3440), .B(n3127), .Z(out[376]) );
  XOR U5033 ( .A(in[65]), .B(n4419), .Z(n3443) );
  XOR U5034 ( .A(in[1310]), .B(n4262), .Z(n3869) );
  XNOR U5035 ( .A(in[1237]), .B(n3128), .Z(n3866) );
  NANDN U5036 ( .A(n3869), .B(n3866), .Z(n3129) );
  XNOR U5037 ( .A(n3443), .B(n3129), .Z(out[377]) );
  XOR U5038 ( .A(in[66]), .B(n4422), .Z(n3446) );
  XOR U5039 ( .A(in[1311]), .B(n4263), .Z(n3873) );
  XNOR U5040 ( .A(in[1238]), .B(n3130), .Z(n3870) );
  NANDN U5041 ( .A(n3873), .B(n3870), .Z(n3131) );
  XNOR U5042 ( .A(n3446), .B(n3131), .Z(out[378]) );
  XOR U5043 ( .A(in[67]), .B(n4425), .Z(n3449) );
  XOR U5044 ( .A(in[1312]), .B(n4266), .Z(n3877) );
  XNOR U5045 ( .A(in[1239]), .B(n3132), .Z(n3874) );
  NANDN U5046 ( .A(n3877), .B(n3874), .Z(n3133) );
  XNOR U5047 ( .A(n3449), .B(n3133), .Z(out[379]) );
  ANDN U5048 ( .B(n3135), .A(n3134), .Z(n3136) );
  XOR U5049 ( .A(n3137), .B(n3136), .Z(out[37]) );
  XOR U5050 ( .A(in[68]), .B(n4428), .Z(n3452) );
  XOR U5051 ( .A(in[1313]), .B(n4269), .Z(n3881) );
  XNOR U5052 ( .A(in[1240]), .B(n3138), .Z(n3878) );
  NANDN U5053 ( .A(n3881), .B(n3878), .Z(n3139) );
  XNOR U5054 ( .A(n3452), .B(n3139), .Z(out[380]) );
  XOR U5055 ( .A(in[69]), .B(n4431), .Z(n3455) );
  XOR U5056 ( .A(in[1314]), .B(n4272), .Z(n3885) );
  XNOR U5057 ( .A(in[1241]), .B(n3140), .Z(n3882) );
  NANDN U5058 ( .A(n3885), .B(n3882), .Z(n3141) );
  XNOR U5059 ( .A(n3455), .B(n3141), .Z(out[381]) );
  XOR U5060 ( .A(in[70]), .B(n4434), .Z(n3462) );
  XOR U5061 ( .A(in[1315]), .B(n3142), .Z(n3889) );
  XNOR U5062 ( .A(in[1242]), .B(n3143), .Z(n3886) );
  NANDN U5063 ( .A(n3889), .B(n3886), .Z(n3144) );
  XOR U5064 ( .A(n3462), .B(n3144), .Z(out[382]) );
  XOR U5065 ( .A(in[71]), .B(n4445), .Z(n3465) );
  XOR U5066 ( .A(in[1316]), .B(n4278), .Z(n3893) );
  XNOR U5067 ( .A(in[1243]), .B(n3145), .Z(n3890) );
  NANDN U5068 ( .A(n3893), .B(n3890), .Z(n3146) );
  XNOR U5069 ( .A(n3465), .B(n3146), .Z(out[383]) );
  XOR U5070 ( .A(in[497]), .B(n4137), .Z(n3467) );
  XOR U5071 ( .A(in[498]), .B(n4141), .Z(n3469) );
  ANDN U5072 ( .B(n3619), .A(n3147), .Z(n3148) );
  XNOR U5073 ( .A(n3469), .B(n3148), .Z(out[385]) );
  XOR U5074 ( .A(in[499]), .B(n4145), .Z(n3471) );
  ANDN U5075 ( .B(n3623), .A(n3149), .Z(n3150) );
  XNOR U5076 ( .A(n3471), .B(n3150), .Z(out[386]) );
  XOR U5077 ( .A(in[500]), .B(n4149), .Z(n3473) );
  ANDN U5078 ( .B(n3627), .A(n3151), .Z(n3152) );
  XNOR U5079 ( .A(n3473), .B(n3152), .Z(out[387]) );
  XOR U5080 ( .A(in[501]), .B(n4153), .Z(n3475) );
  XOR U5081 ( .A(in[502]), .B(n4163), .Z(n3476) );
  NOR U5082 ( .A(n3154), .B(n3153), .Z(n3155) );
  XOR U5083 ( .A(n3156), .B(n3155), .Z(out[38]) );
  XOR U5084 ( .A(in[503]), .B(n4167), .Z(n3477) );
  XOR U5085 ( .A(in[504]), .B(n4171), .Z(n3478) );
  XOR U5086 ( .A(in[505]), .B(n4175), .Z(n3483) );
  XOR U5087 ( .A(in[506]), .B(n3899), .Z(n3484) );
  NOR U5088 ( .A(n3655), .B(n3292), .Z(n3157) );
  XNOR U5089 ( .A(n3484), .B(n3157), .Z(out[393]) );
  XOR U5090 ( .A(in[507]), .B(n3903), .Z(n3486) );
  NOR U5091 ( .A(n3659), .B(n3295), .Z(n3158) );
  XNOR U5092 ( .A(n3486), .B(n3158), .Z(out[394]) );
  XOR U5093 ( .A(in[508]), .B(n3907), .Z(n3488) );
  NOR U5094 ( .A(n3663), .B(n3298), .Z(n3159) );
  XNOR U5095 ( .A(n3488), .B(n3159), .Z(out[395]) );
  XOR U5096 ( .A(in[509]), .B(n3911), .Z(n3490) );
  NOR U5097 ( .A(n3667), .B(n3305), .Z(n3160) );
  XNOR U5098 ( .A(n3490), .B(n3160), .Z(out[396]) );
  XOR U5099 ( .A(in[510]), .B(n3915), .Z(n3492) );
  NOR U5100 ( .A(n3671), .B(n3308), .Z(n3161) );
  XNOR U5101 ( .A(n3492), .B(n3161), .Z(out[397]) );
  XOR U5102 ( .A(in[511]), .B(n3919), .Z(n3494) );
  NOR U5103 ( .A(n3679), .B(n3311), .Z(n3162) );
  XNOR U5104 ( .A(n3494), .B(n3162), .Z(out[398]) );
  XOR U5105 ( .A(in[448]), .B(n3923), .Z(n3496) );
  NOR U5106 ( .A(n3683), .B(n3314), .Z(n3163) );
  XNOR U5107 ( .A(n3496), .B(n3163), .Z(out[399]) );
  ANDN U5108 ( .B(n3165), .A(n3164), .Z(n3166) );
  XOR U5109 ( .A(n3167), .B(n3166), .Z(out[39]) );
  OR U5110 ( .A(n4069), .B(n3168), .Z(n3169) );
  XNOR U5111 ( .A(n4068), .B(n3169), .Z(out[3]) );
  XOR U5112 ( .A(in[449]), .B(n3927), .Z(n3498) );
  NOR U5113 ( .A(n3687), .B(n3317), .Z(n3170) );
  XNOR U5114 ( .A(n3498), .B(n3170), .Z(out[400]) );
  XOR U5115 ( .A(n3171), .B(in[450]), .Z(n3500) );
  NOR U5116 ( .A(n3691), .B(n3320), .Z(n3172) );
  XOR U5117 ( .A(n3500), .B(n3172), .Z(out[401]) );
  XOR U5118 ( .A(n3173), .B(in[451]), .Z(n3505) );
  NOR U5119 ( .A(n3695), .B(n3322), .Z(n3174) );
  XOR U5120 ( .A(n3505), .B(n3174), .Z(out[402]) );
  XOR U5121 ( .A(n3175), .B(in[452]), .Z(n3506) );
  NOR U5122 ( .A(n3699), .B(n3324), .Z(n3176) );
  XOR U5123 ( .A(n3506), .B(n3176), .Z(out[403]) );
  XOR U5124 ( .A(n3177), .B(in[453]), .Z(n3507) );
  NOR U5125 ( .A(n3703), .B(n3326), .Z(n3178) );
  XOR U5126 ( .A(n3507), .B(n3178), .Z(out[404]) );
  XOR U5127 ( .A(n3179), .B(in[454]), .Z(n3508) );
  NOR U5128 ( .A(n3707), .B(n3328), .Z(n3180) );
  XOR U5129 ( .A(n3508), .B(n3180), .Z(out[405]) );
  XOR U5130 ( .A(n3181), .B(in[455]), .Z(n3509) );
  NOR U5131 ( .A(n3711), .B(n3334), .Z(n3182) );
  XOR U5132 ( .A(n3509), .B(n3182), .Z(out[406]) );
  XOR U5133 ( .A(n3183), .B(in[456]), .Z(n3510) );
  NOR U5134 ( .A(n3715), .B(n3336), .Z(n3184) );
  XOR U5135 ( .A(n3510), .B(n3184), .Z(out[407]) );
  XOR U5136 ( .A(in[457]), .B(n3185), .Z(n3511) );
  NOR U5137 ( .A(n3725), .B(n3338), .Z(n3186) );
  XOR U5138 ( .A(n3511), .B(n3186), .Z(out[408]) );
  XOR U5139 ( .A(n3187), .B(in[458]), .Z(n3512) );
  NOR U5140 ( .A(n3729), .B(n3340), .Z(n3188) );
  XOR U5141 ( .A(n3512), .B(n3188), .Z(out[409]) );
  ANDN U5142 ( .B(n3190), .A(n3189), .Z(n3191) );
  XNOR U5143 ( .A(n3192), .B(n3191), .Z(out[40]) );
  XOR U5144 ( .A(n3971), .B(in[459]), .Z(n3513) );
  NOR U5145 ( .A(n3733), .B(n3342), .Z(n3193) );
  XNOR U5146 ( .A(n3513), .B(n3193), .Z(out[410]) );
  XOR U5147 ( .A(in[460]), .B(n3194), .Z(n3515) );
  NOR U5148 ( .A(n3737), .B(n3344), .Z(n3195) );
  XOR U5149 ( .A(n3515), .B(n3195), .Z(out[411]) );
  XOR U5150 ( .A(in[461]), .B(n3196), .Z(n3346) );
  NOR U5151 ( .A(n3197), .B(n3741), .Z(n3198) );
  XOR U5152 ( .A(n3346), .B(n3198), .Z(out[412]) );
  XOR U5153 ( .A(in[462]), .B(n3199), .Z(n3350) );
  NOR U5154 ( .A(n3200), .B(n3745), .Z(n3201) );
  XOR U5155 ( .A(n3350), .B(n3201), .Z(out[413]) );
  XOR U5156 ( .A(in[463]), .B(n3202), .Z(n3353) );
  NOR U5157 ( .A(n3203), .B(n3749), .Z(n3204) );
  XOR U5158 ( .A(n3353), .B(n3204), .Z(out[414]) );
  XOR U5159 ( .A(in[464]), .B(n3205), .Z(n3356) );
  NOR U5160 ( .A(n3206), .B(n3753), .Z(n3207) );
  XOR U5161 ( .A(n3356), .B(n3207), .Z(out[415]) );
  XOR U5162 ( .A(in[465]), .B(n3208), .Z(n3363) );
  NOR U5163 ( .A(n3209), .B(n3757), .Z(n3210) );
  XOR U5164 ( .A(n3363), .B(n3210), .Z(out[416]) );
  XOR U5165 ( .A(in[466]), .B(n3211), .Z(n3366) );
  NOR U5166 ( .A(n3212), .B(n3761), .Z(n3213) );
  XOR U5167 ( .A(n3366), .B(n3213), .Z(out[417]) );
  XOR U5168 ( .A(in[467]), .B(n3214), .Z(n3369) );
  NOR U5169 ( .A(n3215), .B(n3769), .Z(n3216) );
  XOR U5170 ( .A(n3369), .B(n3216), .Z(out[418]) );
  XOR U5171 ( .A(in[468]), .B(n3217), .Z(n3372) );
  NOR U5172 ( .A(n3218), .B(n3773), .Z(n3219) );
  XOR U5173 ( .A(n3372), .B(n3219), .Z(out[419]) );
  AND U5174 ( .A(n3221), .B(n3220), .Z(n3222) );
  XNOR U5175 ( .A(n3223), .B(n3222), .Z(out[41]) );
  XOR U5176 ( .A(in[469]), .B(n4014), .Z(n3540) );
  NOR U5177 ( .A(n3224), .B(n3777), .Z(n3225) );
  XNOR U5178 ( .A(n3540), .B(n3225), .Z(out[420]) );
  XOR U5179 ( .A(in[470]), .B(n4018), .Z(n3542) );
  NOR U5180 ( .A(n3226), .B(n3781), .Z(n3227) );
  XNOR U5181 ( .A(n3542), .B(n3227), .Z(out[421]) );
  XOR U5182 ( .A(in[471]), .B(n4022), .Z(n3549) );
  NOR U5183 ( .A(n3228), .B(n3785), .Z(n3229) );
  XNOR U5184 ( .A(n3549), .B(n3229), .Z(out[422]) );
  XOR U5185 ( .A(in[472]), .B(n4030), .Z(n3552) );
  NOR U5186 ( .A(n3230), .B(n3789), .Z(n3231) );
  XNOR U5187 ( .A(n3552), .B(n3231), .Z(out[423]) );
  XOR U5188 ( .A(in[473]), .B(n4034), .Z(n3555) );
  ANDN U5189 ( .B(n3793), .A(n3232), .Z(n3233) );
  XNOR U5190 ( .A(n3555), .B(n3233), .Z(out[424]) );
  XOR U5191 ( .A(in[474]), .B(n4038), .Z(n3558) );
  ANDN U5192 ( .B(n3797), .A(n3234), .Z(n3235) );
  XNOR U5193 ( .A(n3558), .B(n3235), .Z(out[425]) );
  XOR U5194 ( .A(in[475]), .B(n4042), .Z(n3561) );
  ANDN U5195 ( .B(n3801), .A(n3236), .Z(n3237) );
  XNOR U5196 ( .A(n3561), .B(n3237), .Z(out[426]) );
  XOR U5197 ( .A(in[476]), .B(n4046), .Z(n3564) );
  ANDN U5198 ( .B(n3805), .A(n3238), .Z(n3239) );
  XNOR U5199 ( .A(n3564), .B(n3239), .Z(out[427]) );
  XOR U5200 ( .A(in[477]), .B(n4050), .Z(n3566) );
  ANDN U5201 ( .B(n3813), .A(n3240), .Z(n3241) );
  XNOR U5202 ( .A(n3566), .B(n3241), .Z(out[428]) );
  XOR U5203 ( .A(in[478]), .B(n4054), .Z(n3399) );
  ANDN U5204 ( .B(n3817), .A(n3242), .Z(n3243) );
  XOR U5205 ( .A(n3399), .B(n3243), .Z(out[429]) );
  AND U5206 ( .A(n3245), .B(n3244), .Z(n3246) );
  XNOR U5207 ( .A(n3247), .B(n3246), .Z(out[42]) );
  XOR U5208 ( .A(in[479]), .B(n4058), .Z(n3403) );
  ANDN U5209 ( .B(n3821), .A(n3248), .Z(n3249) );
  XOR U5210 ( .A(n3403), .B(n3249), .Z(out[430]) );
  XOR U5211 ( .A(in[480]), .B(n4062), .Z(n3407) );
  ANDN U5212 ( .B(n3825), .A(n3250), .Z(n3251) );
  XOR U5213 ( .A(n3407), .B(n3251), .Z(out[431]) );
  XOR U5214 ( .A(in[481]), .B(n4066), .Z(n3410) );
  ANDN U5215 ( .B(n3829), .A(n3252), .Z(n3253) );
  XOR U5216 ( .A(n3410), .B(n3253), .Z(out[432]) );
  XOR U5217 ( .A(in[482]), .B(n4074), .Z(n3413) );
  ANDN U5218 ( .B(n3833), .A(n3254), .Z(n3255) );
  XOR U5219 ( .A(n3413), .B(n3255), .Z(out[433]) );
  XOR U5220 ( .A(in[483]), .B(n4078), .Z(n3416) );
  XOR U5221 ( .A(in[484]), .B(n4082), .Z(n3419) );
  XOR U5222 ( .A(in[485]), .B(n4086), .Z(n3586) );
  XOR U5223 ( .A(in[486]), .B(n4089), .Z(n3588) );
  XOR U5224 ( .A(in[487]), .B(n4093), .Z(n3590) );
  XOR U5225 ( .A(in[488]), .B(n4097), .Z(n3592) );
  AND U5226 ( .A(n3257), .B(n3256), .Z(n3258) );
  XNOR U5227 ( .A(n3259), .B(n3258), .Z(out[43]) );
  XOR U5228 ( .A(in[489]), .B(n4101), .Z(n3594) );
  XOR U5229 ( .A(in[490]), .B(n4105), .Z(n3596) );
  XOR U5230 ( .A(in[491]), .B(n4109), .Z(n3602) );
  XOR U5231 ( .A(in[492]), .B(n4117), .Z(n3603) );
  XOR U5232 ( .A(in[493]), .B(n4121), .Z(n3604) );
  XOR U5233 ( .A(in[494]), .B(n4125), .Z(n3606) );
  XOR U5234 ( .A(in[495]), .B(n4129), .Z(n3608) );
  XOR U5235 ( .A(in[496]), .B(n4133), .Z(n3610) );
  XOR U5236 ( .A(in[886]), .B(n3260), .Z(n3613) );
  NAND U5237 ( .A(n3261), .B(n3467), .Z(n3262) );
  XOR U5238 ( .A(n3613), .B(n3262), .Z(out[448]) );
  XOR U5239 ( .A(in[887]), .B(n3263), .Z(n3617) );
  NANDN U5240 ( .A(n3264), .B(n3469), .Z(n3265) );
  XOR U5241 ( .A(n3617), .B(n3265), .Z(out[449]) );
  AND U5242 ( .A(n3267), .B(n3266), .Z(n3268) );
  XNOR U5243 ( .A(n3269), .B(n3268), .Z(out[44]) );
  XOR U5244 ( .A(in[888]), .B(n3270), .Z(n3621) );
  NANDN U5245 ( .A(n3271), .B(n3471), .Z(n3272) );
  XOR U5246 ( .A(n3621), .B(n3272), .Z(out[450]) );
  XOR U5247 ( .A(in[889]), .B(n3273), .Z(n3625) );
  NANDN U5248 ( .A(n3274), .B(n3473), .Z(n3275) );
  XOR U5249 ( .A(n3625), .B(n3275), .Z(out[451]) );
  XOR U5250 ( .A(in[890]), .B(n3276), .Z(n3633) );
  NANDN U5251 ( .A(n3475), .B(n3277), .Z(n3278) );
  XOR U5252 ( .A(n3633), .B(n3278), .Z(out[452]) );
  XOR U5253 ( .A(in[891]), .B(n3279), .Z(n3637) );
  NANDN U5254 ( .A(n3476), .B(n3280), .Z(n3281) );
  XNOR U5255 ( .A(n3637), .B(n3281), .Z(out[453]) );
  XOR U5256 ( .A(in[892]), .B(n3282), .Z(n3641) );
  NANDN U5257 ( .A(n3477), .B(n3283), .Z(n3284) );
  XNOR U5258 ( .A(n3641), .B(n3284), .Z(out[454]) );
  XOR U5259 ( .A(in[893]), .B(n3285), .Z(n3645) );
  NANDN U5260 ( .A(n3478), .B(n3286), .Z(n3287) );
  XNOR U5261 ( .A(n3645), .B(n3287), .Z(out[455]) );
  XOR U5262 ( .A(in[894]), .B(n3288), .Z(n3649) );
  NANDN U5263 ( .A(n3483), .B(n3289), .Z(n3290) );
  XOR U5264 ( .A(n3649), .B(n3290), .Z(out[456]) );
  IV U5265 ( .A(n3291), .Z(n3900) );
  XOR U5266 ( .A(in[895]), .B(n3900), .Z(n3652) );
  NAND U5267 ( .A(n3292), .B(n3484), .Z(n3293) );
  XNOR U5268 ( .A(n3652), .B(n3293), .Z(out[457]) );
  IV U5269 ( .A(n3294), .Z(n3904) );
  XOR U5270 ( .A(in[832]), .B(n3904), .Z(n3656) );
  NAND U5271 ( .A(n3295), .B(n3486), .Z(n3296) );
  XNOR U5272 ( .A(n3656), .B(n3296), .Z(out[458]) );
  IV U5273 ( .A(n3297), .Z(n3908) );
  XOR U5274 ( .A(in[833]), .B(n3908), .Z(n3660) );
  NAND U5275 ( .A(n3298), .B(n3488), .Z(n3299) );
  XNOR U5276 ( .A(n3660), .B(n3299), .Z(out[459]) );
  AND U5277 ( .A(n3301), .B(n3300), .Z(n3302) );
  XNOR U5278 ( .A(n3303), .B(n3302), .Z(out[45]) );
  IV U5279 ( .A(n3304), .Z(n3912) );
  XOR U5280 ( .A(in[834]), .B(n3912), .Z(n3664) );
  NAND U5281 ( .A(n3305), .B(n3490), .Z(n3306) );
  XNOR U5282 ( .A(n3664), .B(n3306), .Z(out[460]) );
  IV U5283 ( .A(n3307), .Z(n3916) );
  XOR U5284 ( .A(in[835]), .B(n3916), .Z(n3668) );
  NAND U5285 ( .A(n3308), .B(n3492), .Z(n3309) );
  XNOR U5286 ( .A(n3668), .B(n3309), .Z(out[461]) );
  IV U5287 ( .A(n3310), .Z(n3920) );
  XOR U5288 ( .A(in[836]), .B(n3920), .Z(n3676) );
  NAND U5289 ( .A(n3311), .B(n3494), .Z(n3312) );
  XNOR U5290 ( .A(n3676), .B(n3312), .Z(out[462]) );
  IV U5291 ( .A(n3313), .Z(n3924) );
  XOR U5292 ( .A(in[837]), .B(n3924), .Z(n3680) );
  NAND U5293 ( .A(n3314), .B(n3496), .Z(n3315) );
  XNOR U5294 ( .A(n3680), .B(n3315), .Z(out[463]) );
  IV U5295 ( .A(n3316), .Z(n3928) );
  XOR U5296 ( .A(in[838]), .B(n3928), .Z(n3684) );
  NAND U5297 ( .A(n3317), .B(n3498), .Z(n3318) );
  XNOR U5298 ( .A(n3684), .B(n3318), .Z(out[464]) );
  XNOR U5299 ( .A(in[839]), .B(n3319), .Z(n3688) );
  NANDN U5300 ( .A(n3500), .B(n3320), .Z(n3321) );
  XNOR U5301 ( .A(n3688), .B(n3321), .Z(out[465]) );
  XNOR U5302 ( .A(in[840]), .B(n3935), .Z(n3692) );
  NANDN U5303 ( .A(n3505), .B(n3322), .Z(n3323) );
  XNOR U5304 ( .A(n3692), .B(n3323), .Z(out[466]) );
  XNOR U5305 ( .A(in[841]), .B(n3942), .Z(n3696) );
  NANDN U5306 ( .A(n3506), .B(n3324), .Z(n3325) );
  XNOR U5307 ( .A(n3696), .B(n3325), .Z(out[467]) );
  XNOR U5308 ( .A(in[842]), .B(n3946), .Z(n3700) );
  NANDN U5309 ( .A(n3507), .B(n3326), .Z(n3327) );
  XNOR U5310 ( .A(n3700), .B(n3327), .Z(out[468]) );
  XNOR U5311 ( .A(in[843]), .B(n3950), .Z(n3704) );
  NANDN U5312 ( .A(n3508), .B(n3328), .Z(n3329) );
  XNOR U5313 ( .A(n3704), .B(n3329), .Z(out[469]) );
  AND U5314 ( .A(n3331), .B(n3330), .Z(n3332) );
  XNOR U5315 ( .A(n3333), .B(n3332), .Z(out[46]) );
  XNOR U5316 ( .A(in[844]), .B(n3954), .Z(n3708) );
  NANDN U5317 ( .A(n3509), .B(n3334), .Z(n3335) );
  XNOR U5318 ( .A(n3708), .B(n3335), .Z(out[470]) );
  XNOR U5319 ( .A(in[845]), .B(n3958), .Z(n3712) );
  NANDN U5320 ( .A(n3510), .B(n3336), .Z(n3337) );
  XNOR U5321 ( .A(n3712), .B(n3337), .Z(out[471]) );
  XNOR U5322 ( .A(in[846]), .B(n3962), .Z(n3722) );
  NANDN U5323 ( .A(n3511), .B(n3338), .Z(n3339) );
  XNOR U5324 ( .A(n3722), .B(n3339), .Z(out[472]) );
  XNOR U5325 ( .A(in[847]), .B(n3966), .Z(n3726) );
  NANDN U5326 ( .A(n3512), .B(n3340), .Z(n3341) );
  XNOR U5327 ( .A(n3726), .B(n3341), .Z(out[473]) );
  XNOR U5328 ( .A(in[848]), .B(n3970), .Z(n3730) );
  NAND U5329 ( .A(n3342), .B(n3513), .Z(n3343) );
  XNOR U5330 ( .A(n3730), .B(n3343), .Z(out[474]) );
  XNOR U5331 ( .A(in[849]), .B(n3974), .Z(n3734) );
  NANDN U5332 ( .A(n3515), .B(n3344), .Z(n3345) );
  XNOR U5333 ( .A(n3734), .B(n3345), .Z(out[475]) );
  XNOR U5334 ( .A(in[850]), .B(n3978), .Z(n3738) );
  IV U5335 ( .A(n3346), .Z(n3520) );
  NANDN U5336 ( .A(n3347), .B(n3520), .Z(n3348) );
  XNOR U5337 ( .A(n3738), .B(n3348), .Z(out[476]) );
  XOR U5338 ( .A(in[851]), .B(n3349), .Z(n3742) );
  IV U5339 ( .A(n3350), .Z(n3522) );
  NANDN U5340 ( .A(n3351), .B(n3522), .Z(n3352) );
  XOR U5341 ( .A(n3742), .B(n3352), .Z(out[477]) );
  XOR U5342 ( .A(in[852]), .B(n3989), .Z(n3524) );
  IV U5343 ( .A(n3353), .Z(n3525) );
  NANDN U5344 ( .A(n3354), .B(n3525), .Z(n3355) );
  XNOR U5345 ( .A(n3524), .B(n3355), .Z(out[478]) );
  XOR U5346 ( .A(in[853]), .B(n3993), .Z(n3750) );
  IV U5347 ( .A(n3356), .Z(n3527) );
  NANDN U5348 ( .A(n3357), .B(n3527), .Z(n3358) );
  XOR U5349 ( .A(n3750), .B(n3358), .Z(out[479]) );
  ANDN U5350 ( .B(n3360), .A(n3359), .Z(n3361) );
  XNOR U5351 ( .A(n3362), .B(n3361), .Z(out[47]) );
  XOR U5352 ( .A(in[854]), .B(n3997), .Z(n3754) );
  IV U5353 ( .A(n3363), .Z(n3529) );
  NANDN U5354 ( .A(n3364), .B(n3529), .Z(n3365) );
  XOR U5355 ( .A(n3754), .B(n3365), .Z(out[480]) );
  XOR U5356 ( .A(in[855]), .B(n4001), .Z(n3531) );
  IV U5357 ( .A(n3366), .Z(n3532) );
  NANDN U5358 ( .A(n3367), .B(n3532), .Z(n3368) );
  XNOR U5359 ( .A(n3531), .B(n3368), .Z(out[481]) );
  XOR U5360 ( .A(in[856]), .B(n4005), .Z(n3534) );
  IV U5361 ( .A(n3369), .Z(n3535) );
  NANDN U5362 ( .A(n3370), .B(n3535), .Z(n3371) );
  XNOR U5363 ( .A(n3534), .B(n3371), .Z(out[482]) );
  XOR U5364 ( .A(in[857]), .B(n4009), .Z(n3537) );
  IV U5365 ( .A(n3372), .Z(n3538) );
  NANDN U5366 ( .A(n3373), .B(n3538), .Z(n3374) );
  XNOR U5367 ( .A(n3537), .B(n3374), .Z(out[483]) );
  XOR U5368 ( .A(in[858]), .B(n4013), .Z(n3774) );
  NANDN U5369 ( .A(n3375), .B(n3540), .Z(n3376) );
  XOR U5370 ( .A(n3774), .B(n3376), .Z(out[484]) );
  XOR U5371 ( .A(in[859]), .B(n4017), .Z(n3778) );
  NANDN U5372 ( .A(n3377), .B(n3542), .Z(n3378) );
  XOR U5373 ( .A(n3778), .B(n3378), .Z(out[485]) );
  XOR U5374 ( .A(in[860]), .B(n4021), .Z(n3548) );
  NANDN U5375 ( .A(n3379), .B(n3549), .Z(n3380) );
  XNOR U5376 ( .A(n3548), .B(n3380), .Z(out[486]) );
  XOR U5377 ( .A(in[861]), .B(n4029), .Z(n3551) );
  NANDN U5378 ( .A(n3381), .B(n3552), .Z(n3382) );
  XNOR U5379 ( .A(n3551), .B(n3382), .Z(out[487]) );
  XOR U5380 ( .A(in[862]), .B(n4033), .Z(n3554) );
  NANDN U5381 ( .A(n3383), .B(n3555), .Z(n3384) );
  XNOR U5382 ( .A(n3554), .B(n3384), .Z(out[488]) );
  XOR U5383 ( .A(in[863]), .B(n4037), .Z(n3557) );
  NANDN U5384 ( .A(n3385), .B(n3558), .Z(n3386) );
  XNOR U5385 ( .A(n3557), .B(n3386), .Z(out[489]) );
  AND U5386 ( .A(n3388), .B(n3387), .Z(n3389) );
  XNOR U5387 ( .A(n3390), .B(n3389), .Z(out[48]) );
  XOR U5388 ( .A(in[864]), .B(n4041), .Z(n3560) );
  NANDN U5389 ( .A(n3391), .B(n3561), .Z(n3392) );
  XNOR U5390 ( .A(n3560), .B(n3392), .Z(out[490]) );
  XOR U5391 ( .A(in[865]), .B(n4045), .Z(n3563) );
  NANDN U5392 ( .A(n3393), .B(n3564), .Z(n3394) );
  XNOR U5393 ( .A(n3563), .B(n3394), .Z(out[491]) );
  XNOR U5394 ( .A(n3395), .B(in[866]), .Z(n3811) );
  NANDN U5395 ( .A(n3396), .B(n3566), .Z(n3397) );
  XNOR U5396 ( .A(n3811), .B(n3397), .Z(out[492]) );
  XNOR U5397 ( .A(n3398), .B(in[867]), .Z(n3815) );
  IV U5398 ( .A(n3399), .Z(n3568) );
  NANDN U5399 ( .A(n3400), .B(n3568), .Z(n3401) );
  XNOR U5400 ( .A(n3815), .B(n3401), .Z(out[493]) );
  XNOR U5401 ( .A(n3402), .B(in[868]), .Z(n3819) );
  IV U5402 ( .A(n3403), .Z(n3570) );
  NANDN U5403 ( .A(n3404), .B(n3570), .Z(n3405) );
  XNOR U5404 ( .A(n3819), .B(n3405), .Z(out[494]) );
  XNOR U5405 ( .A(n3406), .B(in[869]), .Z(n3823) );
  IV U5406 ( .A(n3407), .Z(n3572) );
  NANDN U5407 ( .A(n3408), .B(n3572), .Z(n3409) );
  XNOR U5408 ( .A(n3823), .B(n3409), .Z(out[495]) );
  XOR U5409 ( .A(in[870]), .B(n4065), .Z(n3827) );
  IV U5410 ( .A(n3410), .Z(n3578) );
  NANDN U5411 ( .A(n3411), .B(n3578), .Z(n3412) );
  XOR U5412 ( .A(n3827), .B(n3412), .Z(out[496]) );
  XOR U5413 ( .A(in[871]), .B(n4073), .Z(n3831) );
  IV U5414 ( .A(n3413), .Z(n3580) );
  NANDN U5415 ( .A(n3414), .B(n3580), .Z(n3415) );
  XOR U5416 ( .A(n3831), .B(n3415), .Z(out[497]) );
  XOR U5417 ( .A(in[872]), .B(n4077), .Z(n3835) );
  IV U5418 ( .A(n3416), .Z(n3582) );
  NANDN U5419 ( .A(n3417), .B(n3582), .Z(n3418) );
  XOR U5420 ( .A(n3835), .B(n3418), .Z(out[498]) );
  XOR U5421 ( .A(in[873]), .B(n4081), .Z(n3839) );
  IV U5422 ( .A(n3419), .Z(n3584) );
  NANDN U5423 ( .A(n3420), .B(n3584), .Z(n3421) );
  XOR U5424 ( .A(n3839), .B(n3421), .Z(out[499]) );
  ANDN U5425 ( .B(n3423), .A(n3422), .Z(n3424) );
  XNOR U5426 ( .A(n3425), .B(n3424), .Z(out[49]) );
  OR U5427 ( .A(n4113), .B(n3426), .Z(n3427) );
  XNOR U5428 ( .A(n4112), .B(n3427), .Z(out[4]) );
  XOR U5429 ( .A(in[874]), .B(n4085), .Z(n3843) );
  NAND U5430 ( .A(n3428), .B(n3586), .Z(n3429) );
  XOR U5431 ( .A(n3843), .B(n3429), .Z(out[500]) );
  XOR U5432 ( .A(in[875]), .B(n3430), .Z(n3847) );
  NAND U5433 ( .A(n3431), .B(n3588), .Z(n3432) );
  XOR U5434 ( .A(n3847), .B(n3432), .Z(out[501]) );
  XOR U5435 ( .A(in[876]), .B(n3433), .Z(n3855) );
  NAND U5436 ( .A(n3434), .B(n3590), .Z(n3435) );
  XOR U5437 ( .A(n3855), .B(n3435), .Z(out[502]) );
  XOR U5438 ( .A(in[877]), .B(n3436), .Z(n3859) );
  NAND U5439 ( .A(n3437), .B(n3592), .Z(n3438) );
  XOR U5440 ( .A(n3859), .B(n3438), .Z(out[503]) );
  XOR U5441 ( .A(in[878]), .B(n3439), .Z(n3863) );
  NAND U5442 ( .A(n3440), .B(n3594), .Z(n3441) );
  XOR U5443 ( .A(n3863), .B(n3441), .Z(out[504]) );
  XOR U5444 ( .A(in[879]), .B(n3442), .Z(n3867) );
  NAND U5445 ( .A(n3443), .B(n3596), .Z(n3444) );
  XOR U5446 ( .A(n3867), .B(n3444), .Z(out[505]) );
  XOR U5447 ( .A(in[880]), .B(n3445), .Z(n3871) );
  NANDN U5448 ( .A(n3602), .B(n3446), .Z(n3447) );
  XOR U5449 ( .A(n3871), .B(n3447), .Z(out[506]) );
  XOR U5450 ( .A(in[881]), .B(n3448), .Z(n3875) );
  NANDN U5451 ( .A(n3603), .B(n3449), .Z(n3450) );
  XOR U5452 ( .A(n3875), .B(n3450), .Z(out[507]) );
  XOR U5453 ( .A(in[882]), .B(n3451), .Z(n3879) );
  NAND U5454 ( .A(n3452), .B(n3604), .Z(n3453) );
  XOR U5455 ( .A(n3879), .B(n3453), .Z(out[508]) );
  XOR U5456 ( .A(in[883]), .B(n3454), .Z(n3883) );
  NAND U5457 ( .A(n3455), .B(n3606), .Z(n3456) );
  XOR U5458 ( .A(n3883), .B(n3456), .Z(out[509]) );
  ANDN U5459 ( .B(n3458), .A(n3457), .Z(n3459) );
  XNOR U5460 ( .A(n3460), .B(n3459), .Z(out[50]) );
  XOR U5461 ( .A(in[884]), .B(n3461), .Z(n3887) );
  NANDN U5462 ( .A(n3462), .B(n3608), .Z(n3463) );
  XOR U5463 ( .A(n3887), .B(n3463), .Z(out[510]) );
  XOR U5464 ( .A(in[885]), .B(n3464), .Z(n3891) );
  NAND U5465 ( .A(n3465), .B(n3610), .Z(n3466) );
  XOR U5466 ( .A(n3891), .B(n3466), .Z(out[511]) );
  NANDN U5467 ( .A(n3467), .B(n3613), .Z(n3468) );
  XNOR U5468 ( .A(n3612), .B(n3468), .Z(out[512]) );
  NANDN U5469 ( .A(n3469), .B(n3617), .Z(n3470) );
  XNOR U5470 ( .A(n3616), .B(n3470), .Z(out[513]) );
  NANDN U5471 ( .A(n3471), .B(n3621), .Z(n3472) );
  XNOR U5472 ( .A(n3620), .B(n3472), .Z(out[514]) );
  NANDN U5473 ( .A(n3473), .B(n3625), .Z(n3474) );
  XNOR U5474 ( .A(n3624), .B(n3474), .Z(out[515]) );
  ANDN U5475 ( .B(n3480), .A(n3479), .Z(n3481) );
  XNOR U5476 ( .A(n3482), .B(n3481), .Z(out[51]) );
  OR U5477 ( .A(n3652), .B(n3484), .Z(n3485) );
  XOR U5478 ( .A(n3653), .B(n3485), .Z(out[521]) );
  OR U5479 ( .A(n3656), .B(n3486), .Z(n3487) );
  XOR U5480 ( .A(n3657), .B(n3487), .Z(out[522]) );
  OR U5481 ( .A(n3660), .B(n3488), .Z(n3489) );
  XOR U5482 ( .A(n3661), .B(n3489), .Z(out[523]) );
  OR U5483 ( .A(n3664), .B(n3490), .Z(n3491) );
  XOR U5484 ( .A(n3665), .B(n3491), .Z(out[524]) );
  OR U5485 ( .A(n3668), .B(n3492), .Z(n3493) );
  XOR U5486 ( .A(n3669), .B(n3493), .Z(out[525]) );
  OR U5487 ( .A(n3676), .B(n3494), .Z(n3495) );
  XOR U5488 ( .A(n3677), .B(n3495), .Z(out[526]) );
  OR U5489 ( .A(n3680), .B(n3496), .Z(n3497) );
  XOR U5490 ( .A(n3681), .B(n3497), .Z(out[527]) );
  OR U5491 ( .A(n3684), .B(n3498), .Z(n3499) );
  XOR U5492 ( .A(n3685), .B(n3499), .Z(out[528]) );
  ANDN U5493 ( .B(n3502), .A(n3501), .Z(n3503) );
  XNOR U5494 ( .A(n3504), .B(n3503), .Z(out[52]) );
  OR U5495 ( .A(n3730), .B(n3513), .Z(n3514) );
  XOR U5496 ( .A(n3731), .B(n3514), .Z(out[538]) );
  ANDN U5497 ( .B(n3517), .A(n3516), .Z(n3518) );
  XNOR U5498 ( .A(n3519), .B(n3518), .Z(out[53]) );
  OR U5499 ( .A(n3738), .B(n3520), .Z(n3521) );
  XOR U5500 ( .A(n3739), .B(n3521), .Z(out[540]) );
  NANDN U5501 ( .A(n3522), .B(n3742), .Z(n3523) );
  XOR U5502 ( .A(n3743), .B(n3523), .Z(out[541]) );
  IV U5503 ( .A(n3524), .Z(n3746) );
  NANDN U5504 ( .A(n3525), .B(n3746), .Z(n3526) );
  XOR U5505 ( .A(n3747), .B(n3526), .Z(out[542]) );
  NANDN U5506 ( .A(n3527), .B(n3750), .Z(n3528) );
  XOR U5507 ( .A(n3751), .B(n3528), .Z(out[543]) );
  NANDN U5508 ( .A(n3529), .B(n3754), .Z(n3530) );
  XOR U5509 ( .A(n3755), .B(n3530), .Z(out[544]) );
  IV U5510 ( .A(n3531), .Z(n3758) );
  NANDN U5511 ( .A(n3532), .B(n3758), .Z(n3533) );
  XOR U5512 ( .A(n3759), .B(n3533), .Z(out[545]) );
  IV U5513 ( .A(n3534), .Z(n3766) );
  NANDN U5514 ( .A(n3535), .B(n3766), .Z(n3536) );
  XOR U5515 ( .A(n3767), .B(n3536), .Z(out[546]) );
  IV U5516 ( .A(n3537), .Z(n3770) );
  NANDN U5517 ( .A(n3538), .B(n3770), .Z(n3539) );
  XOR U5518 ( .A(n3771), .B(n3539), .Z(out[547]) );
  NANDN U5519 ( .A(n3540), .B(n3774), .Z(n3541) );
  XOR U5520 ( .A(n3775), .B(n3541), .Z(out[548]) );
  NANDN U5521 ( .A(n3542), .B(n3778), .Z(n3543) );
  XOR U5522 ( .A(n3779), .B(n3543), .Z(out[549]) );
  ANDN U5523 ( .B(n3545), .A(n3544), .Z(n3546) );
  XNOR U5524 ( .A(n3547), .B(n3546), .Z(out[54]) );
  IV U5525 ( .A(n3548), .Z(n3782) );
  NANDN U5526 ( .A(n3549), .B(n3782), .Z(n3550) );
  XOR U5527 ( .A(n3783), .B(n3550), .Z(out[550]) );
  IV U5528 ( .A(n3551), .Z(n3786) );
  NANDN U5529 ( .A(n3552), .B(n3786), .Z(n3553) );
  XOR U5530 ( .A(n3787), .B(n3553), .Z(out[551]) );
  IV U5531 ( .A(n3554), .Z(n3791) );
  NANDN U5532 ( .A(n3555), .B(n3791), .Z(n3556) );
  XNOR U5533 ( .A(n3790), .B(n3556), .Z(out[552]) );
  IV U5534 ( .A(n3557), .Z(n3795) );
  NANDN U5535 ( .A(n3558), .B(n3795), .Z(n3559) );
  XNOR U5536 ( .A(n3794), .B(n3559), .Z(out[553]) );
  IV U5537 ( .A(n3560), .Z(n3799) );
  NANDN U5538 ( .A(n3561), .B(n3799), .Z(n3562) );
  XNOR U5539 ( .A(n3798), .B(n3562), .Z(out[554]) );
  IV U5540 ( .A(n3563), .Z(n3803) );
  NANDN U5541 ( .A(n3564), .B(n3803), .Z(n3565) );
  XNOR U5542 ( .A(n3802), .B(n3565), .Z(out[555]) );
  OR U5543 ( .A(n3811), .B(n3566), .Z(n3567) );
  XNOR U5544 ( .A(n3810), .B(n3567), .Z(out[556]) );
  OR U5545 ( .A(n3815), .B(n3568), .Z(n3569) );
  XNOR U5546 ( .A(n3814), .B(n3569), .Z(out[557]) );
  OR U5547 ( .A(n3819), .B(n3570), .Z(n3571) );
  XNOR U5548 ( .A(n3818), .B(n3571), .Z(out[558]) );
  OR U5549 ( .A(n3823), .B(n3572), .Z(n3573) );
  XNOR U5550 ( .A(n3822), .B(n3573), .Z(out[559]) );
  ANDN U5551 ( .B(n3575), .A(n3574), .Z(n3576) );
  XNOR U5552 ( .A(n3577), .B(n3576), .Z(out[55]) );
  NANDN U5553 ( .A(n3578), .B(n3827), .Z(n3579) );
  XNOR U5554 ( .A(n3826), .B(n3579), .Z(out[560]) );
  NANDN U5555 ( .A(n3580), .B(n3831), .Z(n3581) );
  XNOR U5556 ( .A(n3830), .B(n3581), .Z(out[561]) );
  NANDN U5557 ( .A(n3582), .B(n3835), .Z(n3583) );
  XNOR U5558 ( .A(n3834), .B(n3583), .Z(out[562]) );
  NANDN U5559 ( .A(n3584), .B(n3839), .Z(n3585) );
  XNOR U5560 ( .A(n3838), .B(n3585), .Z(out[563]) );
  NANDN U5561 ( .A(n3586), .B(n3843), .Z(n3587) );
  XNOR U5562 ( .A(n3842), .B(n3587), .Z(out[564]) );
  NANDN U5563 ( .A(n3588), .B(n3847), .Z(n3589) );
  XNOR U5564 ( .A(n3846), .B(n3589), .Z(out[565]) );
  NANDN U5565 ( .A(n3590), .B(n3855), .Z(n3591) );
  XNOR U5566 ( .A(n3854), .B(n3591), .Z(out[566]) );
  NANDN U5567 ( .A(n3592), .B(n3859), .Z(n3593) );
  XNOR U5568 ( .A(n3858), .B(n3593), .Z(out[567]) );
  NANDN U5569 ( .A(n3594), .B(n3863), .Z(n3595) );
  XNOR U5570 ( .A(n3862), .B(n3595), .Z(out[568]) );
  NANDN U5571 ( .A(n3596), .B(n3867), .Z(n3597) );
  XNOR U5572 ( .A(n3866), .B(n3597), .Z(out[569]) );
  ANDN U5573 ( .B(n3599), .A(n3598), .Z(n3600) );
  XNOR U5574 ( .A(n3601), .B(n3600), .Z(out[56]) );
  NANDN U5575 ( .A(n3604), .B(n3879), .Z(n3605) );
  XNOR U5576 ( .A(n3878), .B(n3605), .Z(out[572]) );
  NANDN U5577 ( .A(n3606), .B(n3883), .Z(n3607) );
  XNOR U5578 ( .A(n3882), .B(n3607), .Z(out[573]) );
  NANDN U5579 ( .A(n3608), .B(n3887), .Z(n3609) );
  XNOR U5580 ( .A(n3886), .B(n3609), .Z(out[574]) );
  NANDN U5581 ( .A(n3610), .B(n3891), .Z(n3611) );
  XNOR U5582 ( .A(n3890), .B(n3611), .Z(out[575]) );
  NOR U5583 ( .A(n3613), .B(n3612), .Z(n3614) );
  XOR U5584 ( .A(n3615), .B(n3614), .Z(out[576]) );
  NOR U5585 ( .A(n3617), .B(n3616), .Z(n3618) );
  XOR U5586 ( .A(n3619), .B(n3618), .Z(out[577]) );
  NOR U5587 ( .A(n3621), .B(n3620), .Z(n3622) );
  XOR U5588 ( .A(n3623), .B(n3622), .Z(out[578]) );
  NOR U5589 ( .A(n3625), .B(n3624), .Z(n3626) );
  XOR U5590 ( .A(n3627), .B(n3626), .Z(out[579]) );
  ANDN U5591 ( .B(n3629), .A(n3628), .Z(n3630) );
  XNOR U5592 ( .A(n3631), .B(n3630), .Z(out[57]) );
  NOR U5593 ( .A(n3633), .B(n3632), .Z(n3634) );
  XOR U5594 ( .A(n3635), .B(n3634), .Z(out[580]) );
  ANDN U5595 ( .B(n3637), .A(n3636), .Z(n3638) );
  XOR U5596 ( .A(n3639), .B(n3638), .Z(out[581]) );
  ANDN U5597 ( .B(n3641), .A(n3640), .Z(n3642) );
  XOR U5598 ( .A(n3643), .B(n3642), .Z(out[582]) );
  ANDN U5599 ( .B(n3645), .A(n3644), .Z(n3646) );
  XOR U5600 ( .A(n3647), .B(n3646), .Z(out[583]) );
  NOR U5601 ( .A(n3649), .B(n3648), .Z(n3650) );
  XOR U5602 ( .A(n3651), .B(n3650), .Z(out[584]) );
  AND U5603 ( .A(n3653), .B(n3652), .Z(n3654) );
  XNOR U5604 ( .A(n3655), .B(n3654), .Z(out[585]) );
  AND U5605 ( .A(n3657), .B(n3656), .Z(n3658) );
  XNOR U5606 ( .A(n3659), .B(n3658), .Z(out[586]) );
  AND U5607 ( .A(n3661), .B(n3660), .Z(n3662) );
  XNOR U5608 ( .A(n3663), .B(n3662), .Z(out[587]) );
  AND U5609 ( .A(n3665), .B(n3664), .Z(n3666) );
  XNOR U5610 ( .A(n3667), .B(n3666), .Z(out[588]) );
  AND U5611 ( .A(n3669), .B(n3668), .Z(n3670) );
  XNOR U5612 ( .A(n3671), .B(n3670), .Z(out[589]) );
  ANDN U5613 ( .B(n3673), .A(n3672), .Z(n3674) );
  XNOR U5614 ( .A(n3675), .B(n3674), .Z(out[58]) );
  AND U5615 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U5616 ( .A(n3679), .B(n3678), .Z(out[590]) );
  AND U5617 ( .A(n3681), .B(n3680), .Z(n3682) );
  XNOR U5618 ( .A(n3683), .B(n3682), .Z(out[591]) );
  AND U5619 ( .A(n3685), .B(n3684), .Z(n3686) );
  XNOR U5620 ( .A(n3687), .B(n3686), .Z(out[592]) );
  AND U5621 ( .A(n3689), .B(n3688), .Z(n3690) );
  XNOR U5622 ( .A(n3691), .B(n3690), .Z(out[593]) );
  AND U5623 ( .A(n3693), .B(n3692), .Z(n3694) );
  XNOR U5624 ( .A(n3695), .B(n3694), .Z(out[594]) );
  AND U5625 ( .A(n3697), .B(n3696), .Z(n3698) );
  XNOR U5626 ( .A(n3699), .B(n3698), .Z(out[595]) );
  AND U5627 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR U5628 ( .A(n3703), .B(n3702), .Z(out[596]) );
  AND U5629 ( .A(n3705), .B(n3704), .Z(n3706) );
  XNOR U5630 ( .A(n3707), .B(n3706), .Z(out[597]) );
  AND U5631 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U5632 ( .A(n3711), .B(n3710), .Z(out[598]) );
  AND U5633 ( .A(n3713), .B(n3712), .Z(n3714) );
  XNOR U5634 ( .A(n3715), .B(n3714), .Z(out[599]) );
  ANDN U5635 ( .B(n3717), .A(n3716), .Z(n3718) );
  XNOR U5636 ( .A(n3719), .B(n3718), .Z(out[59]) );
  OR U5637 ( .A(n4157), .B(n3720), .Z(n3721) );
  XNOR U5638 ( .A(n4156), .B(n3721), .Z(out[5]) );
  AND U5639 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U5640 ( .A(n3725), .B(n3724), .Z(out[600]) );
  AND U5641 ( .A(n3727), .B(n3726), .Z(n3728) );
  XNOR U5642 ( .A(n3729), .B(n3728), .Z(out[601]) );
  AND U5643 ( .A(n3731), .B(n3730), .Z(n3732) );
  XNOR U5644 ( .A(n3733), .B(n3732), .Z(out[602]) );
  AND U5645 ( .A(n3735), .B(n3734), .Z(n3736) );
  XNOR U5646 ( .A(n3737), .B(n3736), .Z(out[603]) );
  AND U5647 ( .A(n3739), .B(n3738), .Z(n3740) );
  XNOR U5648 ( .A(n3741), .B(n3740), .Z(out[604]) );
  ANDN U5649 ( .B(n3743), .A(n3742), .Z(n3744) );
  XNOR U5650 ( .A(n3745), .B(n3744), .Z(out[605]) );
  ANDN U5651 ( .B(n3747), .A(n3746), .Z(n3748) );
  XNOR U5652 ( .A(n3749), .B(n3748), .Z(out[606]) );
  ANDN U5653 ( .B(n3751), .A(n3750), .Z(n3752) );
  XNOR U5654 ( .A(n3753), .B(n3752), .Z(out[607]) );
  ANDN U5655 ( .B(n3755), .A(n3754), .Z(n3756) );
  XNOR U5656 ( .A(n3757), .B(n3756), .Z(out[608]) );
  ANDN U5657 ( .B(n3759), .A(n3758), .Z(n3760) );
  XNOR U5658 ( .A(n3761), .B(n3760), .Z(out[609]) );
  ANDN U5659 ( .B(n3763), .A(n3762), .Z(n3764) );
  XNOR U5660 ( .A(n3765), .B(n3764), .Z(out[60]) );
  ANDN U5661 ( .B(n3767), .A(n3766), .Z(n3768) );
  XNOR U5662 ( .A(n3769), .B(n3768), .Z(out[610]) );
  ANDN U5663 ( .B(n3771), .A(n3770), .Z(n3772) );
  XNOR U5664 ( .A(n3773), .B(n3772), .Z(out[611]) );
  ANDN U5665 ( .B(n3775), .A(n3774), .Z(n3776) );
  XNOR U5666 ( .A(n3777), .B(n3776), .Z(out[612]) );
  ANDN U5667 ( .B(n3779), .A(n3778), .Z(n3780) );
  XNOR U5668 ( .A(n3781), .B(n3780), .Z(out[613]) );
  ANDN U5669 ( .B(n3783), .A(n3782), .Z(n3784) );
  XNOR U5670 ( .A(n3785), .B(n3784), .Z(out[614]) );
  ANDN U5671 ( .B(n3787), .A(n3786), .Z(n3788) );
  XNOR U5672 ( .A(n3789), .B(n3788), .Z(out[615]) );
  NOR U5673 ( .A(n3791), .B(n3790), .Z(n3792) );
  XOR U5674 ( .A(n3793), .B(n3792), .Z(out[616]) );
  NOR U5675 ( .A(n3795), .B(n3794), .Z(n3796) );
  XOR U5676 ( .A(n3797), .B(n3796), .Z(out[617]) );
  NOR U5677 ( .A(n3799), .B(n3798), .Z(n3800) );
  XOR U5678 ( .A(n3801), .B(n3800), .Z(out[618]) );
  NOR U5679 ( .A(n3803), .B(n3802), .Z(n3804) );
  XOR U5680 ( .A(n3805), .B(n3804), .Z(out[619]) );
  ANDN U5681 ( .B(n3807), .A(n3806), .Z(n3808) );
  XOR U5682 ( .A(n3809), .B(n3808), .Z(out[61]) );
  ANDN U5683 ( .B(n3811), .A(n3810), .Z(n3812) );
  XOR U5684 ( .A(n3813), .B(n3812), .Z(out[620]) );
  ANDN U5685 ( .B(n3815), .A(n3814), .Z(n3816) );
  XOR U5686 ( .A(n3817), .B(n3816), .Z(out[621]) );
  ANDN U5687 ( .B(n3819), .A(n3818), .Z(n3820) );
  XOR U5688 ( .A(n3821), .B(n3820), .Z(out[622]) );
  ANDN U5689 ( .B(n3823), .A(n3822), .Z(n3824) );
  XOR U5690 ( .A(n3825), .B(n3824), .Z(out[623]) );
  NOR U5691 ( .A(n3827), .B(n3826), .Z(n3828) );
  XOR U5692 ( .A(n3829), .B(n3828), .Z(out[624]) );
  NOR U5693 ( .A(n3831), .B(n3830), .Z(n3832) );
  XOR U5694 ( .A(n3833), .B(n3832), .Z(out[625]) );
  NOR U5695 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U5696 ( .A(n3837), .B(n3836), .Z(out[626]) );
  NOR U5697 ( .A(n3839), .B(n3838), .Z(n3840) );
  XOR U5698 ( .A(n3841), .B(n3840), .Z(out[627]) );
  NOR U5699 ( .A(n3843), .B(n3842), .Z(n3844) );
  XOR U5700 ( .A(n3845), .B(n3844), .Z(out[628]) );
  NOR U5701 ( .A(n3847), .B(n3846), .Z(n3848) );
  XOR U5702 ( .A(n3849), .B(n3848), .Z(out[629]) );
  ANDN U5703 ( .B(n3851), .A(n3850), .Z(n3852) );
  XOR U5704 ( .A(n3853), .B(n3852), .Z(out[62]) );
  NOR U5705 ( .A(n3855), .B(n3854), .Z(n3856) );
  XOR U5706 ( .A(n3857), .B(n3856), .Z(out[630]) );
  NOR U5707 ( .A(n3859), .B(n3858), .Z(n3860) );
  XOR U5708 ( .A(n3861), .B(n3860), .Z(out[631]) );
  NOR U5709 ( .A(n3863), .B(n3862), .Z(n3864) );
  XOR U5710 ( .A(n3865), .B(n3864), .Z(out[632]) );
  NOR U5711 ( .A(n3867), .B(n3866), .Z(n3868) );
  XOR U5712 ( .A(n3869), .B(n3868), .Z(out[633]) );
  NOR U5713 ( .A(n3871), .B(n3870), .Z(n3872) );
  XOR U5714 ( .A(n3873), .B(n3872), .Z(out[634]) );
  NOR U5715 ( .A(n3875), .B(n3874), .Z(n3876) );
  XOR U5716 ( .A(n3877), .B(n3876), .Z(out[635]) );
  NOR U5717 ( .A(n3879), .B(n3878), .Z(n3880) );
  XOR U5718 ( .A(n3881), .B(n3880), .Z(out[636]) );
  NOR U5719 ( .A(n3883), .B(n3882), .Z(n3884) );
  XOR U5720 ( .A(n3885), .B(n3884), .Z(out[637]) );
  NOR U5721 ( .A(n3887), .B(n3886), .Z(n3888) );
  XOR U5722 ( .A(n3889), .B(n3888), .Z(out[638]) );
  NOR U5723 ( .A(n3891), .B(n3890), .Z(n3892) );
  XOR U5724 ( .A(n3893), .B(n3892), .Z(out[639]) );
  ANDN U5725 ( .B(n3895), .A(n3894), .Z(n3896) );
  XOR U5726 ( .A(n3897), .B(n3896), .Z(out[63]) );
  XOR U5727 ( .A(in[302]), .B(n3898), .Z(n4179) );
  IV U5728 ( .A(n4179), .Z(n4336) );
  XOR U5729 ( .A(in[1146]), .B(n3899), .Z(n4709) );
  XOR U5730 ( .A(in[1535]), .B(n3900), .Z(n4711) );
  OR U5731 ( .A(n4709), .B(n4711), .Z(n3901) );
  XOR U5732 ( .A(n4336), .B(n3901), .Z(out[640]) );
  XOR U5733 ( .A(in[303]), .B(n3902), .Z(n4182) );
  IV U5734 ( .A(n4182), .Z(n4338) );
  XOR U5735 ( .A(in[1147]), .B(n3903), .Z(n4713) );
  XOR U5736 ( .A(in[1472]), .B(n3904), .Z(n4715) );
  OR U5737 ( .A(n4713), .B(n4715), .Z(n3905) );
  XOR U5738 ( .A(n4338), .B(n3905), .Z(out[641]) );
  XOR U5739 ( .A(in[304]), .B(n3906), .Z(n4185) );
  IV U5740 ( .A(n4185), .Z(n4344) );
  XOR U5741 ( .A(in[1148]), .B(n3907), .Z(n4717) );
  XOR U5742 ( .A(in[1473]), .B(n3908), .Z(n4719) );
  OR U5743 ( .A(n4717), .B(n4719), .Z(n3909) );
  XOR U5744 ( .A(n4344), .B(n3909), .Z(out[642]) );
  XOR U5745 ( .A(in[305]), .B(n3910), .Z(n4188) );
  IV U5746 ( .A(n4188), .Z(n4346) );
  XOR U5747 ( .A(in[1149]), .B(n3911), .Z(n4721) );
  XOR U5748 ( .A(in[1474]), .B(n3912), .Z(n4723) );
  OR U5749 ( .A(n4721), .B(n4723), .Z(n3913) );
  XOR U5750 ( .A(n4346), .B(n3913), .Z(out[643]) );
  XOR U5751 ( .A(in[306]), .B(n3914), .Z(n4191) );
  IV U5752 ( .A(n4191), .Z(n4348) );
  XOR U5753 ( .A(in[1150]), .B(n3915), .Z(n4733) );
  XOR U5754 ( .A(in[1475]), .B(n3916), .Z(n4735) );
  OR U5755 ( .A(n4733), .B(n4735), .Z(n3917) );
  XOR U5756 ( .A(n4348), .B(n3917), .Z(out[644]) );
  XOR U5757 ( .A(in[307]), .B(n3918), .Z(n4351) );
  XOR U5758 ( .A(in[1151]), .B(n3919), .Z(n4737) );
  XOR U5759 ( .A(in[1476]), .B(n3920), .Z(n4739) );
  OR U5760 ( .A(n4737), .B(n4739), .Z(n3921) );
  XOR U5761 ( .A(n4351), .B(n3921), .Z(out[645]) );
  XOR U5762 ( .A(in[308]), .B(n3922), .Z(n4354) );
  XOR U5763 ( .A(in[1088]), .B(n3923), .Z(n4741) );
  XOR U5764 ( .A(in[1477]), .B(n3924), .Z(n4743) );
  OR U5765 ( .A(n4741), .B(n4743), .Z(n3925) );
  XOR U5766 ( .A(n4354), .B(n3925), .Z(out[646]) );
  XOR U5767 ( .A(in[309]), .B(n3926), .Z(n4357) );
  XOR U5768 ( .A(in[1089]), .B(n3927), .Z(n4745) );
  XOR U5769 ( .A(in[1478]), .B(n3928), .Z(n4747) );
  OR U5770 ( .A(n4745), .B(n4747), .Z(n3929) );
  XOR U5771 ( .A(n4357), .B(n3929), .Z(out[647]) );
  XOR U5772 ( .A(in[310]), .B(n3930), .Z(n4359) );
  XOR U5773 ( .A(in[1479]), .B(n3931), .Z(n4751) );
  XNOR U5774 ( .A(n3932), .B(in[1090]), .Z(n4748) );
  NANDN U5775 ( .A(n4751), .B(n4748), .Z(n3933) );
  XOR U5776 ( .A(n4359), .B(n3933), .Z(out[648]) );
  XOR U5777 ( .A(in[311]), .B(n3934), .Z(n4362) );
  XNOR U5778 ( .A(n3936), .B(in[1091]), .Z(n4752) );
  NANDN U5779 ( .A(n4755), .B(n4752), .Z(n3937) );
  XOR U5780 ( .A(n4362), .B(n3937), .Z(out[649]) );
  XOR U5781 ( .A(in[312]), .B(n3941), .Z(n4365) );
  XNOR U5782 ( .A(n3943), .B(in[1092]), .Z(n4756) );
  NANDN U5783 ( .A(n4759), .B(n4756), .Z(n3944) );
  XOR U5784 ( .A(n4365), .B(n3944), .Z(out[650]) );
  XOR U5785 ( .A(in[313]), .B(n3945), .Z(n4368) );
  XNOR U5786 ( .A(n3947), .B(in[1093]), .Z(n4760) );
  NANDN U5787 ( .A(n4763), .B(n4760), .Z(n3948) );
  XOR U5788 ( .A(n4368), .B(n3948), .Z(out[651]) );
  XOR U5789 ( .A(in[314]), .B(n3949), .Z(n4375) );
  XNOR U5790 ( .A(n3951), .B(in[1094]), .Z(n4764) );
  NANDN U5791 ( .A(n4767), .B(n4764), .Z(n3952) );
  XOR U5792 ( .A(n4375), .B(n3952), .Z(out[652]) );
  XOR U5793 ( .A(in[315]), .B(n3953), .Z(n4206) );
  IV U5794 ( .A(n4206), .Z(n4378) );
  XNOR U5795 ( .A(n3955), .B(in[1095]), .Z(n4768) );
  NANDN U5796 ( .A(n4771), .B(n4768), .Z(n3956) );
  XOR U5797 ( .A(n4378), .B(n3956), .Z(out[653]) );
  XOR U5798 ( .A(in[316]), .B(n3957), .Z(n4209) );
  IV U5799 ( .A(n4209), .Z(n4381) );
  XNOR U5800 ( .A(n3959), .B(in[1096]), .Z(n4776) );
  NANDN U5801 ( .A(n4779), .B(n4776), .Z(n3960) );
  XOR U5802 ( .A(n4381), .B(n3960), .Z(out[654]) );
  XOR U5803 ( .A(in[317]), .B(n3961), .Z(n4212) );
  IV U5804 ( .A(n4212), .Z(n4384) );
  XNOR U5805 ( .A(in[1097]), .B(n3963), .Z(n4780) );
  NANDN U5806 ( .A(n4783), .B(n4780), .Z(n3964) );
  XOR U5807 ( .A(n4384), .B(n3964), .Z(out[655]) );
  XOR U5808 ( .A(in[318]), .B(n3965), .Z(n4217) );
  IV U5809 ( .A(n4217), .Z(n4387) );
  XNOR U5810 ( .A(n3967), .B(in[1098]), .Z(n4784) );
  NANDN U5811 ( .A(n4787), .B(n4784), .Z(n3968) );
  XOR U5812 ( .A(n4387), .B(n3968), .Z(out[656]) );
  XOR U5813 ( .A(in[319]), .B(n3969), .Z(n4220) );
  IV U5814 ( .A(n4220), .Z(n4389) );
  XNOR U5815 ( .A(n3971), .B(in[1099]), .Z(n4788) );
  NANDN U5816 ( .A(n4791), .B(n4788), .Z(n3972) );
  XOR U5817 ( .A(n4389), .B(n3972), .Z(out[657]) );
  XOR U5818 ( .A(in[256]), .B(n3973), .Z(n4223) );
  IV U5819 ( .A(n4223), .Z(n4392) );
  XNOR U5820 ( .A(in[1100]), .B(n3975), .Z(n4792) );
  NANDN U5821 ( .A(n4795), .B(n4792), .Z(n3976) );
  XOR U5822 ( .A(n4392), .B(n3976), .Z(out[658]) );
  XOR U5823 ( .A(in[257]), .B(n3977), .Z(n4226) );
  IV U5824 ( .A(n4226), .Z(n4395) );
  XNOR U5825 ( .A(in[1101]), .B(n3979), .Z(n4796) );
  NANDN U5826 ( .A(n4799), .B(n4796), .Z(n3980) );
  XOR U5827 ( .A(n4395), .B(n3980), .Z(out[659]) );
  XOR U5828 ( .A(in[258]), .B(n3984), .Z(n4229) );
  IV U5829 ( .A(n4229), .Z(n4398) );
  XOR U5830 ( .A(in[1491]), .B(n3985), .Z(n4803) );
  XNOR U5831 ( .A(in[1102]), .B(n3986), .Z(n4800) );
  NANDN U5832 ( .A(n4803), .B(n4800), .Z(n3987) );
  XOR U5833 ( .A(n4398), .B(n3987), .Z(out[660]) );
  XOR U5834 ( .A(in[259]), .B(n3988), .Z(n4232) );
  IV U5835 ( .A(n4232), .Z(n4401) );
  XOR U5836 ( .A(in[1492]), .B(n3989), .Z(n4807) );
  XNOR U5837 ( .A(in[1103]), .B(n3990), .Z(n4804) );
  NANDN U5838 ( .A(n4807), .B(n4804), .Z(n3991) );
  XOR U5839 ( .A(n4401), .B(n3991), .Z(out[661]) );
  XOR U5840 ( .A(in[260]), .B(n3992), .Z(n4408) );
  XOR U5841 ( .A(in[1493]), .B(n3993), .Z(n4235) );
  IV U5842 ( .A(n4235), .Z(n4811) );
  XNOR U5843 ( .A(in[1104]), .B(n3994), .Z(n4808) );
  NANDN U5844 ( .A(n4811), .B(n4808), .Z(n3995) );
  XNOR U5845 ( .A(n4408), .B(n3995), .Z(out[662]) );
  XOR U5846 ( .A(in[261]), .B(n3996), .Z(n4411) );
  XOR U5847 ( .A(in[1494]), .B(n3997), .Z(n4238) );
  IV U5848 ( .A(n4238), .Z(n4815) );
  XNOR U5849 ( .A(in[1105]), .B(n3998), .Z(n4812) );
  NANDN U5850 ( .A(n4815), .B(n4812), .Z(n3999) );
  XNOR U5851 ( .A(n4411), .B(n3999), .Z(out[663]) );
  XOR U5852 ( .A(in[262]), .B(n4000), .Z(n4414) );
  XOR U5853 ( .A(in[1495]), .B(n4001), .Z(n4823) );
  XNOR U5854 ( .A(in[1106]), .B(n4002), .Z(n4820) );
  NANDN U5855 ( .A(n4823), .B(n4820), .Z(n4003) );
  XNOR U5856 ( .A(n4414), .B(n4003), .Z(out[664]) );
  XOR U5857 ( .A(in[263]), .B(n4004), .Z(n4417) );
  XOR U5858 ( .A(in[1496]), .B(n4005), .Z(n4827) );
  XNOR U5859 ( .A(in[1107]), .B(n4006), .Z(n4824) );
  NANDN U5860 ( .A(n4827), .B(n4824), .Z(n4007) );
  XNOR U5861 ( .A(n4417), .B(n4007), .Z(out[665]) );
  XOR U5862 ( .A(in[264]), .B(n4008), .Z(n4420) );
  XOR U5863 ( .A(in[1497]), .B(n4009), .Z(n4831) );
  XNOR U5864 ( .A(in[1108]), .B(n4010), .Z(n4828) );
  NANDN U5865 ( .A(n4831), .B(n4828), .Z(n4011) );
  XNOR U5866 ( .A(n4420), .B(n4011), .Z(out[666]) );
  XOR U5867 ( .A(in[265]), .B(n4012), .Z(n4423) );
  XOR U5868 ( .A(in[1498]), .B(n4013), .Z(n4246) );
  IV U5869 ( .A(n4246), .Z(n4835) );
  XNOR U5870 ( .A(in[1109]), .B(n4014), .Z(n4832) );
  NANDN U5871 ( .A(n4835), .B(n4832), .Z(n4015) );
  XNOR U5872 ( .A(n4423), .B(n4015), .Z(out[667]) );
  XOR U5873 ( .A(in[266]), .B(n4016), .Z(n4426) );
  XOR U5874 ( .A(in[1499]), .B(n4017), .Z(n4249) );
  IV U5875 ( .A(n4249), .Z(n4839) );
  XNOR U5876 ( .A(in[1110]), .B(n4018), .Z(n4836) );
  NANDN U5877 ( .A(n4839), .B(n4836), .Z(n4019) );
  XNOR U5878 ( .A(n4426), .B(n4019), .Z(out[668]) );
  XOR U5879 ( .A(in[267]), .B(n4020), .Z(n4429) );
  XOR U5880 ( .A(in[1500]), .B(n4021), .Z(n4843) );
  XNOR U5881 ( .A(in[1111]), .B(n4022), .Z(n4840) );
  NANDN U5882 ( .A(n4843), .B(n4840), .Z(n4023) );
  XNOR U5883 ( .A(n4429), .B(n4023), .Z(out[669]) );
  ANDN U5884 ( .B(n4025), .A(n4024), .Z(n4026) );
  XOR U5885 ( .A(n4027), .B(n4026), .Z(out[66]) );
  XOR U5886 ( .A(in[268]), .B(n4028), .Z(n4432) );
  XOR U5887 ( .A(in[1501]), .B(n4029), .Z(n4847) );
  XNOR U5888 ( .A(in[1112]), .B(n4030), .Z(n4844) );
  NANDN U5889 ( .A(n4847), .B(n4844), .Z(n4031) );
  XNOR U5890 ( .A(n4432), .B(n4031), .Z(out[670]) );
  XOR U5891 ( .A(in[269]), .B(n4032), .Z(n4435) );
  XOR U5892 ( .A(in[1502]), .B(n4033), .Z(n4851) );
  XNOR U5893 ( .A(in[1113]), .B(n4034), .Z(n4848) );
  NANDN U5894 ( .A(n4851), .B(n4848), .Z(n4035) );
  XNOR U5895 ( .A(n4435), .B(n4035), .Z(out[671]) );
  XOR U5896 ( .A(in[270]), .B(n4036), .Z(n4446) );
  XOR U5897 ( .A(in[1503]), .B(n4037), .Z(n4855) );
  XNOR U5898 ( .A(in[1114]), .B(n4038), .Z(n4852) );
  NANDN U5899 ( .A(n4855), .B(n4852), .Z(n4039) );
  XNOR U5900 ( .A(n4446), .B(n4039), .Z(out[672]) );
  XOR U5901 ( .A(in[271]), .B(n4040), .Z(n4449) );
  XOR U5902 ( .A(in[1504]), .B(n4041), .Z(n4859) );
  XNOR U5903 ( .A(in[1115]), .B(n4042), .Z(n4856) );
  NANDN U5904 ( .A(n4859), .B(n4856), .Z(n4043) );
  XNOR U5905 ( .A(n4449), .B(n4043), .Z(out[673]) );
  XOR U5906 ( .A(in[272]), .B(n4044), .Z(n4452) );
  XOR U5907 ( .A(in[1505]), .B(n4045), .Z(n4867) );
  XNOR U5908 ( .A(in[1116]), .B(n4046), .Z(n4864) );
  NANDN U5909 ( .A(n4867), .B(n4864), .Z(n4047) );
  XNOR U5910 ( .A(n4452), .B(n4047), .Z(out[674]) );
  XNOR U5911 ( .A(in[273]), .B(n4048), .Z(n4455) );
  XOR U5912 ( .A(n4049), .B(in[1506]), .Z(n4871) );
  XNOR U5913 ( .A(in[1117]), .B(n4050), .Z(n4868) );
  NANDN U5914 ( .A(n4871), .B(n4868), .Z(n4051) );
  XNOR U5915 ( .A(n4455), .B(n4051), .Z(out[675]) );
  XOR U5916 ( .A(in[274]), .B(n4052), .Z(n4458) );
  XOR U5917 ( .A(n4053), .B(in[1507]), .Z(n4875) );
  XOR U5918 ( .A(in[1118]), .B(n4054), .Z(n4872) );
  NANDN U5919 ( .A(n4875), .B(n4872), .Z(n4055) );
  XNOR U5920 ( .A(n4458), .B(n4055), .Z(out[676]) );
  XOR U5921 ( .A(in[275]), .B(n4056), .Z(n4461) );
  XOR U5922 ( .A(n4057), .B(in[1508]), .Z(n4879) );
  XOR U5923 ( .A(in[1119]), .B(n4058), .Z(n4876) );
  NANDN U5924 ( .A(n4879), .B(n4876), .Z(n4059) );
  XNOR U5925 ( .A(n4461), .B(n4059), .Z(out[677]) );
  XOR U5926 ( .A(in[276]), .B(n4060), .Z(n4464) );
  XOR U5927 ( .A(n4061), .B(in[1509]), .Z(n4883) );
  XOR U5928 ( .A(in[1120]), .B(n4062), .Z(n4880) );
  NANDN U5929 ( .A(n4883), .B(n4880), .Z(n4063) );
  XNOR U5930 ( .A(n4464), .B(n4063), .Z(out[678]) );
  XOR U5931 ( .A(in[277]), .B(n4064), .Z(n4467) );
  XOR U5932 ( .A(in[1510]), .B(n4065), .Z(n4264) );
  IV U5933 ( .A(n4264), .Z(n4887) );
  XOR U5934 ( .A(in[1121]), .B(n4066), .Z(n4884) );
  NANDN U5935 ( .A(n4887), .B(n4884), .Z(n4067) );
  XNOR U5936 ( .A(n4467), .B(n4067), .Z(out[679]) );
  ANDN U5937 ( .B(n4069), .A(n4068), .Z(n4070) );
  XOR U5938 ( .A(n4071), .B(n4070), .Z(out[67]) );
  XOR U5939 ( .A(in[278]), .B(n4072), .Z(n4470) );
  XOR U5940 ( .A(in[1511]), .B(n4073), .Z(n4267) );
  IV U5941 ( .A(n4267), .Z(n4891) );
  XOR U5942 ( .A(in[1122]), .B(n4074), .Z(n4888) );
  NANDN U5943 ( .A(n4891), .B(n4888), .Z(n4075) );
  XNOR U5944 ( .A(n4470), .B(n4075), .Z(out[680]) );
  XOR U5945 ( .A(in[279]), .B(n4076), .Z(n4473) );
  XOR U5946 ( .A(in[1512]), .B(n4077), .Z(n4270) );
  IV U5947 ( .A(n4270), .Z(n4895) );
  XOR U5948 ( .A(in[1123]), .B(n4078), .Z(n4892) );
  NANDN U5949 ( .A(n4895), .B(n4892), .Z(n4079) );
  XNOR U5950 ( .A(n4473), .B(n4079), .Z(out[681]) );
  XOR U5951 ( .A(in[280]), .B(n4080), .Z(n4480) );
  XOR U5952 ( .A(in[1513]), .B(n4081), .Z(n4273) );
  IV U5953 ( .A(n4273), .Z(n4899) );
  XOR U5954 ( .A(in[1124]), .B(n4082), .Z(n4896) );
  NANDN U5955 ( .A(n4899), .B(n4896), .Z(n4083) );
  XNOR U5956 ( .A(n4480), .B(n4083), .Z(out[682]) );
  XOR U5957 ( .A(in[281]), .B(n4084), .Z(n4483) );
  XOR U5958 ( .A(in[1514]), .B(n4085), .Z(n4276) );
  IV U5959 ( .A(n4276), .Z(n4903) );
  XNOR U5960 ( .A(in[1125]), .B(n4086), .Z(n4900) );
  NANDN U5961 ( .A(n4903), .B(n4900), .Z(n4087) );
  XNOR U5962 ( .A(n4483), .B(n4087), .Z(out[683]) );
  XOR U5963 ( .A(in[282]), .B(n4088), .Z(n4486) );
  XOR U5964 ( .A(in[1126]), .B(n4089), .Z(n4909) );
  XNOR U5965 ( .A(in[1515]), .B(n4090), .Z(n4911) );
  NANDN U5966 ( .A(n4909), .B(n4911), .Z(n4091) );
  XNOR U5967 ( .A(n4486), .B(n4091), .Z(out[684]) );
  XOR U5968 ( .A(in[283]), .B(n4092), .Z(n4489) );
  XOR U5969 ( .A(in[1127]), .B(n4093), .Z(n4913) );
  XNOR U5970 ( .A(in[1516]), .B(n4094), .Z(n4915) );
  NANDN U5971 ( .A(n4913), .B(n4915), .Z(n4095) );
  XNOR U5972 ( .A(n4489), .B(n4095), .Z(out[685]) );
  XOR U5973 ( .A(in[284]), .B(n4096), .Z(n4492) );
  XOR U5974 ( .A(in[1128]), .B(n4097), .Z(n4917) );
  XNOR U5975 ( .A(in[1517]), .B(n4098), .Z(n4919) );
  NANDN U5976 ( .A(n4917), .B(n4919), .Z(n4099) );
  XNOR U5977 ( .A(n4492), .B(n4099), .Z(out[686]) );
  XOR U5978 ( .A(in[285]), .B(n4100), .Z(n4495) );
  XOR U5979 ( .A(in[1129]), .B(n4101), .Z(n4921) );
  XNOR U5980 ( .A(in[1518]), .B(n4102), .Z(n4923) );
  NANDN U5981 ( .A(n4921), .B(n4923), .Z(n4103) );
  XNOR U5982 ( .A(n4495), .B(n4103), .Z(out[687]) );
  XOR U5983 ( .A(in[286]), .B(n4104), .Z(n4498) );
  XOR U5984 ( .A(in[1130]), .B(n4105), .Z(n4925) );
  XNOR U5985 ( .A(in[1519]), .B(n4106), .Z(n4927) );
  NANDN U5986 ( .A(n4925), .B(n4927), .Z(n4107) );
  XNOR U5987 ( .A(n4498), .B(n4107), .Z(out[688]) );
  XOR U5988 ( .A(in[287]), .B(n4108), .Z(n4501) );
  XNOR U5989 ( .A(in[1131]), .B(n4109), .Z(n4929) );
  XNOR U5990 ( .A(in[1520]), .B(n4110), .Z(n4931) );
  NANDN U5991 ( .A(n4929), .B(n4931), .Z(n4111) );
  XNOR U5992 ( .A(n4501), .B(n4111), .Z(out[689]) );
  ANDN U5993 ( .B(n4113), .A(n4112), .Z(n4114) );
  XOR U5994 ( .A(n4115), .B(n4114), .Z(out[68]) );
  XOR U5995 ( .A(in[288]), .B(n4116), .Z(n4504) );
  XNOR U5996 ( .A(in[1132]), .B(n4117), .Z(n4933) );
  XNOR U5997 ( .A(in[1521]), .B(n4118), .Z(n4935) );
  NANDN U5998 ( .A(n4933), .B(n4935), .Z(n4119) );
  XNOR U5999 ( .A(n4504), .B(n4119), .Z(out[690]) );
  XOR U6000 ( .A(in[289]), .B(n4120), .Z(n4507) );
  XOR U6001 ( .A(in[1133]), .B(n4121), .Z(n4937) );
  XNOR U6002 ( .A(in[1522]), .B(n4122), .Z(n4939) );
  NANDN U6003 ( .A(n4937), .B(n4939), .Z(n4123) );
  XNOR U6004 ( .A(n4507), .B(n4123), .Z(out[691]) );
  XNOR U6005 ( .A(in[290]), .B(n4124), .Z(n4514) );
  XOR U6006 ( .A(in[1134]), .B(n4125), .Z(n4941) );
  XNOR U6007 ( .A(in[1523]), .B(n4126), .Z(n4943) );
  NANDN U6008 ( .A(n4941), .B(n4943), .Z(n4127) );
  XNOR U6009 ( .A(n4514), .B(n4127), .Z(out[692]) );
  XOR U6010 ( .A(in[291]), .B(n4128), .Z(n4517) );
  XOR U6011 ( .A(in[1135]), .B(n4129), .Z(n4945) );
  XNOR U6012 ( .A(in[1524]), .B(n4130), .Z(n4947) );
  NANDN U6013 ( .A(n4945), .B(n4947), .Z(n4131) );
  XNOR U6014 ( .A(n4517), .B(n4131), .Z(out[693]) );
  XOR U6015 ( .A(in[292]), .B(n4132), .Z(n4520) );
  XOR U6016 ( .A(in[1136]), .B(n4133), .Z(n4953) );
  XNOR U6017 ( .A(in[1525]), .B(n4134), .Z(n4955) );
  NANDN U6018 ( .A(n4953), .B(n4955), .Z(n4135) );
  XNOR U6019 ( .A(n4520), .B(n4135), .Z(out[694]) );
  XOR U6020 ( .A(in[293]), .B(n4136), .Z(n4305) );
  IV U6021 ( .A(n4305), .Z(n4524) );
  XOR U6022 ( .A(in[1137]), .B(n4137), .Z(n4957) );
  XNOR U6023 ( .A(in[1526]), .B(n4138), .Z(n4959) );
  NANDN U6024 ( .A(n4957), .B(n4959), .Z(n4139) );
  XOR U6025 ( .A(n4524), .B(n4139), .Z(out[695]) );
  XOR U6026 ( .A(in[294]), .B(n4140), .Z(n4312) );
  IV U6027 ( .A(n4312), .Z(n4528) );
  XOR U6028 ( .A(in[1138]), .B(n4141), .Z(n4961) );
  XNOR U6029 ( .A(in[1527]), .B(n4142), .Z(n4963) );
  NANDN U6030 ( .A(n4961), .B(n4963), .Z(n4143) );
  XOR U6031 ( .A(n4528), .B(n4143), .Z(out[696]) );
  XOR U6032 ( .A(in[295]), .B(n4144), .Z(n4315) );
  IV U6033 ( .A(n4315), .Z(n4532) );
  XOR U6034 ( .A(in[1139]), .B(n4145), .Z(n4965) );
  XNOR U6035 ( .A(in[1528]), .B(n4146), .Z(n4967) );
  NANDN U6036 ( .A(n4965), .B(n4967), .Z(n4147) );
  XOR U6037 ( .A(n4532), .B(n4147), .Z(out[697]) );
  XOR U6038 ( .A(in[296]), .B(n4148), .Z(n4318) );
  IV U6039 ( .A(n4318), .Z(n4536) );
  XOR U6040 ( .A(in[1140]), .B(n4149), .Z(n4969) );
  XNOR U6041 ( .A(in[1529]), .B(n4150), .Z(n4971) );
  NANDN U6042 ( .A(n4969), .B(n4971), .Z(n4151) );
  XOR U6043 ( .A(n4536), .B(n4151), .Z(out[698]) );
  XOR U6044 ( .A(in[297]), .B(n4152), .Z(n4321) );
  IV U6045 ( .A(n4321), .Z(n4540) );
  XNOR U6046 ( .A(in[1141]), .B(n4153), .Z(n4973) );
  XNOR U6047 ( .A(in[1530]), .B(n4154), .Z(n4975) );
  NANDN U6048 ( .A(n4973), .B(n4975), .Z(n4155) );
  XOR U6049 ( .A(n4540), .B(n4155), .Z(out[699]) );
  ANDN U6050 ( .B(n4157), .A(n4156), .Z(n4158) );
  XOR U6051 ( .A(n4159), .B(n4158), .Z(out[69]) );
  OR U6052 ( .A(n4195), .B(n4160), .Z(n4161) );
  XNOR U6053 ( .A(n4194), .B(n4161), .Z(out[6]) );
  XOR U6054 ( .A(in[298]), .B(n4162), .Z(n4324) );
  IV U6055 ( .A(n4324), .Z(n4544) );
  XNOR U6056 ( .A(in[1142]), .B(n4163), .Z(n4977) );
  XNOR U6057 ( .A(in[1531]), .B(n4164), .Z(n4979) );
  OR U6058 ( .A(n4977), .B(n4979), .Z(n4165) );
  XOR U6059 ( .A(n4544), .B(n4165), .Z(out[700]) );
  XOR U6060 ( .A(in[299]), .B(n4166), .Z(n4327) );
  IV U6061 ( .A(n4327), .Z(n4547) );
  XNOR U6062 ( .A(in[1143]), .B(n4167), .Z(n4981) );
  XNOR U6063 ( .A(in[1532]), .B(n4168), .Z(n4983) );
  OR U6064 ( .A(n4981), .B(n4983), .Z(n4169) );
  XOR U6065 ( .A(n4547), .B(n4169), .Z(out[701]) );
  XOR U6066 ( .A(in[300]), .B(n4170), .Z(n4330) );
  IV U6067 ( .A(n4330), .Z(n4553) );
  XNOR U6068 ( .A(in[1144]), .B(n4171), .Z(n4985) );
  XNOR U6069 ( .A(in[1533]), .B(n4172), .Z(n4987) );
  OR U6070 ( .A(n4985), .B(n4987), .Z(n4173) );
  XOR U6071 ( .A(n4553), .B(n4173), .Z(out[702]) );
  XOR U6072 ( .A(in[301]), .B(n4174), .Z(n4333) );
  IV U6073 ( .A(n4333), .Z(n4555) );
  XNOR U6074 ( .A(in[1145]), .B(n4175), .Z(n4989) );
  XNOR U6075 ( .A(in[1534]), .B(n4176), .Z(n4991) );
  NANDN U6076 ( .A(n4989), .B(n4991), .Z(n4177) );
  XOR U6077 ( .A(n4555), .B(n4177), .Z(out[703]) );
  XOR U6078 ( .A(in[376]), .B(n4178), .Z(n4556) );
  ANDN U6079 ( .B(n4711), .A(n4179), .Z(n4180) );
  XOR U6080 ( .A(n4556), .B(n4180), .Z(out[704]) );
  XOR U6081 ( .A(in[377]), .B(n4181), .Z(n4559) );
  ANDN U6082 ( .B(n4715), .A(n4182), .Z(n4183) );
  XOR U6083 ( .A(n4559), .B(n4183), .Z(out[705]) );
  XOR U6084 ( .A(in[378]), .B(n4184), .Z(n4562) );
  ANDN U6085 ( .B(n4719), .A(n4185), .Z(n4186) );
  XOR U6086 ( .A(n4562), .B(n4186), .Z(out[706]) );
  XOR U6087 ( .A(in[379]), .B(n4187), .Z(n4565) );
  ANDN U6088 ( .B(n4723), .A(n4188), .Z(n4189) );
  XOR U6089 ( .A(n4565), .B(n4189), .Z(out[707]) );
  XOR U6090 ( .A(in[380]), .B(n4190), .Z(n4568) );
  ANDN U6091 ( .B(n4735), .A(n4191), .Z(n4192) );
  XNOR U6092 ( .A(n4568), .B(n4192), .Z(out[708]) );
  XOR U6093 ( .A(in[381]), .B(n4193), .Z(n4570) );
  ANDN U6094 ( .B(n4195), .A(n4194), .Z(n4196) );
  XOR U6095 ( .A(n4197), .B(n4196), .Z(out[70]) );
  XOR U6096 ( .A(in[382]), .B(n4198), .Z(n4572) );
  XOR U6097 ( .A(in[383]), .B(n4199), .Z(n4574) );
  XOR U6098 ( .A(in[320]), .B(n4200), .Z(n4581) );
  XOR U6099 ( .A(in[321]), .B(n4201), .Z(n4583) );
  XOR U6100 ( .A(in[322]), .B(n4202), .Z(n4585) );
  XOR U6101 ( .A(in[323]), .B(n4203), .Z(n4587) );
  XOR U6102 ( .A(in[324]), .B(n4204), .Z(n4589) );
  XOR U6103 ( .A(in[325]), .B(n4205), .Z(n4591) );
  ANDN U6104 ( .B(n4771), .A(n4206), .Z(n4207) );
  XNOR U6105 ( .A(n4591), .B(n4207), .Z(out[717]) );
  XOR U6106 ( .A(in[326]), .B(n4208), .Z(n4593) );
  ANDN U6107 ( .B(n4779), .A(n4209), .Z(n4210) );
  XNOR U6108 ( .A(n4593), .B(n4210), .Z(out[718]) );
  XOR U6109 ( .A(in[327]), .B(n4211), .Z(n4595) );
  ANDN U6110 ( .B(n4783), .A(n4212), .Z(n4213) );
  XNOR U6111 ( .A(n4595), .B(n4213), .Z(out[719]) );
  ANDN U6112 ( .B(n4442), .A(n4444), .Z(n4214) );
  XOR U6113 ( .A(n4215), .B(n4214), .Z(out[71]) );
  XOR U6114 ( .A(in[328]), .B(n4216), .Z(n4597) );
  ANDN U6115 ( .B(n4787), .A(n4217), .Z(n4218) );
  XOR U6116 ( .A(n4597), .B(n4218), .Z(out[720]) );
  XOR U6117 ( .A(in[329]), .B(n4219), .Z(n4600) );
  ANDN U6118 ( .B(n4791), .A(n4220), .Z(n4221) );
  XNOR U6119 ( .A(n4600), .B(n4221), .Z(out[721]) );
  XOR U6120 ( .A(in[330]), .B(n4222), .Z(n4606) );
  ANDN U6121 ( .B(n4795), .A(n4223), .Z(n4224) );
  XNOR U6122 ( .A(n4606), .B(n4224), .Z(out[722]) );
  XOR U6123 ( .A(in[331]), .B(n4225), .Z(n4608) );
  ANDN U6124 ( .B(n4799), .A(n4226), .Z(n4227) );
  XNOR U6125 ( .A(n4608), .B(n4227), .Z(out[723]) );
  XOR U6126 ( .A(in[332]), .B(n4228), .Z(n4610) );
  ANDN U6127 ( .B(n4803), .A(n4229), .Z(n4230) );
  XNOR U6128 ( .A(n4610), .B(n4230), .Z(out[724]) );
  XOR U6129 ( .A(in[333]), .B(n4231), .Z(n4612) );
  ANDN U6130 ( .B(n4807), .A(n4232), .Z(n4233) );
  XNOR U6131 ( .A(n4612), .B(n4233), .Z(out[725]) );
  XOR U6132 ( .A(in[334]), .B(n4234), .Z(n4614) );
  NOR U6133 ( .A(n4235), .B(n4408), .Z(n4236) );
  XOR U6134 ( .A(n4614), .B(n4236), .Z(out[726]) );
  XOR U6135 ( .A(in[335]), .B(n4237), .Z(n4617) );
  NOR U6136 ( .A(n4238), .B(n4411), .Z(n4239) );
  XOR U6137 ( .A(n4617), .B(n4239), .Z(out[727]) );
  XOR U6138 ( .A(in[336]), .B(n4240), .Z(n4620) );
  XOR U6139 ( .A(in[337]), .B(n4241), .Z(n4623) );
  ANDN U6140 ( .B(n4729), .A(n4731), .Z(n4242) );
  XOR U6141 ( .A(n4243), .B(n4242), .Z(out[72]) );
  XOR U6142 ( .A(in[338]), .B(n4244), .Z(n4626) );
  XOR U6143 ( .A(in[339]), .B(n4245), .Z(n4628) );
  NOR U6144 ( .A(n4246), .B(n4423), .Z(n4247) );
  XNOR U6145 ( .A(n4628), .B(n4247), .Z(out[731]) );
  XOR U6146 ( .A(in[340]), .B(n4248), .Z(n4633) );
  NOR U6147 ( .A(n4249), .B(n4426), .Z(n4250) );
  XOR U6148 ( .A(n4633), .B(n4250), .Z(out[732]) );
  XOR U6149 ( .A(in[341]), .B(n4251), .Z(n4636) );
  XOR U6150 ( .A(in[342]), .B(n4252), .Z(n4639) );
  XOR U6151 ( .A(in[343]), .B(n4253), .Z(n4642) );
  XOR U6152 ( .A(in[344]), .B(n4254), .Z(n4643) );
  XOR U6153 ( .A(in[345]), .B(n4255), .Z(n4646) );
  XOR U6154 ( .A(in[346]), .B(n4256), .Z(n4649) );
  XOR U6155 ( .A(in[347]), .B(n4257), .Z(n4652) );
  ANDN U6156 ( .B(n5160), .A(n5162), .Z(n4258) );
  XOR U6157 ( .A(n4259), .B(n4258), .Z(out[73]) );
  XOR U6158 ( .A(in[348]), .B(n4260), .Z(n4655) );
  XOR U6159 ( .A(in[349]), .B(n4261), .Z(n4658) );
  XOR U6160 ( .A(in[350]), .B(n4262), .Z(n4663) );
  XOR U6161 ( .A(in[351]), .B(n4263), .Z(n4664) );
  NOR U6162 ( .A(n4264), .B(n4467), .Z(n4265) );
  XOR U6163 ( .A(n4664), .B(n4265), .Z(out[743]) );
  XOR U6164 ( .A(in[352]), .B(n4266), .Z(n4665) );
  NOR U6165 ( .A(n4267), .B(n4470), .Z(n4268) );
  XOR U6166 ( .A(n4665), .B(n4268), .Z(out[744]) );
  XOR U6167 ( .A(in[353]), .B(n4269), .Z(n4666) );
  NOR U6168 ( .A(n4270), .B(n4473), .Z(n4271) );
  XOR U6169 ( .A(n4666), .B(n4271), .Z(out[745]) );
  XOR U6170 ( .A(in[354]), .B(n4272), .Z(n4667) );
  NOR U6171 ( .A(n4273), .B(n4480), .Z(n4274) );
  XOR U6172 ( .A(n4667), .B(n4274), .Z(out[746]) );
  XOR U6173 ( .A(in[355]), .B(n4275), .Z(n4668) );
  NOR U6174 ( .A(n4276), .B(n4483), .Z(n4277) );
  XNOR U6175 ( .A(n4668), .B(n4277), .Z(out[747]) );
  XOR U6176 ( .A(in[356]), .B(n4278), .Z(n4670) );
  NOR U6177 ( .A(n4911), .B(n4486), .Z(n4279) );
  XOR U6178 ( .A(n4670), .B(n4279), .Z(out[748]) );
  XOR U6179 ( .A(in[357]), .B(n4280), .Z(n4671) );
  NOR U6180 ( .A(n4915), .B(n4489), .Z(n4281) );
  XOR U6181 ( .A(n4671), .B(n4281), .Z(out[749]) );
  ANDN U6182 ( .B(n4283), .A(n4282), .Z(n4284) );
  XOR U6183 ( .A(n4285), .B(n4284), .Z(out[74]) );
  XOR U6184 ( .A(in[358]), .B(n4286), .Z(n4672) );
  NOR U6185 ( .A(n4919), .B(n4492), .Z(n4287) );
  XOR U6186 ( .A(n4672), .B(n4287), .Z(out[750]) );
  XOR U6187 ( .A(in[359]), .B(n4288), .Z(n4673) );
  NOR U6188 ( .A(n4923), .B(n4495), .Z(n4289) );
  XOR U6189 ( .A(n4673), .B(n4289), .Z(out[751]) );
  XOR U6190 ( .A(in[360]), .B(n4290), .Z(n4677) );
  NOR U6191 ( .A(n4927), .B(n4498), .Z(n4291) );
  XOR U6192 ( .A(n4677), .B(n4291), .Z(out[752]) );
  XOR U6193 ( .A(in[361]), .B(n4292), .Z(n4678) );
  NOR U6194 ( .A(n4931), .B(n4501), .Z(n4293) );
  XOR U6195 ( .A(n4678), .B(n4293), .Z(out[753]) );
  XOR U6196 ( .A(in[362]), .B(n4294), .Z(n4679) );
  NOR U6197 ( .A(n4935), .B(n4504), .Z(n4295) );
  XOR U6198 ( .A(n4679), .B(n4295), .Z(out[754]) );
  XOR U6199 ( .A(in[363]), .B(n4296), .Z(n4680) );
  NOR U6200 ( .A(n4939), .B(n4507), .Z(n4297) );
  XOR U6201 ( .A(n4680), .B(n4297), .Z(out[755]) );
  XOR U6202 ( .A(in[364]), .B(n4298), .Z(n4681) );
  NOR U6203 ( .A(n4943), .B(n4514), .Z(n4299) );
  XOR U6204 ( .A(n4681), .B(n4299), .Z(out[756]) );
  XOR U6205 ( .A(in[365]), .B(n4300), .Z(n4682) );
  NOR U6206 ( .A(n4947), .B(n4517), .Z(n4301) );
  XOR U6207 ( .A(n4682), .B(n4301), .Z(out[757]) );
  XOR U6208 ( .A(in[366]), .B(n4302), .Z(n4683) );
  NOR U6209 ( .A(n4955), .B(n4520), .Z(n4303) );
  XOR U6210 ( .A(n4683), .B(n4303), .Z(out[758]) );
  XOR U6211 ( .A(in[367]), .B(n4304), .Z(n4523) );
  NOR U6212 ( .A(n4305), .B(n4959), .Z(n4306) );
  XOR U6213 ( .A(n4523), .B(n4306), .Z(out[759]) );
  ANDN U6214 ( .B(n4308), .A(n4307), .Z(n4309) );
  XOR U6215 ( .A(n4310), .B(n4309), .Z(out[75]) );
  XOR U6216 ( .A(in[368]), .B(n4311), .Z(n4527) );
  NOR U6217 ( .A(n4312), .B(n4963), .Z(n4313) );
  XOR U6218 ( .A(n4527), .B(n4313), .Z(out[760]) );
  XOR U6219 ( .A(in[369]), .B(n4314), .Z(n4531) );
  NOR U6220 ( .A(n4315), .B(n4967), .Z(n4316) );
  XOR U6221 ( .A(n4531), .B(n4316), .Z(out[761]) );
  XOR U6222 ( .A(in[370]), .B(n4317), .Z(n4535) );
  NOR U6223 ( .A(n4318), .B(n4971), .Z(n4319) );
  XOR U6224 ( .A(n4535), .B(n4319), .Z(out[762]) );
  XOR U6225 ( .A(in[371]), .B(n4320), .Z(n4539) );
  NOR U6226 ( .A(n4321), .B(n4975), .Z(n4322) );
  XOR U6227 ( .A(n4539), .B(n4322), .Z(out[763]) );
  XOR U6228 ( .A(in[372]), .B(n4323), .Z(n4543) );
  ANDN U6229 ( .B(n4979), .A(n4324), .Z(n4325) );
  XOR U6230 ( .A(n4543), .B(n4325), .Z(out[764]) );
  XOR U6231 ( .A(in[373]), .B(n4326), .Z(n4699) );
  ANDN U6232 ( .B(n4983), .A(n4327), .Z(n4328) );
  XOR U6233 ( .A(n4699), .B(n4328), .Z(out[765]) );
  XOR U6234 ( .A(in[374]), .B(n4329), .Z(n4702) );
  ANDN U6235 ( .B(n4987), .A(n4330), .Z(n4331) );
  XOR U6236 ( .A(n4702), .B(n4331), .Z(out[766]) );
  XOR U6237 ( .A(in[375]), .B(n4332), .Z(n4705) );
  NOR U6238 ( .A(n4333), .B(n4991), .Z(n4334) );
  XOR U6239 ( .A(n4705), .B(n4334), .Z(out[767]) );
  XOR U6240 ( .A(in[743]), .B(n4335), .Z(n4557) );
  IV U6241 ( .A(n4557), .Z(n4708) );
  XOR U6242 ( .A(in[744]), .B(n4337), .Z(n4560) );
  IV U6243 ( .A(n4560), .Z(n4712) );
  ANDN U6244 ( .B(n4340), .A(n4339), .Z(n4341) );
  XOR U6245 ( .A(n4342), .B(n4341), .Z(out[76]) );
  XOR U6246 ( .A(in[745]), .B(n4343), .Z(n4563) );
  IV U6247 ( .A(n4563), .Z(n4716) );
  XOR U6248 ( .A(in[746]), .B(n4345), .Z(n4566) );
  IV U6249 ( .A(n4566), .Z(n4720) );
  XNOR U6250 ( .A(in[747]), .B(n4347), .Z(n4732) );
  NANDN U6251 ( .A(n4348), .B(n4568), .Z(n4349) );
  XOR U6252 ( .A(n4732), .B(n4349), .Z(out[772]) );
  XNOR U6253 ( .A(in[748]), .B(n4350), .Z(n4736) );
  NANDN U6254 ( .A(n4351), .B(n4570), .Z(n4352) );
  XOR U6255 ( .A(n4736), .B(n4352), .Z(out[773]) );
  XNOR U6256 ( .A(in[749]), .B(n4353), .Z(n4740) );
  NANDN U6257 ( .A(n4354), .B(n4572), .Z(n4355) );
  XOR U6258 ( .A(n4740), .B(n4355), .Z(out[774]) );
  XOR U6259 ( .A(in[750]), .B(n4356), .Z(n4575) );
  IV U6260 ( .A(n4575), .Z(n4744) );
  XNOR U6261 ( .A(in[751]), .B(n4358), .Z(n4749) );
  NANDN U6262 ( .A(n4359), .B(n4581), .Z(n4360) );
  XOR U6263 ( .A(n4749), .B(n4360), .Z(out[776]) );
  XNOR U6264 ( .A(in[752]), .B(n4361), .Z(n4753) );
  NANDN U6265 ( .A(n4362), .B(n4583), .Z(n4363) );
  XOR U6266 ( .A(n4753), .B(n4363), .Z(out[777]) );
  XNOR U6267 ( .A(in[753]), .B(n4364), .Z(n4757) );
  NANDN U6268 ( .A(n4365), .B(n4585), .Z(n4366) );
  XOR U6269 ( .A(n4757), .B(n4366), .Z(out[778]) );
  XNOR U6270 ( .A(in[754]), .B(n4367), .Z(n4761) );
  NANDN U6271 ( .A(n4368), .B(n4587), .Z(n4369) );
  XOR U6272 ( .A(n4761), .B(n4369), .Z(out[779]) );
  ANDN U6273 ( .B(n4371), .A(n4370), .Z(n4372) );
  XOR U6274 ( .A(n4373), .B(n4372), .Z(out[77]) );
  XNOR U6275 ( .A(in[755]), .B(n4374), .Z(n4765) );
  NANDN U6276 ( .A(n4375), .B(n4589), .Z(n4376) );
  XOR U6277 ( .A(n4765), .B(n4376), .Z(out[780]) );
  XNOR U6278 ( .A(in[756]), .B(n4377), .Z(n4769) );
  NANDN U6279 ( .A(n4378), .B(n4591), .Z(n4379) );
  XOR U6280 ( .A(n4769), .B(n4379), .Z(out[781]) );
  XNOR U6281 ( .A(in[757]), .B(n4380), .Z(n4777) );
  NANDN U6282 ( .A(n4381), .B(n4593), .Z(n4382) );
  XOR U6283 ( .A(n4777), .B(n4382), .Z(out[782]) );
  XNOR U6284 ( .A(in[758]), .B(n4383), .Z(n4781) );
  NANDN U6285 ( .A(n4384), .B(n4595), .Z(n4385) );
  XOR U6286 ( .A(n4781), .B(n4385), .Z(out[783]) );
  XOR U6287 ( .A(in[759]), .B(n4386), .Z(n4598) );
  IV U6288 ( .A(n4598), .Z(n4785) );
  XNOR U6289 ( .A(in[760]), .B(n4388), .Z(n4789) );
  NANDN U6290 ( .A(n4389), .B(n4600), .Z(n4390) );
  XOR U6291 ( .A(n4789), .B(n4390), .Z(out[785]) );
  XNOR U6292 ( .A(in[761]), .B(n4391), .Z(n4793) );
  NANDN U6293 ( .A(n4392), .B(n4606), .Z(n4393) );
  XOR U6294 ( .A(n4793), .B(n4393), .Z(out[786]) );
  XOR U6295 ( .A(in[762]), .B(n4394), .Z(n4797) );
  NANDN U6296 ( .A(n4395), .B(n4608), .Z(n4396) );
  XOR U6297 ( .A(n4797), .B(n4396), .Z(out[787]) );
  XOR U6298 ( .A(in[763]), .B(n4397), .Z(n4801) );
  NANDN U6299 ( .A(n4398), .B(n4610), .Z(n4399) );
  XOR U6300 ( .A(n4801), .B(n4399), .Z(out[788]) );
  XNOR U6301 ( .A(in[764]), .B(n4400), .Z(n4805) );
  NANDN U6302 ( .A(n4401), .B(n4612), .Z(n4402) );
  XOR U6303 ( .A(n4805), .B(n4402), .Z(out[789]) );
  ANDN U6304 ( .B(n4404), .A(n4403), .Z(n4405) );
  XOR U6305 ( .A(n4406), .B(n4405), .Z(out[78]) );
  XOR U6306 ( .A(in[765]), .B(n4407), .Z(n4615) );
  IV U6307 ( .A(n4615), .Z(n4809) );
  NANDN U6308 ( .A(n4614), .B(n4408), .Z(n4409) );
  XOR U6309 ( .A(n4809), .B(n4409), .Z(out[790]) );
  XOR U6310 ( .A(in[766]), .B(n4410), .Z(n4618) );
  IV U6311 ( .A(n4618), .Z(n4813) );
  NANDN U6312 ( .A(n4617), .B(n4411), .Z(n4412) );
  XOR U6313 ( .A(n4813), .B(n4412), .Z(out[791]) );
  XOR U6314 ( .A(in[767]), .B(n4413), .Z(n4621) );
  IV U6315 ( .A(n4621), .Z(n4821) );
  NANDN U6316 ( .A(n4620), .B(n4414), .Z(n4415) );
  XOR U6317 ( .A(n4821), .B(n4415), .Z(out[792]) );
  XOR U6318 ( .A(in[704]), .B(n4416), .Z(n4624) );
  IV U6319 ( .A(n4624), .Z(n4825) );
  NANDN U6320 ( .A(n4623), .B(n4417), .Z(n4418) );
  XOR U6321 ( .A(n4825), .B(n4418), .Z(out[793]) );
  XNOR U6322 ( .A(in[705]), .B(n4419), .Z(n4829) );
  NAND U6323 ( .A(n4420), .B(n4626), .Z(n4421) );
  XOR U6324 ( .A(n4829), .B(n4421), .Z(out[794]) );
  XNOR U6325 ( .A(in[706]), .B(n4422), .Z(n4833) );
  NAND U6326 ( .A(n4423), .B(n4628), .Z(n4424) );
  XOR U6327 ( .A(n4833), .B(n4424), .Z(out[795]) );
  XOR U6328 ( .A(in[707]), .B(n4425), .Z(n4634) );
  IV U6329 ( .A(n4634), .Z(n4837) );
  NANDN U6330 ( .A(n4633), .B(n4426), .Z(n4427) );
  XOR U6331 ( .A(n4837), .B(n4427), .Z(out[796]) );
  XOR U6332 ( .A(in[708]), .B(n4428), .Z(n4637) );
  IV U6333 ( .A(n4637), .Z(n4841) );
  NANDN U6334 ( .A(n4636), .B(n4429), .Z(n4430) );
  XOR U6335 ( .A(n4841), .B(n4430), .Z(out[797]) );
  XOR U6336 ( .A(in[709]), .B(n4431), .Z(n4640) );
  IV U6337 ( .A(n4640), .Z(n4845) );
  NANDN U6338 ( .A(n4639), .B(n4432), .Z(n4433) );
  XOR U6339 ( .A(n4845), .B(n4433), .Z(out[798]) );
  XOR U6340 ( .A(in[710]), .B(n4434), .Z(n4849) );
  NANDN U6341 ( .A(n4642), .B(n4435), .Z(n4436) );
  XOR U6342 ( .A(n4849), .B(n4436), .Z(out[799]) );
  ANDN U6343 ( .B(n4438), .A(n4437), .Z(n4439) );
  XOR U6344 ( .A(n4440), .B(n4439), .Z(out[79]) );
  OR U6345 ( .A(n4442), .B(n4441), .Z(n4443) );
  XNOR U6346 ( .A(n4444), .B(n4443), .Z(out[7]) );
  XOR U6347 ( .A(in[711]), .B(n4445), .Z(n4644) );
  IV U6348 ( .A(n4644), .Z(n4853) );
  NANDN U6349 ( .A(n4643), .B(n4446), .Z(n4447) );
  XOR U6350 ( .A(n4853), .B(n4447), .Z(out[800]) );
  XOR U6351 ( .A(in[712]), .B(n4448), .Z(n4647) );
  IV U6352 ( .A(n4647), .Z(n4857) );
  NANDN U6353 ( .A(n4646), .B(n4449), .Z(n4450) );
  XOR U6354 ( .A(n4857), .B(n4450), .Z(out[801]) );
  XOR U6355 ( .A(in[713]), .B(n4451), .Z(n4650) );
  IV U6356 ( .A(n4650), .Z(n4865) );
  NANDN U6357 ( .A(n4649), .B(n4452), .Z(n4453) );
  XOR U6358 ( .A(n4865), .B(n4453), .Z(out[802]) );
  XOR U6359 ( .A(in[714]), .B(n4454), .Z(n4653) );
  IV U6360 ( .A(n4653), .Z(n4869) );
  NANDN U6361 ( .A(n4652), .B(n4455), .Z(n4456) );
  XOR U6362 ( .A(n4869), .B(n4456), .Z(out[803]) );
  XOR U6363 ( .A(in[715]), .B(n4457), .Z(n4656) );
  IV U6364 ( .A(n4656), .Z(n4873) );
  NANDN U6365 ( .A(n4655), .B(n4458), .Z(n4459) );
  XOR U6366 ( .A(n4873), .B(n4459), .Z(out[804]) );
  XNOR U6367 ( .A(n4460), .B(in[716]), .Z(n4877) );
  NANDN U6368 ( .A(n4658), .B(n4461), .Z(n4462) );
  XNOR U6369 ( .A(n4877), .B(n4462), .Z(out[805]) );
  XNOR U6370 ( .A(n4463), .B(in[717]), .Z(n4881) );
  NANDN U6371 ( .A(n4663), .B(n4464), .Z(n4465) );
  XNOR U6372 ( .A(n4881), .B(n4465), .Z(out[806]) );
  XNOR U6373 ( .A(n4466), .B(in[718]), .Z(n4885) );
  NANDN U6374 ( .A(n4664), .B(n4467), .Z(n4468) );
  XNOR U6375 ( .A(n4885), .B(n4468), .Z(out[807]) );
  XNOR U6376 ( .A(n4469), .B(in[719]), .Z(n4889) );
  NANDN U6377 ( .A(n4665), .B(n4470), .Z(n4471) );
  XNOR U6378 ( .A(n4889), .B(n4471), .Z(out[808]) );
  XNOR U6379 ( .A(n4472), .B(in[720]), .Z(n4893) );
  NANDN U6380 ( .A(n4666), .B(n4473), .Z(n4474) );
  XNOR U6381 ( .A(n4893), .B(n4474), .Z(out[809]) );
  ANDN U6382 ( .B(n4476), .A(n4475), .Z(n4477) );
  XOR U6383 ( .A(n4478), .B(n4477), .Z(out[80]) );
  XNOR U6384 ( .A(n4479), .B(in[721]), .Z(n4897) );
  NANDN U6385 ( .A(n4667), .B(n4480), .Z(n4481) );
  XNOR U6386 ( .A(n4897), .B(n4481), .Z(out[810]) );
  XNOR U6387 ( .A(n4482), .B(in[722]), .Z(n4901) );
  NAND U6388 ( .A(n4483), .B(n4668), .Z(n4484) );
  XNOR U6389 ( .A(n4901), .B(n4484), .Z(out[811]) );
  XNOR U6390 ( .A(n4485), .B(in[723]), .Z(n4908) );
  NANDN U6391 ( .A(n4670), .B(n4486), .Z(n4487) );
  XNOR U6392 ( .A(n4908), .B(n4487), .Z(out[812]) );
  XNOR U6393 ( .A(in[724]), .B(n4488), .Z(n4912) );
  NANDN U6394 ( .A(n4671), .B(n4489), .Z(n4490) );
  XNOR U6395 ( .A(n4912), .B(n4490), .Z(out[813]) );
  XNOR U6396 ( .A(in[725]), .B(n4491), .Z(n4916) );
  NANDN U6397 ( .A(n4672), .B(n4492), .Z(n4493) );
  XNOR U6398 ( .A(n4916), .B(n4493), .Z(out[814]) );
  XNOR U6399 ( .A(in[726]), .B(n4494), .Z(n4920) );
  NANDN U6400 ( .A(n4673), .B(n4495), .Z(n4496) );
  XNOR U6401 ( .A(n4920), .B(n4496), .Z(out[815]) );
  XNOR U6402 ( .A(in[727]), .B(n4497), .Z(n4924) );
  NANDN U6403 ( .A(n4677), .B(n4498), .Z(n4499) );
  XNOR U6404 ( .A(n4924), .B(n4499), .Z(out[816]) );
  XNOR U6405 ( .A(in[728]), .B(n4500), .Z(n4928) );
  NANDN U6406 ( .A(n4678), .B(n4501), .Z(n4502) );
  XNOR U6407 ( .A(n4928), .B(n4502), .Z(out[817]) );
  XNOR U6408 ( .A(in[729]), .B(n4503), .Z(n4932) );
  NANDN U6409 ( .A(n4679), .B(n4504), .Z(n4505) );
  XNOR U6410 ( .A(n4932), .B(n4505), .Z(out[818]) );
  XNOR U6411 ( .A(in[730]), .B(n4506), .Z(n4936) );
  NANDN U6412 ( .A(n4680), .B(n4507), .Z(n4508) );
  XNOR U6413 ( .A(n4936), .B(n4508), .Z(out[819]) );
  ANDN U6414 ( .B(n4510), .A(n4509), .Z(n4511) );
  XOR U6415 ( .A(n4512), .B(n4511), .Z(out[81]) );
  XOR U6416 ( .A(in[731]), .B(n4513), .Z(n4940) );
  NANDN U6417 ( .A(n4681), .B(n4514), .Z(n4515) );
  XNOR U6418 ( .A(n4940), .B(n4515), .Z(out[820]) );
  XOR U6419 ( .A(in[732]), .B(n4516), .Z(n4944) );
  NANDN U6420 ( .A(n4682), .B(n4517), .Z(n4518) );
  XNOR U6421 ( .A(n4944), .B(n4518), .Z(out[821]) );
  XOR U6422 ( .A(in[733]), .B(n4519), .Z(n4952) );
  NANDN U6423 ( .A(n4683), .B(n4520), .Z(n4521) );
  XNOR U6424 ( .A(n4952), .B(n4521), .Z(out[822]) );
  XNOR U6425 ( .A(in[734]), .B(n4522), .Z(n4956) );
  IV U6426 ( .A(n4523), .Z(n4684) );
  NANDN U6427 ( .A(n4524), .B(n4684), .Z(n4525) );
  XNOR U6428 ( .A(n4956), .B(n4525), .Z(out[823]) );
  XNOR U6429 ( .A(in[735]), .B(n4526), .Z(n4960) );
  IV U6430 ( .A(n4527), .Z(n4686) );
  NANDN U6431 ( .A(n4528), .B(n4686), .Z(n4529) );
  XNOR U6432 ( .A(n4960), .B(n4529), .Z(out[824]) );
  XNOR U6433 ( .A(in[736]), .B(n4530), .Z(n4964) );
  IV U6434 ( .A(n4531), .Z(n4688) );
  NANDN U6435 ( .A(n4532), .B(n4688), .Z(n4533) );
  XNOR U6436 ( .A(n4964), .B(n4533), .Z(out[825]) );
  XNOR U6437 ( .A(in[737]), .B(n4534), .Z(n4968) );
  IV U6438 ( .A(n4535), .Z(n4693) );
  NANDN U6439 ( .A(n4536), .B(n4693), .Z(n4537) );
  XNOR U6440 ( .A(n4968), .B(n4537), .Z(out[826]) );
  XNOR U6441 ( .A(in[738]), .B(n4538), .Z(n4972) );
  IV U6442 ( .A(n4539), .Z(n4695) );
  NANDN U6443 ( .A(n4540), .B(n4695), .Z(n4541) );
  XNOR U6444 ( .A(n4972), .B(n4541), .Z(out[827]) );
  XNOR U6445 ( .A(in[739]), .B(n4542), .Z(n4976) );
  IV U6446 ( .A(n4543), .Z(n4697) );
  NANDN U6447 ( .A(n4544), .B(n4697), .Z(n4545) );
  XNOR U6448 ( .A(n4976), .B(n4545), .Z(out[828]) );
  XOR U6449 ( .A(in[740]), .B(n4546), .Z(n4700) );
  IV U6450 ( .A(n4700), .Z(n4980) );
  ANDN U6451 ( .B(n4549), .A(n4548), .Z(n4550) );
  XOR U6452 ( .A(n4551), .B(n4550), .Z(out[82]) );
  XOR U6453 ( .A(in[741]), .B(n4552), .Z(n4703) );
  IV U6454 ( .A(n4703), .Z(n4984) );
  XOR U6455 ( .A(in[742]), .B(n4554), .Z(n4706) );
  IV U6456 ( .A(n4706), .Z(n4988) );
  NANDN U6457 ( .A(n4557), .B(n4556), .Z(n4558) );
  XOR U6458 ( .A(n4709), .B(n4558), .Z(out[832]) );
  NANDN U6459 ( .A(n4560), .B(n4559), .Z(n4561) );
  XOR U6460 ( .A(n4713), .B(n4561), .Z(out[833]) );
  NANDN U6461 ( .A(n4563), .B(n4562), .Z(n4564) );
  XOR U6462 ( .A(n4717), .B(n4564), .Z(out[834]) );
  NANDN U6463 ( .A(n4566), .B(n4565), .Z(n4567) );
  XOR U6464 ( .A(n4721), .B(n4567), .Z(out[835]) );
  NANDN U6465 ( .A(n4568), .B(n4732), .Z(n4569) );
  XOR U6466 ( .A(n4733), .B(n4569), .Z(out[836]) );
  NANDN U6467 ( .A(n4570), .B(n4736), .Z(n4571) );
  XOR U6468 ( .A(n4737), .B(n4571), .Z(out[837]) );
  NANDN U6469 ( .A(n4572), .B(n4740), .Z(n4573) );
  XOR U6470 ( .A(n4741), .B(n4573), .Z(out[838]) );
  NANDN U6471 ( .A(n4575), .B(n4574), .Z(n4576) );
  XOR U6472 ( .A(n4745), .B(n4576), .Z(out[839]) );
  ANDN U6473 ( .B(n4578), .A(n4577), .Z(n4579) );
  XOR U6474 ( .A(n4580), .B(n4579), .Z(out[83]) );
  NANDN U6475 ( .A(n4581), .B(n4749), .Z(n4582) );
  XNOR U6476 ( .A(n4748), .B(n4582), .Z(out[840]) );
  NANDN U6477 ( .A(n4583), .B(n4753), .Z(n4584) );
  XNOR U6478 ( .A(n4752), .B(n4584), .Z(out[841]) );
  NANDN U6479 ( .A(n4585), .B(n4757), .Z(n4586) );
  XNOR U6480 ( .A(n4756), .B(n4586), .Z(out[842]) );
  NANDN U6481 ( .A(n4587), .B(n4761), .Z(n4588) );
  XNOR U6482 ( .A(n4760), .B(n4588), .Z(out[843]) );
  NANDN U6483 ( .A(n4589), .B(n4765), .Z(n4590) );
  XNOR U6484 ( .A(n4764), .B(n4590), .Z(out[844]) );
  NANDN U6485 ( .A(n4591), .B(n4769), .Z(n4592) );
  XNOR U6486 ( .A(n4768), .B(n4592), .Z(out[845]) );
  NANDN U6487 ( .A(n4593), .B(n4777), .Z(n4594) );
  XNOR U6488 ( .A(n4776), .B(n4594), .Z(out[846]) );
  NANDN U6489 ( .A(n4595), .B(n4781), .Z(n4596) );
  XNOR U6490 ( .A(n4780), .B(n4596), .Z(out[847]) );
  NANDN U6491 ( .A(n4598), .B(n4597), .Z(n4599) );
  XNOR U6492 ( .A(n4784), .B(n4599), .Z(out[848]) );
  NANDN U6493 ( .A(n4600), .B(n4789), .Z(n4601) );
  XNOR U6494 ( .A(n4788), .B(n4601), .Z(out[849]) );
  ANDN U6495 ( .B(n4603), .A(n4602), .Z(n4604) );
  XOR U6496 ( .A(n4605), .B(n4604), .Z(out[84]) );
  NANDN U6497 ( .A(n4606), .B(n4793), .Z(n4607) );
  XNOR U6498 ( .A(n4792), .B(n4607), .Z(out[850]) );
  NANDN U6499 ( .A(n4608), .B(n4797), .Z(n4609) );
  XNOR U6500 ( .A(n4796), .B(n4609), .Z(out[851]) );
  NANDN U6501 ( .A(n4610), .B(n4801), .Z(n4611) );
  XNOR U6502 ( .A(n4800), .B(n4611), .Z(out[852]) );
  NANDN U6503 ( .A(n4612), .B(n4805), .Z(n4613) );
  XNOR U6504 ( .A(n4804), .B(n4613), .Z(out[853]) );
  NANDN U6505 ( .A(n4615), .B(n4614), .Z(n4616) );
  XNOR U6506 ( .A(n4808), .B(n4616), .Z(out[854]) );
  NANDN U6507 ( .A(n4618), .B(n4617), .Z(n4619) );
  XNOR U6508 ( .A(n4812), .B(n4619), .Z(out[855]) );
  NANDN U6509 ( .A(n4621), .B(n4620), .Z(n4622) );
  XNOR U6510 ( .A(n4820), .B(n4622), .Z(out[856]) );
  NANDN U6511 ( .A(n4624), .B(n4623), .Z(n4625) );
  XNOR U6512 ( .A(n4824), .B(n4625), .Z(out[857]) );
  NANDN U6513 ( .A(n4626), .B(n4829), .Z(n4627) );
  XNOR U6514 ( .A(n4828), .B(n4627), .Z(out[858]) );
  NANDN U6515 ( .A(n4628), .B(n4833), .Z(n4629) );
  XNOR U6516 ( .A(n4832), .B(n4629), .Z(out[859]) );
  NANDN U6517 ( .A(n4634), .B(n4633), .Z(n4635) );
  XNOR U6518 ( .A(n4836), .B(n4635), .Z(out[860]) );
  NANDN U6519 ( .A(n4637), .B(n4636), .Z(n4638) );
  XNOR U6520 ( .A(n4840), .B(n4638), .Z(out[861]) );
  NANDN U6521 ( .A(n4640), .B(n4639), .Z(n4641) );
  XNOR U6522 ( .A(n4844), .B(n4641), .Z(out[862]) );
  NANDN U6523 ( .A(n4644), .B(n4643), .Z(n4645) );
  XNOR U6524 ( .A(n4852), .B(n4645), .Z(out[864]) );
  NANDN U6525 ( .A(n4647), .B(n4646), .Z(n4648) );
  XNOR U6526 ( .A(n4856), .B(n4648), .Z(out[865]) );
  NANDN U6527 ( .A(n4650), .B(n4649), .Z(n4651) );
  XNOR U6528 ( .A(n4864), .B(n4651), .Z(out[866]) );
  NANDN U6529 ( .A(n4653), .B(n4652), .Z(n4654) );
  XNOR U6530 ( .A(n4868), .B(n4654), .Z(out[867]) );
  NANDN U6531 ( .A(n4656), .B(n4655), .Z(n4657) );
  XNOR U6532 ( .A(n4872), .B(n4657), .Z(out[868]) );
  ANDN U6533 ( .B(n4660), .A(n4659), .Z(n4661) );
  XOR U6534 ( .A(n4662), .B(n4661), .Z(out[86]) );
  OR U6535 ( .A(n4901), .B(n4668), .Z(n4669) );
  XNOR U6536 ( .A(n4900), .B(n4669), .Z(out[875]) );
  OR U6537 ( .A(n4956), .B(n4684), .Z(n4685) );
  XOR U6538 ( .A(n4957), .B(n4685), .Z(out[887]) );
  OR U6539 ( .A(n4960), .B(n4686), .Z(n4687) );
  XOR U6540 ( .A(n4961), .B(n4687), .Z(out[888]) );
  OR U6541 ( .A(n4964), .B(n4688), .Z(n4689) );
  XOR U6542 ( .A(n4965), .B(n4689), .Z(out[889]) );
  OR U6543 ( .A(n4968), .B(n4693), .Z(n4694) );
  XOR U6544 ( .A(n4969), .B(n4694), .Z(out[890]) );
  OR U6545 ( .A(n4972), .B(n4695), .Z(n4696) );
  XOR U6546 ( .A(n4973), .B(n4696), .Z(out[891]) );
  OR U6547 ( .A(n4976), .B(n4697), .Z(n4698) );
  XOR U6548 ( .A(n4977), .B(n4698), .Z(out[892]) );
  NANDN U6549 ( .A(n4700), .B(n4699), .Z(n4701) );
  XOR U6550 ( .A(n4981), .B(n4701), .Z(out[893]) );
  NANDN U6551 ( .A(n4703), .B(n4702), .Z(n4704) );
  XOR U6552 ( .A(n4985), .B(n4704), .Z(out[894]) );
  NANDN U6553 ( .A(n4706), .B(n4705), .Z(n4707) );
  XOR U6554 ( .A(n4989), .B(n4707), .Z(out[895]) );
  ANDN U6555 ( .B(n4709), .A(n4708), .Z(n4710) );
  XOR U6556 ( .A(n4711), .B(n4710), .Z(out[896]) );
  ANDN U6557 ( .B(n4713), .A(n4712), .Z(n4714) );
  XOR U6558 ( .A(n4715), .B(n4714), .Z(out[897]) );
  ANDN U6559 ( .B(n4717), .A(n4716), .Z(n4718) );
  XOR U6560 ( .A(n4719), .B(n4718), .Z(out[898]) );
  ANDN U6561 ( .B(n4721), .A(n4720), .Z(n4722) );
  XOR U6562 ( .A(n4723), .B(n4722), .Z(out[899]) );
  ANDN U6563 ( .B(n4725), .A(n4724), .Z(n4726) );
  XOR U6564 ( .A(n4727), .B(n4726), .Z(out[89]) );
  OR U6565 ( .A(n4729), .B(n4728), .Z(n4730) );
  XNOR U6566 ( .A(n4731), .B(n4730), .Z(out[8]) );
  ANDN U6567 ( .B(n4733), .A(n4732), .Z(n4734) );
  XOR U6568 ( .A(n4735), .B(n4734), .Z(out[900]) );
  ANDN U6569 ( .B(n4737), .A(n4736), .Z(n4738) );
  XOR U6570 ( .A(n4739), .B(n4738), .Z(out[901]) );
  ANDN U6571 ( .B(n4741), .A(n4740), .Z(n4742) );
  XOR U6572 ( .A(n4743), .B(n4742), .Z(out[902]) );
  ANDN U6573 ( .B(n4745), .A(n4744), .Z(n4746) );
  XOR U6574 ( .A(n4747), .B(n4746), .Z(out[903]) );
  NOR U6575 ( .A(n4749), .B(n4748), .Z(n4750) );
  XOR U6576 ( .A(n4751), .B(n4750), .Z(out[904]) );
  NOR U6577 ( .A(n4753), .B(n4752), .Z(n4754) );
  XOR U6578 ( .A(n4755), .B(n4754), .Z(out[905]) );
  NOR U6579 ( .A(n4757), .B(n4756), .Z(n4758) );
  XOR U6580 ( .A(n4759), .B(n4758), .Z(out[906]) );
  NOR U6581 ( .A(n4761), .B(n4760), .Z(n4762) );
  XOR U6582 ( .A(n4763), .B(n4762), .Z(out[907]) );
  NOR U6583 ( .A(n4765), .B(n4764), .Z(n4766) );
  XOR U6584 ( .A(n4767), .B(n4766), .Z(out[908]) );
  NOR U6585 ( .A(n4769), .B(n4768), .Z(n4770) );
  XOR U6586 ( .A(n4771), .B(n4770), .Z(out[909]) );
  ANDN U6587 ( .B(n4773), .A(n4772), .Z(n4774) );
  XOR U6588 ( .A(n4775), .B(n4774), .Z(out[90]) );
  NOR U6589 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U6590 ( .A(n4779), .B(n4778), .Z(out[910]) );
  NOR U6591 ( .A(n4781), .B(n4780), .Z(n4782) );
  XOR U6592 ( .A(n4783), .B(n4782), .Z(out[911]) );
  NOR U6593 ( .A(n4785), .B(n4784), .Z(n4786) );
  XOR U6594 ( .A(n4787), .B(n4786), .Z(out[912]) );
  NOR U6595 ( .A(n4789), .B(n4788), .Z(n4790) );
  XOR U6596 ( .A(n4791), .B(n4790), .Z(out[913]) );
  NOR U6597 ( .A(n4793), .B(n4792), .Z(n4794) );
  XOR U6598 ( .A(n4795), .B(n4794), .Z(out[914]) );
  NOR U6599 ( .A(n4797), .B(n4796), .Z(n4798) );
  XOR U6600 ( .A(n4799), .B(n4798), .Z(out[915]) );
  NOR U6601 ( .A(n4801), .B(n4800), .Z(n4802) );
  XOR U6602 ( .A(n4803), .B(n4802), .Z(out[916]) );
  NOR U6603 ( .A(n4805), .B(n4804), .Z(n4806) );
  XOR U6604 ( .A(n4807), .B(n4806), .Z(out[917]) );
  NOR U6605 ( .A(n4809), .B(n4808), .Z(n4810) );
  XOR U6606 ( .A(n4811), .B(n4810), .Z(out[918]) );
  NOR U6607 ( .A(n4813), .B(n4812), .Z(n4814) );
  XOR U6608 ( .A(n4815), .B(n4814), .Z(out[919]) );
  ANDN U6609 ( .B(n4817), .A(n4816), .Z(n4818) );
  XOR U6610 ( .A(n4819), .B(n4818), .Z(out[91]) );
  NOR U6611 ( .A(n4821), .B(n4820), .Z(n4822) );
  XOR U6612 ( .A(n4823), .B(n4822), .Z(out[920]) );
  NOR U6613 ( .A(n4825), .B(n4824), .Z(n4826) );
  XOR U6614 ( .A(n4827), .B(n4826), .Z(out[921]) );
  NOR U6615 ( .A(n4829), .B(n4828), .Z(n4830) );
  XOR U6616 ( .A(n4831), .B(n4830), .Z(out[922]) );
  NOR U6617 ( .A(n4833), .B(n4832), .Z(n4834) );
  XOR U6618 ( .A(n4835), .B(n4834), .Z(out[923]) );
  NOR U6619 ( .A(n4837), .B(n4836), .Z(n4838) );
  XOR U6620 ( .A(n4839), .B(n4838), .Z(out[924]) );
  NOR U6621 ( .A(n4841), .B(n4840), .Z(n4842) );
  XOR U6622 ( .A(n4843), .B(n4842), .Z(out[925]) );
  NOR U6623 ( .A(n4845), .B(n4844), .Z(n4846) );
  XOR U6624 ( .A(n4847), .B(n4846), .Z(out[926]) );
  NOR U6625 ( .A(n4849), .B(n4848), .Z(n4850) );
  XOR U6626 ( .A(n4851), .B(n4850), .Z(out[927]) );
  NOR U6627 ( .A(n4853), .B(n4852), .Z(n4854) );
  XOR U6628 ( .A(n4855), .B(n4854), .Z(out[928]) );
  NOR U6629 ( .A(n4857), .B(n4856), .Z(n4858) );
  XOR U6630 ( .A(n4859), .B(n4858), .Z(out[929]) );
  AND U6631 ( .A(n4861), .B(n4860), .Z(n4862) );
  XNOR U6632 ( .A(n4863), .B(n4862), .Z(out[92]) );
  NOR U6633 ( .A(n4865), .B(n4864), .Z(n4866) );
  XOR U6634 ( .A(n4867), .B(n4866), .Z(out[930]) );
  NOR U6635 ( .A(n4869), .B(n4868), .Z(n4870) );
  XOR U6636 ( .A(n4871), .B(n4870), .Z(out[931]) );
  NOR U6637 ( .A(n4873), .B(n4872), .Z(n4874) );
  XOR U6638 ( .A(n4875), .B(n4874), .Z(out[932]) );
  ANDN U6639 ( .B(n4877), .A(n4876), .Z(n4878) );
  XOR U6640 ( .A(n4879), .B(n4878), .Z(out[933]) );
  ANDN U6641 ( .B(n4881), .A(n4880), .Z(n4882) );
  XOR U6642 ( .A(n4883), .B(n4882), .Z(out[934]) );
  ANDN U6643 ( .B(n4885), .A(n4884), .Z(n4886) );
  XOR U6644 ( .A(n4887), .B(n4886), .Z(out[935]) );
  ANDN U6645 ( .B(n4889), .A(n4888), .Z(n4890) );
  XOR U6646 ( .A(n4891), .B(n4890), .Z(out[936]) );
  ANDN U6647 ( .B(n4893), .A(n4892), .Z(n4894) );
  XOR U6648 ( .A(n4895), .B(n4894), .Z(out[937]) );
  ANDN U6649 ( .B(n4897), .A(n4896), .Z(n4898) );
  XOR U6650 ( .A(n4899), .B(n4898), .Z(out[938]) );
  ANDN U6651 ( .B(n4901), .A(n4900), .Z(n4902) );
  XOR U6652 ( .A(n4903), .B(n4902), .Z(out[939]) );
  AND U6653 ( .A(n4905), .B(n4904), .Z(n4906) );
  XNOR U6654 ( .A(n4907), .B(n4906), .Z(out[93]) );
  AND U6655 ( .A(n4909), .B(n4908), .Z(n4910) );
  XNOR U6656 ( .A(n4911), .B(n4910), .Z(out[940]) );
  AND U6657 ( .A(n4913), .B(n4912), .Z(n4914) );
  XNOR U6658 ( .A(n4915), .B(n4914), .Z(out[941]) );
  AND U6659 ( .A(n4917), .B(n4916), .Z(n4918) );
  XNOR U6660 ( .A(n4919), .B(n4918), .Z(out[942]) );
  AND U6661 ( .A(n4921), .B(n4920), .Z(n4922) );
  XNOR U6662 ( .A(n4923), .B(n4922), .Z(out[943]) );
  AND U6663 ( .A(n4925), .B(n4924), .Z(n4926) );
  XNOR U6664 ( .A(n4927), .B(n4926), .Z(out[944]) );
  AND U6665 ( .A(n4929), .B(n4928), .Z(n4930) );
  XNOR U6666 ( .A(n4931), .B(n4930), .Z(out[945]) );
  AND U6667 ( .A(n4933), .B(n4932), .Z(n4934) );
  XNOR U6668 ( .A(n4935), .B(n4934), .Z(out[946]) );
  AND U6669 ( .A(n4937), .B(n4936), .Z(n4938) );
  XNOR U6670 ( .A(n4939), .B(n4938), .Z(out[947]) );
  AND U6671 ( .A(n4941), .B(n4940), .Z(n4942) );
  XNOR U6672 ( .A(n4943), .B(n4942), .Z(out[948]) );
  AND U6673 ( .A(n4945), .B(n4944), .Z(n4946) );
  XNOR U6674 ( .A(n4947), .B(n4946), .Z(out[949]) );
  AND U6675 ( .A(n4949), .B(n4948), .Z(n4950) );
  XNOR U6676 ( .A(n4951), .B(n4950), .Z(out[94]) );
  AND U6677 ( .A(n4953), .B(n4952), .Z(n4954) );
  XNOR U6678 ( .A(n4955), .B(n4954), .Z(out[950]) );
  AND U6679 ( .A(n4957), .B(n4956), .Z(n4958) );
  XNOR U6680 ( .A(n4959), .B(n4958), .Z(out[951]) );
  AND U6681 ( .A(n4961), .B(n4960), .Z(n4962) );
  XNOR U6682 ( .A(n4963), .B(n4962), .Z(out[952]) );
  AND U6683 ( .A(n4965), .B(n4964), .Z(n4966) );
  XNOR U6684 ( .A(n4967), .B(n4966), .Z(out[953]) );
  AND U6685 ( .A(n4969), .B(n4968), .Z(n4970) );
  XNOR U6686 ( .A(n4971), .B(n4970), .Z(out[954]) );
  AND U6687 ( .A(n4973), .B(n4972), .Z(n4974) );
  XNOR U6688 ( .A(n4975), .B(n4974), .Z(out[955]) );
  AND U6689 ( .A(n4977), .B(n4976), .Z(n4978) );
  XOR U6690 ( .A(n4979), .B(n4978), .Z(out[956]) );
  ANDN U6691 ( .B(n4981), .A(n4980), .Z(n4982) );
  XOR U6692 ( .A(n4983), .B(n4982), .Z(out[957]) );
  ANDN U6693 ( .B(n4985), .A(n4984), .Z(n4986) );
  XOR U6694 ( .A(n4987), .B(n4986), .Z(out[958]) );
  ANDN U6695 ( .B(n4989), .A(n4988), .Z(n4990) );
  XNOR U6696 ( .A(n4991), .B(n4990), .Z(out[959]) );
  AND U6697 ( .A(n4993), .B(n4992), .Z(n4994) );
  XNOR U6698 ( .A(n4995), .B(n4994), .Z(out[95]) );
  ANDN U6699 ( .B(n4997), .A(n4996), .Z(n4998) );
  XOR U6700 ( .A(n4999), .B(n4998), .Z(out[960]) );
  ANDN U6701 ( .B(n5001), .A(n5000), .Z(n5002) );
  XOR U6702 ( .A(n5003), .B(n5002), .Z(out[961]) );
  ANDN U6703 ( .B(n5005), .A(n5004), .Z(n5006) );
  XOR U6704 ( .A(n5007), .B(n5006), .Z(out[962]) );
  ANDN U6705 ( .B(n5009), .A(n5008), .Z(n5010) );
  XOR U6706 ( .A(n5011), .B(n5010), .Z(out[963]) );
  ANDN U6707 ( .B(n5013), .A(n5012), .Z(n5014) );
  XOR U6708 ( .A(n5015), .B(n5014), .Z(out[964]) );
  ANDN U6709 ( .B(n5017), .A(n5016), .Z(n5018) );
  XOR U6710 ( .A(n5019), .B(n5018), .Z(out[965]) );
  ANDN U6711 ( .B(n5021), .A(n5020), .Z(n5022) );
  XOR U6712 ( .A(n5023), .B(n5022), .Z(out[966]) );
  ANDN U6713 ( .B(n5025), .A(n5024), .Z(n5026) );
  XOR U6714 ( .A(n5027), .B(n5026), .Z(out[967]) );
  ANDN U6715 ( .B(n5029), .A(n5028), .Z(n5030) );
  XOR U6716 ( .A(n5031), .B(n5030), .Z(out[968]) );
  ANDN U6717 ( .B(n5033), .A(n5032), .Z(n5034) );
  XOR U6718 ( .A(n5035), .B(n5034), .Z(out[969]) );
  AND U6719 ( .A(n5037), .B(n5036), .Z(n5038) );
  XNOR U6720 ( .A(n5039), .B(n5038), .Z(out[96]) );
  ANDN U6721 ( .B(n5041), .A(n5040), .Z(n5042) );
  XOR U6722 ( .A(n5043), .B(n5042), .Z(out[970]) );
  ANDN U6723 ( .B(n5045), .A(n5044), .Z(n5046) );
  XOR U6724 ( .A(n5047), .B(n5046), .Z(out[971]) );
  ANDN U6725 ( .B(n5049), .A(n5048), .Z(n5050) );
  XOR U6726 ( .A(n5051), .B(n5050), .Z(out[972]) );
  ANDN U6727 ( .B(n5053), .A(n5052), .Z(n5054) );
  XOR U6728 ( .A(n5055), .B(n5054), .Z(out[973]) );
  ANDN U6729 ( .B(n5057), .A(n5056), .Z(n5058) );
  XOR U6730 ( .A(n5059), .B(n5058), .Z(out[974]) );
  ANDN U6731 ( .B(n5061), .A(n5060), .Z(n5062) );
  XOR U6732 ( .A(n5063), .B(n5062), .Z(out[975]) );
  ANDN U6733 ( .B(n5074), .A(n5073), .Z(n5075) );
  XOR U6734 ( .A(n5076), .B(n5075), .Z(out[979]) );
  AND U6735 ( .A(n5078), .B(n5077), .Z(n5079) );
  XNOR U6736 ( .A(n5080), .B(n5079), .Z(out[97]) );
  ANDN U6737 ( .B(n5106), .A(n5105), .Z(n5107) );
  XOR U6738 ( .A(n5108), .B(n5107), .Z(out[988]) );
  ANDN U6739 ( .B(n5113), .A(n5112), .Z(n5114) );
  XNOR U6740 ( .A(n5115), .B(n5114), .Z(out[98]) );
  ANDN U6741 ( .B(n5120), .A(n5119), .Z(n5121) );
  XOR U6742 ( .A(n5122), .B(n5121), .Z(out[991]) );
  ANDN U6743 ( .B(n5124), .A(n5123), .Z(n5125) );
  XOR U6744 ( .A(n5126), .B(n5125), .Z(out[992]) );
  ANDN U6745 ( .B(n5128), .A(n5127), .Z(n5129) );
  XOR U6746 ( .A(n5130), .B(n5129), .Z(out[993]) );
  ANDN U6747 ( .B(n5132), .A(n5131), .Z(n5133) );
  XOR U6748 ( .A(n5134), .B(n5133), .Z(out[994]) );
  ANDN U6749 ( .B(n5136), .A(n5135), .Z(n5137) );
  XNOR U6750 ( .A(n5138), .B(n5137), .Z(out[995]) );
  ANDN U6751 ( .B(n5140), .A(n5139), .Z(n5141) );
  XNOR U6752 ( .A(n5142), .B(n5141), .Z(out[996]) );
  ANDN U6753 ( .B(n5144), .A(n5143), .Z(n5145) );
  XNOR U6754 ( .A(n5146), .B(n5145), .Z(out[997]) );
  AND U6755 ( .A(n5148), .B(n5147), .Z(n5149) );
  XNOR U6756 ( .A(n5150), .B(n5149), .Z(out[998]) );
  ANDN U6757 ( .B(n5152), .A(n5151), .Z(n5153) );
  XNOR U6758 ( .A(n5154), .B(n5153), .Z(out[999]) );
  ANDN U6759 ( .B(n5156), .A(n5155), .Z(n5157) );
  XNOR U6760 ( .A(n5158), .B(n5157), .Z(out[99]) );
  OR U6761 ( .A(n5160), .B(n5159), .Z(n5161) );
  XNOR U6762 ( .A(n5162), .B(n5161), .Z(out[9]) );
endmodule


module round_3 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_3, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_3 = round_const[3];

  XNOR U1 ( .A(n1413), .B(n1697), .Z(n3185) );
  XNOR U2 ( .A(n1418), .B(n1701), .Z(n3187) );
  XNOR U3 ( .A(n1425), .B(n1719), .Z(n3198) );
  XNOR U4 ( .A(n1431), .B(n1731), .Z(n3206) );
  XNOR U5 ( .A(n1449), .B(n1030), .Z(n2782) );
  XNOR U6 ( .A(n1461), .B(n1084), .Z(n2866) );
  XOR U7 ( .A(n1422), .B(n1380), .Z(n4464) );
  XOR U8 ( .A(n1384), .B(n1424), .Z(n4467) );
  XOR U9 ( .A(n1388), .B(n1426), .Z(n4470) );
  XOR U10 ( .A(n1392), .B(n1428), .Z(n4473) );
  XOR U11 ( .A(n1396), .B(n1430), .Z(n4476) );
  XOR U12 ( .A(n1442), .B(n760), .Z(n4495) );
  XOR U13 ( .A(n775), .B(n1444), .Z(n4498) );
  XOR U14 ( .A(n1446), .B(n790), .Z(n4501) );
  XOR U15 ( .A(n1448), .B(n816), .Z(n4504) );
  XOR U16 ( .A(n1450), .B(n831), .Z(n4507) );
  XOR U17 ( .A(n1454), .B(n846), .Z(n4510) );
  NANDN U18 ( .A(n2853), .B(n3855), .Z(n1) );
  XNOR U19 ( .A(n3020), .B(n1), .Z(out[190]) );
  NANDN U20 ( .A(n2885), .B(n2884), .Z(n2) );
  XNOR U21 ( .A(n4312), .B(n2), .Z(out[267]) );
  NANDN U22 ( .A(n3448), .B(n3875), .Z(n3) );
  XNOR U23 ( .A(n3604), .B(n3), .Z(out[442]) );
  NANDN U24 ( .A(n3451), .B(n3879), .Z(n4) );
  XNOR U25 ( .A(n3605), .B(n4), .Z(out[443]) );
  XNOR U26 ( .A(n1445), .B(n1004), .Z(n2758) );
  XNOR U27 ( .A(n1443), .B(n1752), .Z(n3220) );
  XNOR U28 ( .A(n1405), .B(n1681), .Z(n3177) );
  XNOR U29 ( .A(n1409), .B(n1689), .Z(n3181) );
  XNOR U30 ( .A(n1433), .B(n1735), .Z(n3209) );
  XNOR U31 ( .A(n1467), .B(n1097), .Z(n2890) );
  XNOR U32 ( .A(n1471), .B(n1117), .Z(n2923) );
  XNOR U33 ( .A(n1496), .B(n1231), .Z(n2215) );
  XNOR U34 ( .A(n1477), .B(n1143), .Z(n4060) );
  XNOR U35 ( .A(n1480), .B(n1156), .Z(n4064) );
  XNOR U36 ( .A(n1676), .B(n1677), .Z(n3075) );
  XNOR U37 ( .A(n1696), .B(n1697), .Z(n3087) );
  XNOR U38 ( .A(n1710), .B(n1711), .Z(n3092) );
  XNOR U39 ( .A(n1718), .B(n1719), .Z(n3096) );
  XNOR U40 ( .A(n1722), .B(n1723), .Z(n3098) );
  XNOR U41 ( .A(n1726), .B(n1727), .Z(n3102) );
  XOR U42 ( .A(n1400), .B(n1432), .Z(n4483) );
  XOR U43 ( .A(n730), .B(n1436), .Z(n4489) );
  XOR U44 ( .A(n745), .B(n1440), .Z(n4492) );
  XNOR U45 ( .A(n1458), .B(n876), .Z(n4520) );
  XOR U46 ( .A(n1472), .B(n921), .Z(n4530) );
  XOR U47 ( .A(n1476), .B(n936), .Z(n4534) );
  XOR U48 ( .A(n698), .B(n1481), .Z(n4542) );
  XNOR U49 ( .A(n3944), .B(in[1481]), .Z(n4766) );
  NAND U50 ( .A(n3941), .B(n3940), .Z(n5) );
  XNOR U51 ( .A(n3942), .B(n5), .Z(out[64]) );
  AND U52 ( .A(n4698), .B(n4697), .Z(n6) );
  XNOR U53 ( .A(n4699), .B(n6), .Z(out[88]) );
  NANDN U54 ( .A(n2851), .B(n3811), .Z(n7) );
  XNOR U55 ( .A(n3019), .B(n7), .Z(out[189]) );
  NAND U56 ( .A(n2894), .B(n4410), .Z(n8) );
  XNOR U57 ( .A(n2893), .B(n8), .Z(out[206]) );
  NAND U58 ( .A(n2897), .B(n4444), .Z(n9) );
  XNOR U59 ( .A(n2896), .B(n9), .Z(out[207]) );
  NAND U60 ( .A(n2900), .B(n4482), .Z(n10) );
  XNOR U61 ( .A(n2899), .B(n10), .Z(out[208]) );
  NAND U62 ( .A(n2903), .B(n4516), .Z(n11) );
  XNOR U63 ( .A(n2902), .B(n11), .Z(out[209]) );
  NANDN U64 ( .A(n2887), .B(n2886), .Z(n12) );
  XNOR U65 ( .A(n4344), .B(n12), .Z(out[268]) );
  NANDN U66 ( .A(n2889), .B(n2888), .Z(n13) );
  XNOR U67 ( .A(n4375), .B(n13), .Z(out[269]) );
  NANDN U68 ( .A(n3280), .B(n3637), .Z(n14) );
  XNOR U69 ( .A(n3477), .B(n14), .Z(out[388]) );
  NANDN U70 ( .A(n3283), .B(n3641), .Z(n15) );
  XNOR U71 ( .A(n3478), .B(n15), .Z(out[389]) );
  NANDN U72 ( .A(n3286), .B(n3645), .Z(n16) );
  XNOR U73 ( .A(n3479), .B(n16), .Z(out[390]) );
  NANDN U74 ( .A(n3289), .B(n3649), .Z(n17) );
  XNOR U75 ( .A(n3480), .B(n17), .Z(out[391]) );
  NANDN U76 ( .A(n3292), .B(n3653), .Z(n18) );
  XNOR U77 ( .A(n3485), .B(n18), .Z(out[392]) );
  NAND U78 ( .A(n3839), .B(n3419), .Z(n19) );
  XNOR U79 ( .A(n3418), .B(n19), .Z(out[434]) );
  NAND U80 ( .A(n3843), .B(n3422), .Z(n20) );
  XNOR U81 ( .A(n3421), .B(n20), .Z(out[435]) );
  ANDN U82 ( .B(n3859), .A(n3436), .Z(n21) );
  XNOR U83 ( .A(n3592), .B(n21), .Z(out[438]) );
  ANDN U84 ( .B(n3863), .A(n3439), .Z(n22) );
  XNOR U85 ( .A(n3594), .B(n22), .Z(out[439]) );
  ANDN U86 ( .B(n3871), .A(n3445), .Z(n23) );
  XNOR U87 ( .A(n3598), .B(n23), .Z(out[441]) );
  ANDN U88 ( .B(n3887), .A(n3457), .Z(n24) );
  XNOR U89 ( .A(n3608), .B(n24), .Z(out[445]) );
  ANDN U90 ( .B(n3895), .A(n3467), .Z(n25) );
  XNOR U91 ( .A(n3612), .B(n25), .Z(out[447]) );
  NAND U92 ( .A(n3604), .B(n3873), .Z(n26) );
  XNOR U93 ( .A(n3872), .B(n26), .Z(out[570]) );
  NAND U94 ( .A(n3605), .B(n3877), .Z(n27) );
  XNOR U95 ( .A(n3876), .B(n27), .Z(out[571]) );
  XNOR U96 ( .A(n1441), .B(n1748), .Z(n3217) );
  XNOR U97 ( .A(n1401), .B(n1677), .Z(n3175) );
  XNOR U98 ( .A(n1706), .B(n1346), .Z(n3933) );
  XNOR U99 ( .A(n1411), .B(n1693), .Z(n3183) );
  XNOR U100 ( .A(n1427), .B(n1723), .Z(n3200) );
  XNOR U101 ( .A(n1435), .B(n1739), .Z(n3212) );
  XNOR U102 ( .A(n1447), .B(n1017), .Z(n2775) );
  XNOR U103 ( .A(n1453), .B(n1043), .Z(n2796) );
  XNOR U104 ( .A(n1455), .B(n1056), .Z(n2819) );
  XNOR U105 ( .A(n1457), .B(n1069), .Z(n2842) );
  XNOR U106 ( .A(n1475), .B(n1130), .Z(n4056) );
  XNOR U107 ( .A(n1655), .B(n1656), .Z(n3063) );
  XNOR U108 ( .A(n1486), .B(n1186), .Z(n4076) );
  XNOR U109 ( .A(n1672), .B(n1673), .Z(n3072) );
  XNOR U110 ( .A(n1680), .B(n1681), .Z(n3077) );
  XNOR U111 ( .A(n1684), .B(n1685), .Z(n3081) );
  XNOR U112 ( .A(n1688), .B(n1689), .Z(n3083) );
  XOR U113 ( .A(n1714), .B(n1715), .Z(n3094) );
  XNOR U114 ( .A(n1730), .B(n1731), .Z(n3104) );
  XNOR U115 ( .A(n1439), .B(n1743), .Z(n4004) );
  XOR U116 ( .A(n715), .B(n1434), .Z(n4486) );
  XNOR U117 ( .A(n1456), .B(n861), .Z(n4517) );
  XNOR U118 ( .A(n1462), .B(n891), .Z(n4523) );
  XOR U119 ( .A(n1468), .B(n906), .Z(n4526) );
  XOR U120 ( .A(n1478), .B(n681), .Z(n4538) );
  XOR U121 ( .A(n809), .B(n1484), .Z(n4546) );
  XNOR U122 ( .A(n3937), .B(in[1480]), .Z(n4762) );
  XNOR U123 ( .A(n3948), .B(in[1482]), .Z(n4770) );
  XNOR U124 ( .A(n3952), .B(in[1483]), .Z(n4774) );
  XNOR U125 ( .A(n3956), .B(in[1484]), .Z(n4778) );
  NANDN U126 ( .A(n3984), .B(n3983), .Z(n28) );
  XNOR U127 ( .A(n3985), .B(n28), .Z(out[65]) );
  AND U128 ( .A(n4780), .B(n4779), .Z(n29) );
  XNOR U129 ( .A(n4781), .B(n29), .Z(out[90]) );
  AND U130 ( .A(n4823), .B(n4822), .Z(n30) );
  XNOR U131 ( .A(n4824), .B(n30), .Z(out[91]) );
  NAND U132 ( .A(n2909), .B(n4584), .Z(n31) );
  XNOR U133 ( .A(n2908), .B(n31), .Z(out[211]) );
  NANDN U134 ( .A(n2930), .B(n4734), .Z(n32) );
  XNOR U135 ( .A(n2929), .B(n32), .Z(out[217]) );
  ANDN U136 ( .B(n3847), .A(n3430), .Z(n33) );
  XNOR U137 ( .A(n3588), .B(n33), .Z(out[436]) );
  AND U138 ( .A(n3891), .B(n3464), .Z(n34) );
  XNOR U139 ( .A(n3610), .B(n34), .Z(out[446]) );
  NANDN U140 ( .A(n3639), .B(n3478), .Z(n35) );
  XNOR U141 ( .A(n3638), .B(n35), .Z(out[517]) );
  NANDN U142 ( .A(n3643), .B(n3479), .Z(n36) );
  XNOR U143 ( .A(n3642), .B(n36), .Z(out[518]) );
  NANDN U144 ( .A(n3647), .B(n3480), .Z(n37) );
  XNOR U145 ( .A(n3646), .B(n37), .Z(out[519]) );
  NAND U146 ( .A(n3485), .B(n3651), .Z(n38) );
  XNOR U147 ( .A(n3650), .B(n38), .Z(out[520]) );
  ANDN U148 ( .B(n3508), .A(n3698), .Z(n39) );
  XNOR U149 ( .A(n3699), .B(n39), .Z(out[531]) );
  ANDN U150 ( .B(n3512), .A(n3714), .Z(n40) );
  XNOR U151 ( .A(n3715), .B(n40), .Z(out[535]) );
  ANDN U152 ( .B(n3513), .A(n3724), .Z(n41) );
  XNOR U153 ( .A(n3725), .B(n41), .Z(out[536]) );
  ANDN U154 ( .B(n3514), .A(n3728), .Z(n42) );
  XNOR U155 ( .A(n3729), .B(n42), .Z(out[537]) );
  ANDN U156 ( .B(n3517), .A(n3736), .Z(n43) );
  XNOR U157 ( .A(n3737), .B(n43), .Z(out[539]) );
  NANDN U158 ( .A(n4433), .B(n4848), .Z(n44) );
  XNOR U159 ( .A(n4642), .B(n44), .Z(out[733]) );
  NANDN U160 ( .A(n4436), .B(n4852), .Z(n45) );
  XNOR U161 ( .A(n4645), .B(n45), .Z(out[734]) );
  NANDN U162 ( .A(n4439), .B(n4856), .Z(n46) );
  XNOR U163 ( .A(n4648), .B(n46), .Z(out[735]) );
  NANDN U164 ( .A(n4456), .B(n4872), .Z(n47) );
  XNOR U165 ( .A(n4655), .B(n47), .Z(out[738]) );
  NANDN U166 ( .A(n4882), .B(n4664), .Z(n48) );
  XNOR U167 ( .A(n4881), .B(n48), .Z(out[869]) );
  NANDN U168 ( .A(n4886), .B(n4669), .Z(n49) );
  XNOR U169 ( .A(n4885), .B(n49), .Z(out[870]) );
  NANDN U170 ( .A(n4890), .B(n4670), .Z(n50) );
  XNOR U171 ( .A(n4889), .B(n50), .Z(out[871]) );
  NANDN U172 ( .A(n4898), .B(n4672), .Z(n51) );
  XNOR U173 ( .A(n4897), .B(n51), .Z(out[873]) );
  NANDN U174 ( .A(n4902), .B(n4673), .Z(n52) );
  XNOR U175 ( .A(n4901), .B(n52), .Z(out[874]) );
  ANDN U176 ( .B(n4676), .A(n4913), .Z(n53) );
  XNOR U177 ( .A(n4914), .B(n53), .Z(out[876]) );
  ANDN U178 ( .B(n4677), .A(n4917), .Z(n54) );
  XNOR U179 ( .A(n4918), .B(n54), .Z(out[877]) );
  ANDN U180 ( .B(n4678), .A(n4921), .Z(n55) );
  XNOR U181 ( .A(n4922), .B(n55), .Z(out[878]) );
  ANDN U182 ( .B(n4679), .A(n4925), .Z(n56) );
  XNOR U183 ( .A(n4926), .B(n56), .Z(out[879]) );
  ANDN U184 ( .B(n4684), .A(n4929), .Z(n57) );
  XNOR U185 ( .A(n4930), .B(n57), .Z(out[880]) );
  ANDN U186 ( .B(n4685), .A(n4933), .Z(n58) );
  XNOR U187 ( .A(n4934), .B(n58), .Z(out[881]) );
  ANDN U188 ( .B(n4686), .A(n4937), .Z(n59) );
  XNOR U189 ( .A(n4938), .B(n59), .Z(out[882]) );
  ANDN U190 ( .B(n4687), .A(n4941), .Z(n60) );
  XNOR U191 ( .A(n4942), .B(n60), .Z(out[883]) );
  OR U192 ( .A(n5072), .B(n5073), .Z(n61) );
  XNOR U193 ( .A(n5074), .B(n61), .Z(out[977]) );
  OR U194 ( .A(n5075), .B(n5076), .Z(n62) );
  XNOR U195 ( .A(n5077), .B(n62), .Z(out[978]) );
  NANDN U196 ( .A(n1508), .B(n1914), .Z(n63) );
  XNOR U197 ( .A(n1761), .B(n63), .Z(out[1067]) );
  ANDN U198 ( .B(n5012), .A(n1600), .Z(n64) );
  XNOR U199 ( .A(n1813), .B(n64), .Z(out[1090]) );
  XNOR U200 ( .A(n564), .B(n681), .Z(n4051) );
  XNOR U201 ( .A(n1407), .B(n1685), .Z(n3179) );
  XNOR U202 ( .A(n1715), .B(n1423), .Z(n2296) );
  XNOR U203 ( .A(n1659), .B(n1660), .Z(n3065) );
  XNOR U204 ( .A(n1664), .B(n1665), .Z(n3067) );
  XNOR U205 ( .A(n1216), .B(n1492), .Z(n4084) );
  NANDN U206 ( .A(n2855), .B(n3899), .Z(n65) );
  XNOR U207 ( .A(n3023), .B(n65), .Z(out[191]) );
  NANDN U208 ( .A(n2918), .B(n4668), .Z(n66) );
  XNOR U209 ( .A(n2917), .B(n66), .Z(out[214]) );
  NANDN U210 ( .A(n2921), .B(n4683), .Z(n67) );
  XNOR U211 ( .A(n2920), .B(n67), .Z(out[215]) );
  ANDN U212 ( .B(n2954), .A(n5163), .Z(n68) );
  XNOR U213 ( .A(n3100), .B(n68), .Z(out[227]) );
  NAND U214 ( .A(n2858), .B(n2857), .Z(n69) );
  XNOR U215 ( .A(n3941), .B(n69), .Z(out[256]) );
  AND U216 ( .A(n3019), .B(n3808), .Z(n70) );
  XNOR U217 ( .A(n3809), .B(n70), .Z(out[317]) );
  ANDN U218 ( .B(n3617), .A(n3264), .Z(n71) );
  XNOR U219 ( .A(n3469), .B(n71), .Z(out[384]) );
  ANDN U220 ( .B(n3867), .A(n3442), .Z(n72) );
  XNOR U221 ( .A(n3596), .B(n72), .Z(out[440]) );
  ANDN U222 ( .B(n3883), .A(n3454), .Z(n73) );
  XNOR U223 ( .A(n3606), .B(n73), .Z(out[444]) );
  ANDN U224 ( .B(n3509), .A(n3702), .Z(n74) );
  XNOR U225 ( .A(n3703), .B(n74), .Z(out[532]) );
  ANDN U226 ( .B(n3510), .A(n3706), .Z(n75) );
  XNOR U227 ( .A(n3707), .B(n75), .Z(out[533]) );
  ANDN U228 ( .B(n3511), .A(n3710), .Z(n76) );
  XNOR U229 ( .A(n3711), .B(n76), .Z(out[534]) );
  NAND U230 ( .A(n4754), .B(n4361), .Z(n77) );
  XNOR U231 ( .A(n4578), .B(n77), .Z(out[711]) );
  NANDN U232 ( .A(n4418), .B(n4828), .Z(n78) );
  XNOR U233 ( .A(n4623), .B(n78), .Z(out[728]) );
  NANDN U234 ( .A(n4468), .B(n4888), .Z(n79) );
  XNOR U235 ( .A(n4669), .B(n79), .Z(out[742]) );
  NOR U236 ( .A(n4601), .B(n4391), .Z(n80) );
  XNOR U237 ( .A(n4791), .B(n80), .Z(out[784]) );
  NANDN U238 ( .A(n4894), .B(n4671), .Z(n81) );
  XNOR U239 ( .A(n4893), .B(n81), .Z(out[872]) );
  ANDN U240 ( .B(n4688), .A(n4945), .Z(n82) );
  XNOR U241 ( .A(n4946), .B(n82), .Z(out[884]) );
  ANDN U242 ( .B(n4689), .A(n4949), .Z(n83) );
  XNOR U243 ( .A(n4950), .B(n83), .Z(out[885]) );
  ANDN U244 ( .B(n4690), .A(n4957), .Z(n84) );
  XNOR U245 ( .A(n4958), .B(n84), .Z(out[886]) );
  OR U246 ( .A(n5086), .B(n5087), .Z(n85) );
  XNOR U247 ( .A(n5088), .B(n85), .Z(out[980]) );
  OR U248 ( .A(n5089), .B(n5090), .Z(n86) );
  XNOR U249 ( .A(n5091), .B(n86), .Z(out[981]) );
  OR U250 ( .A(n5092), .B(n5093), .Z(n87) );
  XNOR U251 ( .A(n5094), .B(n87), .Z(out[982]) );
  OR U252 ( .A(n5095), .B(n5096), .Z(n88) );
  XNOR U253 ( .A(n5097), .B(n88), .Z(out[983]) );
  OR U254 ( .A(n5098), .B(n5099), .Z(n89) );
  XNOR U255 ( .A(n5100), .B(n89), .Z(out[984]) );
  OR U256 ( .A(n5101), .B(n5102), .Z(n90) );
  XNOR U257 ( .A(n5103), .B(n90), .Z(out[985]) );
  OR U258 ( .A(n5104), .B(n5105), .Z(n91) );
  XNOR U259 ( .A(n5106), .B(n91), .Z(out[986]) );
  OR U260 ( .A(n5107), .B(n5108), .Z(n92) );
  XNOR U261 ( .A(n5109), .B(n92), .Z(out[987]) );
  OR U262 ( .A(n5114), .B(n5115), .Z(n93) );
  XNOR U263 ( .A(n5116), .B(n93), .Z(out[989]) );
  OR U264 ( .A(n5121), .B(n5122), .Z(n94) );
  XNOR U265 ( .A(n5123), .B(n94), .Z(out[990]) );
  ANDN U266 ( .B(n1902), .A(n1494), .Z(n95) );
  XNOR U267 ( .A(n1755), .B(n95), .Z(out[1064]) );
  ANDN U268 ( .B(n1906), .A(n1498), .Z(n96) );
  XNOR U269 ( .A(n1757), .B(n96), .Z(out[1065]) );
  ANDN U270 ( .B(n1910), .A(n1504), .Z(n97) );
  XNOR U271 ( .A(n1759), .B(n97), .Z(out[1066]) );
  ANDN U272 ( .B(n1920), .A(n1512), .Z(n98) );
  XNOR U273 ( .A(n1762), .B(n98), .Z(out[1068]) );
  ANDN U274 ( .B(n1924), .A(n1516), .Z(n99) );
  XNOR U275 ( .A(n1764), .B(n99), .Z(out[1069]) );
  ANDN U276 ( .B(n1928), .A(n1520), .Z(n100) );
  XNOR U277 ( .A(n1766), .B(n100), .Z(out[1070]) );
  ANDN U278 ( .B(n1932), .A(n1524), .Z(n101) );
  XNOR U279 ( .A(n1768), .B(n101), .Z(out[1071]) );
  ANDN U280 ( .B(n1936), .A(n1528), .Z(n102) );
  XNOR U281 ( .A(n1772), .B(n102), .Z(out[1072]) );
  ANDN U282 ( .B(n1940), .A(n1532), .Z(n103) );
  XNOR U283 ( .A(n1774), .B(n103), .Z(out[1073]) );
  ANDN U284 ( .B(n1944), .A(n1536), .Z(n104) );
  XNOR U285 ( .A(n1776), .B(n104), .Z(out[1074]) );
  ANDN U286 ( .B(n1948), .A(n1540), .Z(n105) );
  XNOR U287 ( .A(n1778), .B(n105), .Z(out[1075]) );
  ANDN U288 ( .B(n1952), .A(n1546), .Z(n106) );
  XNOR U289 ( .A(n1780), .B(n106), .Z(out[1076]) );
  ANDN U290 ( .B(n1956), .A(n1550), .Z(n107) );
  XNOR U291 ( .A(n1782), .B(n107), .Z(out[1077]) );
  ANDN U292 ( .B(n1962), .A(n1554), .Z(n108) );
  XNOR U293 ( .A(n1784), .B(n108), .Z(out[1078]) );
  ANDN U294 ( .B(n1978), .A(n1570), .Z(n109) );
  XNOR U295 ( .A(n1794), .B(n109), .Z(out[1082]) );
  ANDN U296 ( .B(n1982), .A(n1574), .Z(n110) );
  XNOR U297 ( .A(n1796), .B(n110), .Z(out[1083]) );
  ANDN U298 ( .B(n1986), .A(n1578), .Z(n111) );
  XNOR U299 ( .A(n1798), .B(n111), .Z(out[1084]) );
  ANDN U300 ( .B(n1990), .A(n1582), .Z(n112) );
  XNOR U301 ( .A(n1800), .B(n112), .Z(out[1085]) );
  ANDN U302 ( .B(n1994), .A(n1586), .Z(n113) );
  XNOR U303 ( .A(n1802), .B(n113), .Z(out[1086]) );
  AND U304 ( .A(n1998), .B(n1588), .Z(n114) );
  XNOR U305 ( .A(n1804), .B(n114), .Z(out[1087]) );
  ANDN U306 ( .B(n5004), .A(n1592), .Z(n115) );
  XNOR U307 ( .A(n1807), .B(n115), .Z(out[1088]) );
  ANDN U308 ( .B(n5028), .A(n1616), .Z(n116) );
  XNOR U309 ( .A(n1826), .B(n116), .Z(out[1094]) );
  ANDN U310 ( .B(n5040), .A(n1629), .Z(n117) );
  XNOR U311 ( .A(n1831), .B(n117), .Z(out[1097]) );
  ANDN U312 ( .B(n5048), .A(n1633), .Z(n118) );
  XNOR U313 ( .A(n1833), .B(n118), .Z(out[1098]) );
  ANDN U314 ( .B(n5052), .A(n1637), .Z(n119) );
  XNOR U315 ( .A(n1835), .B(n119), .Z(out[1099]) );
  ANDN U316 ( .B(n5056), .A(n1641), .Z(n120) );
  XNOR U317 ( .A(n1837), .B(n120), .Z(out[1100]) );
  ANDN U318 ( .B(n5060), .A(n1645), .Z(n121) );
  XNOR U319 ( .A(n1839), .B(n121), .Z(out[1101]) );
  ANDN U320 ( .B(n5064), .A(n1649), .Z(n122) );
  XNOR U321 ( .A(n1843), .B(n122), .Z(out[1102]) );
  AND U322 ( .A(n5071), .B(n1657), .Z(n123) );
  XNOR U323 ( .A(n1847), .B(n123), .Z(out[1104]) );
  AND U324 ( .A(n5074), .B(n1661), .Z(n124) );
  XNOR U325 ( .A(n1849), .B(n124), .Z(out[1105]) );
  ANDN U326 ( .B(n5113), .A(n1708), .Z(n125) );
  XNOR U327 ( .A(n1873), .B(n125), .Z(out[1116]) );
  ANDN U328 ( .B(n5139), .A(n1732), .Z(n126) );
  XNOR U329 ( .A(n1887), .B(n126), .Z(out[1122]) );
  NANDN U330 ( .A(n1912), .B(n1761), .Z(n127) );
  XNOR U331 ( .A(n1911), .B(n127), .Z(out[1195]) );
  NANDN U332 ( .A(n2239), .B(n2547), .Z(n128) );
  XNOR U333 ( .A(n2379), .B(n128), .Z(out[1371]) );
  ANDN U334 ( .B(n2438), .A(n2437), .Z(n129) );
  XNOR U335 ( .A(n2439), .B(round_const[0]), .Z(n130) );
  XOR U336 ( .A(n129), .B(n130), .Z(out[1536]) );
  ANDN U337 ( .B(n2441), .A(n2440), .Z(n131) );
  XNOR U338 ( .A(n2442), .B(round_const[1]), .Z(n132) );
  XOR U339 ( .A(n131), .B(n132), .Z(out[1537]) );
  XNOR U340 ( .A(n1420), .B(n1707), .Z(n3189) );
  XNOR U341 ( .A(n1429), .B(n1727), .Z(n3203) );
  XNOR U342 ( .A(n1483), .B(n1171), .Z(n4068) );
  XNOR U343 ( .A(n1489), .B(n1201), .Z(n4080) );
  XNOR U344 ( .A(n1692), .B(n1693), .Z(n3085) );
  XNOR U345 ( .A(n1700), .B(n1701), .Z(n3089) );
  XNOR U346 ( .A(n3960), .B(in[1485]), .Z(n4785) );
  XNOR U347 ( .A(n3964), .B(in[1486]), .Z(n4789) );
  XNOR U348 ( .A(n3968), .B(in[1487]), .Z(n4793) );
  XNOR U349 ( .A(n3972), .B(in[1488]), .Z(n4797) );
  XNOR U350 ( .A(n3976), .B(in[1489]), .Z(n4801) );
  XNOR U351 ( .A(n3980), .B(in[1490]), .Z(n4805) );
  NAND U352 ( .A(n2906), .B(n4555), .Z(n133) );
  XNOR U353 ( .A(n2905), .B(n133), .Z(out[210]) );
  NAND U354 ( .A(n2912), .B(n4609), .Z(n134) );
  XNOR U355 ( .A(n2911), .B(n134), .Z(out[212]) );
  NANDN U356 ( .A(n2915), .B(n4638), .Z(n135) );
  XNOR U357 ( .A(n2914), .B(n135), .Z(out[213]) );
  ANDN U358 ( .B(n3851), .A(n3433), .Z(n136) );
  XNOR U359 ( .A(n3590), .B(n136), .Z(out[437]) );
  NAND U360 ( .A(n3477), .B(n3635), .Z(n137) );
  XNOR U361 ( .A(n3634), .B(n137), .Z(out[516]) );
  ANDN U362 ( .B(n3502), .A(n3690), .Z(n138) );
  XNOR U363 ( .A(n3691), .B(n138), .Z(out[529]) );
  ANDN U364 ( .B(n3507), .A(n3694), .Z(n139) );
  XNOR U365 ( .A(n3695), .B(n139), .Z(out[530]) );
  AND U366 ( .A(n4746), .B(n4355), .Z(n140) );
  XNOR U367 ( .A(n4574), .B(n140), .Z(out[709]) );
  AND U368 ( .A(n4750), .B(n4358), .Z(n141) );
  XNOR U369 ( .A(n4576), .B(n141), .Z(out[710]) );
  AND U370 ( .A(n4758), .B(n4363), .Z(n142) );
  XNOR U371 ( .A(n4585), .B(n142), .Z(out[712]) );
  AND U372 ( .A(n4762), .B(n4366), .Z(n143) );
  XNOR U373 ( .A(n4587), .B(n143), .Z(out[713]) );
  AND U374 ( .A(n4766), .B(n4369), .Z(n144) );
  XNOR U375 ( .A(n4589), .B(n144), .Z(out[714]) );
  AND U376 ( .A(n4770), .B(n4372), .Z(n145) );
  XNOR U377 ( .A(n4591), .B(n145), .Z(out[715]) );
  AND U378 ( .A(n4774), .B(n4379), .Z(n146) );
  XNOR U379 ( .A(n4593), .B(n146), .Z(out[716]) );
  ANDN U380 ( .B(n4817), .A(n4412), .Z(n147) );
  XNOR U381 ( .A(n4618), .B(n147), .Z(out[726]) );
  NANDN U382 ( .A(n4450), .B(n4860), .Z(n148) );
  XNOR U383 ( .A(n4649), .B(n148), .Z(out[736]) );
  NANDN U384 ( .A(n4453), .B(n4864), .Z(n149) );
  XNOR U385 ( .A(n4652), .B(n149), .Z(out[737]) );
  NANDN U386 ( .A(n4459), .B(n4876), .Z(n150) );
  XNOR U387 ( .A(n4658), .B(n150), .Z(out[739]) );
  NANDN U388 ( .A(n4462), .B(n4880), .Z(n151) );
  XNOR U389 ( .A(n4661), .B(n151), .Z(out[740]) );
  NANDN U390 ( .A(n4465), .B(n4884), .Z(n152) );
  XNOR U391 ( .A(n4664), .B(n152), .Z(out[741]) );
  NOR U392 ( .A(n4560), .B(n4340), .Z(n153) );
  XNOR U393 ( .A(n4715), .B(n153), .Z(out[768]) );
  NOR U394 ( .A(n4563), .B(n4342), .Z(n154) );
  XNOR U395 ( .A(n4719), .B(n154), .Z(out[769]) );
  NOR U396 ( .A(n4566), .B(n4348), .Z(n155) );
  XNOR U397 ( .A(n4723), .B(n155), .Z(out[770]) );
  NOR U398 ( .A(n4569), .B(n4350), .Z(n156) );
  XNOR U399 ( .A(n4727), .B(n156), .Z(out[771]) );
  NOR U400 ( .A(n4578), .B(n4361), .Z(n157) );
  XNOR U401 ( .A(n4751), .B(n157), .Z(out[775]) );
  NOR U402 ( .A(n4706), .B(n4551), .Z(n158) );
  XNOR U403 ( .A(n4985), .B(n158), .Z(out[829]) );
  NOR U404 ( .A(n4709), .B(n4557), .Z(n159) );
  XNOR U405 ( .A(n4989), .B(n159), .Z(out[830]) );
  NOR U406 ( .A(n4712), .B(n4559), .Z(n160) );
  XNOR U407 ( .A(n4993), .B(n160), .Z(out[831]) );
  NAND U408 ( .A(n4648), .B(n4854), .Z(n161) );
  XNOR U409 ( .A(n4853), .B(n161), .Z(out[863]) );
  OR U410 ( .A(n5069), .B(n5070), .Z(n162) );
  XNOR U411 ( .A(n5071), .B(n162), .Z(out[976]) );
  ANDN U412 ( .B(n5008), .A(n1596), .Z(n163) );
  XNOR U413 ( .A(n1810), .B(n163), .Z(out[1089]) );
  ANDN U414 ( .B(n5016), .A(n1604), .Z(n164) );
  XNOR U415 ( .A(n1816), .B(n164), .Z(out[1091]) );
  ANDN U416 ( .B(n5020), .A(n1608), .Z(n165) );
  XNOR U417 ( .A(n1821), .B(n165), .Z(out[1092]) );
  ANDN U418 ( .B(n5024), .A(n1612), .Z(n166) );
  XNOR U419 ( .A(n1824), .B(n166), .Z(out[1093]) );
  ANDN U420 ( .B(n5032), .A(n1620), .Z(n167) );
  XNOR U421 ( .A(n1827), .B(n167), .Z(out[1095]) );
  ANDN U422 ( .B(n5036), .A(n1625), .Z(n168) );
  XNOR U423 ( .A(n1829), .B(n168), .Z(out[1096]) );
  AND U424 ( .A(n5068), .B(n1653), .Z(n169) );
  XNOR U425 ( .A(n1845), .B(n169), .Z(out[1103]) );
  AND U426 ( .A(n5077), .B(n1666), .Z(n170) );
  XNOR U427 ( .A(n1851), .B(n170), .Z(out[1106]) );
  ANDN U428 ( .B(n5081), .A(n1670), .Z(n171) );
  XNOR U429 ( .A(n1853), .B(n171), .Z(out[1107]) );
  ANDN U430 ( .B(n5088), .A(n1674), .Z(n172) );
  XNOR U431 ( .A(n1855), .B(n172), .Z(out[1108]) );
  ANDN U432 ( .B(n5091), .A(n1678), .Z(n173) );
  XNOR U433 ( .A(n1857), .B(n173), .Z(out[1109]) );
  ANDN U434 ( .B(n5094), .A(n1682), .Z(n174) );
  XNOR U435 ( .A(n1859), .B(n174), .Z(out[1110]) );
  ANDN U436 ( .B(n5097), .A(n1686), .Z(n175) );
  XNOR U437 ( .A(n1861), .B(n175), .Z(out[1111]) );
  ANDN U438 ( .B(n5100), .A(n1690), .Z(n176) );
  XNOR U439 ( .A(n1865), .B(n176), .Z(out[1112]) );
  ANDN U440 ( .B(n5103), .A(n1694), .Z(n177) );
  XNOR U441 ( .A(n1867), .B(n177), .Z(out[1113]) );
  ANDN U442 ( .B(n5106), .A(n1698), .Z(n178) );
  XNOR U443 ( .A(n1869), .B(n178), .Z(out[1114]) );
  ANDN U444 ( .B(n5116), .A(n1712), .Z(n179) );
  XNOR U445 ( .A(n1875), .B(n179), .Z(out[1117]) );
  OR U446 ( .A(n5026), .B(n1826), .Z(n180) );
  XNOR U447 ( .A(n5025), .B(n180), .Z(out[1222]) );
  ANDN U448 ( .B(n2518), .A(n2224), .Z(n181) );
  XNOR U449 ( .A(n2365), .B(n181), .Z(out[1364]) );
  ANDN U450 ( .B(n2526), .A(n2229), .Z(n182) );
  XNOR U451 ( .A(n2369), .B(n182), .Z(out[1366]) );
  ANDN U452 ( .B(n2530), .A(n2231), .Z(n183) );
  XNOR U453 ( .A(n2371), .B(n183), .Z(out[1367]) );
  ANDN U454 ( .B(n2535), .A(n2233), .Z(n184) );
  XNOR U455 ( .A(n2373), .B(n184), .Z(out[1368]) );
  ANDN U456 ( .B(n2539), .A(n2235), .Z(n185) );
  XNOR U457 ( .A(n2375), .B(n185), .Z(out[1369]) );
  ANDN U458 ( .B(n2543), .A(n2237), .Z(n186) );
  XNOR U459 ( .A(n2377), .B(n186), .Z(out[1370]) );
  ANDN U460 ( .B(n2551), .A(n2241), .Z(n187) );
  XNOR U461 ( .A(n2382), .B(n187), .Z(out[1372]) );
  ANDN U462 ( .B(n2555), .A(n2243), .Z(n188) );
  XNOR U463 ( .A(n2384), .B(n188), .Z(out[1373]) );
  ANDN U464 ( .B(n2559), .A(n2245), .Z(n189) );
  XNOR U465 ( .A(n2386), .B(n189), .Z(out[1374]) );
  ANDN U466 ( .B(n2562), .A(n2247), .Z(n190) );
  XNOR U467 ( .A(n2388), .B(n190), .Z(out[1375]) );
  ANDN U468 ( .B(n2568), .A(n2250), .Z(n191) );
  XNOR U469 ( .A(n2390), .B(n191), .Z(out[1376]) );
  ANDN U470 ( .B(n2648), .A(n2289), .Z(n192) );
  XNOR U471 ( .A(n2412), .B(n192), .Z(out[1395]) );
  ANDN U472 ( .B(n2652), .A(n2292), .Z(n193) );
  XNOR U473 ( .A(n2414), .B(n193), .Z(out[1396]) );
  ANDN U474 ( .B(n2656), .A(n2294), .Z(n194) );
  XNOR U475 ( .A(n2416), .B(n194), .Z(out[1397]) );
  ANDN U476 ( .B(n2674), .A(n2303), .Z(n195) );
  XNOR U477 ( .A(n2421), .B(n195), .Z(out[1401]) );
  ANDN U478 ( .B(n2678), .A(n2305), .Z(n196) );
  XNOR U479 ( .A(n2424), .B(n196), .Z(out[1402]) );
  NAND U480 ( .A(n2495), .B(n2355), .Z(n197) );
  XNOR U481 ( .A(n2494), .B(n197), .Z(out[1487]) );
  NAND U482 ( .A(n2500), .B(n2357), .Z(n198) );
  XNOR U483 ( .A(n2499), .B(n198), .Z(out[1488]) );
  NAND U484 ( .A(n2544), .B(n2379), .Z(n199) );
  XNOR U485 ( .A(n2545), .B(n199), .Z(out[1499]) );
  NAND U486 ( .A(n2569), .B(n2392), .Z(n200) );
  XNOR U487 ( .A(n2570), .B(n200), .Z(out[1505]) );
  NAND U488 ( .A(n2575), .B(n2393), .Z(n201) );
  XNOR U489 ( .A(n2576), .B(n201), .Z(out[1506]) );
  NAND U490 ( .A(n2579), .B(n2394), .Z(n202) );
  XNOR U491 ( .A(n2580), .B(n202), .Z(out[1507]) );
  NAND U492 ( .A(n2583), .B(n2395), .Z(n203) );
  XNOR U493 ( .A(n2584), .B(n203), .Z(out[1508]) );
  NAND U494 ( .A(n2587), .B(n2396), .Z(n204) );
  XNOR U495 ( .A(n2588), .B(n204), .Z(out[1509]) );
  NAND U496 ( .A(n2591), .B(n2398), .Z(n205) );
  XNOR U497 ( .A(n2592), .B(n205), .Z(out[1510]) );
  AND U498 ( .A(n2595), .B(n2399), .Z(n206) );
  XNOR U499 ( .A(n2596), .B(n206), .Z(out[1511]) );
  AND U500 ( .A(n2599), .B(n2400), .Z(n207) );
  XNOR U501 ( .A(n2600), .B(n207), .Z(out[1512]) );
  AND U502 ( .A(n2603), .B(n2401), .Z(n208) );
  XNOR U503 ( .A(n2604), .B(n208), .Z(out[1513]) );
  NAND U504 ( .A(n2607), .B(n2402), .Z(n209) );
  XNOR U505 ( .A(n2608), .B(n209), .Z(out[1514]) );
  AND U506 ( .A(n2611), .B(n2403), .Z(n210) );
  XNOR U507 ( .A(n2612), .B(n210), .Z(out[1515]) );
  AND U508 ( .A(n2617), .B(n2404), .Z(n211) );
  XNOR U509 ( .A(n2618), .B(n211), .Z(out[1516]) );
  ANDN U510 ( .B(n2405), .A(n2621), .Z(n212) );
  XNOR U511 ( .A(n2622), .B(n212), .Z(out[1517]) );
  AND U512 ( .A(n2625), .B(n2406), .Z(n213) );
  XNOR U513 ( .A(n2626), .B(n213), .Z(out[1518]) );
  AND U514 ( .A(n2629), .B(n2407), .Z(n214) );
  XNOR U515 ( .A(n2630), .B(n214), .Z(out[1519]) );
  AND U516 ( .A(n2633), .B(n2409), .Z(n215) );
  XNOR U517 ( .A(n2634), .B(n215), .Z(out[1520]) );
  AND U518 ( .A(n2637), .B(n2410), .Z(n216) );
  XNOR U519 ( .A(n2638), .B(n216), .Z(out[1521]) );
  AND U520 ( .A(n2641), .B(n2411), .Z(n217) );
  XNOR U521 ( .A(n2642), .B(n217), .Z(out[1522]) );
  AND U522 ( .A(n2659), .B(n2418), .Z(n218) );
  XNOR U523 ( .A(n2660), .B(n218), .Z(out[1526]) );
  AND U524 ( .A(n2663), .B(n2419), .Z(n219) );
  XNOR U525 ( .A(n2664), .B(n219), .Z(out[1527]) );
  AND U526 ( .A(n2667), .B(n2420), .Z(n220) );
  XNOR U527 ( .A(n2668), .B(n220), .Z(out[1528]) );
  ANDN U528 ( .B(n2471), .A(n2470), .Z(n221) );
  XNOR U529 ( .A(n2469), .B(n221), .Z(out[1544]) );
  ANDN U530 ( .B(n2474), .A(n2473), .Z(n222) );
  XNOR U531 ( .A(n2472), .B(n222), .Z(out[1545]) );
  ANDN U532 ( .B(n2477), .A(n2476), .Z(n223) );
  XNOR U533 ( .A(n2475), .B(n223), .Z(out[1546]) );
  ANDN U534 ( .B(n2488), .A(n2487), .Z(n224) );
  XNOR U535 ( .A(n2486), .B(n224), .Z(out[1549]) );
  ANDN U536 ( .B(n2696), .A(n2695), .Z(n225) );
  XNOR U537 ( .A(n2697), .B(round_const_63), .Z(n226) );
  XOR U538 ( .A(n225), .B(n226), .Z(out[1599]) );
  XNOR U539 ( .A(in[1162]), .B(n838), .Z(n227) );
  XOR U540 ( .A(in[1469]), .B(in[509]), .Z(n229) );
  XNOR U541 ( .A(in[829]), .B(in[189]), .Z(n228) );
  XNOR U542 ( .A(n229), .B(n228), .Z(n230) );
  XNOR U543 ( .A(in[1149]), .B(n230), .Z(n1099) );
  XOR U544 ( .A(in[1598]), .B(in[638]), .Z(n232) );
  XNOR U545 ( .A(in[958]), .B(in[318]), .Z(n231) );
  XNOR U546 ( .A(n232), .B(n231), .Z(n233) );
  XNOR U547 ( .A(in[1278]), .B(n233), .Z(n1669) );
  XNOR U548 ( .A(n1099), .B(n1669), .Z(n3291) );
  XOR U549 ( .A(in[254]), .B(n3291), .Z(n3940) );
  XOR U550 ( .A(in[1345]), .B(in[65]), .Z(n235) );
  XNOR U551 ( .A(in[1025]), .B(in[385]), .Z(n234) );
  XNOR U552 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U553 ( .A(in[705]), .B(n236), .Z(n1677) );
  XOR U554 ( .A(in[1474]), .B(in[514]), .Z(n238) );
  XNOR U555 ( .A(in[834]), .B(in[194]), .Z(n237) );
  XNOR U556 ( .A(n238), .B(n237), .Z(n239) );
  XOR U557 ( .A(in[1154]), .B(n239), .Z(n1401) );
  XOR U558 ( .A(in[1410]), .B(n3175), .Z(n3941) );
  XOR U559 ( .A(in[137]), .B(in[457]), .Z(n241) );
  XNOR U560 ( .A(in[777]), .B(in[1417]), .Z(n240) );
  XNOR U561 ( .A(n241), .B(n240), .Z(n242) );
  XNOR U562 ( .A(in[1097]), .B(n242), .Z(n1358) );
  XOR U563 ( .A(in[328]), .B(in[8]), .Z(n244) );
  XNOR U564 ( .A(in[968]), .B(in[648]), .Z(n243) );
  XNOR U565 ( .A(n244), .B(n243), .Z(n245) );
  XNOR U566 ( .A(in[1288]), .B(n245), .Z(n1414) );
  XOR U567 ( .A(n1358), .B(n1414), .Z(n4455) );
  XNOR U568 ( .A(in[1033]), .B(n4455), .Z(n2858) );
  OR U569 ( .A(n3941), .B(n2858), .Z(n246) );
  XOR U570 ( .A(n3940), .B(n246), .Z(out[0]) );
  XOR U571 ( .A(in[1386]), .B(in[106]), .Z(n248) );
  XNOR U572 ( .A(in[1066]), .B(in[746]), .Z(n247) );
  XNOR U573 ( .A(n248), .B(n247), .Z(n249) );
  XNOR U574 ( .A(in[426]), .B(n249), .Z(n702) );
  XOR U575 ( .A(in[1515]), .B(in[555]), .Z(n251) );
  XNOR U576 ( .A(in[875]), .B(in[235]), .Z(n250) );
  XNOR U577 ( .A(n251), .B(n250), .Z(n252) );
  XNOR U578 ( .A(in[1195]), .B(n252), .Z(n1523) );
  XOR U579 ( .A(n702), .B(n1523), .Z(n4111) );
  XOR U580 ( .A(in[171]), .B(n4111), .Z(n1494) );
  XOR U581 ( .A(in[140]), .B(in[460]), .Z(n254) );
  XNOR U582 ( .A(in[1100]), .B(in[1420]), .Z(n253) );
  XNOR U583 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U584 ( .A(in[780]), .B(n255), .Z(n1380) );
  XOR U585 ( .A(in[971]), .B(in[1291]), .Z(n257) );
  XNOR U586 ( .A(in[11]), .B(in[331]), .Z(n256) );
  XNOR U587 ( .A(n257), .B(n256), .Z(n258) );
  XOR U588 ( .A(in[651]), .B(n258), .Z(n1422) );
  XNOR U589 ( .A(in[1356]), .B(n4464), .Z(n1902) );
  XOR U590 ( .A(in[1364]), .B(in[724]), .Z(n260) );
  XNOR U591 ( .A(in[84]), .B(in[404]), .Z(n259) );
  XNOR U592 ( .A(n260), .B(n259), .Z(n261) );
  XNOR U593 ( .A(in[1044]), .B(n261), .Z(n1004) );
  XOR U594 ( .A(in[1555]), .B(in[595]), .Z(n263) );
  XNOR U595 ( .A(in[915]), .B(in[275]), .Z(n262) );
  XNOR U596 ( .A(n263), .B(n262), .Z(n264) );
  XNOR U597 ( .A(in[1235]), .B(n264), .Z(n716) );
  XOR U598 ( .A(n1004), .B(n716), .Z(n4252) );
  XOR U599 ( .A(in[980]), .B(n4252), .Z(n1899) );
  NANDN U600 ( .A(n1902), .B(n1899), .Z(n265) );
  XNOR U601 ( .A(n1494), .B(n265), .Z(out[1000]) );
  XOR U602 ( .A(in[1387]), .B(in[107]), .Z(n267) );
  XNOR U603 ( .A(in[1067]), .B(in[747]), .Z(n266) );
  XNOR U604 ( .A(n267), .B(n266), .Z(n268) );
  XNOR U605 ( .A(in[427]), .B(n268), .Z(n713) );
  XOR U606 ( .A(in[1516]), .B(in[556]), .Z(n270) );
  XNOR U607 ( .A(in[876]), .B(in[236]), .Z(n269) );
  XNOR U608 ( .A(n270), .B(n269), .Z(n271) );
  XNOR U609 ( .A(in[1196]), .B(n271), .Z(n1527) );
  XOR U610 ( .A(n713), .B(n1527), .Z(n4119) );
  XOR U611 ( .A(in[172]), .B(n4119), .Z(n1498) );
  XOR U612 ( .A(in[972]), .B(in[12]), .Z(n273) );
  XNOR U613 ( .A(in[1292]), .B(in[332]), .Z(n272) );
  XNOR U614 ( .A(n273), .B(n272), .Z(n274) );
  XNOR U615 ( .A(in[652]), .B(n274), .Z(n1424) );
  XOR U616 ( .A(in[141]), .B(in[461]), .Z(n276) );
  XNOR U617 ( .A(in[1101]), .B(in[1421]), .Z(n275) );
  XNOR U618 ( .A(n276), .B(n275), .Z(n277) );
  XOR U619 ( .A(in[781]), .B(n277), .Z(n1384) );
  XNOR U620 ( .A(in[1357]), .B(n4467), .Z(n1906) );
  XOR U621 ( .A(in[1365]), .B(in[725]), .Z(n279) );
  XNOR U622 ( .A(in[85]), .B(in[405]), .Z(n278) );
  XNOR U623 ( .A(n279), .B(n278), .Z(n280) );
  XNOR U624 ( .A(in[1045]), .B(n280), .Z(n1017) );
  XOR U625 ( .A(in[1556]), .B(in[596]), .Z(n282) );
  XNOR U626 ( .A(in[916]), .B(in[276]), .Z(n281) );
  XNOR U627 ( .A(n282), .B(n281), .Z(n283) );
  XNOR U628 ( .A(in[1236]), .B(n283), .Z(n731) );
  XOR U629 ( .A(n1017), .B(n731), .Z(n4255) );
  XOR U630 ( .A(in[981]), .B(n4255), .Z(n1903) );
  NANDN U631 ( .A(n1906), .B(n1903), .Z(n284) );
  XNOR U632 ( .A(n1498), .B(n284), .Z(out[1001]) );
  XOR U633 ( .A(in[1388]), .B(in[108]), .Z(n286) );
  XNOR U634 ( .A(in[1068]), .B(in[748]), .Z(n285) );
  XNOR U635 ( .A(n286), .B(n285), .Z(n287) );
  XNOR U636 ( .A(in[428]), .B(n287), .Z(n1591) );
  XOR U637 ( .A(in[1517]), .B(in[557]), .Z(n289) );
  XNOR U638 ( .A(in[877]), .B(in[237]), .Z(n288) );
  XNOR U639 ( .A(n289), .B(n288), .Z(n290) );
  XNOR U640 ( .A(in[1197]), .B(n290), .Z(n1531) );
  XOR U641 ( .A(n1591), .B(n1531), .Z(n1363) );
  XOR U642 ( .A(in[173]), .B(n1363), .Z(n1504) );
  XOR U643 ( .A(in[973]), .B(in[13]), .Z(n292) );
  XNOR U644 ( .A(in[1293]), .B(in[333]), .Z(n291) );
  XNOR U645 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U646 ( .A(in[653]), .B(n293), .Z(n1426) );
  XOR U647 ( .A(in[142]), .B(in[1422]), .Z(n295) );
  XNOR U648 ( .A(in[1102]), .B(in[782]), .Z(n294) );
  XNOR U649 ( .A(n295), .B(n294), .Z(n296) );
  XOR U650 ( .A(in[462]), .B(n296), .Z(n1388) );
  XNOR U651 ( .A(in[1358]), .B(n4470), .Z(n1910) );
  XOR U652 ( .A(in[1366]), .B(in[726]), .Z(n298) );
  XNOR U653 ( .A(in[86]), .B(in[406]), .Z(n297) );
  XNOR U654 ( .A(n298), .B(n297), .Z(n299) );
  XNOR U655 ( .A(in[1046]), .B(n299), .Z(n1030) );
  XOR U656 ( .A(in[1557]), .B(in[597]), .Z(n301) );
  XNOR U657 ( .A(in[917]), .B(in[277]), .Z(n300) );
  XNOR U658 ( .A(n301), .B(n300), .Z(n302) );
  XNOR U659 ( .A(in[1237]), .B(n302), .Z(n746) );
  XOR U660 ( .A(n1030), .B(n746), .Z(n4256) );
  XOR U661 ( .A(in[982]), .B(n4256), .Z(n1907) );
  NANDN U662 ( .A(n1910), .B(n1907), .Z(n303) );
  XNOR U663 ( .A(n1504), .B(n303), .Z(out[1002]) );
  XOR U664 ( .A(in[1389]), .B(in[109]), .Z(n305) );
  XNOR U665 ( .A(in[1069]), .B(in[749]), .Z(n304) );
  XNOR U666 ( .A(n305), .B(n304), .Z(n306) );
  XNOR U667 ( .A(in[429]), .B(n306), .Z(n1595) );
  XOR U668 ( .A(in[1518]), .B(in[558]), .Z(n308) );
  XNOR U669 ( .A(in[878]), .B(in[238]), .Z(n307) );
  XNOR U670 ( .A(n308), .B(n307), .Z(n309) );
  XNOR U671 ( .A(in[1198]), .B(n309), .Z(n1535) );
  XOR U672 ( .A(n1595), .B(n1535), .Z(n1403) );
  XOR U673 ( .A(in[174]), .B(n1403), .Z(n1508) );
  XOR U674 ( .A(in[974]), .B(in[14]), .Z(n311) );
  XNOR U675 ( .A(in[1294]), .B(in[334]), .Z(n310) );
  XNOR U676 ( .A(n311), .B(n310), .Z(n312) );
  XNOR U677 ( .A(in[654]), .B(n312), .Z(n1428) );
  XOR U678 ( .A(in[143]), .B(in[1423]), .Z(n314) );
  XNOR U679 ( .A(in[1103]), .B(in[783]), .Z(n313) );
  XNOR U680 ( .A(n314), .B(n313), .Z(n315) );
  XOR U681 ( .A(in[463]), .B(n315), .Z(n1392) );
  XNOR U682 ( .A(in[1359]), .B(n4473), .Z(n1914) );
  XOR U683 ( .A(in[1367]), .B(in[727]), .Z(n317) );
  XNOR U684 ( .A(in[87]), .B(in[407]), .Z(n316) );
  XNOR U685 ( .A(n317), .B(n316), .Z(n318) );
  XNOR U686 ( .A(in[1047]), .B(n318), .Z(n1043) );
  XOR U687 ( .A(in[1558]), .B(in[598]), .Z(n320) );
  XNOR U688 ( .A(in[918]), .B(in[278]), .Z(n319) );
  XNOR U689 ( .A(n320), .B(n319), .Z(n321) );
  XNOR U690 ( .A(in[1238]), .B(n321), .Z(n761) );
  XOR U691 ( .A(n1043), .B(n761), .Z(n4257) );
  XOR U692 ( .A(in[983]), .B(n4257), .Z(n1911) );
  NANDN U693 ( .A(n1914), .B(n1911), .Z(n322) );
  XNOR U694 ( .A(n1508), .B(n322), .Z(out[1003]) );
  XOR U695 ( .A(in[1390]), .B(in[110]), .Z(n324) );
  XNOR U696 ( .A(in[1070]), .B(in[750]), .Z(n323) );
  XNOR U697 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U698 ( .A(in[430]), .B(n325), .Z(n1599) );
  XOR U699 ( .A(in[1519]), .B(in[559]), .Z(n327) );
  XNOR U700 ( .A(in[879]), .B(in[239]), .Z(n326) );
  XNOR U701 ( .A(n327), .B(n326), .Z(n328) );
  XNOR U702 ( .A(in[1199]), .B(n328), .Z(n1539) );
  XOR U703 ( .A(n1599), .B(n1539), .Z(n1415) );
  XOR U704 ( .A(in[175]), .B(n1415), .Z(n1512) );
  XOR U705 ( .A(in[975]), .B(in[15]), .Z(n330) );
  XNOR U706 ( .A(in[1295]), .B(in[335]), .Z(n329) );
  XNOR U707 ( .A(n330), .B(n329), .Z(n331) );
  XNOR U708 ( .A(in[655]), .B(n331), .Z(n1430) );
  XOR U709 ( .A(in[144]), .B(in[1424]), .Z(n333) );
  XNOR U710 ( .A(in[1104]), .B(in[784]), .Z(n332) );
  XNOR U711 ( .A(n333), .B(n332), .Z(n334) );
  XOR U712 ( .A(in[464]), .B(n334), .Z(n1396) );
  XNOR U713 ( .A(in[1360]), .B(n4476), .Z(n1920) );
  XOR U714 ( .A(in[1368]), .B(in[728]), .Z(n336) );
  XNOR U715 ( .A(in[88]), .B(in[408]), .Z(n335) );
  XNOR U716 ( .A(n336), .B(n335), .Z(n337) );
  XNOR U717 ( .A(in[1048]), .B(n337), .Z(n1056) );
  XOR U718 ( .A(in[1559]), .B(in[599]), .Z(n339) );
  XNOR U719 ( .A(in[919]), .B(in[279]), .Z(n338) );
  XNOR U720 ( .A(n339), .B(n338), .Z(n340) );
  XNOR U721 ( .A(in[1239]), .B(n340), .Z(n776) );
  XOR U722 ( .A(n1056), .B(n776), .Z(n4258) );
  XOR U723 ( .A(in[984]), .B(n4258), .Z(n1917) );
  NANDN U724 ( .A(n1920), .B(n1917), .Z(n341) );
  XNOR U725 ( .A(n1512), .B(n341), .Z(out[1004]) );
  XOR U726 ( .A(in[1391]), .B(in[111]), .Z(n343) );
  XNOR U727 ( .A(in[1071]), .B(in[751]), .Z(n342) );
  XNOR U728 ( .A(n343), .B(n342), .Z(n344) );
  XNOR U729 ( .A(in[431]), .B(n344), .Z(n1603) );
  XOR U730 ( .A(in[1520]), .B(in[560]), .Z(n346) );
  XNOR U731 ( .A(in[880]), .B(in[240]), .Z(n345) );
  XNOR U732 ( .A(n346), .B(n345), .Z(n347) );
  XNOR U733 ( .A(in[1200]), .B(n347), .Z(n1545) );
  XOR U734 ( .A(n1603), .B(n1545), .Z(n1437) );
  XOR U735 ( .A(in[176]), .B(n1437), .Z(n1516) );
  XOR U736 ( .A(in[976]), .B(in[16]), .Z(n349) );
  XNOR U737 ( .A(in[1296]), .B(in[336]), .Z(n348) );
  XNOR U738 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U739 ( .A(in[656]), .B(n350), .Z(n1432) );
  XOR U740 ( .A(in[145]), .B(in[1425]), .Z(n352) );
  XNOR U741 ( .A(in[1105]), .B(in[785]), .Z(n351) );
  XNOR U742 ( .A(n352), .B(n351), .Z(n353) );
  XOR U743 ( .A(in[465]), .B(n353), .Z(n1400) );
  XNOR U744 ( .A(in[1361]), .B(n4483), .Z(n1924) );
  XOR U745 ( .A(in[1369]), .B(in[729]), .Z(n355) );
  XNOR U746 ( .A(in[89]), .B(in[409]), .Z(n354) );
  XNOR U747 ( .A(n355), .B(n354), .Z(n356) );
  XNOR U748 ( .A(in[1049]), .B(n356), .Z(n1069) );
  XOR U749 ( .A(in[1560]), .B(in[600]), .Z(n358) );
  XNOR U750 ( .A(in[920]), .B(in[280]), .Z(n357) );
  XNOR U751 ( .A(n358), .B(n357), .Z(n359) );
  XNOR U752 ( .A(in[1240]), .B(n359), .Z(n791) );
  XOR U753 ( .A(n1069), .B(n791), .Z(n4259) );
  XOR U754 ( .A(in[985]), .B(n4259), .Z(n1921) );
  NANDN U755 ( .A(n1924), .B(n1921), .Z(n360) );
  XNOR U756 ( .A(n1516), .B(n360), .Z(out[1005]) );
  XOR U757 ( .A(in[1392]), .B(in[112]), .Z(n362) );
  XNOR U758 ( .A(in[1072]), .B(in[752]), .Z(n361) );
  XNOR U759 ( .A(n362), .B(n361), .Z(n363) );
  XNOR U760 ( .A(in[432]), .B(n363), .Z(n1607) );
  XOR U761 ( .A(in[1521]), .B(in[561]), .Z(n365) );
  XNOR U762 ( .A(in[881]), .B(in[241]), .Z(n364) );
  XNOR U763 ( .A(n365), .B(n364), .Z(n366) );
  XNOR U764 ( .A(in[1201]), .B(n366), .Z(n1549) );
  XOR U765 ( .A(n1607), .B(n1549), .Z(n1465) );
  XOR U766 ( .A(in[177]), .B(n1465), .Z(n1520) );
  XOR U767 ( .A(in[17]), .B(in[657]), .Z(n368) );
  XNOR U768 ( .A(in[977]), .B(in[337]), .Z(n367) );
  XNOR U769 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U770 ( .A(in[1297]), .B(n369), .Z(n1434) );
  XOR U771 ( .A(in[1426]), .B(in[466]), .Z(n371) );
  XNOR U772 ( .A(in[786]), .B(in[146]), .Z(n370) );
  XNOR U773 ( .A(n371), .B(n370), .Z(n372) );
  XOR U774 ( .A(in[1106]), .B(n372), .Z(n715) );
  XNOR U775 ( .A(n4486), .B(in[1362]), .Z(n1928) );
  XOR U776 ( .A(in[1370]), .B(in[730]), .Z(n374) );
  XNOR U777 ( .A(in[90]), .B(in[410]), .Z(n373) );
  XNOR U778 ( .A(n374), .B(n373), .Z(n375) );
  XNOR U779 ( .A(in[1050]), .B(n375), .Z(n1084) );
  XOR U780 ( .A(in[1561]), .B(in[601]), .Z(n377) );
  XNOR U781 ( .A(in[921]), .B(in[281]), .Z(n376) );
  XNOR U782 ( .A(n377), .B(n376), .Z(n378) );
  XNOR U783 ( .A(in[1241]), .B(n378), .Z(n817) );
  XOR U784 ( .A(n1084), .B(n817), .Z(n4260) );
  XOR U785 ( .A(in[986]), .B(n4260), .Z(n1925) );
  NANDN U786 ( .A(n1928), .B(n1925), .Z(n379) );
  XNOR U787 ( .A(n1520), .B(n379), .Z(out[1006]) );
  XOR U788 ( .A(in[1393]), .B(in[113]), .Z(n381) );
  XNOR U789 ( .A(in[1073]), .B(in[753]), .Z(n380) );
  XNOR U790 ( .A(n381), .B(n380), .Z(n382) );
  XNOR U791 ( .A(in[433]), .B(n382), .Z(n1611) );
  XOR U792 ( .A(in[1522]), .B(in[562]), .Z(n384) );
  XNOR U793 ( .A(in[882]), .B(in[242]), .Z(n383) );
  XNOR U794 ( .A(n384), .B(n383), .Z(n385) );
  XNOR U795 ( .A(in[1202]), .B(n385), .Z(n1553) );
  XOR U796 ( .A(n1611), .B(n1553), .Z(n1500) );
  XOR U797 ( .A(in[178]), .B(n1500), .Z(n1524) );
  XOR U798 ( .A(in[978]), .B(in[18]), .Z(n387) );
  XNOR U799 ( .A(in[1298]), .B(in[338]), .Z(n386) );
  XNOR U800 ( .A(n387), .B(n386), .Z(n388) );
  XNOR U801 ( .A(in[658]), .B(n388), .Z(n1436) );
  XOR U802 ( .A(in[147]), .B(in[1427]), .Z(n390) );
  XNOR U803 ( .A(in[1107]), .B(in[787]), .Z(n389) );
  XNOR U804 ( .A(n390), .B(n389), .Z(n391) );
  XOR U805 ( .A(in[467]), .B(n391), .Z(n730) );
  XNOR U806 ( .A(in[1363]), .B(n4489), .Z(n1932) );
  XOR U807 ( .A(in[1371]), .B(in[731]), .Z(n393) );
  XNOR U808 ( .A(in[91]), .B(in[411]), .Z(n392) );
  XNOR U809 ( .A(n393), .B(n392), .Z(n394) );
  XNOR U810 ( .A(in[1051]), .B(n394), .Z(n1097) );
  XOR U811 ( .A(in[1562]), .B(in[602]), .Z(n396) );
  XNOR U812 ( .A(in[922]), .B(in[282]), .Z(n395) );
  XNOR U813 ( .A(n396), .B(n395), .Z(n397) );
  XNOR U814 ( .A(in[1242]), .B(n397), .Z(n832) );
  XOR U815 ( .A(n1097), .B(n832), .Z(n4261) );
  XOR U816 ( .A(in[987]), .B(n4261), .Z(n1929) );
  NANDN U817 ( .A(n1932), .B(n1929), .Z(n398) );
  XNOR U818 ( .A(n1524), .B(n398), .Z(out[1007]) );
  XOR U819 ( .A(in[1394]), .B(in[114]), .Z(n400) );
  XNOR U820 ( .A(in[1074]), .B(in[754]), .Z(n399) );
  XNOR U821 ( .A(n400), .B(n399), .Z(n401) );
  XNOR U822 ( .A(in[434]), .B(n401), .Z(n1615) );
  XOR U823 ( .A(in[1523]), .B(in[563]), .Z(n403) );
  XNOR U824 ( .A(in[883]), .B(in[243]), .Z(n402) );
  XNOR U825 ( .A(n403), .B(n402), .Z(n404) );
  XNOR U826 ( .A(in[1203]), .B(n404), .Z(n1557) );
  XOR U827 ( .A(n1615), .B(n1557), .Z(n1542) );
  XOR U828 ( .A(in[179]), .B(n1542), .Z(n1528) );
  XOR U829 ( .A(in[979]), .B(in[19]), .Z(n406) );
  XNOR U830 ( .A(in[1299]), .B(in[339]), .Z(n405) );
  XNOR U831 ( .A(n406), .B(n405), .Z(n407) );
  XNOR U832 ( .A(in[659]), .B(n407), .Z(n1440) );
  XOR U833 ( .A(in[148]), .B(in[1428]), .Z(n409) );
  XNOR U834 ( .A(in[1108]), .B(in[788]), .Z(n408) );
  XNOR U835 ( .A(n409), .B(n408), .Z(n410) );
  XOR U836 ( .A(in[468]), .B(n410), .Z(n745) );
  XNOR U837 ( .A(in[1364]), .B(n4492), .Z(n1936) );
  XOR U838 ( .A(in[1372]), .B(in[732]), .Z(n412) );
  XNOR U839 ( .A(in[92]), .B(in[412]), .Z(n411) );
  XNOR U840 ( .A(n412), .B(n411), .Z(n413) );
  XNOR U841 ( .A(in[1052]), .B(n413), .Z(n1117) );
  XOR U842 ( .A(in[1563]), .B(in[603]), .Z(n415) );
  XNOR U843 ( .A(in[923]), .B(in[283]), .Z(n414) );
  XNOR U844 ( .A(n415), .B(n414), .Z(n416) );
  XNOR U845 ( .A(in[1243]), .B(n416), .Z(n847) );
  XOR U846 ( .A(n1117), .B(n847), .Z(n4264) );
  XOR U847 ( .A(in[988]), .B(n4264), .Z(n1933) );
  NANDN U848 ( .A(n1936), .B(n1933), .Z(n417) );
  XNOR U849 ( .A(n1528), .B(n417), .Z(out[1008]) );
  XOR U850 ( .A(in[1395]), .B(in[115]), .Z(n419) );
  XNOR U851 ( .A(in[1075]), .B(in[755]), .Z(n418) );
  XNOR U852 ( .A(n419), .B(n418), .Z(n420) );
  XNOR U853 ( .A(in[435]), .B(n420), .Z(n1619) );
  XOR U854 ( .A(in[1524]), .B(in[564]), .Z(n422) );
  XNOR U855 ( .A(in[884]), .B(in[244]), .Z(n421) );
  XNOR U856 ( .A(n422), .B(n421), .Z(n423) );
  XNOR U857 ( .A(in[1204]), .B(n423), .Z(n1561) );
  XOR U858 ( .A(n1619), .B(n1561), .Z(n1584) );
  XOR U859 ( .A(in[180]), .B(n1584), .Z(n1532) );
  XOR U860 ( .A(in[149]), .B(in[1429]), .Z(n425) );
  XNOR U861 ( .A(in[1109]), .B(in[789]), .Z(n424) );
  XNOR U862 ( .A(n425), .B(n424), .Z(n426) );
  XNOR U863 ( .A(in[469]), .B(n426), .Z(n760) );
  XOR U864 ( .A(in[340]), .B(in[660]), .Z(n428) );
  XNOR U865 ( .A(in[20]), .B(in[1300]), .Z(n427) );
  XNOR U866 ( .A(n428), .B(n427), .Z(n429) );
  XOR U867 ( .A(in[980]), .B(n429), .Z(n1442) );
  XNOR U868 ( .A(in[1365]), .B(n4495), .Z(n1940) );
  XOR U869 ( .A(in[1373]), .B(in[733]), .Z(n431) );
  XNOR U870 ( .A(in[93]), .B(in[413]), .Z(n430) );
  XNOR U871 ( .A(n431), .B(n430), .Z(n432) );
  XNOR U872 ( .A(in[1053]), .B(n432), .Z(n1130) );
  XOR U873 ( .A(in[1564]), .B(in[604]), .Z(n434) );
  XNOR U874 ( .A(in[924]), .B(in[284]), .Z(n433) );
  XNOR U875 ( .A(n434), .B(n433), .Z(n435) );
  XNOR U876 ( .A(in[1244]), .B(n435), .Z(n862) );
  XOR U877 ( .A(n1130), .B(n862), .Z(n4265) );
  XOR U878 ( .A(in[989]), .B(n4265), .Z(n1937) );
  NANDN U879 ( .A(n1940), .B(n1937), .Z(n436) );
  XNOR U880 ( .A(n1532), .B(n436), .Z(out[1009]) );
  XOR U881 ( .A(in[1339]), .B(in[59]), .Z(n438) );
  XNOR U882 ( .A(in[699]), .B(in[379]), .Z(n437) );
  XNOR U883 ( .A(n438), .B(n437), .Z(n439) );
  XNOR U884 ( .A(in[1019]), .B(n439), .Z(n1088) );
  XOR U885 ( .A(in[1530]), .B(in[570]), .Z(n441) );
  XNOR U886 ( .A(in[1210]), .B(in[250]), .Z(n440) );
  XNOR U887 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U888 ( .A(in[890]), .B(n442), .Z(n554) );
  XOR U889 ( .A(n1088), .B(n554), .Z(n3955) );
  XOR U890 ( .A(in[635]), .B(n3955), .Z(n2706) );
  IV U891 ( .A(n2706), .Z(n2792) );
  XOR U892 ( .A(in[161]), .B(in[1441]), .Z(n444) );
  XNOR U893 ( .A(in[801]), .B(in[1121]), .Z(n443) );
  XNOR U894 ( .A(n444), .B(n443), .Z(n445) );
  XNOR U895 ( .A(in[481]), .B(n445), .Z(n681) );
  XOR U896 ( .A(in[1570]), .B(in[610]), .Z(n447) );
  XNOR U897 ( .A(in[930]), .B(in[290]), .Z(n446) );
  XNOR U898 ( .A(n447), .B(n446), .Z(n448) );
  XOR U899 ( .A(in[1250]), .B(n448), .Z(n564) );
  XOR U900 ( .A(in[226]), .B(n4051), .Z(n3117) );
  XOR U901 ( .A(in[1061]), .B(in[421]), .Z(n450) );
  XNOR U902 ( .A(in[741]), .B(in[1381]), .Z(n449) );
  XNOR U903 ( .A(n450), .B(n449), .Z(n451) );
  XNOR U904 ( .A(in[101]), .B(n451), .Z(n600) );
  XOR U905 ( .A(in[1510]), .B(in[550]), .Z(n453) );
  XNOR U906 ( .A(in[870]), .B(in[230]), .Z(n452) );
  XNOR U907 ( .A(n453), .B(n452), .Z(n454) );
  XNOR U908 ( .A(in[1190]), .B(n454), .Z(n1503) );
  XNOR U909 ( .A(n600), .B(n1503), .Z(n4091) );
  IV U910 ( .A(n4091), .Z(n1243) );
  XOR U911 ( .A(in[1446]), .B(n1243), .Z(n3114) );
  NANDN U912 ( .A(n3117), .B(n3114), .Z(n455) );
  XOR U913 ( .A(n2792), .B(n455), .Z(out[100]) );
  XOR U914 ( .A(in[1396]), .B(in[116]), .Z(n457) );
  XNOR U915 ( .A(in[1076]), .B(in[756]), .Z(n456) );
  XNOR U916 ( .A(n457), .B(n456), .Z(n458) );
  XNOR U917 ( .A(in[436]), .B(n458), .Z(n1624) );
  XOR U918 ( .A(in[1525]), .B(in[565]), .Z(n460) );
  XNOR U919 ( .A(in[885]), .B(in[245]), .Z(n459) );
  XNOR U920 ( .A(n460), .B(n459), .Z(n461) );
  XNOR U921 ( .A(in[1205]), .B(n461), .Z(n1565) );
  XOR U922 ( .A(n1624), .B(n1565), .Z(n4155) );
  XOR U923 ( .A(in[181]), .B(n4155), .Z(n1536) );
  XOR U924 ( .A(in[341]), .B(in[661]), .Z(n463) );
  XNOR U925 ( .A(in[21]), .B(in[1301]), .Z(n462) );
  XNOR U926 ( .A(n463), .B(n462), .Z(n464) );
  XNOR U927 ( .A(in[981]), .B(n464), .Z(n1444) );
  XOR U928 ( .A(in[150]), .B(in[1430]), .Z(n466) );
  XNOR U929 ( .A(in[1110]), .B(in[790]), .Z(n465) );
  XNOR U930 ( .A(n466), .B(n465), .Z(n467) );
  XOR U931 ( .A(in[470]), .B(n467), .Z(n775) );
  XNOR U932 ( .A(in[1366]), .B(n4498), .Z(n1944) );
  XOR U933 ( .A(in[1374]), .B(in[734]), .Z(n469) );
  XNOR U934 ( .A(in[94]), .B(in[414]), .Z(n468) );
  XNOR U935 ( .A(n469), .B(n468), .Z(n470) );
  XNOR U936 ( .A(in[1054]), .B(n470), .Z(n1143) );
  XOR U937 ( .A(in[1565]), .B(in[605]), .Z(n472) );
  XNOR U938 ( .A(in[925]), .B(in[285]), .Z(n471) );
  XNOR U939 ( .A(n472), .B(n471), .Z(n473) );
  XNOR U940 ( .A(in[1245]), .B(n473), .Z(n877) );
  XOR U941 ( .A(n1143), .B(n877), .Z(n4266) );
  XOR U942 ( .A(in[990]), .B(n4266), .Z(n1941) );
  NANDN U943 ( .A(n1944), .B(n1941), .Z(n474) );
  XNOR U944 ( .A(n1536), .B(n474), .Z(out[1010]) );
  XOR U945 ( .A(in[1526]), .B(in[566]), .Z(n476) );
  XNOR U946 ( .A(in[886]), .B(in[246]), .Z(n475) );
  XNOR U947 ( .A(n476), .B(n475), .Z(n477) );
  XNOR U948 ( .A(in[1206]), .B(n477), .Z(n1569) );
  XOR U949 ( .A(in[1397]), .B(in[117]), .Z(n479) );
  XNOR U950 ( .A(in[1077]), .B(in[757]), .Z(n478) );
  XNOR U951 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U952 ( .A(in[437]), .B(n480), .Z(n1628) );
  XOR U953 ( .A(n1569), .B(n1628), .Z(n4165) );
  XOR U954 ( .A(in[182]), .B(n4165), .Z(n1540) );
  XOR U955 ( .A(in[151]), .B(in[1431]), .Z(n482) );
  XNOR U956 ( .A(in[1111]), .B(in[791]), .Z(n481) );
  XNOR U957 ( .A(n482), .B(n481), .Z(n483) );
  XNOR U958 ( .A(in[471]), .B(n483), .Z(n790) );
  XOR U959 ( .A(in[342]), .B(in[662]), .Z(n485) );
  XNOR U960 ( .A(in[22]), .B(in[1302]), .Z(n484) );
  XNOR U961 ( .A(n485), .B(n484), .Z(n486) );
  XOR U962 ( .A(in[982]), .B(n486), .Z(n1446) );
  XNOR U963 ( .A(in[1367]), .B(n4501), .Z(n1948) );
  XOR U964 ( .A(in[1375]), .B(in[735]), .Z(n488) );
  XNOR U965 ( .A(in[95]), .B(in[415]), .Z(n487) );
  XNOR U966 ( .A(n488), .B(n487), .Z(n489) );
  XNOR U967 ( .A(in[1055]), .B(n489), .Z(n1156) );
  XOR U968 ( .A(in[1566]), .B(in[606]), .Z(n491) );
  XNOR U969 ( .A(in[926]), .B(in[286]), .Z(n490) );
  XNOR U970 ( .A(n491), .B(n490), .Z(n492) );
  XNOR U971 ( .A(in[1246]), .B(n492), .Z(n892) );
  XOR U972 ( .A(n1156), .B(n892), .Z(n4267) );
  XOR U973 ( .A(in[991]), .B(n4267), .Z(n1945) );
  NANDN U974 ( .A(n1948), .B(n1945), .Z(n493) );
  XNOR U975 ( .A(n1540), .B(n493), .Z(out[1011]) );
  XOR U976 ( .A(in[1527]), .B(in[567]), .Z(n495) );
  XNOR U977 ( .A(in[887]), .B(in[247]), .Z(n494) );
  XNOR U978 ( .A(n495), .B(n494), .Z(n496) );
  XNOR U979 ( .A(in[1207]), .B(n496), .Z(n1573) );
  XOR U980 ( .A(in[1398]), .B(in[118]), .Z(n498) );
  XNOR U981 ( .A(in[1078]), .B(in[758]), .Z(n497) );
  XNOR U982 ( .A(n498), .B(n497), .Z(n499) );
  XNOR U983 ( .A(in[438]), .B(n499), .Z(n1632) );
  XOR U984 ( .A(n1573), .B(n1632), .Z(n4169) );
  XOR U985 ( .A(in[183]), .B(n4169), .Z(n1546) );
  XOR U986 ( .A(in[152]), .B(in[1432]), .Z(n501) );
  XNOR U987 ( .A(in[1112]), .B(in[792]), .Z(n500) );
  XNOR U988 ( .A(n501), .B(n500), .Z(n502) );
  XNOR U989 ( .A(in[472]), .B(n502), .Z(n816) );
  XOR U990 ( .A(in[343]), .B(in[663]), .Z(n504) );
  XNOR U991 ( .A(in[23]), .B(in[1303]), .Z(n503) );
  XNOR U992 ( .A(n504), .B(n503), .Z(n505) );
  XOR U993 ( .A(in[983]), .B(n505), .Z(n1448) );
  XNOR U994 ( .A(in[1368]), .B(n4504), .Z(n1952) );
  XOR U995 ( .A(in[1376]), .B(in[736]), .Z(n507) );
  XNOR U996 ( .A(in[96]), .B(in[416]), .Z(n506) );
  XNOR U997 ( .A(n507), .B(n506), .Z(n508) );
  XNOR U998 ( .A(in[1056]), .B(n508), .Z(n1171) );
  XOR U999 ( .A(in[1567]), .B(in[607]), .Z(n510) );
  XNOR U1000 ( .A(in[927]), .B(in[287]), .Z(n509) );
  XNOR U1001 ( .A(n510), .B(n509), .Z(n511) );
  XNOR U1002 ( .A(in[1247]), .B(n511), .Z(n907) );
  XOR U1003 ( .A(n1171), .B(n907), .Z(n4270) );
  XOR U1004 ( .A(in[992]), .B(n4270), .Z(n1949) );
  NANDN U1005 ( .A(n1952), .B(n1949), .Z(n512) );
  XNOR U1006 ( .A(n1546), .B(n512), .Z(out[1012]) );
  XOR U1007 ( .A(in[1528]), .B(in[568]), .Z(n514) );
  XNOR U1008 ( .A(in[888]), .B(in[248]), .Z(n513) );
  XNOR U1009 ( .A(n514), .B(n513), .Z(n515) );
  XNOR U1010 ( .A(in[1208]), .B(n515), .Z(n1577) );
  XOR U1011 ( .A(in[1399]), .B(in[119]), .Z(n517) );
  XNOR U1012 ( .A(in[1079]), .B(in[759]), .Z(n516) );
  XNOR U1013 ( .A(n517), .B(n516), .Z(n518) );
  XNOR U1014 ( .A(in[439]), .B(n518), .Z(n1636) );
  XOR U1015 ( .A(n1577), .B(n1636), .Z(n4173) );
  XOR U1016 ( .A(in[184]), .B(n4173), .Z(n1550) );
  XOR U1017 ( .A(in[153]), .B(in[1433]), .Z(n520) );
  XNOR U1018 ( .A(in[1113]), .B(in[793]), .Z(n519) );
  XNOR U1019 ( .A(n520), .B(n519), .Z(n521) );
  XNOR U1020 ( .A(in[473]), .B(n521), .Z(n831) );
  XOR U1021 ( .A(in[344]), .B(in[664]), .Z(n523) );
  XNOR U1022 ( .A(in[24]), .B(in[1304]), .Z(n522) );
  XNOR U1023 ( .A(n523), .B(n522), .Z(n524) );
  XOR U1024 ( .A(in[984]), .B(n524), .Z(n1450) );
  XNOR U1025 ( .A(in[1369]), .B(n4507), .Z(n1956) );
  XOR U1026 ( .A(in[1377]), .B(in[737]), .Z(n526) );
  XNOR U1027 ( .A(in[97]), .B(in[417]), .Z(n525) );
  XNOR U1028 ( .A(n526), .B(n525), .Z(n527) );
  XNOR U1029 ( .A(in[1057]), .B(n527), .Z(n1186) );
  XOR U1030 ( .A(in[1568]), .B(in[608]), .Z(n529) );
  XNOR U1031 ( .A(in[928]), .B(in[288]), .Z(n528) );
  XNOR U1032 ( .A(n529), .B(n528), .Z(n530) );
  XNOR U1033 ( .A(in[1248]), .B(n530), .Z(n922) );
  XOR U1034 ( .A(n1186), .B(n922), .Z(n4273) );
  XOR U1035 ( .A(in[993]), .B(n4273), .Z(n1953) );
  NANDN U1036 ( .A(n1956), .B(n1953), .Z(n531) );
  XNOR U1037 ( .A(n1550), .B(n531), .Z(out[1013]) );
  XOR U1038 ( .A(in[1529]), .B(in[569]), .Z(n533) );
  XNOR U1039 ( .A(in[889]), .B(in[249]), .Z(n532) );
  XNOR U1040 ( .A(n533), .B(n532), .Z(n534) );
  XNOR U1041 ( .A(in[1209]), .B(n534), .Z(n1581) );
  XOR U1042 ( .A(in[1400]), .B(in[120]), .Z(n536) );
  XNOR U1043 ( .A(in[1080]), .B(in[760]), .Z(n535) );
  XNOR U1044 ( .A(n536), .B(n535), .Z(n537) );
  XNOR U1045 ( .A(in[440]), .B(n537), .Z(n1640) );
  XOR U1046 ( .A(n1581), .B(n1640), .Z(n4177) );
  XOR U1047 ( .A(in[185]), .B(n4177), .Z(n1554) );
  XOR U1048 ( .A(in[154]), .B(in[1434]), .Z(n539) );
  XNOR U1049 ( .A(in[1114]), .B(in[794]), .Z(n538) );
  XNOR U1050 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U1051 ( .A(in[474]), .B(n540), .Z(n846) );
  XOR U1052 ( .A(in[345]), .B(in[665]), .Z(n542) );
  XNOR U1053 ( .A(in[25]), .B(in[1305]), .Z(n541) );
  XNOR U1054 ( .A(n542), .B(n541), .Z(n543) );
  XOR U1055 ( .A(in[985]), .B(n543), .Z(n1454) );
  XNOR U1056 ( .A(in[1370]), .B(n4510), .Z(n1962) );
  XOR U1057 ( .A(in[1569]), .B(in[609]), .Z(n545) );
  XNOR U1058 ( .A(in[929]), .B(in[289]), .Z(n544) );
  XNOR U1059 ( .A(n545), .B(n544), .Z(n546) );
  XNOR U1060 ( .A(in[1249]), .B(n546), .Z(n937) );
  XOR U1061 ( .A(in[1378]), .B(in[738]), .Z(n548) );
  XNOR U1062 ( .A(in[98]), .B(in[418]), .Z(n547) );
  XNOR U1063 ( .A(n548), .B(n547), .Z(n549) );
  XNOR U1064 ( .A(in[1058]), .B(n549), .Z(n1201) );
  XOR U1065 ( .A(n937), .B(n1201), .Z(n4276) );
  XOR U1066 ( .A(in[994]), .B(n4276), .Z(n1959) );
  NANDN U1067 ( .A(n1962), .B(n1959), .Z(n550) );
  XNOR U1068 ( .A(n1554), .B(n550), .Z(out[1014]) );
  XOR U1069 ( .A(in[1401]), .B(in[121]), .Z(n552) );
  XNOR U1070 ( .A(in[1081]), .B(in[761]), .Z(n551) );
  XNOR U1071 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U1072 ( .A(in[441]), .B(n553), .Z(n1644) );
  XOR U1073 ( .A(n554), .B(n1644), .Z(n1792) );
  XOR U1074 ( .A(in[186]), .B(n1792), .Z(n1558) );
  XOR U1075 ( .A(in[155]), .B(in[1435]), .Z(n556) );
  XNOR U1076 ( .A(in[1115]), .B(in[795]), .Z(n555) );
  XNOR U1077 ( .A(n556), .B(n555), .Z(n557) );
  XNOR U1078 ( .A(in[475]), .B(n557), .Z(n861) );
  XOR U1079 ( .A(in[346]), .B(in[666]), .Z(n559) );
  XNOR U1080 ( .A(in[26]), .B(in[1306]), .Z(n558) );
  XNOR U1081 ( .A(n559), .B(n558), .Z(n560) );
  XOR U1082 ( .A(in[986]), .B(n560), .Z(n1456) );
  IV U1083 ( .A(n4517), .Z(n2742) );
  XOR U1084 ( .A(in[1371]), .B(n2742), .Z(n1359) );
  IV U1085 ( .A(n1359), .Z(n1966) );
  XOR U1086 ( .A(in[1379]), .B(in[739]), .Z(n562) );
  XNOR U1087 ( .A(in[99]), .B(in[419]), .Z(n561) );
  XNOR U1088 ( .A(n562), .B(n561), .Z(n563) );
  XOR U1089 ( .A(in[1059]), .B(n563), .Z(n1216) );
  XNOR U1090 ( .A(n564), .B(n1216), .Z(n4279) );
  XNOR U1091 ( .A(in[995]), .B(n4279), .Z(n1963) );
  NANDN U1092 ( .A(n1966), .B(n1963), .Z(n565) );
  XNOR U1093 ( .A(n1558), .B(n565), .Z(out[1015]) );
  XOR U1094 ( .A(in[1402]), .B(in[122]), .Z(n567) );
  XNOR U1095 ( .A(in[1082]), .B(in[762]), .Z(n566) );
  XNOR U1096 ( .A(n567), .B(n566), .Z(n568) );
  XNOR U1097 ( .A(in[442]), .B(n568), .Z(n1648) );
  XOR U1098 ( .A(in[1531]), .B(in[571]), .Z(n570) );
  XNOR U1099 ( .A(in[1211]), .B(in[251]), .Z(n569) );
  XNOR U1100 ( .A(n570), .B(n569), .Z(n571) );
  XNOR U1101 ( .A(in[891]), .B(n571), .Z(n643) );
  XOR U1102 ( .A(n1648), .B(n643), .Z(n1818) );
  XOR U1103 ( .A(in[187]), .B(n1818), .Z(n1562) );
  XOR U1104 ( .A(in[156]), .B(in[1436]), .Z(n573) );
  XNOR U1105 ( .A(in[1116]), .B(in[796]), .Z(n572) );
  XNOR U1106 ( .A(n573), .B(n572), .Z(n574) );
  XNOR U1107 ( .A(in[476]), .B(n574), .Z(n876) );
  XOR U1108 ( .A(in[347]), .B(in[667]), .Z(n576) );
  XNOR U1109 ( .A(in[27]), .B(in[1307]), .Z(n575) );
  XNOR U1110 ( .A(n576), .B(n575), .Z(n577) );
  XOR U1111 ( .A(in[987]), .B(n577), .Z(n1458) );
  IV U1112 ( .A(n4520), .Z(n2759) );
  XOR U1113 ( .A(in[1372]), .B(n2759), .Z(n1369) );
  IV U1114 ( .A(n1369), .Z(n1970) );
  XOR U1115 ( .A(in[1060]), .B(in[420]), .Z(n579) );
  XNOR U1116 ( .A(in[740]), .B(in[1380]), .Z(n578) );
  XNOR U1117 ( .A(n579), .B(n578), .Z(n580) );
  XNOR U1118 ( .A(in[100]), .B(n580), .Z(n1231) );
  XOR U1119 ( .A(in[1571]), .B(in[611]), .Z(n582) );
  XNOR U1120 ( .A(in[931]), .B(in[291]), .Z(n581) );
  XNOR U1121 ( .A(n582), .B(n581), .Z(n583) );
  XNOR U1122 ( .A(in[1251]), .B(n583), .Z(n647) );
  XOR U1123 ( .A(n1231), .B(n647), .Z(n4282) );
  XOR U1124 ( .A(in[996]), .B(n4282), .Z(n1967) );
  NANDN U1125 ( .A(n1970), .B(n1967), .Z(n584) );
  XNOR U1126 ( .A(n1562), .B(n584), .Z(out[1016]) );
  XOR U1127 ( .A(in[1403]), .B(in[123]), .Z(n586) );
  XNOR U1128 ( .A(in[1083]), .B(in[763]), .Z(n585) );
  XNOR U1129 ( .A(n586), .B(n585), .Z(n587) );
  XNOR U1130 ( .A(in[443]), .B(n587), .Z(n1652) );
  XOR U1131 ( .A(in[1532]), .B(in[572]), .Z(n589) );
  XNOR U1132 ( .A(in[1212]), .B(in[252]), .Z(n588) );
  XNOR U1133 ( .A(n589), .B(n588), .Z(n590) );
  XNOR U1134 ( .A(in[892]), .B(n590), .Z(n808) );
  XOR U1135 ( .A(n1652), .B(n808), .Z(n1841) );
  XOR U1136 ( .A(in[188]), .B(n1841), .Z(n1566) );
  XOR U1137 ( .A(in[157]), .B(in[1437]), .Z(n592) );
  XNOR U1138 ( .A(in[1117]), .B(in[797]), .Z(n591) );
  XNOR U1139 ( .A(n592), .B(n591), .Z(n593) );
  XNOR U1140 ( .A(in[477]), .B(n593), .Z(n891) );
  XOR U1141 ( .A(in[348]), .B(in[668]), .Z(n595) );
  XNOR U1142 ( .A(in[28]), .B(in[1308]), .Z(n594) );
  XNOR U1143 ( .A(n595), .B(n594), .Z(n596) );
  XOR U1144 ( .A(in[988]), .B(n596), .Z(n1462) );
  IV U1145 ( .A(n4523), .Z(n2776) );
  XOR U1146 ( .A(in[1373]), .B(n2776), .Z(n1375) );
  IV U1147 ( .A(n1375), .Z(n1974) );
  XOR U1148 ( .A(in[1572]), .B(in[612]), .Z(n598) );
  XNOR U1149 ( .A(in[932]), .B(in[292]), .Z(n597) );
  XNOR U1150 ( .A(n598), .B(n597), .Z(n599) );
  XNOR U1151 ( .A(in[1252]), .B(n599), .Z(n810) );
  XOR U1152 ( .A(n600), .B(n810), .Z(n4284) );
  XOR U1153 ( .A(in[997]), .B(n4284), .Z(n1971) );
  NANDN U1154 ( .A(n1974), .B(n1971), .Z(n601) );
  XNOR U1155 ( .A(n1566), .B(n601), .Z(out[1017]) );
  XOR U1156 ( .A(in[1404]), .B(in[124]), .Z(n603) );
  XNOR U1157 ( .A(in[1084]), .B(in[764]), .Z(n602) );
  XNOR U1158 ( .A(n603), .B(n602), .Z(n604) );
  XNOR U1159 ( .A(in[444]), .B(n604), .Z(n1656) );
  XOR U1160 ( .A(in[1533]), .B(in[573]), .Z(n606) );
  XNOR U1161 ( .A(in[1213]), .B(in[253]), .Z(n605) );
  XNOR U1162 ( .A(n606), .B(n605), .Z(n607) );
  XNOR U1163 ( .A(in[893]), .B(n607), .Z(n967) );
  XOR U1164 ( .A(n1656), .B(n967), .Z(n1863) );
  XOR U1165 ( .A(in[189]), .B(n1863), .Z(n1570) );
  XOR U1166 ( .A(in[158]), .B(in[1438]), .Z(n609) );
  XNOR U1167 ( .A(in[1118]), .B(in[798]), .Z(n608) );
  XNOR U1168 ( .A(n609), .B(n608), .Z(n610) );
  XNOR U1169 ( .A(in[478]), .B(n610), .Z(n906) );
  XOR U1170 ( .A(in[349]), .B(in[669]), .Z(n612) );
  XNOR U1171 ( .A(in[29]), .B(in[1309]), .Z(n611) );
  XNOR U1172 ( .A(n612), .B(n611), .Z(n613) );
  XOR U1173 ( .A(in[989]), .B(n613), .Z(n1468) );
  XNOR U1174 ( .A(in[1374]), .B(n4526), .Z(n1978) );
  XOR U1175 ( .A(in[1062]), .B(in[422]), .Z(n615) );
  XNOR U1176 ( .A(in[742]), .B(in[1382]), .Z(n614) );
  XNOR U1177 ( .A(n615), .B(n614), .Z(n616) );
  XNOR U1178 ( .A(in[102]), .B(n616), .Z(n651) );
  XOR U1179 ( .A(in[1573]), .B(in[613]), .Z(n618) );
  XNOR U1180 ( .A(in[933]), .B(in[293]), .Z(n617) );
  XNOR U1181 ( .A(n618), .B(n617), .Z(n619) );
  XNOR U1182 ( .A(in[1253]), .B(n619), .Z(n969) );
  XOR U1183 ( .A(n651), .B(n969), .Z(n4290) );
  XOR U1184 ( .A(in[998]), .B(n4290), .Z(n1975) );
  NANDN U1185 ( .A(n1978), .B(n1975), .Z(n620) );
  XNOR U1186 ( .A(n1570), .B(n620), .Z(out[1018]) );
  XOR U1187 ( .A(in[1405]), .B(in[125]), .Z(n622) );
  XNOR U1188 ( .A(in[1085]), .B(in[765]), .Z(n621) );
  XNOR U1189 ( .A(n622), .B(n621), .Z(n623) );
  XNOR U1190 ( .A(in[445]), .B(n623), .Z(n1660) );
  XOR U1191 ( .A(in[1534]), .B(in[894]), .Z(n625) );
  XNOR U1192 ( .A(in[574]), .B(in[1214]), .Z(n624) );
  XNOR U1193 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1194 ( .A(in[254]), .B(n626), .Z(n1104) );
  XOR U1195 ( .A(n1660), .B(n1104), .Z(n1885) );
  XOR U1196 ( .A(in[190]), .B(n1885), .Z(n1574) );
  XOR U1197 ( .A(in[1439]), .B(in[479]), .Z(n628) );
  XNOR U1198 ( .A(in[799]), .B(in[159]), .Z(n627) );
  XNOR U1199 ( .A(n628), .B(n627), .Z(n629) );
  XNOR U1200 ( .A(in[1119]), .B(n629), .Z(n921) );
  XOR U1201 ( .A(in[350]), .B(in[670]), .Z(n631) );
  XNOR U1202 ( .A(in[30]), .B(in[1310]), .Z(n630) );
  XNOR U1203 ( .A(n631), .B(n630), .Z(n632) );
  XOR U1204 ( .A(in[990]), .B(n632), .Z(n1472) );
  XNOR U1205 ( .A(in[1375]), .B(n4530), .Z(n1982) );
  XOR U1206 ( .A(in[1063]), .B(in[423]), .Z(n634) );
  XNOR U1207 ( .A(in[743]), .B(in[1383]), .Z(n633) );
  XNOR U1208 ( .A(n634), .B(n633), .Z(n635) );
  XNOR U1209 ( .A(in[103]), .B(n635), .Z(n814) );
  XOR U1210 ( .A(in[1574]), .B(in[614]), .Z(n637) );
  XNOR U1211 ( .A(in[934]), .B(in[294]), .Z(n636) );
  XNOR U1212 ( .A(n637), .B(n636), .Z(n638) );
  XNOR U1213 ( .A(in[1254]), .B(n638), .Z(n1013) );
  XOR U1214 ( .A(n814), .B(n1013), .Z(n4292) );
  XOR U1215 ( .A(in[999]), .B(n4292), .Z(n1979) );
  NANDN U1216 ( .A(n1982), .B(n1979), .Z(n639) );
  XNOR U1217 ( .A(n1574), .B(n639), .Z(out[1019]) );
  XOR U1218 ( .A(in[1340]), .B(in[60]), .Z(n641) );
  XNOR U1219 ( .A(in[700]), .B(in[380]), .Z(n640) );
  XNOR U1220 ( .A(n641), .B(n640), .Z(n642) );
  XNOR U1221 ( .A(in[1020]), .B(n642), .Z(n1098) );
  XOR U1222 ( .A(n643), .B(n1098), .Z(n3959) );
  XOR U1223 ( .A(in[636]), .B(n3959), .Z(n2708) );
  IV U1224 ( .A(n2708), .Z(n2794) );
  XOR U1225 ( .A(in[162]), .B(in[1442]), .Z(n645) );
  XNOR U1226 ( .A(in[802]), .B(in[1122]), .Z(n644) );
  XNOR U1227 ( .A(n645), .B(n644), .Z(n646) );
  XOR U1228 ( .A(in[482]), .B(n646), .Z(n698) );
  XOR U1229 ( .A(n647), .B(n698), .Z(n3400) );
  IV U1230 ( .A(n3400), .Z(n4055) );
  XOR U1231 ( .A(in[227]), .B(n4055), .Z(n3141) );
  XOR U1232 ( .A(in[1511]), .B(in[551]), .Z(n649) );
  XNOR U1233 ( .A(in[871]), .B(in[231]), .Z(n648) );
  XNOR U1234 ( .A(n649), .B(n648), .Z(n650) );
  XNOR U1235 ( .A(in[1191]), .B(n650), .Z(n1507) );
  XNOR U1236 ( .A(n651), .B(n1507), .Z(n4095) );
  IV U1237 ( .A(n4095), .Z(n1258) );
  XOR U1238 ( .A(in[1447]), .B(n1258), .Z(n3138) );
  NANDN U1239 ( .A(n3141), .B(n3138), .Z(n652) );
  XOR U1240 ( .A(n2794), .B(n652), .Z(out[101]) );
  XOR U1241 ( .A(in[1406]), .B(in[126]), .Z(n654) );
  XNOR U1242 ( .A(in[1086]), .B(in[766]), .Z(n653) );
  XNOR U1243 ( .A(n654), .B(n653), .Z(n655) );
  XNOR U1244 ( .A(in[446]), .B(n655), .Z(n1665) );
  XOR U1245 ( .A(in[1535]), .B(in[575]), .Z(n657) );
  XNOR U1246 ( .A(in[895]), .B(in[255]), .Z(n656) );
  XNOR U1247 ( .A(n657), .B(n656), .Z(n658) );
  XNOR U1248 ( .A(in[1215]), .B(n658), .Z(n1252) );
  XOR U1249 ( .A(n1665), .B(n1252), .Z(n1915) );
  XOR U1250 ( .A(in[191]), .B(n1915), .Z(n1578) );
  XOR U1251 ( .A(in[1440]), .B(in[480]), .Z(n660) );
  XNOR U1252 ( .A(in[800]), .B(in[160]), .Z(n659) );
  XNOR U1253 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U1254 ( .A(in[1120]), .B(n661), .Z(n936) );
  XOR U1255 ( .A(in[351]), .B(in[671]), .Z(n663) );
  XNOR U1256 ( .A(in[31]), .B(in[1311]), .Z(n662) );
  XNOR U1257 ( .A(n663), .B(n662), .Z(n664) );
  XOR U1258 ( .A(in[991]), .B(n664), .Z(n1476) );
  XNOR U1259 ( .A(in[1376]), .B(n4534), .Z(n1986) );
  XOR U1260 ( .A(in[1064]), .B(in[424]), .Z(n666) );
  XNOR U1261 ( .A(in[744]), .B(in[1384]), .Z(n665) );
  XNOR U1262 ( .A(n666), .B(n665), .Z(n667) );
  XNOR U1263 ( .A(in[104]), .B(n667), .Z(n973) );
  XOR U1264 ( .A(in[1575]), .B(in[615]), .Z(n669) );
  XNOR U1265 ( .A(in[935]), .B(in[295]), .Z(n668) );
  XNOR U1266 ( .A(n669), .B(n668), .Z(n670) );
  XNOR U1267 ( .A(in[1255]), .B(n670), .Z(n1026) );
  XOR U1268 ( .A(n973), .B(n1026), .Z(n4294) );
  XOR U1269 ( .A(in[1000]), .B(n4294), .Z(n1983) );
  NANDN U1270 ( .A(n1986), .B(n1983), .Z(n671) );
  XNOR U1271 ( .A(n1578), .B(n671), .Z(out[1020]) );
  XOR U1272 ( .A(in[1407]), .B(in[127]), .Z(n673) );
  XNOR U1273 ( .A(in[1087]), .B(in[767]), .Z(n672) );
  XNOR U1274 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U1275 ( .A(in[447]), .B(n674), .Z(n1668) );
  XOR U1276 ( .A(in[1472]), .B(in[512]), .Z(n676) );
  XNOR U1277 ( .A(in[832]), .B(in[192]), .Z(n675) );
  XNOR U1278 ( .A(n676), .B(n675), .Z(n677) );
  XNOR U1279 ( .A(in[1152]), .B(n677), .Z(n1317) );
  XOR U1280 ( .A(n1668), .B(n1317), .Z(n1957) );
  XOR U1281 ( .A(in[128]), .B(n1957), .Z(n1582) );
  XOR U1282 ( .A(in[352]), .B(in[672]), .Z(n679) );
  XNOR U1283 ( .A(in[32]), .B(in[1312]), .Z(n678) );
  XNOR U1284 ( .A(n679), .B(n678), .Z(n680) );
  XOR U1285 ( .A(in[992]), .B(n680), .Z(n1478) );
  XNOR U1286 ( .A(in[1377]), .B(n4538), .Z(n1990) );
  XOR U1287 ( .A(in[1065]), .B(in[425]), .Z(n683) );
  XNOR U1288 ( .A(in[745]), .B(in[1385]), .Z(n682) );
  XNOR U1289 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U1290 ( .A(in[105]), .B(n684), .Z(n1108) );
  XOR U1291 ( .A(in[1576]), .B(in[616]), .Z(n686) );
  XNOR U1292 ( .A(in[936]), .B(in[296]), .Z(n685) );
  XNOR U1293 ( .A(n686), .B(n685), .Z(n687) );
  XNOR U1294 ( .A(in[1256]), .B(n687), .Z(n1039) );
  XOR U1295 ( .A(n1108), .B(n1039), .Z(n4296) );
  XOR U1296 ( .A(in[1001]), .B(n4296), .Z(n1987) );
  NANDN U1297 ( .A(n1990), .B(n1987), .Z(n688) );
  XNOR U1298 ( .A(n1582), .B(n688), .Z(out[1021]) );
  XOR U1299 ( .A(in[1344]), .B(in[64]), .Z(n690) );
  XNOR U1300 ( .A(in[1024]), .B(in[384]), .Z(n689) );
  XNOR U1301 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U1302 ( .A(in[704]), .B(n691), .Z(n1673) );
  XOR U1303 ( .A(in[1473]), .B(in[513]), .Z(n693) );
  XNOR U1304 ( .A(in[833]), .B(in[193]), .Z(n692) );
  XNOR U1305 ( .A(n693), .B(n692), .Z(n694) );
  XNOR U1306 ( .A(in[1153]), .B(n694), .Z(n1362) );
  XOR U1307 ( .A(n1673), .B(n1362), .Z(n1999) );
  XOR U1308 ( .A(in[129]), .B(n1999), .Z(n1586) );
  XOR U1309 ( .A(in[353]), .B(in[673]), .Z(n696) );
  XNOR U1310 ( .A(in[33]), .B(in[1313]), .Z(n695) );
  XNOR U1311 ( .A(n696), .B(n695), .Z(n697) );
  XNOR U1312 ( .A(in[993]), .B(n697), .Z(n1481) );
  XNOR U1313 ( .A(in[1378]), .B(n4542), .Z(n1994) );
  XOR U1314 ( .A(in[1577]), .B(in[617]), .Z(n700) );
  XNOR U1315 ( .A(in[937]), .B(in[297]), .Z(n699) );
  XNOR U1316 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1317 ( .A(in[1257]), .B(n701), .Z(n1052) );
  XOR U1318 ( .A(n702), .B(n1052), .Z(n4298) );
  XOR U1319 ( .A(in[1002]), .B(n4298), .Z(n1991) );
  NANDN U1320 ( .A(n1994), .B(n1991), .Z(n703) );
  XNOR U1321 ( .A(n1586), .B(n703), .Z(out[1022]) );
  IV U1322 ( .A(n3175), .Z(n3934) );
  XOR U1323 ( .A(n3934), .B(in[130]), .Z(n1588) );
  XOR U1324 ( .A(in[354]), .B(in[674]), .Z(n705) );
  XNOR U1325 ( .A(in[34]), .B(in[1314]), .Z(n704) );
  XNOR U1326 ( .A(n705), .B(n704), .Z(n706) );
  XNOR U1327 ( .A(in[994]), .B(n706), .Z(n1484) );
  XOR U1328 ( .A(in[163]), .B(in[1443]), .Z(n708) );
  XNOR U1329 ( .A(in[803]), .B(in[1123]), .Z(n707) );
  XNOR U1330 ( .A(n708), .B(n707), .Z(n709) );
  XOR U1331 ( .A(in[483]), .B(n709), .Z(n809) );
  XNOR U1332 ( .A(in[1379]), .B(n4546), .Z(n1998) );
  XOR U1333 ( .A(in[1578]), .B(in[618]), .Z(n711) );
  XNOR U1334 ( .A(in[938]), .B(in[298]), .Z(n710) );
  XNOR U1335 ( .A(n711), .B(n710), .Z(n712) );
  XNOR U1336 ( .A(in[1258]), .B(n712), .Z(n1065) );
  XOR U1337 ( .A(n713), .B(n1065), .Z(n4300) );
  XOR U1338 ( .A(in[1003]), .B(n4300), .Z(n1995) );
  NANDN U1339 ( .A(n1998), .B(n1995), .Z(n714) );
  XOR U1340 ( .A(n1588), .B(n714), .Z(out[1023]) );
  XNOR U1341 ( .A(n716), .B(n715), .Z(n3987) );
  XOR U1342 ( .A(in[531]), .B(n3987), .Z(n1592) );
  XOR U1343 ( .A(in[35]), .B(in[675]), .Z(n718) );
  XNOR U1344 ( .A(in[355]), .B(in[1315]), .Z(n717) );
  XNOR U1345 ( .A(n718), .B(n717), .Z(n719) );
  XNOR U1346 ( .A(in[995]), .B(n719), .Z(n1487) );
  XOR U1347 ( .A(in[164]), .B(in[1444]), .Z(n721) );
  XNOR U1348 ( .A(in[804]), .B(in[1124]), .Z(n720) );
  XNOR U1349 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U1350 ( .A(in[484]), .B(n722), .Z(n968) );
  XOR U1351 ( .A(n1487), .B(n968), .Z(n4550) );
  XNOR U1352 ( .A(in[1380]), .B(n4550), .Z(n5002) );
  XOR U1353 ( .A(in[1346]), .B(in[66]), .Z(n724) );
  XNOR U1354 ( .A(in[1026]), .B(in[386]), .Z(n723) );
  XNOR U1355 ( .A(n724), .B(n723), .Z(n725) );
  XNOR U1356 ( .A(in[706]), .B(n725), .Z(n1681) );
  XOR U1357 ( .A(in[1475]), .B(in[515]), .Z(n727) );
  XNOR U1358 ( .A(in[835]), .B(in[195]), .Z(n726) );
  XNOR U1359 ( .A(n727), .B(n726), .Z(n728) );
  XOR U1360 ( .A(in[1155]), .B(n728), .Z(n1405) );
  XOR U1361 ( .A(in[131]), .B(n3177), .Z(n5004) );
  OR U1362 ( .A(n5002), .B(n5004), .Z(n729) );
  XNOR U1363 ( .A(n1592), .B(n729), .Z(out[1024]) );
  XNOR U1364 ( .A(n731), .B(n730), .Z(n3991) );
  XOR U1365 ( .A(in[532]), .B(n3991), .Z(n1596) );
  XOR U1366 ( .A(in[1445]), .B(in[165]), .Z(n733) );
  XNOR U1367 ( .A(in[805]), .B(in[1125]), .Z(n732) );
  XNOR U1368 ( .A(n733), .B(n732), .Z(n734) );
  XNOR U1369 ( .A(in[485]), .B(n734), .Z(n1012) );
  XOR U1370 ( .A(in[36]), .B(in[676]), .Z(n736) );
  XNOR U1371 ( .A(in[356]), .B(in[1316]), .Z(n735) );
  XNOR U1372 ( .A(n736), .B(n735), .Z(n737) );
  XNOR U1373 ( .A(in[996]), .B(n737), .Z(n1490) );
  XOR U1374 ( .A(n1012), .B(n1490), .Z(n4556) );
  XNOR U1375 ( .A(in[1381]), .B(n4556), .Z(n5006) );
  XOR U1376 ( .A(in[1347]), .B(in[67]), .Z(n739) );
  XNOR U1377 ( .A(in[1027]), .B(in[387]), .Z(n738) );
  XNOR U1378 ( .A(n739), .B(n738), .Z(n740) );
  XNOR U1379 ( .A(in[707]), .B(n740), .Z(n1685) );
  XOR U1380 ( .A(in[1476]), .B(in[516]), .Z(n742) );
  XNOR U1381 ( .A(in[836]), .B(in[196]), .Z(n741) );
  XNOR U1382 ( .A(n742), .B(n741), .Z(n743) );
  XOR U1383 ( .A(in[1156]), .B(n743), .Z(n1407) );
  XOR U1384 ( .A(in[132]), .B(n3179), .Z(n5008) );
  OR U1385 ( .A(n5006), .B(n5008), .Z(n744) );
  XNOR U1386 ( .A(n1596), .B(n744), .Z(out[1025]) );
  XNOR U1387 ( .A(n746), .B(n745), .Z(n3995) );
  XOR U1388 ( .A(in[533]), .B(n3995), .Z(n1600) );
  XOR U1389 ( .A(in[166]), .B(in[806]), .Z(n748) );
  XNOR U1390 ( .A(in[1126]), .B(in[486]), .Z(n747) );
  XNOR U1391 ( .A(n748), .B(n747), .Z(n749) );
  XNOR U1392 ( .A(in[1446]), .B(n749), .Z(n1025) );
  XOR U1393 ( .A(in[37]), .B(in[677]), .Z(n751) );
  XNOR U1394 ( .A(in[357]), .B(in[1317]), .Z(n750) );
  XNOR U1395 ( .A(n751), .B(n750), .Z(n752) );
  XNOR U1396 ( .A(in[997]), .B(n752), .Z(n1493) );
  XOR U1397 ( .A(n1025), .B(n1493), .Z(n4558) );
  XNOR U1398 ( .A(in[1382]), .B(n4558), .Z(n5010) );
  XOR U1399 ( .A(in[1348]), .B(in[68]), .Z(n754) );
  XNOR U1400 ( .A(in[1028]), .B(in[388]), .Z(n753) );
  XNOR U1401 ( .A(n754), .B(n753), .Z(n755) );
  XNOR U1402 ( .A(in[708]), .B(n755), .Z(n1689) );
  XOR U1403 ( .A(in[1477]), .B(in[517]), .Z(n757) );
  XNOR U1404 ( .A(in[837]), .B(in[197]), .Z(n756) );
  XNOR U1405 ( .A(n757), .B(n756), .Z(n758) );
  XOR U1406 ( .A(in[1157]), .B(n758), .Z(n1409) );
  XOR U1407 ( .A(in[133]), .B(n3181), .Z(n5012) );
  OR U1408 ( .A(n5010), .B(n5012), .Z(n759) );
  XNOR U1409 ( .A(n1600), .B(n759), .Z(out[1026]) );
  XOR U1410 ( .A(n761), .B(n760), .Z(n2003) );
  XOR U1411 ( .A(in[534]), .B(n2003), .Z(n1604) );
  XOR U1412 ( .A(in[38]), .B(in[678]), .Z(n763) );
  XNOR U1413 ( .A(in[358]), .B(in[1318]), .Z(n762) );
  XNOR U1414 ( .A(n763), .B(n762), .Z(n764) );
  XNOR U1415 ( .A(in[998]), .B(n764), .Z(n1497) );
  XOR U1416 ( .A(in[167]), .B(in[807]), .Z(n766) );
  XNOR U1417 ( .A(in[1127]), .B(in[487]), .Z(n765) );
  XNOR U1418 ( .A(n766), .B(n765), .Z(n767) );
  XNOR U1419 ( .A(in[1447]), .B(n767), .Z(n1038) );
  XOR U1420 ( .A(n1497), .B(n1038), .Z(n4339) );
  XNOR U1421 ( .A(in[1383]), .B(n4339), .Z(n5014) );
  XOR U1422 ( .A(in[1349]), .B(in[69]), .Z(n769) );
  XNOR U1423 ( .A(in[1029]), .B(in[389]), .Z(n768) );
  XNOR U1424 ( .A(n769), .B(n768), .Z(n770) );
  XNOR U1425 ( .A(in[709]), .B(n770), .Z(n1693) );
  XOR U1426 ( .A(in[1478]), .B(in[518]), .Z(n772) );
  XNOR U1427 ( .A(in[838]), .B(in[198]), .Z(n771) );
  XNOR U1428 ( .A(n772), .B(n771), .Z(n773) );
  XOR U1429 ( .A(in[1158]), .B(n773), .Z(n1411) );
  XOR U1430 ( .A(in[134]), .B(n3183), .Z(n5016) );
  OR U1431 ( .A(n5014), .B(n5016), .Z(n774) );
  XNOR U1432 ( .A(n1604), .B(n774), .Z(out[1027]) );
  XNOR U1433 ( .A(n776), .B(n775), .Z(n4003) );
  XOR U1434 ( .A(in[535]), .B(n4003), .Z(n1608) );
  XOR U1435 ( .A(in[39]), .B(in[679]), .Z(n778) );
  XNOR U1436 ( .A(in[359]), .B(in[1319]), .Z(n777) );
  XNOR U1437 ( .A(n778), .B(n777), .Z(n779) );
  XNOR U1438 ( .A(in[999]), .B(n779), .Z(n1502) );
  XOR U1439 ( .A(in[168]), .B(in[1448]), .Z(n781) );
  XNOR U1440 ( .A(in[1128]), .B(in[808]), .Z(n780) );
  XNOR U1441 ( .A(n781), .B(n780), .Z(n782) );
  XNOR U1442 ( .A(in[488]), .B(n782), .Z(n1051) );
  XOR U1443 ( .A(n1502), .B(n1051), .Z(n4341) );
  XNOR U1444 ( .A(in[1384]), .B(n4341), .Z(n5018) );
  XOR U1445 ( .A(in[1350]), .B(in[70]), .Z(n784) );
  XNOR U1446 ( .A(in[1030]), .B(in[390]), .Z(n783) );
  XNOR U1447 ( .A(n784), .B(n783), .Z(n785) );
  XNOR U1448 ( .A(in[710]), .B(n785), .Z(n1697) );
  XOR U1449 ( .A(in[199]), .B(in[1479]), .Z(n787) );
  XNOR U1450 ( .A(in[1159]), .B(in[839]), .Z(n786) );
  XNOR U1451 ( .A(n787), .B(n786), .Z(n788) );
  XOR U1452 ( .A(in[519]), .B(n788), .Z(n1413) );
  XOR U1453 ( .A(in[135]), .B(n3185), .Z(n5020) );
  OR U1454 ( .A(n5018), .B(n5020), .Z(n789) );
  XNOR U1455 ( .A(n1608), .B(n789), .Z(out[1028]) );
  XOR U1456 ( .A(n791), .B(n790), .Z(n2006) );
  XOR U1457 ( .A(in[536]), .B(n2006), .Z(n1612) );
  XOR U1458 ( .A(in[680]), .B(in[1320]), .Z(n793) );
  XNOR U1459 ( .A(in[40]), .B(in[360]), .Z(n792) );
  XNOR U1460 ( .A(n793), .B(n792), .Z(n794) );
  XNOR U1461 ( .A(in[1000]), .B(n794), .Z(n1506) );
  XOR U1462 ( .A(in[169]), .B(in[1449]), .Z(n796) );
  XNOR U1463 ( .A(in[1129]), .B(in[809]), .Z(n795) );
  XNOR U1464 ( .A(n796), .B(n795), .Z(n797) );
  XNOR U1465 ( .A(in[489]), .B(n797), .Z(n1064) );
  XOR U1466 ( .A(n1506), .B(n1064), .Z(n4347) );
  XNOR U1467 ( .A(in[1385]), .B(n4347), .Z(n5022) );
  XOR U1468 ( .A(in[1351]), .B(in[711]), .Z(n799) );
  XNOR U1469 ( .A(in[1031]), .B(in[391]), .Z(n798) );
  XNOR U1470 ( .A(n799), .B(n798), .Z(n800) );
  XNOR U1471 ( .A(in[71]), .B(n800), .Z(n1701) );
  XOR U1472 ( .A(in[1480]), .B(in[520]), .Z(n802) );
  XNOR U1473 ( .A(in[840]), .B(in[200]), .Z(n801) );
  XNOR U1474 ( .A(n802), .B(n801), .Z(n803) );
  XOR U1475 ( .A(in[1160]), .B(n803), .Z(n1418) );
  XOR U1476 ( .A(in[136]), .B(n3187), .Z(n5024) );
  OR U1477 ( .A(n5022), .B(n5024), .Z(n804) );
  XNOR U1478 ( .A(n1612), .B(n804), .Z(out[1029]) );
  XOR U1479 ( .A(in[1341]), .B(in[61]), .Z(n806) );
  XNOR U1480 ( .A(in[701]), .B(in[381]), .Z(n805) );
  XNOR U1481 ( .A(n806), .B(n805), .Z(n807) );
  XNOR U1482 ( .A(in[1021]), .B(n807), .Z(n1121) );
  XOR U1483 ( .A(n808), .B(n1121), .Z(n3963) );
  XOR U1484 ( .A(in[637]), .B(n3963), .Z(n2710) );
  IV U1485 ( .A(n2710), .Z(n2799) );
  XOR U1486 ( .A(n810), .B(n809), .Z(n3404) );
  IV U1487 ( .A(n3404), .Z(n4059) );
  XOR U1488 ( .A(in[228]), .B(n4059), .Z(n3160) );
  XOR U1489 ( .A(in[1512]), .B(in[552]), .Z(n812) );
  XNOR U1490 ( .A(in[872]), .B(in[232]), .Z(n811) );
  XNOR U1491 ( .A(n812), .B(n811), .Z(n813) );
  XNOR U1492 ( .A(in[1192]), .B(n813), .Z(n1511) );
  XNOR U1493 ( .A(n814), .B(n1511), .Z(n4099) );
  IV U1494 ( .A(n4099), .Z(n1270) );
  XOR U1495 ( .A(in[1448]), .B(n1270), .Z(n3158) );
  NANDN U1496 ( .A(n3160), .B(n3158), .Z(n815) );
  XOR U1497 ( .A(n2799), .B(n815), .Z(out[102]) );
  XOR U1498 ( .A(n817), .B(n816), .Z(n2009) );
  XOR U1499 ( .A(in[537]), .B(n2009), .Z(n1616) );
  XOR U1500 ( .A(in[1352]), .B(in[712]), .Z(n819) );
  XNOR U1501 ( .A(in[1032]), .B(in[392]), .Z(n818) );
  XNOR U1502 ( .A(n819), .B(n818), .Z(n820) );
  XNOR U1503 ( .A(in[72]), .B(n820), .Z(n1707) );
  XOR U1504 ( .A(in[1481]), .B(in[521]), .Z(n822) );
  XNOR U1505 ( .A(in[841]), .B(in[201]), .Z(n821) );
  XNOR U1506 ( .A(n822), .B(n821), .Z(n823) );
  XOR U1507 ( .A(in[1161]), .B(n823), .Z(n1420) );
  XOR U1508 ( .A(in[137]), .B(n3189), .Z(n5028) );
  XOR U1509 ( .A(in[170]), .B(in[1450]), .Z(n825) );
  XNOR U1510 ( .A(in[1130]), .B(in[810]), .Z(n824) );
  XNOR U1511 ( .A(n825), .B(n824), .Z(n826) );
  XNOR U1512 ( .A(in[490]), .B(n826), .Z(n1080) );
  XOR U1513 ( .A(in[681]), .B(in[1321]), .Z(n828) );
  XNOR U1514 ( .A(in[41]), .B(in[361]), .Z(n827) );
  XNOR U1515 ( .A(n828), .B(n827), .Z(n829) );
  XNOR U1516 ( .A(in[1001]), .B(n829), .Z(n1510) );
  XOR U1517 ( .A(n1080), .B(n1510), .Z(n4349) );
  XOR U1518 ( .A(in[1386]), .B(n4349), .Z(n5025) );
  NANDN U1519 ( .A(n5028), .B(n5025), .Z(n830) );
  XNOR U1520 ( .A(n1616), .B(n830), .Z(out[1030]) );
  XOR U1521 ( .A(n832), .B(n831), .Z(n2012) );
  XOR U1522 ( .A(in[538]), .B(n2012), .Z(n1620) );
  XOR U1523 ( .A(in[1353]), .B(in[393]), .Z(n834) );
  XNOR U1524 ( .A(in[713]), .B(in[73]), .Z(n833) );
  XNOR U1525 ( .A(n834), .B(n833), .Z(n835) );
  XNOR U1526 ( .A(in[1033]), .B(n835), .Z(n1711) );
  XOR U1527 ( .A(in[1482]), .B(in[522]), .Z(n837) );
  XNOR U1528 ( .A(in[842]), .B(in[202]), .Z(n836) );
  XNOR U1529 ( .A(n837), .B(n836), .Z(n838) );
  XOR U1530 ( .A(n1711), .B(n227), .Z(n3191) );
  XOR U1531 ( .A(in[138]), .B(n3191), .Z(n5032) );
  XOR U1532 ( .A(in[811]), .B(in[491]), .Z(n840) );
  XNOR U1533 ( .A(in[1451]), .B(in[1131]), .Z(n839) );
  XNOR U1534 ( .A(n840), .B(n839), .Z(n841) );
  XNOR U1535 ( .A(in[171]), .B(n841), .Z(n1093) );
  XOR U1536 ( .A(in[682]), .B(in[1322]), .Z(n843) );
  XNOR U1537 ( .A(in[42]), .B(in[362]), .Z(n842) );
  XNOR U1538 ( .A(n843), .B(n842), .Z(n844) );
  XNOR U1539 ( .A(in[1002]), .B(n844), .Z(n1515) );
  XOR U1540 ( .A(n1093), .B(n1515), .Z(n4351) );
  XOR U1541 ( .A(in[1387]), .B(n4351), .Z(n5029) );
  NANDN U1542 ( .A(n5032), .B(n5029), .Z(n845) );
  XNOR U1543 ( .A(n1620), .B(n845), .Z(out[1031]) );
  XOR U1544 ( .A(n847), .B(n846), .Z(n2015) );
  XOR U1545 ( .A(in[539]), .B(n2015), .Z(n1625) );
  XOR U1546 ( .A(in[1483]), .B(in[523]), .Z(n849) );
  XNOR U1547 ( .A(in[843]), .B(in[203]), .Z(n848) );
  XNOR U1548 ( .A(n849), .B(n848), .Z(n850) );
  XNOR U1549 ( .A(in[1163]), .B(n850), .Z(n1423) );
  XOR U1550 ( .A(in[1354]), .B(in[714]), .Z(n852) );
  XNOR U1551 ( .A(in[74]), .B(in[394]), .Z(n851) );
  XNOR U1552 ( .A(n852), .B(n851), .Z(n853) );
  XOR U1553 ( .A(in[1034]), .B(n853), .Z(n1715) );
  XOR U1554 ( .A(n2296), .B(in[139]), .Z(n5036) );
  XOR U1555 ( .A(in[683]), .B(in[1323]), .Z(n855) );
  XNOR U1556 ( .A(in[43]), .B(in[363]), .Z(n854) );
  XNOR U1557 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U1558 ( .A(in[1003]), .B(n856), .Z(n1519) );
  XOR U1559 ( .A(in[812]), .B(in[492]), .Z(n858) );
  XNOR U1560 ( .A(in[1452]), .B(in[1132]), .Z(n857) );
  XNOR U1561 ( .A(n858), .B(n857), .Z(n859) );
  XNOR U1562 ( .A(in[172]), .B(n859), .Z(n1113) );
  XOR U1563 ( .A(n1519), .B(n1113), .Z(n4354) );
  XOR U1564 ( .A(in[1388]), .B(n4354), .Z(n5033) );
  NANDN U1565 ( .A(n5036), .B(n5033), .Z(n860) );
  XNOR U1566 ( .A(n1625), .B(n860), .Z(out[1032]) );
  XOR U1567 ( .A(n862), .B(n861), .Z(n4023) );
  XOR U1568 ( .A(in[540]), .B(n4023), .Z(n1629) );
  XOR U1569 ( .A(in[1355]), .B(in[715]), .Z(n864) );
  XNOR U1570 ( .A(in[1035]), .B(in[395]), .Z(n863) );
  XNOR U1571 ( .A(n864), .B(n863), .Z(n865) );
  XNOR U1572 ( .A(in[75]), .B(n865), .Z(n1719) );
  XOR U1573 ( .A(in[1484]), .B(in[524]), .Z(n867) );
  XNOR U1574 ( .A(in[844]), .B(in[204]), .Z(n866) );
  XNOR U1575 ( .A(n867), .B(n866), .Z(n868) );
  XOR U1576 ( .A(in[1164]), .B(n868), .Z(n1425) );
  XOR U1577 ( .A(in[140]), .B(n3198), .Z(n5040) );
  XOR U1578 ( .A(in[1324]), .B(in[44]), .Z(n870) );
  XNOR U1579 ( .A(in[684]), .B(in[364]), .Z(n869) );
  XNOR U1580 ( .A(n870), .B(n869), .Z(n871) );
  XNOR U1581 ( .A(in[1004]), .B(n871), .Z(n1522) );
  XOR U1582 ( .A(in[813]), .B(in[493]), .Z(n873) );
  XNOR U1583 ( .A(in[1453]), .B(in[1133]), .Z(n872) );
  XNOR U1584 ( .A(n873), .B(n872), .Z(n874) );
  XNOR U1585 ( .A(in[173]), .B(n874), .Z(n1126) );
  XOR U1586 ( .A(n1522), .B(n1126), .Z(n4357) );
  XOR U1587 ( .A(in[1389]), .B(n4357), .Z(n5037) );
  NANDN U1588 ( .A(n5040), .B(n5037), .Z(n875) );
  XNOR U1589 ( .A(n1629), .B(n875), .Z(out[1033]) );
  XOR U1590 ( .A(n877), .B(n876), .Z(n4031) );
  XOR U1591 ( .A(in[541]), .B(n4031), .Z(n1633) );
  XOR U1592 ( .A(in[76]), .B(in[1036]), .Z(n879) );
  XNOR U1593 ( .A(in[716]), .B(in[396]), .Z(n878) );
  XNOR U1594 ( .A(n879), .B(n878), .Z(n880) );
  XNOR U1595 ( .A(in[1356]), .B(n880), .Z(n1723) );
  XOR U1596 ( .A(in[1485]), .B(in[525]), .Z(n882) );
  XNOR U1597 ( .A(in[845]), .B(in[205]), .Z(n881) );
  XNOR U1598 ( .A(n882), .B(n881), .Z(n883) );
  XOR U1599 ( .A(in[1165]), .B(n883), .Z(n1427) );
  XOR U1600 ( .A(in[141]), .B(n3200), .Z(n5048) );
  XOR U1601 ( .A(in[814]), .B(in[494]), .Z(n885) );
  XNOR U1602 ( .A(in[1454]), .B(in[1134]), .Z(n884) );
  XNOR U1603 ( .A(n885), .B(n884), .Z(n886) );
  XNOR U1604 ( .A(in[174]), .B(n886), .Z(n1139) );
  XOR U1605 ( .A(in[1325]), .B(in[45]), .Z(n888) );
  XNOR U1606 ( .A(in[685]), .B(in[365]), .Z(n887) );
  XNOR U1607 ( .A(n888), .B(n887), .Z(n889) );
  XNOR U1608 ( .A(in[1005]), .B(n889), .Z(n1526) );
  XOR U1609 ( .A(n1139), .B(n1526), .Z(n4360) );
  XOR U1610 ( .A(in[1390]), .B(n4360), .Z(n5045) );
  NANDN U1611 ( .A(n5048), .B(n5045), .Z(n890) );
  XNOR U1612 ( .A(n1633), .B(n890), .Z(out[1034]) );
  XOR U1613 ( .A(n892), .B(n891), .Z(n4035) );
  XOR U1614 ( .A(in[542]), .B(n4035), .Z(n1637) );
  XOR U1615 ( .A(in[77]), .B(in[1037]), .Z(n894) );
  XNOR U1616 ( .A(in[717]), .B(in[397]), .Z(n893) );
  XNOR U1617 ( .A(n894), .B(n893), .Z(n895) );
  XNOR U1618 ( .A(in[1357]), .B(n895), .Z(n1727) );
  XOR U1619 ( .A(in[1486]), .B(in[526]), .Z(n897) );
  XNOR U1620 ( .A(in[846]), .B(in[206]), .Z(n896) );
  XNOR U1621 ( .A(n897), .B(n896), .Z(n898) );
  XOR U1622 ( .A(in[1166]), .B(n898), .Z(n1429) );
  XOR U1623 ( .A(in[142]), .B(n3203), .Z(n5052) );
  XOR U1624 ( .A(in[815]), .B(in[495]), .Z(n900) );
  XNOR U1625 ( .A(in[1455]), .B(in[1135]), .Z(n899) );
  XNOR U1626 ( .A(n900), .B(n899), .Z(n901) );
  XNOR U1627 ( .A(in[175]), .B(n901), .Z(n1152) );
  XOR U1628 ( .A(in[1326]), .B(in[46]), .Z(n903) );
  XNOR U1629 ( .A(in[686]), .B(in[366]), .Z(n902) );
  XNOR U1630 ( .A(n903), .B(n902), .Z(n904) );
  XNOR U1631 ( .A(in[1006]), .B(n904), .Z(n1530) );
  XOR U1632 ( .A(n1152), .B(n1530), .Z(n4362) );
  XOR U1633 ( .A(in[1391]), .B(n4362), .Z(n5049) );
  NANDN U1634 ( .A(n5052), .B(n5049), .Z(n905) );
  XNOR U1635 ( .A(n1637), .B(n905), .Z(out[1035]) );
  XOR U1636 ( .A(n907), .B(n906), .Z(n4039) );
  XOR U1637 ( .A(in[543]), .B(n4039), .Z(n1641) );
  XOR U1638 ( .A(in[78]), .B(in[1038]), .Z(n909) );
  XNOR U1639 ( .A(in[718]), .B(in[398]), .Z(n908) );
  XNOR U1640 ( .A(n909), .B(n908), .Z(n910) );
  XNOR U1641 ( .A(in[1358]), .B(n910), .Z(n1731) );
  XOR U1642 ( .A(in[1487]), .B(in[527]), .Z(n912) );
  XNOR U1643 ( .A(in[847]), .B(in[207]), .Z(n911) );
  XNOR U1644 ( .A(n912), .B(n911), .Z(n913) );
  XOR U1645 ( .A(in[1167]), .B(n913), .Z(n1431) );
  XOR U1646 ( .A(in[143]), .B(n3206), .Z(n5056) );
  XOR U1647 ( .A(in[816]), .B(in[496]), .Z(n915) );
  XNOR U1648 ( .A(in[1456]), .B(in[1136]), .Z(n914) );
  XNOR U1649 ( .A(n915), .B(n914), .Z(n916) );
  XNOR U1650 ( .A(in[176]), .B(n916), .Z(n1167) );
  XOR U1651 ( .A(in[1327]), .B(in[47]), .Z(n918) );
  XNOR U1652 ( .A(in[687]), .B(in[367]), .Z(n917) );
  XNOR U1653 ( .A(n918), .B(n917), .Z(n919) );
  XNOR U1654 ( .A(in[1007]), .B(n919), .Z(n1534) );
  XOR U1655 ( .A(n1167), .B(n1534), .Z(n4365) );
  XOR U1656 ( .A(in[1392]), .B(n4365), .Z(n5053) );
  NANDN U1657 ( .A(n5056), .B(n5053), .Z(n920) );
  XNOR U1658 ( .A(n1641), .B(n920), .Z(out[1036]) );
  XOR U1659 ( .A(n922), .B(n921), .Z(n4043) );
  XOR U1660 ( .A(in[544]), .B(n4043), .Z(n1645) );
  XOR U1661 ( .A(in[79]), .B(in[1039]), .Z(n924) );
  XNOR U1662 ( .A(in[719]), .B(in[399]), .Z(n923) );
  XNOR U1663 ( .A(n924), .B(n923), .Z(n925) );
  XNOR U1664 ( .A(in[1359]), .B(n925), .Z(n1735) );
  XOR U1665 ( .A(in[1488]), .B(in[528]), .Z(n927) );
  XNOR U1666 ( .A(in[848]), .B(in[208]), .Z(n926) );
  XNOR U1667 ( .A(n927), .B(n926), .Z(n928) );
  XOR U1668 ( .A(in[1168]), .B(n928), .Z(n1433) );
  XOR U1669 ( .A(in[144]), .B(n3209), .Z(n5060) );
  XOR U1670 ( .A(in[1328]), .B(in[48]), .Z(n930) );
  XNOR U1671 ( .A(in[688]), .B(in[368]), .Z(n929) );
  XNOR U1672 ( .A(n930), .B(n929), .Z(n931) );
  XNOR U1673 ( .A(in[1008]), .B(n931), .Z(n1538) );
  XOR U1674 ( .A(in[817]), .B(in[497]), .Z(n933) );
  XNOR U1675 ( .A(in[1457]), .B(in[1137]), .Z(n932) );
  XNOR U1676 ( .A(n933), .B(n932), .Z(n934) );
  XNOR U1677 ( .A(in[177]), .B(n934), .Z(n1182) );
  XOR U1678 ( .A(n1538), .B(n1182), .Z(n4368) );
  XOR U1679 ( .A(in[1393]), .B(n4368), .Z(n5057) );
  NANDN U1680 ( .A(n5060), .B(n5057), .Z(n935) );
  XNOR U1681 ( .A(n1645), .B(n935), .Z(out[1037]) );
  XOR U1682 ( .A(n937), .B(n936), .Z(n4047) );
  XOR U1683 ( .A(in[545]), .B(n4047), .Z(n1649) );
  XOR U1684 ( .A(in[80]), .B(in[1040]), .Z(n939) );
  XNOR U1685 ( .A(in[720]), .B(in[400]), .Z(n938) );
  XNOR U1686 ( .A(n939), .B(n938), .Z(n940) );
  XNOR U1687 ( .A(in[1360]), .B(n940), .Z(n1739) );
  XOR U1688 ( .A(in[1489]), .B(in[529]), .Z(n942) );
  XNOR U1689 ( .A(in[849]), .B(in[209]), .Z(n941) );
  XNOR U1690 ( .A(n942), .B(n941), .Z(n943) );
  XOR U1691 ( .A(in[1169]), .B(n943), .Z(n1435) );
  XOR U1692 ( .A(in[145]), .B(n3212), .Z(n5064) );
  XOR U1693 ( .A(in[1329]), .B(in[49]), .Z(n945) );
  XNOR U1694 ( .A(in[689]), .B(in[369]), .Z(n944) );
  XNOR U1695 ( .A(n945), .B(n944), .Z(n946) );
  XNOR U1696 ( .A(in[1009]), .B(n946), .Z(n1544) );
  XOR U1697 ( .A(in[818]), .B(in[498]), .Z(n948) );
  XNOR U1698 ( .A(in[1458]), .B(in[1138]), .Z(n947) );
  XNOR U1699 ( .A(n948), .B(n947), .Z(n949) );
  XNOR U1700 ( .A(in[178]), .B(n949), .Z(n1197) );
  XOR U1701 ( .A(n1544), .B(n1197), .Z(n4371) );
  XOR U1702 ( .A(in[1394]), .B(n4371), .Z(n5061) );
  NANDN U1703 ( .A(n5064), .B(n5061), .Z(n950) );
  XNOR U1704 ( .A(n1649), .B(n950), .Z(out[1038]) );
  IV U1705 ( .A(n4051), .Z(n3397) );
  XOR U1706 ( .A(n3397), .B(in[546]), .Z(n1653) );
  XOR U1707 ( .A(in[81]), .B(in[1041]), .Z(n952) );
  XNOR U1708 ( .A(in[721]), .B(in[401]), .Z(n951) );
  XNOR U1709 ( .A(n952), .B(n951), .Z(n953) );
  XNOR U1710 ( .A(in[1361]), .B(n953), .Z(n1743) );
  XOR U1711 ( .A(in[1490]), .B(in[530]), .Z(n955) );
  XNOR U1712 ( .A(in[850]), .B(in[210]), .Z(n954) );
  XNOR U1713 ( .A(n955), .B(n954), .Z(n956) );
  XOR U1714 ( .A(in[1170]), .B(n956), .Z(n1439) );
  XOR U1715 ( .A(in[146]), .B(n4004), .Z(n5068) );
  XOR U1716 ( .A(in[819]), .B(in[499]), .Z(n958) );
  XNOR U1717 ( .A(in[1459]), .B(in[1139]), .Z(n957) );
  XNOR U1718 ( .A(n958), .B(n957), .Z(n959) );
  XNOR U1719 ( .A(in[179]), .B(n959), .Z(n1212) );
  XOR U1720 ( .A(in[1330]), .B(in[50]), .Z(n961) );
  XNOR U1721 ( .A(in[690]), .B(in[370]), .Z(n960) );
  XNOR U1722 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U1723 ( .A(in[1010]), .B(n962), .Z(n1548) );
  XOR U1724 ( .A(n1212), .B(n1548), .Z(n4378) );
  XOR U1725 ( .A(in[1395]), .B(n4378), .Z(n5065) );
  NANDN U1726 ( .A(n5068), .B(n5065), .Z(n963) );
  XOR U1727 ( .A(n1653), .B(n963), .Z(out[1039]) );
  XOR U1728 ( .A(in[1342]), .B(in[62]), .Z(n965) );
  XNOR U1729 ( .A(in[702]), .B(in[382]), .Z(n964) );
  XNOR U1730 ( .A(n965), .B(n964), .Z(n966) );
  XNOR U1731 ( .A(in[1022]), .B(n966), .Z(n1134) );
  XOR U1732 ( .A(n967), .B(n1134), .Z(n3967) );
  XOR U1733 ( .A(in[638]), .B(n3967), .Z(n2712) );
  IV U1734 ( .A(n2712), .Z(n2801) );
  XOR U1735 ( .A(n969), .B(n968), .Z(n4063) );
  XOR U1736 ( .A(in[229]), .B(n4063), .Z(n3171) );
  XOR U1737 ( .A(in[1513]), .B(in[553]), .Z(n971) );
  XNOR U1738 ( .A(in[873]), .B(in[233]), .Z(n970) );
  XNOR U1739 ( .A(n971), .B(n970), .Z(n972) );
  XNOR U1740 ( .A(in[1193]), .B(n972), .Z(n1514) );
  XNOR U1741 ( .A(n973), .B(n1514), .Z(n4103) );
  IV U1742 ( .A(n4103), .Z(n1282) );
  XOR U1743 ( .A(in[1449]), .B(n1282), .Z(n3168) );
  NANDN U1744 ( .A(n3171), .B(n3168), .Z(n974) );
  XOR U1745 ( .A(n2801), .B(n974), .Z(out[103]) );
  XOR U1746 ( .A(n3400), .B(in[547]), .Z(n1657) );
  XOR U1747 ( .A(in[1042]), .B(in[402]), .Z(n976) );
  XNOR U1748 ( .A(in[722]), .B(in[82]), .Z(n975) );
  XNOR U1749 ( .A(n976), .B(n975), .Z(n977) );
  XNOR U1750 ( .A(in[1362]), .B(n977), .Z(n1748) );
  XOR U1751 ( .A(in[851]), .B(in[1171]), .Z(n979) );
  XNOR U1752 ( .A(in[1491]), .B(in[211]), .Z(n978) );
  XNOR U1753 ( .A(n979), .B(n978), .Z(n980) );
  XOR U1754 ( .A(in[531]), .B(n980), .Z(n1441) );
  IV U1755 ( .A(n3217), .Z(n4008) );
  XNOR U1756 ( .A(in[147]), .B(n4008), .Z(n5071) );
  XOR U1757 ( .A(in[820]), .B(in[500]), .Z(n982) );
  XNOR U1758 ( .A(in[1460]), .B(in[1140]), .Z(n981) );
  XNOR U1759 ( .A(n982), .B(n981), .Z(n983) );
  XNOR U1760 ( .A(in[180]), .B(n983), .Z(n1227) );
  XOR U1761 ( .A(in[1331]), .B(in[51]), .Z(n985) );
  XNOR U1762 ( .A(in[691]), .B(in[371]), .Z(n984) );
  XNOR U1763 ( .A(n985), .B(n984), .Z(n986) );
  XNOR U1764 ( .A(in[1011]), .B(n986), .Z(n1552) );
  XOR U1765 ( .A(n1227), .B(n1552), .Z(n4381) );
  XOR U1766 ( .A(in[1396]), .B(n4381), .Z(n5070) );
  NANDN U1767 ( .A(n5071), .B(n5070), .Z(n987) );
  XOR U1768 ( .A(n1657), .B(n987), .Z(out[1040]) );
  XOR U1769 ( .A(n3404), .B(in[548]), .Z(n1661) );
  XOR U1770 ( .A(in[83]), .B(in[1043]), .Z(n989) );
  XNOR U1771 ( .A(in[723]), .B(in[403]), .Z(n988) );
  XNOR U1772 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U1773 ( .A(in[1363]), .B(n990), .Z(n1752) );
  XOR U1774 ( .A(in[852]), .B(in[1172]), .Z(n992) );
  XNOR U1775 ( .A(in[1492]), .B(in[212]), .Z(n991) );
  XNOR U1776 ( .A(n992), .B(n991), .Z(n993) );
  XOR U1777 ( .A(in[532]), .B(n993), .Z(n1443) );
  IV U1778 ( .A(n3220), .Z(n4012) );
  XNOR U1779 ( .A(in[148]), .B(n4012), .Z(n5074) );
  XOR U1780 ( .A(in[1332]), .B(in[52]), .Z(n995) );
  XNOR U1781 ( .A(in[692]), .B(in[372]), .Z(n994) );
  XNOR U1782 ( .A(n995), .B(n994), .Z(n996) );
  XNOR U1783 ( .A(in[1012]), .B(n996), .Z(n1556) );
  XOR U1784 ( .A(in[821]), .B(in[501]), .Z(n998) );
  XNOR U1785 ( .A(in[1461]), .B(in[1141]), .Z(n997) );
  XNOR U1786 ( .A(n998), .B(n997), .Z(n999) );
  XNOR U1787 ( .A(in[181]), .B(n999), .Z(n1242) );
  XOR U1788 ( .A(n1556), .B(n1242), .Z(n4384) );
  XOR U1789 ( .A(in[1397]), .B(n4384), .Z(n5073) );
  NANDN U1790 ( .A(n5074), .B(n5073), .Z(n1000) );
  XOR U1791 ( .A(n1661), .B(n1000), .Z(out[1041]) );
  IV U1792 ( .A(n4063), .Z(n3408) );
  XOR U1793 ( .A(n3408), .B(in[549]), .Z(n1666) );
  XOR U1794 ( .A(in[853]), .B(in[1173]), .Z(n1002) );
  XNOR U1795 ( .A(in[1493]), .B(in[213]), .Z(n1001) );
  XNOR U1796 ( .A(n1002), .B(n1001), .Z(n1003) );
  XOR U1797 ( .A(in[533]), .B(n1003), .Z(n1445) );
  IV U1798 ( .A(n2758), .Z(n4016) );
  XNOR U1799 ( .A(in[149]), .B(n4016), .Z(n5077) );
  XOR U1800 ( .A(in[1333]), .B(in[53]), .Z(n1006) );
  XNOR U1801 ( .A(in[693]), .B(in[373]), .Z(n1005) );
  XNOR U1802 ( .A(n1006), .B(n1005), .Z(n1007) );
  XNOR U1803 ( .A(in[1013]), .B(n1007), .Z(n1560) );
  XOR U1804 ( .A(in[822]), .B(in[502]), .Z(n1009) );
  XNOR U1805 ( .A(in[1462]), .B(in[1142]), .Z(n1008) );
  XNOR U1806 ( .A(n1009), .B(n1008), .Z(n1010) );
  XNOR U1807 ( .A(in[182]), .B(n1010), .Z(n1257) );
  XOR U1808 ( .A(n1560), .B(n1257), .Z(n4387) );
  XOR U1809 ( .A(in[1398]), .B(n4387), .Z(n5076) );
  NANDN U1810 ( .A(n5077), .B(n5076), .Z(n1011) );
  XOR U1811 ( .A(n1666), .B(n1011), .Z(out[1042]) );
  XOR U1812 ( .A(n1013), .B(n1012), .Z(n2033) );
  XOR U1813 ( .A(in[550]), .B(n2033), .Z(n1670) );
  XOR U1814 ( .A(in[854]), .B(in[1174]), .Z(n1015) );
  XNOR U1815 ( .A(in[1494]), .B(in[214]), .Z(n1014) );
  XNOR U1816 ( .A(n1015), .B(n1014), .Z(n1016) );
  XOR U1817 ( .A(in[534]), .B(n1016), .Z(n1447) );
  XOR U1818 ( .A(in[150]), .B(n2775), .Z(n5081) );
  XOR U1819 ( .A(in[1334]), .B(in[54]), .Z(n1019) );
  XNOR U1820 ( .A(in[694]), .B(in[374]), .Z(n1018) );
  XNOR U1821 ( .A(n1019), .B(n1018), .Z(n1020) );
  XNOR U1822 ( .A(in[1014]), .B(n1020), .Z(n1564) );
  XOR U1823 ( .A(in[823]), .B(in[503]), .Z(n1022) );
  XNOR U1824 ( .A(in[1463]), .B(in[1143]), .Z(n1021) );
  XNOR U1825 ( .A(n1022), .B(n1021), .Z(n1023) );
  XNOR U1826 ( .A(in[183]), .B(n1023), .Z(n1269) );
  XOR U1827 ( .A(n1564), .B(n1269), .Z(n4390) );
  XOR U1828 ( .A(in[1399]), .B(n4390), .Z(n5078) );
  NANDN U1829 ( .A(n5081), .B(n5078), .Z(n1024) );
  XNOR U1830 ( .A(n1670), .B(n1024), .Z(out[1043]) );
  XOR U1831 ( .A(n1026), .B(n1025), .Z(n2035) );
  XOR U1832 ( .A(in[551]), .B(n2035), .Z(n1674) );
  XOR U1833 ( .A(in[855]), .B(in[1175]), .Z(n1028) );
  XNOR U1834 ( .A(in[1495]), .B(in[215]), .Z(n1027) );
  XNOR U1835 ( .A(n1028), .B(n1027), .Z(n1029) );
  XOR U1836 ( .A(in[535]), .B(n1029), .Z(n1449) );
  XOR U1837 ( .A(in[151]), .B(n2782), .Z(n5088) );
  XOR U1838 ( .A(in[1335]), .B(in[55]), .Z(n1032) );
  XNOR U1839 ( .A(in[695]), .B(in[375]), .Z(n1031) );
  XNOR U1840 ( .A(n1032), .B(n1031), .Z(n1033) );
  XNOR U1841 ( .A(in[1015]), .B(n1033), .Z(n1568) );
  XOR U1842 ( .A(in[824]), .B(in[504]), .Z(n1035) );
  XNOR U1843 ( .A(in[1464]), .B(in[1144]), .Z(n1034) );
  XNOR U1844 ( .A(n1035), .B(n1034), .Z(n1036) );
  XNOR U1845 ( .A(in[184]), .B(n1036), .Z(n1275) );
  XOR U1846 ( .A(n1568), .B(n1275), .Z(n4392) );
  XOR U1847 ( .A(in[1400]), .B(n4392), .Z(n5087) );
  NANDN U1848 ( .A(n5088), .B(n5087), .Z(n1037) );
  XNOR U1849 ( .A(n1674), .B(n1037), .Z(out[1044]) );
  XOR U1850 ( .A(n1039), .B(n1038), .Z(n2039) );
  XOR U1851 ( .A(in[552]), .B(n2039), .Z(n1678) );
  XOR U1852 ( .A(in[856]), .B(in[1176]), .Z(n1041) );
  XNOR U1853 ( .A(in[1496]), .B(in[216]), .Z(n1040) );
  XNOR U1854 ( .A(n1041), .B(n1040), .Z(n1042) );
  XOR U1855 ( .A(in[536]), .B(n1042), .Z(n1453) );
  XOR U1856 ( .A(in[152]), .B(n2796), .Z(n5091) );
  XOR U1857 ( .A(in[825]), .B(in[505]), .Z(n1045) );
  XNOR U1858 ( .A(in[1465]), .B(in[1145]), .Z(n1044) );
  XNOR U1859 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U1860 ( .A(in[185]), .B(n1046), .Z(n1287) );
  XOR U1861 ( .A(in[1336]), .B(in[56]), .Z(n1048) );
  XNOR U1862 ( .A(in[696]), .B(in[376]), .Z(n1047) );
  XNOR U1863 ( .A(n1048), .B(n1047), .Z(n1049) );
  XNOR U1864 ( .A(in[1016]), .B(n1049), .Z(n1572) );
  XOR U1865 ( .A(n1287), .B(n1572), .Z(n4395) );
  XOR U1866 ( .A(in[1401]), .B(n4395), .Z(n5090) );
  NANDN U1867 ( .A(n5091), .B(n5090), .Z(n1050) );
  XNOR U1868 ( .A(n1678), .B(n1050), .Z(out[1045]) );
  XOR U1869 ( .A(n1052), .B(n1051), .Z(n2041) );
  XOR U1870 ( .A(in[553]), .B(n2041), .Z(n1682) );
  XOR U1871 ( .A(in[857]), .B(in[1177]), .Z(n1054) );
  XNOR U1872 ( .A(in[1497]), .B(in[217]), .Z(n1053) );
  XNOR U1873 ( .A(n1054), .B(n1053), .Z(n1055) );
  XOR U1874 ( .A(in[537]), .B(n1055), .Z(n1455) );
  XOR U1875 ( .A(in[153]), .B(n2819), .Z(n5094) );
  XOR U1876 ( .A(in[1337]), .B(in[57]), .Z(n1058) );
  XNOR U1877 ( .A(in[697]), .B(in[377]), .Z(n1057) );
  XNOR U1878 ( .A(n1058), .B(n1057), .Z(n1059) );
  XNOR U1879 ( .A(in[1017]), .B(n1059), .Z(n1576) );
  XOR U1880 ( .A(in[826]), .B(in[506]), .Z(n1061) );
  XNOR U1881 ( .A(in[1466]), .B(in[1146]), .Z(n1060) );
  XNOR U1882 ( .A(n1061), .B(n1060), .Z(n1062) );
  XNOR U1883 ( .A(in[186]), .B(n1062), .Z(n1299) );
  XOR U1884 ( .A(n1576), .B(n1299), .Z(n2112) );
  IV U1885 ( .A(n2112), .Z(n4398) );
  XNOR U1886 ( .A(in[1402]), .B(n4398), .Z(n5093) );
  NANDN U1887 ( .A(n5094), .B(n5093), .Z(n1063) );
  XNOR U1888 ( .A(n1682), .B(n1063), .Z(out[1046]) );
  XOR U1889 ( .A(n1065), .B(n1064), .Z(n2043) );
  XOR U1890 ( .A(in[554]), .B(n2043), .Z(n1686) );
  XOR U1891 ( .A(in[858]), .B(in[1178]), .Z(n1067) );
  XNOR U1892 ( .A(in[1498]), .B(in[218]), .Z(n1066) );
  XNOR U1893 ( .A(n1067), .B(n1066), .Z(n1068) );
  XOR U1894 ( .A(in[538]), .B(n1068), .Z(n1457) );
  XOR U1895 ( .A(in[154]), .B(n2842), .Z(n5097) );
  XOR U1896 ( .A(in[1338]), .B(in[58]), .Z(n1071) );
  XNOR U1897 ( .A(in[698]), .B(in[378]), .Z(n1070) );
  XNOR U1898 ( .A(n1071), .B(n1070), .Z(n1072) );
  XNOR U1899 ( .A(in[1018]), .B(n1072), .Z(n1580) );
  XOR U1900 ( .A(in[827]), .B(in[507]), .Z(n1074) );
  XNOR U1901 ( .A(in[1467]), .B(in[1147]), .Z(n1073) );
  XNOR U1902 ( .A(n1074), .B(n1073), .Z(n1075) );
  XNOR U1903 ( .A(in[187]), .B(n1075), .Z(n1303) );
  XOR U1904 ( .A(n1580), .B(n1303), .Z(n2116) );
  IV U1905 ( .A(n2116), .Z(n4401) );
  XNOR U1906 ( .A(in[1403]), .B(n4401), .Z(n5096) );
  NANDN U1907 ( .A(n5097), .B(n5096), .Z(n1076) );
  XNOR U1908 ( .A(n1686), .B(n1076), .Z(out[1047]) );
  XOR U1909 ( .A(in[1579]), .B(in[619]), .Z(n1078) );
  XNOR U1910 ( .A(in[939]), .B(in[299]), .Z(n1077) );
  XNOR U1911 ( .A(n1078), .B(n1077), .Z(n1079) );
  XNOR U1912 ( .A(in[1259]), .B(n1079), .Z(n1590) );
  XNOR U1913 ( .A(n1080), .B(n1590), .Z(n3432) );
  IV U1914 ( .A(n3432), .Z(n4092) );
  XOR U1915 ( .A(in[555]), .B(n4092), .Z(n1690) );
  XOR U1916 ( .A(in[859]), .B(in[1179]), .Z(n1082) );
  XNOR U1917 ( .A(in[1499]), .B(in[219]), .Z(n1081) );
  XNOR U1918 ( .A(n1082), .B(n1081), .Z(n1083) );
  XOR U1919 ( .A(in[539]), .B(n1083), .Z(n1461) );
  XOR U1920 ( .A(in[155]), .B(n2866), .Z(n5100) );
  XOR U1921 ( .A(in[828]), .B(in[508]), .Z(n1086) );
  XNOR U1922 ( .A(in[1468]), .B(in[1148]), .Z(n1085) );
  XNOR U1923 ( .A(n1086), .B(n1085), .Z(n1087) );
  XNOR U1924 ( .A(in[188]), .B(n1087), .Z(n1307) );
  XOR U1925 ( .A(n1088), .B(n1307), .Z(n4404) );
  XOR U1926 ( .A(in[1404]), .B(n4404), .Z(n5099) );
  NANDN U1927 ( .A(n5100), .B(n5099), .Z(n1089) );
  XNOR U1928 ( .A(n1690), .B(n1089), .Z(out[1048]) );
  XOR U1929 ( .A(in[1580]), .B(in[620]), .Z(n1091) );
  XNOR U1930 ( .A(in[940]), .B(in[300]), .Z(n1090) );
  XNOR U1931 ( .A(n1091), .B(n1090), .Z(n1092) );
  XNOR U1932 ( .A(in[1260]), .B(n1092), .Z(n1594) );
  XNOR U1933 ( .A(n1093), .B(n1594), .Z(n3435) );
  IV U1934 ( .A(n3435), .Z(n4096) );
  XOR U1935 ( .A(in[556]), .B(n4096), .Z(n1694) );
  XOR U1936 ( .A(in[860]), .B(in[1180]), .Z(n1095) );
  XNOR U1937 ( .A(in[1500]), .B(in[220]), .Z(n1094) );
  XNOR U1938 ( .A(n1095), .B(n1094), .Z(n1096) );
  XOR U1939 ( .A(in[540]), .B(n1096), .Z(n1467) );
  XOR U1940 ( .A(in[156]), .B(n2890), .Z(n5103) );
  XOR U1941 ( .A(n1099), .B(n1098), .Z(n4411) );
  XOR U1942 ( .A(in[1405]), .B(n4411), .Z(n5102) );
  NANDN U1943 ( .A(n5103), .B(n5102), .Z(n1100) );
  XNOR U1944 ( .A(n1694), .B(n1100), .Z(out[1049]) );
  XOR U1945 ( .A(in[1343]), .B(in[63]), .Z(n1102) );
  XNOR U1946 ( .A(in[703]), .B(in[383]), .Z(n1101) );
  XNOR U1947 ( .A(n1102), .B(n1101), .Z(n1103) );
  XNOR U1948 ( .A(in[1023]), .B(n1103), .Z(n1147) );
  XOR U1949 ( .A(n1104), .B(n1147), .Z(n3971) );
  XOR U1950 ( .A(in[639]), .B(n3971), .Z(n2714) );
  IV U1951 ( .A(n2714), .Z(n2803) );
  XNOR U1952 ( .A(in[230]), .B(n2033), .Z(n3196) );
  XOR U1953 ( .A(in[874]), .B(in[1194]), .Z(n1106) );
  XNOR U1954 ( .A(in[1514]), .B(in[234]), .Z(n1105) );
  XNOR U1955 ( .A(n1106), .B(n1105), .Z(n1107) );
  XNOR U1956 ( .A(in[554]), .B(n1107), .Z(n1518) );
  XNOR U1957 ( .A(n1108), .B(n1518), .Z(n4107) );
  IV U1958 ( .A(n4107), .Z(n1288) );
  XOR U1959 ( .A(in[1450]), .B(n1288), .Z(n3193) );
  NAND U1960 ( .A(n3196), .B(n3193), .Z(n1109) );
  XOR U1961 ( .A(n2803), .B(n1109), .Z(out[104]) );
  XOR U1962 ( .A(in[1581]), .B(in[621]), .Z(n1111) );
  XNOR U1963 ( .A(in[941]), .B(in[301]), .Z(n1110) );
  XNOR U1964 ( .A(n1111), .B(n1110), .Z(n1112) );
  XNOR U1965 ( .A(in[1261]), .B(n1112), .Z(n1598) );
  XNOR U1966 ( .A(n1113), .B(n1598), .Z(n3438) );
  IV U1967 ( .A(n3438), .Z(n4100) );
  XOR U1968 ( .A(in[557]), .B(n4100), .Z(n1698) );
  XOR U1969 ( .A(in[861]), .B(in[1181]), .Z(n1115) );
  XNOR U1970 ( .A(in[1501]), .B(in[221]), .Z(n1114) );
  XNOR U1971 ( .A(n1115), .B(n1114), .Z(n1116) );
  XOR U1972 ( .A(in[541]), .B(n1116), .Z(n1471) );
  XOR U1973 ( .A(in[157]), .B(n2923), .Z(n5106) );
  XOR U1974 ( .A(in[830]), .B(in[510]), .Z(n1119) );
  XNOR U1975 ( .A(in[1470]), .B(in[1150]), .Z(n1118) );
  XNOR U1976 ( .A(n1119), .B(n1118), .Z(n1120) );
  XNOR U1977 ( .A(in[190]), .B(n1120), .Z(n1311) );
  XOR U1978 ( .A(n1121), .B(n1311), .Z(n4414) );
  XOR U1979 ( .A(in[1406]), .B(n4414), .Z(n5105) );
  NANDN U1980 ( .A(n5106), .B(n5105), .Z(n1122) );
  XNOR U1981 ( .A(n1698), .B(n1122), .Z(out[1050]) );
  XOR U1982 ( .A(in[1582]), .B(in[622]), .Z(n1124) );
  XNOR U1983 ( .A(in[942]), .B(in[302]), .Z(n1123) );
  XNOR U1984 ( .A(n1124), .B(n1123), .Z(n1125) );
  XNOR U1985 ( .A(in[1262]), .B(n1125), .Z(n1602) );
  XNOR U1986 ( .A(n1126), .B(n1602), .Z(n3441) );
  IV U1987 ( .A(n3441), .Z(n4104) );
  XOR U1988 ( .A(in[558]), .B(n4104), .Z(n1702) );
  XOR U1989 ( .A(in[862]), .B(in[1182]), .Z(n1128) );
  XNOR U1990 ( .A(in[1502]), .B(in[222]), .Z(n1127) );
  XNOR U1991 ( .A(n1128), .B(n1127), .Z(n1129) );
  XOR U1992 ( .A(in[542]), .B(n1129), .Z(n1475) );
  XNOR U1993 ( .A(in[158]), .B(n4056), .Z(n1451) );
  IV U1994 ( .A(n1451), .Z(n5109) );
  XOR U1995 ( .A(in[831]), .B(in[511]), .Z(n1132) );
  XNOR U1996 ( .A(in[1471]), .B(in[1151]), .Z(n1131) );
  XNOR U1997 ( .A(n1132), .B(n1131), .Z(n1133) );
  XNOR U1998 ( .A(in[191]), .B(n1133), .Z(n1315) );
  XOR U1999 ( .A(n1134), .B(n1315), .Z(n4417) );
  XOR U2000 ( .A(in[1407]), .B(n4417), .Z(n5108) );
  NANDN U2001 ( .A(n5109), .B(n5108), .Z(n1135) );
  XNOR U2002 ( .A(n1702), .B(n1135), .Z(out[1051]) );
  XOR U2003 ( .A(in[1583]), .B(in[623]), .Z(n1137) );
  XNOR U2004 ( .A(in[943]), .B(in[303]), .Z(n1136) );
  XNOR U2005 ( .A(n1137), .B(n1136), .Z(n1138) );
  XNOR U2006 ( .A(in[1263]), .B(n1138), .Z(n1606) );
  XNOR U2007 ( .A(n1139), .B(n1606), .Z(n3444) );
  IV U2008 ( .A(n3444), .Z(n4108) );
  XOR U2009 ( .A(in[559]), .B(n4108), .Z(n1708) );
  XOR U2010 ( .A(in[863]), .B(in[1183]), .Z(n1141) );
  XNOR U2011 ( .A(in[1503]), .B(in[223]), .Z(n1140) );
  XNOR U2012 ( .A(n1141), .B(n1140), .Z(n1142) );
  XOR U2013 ( .A(in[543]), .B(n1142), .Z(n1477) );
  XOR U2014 ( .A(in[159]), .B(n4060), .Z(n5113) );
  XOR U2015 ( .A(in[768]), .B(in[1088]), .Z(n1145) );
  XNOR U2016 ( .A(in[448]), .B(in[1408]), .Z(n1144) );
  XNOR U2017 ( .A(n1145), .B(n1144), .Z(n1146) );
  XNOR U2018 ( .A(in[128]), .B(n1146), .Z(n1322) );
  XOR U2019 ( .A(n1147), .B(n1322), .Z(n4420) );
  XOR U2020 ( .A(in[1344]), .B(n4420), .Z(n5110) );
  NANDN U2021 ( .A(n5113), .B(n5110), .Z(n1148) );
  XNOR U2022 ( .A(n1708), .B(n1148), .Z(out[1052]) );
  XOR U2023 ( .A(in[1584]), .B(in[624]), .Z(n1150) );
  XNOR U2024 ( .A(in[944]), .B(in[304]), .Z(n1149) );
  XNOR U2025 ( .A(n1150), .B(n1149), .Z(n1151) );
  XNOR U2026 ( .A(in[1264]), .B(n1151), .Z(n1610) );
  XNOR U2027 ( .A(n1152), .B(n1610), .Z(n3447) );
  IV U2028 ( .A(n3447), .Z(n4112) );
  XOR U2029 ( .A(in[560]), .B(n4112), .Z(n1712) );
  XOR U2030 ( .A(in[224]), .B(in[864]), .Z(n1154) );
  XNOR U2031 ( .A(in[1184]), .B(in[1504]), .Z(n1153) );
  XNOR U2032 ( .A(n1154), .B(n1153), .Z(n1155) );
  XOR U2033 ( .A(in[544]), .B(n1155), .Z(n1480) );
  XOR U2034 ( .A(in[160]), .B(n4064), .Z(n5116) );
  XOR U2035 ( .A(in[1280]), .B(in[640]), .Z(n1158) );
  XNOR U2036 ( .A(in[960]), .B(in[320]), .Z(n1157) );
  XNOR U2037 ( .A(n1158), .B(n1157), .Z(n1159) );
  XNOR U2038 ( .A(in[0]), .B(n1159), .Z(n1251) );
  XOR U2039 ( .A(in[769]), .B(in[1089]), .Z(n1161) );
  XNOR U2040 ( .A(in[449]), .B(in[1409]), .Z(n1160) );
  XNOR U2041 ( .A(n1161), .B(n1160), .Z(n1162) );
  XNOR U2042 ( .A(in[129]), .B(n1162), .Z(n1326) );
  XOR U2043 ( .A(n1251), .B(n1326), .Z(n4423) );
  XOR U2044 ( .A(in[1345]), .B(n4423), .Z(n5115) );
  NANDN U2045 ( .A(n5116), .B(n5115), .Z(n1163) );
  XNOR U2046 ( .A(n1712), .B(n1163), .Z(out[1053]) );
  XOR U2047 ( .A(in[1585]), .B(in[625]), .Z(n1165) );
  XNOR U2048 ( .A(in[945]), .B(in[305]), .Z(n1164) );
  XNOR U2049 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U2050 ( .A(in[1265]), .B(n1166), .Z(n1614) );
  XNOR U2051 ( .A(n1167), .B(n1614), .Z(n3450) );
  IV U2052 ( .A(n3450), .Z(n4120) );
  XOR U2053 ( .A(in[561]), .B(n4120), .Z(n1716) );
  XOR U2054 ( .A(in[225]), .B(in[865]), .Z(n1169) );
  XNOR U2055 ( .A(in[1185]), .B(in[1505]), .Z(n1168) );
  XNOR U2056 ( .A(n1169), .B(n1168), .Z(n1170) );
  XOR U2057 ( .A(in[545]), .B(n1170), .Z(n1483) );
  XNOR U2058 ( .A(in[161]), .B(n4068), .Z(n1459) );
  IV U2059 ( .A(n1459), .Z(n5123) );
  XOR U2060 ( .A(in[1]), .B(in[641]), .Z(n1173) );
  XNOR U2061 ( .A(in[961]), .B(in[321]), .Z(n1172) );
  XNOR U2062 ( .A(n1173), .B(n1172), .Z(n1174) );
  XNOR U2063 ( .A(in[1281]), .B(n1174), .Z(n1316) );
  XOR U2064 ( .A(in[1090]), .B(in[450]), .Z(n1176) );
  XNOR U2065 ( .A(in[130]), .B(in[770]), .Z(n1175) );
  XNOR U2066 ( .A(n1176), .B(n1175), .Z(n1177) );
  XNOR U2067 ( .A(in[1410]), .B(n1177), .Z(n1330) );
  XOR U2068 ( .A(n1316), .B(n1330), .Z(n4426) );
  XOR U2069 ( .A(in[1346]), .B(n4426), .Z(n5122) );
  NANDN U2070 ( .A(n5123), .B(n5122), .Z(n1178) );
  XNOR U2071 ( .A(n1716), .B(n1178), .Z(out[1054]) );
  XOR U2072 ( .A(in[1586]), .B(in[626]), .Z(n1180) );
  XNOR U2073 ( .A(in[946]), .B(in[306]), .Z(n1179) );
  XNOR U2074 ( .A(n1180), .B(n1179), .Z(n1181) );
  XNOR U2075 ( .A(in[1266]), .B(n1181), .Z(n1618) );
  XNOR U2076 ( .A(n1182), .B(n1618), .Z(n3453) );
  IV U2077 ( .A(n3453), .Z(n4124) );
  XOR U2078 ( .A(in[562]), .B(n4124), .Z(n1720) );
  XOR U2079 ( .A(in[1186]), .B(in[1506]), .Z(n1184) );
  XNOR U2080 ( .A(in[546]), .B(in[866]), .Z(n1183) );
  XNOR U2081 ( .A(n1184), .B(n1183), .Z(n1185) );
  XOR U2082 ( .A(in[226]), .B(n1185), .Z(n1486) );
  XNOR U2083 ( .A(in[162]), .B(n4076), .Z(n1463) );
  IV U2084 ( .A(n1463), .Z(n5127) );
  XOR U2085 ( .A(in[771]), .B(in[1091]), .Z(n1188) );
  XNOR U2086 ( .A(in[451]), .B(in[1411]), .Z(n1187) );
  XNOR U2087 ( .A(n1188), .B(n1187), .Z(n1189) );
  XNOR U2088 ( .A(in[131]), .B(n1189), .Z(n1334) );
  XOR U2089 ( .A(in[2]), .B(in[642]), .Z(n1191) );
  XNOR U2090 ( .A(in[962]), .B(in[322]), .Z(n1190) );
  XNOR U2091 ( .A(n1191), .B(n1190), .Z(n1192) );
  XNOR U2092 ( .A(in[1282]), .B(n1192), .Z(n1361) );
  XOR U2093 ( .A(n1334), .B(n1361), .Z(n4429) );
  XOR U2094 ( .A(in[1347]), .B(n4429), .Z(n5124) );
  NANDN U2095 ( .A(n5127), .B(n5124), .Z(n1193) );
  XNOR U2096 ( .A(n1720), .B(n1193), .Z(out[1055]) );
  XOR U2097 ( .A(in[1587]), .B(in[627]), .Z(n1195) );
  XNOR U2098 ( .A(in[947]), .B(in[307]), .Z(n1194) );
  XNOR U2099 ( .A(n1195), .B(n1194), .Z(n1196) );
  XNOR U2100 ( .A(in[1267]), .B(n1196), .Z(n1623) );
  XNOR U2101 ( .A(n1197), .B(n1623), .Z(n3456) );
  IV U2102 ( .A(n3456), .Z(n4128) );
  XOR U2103 ( .A(in[563]), .B(n4128), .Z(n1724) );
  XOR U2104 ( .A(in[1187]), .B(in[1507]), .Z(n1199) );
  XNOR U2105 ( .A(in[547]), .B(in[867]), .Z(n1198) );
  XNOR U2106 ( .A(n1199), .B(n1198), .Z(n1200) );
  XOR U2107 ( .A(in[227]), .B(n1200), .Z(n1489) );
  XNOR U2108 ( .A(in[163]), .B(n4080), .Z(n1469) );
  IV U2109 ( .A(n1469), .Z(n5131) );
  XOR U2110 ( .A(in[772]), .B(in[1092]), .Z(n1203) );
  XNOR U2111 ( .A(in[452]), .B(in[1412]), .Z(n1202) );
  XNOR U2112 ( .A(n1203), .B(n1202), .Z(n1204) );
  XNOR U2113 ( .A(in[132]), .B(n1204), .Z(n1338) );
  XOR U2114 ( .A(in[323]), .B(in[643]), .Z(n1206) );
  XNOR U2115 ( .A(in[963]), .B(in[3]), .Z(n1205) );
  XNOR U2116 ( .A(n1206), .B(n1205), .Z(n1207) );
  XNOR U2117 ( .A(in[1283]), .B(n1207), .Z(n1402) );
  XOR U2118 ( .A(n1338), .B(n1402), .Z(n4432) );
  XOR U2119 ( .A(in[1348]), .B(n4432), .Z(n5128) );
  NANDN U2120 ( .A(n5131), .B(n5128), .Z(n1208) );
  XNOR U2121 ( .A(n1724), .B(n1208), .Z(out[1056]) );
  XOR U2122 ( .A(in[1588]), .B(in[628]), .Z(n1210) );
  XNOR U2123 ( .A(in[948]), .B(in[308]), .Z(n1209) );
  XNOR U2124 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U2125 ( .A(in[1268]), .B(n1211), .Z(n1627) );
  XNOR U2126 ( .A(n1212), .B(n1627), .Z(n3463) );
  IV U2127 ( .A(n3463), .Z(n4132) );
  XOR U2128 ( .A(in[564]), .B(n4132), .Z(n1728) );
  XOR U2129 ( .A(in[1188]), .B(in[1508]), .Z(n1214) );
  XNOR U2130 ( .A(in[548]), .B(in[868]), .Z(n1213) );
  XNOR U2131 ( .A(n1214), .B(n1213), .Z(n1215) );
  XNOR U2132 ( .A(in[228]), .B(n1215), .Z(n1492) );
  XNOR U2133 ( .A(in[164]), .B(n4084), .Z(n1473) );
  IV U2134 ( .A(n1473), .Z(n5135) );
  XOR U2135 ( .A(in[324]), .B(in[644]), .Z(n1218) );
  XNOR U2136 ( .A(in[964]), .B(in[4]), .Z(n1217) );
  XNOR U2137 ( .A(n1218), .B(n1217), .Z(n1219) );
  XNOR U2138 ( .A(in[1284]), .B(n1219), .Z(n1406) );
  XOR U2139 ( .A(in[773]), .B(in[1093]), .Z(n1221) );
  XNOR U2140 ( .A(in[453]), .B(in[1413]), .Z(n1220) );
  XNOR U2141 ( .A(n1221), .B(n1220), .Z(n1222) );
  XNOR U2142 ( .A(in[133]), .B(n1222), .Z(n1342) );
  XOR U2143 ( .A(n1406), .B(n1342), .Z(n4435) );
  XOR U2144 ( .A(in[1349]), .B(n4435), .Z(n5132) );
  NANDN U2145 ( .A(n5135), .B(n5132), .Z(n1223) );
  XNOR U2146 ( .A(n1728), .B(n1223), .Z(out[1057]) );
  XOR U2147 ( .A(in[1589]), .B(in[629]), .Z(n1225) );
  XNOR U2148 ( .A(in[949]), .B(in[309]), .Z(n1224) );
  XNOR U2149 ( .A(n1225), .B(n1224), .Z(n1226) );
  XNOR U2150 ( .A(in[1269]), .B(n1226), .Z(n1631) );
  XNOR U2151 ( .A(n1227), .B(n1631), .Z(n3466) );
  IV U2152 ( .A(n3466), .Z(n4136) );
  XOR U2153 ( .A(in[565]), .B(n4136), .Z(n1732) );
  XOR U2154 ( .A(in[1189]), .B(in[1509]), .Z(n1229) );
  XNOR U2155 ( .A(in[549]), .B(in[869]), .Z(n1228) );
  XNOR U2156 ( .A(n1229), .B(n1228), .Z(n1230) );
  XOR U2157 ( .A(in[229]), .B(n1230), .Z(n1496) );
  XOR U2158 ( .A(in[165]), .B(n2215), .Z(n5139) );
  XOR U2159 ( .A(in[774]), .B(in[1094]), .Z(n1233) );
  XNOR U2160 ( .A(in[454]), .B(in[1414]), .Z(n1232) );
  XNOR U2161 ( .A(n1233), .B(n1232), .Z(n1234) );
  XNOR U2162 ( .A(in[134]), .B(n1234), .Z(n1346) );
  XOR U2163 ( .A(in[325]), .B(in[645]), .Z(n1236) );
  XNOR U2164 ( .A(in[965]), .B(in[5]), .Z(n1235) );
  XNOR U2165 ( .A(n1236), .B(n1235), .Z(n1237) );
  XNOR U2166 ( .A(in[1285]), .B(n1237), .Z(n1408) );
  XOR U2167 ( .A(n1346), .B(n1408), .Z(n2128) );
  IV U2168 ( .A(n2128), .Z(n4438) );
  XNOR U2169 ( .A(in[1350]), .B(n4438), .Z(n5136) );
  NANDN U2170 ( .A(n5139), .B(n5136), .Z(n1238) );
  XNOR U2171 ( .A(n1732), .B(n1238), .Z(out[1058]) );
  XOR U2172 ( .A(in[1590]), .B(in[630]), .Z(n1240) );
  XNOR U2173 ( .A(in[950]), .B(in[310]), .Z(n1239) );
  XNOR U2174 ( .A(n1240), .B(n1239), .Z(n1241) );
  XNOR U2175 ( .A(in[1270]), .B(n1241), .Z(n1635) );
  XNOR U2176 ( .A(n1242), .B(n1635), .Z(n3263) );
  IV U2177 ( .A(n3263), .Z(n4140) );
  XOR U2178 ( .A(in[566]), .B(n4140), .Z(n1736) );
  XNOR U2179 ( .A(in[166]), .B(n1243), .Z(n5143) );
  XOR U2180 ( .A(in[775]), .B(in[1095]), .Z(n1245) );
  XNOR U2181 ( .A(in[455]), .B(in[1415]), .Z(n1244) );
  XNOR U2182 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U2183 ( .A(in[135]), .B(n1246), .Z(n1350) );
  XOR U2184 ( .A(in[326]), .B(in[6]), .Z(n1248) );
  XNOR U2185 ( .A(in[966]), .B(in[646]), .Z(n1247) );
  XNOR U2186 ( .A(n1248), .B(n1247), .Z(n1249) );
  XNOR U2187 ( .A(in[1286]), .B(n1249), .Z(n1410) );
  XOR U2188 ( .A(n1350), .B(n1410), .Z(n4449) );
  XOR U2189 ( .A(in[1351]), .B(n4449), .Z(n5140) );
  NAND U2190 ( .A(n5143), .B(n5140), .Z(n1250) );
  XNOR U2191 ( .A(n1736), .B(n1250), .Z(out[1059]) );
  XOR U2192 ( .A(n1252), .B(n1251), .Z(n3975) );
  XOR U2193 ( .A(in[576]), .B(n3975), .Z(n2716) );
  IV U2194 ( .A(n2716), .Z(n2805) );
  XNOR U2195 ( .A(in[1451]), .B(n4111), .Z(n3224) );
  XNOR U2196 ( .A(in[231]), .B(n2035), .Z(n3226) );
  NANDN U2197 ( .A(n3224), .B(n3226), .Z(n1253) );
  XOR U2198 ( .A(n2805), .B(n1253), .Z(out[105]) );
  XOR U2199 ( .A(in[1591]), .B(in[631]), .Z(n1255) );
  XNOR U2200 ( .A(in[951]), .B(in[311]), .Z(n1254) );
  XNOR U2201 ( .A(n1255), .B(n1254), .Z(n1256) );
  XNOR U2202 ( .A(in[1271]), .B(n1256), .Z(n1639) );
  XNOR U2203 ( .A(n1257), .B(n1639), .Z(n3266) );
  IV U2204 ( .A(n3266), .Z(n4144) );
  XOR U2205 ( .A(in[567]), .B(n4144), .Z(n1740) );
  XNOR U2206 ( .A(in[167]), .B(n1258), .Z(n5147) );
  XOR U2207 ( .A(in[327]), .B(in[7]), .Z(n1260) );
  XNOR U2208 ( .A(in[967]), .B(in[647]), .Z(n1259) );
  XNOR U2209 ( .A(n1260), .B(n1259), .Z(n1261) );
  XNOR U2210 ( .A(in[1287]), .B(n1261), .Z(n1412) );
  XOR U2211 ( .A(in[776]), .B(in[1096]), .Z(n1263) );
  XNOR U2212 ( .A(in[456]), .B(in[1416]), .Z(n1262) );
  XNOR U2213 ( .A(n1263), .B(n1262), .Z(n1264) );
  XNOR U2214 ( .A(in[136]), .B(n1264), .Z(n1354) );
  XOR U2215 ( .A(n1412), .B(n1354), .Z(n4452) );
  XOR U2216 ( .A(in[1352]), .B(n4452), .Z(n5144) );
  NAND U2217 ( .A(n5147), .B(n5144), .Z(n1265) );
  XNOR U2218 ( .A(n1740), .B(n1265), .Z(out[1060]) );
  XOR U2219 ( .A(in[632]), .B(in[1592]), .Z(n1267) );
  XNOR U2220 ( .A(in[1272]), .B(in[312]), .Z(n1266) );
  XNOR U2221 ( .A(n1267), .B(n1266), .Z(n1268) );
  XNOR U2222 ( .A(in[952]), .B(n1268), .Z(n1643) );
  XNOR U2223 ( .A(n1269), .B(n1643), .Z(n3273) );
  IV U2224 ( .A(n3273), .Z(n4148) );
  XOR U2225 ( .A(in[568]), .B(n4148), .Z(n1744) );
  XNOR U2226 ( .A(in[168]), .B(n1270), .Z(n5151) );
  XOR U2227 ( .A(in[1353]), .B(n4455), .Z(n5148) );
  NAND U2228 ( .A(n5151), .B(n5148), .Z(n1271) );
  XNOR U2229 ( .A(n1744), .B(n1271), .Z(out[1061]) );
  XOR U2230 ( .A(in[633]), .B(in[1593]), .Z(n1273) );
  XNOR U2231 ( .A(in[1273]), .B(in[313]), .Z(n1272) );
  XNOR U2232 ( .A(n1273), .B(n1272), .Z(n1274) );
  XNOR U2233 ( .A(in[953]), .B(n1274), .Z(n1647) );
  XNOR U2234 ( .A(n1275), .B(n1647), .Z(n3276) );
  IV U2235 ( .A(n3276), .Z(n4152) );
  XOR U2236 ( .A(in[569]), .B(n4152), .Z(n1749) );
  XOR U2237 ( .A(in[778]), .B(in[1098]), .Z(n1277) );
  XNOR U2238 ( .A(in[458]), .B(in[1418]), .Z(n1276) );
  XNOR U2239 ( .A(n1277), .B(n1276), .Z(n1278) );
  XNOR U2240 ( .A(in[138]), .B(n1278), .Z(n1368) );
  XOR U2241 ( .A(in[329]), .B(in[969]), .Z(n1280) );
  XNOR U2242 ( .A(in[9]), .B(in[649]), .Z(n1279) );
  XNOR U2243 ( .A(n1280), .B(n1279), .Z(n1281) );
  XNOR U2244 ( .A(in[1289]), .B(n1281), .Z(n1419) );
  XOR U2245 ( .A(n1368), .B(n1419), .Z(n4458) );
  XNOR U2246 ( .A(in[1354]), .B(n4458), .Z(n5153) );
  XNOR U2247 ( .A(in[169]), .B(n1282), .Z(n5155) );
  NANDN U2248 ( .A(n5153), .B(n5155), .Z(n1283) );
  XNOR U2249 ( .A(n1749), .B(n1283), .Z(out[1062]) );
  XOR U2250 ( .A(in[634]), .B(in[1594]), .Z(n1285) );
  XNOR U2251 ( .A(in[1274]), .B(in[314]), .Z(n1284) );
  XNOR U2252 ( .A(n1285), .B(n1284), .Z(n1286) );
  XNOR U2253 ( .A(in[954]), .B(n1286), .Z(n1651) );
  XNOR U2254 ( .A(n1287), .B(n1651), .Z(n3279) );
  IV U2255 ( .A(n3279), .Z(n4156) );
  XOR U2256 ( .A(in[570]), .B(n4156), .Z(n1753) );
  XNOR U2257 ( .A(in[170]), .B(n1288), .Z(n5159) );
  XOR U2258 ( .A(in[1290]), .B(in[650]), .Z(n1290) );
  XNOR U2259 ( .A(in[970]), .B(in[330]), .Z(n1289) );
  XNOR U2260 ( .A(n1290), .B(n1289), .Z(n1291) );
  XNOR U2261 ( .A(in[10]), .B(n1291), .Z(n1421) );
  XOR U2262 ( .A(in[1419]), .B(in[779]), .Z(n1293) );
  XNOR U2263 ( .A(in[1099]), .B(in[459]), .Z(n1292) );
  XNOR U2264 ( .A(n1293), .B(n1292), .Z(n1294) );
  XNOR U2265 ( .A(in[139]), .B(n1294), .Z(n1374) );
  XOR U2266 ( .A(n1421), .B(n1374), .Z(n4461) );
  XOR U2267 ( .A(in[1355]), .B(n4461), .Z(n5156) );
  NAND U2268 ( .A(n5159), .B(n5156), .Z(n1295) );
  XNOR U2269 ( .A(n1753), .B(n1295), .Z(out[1063]) );
  XOR U2270 ( .A(in[955]), .B(in[1275]), .Z(n1297) );
  XNOR U2271 ( .A(in[1595]), .B(in[315]), .Z(n1296) );
  XNOR U2272 ( .A(n1297), .B(n1296), .Z(n1298) );
  XOR U2273 ( .A(in[635]), .B(n1298), .Z(n1655) );
  XOR U2274 ( .A(n1299), .B(n1655), .Z(n4166) );
  XOR U2275 ( .A(in[571]), .B(n4166), .Z(n1755) );
  XOR U2276 ( .A(in[956]), .B(in[1276]), .Z(n1301) );
  XNOR U2277 ( .A(in[1596]), .B(in[316]), .Z(n1300) );
  XNOR U2278 ( .A(n1301), .B(n1300), .Z(n1302) );
  XOR U2279 ( .A(in[636]), .B(n1302), .Z(n1659) );
  XOR U2280 ( .A(n1303), .B(n1659), .Z(n4170) );
  XOR U2281 ( .A(in[572]), .B(n4170), .Z(n1757) );
  XOR U2282 ( .A(in[957]), .B(in[1277]), .Z(n1305) );
  XNOR U2283 ( .A(in[1597]), .B(in[317]), .Z(n1304) );
  XNOR U2284 ( .A(n1305), .B(n1304), .Z(n1306) );
  XOR U2285 ( .A(in[637]), .B(n1306), .Z(n1664) );
  XOR U2286 ( .A(n1307), .B(n1664), .Z(n4174) );
  XOR U2287 ( .A(in[573]), .B(n4174), .Z(n1759) );
  IV U2288 ( .A(n3291), .Z(n4178) );
  XOR U2289 ( .A(in[574]), .B(n4178), .Z(n1761) );
  XOR U2290 ( .A(in[959]), .B(in[1279]), .Z(n1309) );
  XNOR U2291 ( .A(in[1599]), .B(in[319]), .Z(n1308) );
  XNOR U2292 ( .A(n1309), .B(n1308), .Z(n1310) );
  XOR U2293 ( .A(in[639]), .B(n1310), .Z(n1672) );
  XOR U2294 ( .A(n1311), .B(n1672), .Z(n3294) );
  XOR U2295 ( .A(in[575]), .B(n3294), .Z(n1762) );
  XOR U2296 ( .A(in[896]), .B(in[1216]), .Z(n1313) );
  XNOR U2297 ( .A(in[1536]), .B(in[256]), .Z(n1312) );
  XNOR U2298 ( .A(n1313), .B(n1312), .Z(n1314) );
  XOR U2299 ( .A(in[576]), .B(n1314), .Z(n1676) );
  XOR U2300 ( .A(n1315), .B(n1676), .Z(n3297) );
  XOR U2301 ( .A(in[512]), .B(n3297), .Z(n1764) );
  XOR U2302 ( .A(n1317), .B(n1316), .Z(n3979) );
  XOR U2303 ( .A(in[577]), .B(n3979), .Z(n2719) );
  IV U2304 ( .A(n2719), .Z(n2807) );
  XNOR U2305 ( .A(in[1452]), .B(n4119), .Z(n3248) );
  XNOR U2306 ( .A(in[232]), .B(n2039), .Z(n3250) );
  NANDN U2307 ( .A(n3248), .B(n3250), .Z(n1318) );
  XOR U2308 ( .A(n2807), .B(n1318), .Z(out[106]) );
  XOR U2309 ( .A(in[897]), .B(in[1217]), .Z(n1320) );
  XNOR U2310 ( .A(in[1537]), .B(in[257]), .Z(n1319) );
  XNOR U2311 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U2312 ( .A(in[577]), .B(n1321), .Z(n1680) );
  XOR U2313 ( .A(n1322), .B(n1680), .Z(n3300) );
  XOR U2314 ( .A(in[513]), .B(n3300), .Z(n1766) );
  XOR U2315 ( .A(in[1538]), .B(in[578]), .Z(n1324) );
  XNOR U2316 ( .A(in[898]), .B(in[258]), .Z(n1323) );
  XNOR U2317 ( .A(n1324), .B(n1323), .Z(n1325) );
  XOR U2318 ( .A(in[1218]), .B(n1325), .Z(n1684) );
  XOR U2319 ( .A(n1326), .B(n1684), .Z(n3307) );
  XOR U2320 ( .A(in[514]), .B(n3307), .Z(n1768) );
  XOR U2321 ( .A(in[1539]), .B(in[579]), .Z(n1328) );
  XNOR U2322 ( .A(in[899]), .B(in[259]), .Z(n1327) );
  XNOR U2323 ( .A(n1328), .B(n1327), .Z(n1329) );
  XOR U2324 ( .A(in[1219]), .B(n1329), .Z(n1688) );
  XOR U2325 ( .A(n1330), .B(n1688), .Z(n3310) );
  XOR U2326 ( .A(in[515]), .B(n3310), .Z(n1772) );
  XOR U2327 ( .A(in[1540]), .B(in[580]), .Z(n1332) );
  XNOR U2328 ( .A(in[900]), .B(in[260]), .Z(n1331) );
  XNOR U2329 ( .A(n1332), .B(n1331), .Z(n1333) );
  XOR U2330 ( .A(in[1220]), .B(n1333), .Z(n1692) );
  XOR U2331 ( .A(n1334), .B(n1692), .Z(n3313) );
  XOR U2332 ( .A(in[516]), .B(n3313), .Z(n1774) );
  XOR U2333 ( .A(in[1541]), .B(in[581]), .Z(n1336) );
  XNOR U2334 ( .A(in[901]), .B(in[261]), .Z(n1335) );
  XNOR U2335 ( .A(n1336), .B(n1335), .Z(n1337) );
  XOR U2336 ( .A(in[1221]), .B(n1337), .Z(n1696) );
  XOR U2337 ( .A(n1338), .B(n1696), .Z(n3316) );
  XOR U2338 ( .A(in[517]), .B(n3316), .Z(n1776) );
  XOR U2339 ( .A(in[1542]), .B(in[582]), .Z(n1340) );
  XNOR U2340 ( .A(in[902]), .B(in[262]), .Z(n1339) );
  XNOR U2341 ( .A(n1340), .B(n1339), .Z(n1341) );
  XOR U2342 ( .A(in[1222]), .B(n1341), .Z(n1700) );
  XOR U2343 ( .A(n1342), .B(n1700), .Z(n3319) );
  XOR U2344 ( .A(in[518]), .B(n3319), .Z(n1778) );
  XOR U2345 ( .A(in[1543]), .B(in[583]), .Z(n1344) );
  XNOR U2346 ( .A(in[903]), .B(in[263]), .Z(n1343) );
  XNOR U2347 ( .A(n1344), .B(n1343), .Z(n1345) );
  XOR U2348 ( .A(in[1223]), .B(n1345), .Z(n1706) );
  IV U2349 ( .A(n3933), .Z(n3322) );
  XOR U2350 ( .A(in[519]), .B(n3322), .Z(n1780) );
  XOR U2351 ( .A(in[1544]), .B(in[584]), .Z(n1348) );
  XNOR U2352 ( .A(in[904]), .B(in[264]), .Z(n1347) );
  XNOR U2353 ( .A(n1348), .B(n1347), .Z(n1349) );
  XOR U2354 ( .A(in[1224]), .B(n1349), .Z(n1710) );
  XOR U2355 ( .A(n1350), .B(n1710), .Z(n3937) );
  XOR U2356 ( .A(in[520]), .B(n3937), .Z(n1782) );
  XOR U2357 ( .A(in[1545]), .B(in[585]), .Z(n1352) );
  XNOR U2358 ( .A(in[905]), .B(in[265]), .Z(n1351) );
  XNOR U2359 ( .A(n1352), .B(n1351), .Z(n1353) );
  XOR U2360 ( .A(in[1225]), .B(n1353), .Z(n1714) );
  XOR U2361 ( .A(n1354), .B(n1714), .Z(n3944) );
  XOR U2362 ( .A(in[521]), .B(n3944), .Z(n1784) );
  XOR U2363 ( .A(in[1546]), .B(in[586]), .Z(n1356) );
  XNOR U2364 ( .A(in[906]), .B(in[266]), .Z(n1355) );
  XNOR U2365 ( .A(n1356), .B(n1355), .Z(n1357) );
  XOR U2366 ( .A(in[1226]), .B(n1357), .Z(n1718) );
  XOR U2367 ( .A(n1358), .B(n1718), .Z(n3948) );
  XOR U2368 ( .A(in[522]), .B(n3948), .Z(n1786) );
  NOR U2369 ( .A(n1359), .B(n1558), .Z(n1360) );
  XNOR U2370 ( .A(n1786), .B(n1360), .Z(out[1079]) );
  XOR U2371 ( .A(n1362), .B(n1361), .Z(n3986) );
  XOR U2372 ( .A(in[578]), .B(n3986), .Z(n2721) );
  IV U2373 ( .A(n2721), .Z(n2809) );
  IV U2374 ( .A(n1363), .Z(n4123) );
  XOR U2375 ( .A(in[1453]), .B(n4123), .Z(n3260) );
  XNOR U2376 ( .A(in[233]), .B(n2041), .Z(n3262) );
  NANDN U2377 ( .A(n3260), .B(n3262), .Z(n1364) );
  XOR U2378 ( .A(n2809), .B(n1364), .Z(out[107]) );
  XOR U2379 ( .A(in[1547]), .B(in[587]), .Z(n1366) );
  XNOR U2380 ( .A(in[907]), .B(in[267]), .Z(n1365) );
  XNOR U2381 ( .A(n1366), .B(n1365), .Z(n1367) );
  XOR U2382 ( .A(in[1227]), .B(n1367), .Z(n1722) );
  XOR U2383 ( .A(n1368), .B(n1722), .Z(n3952) );
  XOR U2384 ( .A(in[523]), .B(n3952), .Z(n1788) );
  NOR U2385 ( .A(n1369), .B(n1562), .Z(n1370) );
  XNOR U2386 ( .A(n1788), .B(n1370), .Z(out[1080]) );
  XOR U2387 ( .A(in[1548]), .B(in[588]), .Z(n1372) );
  XNOR U2388 ( .A(in[908]), .B(in[268]), .Z(n1371) );
  XNOR U2389 ( .A(n1372), .B(n1371), .Z(n1373) );
  XOR U2390 ( .A(in[1228]), .B(n1373), .Z(n1726) );
  XOR U2391 ( .A(n1374), .B(n1726), .Z(n3956) );
  XOR U2392 ( .A(in[524]), .B(n3956), .Z(n1790) );
  NOR U2393 ( .A(n1375), .B(n1566), .Z(n1376) );
  XNOR U2394 ( .A(n1790), .B(n1376), .Z(out[1081]) );
  XOR U2395 ( .A(in[1549]), .B(in[589]), .Z(n1378) );
  XNOR U2396 ( .A(in[909]), .B(in[269]), .Z(n1377) );
  XNOR U2397 ( .A(n1378), .B(n1377), .Z(n1379) );
  XOR U2398 ( .A(in[1229]), .B(n1379), .Z(n1730) );
  XOR U2399 ( .A(n1380), .B(n1730), .Z(n3960) );
  XOR U2400 ( .A(in[525]), .B(n3960), .Z(n1794) );
  XOR U2401 ( .A(in[1550]), .B(in[590]), .Z(n1382) );
  XNOR U2402 ( .A(in[910]), .B(in[270]), .Z(n1381) );
  XNOR U2403 ( .A(n1382), .B(n1381), .Z(n1383) );
  XNOR U2404 ( .A(in[1230]), .B(n1383), .Z(n1734) );
  XOR U2405 ( .A(n1734), .B(n1384), .Z(n3964) );
  XOR U2406 ( .A(in[526]), .B(n3964), .Z(n1796) );
  XOR U2407 ( .A(in[1551]), .B(in[591]), .Z(n1386) );
  XNOR U2408 ( .A(in[911]), .B(in[271]), .Z(n1385) );
  XNOR U2409 ( .A(n1386), .B(n1385), .Z(n1387) );
  XNOR U2410 ( .A(in[1231]), .B(n1387), .Z(n1738) );
  XOR U2411 ( .A(n1738), .B(n1388), .Z(n3968) );
  XOR U2412 ( .A(in[527]), .B(n3968), .Z(n1798) );
  XOR U2413 ( .A(in[1552]), .B(in[592]), .Z(n1390) );
  XNOR U2414 ( .A(in[912]), .B(in[272]), .Z(n1389) );
  XNOR U2415 ( .A(n1390), .B(n1389), .Z(n1391) );
  XNOR U2416 ( .A(in[1232]), .B(n1391), .Z(n1742) );
  XOR U2417 ( .A(n1742), .B(n1392), .Z(n3972) );
  XOR U2418 ( .A(in[528]), .B(n3972), .Z(n1800) );
  XOR U2419 ( .A(in[1553]), .B(in[593]), .Z(n1394) );
  XNOR U2420 ( .A(in[913]), .B(in[273]), .Z(n1393) );
  XNOR U2421 ( .A(n1394), .B(n1393), .Z(n1395) );
  XNOR U2422 ( .A(in[1233]), .B(n1395), .Z(n1747) );
  XOR U2423 ( .A(n1747), .B(n1396), .Z(n3976) );
  XOR U2424 ( .A(in[529]), .B(n3976), .Z(n1802) );
  XOR U2425 ( .A(in[1554]), .B(in[594]), .Z(n1398) );
  XNOR U2426 ( .A(in[914]), .B(in[274]), .Z(n1397) );
  XNOR U2427 ( .A(n1398), .B(n1397), .Z(n1399) );
  XNOR U2428 ( .A(in[1234]), .B(n1399), .Z(n1751) );
  XOR U2429 ( .A(n1751), .B(n1400), .Z(n3980) );
  XOR U2430 ( .A(in[530]), .B(n3980), .Z(n1804) );
  XNOR U2431 ( .A(in[957]), .B(n3963), .Z(n1807) );
  XNOR U2432 ( .A(in[958]), .B(n3967), .Z(n1810) );
  XNOR U2433 ( .A(n1402), .B(n1401), .Z(n3990) );
  XOR U2434 ( .A(in[579]), .B(n3990), .Z(n2723) );
  IV U2435 ( .A(n2723), .Z(n2811) );
  IV U2436 ( .A(n1403), .Z(n4127) );
  XOR U2437 ( .A(in[1454]), .B(n4127), .Z(n3270) );
  XNOR U2438 ( .A(in[234]), .B(n2043), .Z(n3272) );
  NANDN U2439 ( .A(n3270), .B(n3272), .Z(n1404) );
  XOR U2440 ( .A(n2811), .B(n1404), .Z(out[108]) );
  XNOR U2441 ( .A(in[959]), .B(n3971), .Z(n1813) );
  XNOR U2442 ( .A(in[896]), .B(n3975), .Z(n1816) );
  XNOR U2443 ( .A(in[897]), .B(n3979), .Z(n1821) );
  XNOR U2444 ( .A(in[898]), .B(n3986), .Z(n1824) );
  XNOR U2445 ( .A(in[899]), .B(n3990), .Z(n1826) );
  XOR U2446 ( .A(n1406), .B(n1405), .Z(n2007) );
  XOR U2447 ( .A(in[900]), .B(n2007), .Z(n1827) );
  XOR U2448 ( .A(n1408), .B(n1407), .Z(n2010) );
  XOR U2449 ( .A(in[901]), .B(n2010), .Z(n1829) );
  XOR U2450 ( .A(n1410), .B(n1409), .Z(n2013) );
  XOR U2451 ( .A(in[902]), .B(n2013), .Z(n1831) );
  XOR U2452 ( .A(n1412), .B(n1411), .Z(n2016) );
  XOR U2453 ( .A(in[903]), .B(n2016), .Z(n1833) );
  XOR U2454 ( .A(n1414), .B(n1413), .Z(n2018) );
  XOR U2455 ( .A(in[904]), .B(n2018), .Z(n1835) );
  IV U2456 ( .A(n2007), .Z(n3994) );
  XOR U2457 ( .A(in[580]), .B(n3994), .Z(n2813) );
  IV U2458 ( .A(n1415), .Z(n4131) );
  XOR U2459 ( .A(in[1455]), .B(n4131), .Z(n3304) );
  XNOR U2460 ( .A(in[235]), .B(n4092), .Z(n3306) );
  NANDN U2461 ( .A(n3304), .B(n3306), .Z(n1416) );
  XNOR U2462 ( .A(n2813), .B(n1416), .Z(out[109]) );
  XNOR U2463 ( .A(in[200]), .B(n3937), .Z(n4286) );
  XOR U2464 ( .A(in[1420]), .B(n3198), .Z(n4287) );
  XNOR U2465 ( .A(n4489), .B(in[1043]), .Z(n2881) );
  NANDN U2466 ( .A(n4287), .B(n2881), .Z(n1417) );
  XNOR U2467 ( .A(n4286), .B(n1417), .Z(out[10]) );
  XOR U2468 ( .A(n1419), .B(n1418), .Z(n2020) );
  XOR U2469 ( .A(in[905]), .B(n2020), .Z(n1837) );
  XOR U2470 ( .A(n1421), .B(n1420), .Z(n2023) );
  XOR U2471 ( .A(in[906]), .B(n2023), .Z(n1839) );
  XOR U2472 ( .A(n1422), .B(n227), .Z(n4022) );
  XOR U2473 ( .A(in[907]), .B(n4022), .Z(n1843) );
  XNOR U2474 ( .A(n1424), .B(n1423), .Z(n1704) );
  XOR U2475 ( .A(in[908]), .B(n1704), .Z(n1845) );
  XOR U2476 ( .A(n1426), .B(n1425), .Z(n2027) );
  XOR U2477 ( .A(in[909]), .B(n2027), .Z(n1847) );
  XOR U2478 ( .A(n1428), .B(n1427), .Z(n3118) );
  XOR U2479 ( .A(in[910]), .B(n3118), .Z(n1849) );
  XOR U2480 ( .A(n1430), .B(n1429), .Z(n3120) );
  XOR U2481 ( .A(in[911]), .B(n3120), .Z(n1851) );
  XOR U2482 ( .A(n1432), .B(n1431), .Z(n3122) );
  XOR U2483 ( .A(in[912]), .B(n3122), .Z(n1853) );
  XOR U2484 ( .A(n1434), .B(n1433), .Z(n3124) );
  XOR U2485 ( .A(in[913]), .B(n3124), .Z(n1855) );
  XOR U2486 ( .A(n1436), .B(n1435), .Z(n3126) );
  XOR U2487 ( .A(in[914]), .B(n3126), .Z(n1857) );
  IV U2488 ( .A(n2010), .Z(n3998) );
  XOR U2489 ( .A(in[581]), .B(n3998), .Z(n2815) );
  IV U2490 ( .A(n1437), .Z(n4135) );
  XOR U2491 ( .A(in[1456]), .B(n4135), .Z(n3334) );
  XNOR U2492 ( .A(in[236]), .B(n4096), .Z(n3336) );
  NANDN U2493 ( .A(n3334), .B(n3336), .Z(n1438) );
  XNOR U2494 ( .A(n2815), .B(n1438), .Z(out[110]) );
  XOR U2495 ( .A(n1440), .B(n1439), .Z(n3128) );
  XOR U2496 ( .A(in[915]), .B(n3128), .Z(n1859) );
  XNOR U2497 ( .A(n1442), .B(n1441), .Z(n3130) );
  XOR U2498 ( .A(in[916]), .B(n3130), .Z(n1861) );
  XOR U2499 ( .A(n1444), .B(n1443), .Z(n3132) );
  XOR U2500 ( .A(in[917]), .B(n3132), .Z(n1865) );
  XNOR U2501 ( .A(n1446), .B(n1445), .Z(n3134) );
  XOR U2502 ( .A(in[918]), .B(n3134), .Z(n1867) );
  XNOR U2503 ( .A(n1448), .B(n1447), .Z(n3136) );
  XOR U2504 ( .A(in[919]), .B(n3136), .Z(n1869) );
  XNOR U2505 ( .A(n1450), .B(n1449), .Z(n3142) );
  XOR U2506 ( .A(in[920]), .B(n3142), .Z(n1871) );
  NOR U2507 ( .A(n1451), .B(n1702), .Z(n1452) );
  XNOR U2508 ( .A(n1871), .B(n1452), .Z(out[1115]) );
  XNOR U2509 ( .A(n1454), .B(n1453), .Z(n3144) );
  XOR U2510 ( .A(in[921]), .B(n3144), .Z(n1873) );
  XNOR U2511 ( .A(n1456), .B(n1455), .Z(n3147) );
  XOR U2512 ( .A(in[922]), .B(n3147), .Z(n1875) );
  XNOR U2513 ( .A(n1458), .B(n1457), .Z(n3149) );
  XOR U2514 ( .A(in[923]), .B(n3149), .Z(n1877) );
  NOR U2515 ( .A(n1459), .B(n1716), .Z(n1460) );
  XNOR U2516 ( .A(n1877), .B(n1460), .Z(out[1118]) );
  XNOR U2517 ( .A(n1462), .B(n1461), .Z(n3028) );
  XOR U2518 ( .A(in[924]), .B(n3028), .Z(n1879) );
  NOR U2519 ( .A(n1463), .B(n1720), .Z(n1464) );
  XNOR U2520 ( .A(n1879), .B(n1464), .Z(out[1119]) );
  IV U2521 ( .A(n2013), .Z(n4002) );
  XOR U2522 ( .A(in[582]), .B(n4002), .Z(n2817) );
  IV U2523 ( .A(n1465), .Z(n4139) );
  XOR U2524 ( .A(in[1457]), .B(n4139), .Z(n3362) );
  XNOR U2525 ( .A(in[237]), .B(n4100), .Z(n3364) );
  NANDN U2526 ( .A(n3362), .B(n3364), .Z(n1466) );
  XNOR U2527 ( .A(n2817), .B(n1466), .Z(out[111]) );
  XNOR U2528 ( .A(n1468), .B(n1467), .Z(n3030) );
  XOR U2529 ( .A(in[925]), .B(n3030), .Z(n1881) );
  NOR U2530 ( .A(n1469), .B(n1724), .Z(n1470) );
  XNOR U2531 ( .A(n1881), .B(n1470), .Z(out[1120]) );
  XNOR U2532 ( .A(n1472), .B(n1471), .Z(n3032) );
  XOR U2533 ( .A(in[926]), .B(n3032), .Z(n1883) );
  NOR U2534 ( .A(n1473), .B(n1728), .Z(n1474) );
  XNOR U2535 ( .A(n1883), .B(n1474), .Z(out[1121]) );
  XNOR U2536 ( .A(n1476), .B(n1475), .Z(n3034) );
  XOR U2537 ( .A(in[927]), .B(n3034), .Z(n1887) );
  XNOR U2538 ( .A(n1478), .B(n1477), .Z(n3036) );
  XOR U2539 ( .A(in[928]), .B(n3036), .Z(n1889) );
  NOR U2540 ( .A(n5143), .B(n1736), .Z(n1479) );
  XNOR U2541 ( .A(n1889), .B(n1479), .Z(out[1123]) );
  XOR U2542 ( .A(n1481), .B(n1480), .Z(n3038) );
  XOR U2543 ( .A(in[929]), .B(n3038), .Z(n1891) );
  NOR U2544 ( .A(n5147), .B(n1740), .Z(n1482) );
  XNOR U2545 ( .A(n1891), .B(n1482), .Z(out[1124]) );
  XOR U2546 ( .A(n1484), .B(n1483), .Z(n2168) );
  XOR U2547 ( .A(in[930]), .B(n2168), .Z(n1893) );
  NOR U2548 ( .A(n5151), .B(n1744), .Z(n1485) );
  XNOR U2549 ( .A(n1893), .B(n1485), .Z(out[1125]) );
  XOR U2550 ( .A(n1487), .B(n1486), .Z(n3041) );
  XOR U2551 ( .A(in[931]), .B(n3041), .Z(n1895) );
  NOR U2552 ( .A(n5155), .B(n1749), .Z(n1488) );
  XNOR U2553 ( .A(n1895), .B(n1488), .Z(out[1126]) );
  XOR U2554 ( .A(n1490), .B(n1489), .Z(n3043) );
  XOR U2555 ( .A(in[932]), .B(n3043), .Z(n1897) );
  NOR U2556 ( .A(n5159), .B(n1753), .Z(n1491) );
  XNOR U2557 ( .A(n1897), .B(n1491), .Z(out[1127]) );
  XOR U2558 ( .A(n1493), .B(n1492), .Z(n4138) );
  XOR U2559 ( .A(in[933]), .B(n4138), .Z(n1900) );
  NAND U2560 ( .A(n1494), .B(n1755), .Z(n1495) );
  XNOR U2561 ( .A(n1900), .B(n1495), .Z(out[1128]) );
  XNOR U2562 ( .A(n1497), .B(n1496), .Z(n4142) );
  XOR U2563 ( .A(in[934]), .B(n4142), .Z(n1904) );
  NAND U2564 ( .A(n1498), .B(n1757), .Z(n1499) );
  XNOR U2565 ( .A(n1904), .B(n1499), .Z(out[1129]) );
  IV U2566 ( .A(n2016), .Z(n4006) );
  XOR U2567 ( .A(in[583]), .B(n4006), .Z(n2822) );
  IV U2568 ( .A(n1500), .Z(n4143) );
  XOR U2569 ( .A(in[1458]), .B(n4143), .Z(n3390) );
  XNOR U2570 ( .A(in[238]), .B(n4104), .Z(n3392) );
  NANDN U2571 ( .A(n3390), .B(n3392), .Z(n1501) );
  XNOR U2572 ( .A(n2822), .B(n1501), .Z(out[112]) );
  XOR U2573 ( .A(n1503), .B(n1502), .Z(n4146) );
  XOR U2574 ( .A(in[935]), .B(n4146), .Z(n1908) );
  NAND U2575 ( .A(n1504), .B(n1759), .Z(n1505) );
  XNOR U2576 ( .A(n1908), .B(n1505), .Z(out[1130]) );
  XOR U2577 ( .A(n1507), .B(n1506), .Z(n4150) );
  XOR U2578 ( .A(in[936]), .B(n4150), .Z(n1912) );
  NANDN U2579 ( .A(n1761), .B(n1508), .Z(n1509) );
  XNOR U2580 ( .A(n1912), .B(n1509), .Z(out[1131]) );
  XOR U2581 ( .A(n1511), .B(n1510), .Z(n4154) );
  XOR U2582 ( .A(in[937]), .B(n4154), .Z(n1918) );
  NAND U2583 ( .A(n1512), .B(n1762), .Z(n1513) );
  XNOR U2584 ( .A(n1918), .B(n1513), .Z(out[1132]) );
  XOR U2585 ( .A(n1515), .B(n1514), .Z(n4164) );
  XOR U2586 ( .A(in[938]), .B(n4164), .Z(n1922) );
  NAND U2587 ( .A(n1516), .B(n1764), .Z(n1517) );
  XNOR U2588 ( .A(n1922), .B(n1517), .Z(out[1133]) );
  XOR U2589 ( .A(n1519), .B(n1518), .Z(n4168) );
  XOR U2590 ( .A(in[939]), .B(n4168), .Z(n1926) );
  NAND U2591 ( .A(n1520), .B(n1766), .Z(n1521) );
  XNOR U2592 ( .A(n1926), .B(n1521), .Z(out[1134]) );
  XOR U2593 ( .A(n1523), .B(n1522), .Z(n4172) );
  XOR U2594 ( .A(in[940]), .B(n4172), .Z(n1930) );
  NAND U2595 ( .A(n1524), .B(n1768), .Z(n1525) );
  XNOR U2596 ( .A(n1930), .B(n1525), .Z(out[1135]) );
  XOR U2597 ( .A(n1527), .B(n1526), .Z(n4176) );
  XOR U2598 ( .A(in[941]), .B(n4176), .Z(n1934) );
  NAND U2599 ( .A(n1528), .B(n1772), .Z(n1529) );
  XNOR U2600 ( .A(n1934), .B(n1529), .Z(out[1136]) );
  XOR U2601 ( .A(n1531), .B(n1530), .Z(n3900) );
  XOR U2602 ( .A(in[942]), .B(n3900), .Z(n1938) );
  NAND U2603 ( .A(n1532), .B(n1774), .Z(n1533) );
  XNOR U2604 ( .A(n1938), .B(n1533), .Z(out[1137]) );
  XOR U2605 ( .A(n1535), .B(n1534), .Z(n3904) );
  XOR U2606 ( .A(in[943]), .B(n3904), .Z(n1942) );
  NAND U2607 ( .A(n1536), .B(n1776), .Z(n1537) );
  XNOR U2608 ( .A(n1942), .B(n1537), .Z(out[1138]) );
  XOR U2609 ( .A(n1539), .B(n1538), .Z(n3908) );
  XOR U2610 ( .A(in[944]), .B(n3908), .Z(n1946) );
  NAND U2611 ( .A(n1540), .B(n1778), .Z(n1541) );
  XNOR U2612 ( .A(n1946), .B(n1541), .Z(out[1139]) );
  IV U2613 ( .A(n2018), .Z(n4010) );
  XOR U2614 ( .A(in[584]), .B(n4010), .Z(n2824) );
  IV U2615 ( .A(n1542), .Z(n4147) );
  XOR U2616 ( .A(in[1459]), .B(n4147), .Z(n3425) );
  XNOR U2617 ( .A(in[239]), .B(n4108), .Z(n3427) );
  NANDN U2618 ( .A(n3425), .B(n3427), .Z(n1543) );
  XNOR U2619 ( .A(n2824), .B(n1543), .Z(out[113]) );
  XOR U2620 ( .A(n1545), .B(n1544), .Z(n3912) );
  XOR U2621 ( .A(in[945]), .B(n3912), .Z(n1950) );
  NAND U2622 ( .A(n1546), .B(n1780), .Z(n1547) );
  XNOR U2623 ( .A(n1950), .B(n1547), .Z(out[1140]) );
  XOR U2624 ( .A(n1549), .B(n1548), .Z(n3916) );
  XOR U2625 ( .A(in[946]), .B(n3916), .Z(n1954) );
  NAND U2626 ( .A(n1550), .B(n1782), .Z(n1551) );
  XNOR U2627 ( .A(n1954), .B(n1551), .Z(out[1141]) );
  XNOR U2628 ( .A(n1553), .B(n1552), .Z(n3920) );
  IV U2629 ( .A(n3920), .Z(n2573) );
  XOR U2630 ( .A(in[947]), .B(n2573), .Z(n1960) );
  NAND U2631 ( .A(n1554), .B(n1784), .Z(n1555) );
  XNOR U2632 ( .A(n1960), .B(n1555), .Z(out[1142]) );
  XNOR U2633 ( .A(n1557), .B(n1556), .Z(n3924) );
  IV U2634 ( .A(n3924), .Z(n2615) );
  XOR U2635 ( .A(in[948]), .B(n2615), .Z(n1964) );
  NAND U2636 ( .A(n1558), .B(n1786), .Z(n1559) );
  XNOR U2637 ( .A(n1964), .B(n1559), .Z(out[1143]) );
  XNOR U2638 ( .A(n1561), .B(n1560), .Z(n3928) );
  IV U2639 ( .A(n3928), .Z(n2657) );
  XOR U2640 ( .A(in[949]), .B(n2657), .Z(n1968) );
  NAND U2641 ( .A(n1562), .B(n1788), .Z(n1563) );
  XNOR U2642 ( .A(n1968), .B(n1563), .Z(out[1144]) );
  XOR U2643 ( .A(n1565), .B(n1564), .Z(n3069) );
  XOR U2644 ( .A(in[950]), .B(n3069), .Z(n1972) );
  NAND U2645 ( .A(n1566), .B(n1790), .Z(n1567) );
  XNOR U2646 ( .A(n1972), .B(n1567), .Z(out[1145]) );
  XOR U2647 ( .A(n1569), .B(n1568), .Z(n3071) );
  XOR U2648 ( .A(in[951]), .B(n3071), .Z(n1976) );
  NAND U2649 ( .A(n1570), .B(n1794), .Z(n1571) );
  XNOR U2650 ( .A(n1976), .B(n1571), .Z(out[1146]) );
  XOR U2651 ( .A(n1573), .B(n1572), .Z(n3074) );
  XOR U2652 ( .A(in[952]), .B(n3074), .Z(n1980) );
  NAND U2653 ( .A(n1574), .B(n1796), .Z(n1575) );
  XNOR U2654 ( .A(n1980), .B(n1575), .Z(out[1147]) );
  XNOR U2655 ( .A(n1577), .B(n1576), .Z(n3947) );
  IV U2656 ( .A(n3947), .Z(n2702) );
  XOR U2657 ( .A(in[953]), .B(n2702), .Z(n1984) );
  NAND U2658 ( .A(n1578), .B(n1798), .Z(n1579) );
  XNOR U2659 ( .A(n1984), .B(n1579), .Z(out[1148]) );
  XNOR U2660 ( .A(n1581), .B(n1580), .Z(n3951) );
  IV U2661 ( .A(n3951), .Z(n2704) );
  XOR U2662 ( .A(in[954]), .B(n2704), .Z(n1988) );
  NAND U2663 ( .A(n1582), .B(n1800), .Z(n1583) );
  XNOR U2664 ( .A(n1988), .B(n1583), .Z(out[1149]) );
  IV U2665 ( .A(n2020), .Z(n4014) );
  XOR U2666 ( .A(in[585]), .B(n4014), .Z(n2826) );
  IV U2667 ( .A(n1584), .Z(n4151) );
  XOR U2668 ( .A(in[1460]), .B(n4151), .Z(n3460) );
  XNOR U2669 ( .A(in[240]), .B(n4112), .Z(n3462) );
  NANDN U2670 ( .A(n3460), .B(n3462), .Z(n1585) );
  XNOR U2671 ( .A(n2826), .B(n1585), .Z(out[114]) );
  XOR U2672 ( .A(in[955]), .B(n3955), .Z(n1992) );
  NAND U2673 ( .A(n1586), .B(n1802), .Z(n1587) );
  XNOR U2674 ( .A(n1992), .B(n1587), .Z(out[1150]) );
  XOR U2675 ( .A(in[956]), .B(n3959), .Z(n1996) );
  NANDN U2676 ( .A(n1588), .B(n1804), .Z(n1589) );
  XNOR U2677 ( .A(n1996), .B(n1589), .Z(out[1151]) );
  XOR U2678 ( .A(n1591), .B(n1590), .Z(n4302) );
  XOR U2679 ( .A(in[1004]), .B(n4302), .Z(n1806) );
  NAND U2680 ( .A(n1592), .B(n1807), .Z(n1593) );
  XNOR U2681 ( .A(n1806), .B(n1593), .Z(out[1152]) );
  XOR U2682 ( .A(n1595), .B(n1594), .Z(n4304) );
  XOR U2683 ( .A(in[1005]), .B(n4304), .Z(n1809) );
  NAND U2684 ( .A(n1596), .B(n1810), .Z(n1597) );
  XNOR U2685 ( .A(n1809), .B(n1597), .Z(out[1153]) );
  XOR U2686 ( .A(n1599), .B(n1598), .Z(n4306) );
  XOR U2687 ( .A(in[1006]), .B(n4306), .Z(n1812) );
  NAND U2688 ( .A(n1600), .B(n1813), .Z(n1601) );
  XNOR U2689 ( .A(n1812), .B(n1601), .Z(out[1154]) );
  XOR U2690 ( .A(n1603), .B(n1602), .Z(n4308) );
  XOR U2691 ( .A(in[1007]), .B(n4308), .Z(n1815) );
  NAND U2692 ( .A(n1604), .B(n1816), .Z(n1605) );
  XNOR U2693 ( .A(n1815), .B(n1605), .Z(out[1155]) );
  XOR U2694 ( .A(n1607), .B(n1606), .Z(n4315) );
  XOR U2695 ( .A(in[1008]), .B(n4315), .Z(n1820) );
  NAND U2696 ( .A(n1608), .B(n1821), .Z(n1609) );
  XNOR U2697 ( .A(n1820), .B(n1609), .Z(out[1156]) );
  XOR U2698 ( .A(n1611), .B(n1610), .Z(n4318) );
  XOR U2699 ( .A(in[1009]), .B(n4318), .Z(n1823) );
  NAND U2700 ( .A(n1612), .B(n1824), .Z(n1613) );
  XNOR U2701 ( .A(n1823), .B(n1613), .Z(out[1157]) );
  XOR U2702 ( .A(n1615), .B(n1614), .Z(n4321) );
  XOR U2703 ( .A(in[1010]), .B(n4321), .Z(n5026) );
  NAND U2704 ( .A(n1616), .B(n1826), .Z(n1617) );
  XNOR U2705 ( .A(n5026), .B(n1617), .Z(out[1158]) );
  XOR U2706 ( .A(n1619), .B(n1618), .Z(n4324) );
  XOR U2707 ( .A(in[1011]), .B(n4324), .Z(n5030) );
  NAND U2708 ( .A(n1620), .B(n1827), .Z(n1621) );
  XNOR U2709 ( .A(n5030), .B(n1621), .Z(out[1159]) );
  IV U2710 ( .A(n2023), .Z(n4018) );
  XOR U2711 ( .A(in[586]), .B(n4018), .Z(n2828) );
  XNOR U2712 ( .A(in[1461]), .B(n4155), .Z(n3482) );
  XNOR U2713 ( .A(in[241]), .B(n4120), .Z(n3484) );
  NANDN U2714 ( .A(n3482), .B(n3484), .Z(n1622) );
  XNOR U2715 ( .A(n2828), .B(n1622), .Z(out[115]) );
  XOR U2716 ( .A(n1624), .B(n1623), .Z(n4327) );
  XOR U2717 ( .A(in[1012]), .B(n4327), .Z(n5034) );
  NAND U2718 ( .A(n1625), .B(n1829), .Z(n1626) );
  XNOR U2719 ( .A(n5034), .B(n1626), .Z(out[1160]) );
  XOR U2720 ( .A(n1628), .B(n1627), .Z(n4330) );
  XOR U2721 ( .A(in[1013]), .B(n4330), .Z(n5038) );
  NAND U2722 ( .A(n1629), .B(n1831), .Z(n1630) );
  XNOR U2723 ( .A(n5038), .B(n1630), .Z(out[1161]) );
  XOR U2724 ( .A(n1632), .B(n1631), .Z(n4333) );
  XOR U2725 ( .A(in[1014]), .B(n4333), .Z(n5046) );
  NAND U2726 ( .A(n1633), .B(n1833), .Z(n1634) );
  XNOR U2727 ( .A(n5046), .B(n1634), .Z(out[1162]) );
  XOR U2728 ( .A(n1636), .B(n1635), .Z(n4336) );
  XOR U2729 ( .A(in[1015]), .B(n4336), .Z(n5050) );
  NAND U2730 ( .A(n1637), .B(n1835), .Z(n1638) );
  XNOR U2731 ( .A(n5050), .B(n1638), .Z(out[1163]) );
  XOR U2732 ( .A(n1640), .B(n1639), .Z(n4180) );
  XOR U2733 ( .A(in[1016]), .B(n4180), .Z(n5054) );
  NAND U2734 ( .A(n1641), .B(n1837), .Z(n1642) );
  XNOR U2735 ( .A(n5054), .B(n1642), .Z(out[1164]) );
  XOR U2736 ( .A(n1644), .B(n1643), .Z(n4183) );
  XOR U2737 ( .A(in[1017]), .B(n4183), .Z(n5058) );
  NAND U2738 ( .A(n1645), .B(n1839), .Z(n1646) );
  XNOR U2739 ( .A(n5058), .B(n1646), .Z(out[1165]) );
  XOR U2740 ( .A(n1648), .B(n1647), .Z(n4186) );
  XOR U2741 ( .A(in[1018]), .B(n4186), .Z(n5062) );
  NAND U2742 ( .A(n1649), .B(n1843), .Z(n1650) );
  XNOR U2743 ( .A(n5062), .B(n1650), .Z(out[1166]) );
  XOR U2744 ( .A(n1652), .B(n1651), .Z(n4189) );
  XOR U2745 ( .A(in[1019]), .B(n4189), .Z(n5066) );
  NANDN U2746 ( .A(n1653), .B(n1845), .Z(n1654) );
  XNOR U2747 ( .A(n5066), .B(n1654), .Z(out[1167]) );
  IV U2748 ( .A(n3063), .Z(n4192) );
  XOR U2749 ( .A(in[1020]), .B(n4192), .Z(n5069) );
  NANDN U2750 ( .A(n1657), .B(n1847), .Z(n1658) );
  XOR U2751 ( .A(n5069), .B(n1658), .Z(out[1168]) );
  IV U2752 ( .A(n3065), .Z(n4195) );
  XOR U2753 ( .A(in[1021]), .B(n4195), .Z(n5072) );
  NANDN U2754 ( .A(n1661), .B(n1849), .Z(n1662) );
  XOR U2755 ( .A(n5072), .B(n1662), .Z(out[1169]) );
  XNOR U2756 ( .A(in[587]), .B(n4022), .Z(n2830) );
  XNOR U2757 ( .A(in[1462]), .B(n4165), .Z(n3504) );
  XNOR U2758 ( .A(in[242]), .B(n4124), .Z(n3506) );
  NANDN U2759 ( .A(n3504), .B(n3506), .Z(n1663) );
  XNOR U2760 ( .A(n2830), .B(n1663), .Z(out[116]) );
  IV U2761 ( .A(n3067), .Z(n4200) );
  XOR U2762 ( .A(in[1022]), .B(n4200), .Z(n5075) );
  NANDN U2763 ( .A(n1666), .B(n1851), .Z(n1667) );
  XOR U2764 ( .A(n5075), .B(n1667), .Z(out[1170]) );
  XOR U2765 ( .A(n1669), .B(n1668), .Z(n4201) );
  XOR U2766 ( .A(in[1023]), .B(n4201), .Z(n5079) );
  NAND U2767 ( .A(n1670), .B(n1853), .Z(n1671) );
  XNOR U2768 ( .A(n5079), .B(n1671), .Z(out[1171]) );
  IV U2769 ( .A(n3072), .Z(n4202) );
  XOR U2770 ( .A(in[960]), .B(n4202), .Z(n5086) );
  NAND U2771 ( .A(n1674), .B(n1855), .Z(n1675) );
  XOR U2772 ( .A(n5086), .B(n1675), .Z(out[1172]) );
  IV U2773 ( .A(n3075), .Z(n4203) );
  XOR U2774 ( .A(in[961]), .B(n4203), .Z(n5089) );
  NAND U2775 ( .A(n1678), .B(n1857), .Z(n1679) );
  XOR U2776 ( .A(n5089), .B(n1679), .Z(out[1173]) );
  IV U2777 ( .A(n3077), .Z(n4204) );
  XOR U2778 ( .A(in[962]), .B(n4204), .Z(n5092) );
  NAND U2779 ( .A(n1682), .B(n1859), .Z(n1683) );
  XOR U2780 ( .A(n5092), .B(n1683), .Z(out[1174]) );
  IV U2781 ( .A(n3081), .Z(n4205) );
  XOR U2782 ( .A(in[963]), .B(n4205), .Z(n5095) );
  NAND U2783 ( .A(n1686), .B(n1861), .Z(n1687) );
  XOR U2784 ( .A(n5095), .B(n1687), .Z(out[1175]) );
  IV U2785 ( .A(n3083), .Z(n4206) );
  XOR U2786 ( .A(in[964]), .B(n4206), .Z(n5098) );
  NAND U2787 ( .A(n1690), .B(n1865), .Z(n1691) );
  XOR U2788 ( .A(n5098), .B(n1691), .Z(out[1176]) );
  IV U2789 ( .A(n3085), .Z(n4207) );
  XOR U2790 ( .A(in[965]), .B(n4207), .Z(n5101) );
  NAND U2791 ( .A(n1694), .B(n1867), .Z(n1695) );
  XOR U2792 ( .A(n5101), .B(n1695), .Z(out[1177]) );
  IV U2793 ( .A(n3087), .Z(n4210) );
  XOR U2794 ( .A(in[966]), .B(n4210), .Z(n5104) );
  NAND U2795 ( .A(n1698), .B(n1869), .Z(n1699) );
  XOR U2796 ( .A(n5104), .B(n1699), .Z(out[1178]) );
  IV U2797 ( .A(n3089), .Z(n4213) );
  XOR U2798 ( .A(in[967]), .B(n4213), .Z(n5107) );
  NAND U2799 ( .A(n1702), .B(n1871), .Z(n1703) );
  XOR U2800 ( .A(n5107), .B(n1703), .Z(out[1179]) );
  IV U2801 ( .A(n1704), .Z(n4030) );
  XOR U2802 ( .A(in[588]), .B(n4030), .Z(n2832) );
  XNOR U2803 ( .A(in[1463]), .B(n4169), .Z(n3519) );
  XNOR U2804 ( .A(in[243]), .B(n4128), .Z(n3521) );
  NANDN U2805 ( .A(n3519), .B(n3521), .Z(n1705) );
  XNOR U2806 ( .A(n2832), .B(n1705), .Z(out[117]) );
  XNOR U2807 ( .A(n1707), .B(n1706), .Z(n4218) );
  XOR U2808 ( .A(in[968]), .B(n4218), .Z(n5111) );
  NAND U2809 ( .A(n1708), .B(n1873), .Z(n1709) );
  XNOR U2810 ( .A(n5111), .B(n1709), .Z(out[1180]) );
  IV U2811 ( .A(n3092), .Z(n4221) );
  XOR U2812 ( .A(in[969]), .B(n4221), .Z(n5114) );
  NAND U2813 ( .A(n1712), .B(n1875), .Z(n1713) );
  XOR U2814 ( .A(n5114), .B(n1713), .Z(out[1181]) );
  IV U2815 ( .A(n3094), .Z(n4224) );
  XOR U2816 ( .A(in[970]), .B(n4224), .Z(n5121) );
  NAND U2817 ( .A(n1716), .B(n1877), .Z(n1717) );
  XOR U2818 ( .A(n5121), .B(n1717), .Z(out[1182]) );
  XOR U2819 ( .A(in[971]), .B(n3096), .Z(n5125) );
  NAND U2820 ( .A(n1720), .B(n1879), .Z(n1721) );
  XNOR U2821 ( .A(n5125), .B(n1721), .Z(out[1183]) );
  XOR U2822 ( .A(in[972]), .B(n3098), .Z(n5129) );
  NAND U2823 ( .A(n1724), .B(n1881), .Z(n1725) );
  XNOR U2824 ( .A(n5129), .B(n1725), .Z(out[1184]) );
  XOR U2825 ( .A(in[973]), .B(n3102), .Z(n5133) );
  NAND U2826 ( .A(n1728), .B(n1883), .Z(n1729) );
  XNOR U2827 ( .A(n5133), .B(n1729), .Z(out[1185]) );
  XOR U2828 ( .A(in[974]), .B(n3104), .Z(n5137) );
  NAND U2829 ( .A(n1732), .B(n1887), .Z(n1733) );
  XNOR U2830 ( .A(n5137), .B(n1733), .Z(out[1186]) );
  XOR U2831 ( .A(n1735), .B(n1734), .Z(n4237) );
  XOR U2832 ( .A(in[975]), .B(n4237), .Z(n5141) );
  NAND U2833 ( .A(n1736), .B(n1889), .Z(n1737) );
  XNOR U2834 ( .A(n5141), .B(n1737), .Z(out[1187]) );
  XOR U2835 ( .A(n1739), .B(n1738), .Z(n4240) );
  XOR U2836 ( .A(in[976]), .B(n4240), .Z(n5145) );
  NAND U2837 ( .A(n1740), .B(n1891), .Z(n1741) );
  XNOR U2838 ( .A(n5145), .B(n1741), .Z(out[1188]) );
  XOR U2839 ( .A(n1743), .B(n1742), .Z(n4241) );
  XOR U2840 ( .A(in[977]), .B(n4241), .Z(n5149) );
  NAND U2841 ( .A(n1744), .B(n1893), .Z(n1745) );
  XNOR U2842 ( .A(n5149), .B(n1745), .Z(out[1189]) );
  IV U2843 ( .A(n2027), .Z(n4034) );
  XOR U2844 ( .A(in[589]), .B(n4034), .Z(n2834) );
  XNOR U2845 ( .A(in[1464]), .B(n4173), .Z(n3547) );
  XNOR U2846 ( .A(in[244]), .B(n4132), .Z(n3549) );
  NANDN U2847 ( .A(n3547), .B(n3549), .Z(n1746) );
  XNOR U2848 ( .A(n2834), .B(n1746), .Z(out[118]) );
  XOR U2849 ( .A(n1748), .B(n1747), .Z(n4246) );
  XOR U2850 ( .A(in[978]), .B(n4246), .Z(n5152) );
  NAND U2851 ( .A(n1749), .B(n1895), .Z(n1750) );
  XNOR U2852 ( .A(n5152), .B(n1750), .Z(out[1190]) );
  XOR U2853 ( .A(n1752), .B(n1751), .Z(n4249) );
  XOR U2854 ( .A(in[979]), .B(n4249), .Z(n5157) );
  NAND U2855 ( .A(n1753), .B(n1897), .Z(n1754) );
  XNOR U2856 ( .A(n5157), .B(n1754), .Z(out[1191]) );
  OR U2857 ( .A(n1900), .B(n1755), .Z(n1756) );
  XNOR U2858 ( .A(n1899), .B(n1756), .Z(out[1192]) );
  OR U2859 ( .A(n1904), .B(n1757), .Z(n1758) );
  XNOR U2860 ( .A(n1903), .B(n1758), .Z(out[1193]) );
  OR U2861 ( .A(n1908), .B(n1759), .Z(n1760) );
  XNOR U2862 ( .A(n1907), .B(n1760), .Z(out[1194]) );
  OR U2863 ( .A(n1918), .B(n1762), .Z(n1763) );
  XNOR U2864 ( .A(n1917), .B(n1763), .Z(out[1196]) );
  OR U2865 ( .A(n1922), .B(n1764), .Z(n1765) );
  XNOR U2866 ( .A(n1921), .B(n1765), .Z(out[1197]) );
  OR U2867 ( .A(n1926), .B(n1766), .Z(n1767) );
  XNOR U2868 ( .A(n1925), .B(n1767), .Z(out[1198]) );
  OR U2869 ( .A(n1930), .B(n1768), .Z(n1769) );
  XNOR U2870 ( .A(n1929), .B(n1769), .Z(out[1199]) );
  IV U2871 ( .A(n3118), .Z(n4038) );
  XOR U2872 ( .A(in[590]), .B(n4038), .Z(n2836) );
  XNOR U2873 ( .A(in[1465]), .B(n4177), .Z(n3577) );
  XNOR U2874 ( .A(in[245]), .B(n4136), .Z(n3579) );
  NANDN U2875 ( .A(n3577), .B(n3579), .Z(n1770) );
  XNOR U2876 ( .A(n2836), .B(n1770), .Z(out[119]) );
  XNOR U2877 ( .A(in[201]), .B(n3944), .Z(n4311) );
  XOR U2878 ( .A(in[1421]), .B(n3200), .Z(n4312) );
  XNOR U2879 ( .A(in[1044]), .B(n4492), .Z(n2885) );
  NANDN U2880 ( .A(n4312), .B(n2885), .Z(n1771) );
  XNOR U2881 ( .A(n4311), .B(n1771), .Z(out[11]) );
  OR U2882 ( .A(n1934), .B(n1772), .Z(n1773) );
  XNOR U2883 ( .A(n1933), .B(n1773), .Z(out[1200]) );
  OR U2884 ( .A(n1938), .B(n1774), .Z(n1775) );
  XNOR U2885 ( .A(n1937), .B(n1775), .Z(out[1201]) );
  OR U2886 ( .A(n1942), .B(n1776), .Z(n1777) );
  XNOR U2887 ( .A(n1941), .B(n1777), .Z(out[1202]) );
  OR U2888 ( .A(n1946), .B(n1778), .Z(n1779) );
  XNOR U2889 ( .A(n1945), .B(n1779), .Z(out[1203]) );
  OR U2890 ( .A(n1950), .B(n1780), .Z(n1781) );
  XNOR U2891 ( .A(n1949), .B(n1781), .Z(out[1204]) );
  OR U2892 ( .A(n1954), .B(n1782), .Z(n1783) );
  XNOR U2893 ( .A(n1953), .B(n1783), .Z(out[1205]) );
  OR U2894 ( .A(n1960), .B(n1784), .Z(n1785) );
  XNOR U2895 ( .A(n1959), .B(n1785), .Z(out[1206]) );
  OR U2896 ( .A(n1964), .B(n1786), .Z(n1787) );
  XNOR U2897 ( .A(n1963), .B(n1787), .Z(out[1207]) );
  OR U2898 ( .A(n1968), .B(n1788), .Z(n1789) );
  XNOR U2899 ( .A(n1967), .B(n1789), .Z(out[1208]) );
  OR U2900 ( .A(n1972), .B(n1790), .Z(n1791) );
  XNOR U2901 ( .A(n1971), .B(n1791), .Z(out[1209]) );
  IV U2902 ( .A(n3120), .Z(n4042) );
  XOR U2903 ( .A(in[591]), .B(n4042), .Z(n2838) );
  IV U2904 ( .A(n1792), .Z(n3901) );
  XOR U2905 ( .A(in[1466]), .B(n3901), .Z(n3601) );
  XNOR U2906 ( .A(in[246]), .B(n4140), .Z(n3603) );
  NANDN U2907 ( .A(n3601), .B(n3603), .Z(n1793) );
  XNOR U2908 ( .A(n2838), .B(n1793), .Z(out[120]) );
  OR U2909 ( .A(n1976), .B(n1794), .Z(n1795) );
  XNOR U2910 ( .A(n1975), .B(n1795), .Z(out[1210]) );
  OR U2911 ( .A(n1980), .B(n1796), .Z(n1797) );
  XNOR U2912 ( .A(n1979), .B(n1797), .Z(out[1211]) );
  OR U2913 ( .A(n1984), .B(n1798), .Z(n1799) );
  XNOR U2914 ( .A(n1983), .B(n1799), .Z(out[1212]) );
  OR U2915 ( .A(n1988), .B(n1800), .Z(n1801) );
  XNOR U2916 ( .A(n1987), .B(n1801), .Z(out[1213]) );
  OR U2917 ( .A(n1992), .B(n1802), .Z(n1803) );
  XNOR U2918 ( .A(n1991), .B(n1803), .Z(out[1214]) );
  OR U2919 ( .A(n1996), .B(n1804), .Z(n1805) );
  XNOR U2920 ( .A(n1995), .B(n1805), .Z(out[1215]) );
  IV U2921 ( .A(n1806), .Z(n5001) );
  NANDN U2922 ( .A(n1807), .B(n5001), .Z(n1808) );
  XOR U2923 ( .A(n5002), .B(n1808), .Z(out[1216]) );
  IV U2924 ( .A(n1809), .Z(n5005) );
  NANDN U2925 ( .A(n1810), .B(n5005), .Z(n1811) );
  XOR U2926 ( .A(n5006), .B(n1811), .Z(out[1217]) );
  IV U2927 ( .A(n1812), .Z(n5009) );
  NANDN U2928 ( .A(n1813), .B(n5009), .Z(n1814) );
  XOR U2929 ( .A(n5010), .B(n1814), .Z(out[1218]) );
  IV U2930 ( .A(n1815), .Z(n5013) );
  NANDN U2931 ( .A(n1816), .B(n5013), .Z(n1817) );
  XOR U2932 ( .A(n5014), .B(n1817), .Z(out[1219]) );
  IV U2933 ( .A(n3122), .Z(n4046) );
  XOR U2934 ( .A(in[592]), .B(n4046), .Z(n2840) );
  IV U2935 ( .A(n1818), .Z(n3905) );
  XOR U2936 ( .A(in[1467]), .B(n3905), .Z(n3631) );
  XNOR U2937 ( .A(in[247]), .B(n4144), .Z(n3633) );
  NANDN U2938 ( .A(n3631), .B(n3633), .Z(n1819) );
  XNOR U2939 ( .A(n2840), .B(n1819), .Z(out[121]) );
  IV U2940 ( .A(n1820), .Z(n5017) );
  NANDN U2941 ( .A(n1821), .B(n5017), .Z(n1822) );
  XOR U2942 ( .A(n5018), .B(n1822), .Z(out[1220]) );
  IV U2943 ( .A(n1823), .Z(n5021) );
  NANDN U2944 ( .A(n1824), .B(n5021), .Z(n1825) );
  XOR U2945 ( .A(n5022), .B(n1825), .Z(out[1221]) );
  OR U2946 ( .A(n5030), .B(n1827), .Z(n1828) );
  XNOR U2947 ( .A(n5029), .B(n1828), .Z(out[1223]) );
  OR U2948 ( .A(n5034), .B(n1829), .Z(n1830) );
  XNOR U2949 ( .A(n5033), .B(n1830), .Z(out[1224]) );
  OR U2950 ( .A(n5038), .B(n1831), .Z(n1832) );
  XNOR U2951 ( .A(n5037), .B(n1832), .Z(out[1225]) );
  OR U2952 ( .A(n5046), .B(n1833), .Z(n1834) );
  XNOR U2953 ( .A(n5045), .B(n1834), .Z(out[1226]) );
  OR U2954 ( .A(n5050), .B(n1835), .Z(n1836) );
  XNOR U2955 ( .A(n5049), .B(n1836), .Z(out[1227]) );
  OR U2956 ( .A(n5054), .B(n1837), .Z(n1838) );
  XNOR U2957 ( .A(n5053), .B(n1838), .Z(out[1228]) );
  OR U2958 ( .A(n5058), .B(n1839), .Z(n1840) );
  XNOR U2959 ( .A(n5057), .B(n1840), .Z(out[1229]) );
  IV U2960 ( .A(n3124), .Z(n4050) );
  XOR U2961 ( .A(in[593]), .B(n4050), .Z(n2845) );
  IV U2962 ( .A(n1841), .Z(n3909) );
  XOR U2963 ( .A(in[1468]), .B(n3909), .Z(n3675) );
  XNOR U2964 ( .A(in[248]), .B(n4148), .Z(n3677) );
  NANDN U2965 ( .A(n3675), .B(n3677), .Z(n1842) );
  XNOR U2966 ( .A(n2845), .B(n1842), .Z(out[122]) );
  OR U2967 ( .A(n5062), .B(n1843), .Z(n1844) );
  XNOR U2968 ( .A(n5061), .B(n1844), .Z(out[1230]) );
  OR U2969 ( .A(n5066), .B(n1845), .Z(n1846) );
  XNOR U2970 ( .A(n5065), .B(n1846), .Z(out[1231]) );
  NANDN U2971 ( .A(n1847), .B(n5069), .Z(n1848) );
  XNOR U2972 ( .A(n5070), .B(n1848), .Z(out[1232]) );
  NANDN U2973 ( .A(n1849), .B(n5072), .Z(n1850) );
  XNOR U2974 ( .A(n5073), .B(n1850), .Z(out[1233]) );
  NANDN U2975 ( .A(n1851), .B(n5075), .Z(n1852) );
  XNOR U2976 ( .A(n5076), .B(n1852), .Z(out[1234]) );
  OR U2977 ( .A(n5079), .B(n1853), .Z(n1854) );
  XNOR U2978 ( .A(n5078), .B(n1854), .Z(out[1235]) );
  NANDN U2979 ( .A(n1855), .B(n5086), .Z(n1856) );
  XNOR U2980 ( .A(n5087), .B(n1856), .Z(out[1236]) );
  NANDN U2981 ( .A(n1857), .B(n5089), .Z(n1858) );
  XNOR U2982 ( .A(n5090), .B(n1858), .Z(out[1237]) );
  NANDN U2983 ( .A(n1859), .B(n5092), .Z(n1860) );
  XNOR U2984 ( .A(n5093), .B(n1860), .Z(out[1238]) );
  NANDN U2985 ( .A(n1861), .B(n5095), .Z(n1862) );
  XNOR U2986 ( .A(n5096), .B(n1862), .Z(out[1239]) );
  IV U2987 ( .A(n3126), .Z(n4054) );
  XOR U2988 ( .A(in[594]), .B(n4054), .Z(n2847) );
  IV U2989 ( .A(n1863), .Z(n3913) );
  XOR U2990 ( .A(in[1469]), .B(n3913), .Z(n3719) );
  XNOR U2991 ( .A(in[249]), .B(n4152), .Z(n3721) );
  NANDN U2992 ( .A(n3719), .B(n3721), .Z(n1864) );
  XNOR U2993 ( .A(n2847), .B(n1864), .Z(out[123]) );
  NANDN U2994 ( .A(n1865), .B(n5098), .Z(n1866) );
  XNOR U2995 ( .A(n5099), .B(n1866), .Z(out[1240]) );
  NANDN U2996 ( .A(n1867), .B(n5101), .Z(n1868) );
  XNOR U2997 ( .A(n5102), .B(n1868), .Z(out[1241]) );
  NANDN U2998 ( .A(n1869), .B(n5104), .Z(n1870) );
  XNOR U2999 ( .A(n5105), .B(n1870), .Z(out[1242]) );
  NANDN U3000 ( .A(n1871), .B(n5107), .Z(n1872) );
  XNOR U3001 ( .A(n5108), .B(n1872), .Z(out[1243]) );
  OR U3002 ( .A(n5111), .B(n1873), .Z(n1874) );
  XNOR U3003 ( .A(n5110), .B(n1874), .Z(out[1244]) );
  NANDN U3004 ( .A(n1875), .B(n5114), .Z(n1876) );
  XNOR U3005 ( .A(n5115), .B(n1876), .Z(out[1245]) );
  NANDN U3006 ( .A(n1877), .B(n5121), .Z(n1878) );
  XNOR U3007 ( .A(n5122), .B(n1878), .Z(out[1246]) );
  OR U3008 ( .A(n5125), .B(n1879), .Z(n1880) );
  XNOR U3009 ( .A(n5124), .B(n1880), .Z(out[1247]) );
  OR U3010 ( .A(n5129), .B(n1881), .Z(n1882) );
  XNOR U3011 ( .A(n5128), .B(n1882), .Z(out[1248]) );
  OR U3012 ( .A(n5133), .B(n1883), .Z(n1884) );
  XNOR U3013 ( .A(n5132), .B(n1884), .Z(out[1249]) );
  IV U3014 ( .A(n3128), .Z(n4058) );
  XOR U3015 ( .A(in[595]), .B(n4058), .Z(n2849) );
  IV U3016 ( .A(n1885), .Z(n3917) );
  XOR U3017 ( .A(in[1470]), .B(n3917), .Z(n3765) );
  XNOR U3018 ( .A(in[250]), .B(n4156), .Z(n3767) );
  NANDN U3019 ( .A(n3765), .B(n3767), .Z(n1886) );
  XNOR U3020 ( .A(n2849), .B(n1886), .Z(out[124]) );
  OR U3021 ( .A(n5137), .B(n1887), .Z(n1888) );
  XNOR U3022 ( .A(n5136), .B(n1888), .Z(out[1250]) );
  OR U3023 ( .A(n5141), .B(n1889), .Z(n1890) );
  XNOR U3024 ( .A(n5140), .B(n1890), .Z(out[1251]) );
  OR U3025 ( .A(n5145), .B(n1891), .Z(n1892) );
  XNOR U3026 ( .A(n5144), .B(n1892), .Z(out[1252]) );
  OR U3027 ( .A(n5149), .B(n1893), .Z(n1894) );
  XNOR U3028 ( .A(n5148), .B(n1894), .Z(out[1253]) );
  OR U3029 ( .A(n5152), .B(n1895), .Z(n1896) );
  XOR U3030 ( .A(n5153), .B(n1896), .Z(out[1254]) );
  OR U3031 ( .A(n5157), .B(n1897), .Z(n1898) );
  XNOR U3032 ( .A(n5156), .B(n1898), .Z(out[1255]) );
  ANDN U3033 ( .B(n1900), .A(n1899), .Z(n1901) );
  XOR U3034 ( .A(n1902), .B(n1901), .Z(out[1256]) );
  ANDN U3035 ( .B(n1904), .A(n1903), .Z(n1905) );
  XOR U3036 ( .A(n1906), .B(n1905), .Z(out[1257]) );
  ANDN U3037 ( .B(n1908), .A(n1907), .Z(n1909) );
  XOR U3038 ( .A(n1910), .B(n1909), .Z(out[1258]) );
  ANDN U3039 ( .B(n1912), .A(n1911), .Z(n1913) );
  XOR U3040 ( .A(n1914), .B(n1913), .Z(out[1259]) );
  IV U3041 ( .A(n3130), .Z(n4062) );
  XOR U3042 ( .A(in[596]), .B(n4062), .Z(n2851) );
  IV U3043 ( .A(n1915), .Z(n3921) );
  XOR U3044 ( .A(in[1471]), .B(n3921), .Z(n3809) );
  IV U3045 ( .A(n4166), .Z(n3282) );
  XOR U3046 ( .A(in[251]), .B(n3282), .Z(n3811) );
  OR U3047 ( .A(n3809), .B(n3811), .Z(n1916) );
  XNOR U3048 ( .A(n2851), .B(n1916), .Z(out[125]) );
  ANDN U3049 ( .B(n1918), .A(n1917), .Z(n1919) );
  XOR U3050 ( .A(n1920), .B(n1919), .Z(out[1260]) );
  ANDN U3051 ( .B(n1922), .A(n1921), .Z(n1923) );
  XOR U3052 ( .A(n1924), .B(n1923), .Z(out[1261]) );
  ANDN U3053 ( .B(n1926), .A(n1925), .Z(n1927) );
  XOR U3054 ( .A(n1928), .B(n1927), .Z(out[1262]) );
  ANDN U3055 ( .B(n1930), .A(n1929), .Z(n1931) );
  XOR U3056 ( .A(n1932), .B(n1931), .Z(out[1263]) );
  ANDN U3057 ( .B(n1934), .A(n1933), .Z(n1935) );
  XOR U3058 ( .A(n1936), .B(n1935), .Z(out[1264]) );
  ANDN U3059 ( .B(n1938), .A(n1937), .Z(n1939) );
  XOR U3060 ( .A(n1940), .B(n1939), .Z(out[1265]) );
  ANDN U3061 ( .B(n1942), .A(n1941), .Z(n1943) );
  XOR U3062 ( .A(n1944), .B(n1943), .Z(out[1266]) );
  ANDN U3063 ( .B(n1946), .A(n1945), .Z(n1947) );
  XOR U3064 ( .A(n1948), .B(n1947), .Z(out[1267]) );
  ANDN U3065 ( .B(n1950), .A(n1949), .Z(n1951) );
  XOR U3066 ( .A(n1952), .B(n1951), .Z(out[1268]) );
  ANDN U3067 ( .B(n1954), .A(n1953), .Z(n1955) );
  XOR U3068 ( .A(n1956), .B(n1955), .Z(out[1269]) );
  IV U3069 ( .A(n3132), .Z(n4066) );
  XOR U3070 ( .A(in[597]), .B(n4066), .Z(n2853) );
  IV U3071 ( .A(n1957), .Z(n3925) );
  XOR U3072 ( .A(in[1408]), .B(n3925), .Z(n3853) );
  IV U3073 ( .A(n4170), .Z(n3285) );
  XOR U3074 ( .A(in[252]), .B(n3285), .Z(n3855) );
  OR U3075 ( .A(n3853), .B(n3855), .Z(n1958) );
  XNOR U3076 ( .A(n2853), .B(n1958), .Z(out[126]) );
  ANDN U3077 ( .B(n1960), .A(n1959), .Z(n1961) );
  XOR U3078 ( .A(n1962), .B(n1961), .Z(out[1270]) );
  ANDN U3079 ( .B(n1964), .A(n1963), .Z(n1965) );
  XOR U3080 ( .A(n1966), .B(n1965), .Z(out[1271]) );
  ANDN U3081 ( .B(n1968), .A(n1967), .Z(n1969) );
  XOR U3082 ( .A(n1970), .B(n1969), .Z(out[1272]) );
  ANDN U3083 ( .B(n1972), .A(n1971), .Z(n1973) );
  XOR U3084 ( .A(n1974), .B(n1973), .Z(out[1273]) );
  ANDN U3085 ( .B(n1976), .A(n1975), .Z(n1977) );
  XOR U3086 ( .A(n1978), .B(n1977), .Z(out[1274]) );
  ANDN U3087 ( .B(n1980), .A(n1979), .Z(n1981) );
  XOR U3088 ( .A(n1982), .B(n1981), .Z(out[1275]) );
  ANDN U3089 ( .B(n1984), .A(n1983), .Z(n1985) );
  XOR U3090 ( .A(n1986), .B(n1985), .Z(out[1276]) );
  ANDN U3091 ( .B(n1988), .A(n1987), .Z(n1989) );
  XOR U3092 ( .A(n1990), .B(n1989), .Z(out[1277]) );
  ANDN U3093 ( .B(n1992), .A(n1991), .Z(n1993) );
  XOR U3094 ( .A(n1994), .B(n1993), .Z(out[1278]) );
  ANDN U3095 ( .B(n1996), .A(n1995), .Z(n1997) );
  XOR U3096 ( .A(n1998), .B(n1997), .Z(out[1279]) );
  IV U3097 ( .A(n3134), .Z(n4074) );
  XOR U3098 ( .A(in[598]), .B(n4074), .Z(n2855) );
  IV U3099 ( .A(n1999), .Z(n3929) );
  XOR U3100 ( .A(in[1409]), .B(n3929), .Z(n3897) );
  IV U3101 ( .A(n4174), .Z(n3288) );
  XOR U3102 ( .A(in[253]), .B(n3288), .Z(n3899) );
  OR U3103 ( .A(n3897), .B(n3899), .Z(n2000) );
  XNOR U3104 ( .A(n2855), .B(n2000), .Z(out[127]) );
  XOR U3105 ( .A(in[50]), .B(n4321), .Z(n2181) );
  XNOR U3106 ( .A(in[1172]), .B(n3991), .Z(n2438) );
  XNOR U3107 ( .A(in[1536]), .B(n3975), .Z(n2439) );
  NANDN U3108 ( .A(n2438), .B(n2439), .Z(n2001) );
  XNOR U3109 ( .A(n2181), .B(n2001), .Z(out[1280]) );
  XOR U3110 ( .A(in[51]), .B(n4324), .Z(n2183) );
  XNOR U3111 ( .A(in[1173]), .B(n3995), .Z(n2441) );
  XNOR U3112 ( .A(in[1537]), .B(n3979), .Z(n2442) );
  NANDN U3113 ( .A(n2441), .B(n2442), .Z(n2002) );
  XNOR U3114 ( .A(n2183), .B(n2002), .Z(out[1281]) );
  XOR U3115 ( .A(in[52]), .B(n4327), .Z(n2186) );
  IV U3116 ( .A(n2003), .Z(n3999) );
  XOR U3117 ( .A(in[1174]), .B(n3999), .Z(n2444) );
  XNOR U3118 ( .A(in[1538]), .B(n3986), .Z(n2092) );
  IV U3119 ( .A(n2092), .Z(n2446) );
  OR U3120 ( .A(n2444), .B(n2446), .Z(n2004) );
  XNOR U3121 ( .A(n2186), .B(n2004), .Z(out[1282]) );
  XOR U3122 ( .A(in[53]), .B(n4330), .Z(n2188) );
  XNOR U3123 ( .A(in[1175]), .B(n4003), .Z(n2448) );
  XNOR U3124 ( .A(in[1539]), .B(n3990), .Z(n2449) );
  NANDN U3125 ( .A(n2448), .B(n2449), .Z(n2005) );
  XNOR U3126 ( .A(n2188), .B(n2005), .Z(out[1283]) );
  XOR U3127 ( .A(in[54]), .B(n4333), .Z(n2190) );
  IV U3128 ( .A(n2006), .Z(n4007) );
  XOR U3129 ( .A(in[1176]), .B(n4007), .Z(n2454) );
  XOR U3130 ( .A(in[1540]), .B(n2007), .Z(n2095) );
  IV U3131 ( .A(n2095), .Z(n2456) );
  OR U3132 ( .A(n2454), .B(n2456), .Z(n2008) );
  XNOR U3133 ( .A(n2190), .B(n2008), .Z(out[1284]) );
  XOR U3134 ( .A(in[55]), .B(n4336), .Z(n2192) );
  IV U3135 ( .A(n2009), .Z(n4011) );
  XOR U3136 ( .A(in[1177]), .B(n4011), .Z(n2458) );
  XOR U3137 ( .A(in[1541]), .B(n2010), .Z(n2097) );
  IV U3138 ( .A(n2097), .Z(n2460) );
  OR U3139 ( .A(n2458), .B(n2460), .Z(n2011) );
  XNOR U3140 ( .A(n2192), .B(n2011), .Z(out[1285]) );
  XOR U3141 ( .A(in[56]), .B(n4180), .Z(n2194) );
  IV U3142 ( .A(n2012), .Z(n4015) );
  XOR U3143 ( .A(in[1178]), .B(n4015), .Z(n2462) );
  XOR U3144 ( .A(in[1542]), .B(n2013), .Z(n2100) );
  IV U3145 ( .A(n2100), .Z(n2464) );
  OR U3146 ( .A(n2462), .B(n2464), .Z(n2014) );
  XNOR U3147 ( .A(n2194), .B(n2014), .Z(out[1286]) );
  XOR U3148 ( .A(in[57]), .B(n4183), .Z(n2196) );
  IV U3149 ( .A(n2015), .Z(n4019) );
  XOR U3150 ( .A(in[1179]), .B(n4019), .Z(n2466) );
  XOR U3151 ( .A(in[1543]), .B(n2016), .Z(n2102) );
  IV U3152 ( .A(n2102), .Z(n2468) );
  OR U3153 ( .A(n2466), .B(n2468), .Z(n2017) );
  XNOR U3154 ( .A(n2196), .B(n2017), .Z(out[1287]) );
  XOR U3155 ( .A(in[58]), .B(n4186), .Z(n2198) );
  XNOR U3156 ( .A(in[1180]), .B(n4023), .Z(n2471) );
  XOR U3157 ( .A(in[1544]), .B(n2018), .Z(n2469) );
  NANDN U3158 ( .A(n2471), .B(n2469), .Z(n2019) );
  XNOR U3159 ( .A(n2198), .B(n2019), .Z(out[1288]) );
  XOR U3160 ( .A(in[59]), .B(n4189), .Z(n2200) );
  XNOR U3161 ( .A(in[1181]), .B(n4031), .Z(n2474) );
  XOR U3162 ( .A(in[1545]), .B(n2020), .Z(n2472) );
  NANDN U3163 ( .A(n2474), .B(n2472), .Z(n2021) );
  XNOR U3164 ( .A(n2200), .B(n2021), .Z(out[1289]) );
  XOR U3165 ( .A(in[665]), .B(n4259), .Z(n2857) );
  IV U3166 ( .A(n3136), .Z(n4078) );
  XOR U3167 ( .A(in[599]), .B(n4078), .Z(n3942) );
  OR U3168 ( .A(n3942), .B(n3940), .Z(n2022) );
  XNOR U3169 ( .A(n2857), .B(n2022), .Z(out[128]) );
  XOR U3170 ( .A(in[60]), .B(n3063), .Z(n2202) );
  XNOR U3171 ( .A(in[1182]), .B(n4035), .Z(n2477) );
  XOR U3172 ( .A(in[1546]), .B(n2023), .Z(n2475) );
  NANDN U3173 ( .A(n2477), .B(n2475), .Z(n2024) );
  XNOR U3174 ( .A(n2202), .B(n2024), .Z(out[1290]) );
  XOR U3175 ( .A(in[61]), .B(n3065), .Z(n2204) );
  XNOR U3176 ( .A(in[1183]), .B(n4039), .Z(n2479) );
  XOR U3177 ( .A(in[1547]), .B(n4022), .Z(n2481) );
  NANDN U3178 ( .A(n2479), .B(n2481), .Z(n2025) );
  XNOR U3179 ( .A(n2204), .B(n2025), .Z(out[1291]) );
  XOR U3180 ( .A(in[62]), .B(n3067), .Z(n2207) );
  XNOR U3181 ( .A(in[1184]), .B(n4043), .Z(n2483) );
  XNOR U3182 ( .A(in[1548]), .B(n4030), .Z(n2485) );
  NANDN U3183 ( .A(n2483), .B(n2485), .Z(n2026) );
  XNOR U3184 ( .A(n2207), .B(n2026), .Z(out[1292]) );
  XOR U3185 ( .A(in[63]), .B(n4201), .Z(n2209) );
  XNOR U3186 ( .A(in[1185]), .B(n4047), .Z(n2488) );
  XOR U3187 ( .A(in[1549]), .B(n2027), .Z(n2486) );
  NANDN U3188 ( .A(n2488), .B(n2486), .Z(n2028) );
  XNOR U3189 ( .A(n2209), .B(n2028), .Z(out[1293]) );
  XOR U3190 ( .A(in[0]), .B(n3072), .Z(n2211) );
  XOR U3191 ( .A(in[1550]), .B(n3118), .Z(n2110) );
  IV U3192 ( .A(n2110), .Z(n2493) );
  XNOR U3193 ( .A(n3397), .B(in[1186]), .Z(n2490) );
  NANDN U3194 ( .A(n2493), .B(n2490), .Z(n2029) );
  XNOR U3195 ( .A(n2211), .B(n2029), .Z(out[1294]) );
  XOR U3196 ( .A(in[1]), .B(n3075), .Z(n2213) );
  XOR U3197 ( .A(in[1551]), .B(n3120), .Z(n2113) );
  IV U3198 ( .A(n2113), .Z(n2496) );
  XNOR U3199 ( .A(n3400), .B(in[1187]), .Z(n2494) );
  NANDN U3200 ( .A(n2496), .B(n2494), .Z(n2030) );
  XNOR U3201 ( .A(n2213), .B(n2030), .Z(out[1295]) );
  XOR U3202 ( .A(in[2]), .B(n3077), .Z(n2216) );
  XOR U3203 ( .A(in[1552]), .B(n3122), .Z(n2117) );
  IV U3204 ( .A(n2117), .Z(n2502) );
  XNOR U3205 ( .A(n3404), .B(in[1188]), .Z(n2499) );
  NANDN U3206 ( .A(n2502), .B(n2499), .Z(n2031) );
  XNOR U3207 ( .A(n2216), .B(n2031), .Z(out[1296]) );
  XOR U3208 ( .A(in[3]), .B(n3081), .Z(n2218) );
  XOR U3209 ( .A(n3408), .B(in[1189]), .Z(n2504) );
  XOR U3210 ( .A(in[1553]), .B(n3124), .Z(n2119) );
  IV U3211 ( .A(n2119), .Z(n2506) );
  OR U3212 ( .A(n2504), .B(n2506), .Z(n2032) );
  XNOR U3213 ( .A(n2218), .B(n2032), .Z(out[1297]) );
  XOR U3214 ( .A(in[4]), .B(n3083), .Z(n2220) );
  IV U3215 ( .A(n2033), .Z(n4067) );
  XOR U3216 ( .A(in[1190]), .B(n4067), .Z(n2508) );
  XOR U3217 ( .A(in[1554]), .B(n3126), .Z(n2121) );
  IV U3218 ( .A(n2121), .Z(n2510) );
  OR U3219 ( .A(n2508), .B(n2510), .Z(n2034) );
  XNOR U3220 ( .A(n2220), .B(n2034), .Z(out[1298]) );
  XOR U3221 ( .A(in[5]), .B(n3085), .Z(n2222) );
  IV U3222 ( .A(n2035), .Z(n4075) );
  XOR U3223 ( .A(in[1191]), .B(n4075), .Z(n2512) );
  XOR U3224 ( .A(in[1555]), .B(n3128), .Z(n2123) );
  IV U3225 ( .A(n2123), .Z(n2514) );
  OR U3226 ( .A(n2512), .B(n2514), .Z(n2036) );
  XNOR U3227 ( .A(n2222), .B(n2036), .Z(out[1299]) );
  XOR U3228 ( .A(in[666]), .B(n4260), .Z(n2860) );
  IV U3229 ( .A(n3142), .Z(n4082) );
  XOR U3230 ( .A(in[600]), .B(n4082), .Z(n3985) );
  XNOR U3231 ( .A(in[255]), .B(n3294), .Z(n3984) );
  NANDN U3232 ( .A(n3985), .B(n3984), .Z(n2037) );
  XNOR U3233 ( .A(n2860), .B(n2037), .Z(out[129]) );
  XNOR U3234 ( .A(in[202]), .B(n3948), .Z(n4343) );
  XOR U3235 ( .A(in[1422]), .B(n3203), .Z(n4344) );
  XNOR U3236 ( .A(in[1045]), .B(n4495), .Z(n2887) );
  NANDN U3237 ( .A(n4344), .B(n2887), .Z(n2038) );
  XNOR U3238 ( .A(n4343), .B(n2038), .Z(out[12]) );
  XOR U3239 ( .A(in[6]), .B(n3087), .Z(n2224) );
  IV U3240 ( .A(n2039), .Z(n4079) );
  XOR U3241 ( .A(in[1192]), .B(n4079), .Z(n2516) );
  XOR U3242 ( .A(in[1556]), .B(n4062), .Z(n2518) );
  OR U3243 ( .A(n2516), .B(n2518), .Z(n2040) );
  XNOR U3244 ( .A(n2224), .B(n2040), .Z(out[1300]) );
  XOR U3245 ( .A(in[7]), .B(n3089), .Z(n2226) );
  IV U3246 ( .A(n2041), .Z(n4083) );
  XOR U3247 ( .A(in[1193]), .B(n4083), .Z(n2520) );
  XOR U3248 ( .A(in[1557]), .B(n3132), .Z(n2125) );
  IV U3249 ( .A(n2125), .Z(n2522) );
  OR U3250 ( .A(n2520), .B(n2522), .Z(n2042) );
  XNOR U3251 ( .A(n2226), .B(n2042), .Z(out[1301]) );
  XOR U3252 ( .A(in[8]), .B(n4218), .Z(n2229) );
  IV U3253 ( .A(n2043), .Z(n4087) );
  XOR U3254 ( .A(in[1194]), .B(n4087), .Z(n2524) );
  XOR U3255 ( .A(in[1558]), .B(n4074), .Z(n2526) );
  OR U3256 ( .A(n2524), .B(n2526), .Z(n2044) );
  XNOR U3257 ( .A(n2229), .B(n2044), .Z(out[1302]) );
  XOR U3258 ( .A(in[9]), .B(n3092), .Z(n2231) );
  XOR U3259 ( .A(in[1559]), .B(n4078), .Z(n2530) );
  XOR U3260 ( .A(in[1195]), .B(n4092), .Z(n2528) );
  NANDN U3261 ( .A(n2530), .B(n2528), .Z(n2045) );
  XNOR U3262 ( .A(n2231), .B(n2045), .Z(out[1303]) );
  XOR U3263 ( .A(in[10]), .B(n3094), .Z(n2233) );
  XOR U3264 ( .A(in[1560]), .B(n4082), .Z(n2535) );
  XOR U3265 ( .A(in[1196]), .B(n4096), .Z(n2533) );
  NANDN U3266 ( .A(n2535), .B(n2533), .Z(n2046) );
  XNOR U3267 ( .A(n2233), .B(n2046), .Z(out[1304]) );
  XOR U3268 ( .A(in[11]), .B(n3096), .Z(n2235) );
  IV U3269 ( .A(n3144), .Z(n4086) );
  XOR U3270 ( .A(in[1561]), .B(n4086), .Z(n2539) );
  XOR U3271 ( .A(in[1197]), .B(n4100), .Z(n2537) );
  NANDN U3272 ( .A(n2539), .B(n2537), .Z(n2047) );
  XNOR U3273 ( .A(n2235), .B(n2047), .Z(out[1305]) );
  XOR U3274 ( .A(in[12]), .B(n3098), .Z(n2237) );
  IV U3275 ( .A(n3147), .Z(n4090) );
  XOR U3276 ( .A(in[1562]), .B(n4090), .Z(n2543) );
  XOR U3277 ( .A(in[1198]), .B(n4104), .Z(n2541) );
  NANDN U3278 ( .A(n2543), .B(n2541), .Z(n2048) );
  XNOR U3279 ( .A(n2237), .B(n2048), .Z(out[1306]) );
  XOR U3280 ( .A(in[13]), .B(n3102), .Z(n2239) );
  IV U3281 ( .A(n3149), .Z(n4094) );
  XOR U3282 ( .A(in[1563]), .B(n4094), .Z(n2547) );
  XOR U3283 ( .A(in[1199]), .B(n4108), .Z(n2545) );
  NANDN U3284 ( .A(n2547), .B(n2545), .Z(n2049) );
  XNOR U3285 ( .A(n2239), .B(n2049), .Z(out[1307]) );
  XOR U3286 ( .A(in[14]), .B(n3104), .Z(n2241) );
  IV U3287 ( .A(n3028), .Z(n4098) );
  XOR U3288 ( .A(in[1564]), .B(n4098), .Z(n2551) );
  XOR U3289 ( .A(in[1200]), .B(n4112), .Z(n2549) );
  NANDN U3290 ( .A(n2551), .B(n2549), .Z(n2050) );
  XNOR U3291 ( .A(n2241), .B(n2050), .Z(out[1308]) );
  XOR U3292 ( .A(in[15]), .B(n4237), .Z(n2243) );
  IV U3293 ( .A(n3030), .Z(n4102) );
  XOR U3294 ( .A(in[1565]), .B(n4102), .Z(n2555) );
  XOR U3295 ( .A(in[1201]), .B(n4120), .Z(n2553) );
  NANDN U3296 ( .A(n2555), .B(n2553), .Z(n2051) );
  XNOR U3297 ( .A(n2243), .B(n2051), .Z(out[1309]) );
  XOR U3298 ( .A(in[667]), .B(n4261), .Z(n2746) );
  IV U3299 ( .A(n2746), .Z(n2862) );
  XOR U3300 ( .A(in[601]), .B(n4086), .Z(n4029) );
  XNOR U3301 ( .A(in[192]), .B(n3297), .Z(n4026) );
  NANDN U3302 ( .A(n4029), .B(n4026), .Z(n2052) );
  XOR U3303 ( .A(n2862), .B(n2052), .Z(out[130]) );
  XOR U3304 ( .A(in[16]), .B(n4240), .Z(n2245) );
  IV U3305 ( .A(n3032), .Z(n4106) );
  XOR U3306 ( .A(in[1566]), .B(n4106), .Z(n2559) );
  XOR U3307 ( .A(in[1202]), .B(n4124), .Z(n2557) );
  NANDN U3308 ( .A(n2559), .B(n2557), .Z(n2053) );
  XNOR U3309 ( .A(n2245), .B(n2053), .Z(out[1310]) );
  XOR U3310 ( .A(in[17]), .B(n4241), .Z(n2247) );
  IV U3311 ( .A(n3034), .Z(n4110) );
  XOR U3312 ( .A(in[1567]), .B(n4110), .Z(n2562) );
  XOR U3313 ( .A(in[1203]), .B(n4128), .Z(n2561) );
  NANDN U3314 ( .A(n2562), .B(n2561), .Z(n2054) );
  XNOR U3315 ( .A(n2247), .B(n2054), .Z(out[1311]) );
  XOR U3316 ( .A(in[18]), .B(n4246), .Z(n2250) );
  IV U3317 ( .A(n3036), .Z(n4118) );
  XOR U3318 ( .A(in[1568]), .B(n4118), .Z(n2568) );
  XOR U3319 ( .A(in[1204]), .B(n4132), .Z(n2566) );
  NANDN U3320 ( .A(n2568), .B(n2566), .Z(n2055) );
  XNOR U3321 ( .A(n2250), .B(n2055), .Z(out[1312]) );
  XOR U3322 ( .A(in[19]), .B(n4249), .Z(n2252) );
  XOR U3323 ( .A(in[1569]), .B(n3038), .Z(n2129) );
  IV U3324 ( .A(n2129), .Z(n2572) );
  XOR U3325 ( .A(in[1205]), .B(n4136), .Z(n2570) );
  NANDN U3326 ( .A(n2572), .B(n2570), .Z(n2056) );
  XNOR U3327 ( .A(n2252), .B(n2056), .Z(out[1313]) );
  XOR U3328 ( .A(in[20]), .B(n4252), .Z(n2254) );
  XOR U3329 ( .A(in[1570]), .B(n2168), .Z(n2131) );
  IV U3330 ( .A(n2131), .Z(n2578) );
  XOR U3331 ( .A(in[1206]), .B(n4140), .Z(n2576) );
  NANDN U3332 ( .A(n2578), .B(n2576), .Z(n2057) );
  XNOR U3333 ( .A(n2254), .B(n2057), .Z(out[1314]) );
  XOR U3334 ( .A(in[21]), .B(n4255), .Z(n2256) );
  XOR U3335 ( .A(in[1571]), .B(n3041), .Z(n2133) );
  IV U3336 ( .A(n2133), .Z(n2582) );
  XOR U3337 ( .A(in[1207]), .B(n4144), .Z(n2580) );
  NANDN U3338 ( .A(n2582), .B(n2580), .Z(n2058) );
  XNOR U3339 ( .A(n2256), .B(n2058), .Z(out[1315]) );
  XOR U3340 ( .A(in[22]), .B(n4256), .Z(n2258) );
  XOR U3341 ( .A(in[1572]), .B(n3043), .Z(n2136) );
  IV U3342 ( .A(n2136), .Z(n2586) );
  XOR U3343 ( .A(in[1208]), .B(n4148), .Z(n2584) );
  NANDN U3344 ( .A(n2586), .B(n2584), .Z(n2059) );
  XNOR U3345 ( .A(n2258), .B(n2059), .Z(out[1316]) );
  XOR U3346 ( .A(in[23]), .B(n4257), .Z(n2260) );
  XNOR U3347 ( .A(in[1573]), .B(n4138), .Z(n2138) );
  IV U3348 ( .A(n2138), .Z(n2590) );
  XOR U3349 ( .A(in[1209]), .B(n4152), .Z(n2588) );
  NANDN U3350 ( .A(n2590), .B(n2588), .Z(n2060) );
  XNOR U3351 ( .A(n2260), .B(n2060), .Z(out[1317]) );
  XOR U3352 ( .A(in[24]), .B(n4258), .Z(n2262) );
  XNOR U3353 ( .A(in[1574]), .B(n4142), .Z(n2594) );
  XOR U3354 ( .A(in[1210]), .B(n4156), .Z(n2592) );
  NAND U3355 ( .A(n2594), .B(n2592), .Z(n2061) );
  XNOR U3356 ( .A(n2262), .B(n2061), .Z(out[1318]) );
  XOR U3357 ( .A(in[25]), .B(n4259), .Z(n2264) );
  XOR U3358 ( .A(in[1211]), .B(n4166), .Z(n2596) );
  XNOR U3359 ( .A(in[1575]), .B(n4146), .Z(n2141) );
  IV U3360 ( .A(n2141), .Z(n2598) );
  OR U3361 ( .A(n2596), .B(n2598), .Z(n2062) );
  XNOR U3362 ( .A(n2264), .B(n2062), .Z(out[1319]) );
  XOR U3363 ( .A(in[668]), .B(n4264), .Z(n2748) );
  IV U3364 ( .A(n2748), .Z(n2864) );
  XOR U3365 ( .A(in[602]), .B(n4090), .Z(n4073) );
  XNOR U3366 ( .A(in[193]), .B(n3300), .Z(n4070) );
  NANDN U3367 ( .A(n4073), .B(n4070), .Z(n2063) );
  XOR U3368 ( .A(n2864), .B(n2063), .Z(out[131]) );
  XOR U3369 ( .A(in[26]), .B(n4260), .Z(n2266) );
  XOR U3370 ( .A(in[1212]), .B(n4170), .Z(n2600) );
  XNOR U3371 ( .A(in[1576]), .B(n4150), .Z(n2143) );
  IV U3372 ( .A(n2143), .Z(n2602) );
  OR U3373 ( .A(n2600), .B(n2602), .Z(n2064) );
  XNOR U3374 ( .A(n2266), .B(n2064), .Z(out[1320]) );
  XOR U3375 ( .A(in[27]), .B(n4261), .Z(n2268) );
  XOR U3376 ( .A(in[1213]), .B(n4174), .Z(n2604) );
  XNOR U3377 ( .A(in[1577]), .B(n4154), .Z(n2145) );
  IV U3378 ( .A(n2145), .Z(n2606) );
  OR U3379 ( .A(n2604), .B(n2606), .Z(n2065) );
  XNOR U3380 ( .A(n2268), .B(n2065), .Z(out[1321]) );
  XOR U3381 ( .A(in[28]), .B(n4264), .Z(n2271) );
  XNOR U3382 ( .A(in[1578]), .B(n4164), .Z(n2147) );
  IV U3383 ( .A(n2147), .Z(n2610) );
  XOR U3384 ( .A(in[1214]), .B(n4178), .Z(n2608) );
  NANDN U3385 ( .A(n2610), .B(n2608), .Z(n2066) );
  XNOR U3386 ( .A(n2271), .B(n2066), .Z(out[1322]) );
  XOR U3387 ( .A(in[29]), .B(n4265), .Z(n2273) );
  XOR U3388 ( .A(in[1215]), .B(n3294), .Z(n2612) );
  XNOR U3389 ( .A(in[1579]), .B(n4168), .Z(n2149) );
  IV U3390 ( .A(n2149), .Z(n2614) );
  OR U3391 ( .A(n2612), .B(n2614), .Z(n2067) );
  XNOR U3392 ( .A(n2273), .B(n2067), .Z(out[1323]) );
  XOR U3393 ( .A(in[30]), .B(n4266), .Z(n2275) );
  XOR U3394 ( .A(in[1152]), .B(n3297), .Z(n2618) );
  XNOR U3395 ( .A(in[1580]), .B(n4172), .Z(n2151) );
  IV U3396 ( .A(n2151), .Z(n2620) );
  OR U3397 ( .A(n2618), .B(n2620), .Z(n2068) );
  XNOR U3398 ( .A(n2275), .B(n2068), .Z(out[1324]) );
  XOR U3399 ( .A(in[31]), .B(n4267), .Z(n2277) );
  XOR U3400 ( .A(in[1153]), .B(n3300), .Z(n2622) );
  XNOR U3401 ( .A(in[1581]), .B(n4176), .Z(n2153) );
  IV U3402 ( .A(n2153), .Z(n2624) );
  OR U3403 ( .A(n2622), .B(n2624), .Z(n2069) );
  XNOR U3404 ( .A(n2277), .B(n2069), .Z(out[1325]) );
  XOR U3405 ( .A(in[32]), .B(n4270), .Z(n2279) );
  XOR U3406 ( .A(in[1154]), .B(n3307), .Z(n2626) );
  XNOR U3407 ( .A(in[1582]), .B(n3900), .Z(n2156) );
  IV U3408 ( .A(n2156), .Z(n2628) );
  OR U3409 ( .A(n2626), .B(n2628), .Z(n2070) );
  XNOR U3410 ( .A(n2279), .B(n2070), .Z(out[1326]) );
  XOR U3411 ( .A(in[33]), .B(n4273), .Z(n2281) );
  XOR U3412 ( .A(in[1155]), .B(n3310), .Z(n2630) );
  XNOR U3413 ( .A(in[1583]), .B(n3904), .Z(n2158) );
  IV U3414 ( .A(n2158), .Z(n2632) );
  OR U3415 ( .A(n2630), .B(n2632), .Z(n2071) );
  XNOR U3416 ( .A(n2281), .B(n2071), .Z(out[1327]) );
  XOR U3417 ( .A(in[34]), .B(n4276), .Z(n2283) );
  XOR U3418 ( .A(in[1156]), .B(n3313), .Z(n2634) );
  XNOR U3419 ( .A(in[1584]), .B(n3908), .Z(n2160) );
  IV U3420 ( .A(n2160), .Z(n2636) );
  OR U3421 ( .A(n2634), .B(n2636), .Z(n2072) );
  XNOR U3422 ( .A(n2283), .B(n2072), .Z(out[1328]) );
  IV U3423 ( .A(n4279), .Z(n3146) );
  XOR U3424 ( .A(in[35]), .B(n3146), .Z(n2285) );
  XOR U3425 ( .A(in[1157]), .B(n3316), .Z(n2638) );
  XNOR U3426 ( .A(in[1585]), .B(n3912), .Z(n2162) );
  IV U3427 ( .A(n2162), .Z(n2640) );
  OR U3428 ( .A(n2638), .B(n2640), .Z(n2073) );
  XNOR U3429 ( .A(n2285), .B(n2073), .Z(out[1329]) );
  XOR U3430 ( .A(in[669]), .B(n4265), .Z(n2750) );
  IV U3431 ( .A(n2750), .Z(n2869) );
  XOR U3432 ( .A(in[603]), .B(n4094), .Z(n4117) );
  XNOR U3433 ( .A(in[194]), .B(n3307), .Z(n4114) );
  NANDN U3434 ( .A(n4117), .B(n4114), .Z(n2074) );
  XOR U3435 ( .A(n2869), .B(n2074), .Z(out[132]) );
  XOR U3436 ( .A(in[36]), .B(n4282), .Z(n2287) );
  XOR U3437 ( .A(in[1158]), .B(n3319), .Z(n2642) );
  XNOR U3438 ( .A(in[1586]), .B(n3916), .Z(n2164) );
  IV U3439 ( .A(n2164), .Z(n2644) );
  OR U3440 ( .A(n2642), .B(n2644), .Z(n2075) );
  XNOR U3441 ( .A(n2287), .B(n2075), .Z(out[1330]) );
  XOR U3442 ( .A(in[37]), .B(n4284), .Z(n2289) );
  XOR U3443 ( .A(in[1159]), .B(n3322), .Z(n2646) );
  XOR U3444 ( .A(in[1587]), .B(n2573), .Z(n2648) );
  OR U3445 ( .A(n2646), .B(n2648), .Z(n2076) );
  XNOR U3446 ( .A(n2289), .B(n2076), .Z(out[1331]) );
  XOR U3447 ( .A(in[38]), .B(n4290), .Z(n2292) );
  XOR U3448 ( .A(in[1160]), .B(n3937), .Z(n2650) );
  XOR U3449 ( .A(in[1588]), .B(n2615), .Z(n2652) );
  OR U3450 ( .A(n2650), .B(n2652), .Z(n2077) );
  XNOR U3451 ( .A(n2292), .B(n2077), .Z(out[1332]) );
  XOR U3452 ( .A(in[39]), .B(n4292), .Z(n2294) );
  XOR U3453 ( .A(in[1161]), .B(n3944), .Z(n2654) );
  XOR U3454 ( .A(in[1589]), .B(n2657), .Z(n2656) );
  OR U3455 ( .A(n2654), .B(n2656), .Z(n2078) );
  XNOR U3456 ( .A(n2294), .B(n2078), .Z(out[1333]) );
  XOR U3457 ( .A(in[40]), .B(n4294), .Z(n2297) );
  XOR U3458 ( .A(in[1162]), .B(n3948), .Z(n2660) );
  XNOR U3459 ( .A(in[1590]), .B(n3069), .Z(n2662) );
  NANDN U3460 ( .A(n2660), .B(n2662), .Z(n2079) );
  XNOR U3461 ( .A(n2297), .B(n2079), .Z(out[1334]) );
  XOR U3462 ( .A(in[41]), .B(n4296), .Z(n2299) );
  XOR U3463 ( .A(in[1163]), .B(n3952), .Z(n2664) );
  XNOR U3464 ( .A(in[1591]), .B(n3071), .Z(n2666) );
  NANDN U3465 ( .A(n2664), .B(n2666), .Z(n2080) );
  XNOR U3466 ( .A(n2299), .B(n2080), .Z(out[1335]) );
  XOR U3467 ( .A(in[42]), .B(n4298), .Z(n2301) );
  XOR U3468 ( .A(in[1164]), .B(n3956), .Z(n2668) );
  XNOR U3469 ( .A(in[1592]), .B(n3074), .Z(n2670) );
  NANDN U3470 ( .A(n2668), .B(n2670), .Z(n2081) );
  XNOR U3471 ( .A(n2301), .B(n2081), .Z(out[1336]) );
  XOR U3472 ( .A(in[43]), .B(n4300), .Z(n2303) );
  XOR U3473 ( .A(in[1165]), .B(n3960), .Z(n2672) );
  XOR U3474 ( .A(in[1593]), .B(n2702), .Z(n2674) );
  OR U3475 ( .A(n2672), .B(n2674), .Z(n2082) );
  XNOR U3476 ( .A(n2303), .B(n2082), .Z(out[1337]) );
  XOR U3477 ( .A(in[44]), .B(n4302), .Z(n2305) );
  XOR U3478 ( .A(in[1166]), .B(n3964), .Z(n2676) );
  XOR U3479 ( .A(in[1594]), .B(n2704), .Z(n2678) );
  OR U3480 ( .A(n2676), .B(n2678), .Z(n2083) );
  XNOR U3481 ( .A(n2305), .B(n2083), .Z(out[1338]) );
  XOR U3482 ( .A(in[45]), .B(n4304), .Z(n2307) );
  XOR U3483 ( .A(in[1167]), .B(n3968), .Z(n2680) );
  XNOR U3484 ( .A(in[1595]), .B(n3955), .Z(n2172) );
  IV U3485 ( .A(n2172), .Z(n2682) );
  OR U3486 ( .A(n2680), .B(n2682), .Z(n2084) );
  XNOR U3487 ( .A(n2307), .B(n2084), .Z(out[1339]) );
  XOR U3488 ( .A(in[670]), .B(n4266), .Z(n2752) );
  IV U3489 ( .A(n2752), .Z(n2871) );
  XOR U3490 ( .A(in[604]), .B(n4098), .Z(n4161) );
  XNOR U3491 ( .A(in[195]), .B(n3310), .Z(n4158) );
  NANDN U3492 ( .A(n4161), .B(n4158), .Z(n2085) );
  XOR U3493 ( .A(n2871), .B(n2085), .Z(out[133]) );
  XOR U3494 ( .A(in[46]), .B(n4306), .Z(n2309) );
  XOR U3495 ( .A(in[1168]), .B(n3972), .Z(n2684) );
  XNOR U3496 ( .A(in[1596]), .B(n3959), .Z(n2174) );
  IV U3497 ( .A(n2174), .Z(n2686) );
  OR U3498 ( .A(n2684), .B(n2686), .Z(n2086) );
  XNOR U3499 ( .A(n2309), .B(n2086), .Z(out[1340]) );
  XOR U3500 ( .A(in[47]), .B(n4308), .Z(n2311) );
  XOR U3501 ( .A(in[1169]), .B(n3976), .Z(n2688) );
  XNOR U3502 ( .A(in[1597]), .B(n3963), .Z(n2176) );
  IV U3503 ( .A(n2176), .Z(n2690) );
  OR U3504 ( .A(n2688), .B(n2690), .Z(n2087) );
  XNOR U3505 ( .A(n2311), .B(n2087), .Z(out[1341]) );
  XOR U3506 ( .A(in[48]), .B(n4315), .Z(n2314) );
  XOR U3507 ( .A(in[1170]), .B(n3980), .Z(n2692) );
  XNOR U3508 ( .A(in[1598]), .B(n3967), .Z(n2178) );
  IV U3509 ( .A(n2178), .Z(n2694) );
  OR U3510 ( .A(n2692), .B(n2694), .Z(n2088) );
  XNOR U3511 ( .A(n2314), .B(n2088), .Z(out[1342]) );
  XOR U3512 ( .A(in[49]), .B(n4318), .Z(n2316) );
  XNOR U3513 ( .A(in[1171]), .B(n3987), .Z(n2696) );
  XNOR U3514 ( .A(in[1599]), .B(n3971), .Z(n2697) );
  NANDN U3515 ( .A(n2696), .B(n2697), .Z(n2089) );
  XNOR U3516 ( .A(n2316), .B(n2089), .Z(out[1343]) );
  XNOR U3517 ( .A(in[427]), .B(n4351), .Z(n2318) );
  NOR U3518 ( .A(n2439), .B(n2181), .Z(n2090) );
  XNOR U3519 ( .A(n2318), .B(n2090), .Z(out[1344]) );
  XNOR U3520 ( .A(in[428]), .B(n4354), .Z(n2320) );
  NOR U3521 ( .A(n2442), .B(n2183), .Z(n2091) );
  XNOR U3522 ( .A(n2320), .B(n2091), .Z(out[1345]) );
  XNOR U3523 ( .A(in[429]), .B(n4357), .Z(n2322) );
  NOR U3524 ( .A(n2092), .B(n2186), .Z(n2093) );
  XNOR U3525 ( .A(n2322), .B(n2093), .Z(out[1346]) );
  XNOR U3526 ( .A(in[430]), .B(n4360), .Z(n2324) );
  NOR U3527 ( .A(n2449), .B(n2188), .Z(n2094) );
  XNOR U3528 ( .A(n2324), .B(n2094), .Z(out[1347]) );
  XNOR U3529 ( .A(in[431]), .B(n4362), .Z(n2326) );
  NOR U3530 ( .A(n2095), .B(n2190), .Z(n2096) );
  XNOR U3531 ( .A(n2326), .B(n2096), .Z(out[1348]) );
  XNOR U3532 ( .A(in[432]), .B(n4365), .Z(n2328) );
  NOR U3533 ( .A(n2097), .B(n2192), .Z(n2098) );
  XNOR U3534 ( .A(n2328), .B(n2098), .Z(out[1349]) );
  XOR U3535 ( .A(in[671]), .B(n4267), .Z(n2754) );
  IV U3536 ( .A(n2754), .Z(n2873) );
  XOR U3537 ( .A(in[605]), .B(n4102), .Z(n4199) );
  XNOR U3538 ( .A(in[196]), .B(n3313), .Z(n4196) );
  NANDN U3539 ( .A(n4199), .B(n4196), .Z(n2099) );
  XOR U3540 ( .A(n2873), .B(n2099), .Z(out[134]) );
  XNOR U3541 ( .A(in[433]), .B(n4368), .Z(n2330) );
  NOR U3542 ( .A(n2100), .B(n2194), .Z(n2101) );
  XNOR U3543 ( .A(n2330), .B(n2101), .Z(out[1350]) );
  XNOR U3544 ( .A(in[434]), .B(n4371), .Z(n2332) );
  NOR U3545 ( .A(n2102), .B(n2196), .Z(n2103) );
  XNOR U3546 ( .A(n2332), .B(n2103), .Z(out[1351]) );
  XNOR U3547 ( .A(in[435]), .B(n4378), .Z(n2335) );
  NOR U3548 ( .A(n2469), .B(n2198), .Z(n2104) );
  XNOR U3549 ( .A(n2335), .B(n2104), .Z(out[1352]) );
  XNOR U3550 ( .A(in[436]), .B(n4381), .Z(n2338) );
  NOR U3551 ( .A(n2472), .B(n2200), .Z(n2105) );
  XNOR U3552 ( .A(n2338), .B(n2105), .Z(out[1353]) );
  XNOR U3553 ( .A(in[437]), .B(n4384), .Z(n2341) );
  NOR U3554 ( .A(n2475), .B(n2202), .Z(n2106) );
  XNOR U3555 ( .A(n2341), .B(n2106), .Z(out[1354]) );
  XNOR U3556 ( .A(in[438]), .B(n4387), .Z(n2344) );
  NOR U3557 ( .A(n2481), .B(n2204), .Z(n2107) );
  XNOR U3558 ( .A(n2344), .B(n2107), .Z(out[1355]) );
  XNOR U3559 ( .A(in[439]), .B(n4390), .Z(n2347) );
  NOR U3560 ( .A(n2485), .B(n2207), .Z(n2108) );
  XNOR U3561 ( .A(n2347), .B(n2108), .Z(out[1356]) );
  XNOR U3562 ( .A(in[440]), .B(n4392), .Z(n2350) );
  NOR U3563 ( .A(n2486), .B(n2209), .Z(n2109) );
  XNOR U3564 ( .A(n2350), .B(n2109), .Z(out[1357]) );
  XNOR U3565 ( .A(in[441]), .B(n4395), .Z(n2353) );
  NOR U3566 ( .A(n2110), .B(n2211), .Z(n2111) );
  XNOR U3567 ( .A(n2353), .B(n2111), .Z(out[1358]) );
  XOR U3568 ( .A(in[442]), .B(n2112), .Z(n2355) );
  NOR U3569 ( .A(n2113), .B(n2213), .Z(n2114) );
  XOR U3570 ( .A(n2355), .B(n2114), .Z(out[1359]) );
  XOR U3571 ( .A(in[672]), .B(n4270), .Z(n2756) );
  IV U3572 ( .A(n2756), .Z(n2875) );
  XOR U3573 ( .A(in[606]), .B(n4106), .Z(n4217) );
  XNOR U3574 ( .A(in[197]), .B(n3316), .Z(n4448) );
  NANDN U3575 ( .A(n4217), .B(n4448), .Z(n2115) );
  XOR U3576 ( .A(n2875), .B(n2115), .Z(out[135]) );
  XOR U3577 ( .A(in[443]), .B(n2116), .Z(n2357) );
  NOR U3578 ( .A(n2117), .B(n2216), .Z(n2118) );
  XOR U3579 ( .A(n2357), .B(n2118), .Z(out[1360]) );
  XNOR U3580 ( .A(in[444]), .B(n4404), .Z(n2358) );
  NOR U3581 ( .A(n2119), .B(n2218), .Z(n2120) );
  XNOR U3582 ( .A(n2358), .B(n2120), .Z(out[1361]) );
  XNOR U3583 ( .A(in[445]), .B(n4411), .Z(n2361) );
  NOR U3584 ( .A(n2121), .B(n2220), .Z(n2122) );
  XNOR U3585 ( .A(n2361), .B(n2122), .Z(out[1362]) );
  XNOR U3586 ( .A(in[446]), .B(n4414), .Z(n2363) );
  NOR U3587 ( .A(n2123), .B(n2222), .Z(n2124) );
  XNOR U3588 ( .A(n2363), .B(n2124), .Z(out[1363]) );
  XNOR U3589 ( .A(in[447]), .B(n4417), .Z(n2365) );
  XNOR U3590 ( .A(in[384]), .B(n4420), .Z(n2367) );
  NOR U3591 ( .A(n2125), .B(n2226), .Z(n2126) );
  XNOR U3592 ( .A(n2367), .B(n2126), .Z(out[1365]) );
  XNOR U3593 ( .A(in[385]), .B(n4423), .Z(n2369) );
  XNOR U3594 ( .A(in[386]), .B(n4426), .Z(n2371) );
  XNOR U3595 ( .A(in[387]), .B(n4429), .Z(n2373) );
  XNOR U3596 ( .A(in[388]), .B(n4432), .Z(n2375) );
  XOR U3597 ( .A(in[673]), .B(n4273), .Z(n2763) );
  IV U3598 ( .A(n2763), .Z(n2877) );
  XOR U3599 ( .A(in[607]), .B(n4110), .Z(n4245) );
  XNOR U3600 ( .A(in[198]), .B(n3319), .Z(n4738) );
  NANDN U3601 ( .A(n4245), .B(n4738), .Z(n2127) );
  XOR U3602 ( .A(n2877), .B(n2127), .Z(out[136]) );
  XNOR U3603 ( .A(in[389]), .B(n4435), .Z(n2377) );
  XOR U3604 ( .A(in[390]), .B(n2128), .Z(n2379) );
  XNOR U3605 ( .A(in[391]), .B(n4449), .Z(n2382) );
  XNOR U3606 ( .A(in[392]), .B(n4452), .Z(n2384) );
  XNOR U3607 ( .A(in[393]), .B(n4455), .Z(n2386) );
  XNOR U3608 ( .A(in[394]), .B(n4458), .Z(n2388) );
  XNOR U3609 ( .A(in[395]), .B(n4461), .Z(n2390) );
  XNOR U3610 ( .A(n4464), .B(in[396]), .Z(n2392) );
  NOR U3611 ( .A(n2129), .B(n2252), .Z(n2130) );
  XOR U3612 ( .A(n2392), .B(n2130), .Z(out[1377]) );
  XNOR U3613 ( .A(n4467), .B(in[397]), .Z(n2393) );
  NOR U3614 ( .A(n2131), .B(n2254), .Z(n2132) );
  XOR U3615 ( .A(n2393), .B(n2132), .Z(out[1378]) );
  XNOR U3616 ( .A(n4470), .B(in[398]), .Z(n2394) );
  NOR U3617 ( .A(n2133), .B(n2256), .Z(n2134) );
  XOR U3618 ( .A(n2394), .B(n2134), .Z(out[1379]) );
  XOR U3619 ( .A(in[674]), .B(n4276), .Z(n2765) );
  IV U3620 ( .A(n2765), .Z(n2879) );
  XOR U3621 ( .A(in[608]), .B(n4118), .Z(n4263) );
  XNOR U3622 ( .A(in[199]), .B(n3322), .Z(n5167) );
  NANDN U3623 ( .A(n4263), .B(n5167), .Z(n2135) );
  XOR U3624 ( .A(n2879), .B(n2135), .Z(out[137]) );
  XNOR U3625 ( .A(n4473), .B(in[399]), .Z(n2395) );
  NOR U3626 ( .A(n2136), .B(n2258), .Z(n2137) );
  XOR U3627 ( .A(n2395), .B(n2137), .Z(out[1380]) );
  XNOR U3628 ( .A(n4476), .B(in[400]), .Z(n2396) );
  NOR U3629 ( .A(n2138), .B(n2260), .Z(n2139) );
  XOR U3630 ( .A(n2396), .B(n2139), .Z(out[1381]) );
  XNOR U3631 ( .A(n4483), .B(in[401]), .Z(n2398) );
  NOR U3632 ( .A(n2594), .B(n2262), .Z(n2140) );
  XOR U3633 ( .A(n2398), .B(n2140), .Z(out[1382]) );
  XNOR U3634 ( .A(n4486), .B(in[402]), .Z(n2399) );
  NOR U3635 ( .A(n2141), .B(n2264), .Z(n2142) );
  XOR U3636 ( .A(n2399), .B(n2142), .Z(out[1383]) );
  XNOR U3637 ( .A(n4489), .B(in[403]), .Z(n2400) );
  NOR U3638 ( .A(n2143), .B(n2266), .Z(n2144) );
  XOR U3639 ( .A(n2400), .B(n2144), .Z(out[1384]) );
  XNOR U3640 ( .A(in[404]), .B(n4492), .Z(n2401) );
  NOR U3641 ( .A(n2145), .B(n2268), .Z(n2146) );
  XOR U3642 ( .A(n2401), .B(n2146), .Z(out[1385]) );
  XNOR U3643 ( .A(in[405]), .B(n4495), .Z(n2402) );
  NOR U3644 ( .A(n2147), .B(n2271), .Z(n2148) );
  XOR U3645 ( .A(n2402), .B(n2148), .Z(out[1386]) );
  XNOR U3646 ( .A(in[406]), .B(n4498), .Z(n2403) );
  NOR U3647 ( .A(n2149), .B(n2273), .Z(n2150) );
  XOR U3648 ( .A(n2403), .B(n2150), .Z(out[1387]) );
  XNOR U3649 ( .A(in[407]), .B(n4501), .Z(n2404) );
  NOR U3650 ( .A(n2151), .B(n2275), .Z(n2152) );
  XOR U3651 ( .A(n2404), .B(n2152), .Z(out[1388]) );
  XNOR U3652 ( .A(in[408]), .B(n4504), .Z(n2405) );
  NOR U3653 ( .A(n2153), .B(n2277), .Z(n2154) );
  XOR U3654 ( .A(n2405), .B(n2154), .Z(out[1389]) );
  XOR U3655 ( .A(in[675]), .B(n4279), .Z(n2882) );
  IV U3656 ( .A(n3038), .Z(n4122) );
  XOR U3657 ( .A(in[609]), .B(n4122), .Z(n4289) );
  NANDN U3658 ( .A(n4289), .B(n4286), .Z(n2155) );
  XOR U3659 ( .A(n2882), .B(n2155), .Z(out[138]) );
  XNOR U3660 ( .A(in[409]), .B(n4507), .Z(n2406) );
  NOR U3661 ( .A(n2156), .B(n2279), .Z(n2157) );
  XOR U3662 ( .A(n2406), .B(n2157), .Z(out[1390]) );
  XNOR U3663 ( .A(in[410]), .B(n4510), .Z(n2407) );
  NOR U3664 ( .A(n2158), .B(n2281), .Z(n2159) );
  XOR U3665 ( .A(n2407), .B(n2159), .Z(out[1391]) );
  XOR U3666 ( .A(in[411]), .B(n4517), .Z(n2409) );
  NOR U3667 ( .A(n2160), .B(n2283), .Z(n2161) );
  XOR U3668 ( .A(n2409), .B(n2161), .Z(out[1392]) );
  XOR U3669 ( .A(in[412]), .B(n4520), .Z(n2410) );
  NOR U3670 ( .A(n2162), .B(n2285), .Z(n2163) );
  XOR U3671 ( .A(n2410), .B(n2163), .Z(out[1393]) );
  XOR U3672 ( .A(in[413]), .B(n4523), .Z(n2411) );
  NOR U3673 ( .A(n2164), .B(n2287), .Z(n2165) );
  XOR U3674 ( .A(n2411), .B(n2165), .Z(out[1394]) );
  XOR U3675 ( .A(in[414]), .B(n4526), .Z(n2412) );
  XOR U3676 ( .A(in[415]), .B(n4530), .Z(n2414) );
  XOR U3677 ( .A(in[416]), .B(n4534), .Z(n2416) );
  XNOR U3678 ( .A(in[417]), .B(n4538), .Z(n2418) );
  NOR U3679 ( .A(n2662), .B(n2297), .Z(n2166) );
  XOR U3680 ( .A(n2418), .B(n2166), .Z(out[1398]) );
  XNOR U3681 ( .A(in[418]), .B(n4542), .Z(n2419) );
  NOR U3682 ( .A(n2666), .B(n2299), .Z(n2167) );
  XOR U3683 ( .A(n2419), .B(n2167), .Z(out[1399]) );
  XOR U3684 ( .A(in[676]), .B(n4282), .Z(n2884) );
  IV U3685 ( .A(n2168), .Z(n4126) );
  XOR U3686 ( .A(in[610]), .B(n4126), .Z(n4314) );
  NANDN U3687 ( .A(n4314), .B(n4311), .Z(n2169) );
  XNOR U3688 ( .A(n2884), .B(n2169), .Z(out[139]) );
  XNOR U3689 ( .A(in[203]), .B(n3952), .Z(n4374) );
  XOR U3690 ( .A(in[1423]), .B(n3206), .Z(n4375) );
  XNOR U3691 ( .A(in[1046]), .B(n4498), .Z(n2889) );
  NANDN U3692 ( .A(n4375), .B(n2889), .Z(n2170) );
  XNOR U3693 ( .A(n4374), .B(n2170), .Z(out[13]) );
  XNOR U3694 ( .A(in[419]), .B(n4546), .Z(n2420) );
  NOR U3695 ( .A(n2670), .B(n2301), .Z(n2171) );
  XOR U3696 ( .A(n2420), .B(n2171), .Z(out[1400]) );
  XNOR U3697 ( .A(in[420]), .B(n4550), .Z(n2421) );
  XNOR U3698 ( .A(in[421]), .B(n4556), .Z(n2424) );
  XNOR U3699 ( .A(in[422]), .B(n4558), .Z(n2426) );
  NOR U3700 ( .A(n2172), .B(n2307), .Z(n2173) );
  XNOR U3701 ( .A(n2426), .B(n2173), .Z(out[1403]) );
  XNOR U3702 ( .A(in[423]), .B(n4339), .Z(n2428) );
  NOR U3703 ( .A(n2174), .B(n2309), .Z(n2175) );
  XNOR U3704 ( .A(n2428), .B(n2175), .Z(out[1404]) );
  XNOR U3705 ( .A(in[424]), .B(n4341), .Z(n2431) );
  NOR U3706 ( .A(n2176), .B(n2311), .Z(n2177) );
  XNOR U3707 ( .A(n2431), .B(n2177), .Z(out[1405]) );
  XNOR U3708 ( .A(in[425]), .B(n4347), .Z(n2433) );
  NOR U3709 ( .A(n2178), .B(n2314), .Z(n2179) );
  XNOR U3710 ( .A(n2433), .B(n2179), .Z(out[1406]) );
  XNOR U3711 ( .A(in[426]), .B(n4349), .Z(n2435) );
  NOR U3712 ( .A(n2697), .B(n2316), .Z(n2180) );
  XNOR U3713 ( .A(n2435), .B(n2180), .Z(out[1407]) );
  XOR U3714 ( .A(in[789]), .B(n4016), .Z(n2437) );
  NAND U3715 ( .A(n2181), .B(n2318), .Z(n2182) );
  XOR U3716 ( .A(n2437), .B(n2182), .Z(out[1408]) );
  IV U3717 ( .A(n2775), .Z(n4020) );
  XOR U3718 ( .A(in[790]), .B(n4020), .Z(n2440) );
  NAND U3719 ( .A(n2183), .B(n2320), .Z(n2184) );
  XOR U3720 ( .A(n2440), .B(n2184), .Z(out[1409]) );
  XOR U3721 ( .A(in[677]), .B(n4284), .Z(n2886) );
  IV U3722 ( .A(n3041), .Z(n4130) );
  XOR U3723 ( .A(in[611]), .B(n4130), .Z(n4346) );
  NANDN U3724 ( .A(n4346), .B(n4343), .Z(n2185) );
  XNOR U3725 ( .A(n2886), .B(n2185), .Z(out[140]) );
  IV U3726 ( .A(n2782), .Z(n4024) );
  XOR U3727 ( .A(in[791]), .B(n4024), .Z(n2443) );
  NAND U3728 ( .A(n2186), .B(n2322), .Z(n2187) );
  XOR U3729 ( .A(n2443), .B(n2187), .Z(out[1410]) );
  IV U3730 ( .A(n2796), .Z(n4032) );
  XOR U3731 ( .A(in[792]), .B(n4032), .Z(n2447) );
  NAND U3732 ( .A(n2188), .B(n2324), .Z(n2189) );
  XOR U3733 ( .A(n2447), .B(n2189), .Z(out[1411]) );
  IV U3734 ( .A(n2819), .Z(n4036) );
  XOR U3735 ( .A(in[793]), .B(n4036), .Z(n2453) );
  NAND U3736 ( .A(n2190), .B(n2326), .Z(n2191) );
  XOR U3737 ( .A(n2453), .B(n2191), .Z(out[1412]) );
  IV U3738 ( .A(n2842), .Z(n4040) );
  XOR U3739 ( .A(in[794]), .B(n4040), .Z(n2457) );
  NAND U3740 ( .A(n2192), .B(n2328), .Z(n2193) );
  XOR U3741 ( .A(n2457), .B(n2193), .Z(out[1413]) );
  IV U3742 ( .A(n2866), .Z(n4044) );
  XOR U3743 ( .A(in[795]), .B(n4044), .Z(n2461) );
  NAND U3744 ( .A(n2194), .B(n2330), .Z(n2195) );
  XOR U3745 ( .A(n2461), .B(n2195), .Z(out[1414]) );
  IV U3746 ( .A(n2890), .Z(n4048) );
  XOR U3747 ( .A(in[796]), .B(n4048), .Z(n2465) );
  NAND U3748 ( .A(n2196), .B(n2332), .Z(n2197) );
  XOR U3749 ( .A(n2465), .B(n2197), .Z(out[1415]) );
  IV U3750 ( .A(n2923), .Z(n4052) );
  XOR U3751 ( .A(in[797]), .B(n4052), .Z(n2470) );
  NAND U3752 ( .A(n2198), .B(n2335), .Z(n2199) );
  XOR U3753 ( .A(n2470), .B(n2199), .Z(out[1416]) );
  XOR U3754 ( .A(in[798]), .B(n4056), .Z(n2337) );
  NAND U3755 ( .A(n2200), .B(n2338), .Z(n2201) );
  XNOR U3756 ( .A(n2337), .B(n2201), .Z(out[1417]) );
  XOR U3757 ( .A(in[799]), .B(n4060), .Z(n2340) );
  NAND U3758 ( .A(n2202), .B(n2341), .Z(n2203) );
  XNOR U3759 ( .A(n2340), .B(n2203), .Z(out[1418]) );
  XOR U3760 ( .A(in[800]), .B(n4064), .Z(n2343) );
  NAND U3761 ( .A(n2204), .B(n2344), .Z(n2205) );
  XNOR U3762 ( .A(n2343), .B(n2205), .Z(out[1419]) );
  XOR U3763 ( .A(in[678]), .B(n4290), .Z(n2888) );
  IV U3764 ( .A(n3043), .Z(n4134) );
  XOR U3765 ( .A(in[612]), .B(n4134), .Z(n4377) );
  NANDN U3766 ( .A(n4377), .B(n4374), .Z(n2206) );
  XNOR U3767 ( .A(n2888), .B(n2206), .Z(out[141]) );
  XOR U3768 ( .A(in[801]), .B(n4068), .Z(n2346) );
  NAND U3769 ( .A(n2207), .B(n2347), .Z(n2208) );
  XNOR U3770 ( .A(n2346), .B(n2208), .Z(out[1420]) );
  XOR U3771 ( .A(in[802]), .B(n4076), .Z(n2349) );
  NAND U3772 ( .A(n2209), .B(n2350), .Z(n2210) );
  XNOR U3773 ( .A(n2349), .B(n2210), .Z(out[1421]) );
  XOR U3774 ( .A(in[803]), .B(n4080), .Z(n2352) );
  NAND U3775 ( .A(n2211), .B(n2353), .Z(n2212) );
  XNOR U3776 ( .A(n2352), .B(n2212), .Z(out[1422]) );
  XOR U3777 ( .A(in[804]), .B(n4084), .Z(n2356) );
  NANDN U3778 ( .A(n2355), .B(n2213), .Z(n2214) );
  XNOR U3779 ( .A(n2356), .B(n2214), .Z(out[1423]) );
  IV U3780 ( .A(n2215), .Z(n4088) );
  XOR U3781 ( .A(in[805]), .B(n4088), .Z(n2500) );
  NANDN U3782 ( .A(n2357), .B(n2216), .Z(n2217) );
  XOR U3783 ( .A(n2500), .B(n2217), .Z(out[1424]) );
  XNOR U3784 ( .A(in[806]), .B(n4091), .Z(n2503) );
  NAND U3785 ( .A(n2218), .B(n2358), .Z(n2219) );
  XNOR U3786 ( .A(n2503), .B(n2219), .Z(out[1425]) );
  XNOR U3787 ( .A(in[807]), .B(n4095), .Z(n2507) );
  NAND U3788 ( .A(n2220), .B(n2361), .Z(n2221) );
  XNOR U3789 ( .A(n2507), .B(n2221), .Z(out[1426]) );
  XNOR U3790 ( .A(in[808]), .B(n4099), .Z(n2511) );
  NAND U3791 ( .A(n2222), .B(n2363), .Z(n2223) );
  XNOR U3792 ( .A(n2511), .B(n2223), .Z(out[1427]) );
  XNOR U3793 ( .A(in[809]), .B(n4103), .Z(n2515) );
  NAND U3794 ( .A(n2224), .B(n2365), .Z(n2225) );
  XNOR U3795 ( .A(n2515), .B(n2225), .Z(out[1428]) );
  XNOR U3796 ( .A(in[810]), .B(n4107), .Z(n2519) );
  NAND U3797 ( .A(n2226), .B(n2367), .Z(n2227) );
  XNOR U3798 ( .A(n2519), .B(n2227), .Z(out[1429]) );
  XOR U3799 ( .A(in[679]), .B(n4292), .Z(n2771) );
  XOR U3800 ( .A(in[613]), .B(n4138), .Z(n4410) );
  XNOR U3801 ( .A(in[204]), .B(n3956), .Z(n4407) );
  NANDN U3802 ( .A(n4410), .B(n4407), .Z(n2228) );
  XNOR U3803 ( .A(n2771), .B(n2228), .Z(out[142]) );
  XNOR U3804 ( .A(in[811]), .B(n4111), .Z(n2523) );
  NAND U3805 ( .A(n2229), .B(n2369), .Z(n2230) );
  XOR U3806 ( .A(n2523), .B(n2230), .Z(out[1430]) );
  XNOR U3807 ( .A(in[812]), .B(n4119), .Z(n2527) );
  NAND U3808 ( .A(n2231), .B(n2371), .Z(n2232) );
  XOR U3809 ( .A(n2527), .B(n2232), .Z(out[1431]) );
  XOR U3810 ( .A(in[813]), .B(n4123), .Z(n2532) );
  NAND U3811 ( .A(n2233), .B(n2373), .Z(n2234) );
  XOR U3812 ( .A(n2532), .B(n2234), .Z(out[1432]) );
  XOR U3813 ( .A(in[814]), .B(n4127), .Z(n2536) );
  NAND U3814 ( .A(n2235), .B(n2375), .Z(n2236) );
  XOR U3815 ( .A(n2536), .B(n2236), .Z(out[1433]) );
  XOR U3816 ( .A(in[815]), .B(n4131), .Z(n2540) );
  NAND U3817 ( .A(n2237), .B(n2377), .Z(n2238) );
  XOR U3818 ( .A(n2540), .B(n2238), .Z(out[1434]) );
  XOR U3819 ( .A(in[816]), .B(n4135), .Z(n2544) );
  NANDN U3820 ( .A(n2379), .B(n2239), .Z(n2240) );
  XOR U3821 ( .A(n2544), .B(n2240), .Z(out[1435]) );
  XOR U3822 ( .A(in[817]), .B(n4139), .Z(n2548) );
  NAND U3823 ( .A(n2241), .B(n2382), .Z(n2242) );
  XOR U3824 ( .A(n2548), .B(n2242), .Z(out[1436]) );
  XOR U3825 ( .A(in[818]), .B(n4143), .Z(n2552) );
  NAND U3826 ( .A(n2243), .B(n2384), .Z(n2244) );
  XOR U3827 ( .A(n2552), .B(n2244), .Z(out[1437]) );
  XOR U3828 ( .A(in[819]), .B(n4147), .Z(n2556) );
  NAND U3829 ( .A(n2245), .B(n2386), .Z(n2246) );
  XOR U3830 ( .A(n2556), .B(n2246), .Z(out[1438]) );
  XOR U3831 ( .A(in[820]), .B(n4151), .Z(n2560) );
  NAND U3832 ( .A(n2247), .B(n2388), .Z(n2248) );
  XOR U3833 ( .A(n2560), .B(n2248), .Z(out[1439]) );
  XOR U3834 ( .A(in[680]), .B(n4294), .Z(n2772) );
  XOR U3835 ( .A(in[614]), .B(n4142), .Z(n4444) );
  XNOR U3836 ( .A(in[205]), .B(n3960), .Z(n4441) );
  NANDN U3837 ( .A(n4444), .B(n4441), .Z(n2249) );
  XNOR U3838 ( .A(n2772), .B(n2249), .Z(out[143]) );
  XNOR U3839 ( .A(in[821]), .B(n4155), .Z(n2565) );
  NAND U3840 ( .A(n2250), .B(n2390), .Z(n2251) );
  XOR U3841 ( .A(n2565), .B(n2251), .Z(out[1440]) );
  XNOR U3842 ( .A(in[822]), .B(n4165), .Z(n2569) );
  NANDN U3843 ( .A(n2392), .B(n2252), .Z(n2253) );
  XOR U3844 ( .A(n2569), .B(n2253), .Z(out[1441]) );
  XNOR U3845 ( .A(in[823]), .B(n4169), .Z(n2575) );
  NANDN U3846 ( .A(n2393), .B(n2254), .Z(n2255) );
  XOR U3847 ( .A(n2575), .B(n2255), .Z(out[1442]) );
  XNOR U3848 ( .A(in[824]), .B(n4173), .Z(n2579) );
  NANDN U3849 ( .A(n2394), .B(n2256), .Z(n2257) );
  XOR U3850 ( .A(n2579), .B(n2257), .Z(out[1443]) );
  XNOR U3851 ( .A(in[825]), .B(n4177), .Z(n2583) );
  NANDN U3852 ( .A(n2395), .B(n2258), .Z(n2259) );
  XOR U3853 ( .A(n2583), .B(n2259), .Z(out[1444]) );
  XOR U3854 ( .A(in[826]), .B(n3901), .Z(n2587) );
  NANDN U3855 ( .A(n2396), .B(n2260), .Z(n2261) );
  XOR U3856 ( .A(n2587), .B(n2261), .Z(out[1445]) );
  XOR U3857 ( .A(in[827]), .B(n3905), .Z(n2591) );
  NANDN U3858 ( .A(n2398), .B(n2262), .Z(n2263) );
  XOR U3859 ( .A(n2591), .B(n2263), .Z(out[1446]) );
  XOR U3860 ( .A(in[828]), .B(n3909), .Z(n2595) );
  NANDN U3861 ( .A(n2399), .B(n2264), .Z(n2265) );
  XOR U3862 ( .A(n2595), .B(n2265), .Z(out[1447]) );
  XOR U3863 ( .A(in[829]), .B(n3913), .Z(n2599) );
  NANDN U3864 ( .A(n2400), .B(n2266), .Z(n2267) );
  XOR U3865 ( .A(n2599), .B(n2267), .Z(out[1448]) );
  XOR U3866 ( .A(in[830]), .B(n3917), .Z(n2603) );
  NANDN U3867 ( .A(n2401), .B(n2268), .Z(n2269) );
  XOR U3868 ( .A(n2603), .B(n2269), .Z(out[1449]) );
  XOR U3869 ( .A(in[681]), .B(n4296), .Z(n2773) );
  XOR U3870 ( .A(in[615]), .B(n4146), .Z(n4482) );
  XNOR U3871 ( .A(in[206]), .B(n3964), .Z(n4479) );
  NANDN U3872 ( .A(n4482), .B(n4479), .Z(n2270) );
  XNOR U3873 ( .A(n2773), .B(n2270), .Z(out[144]) );
  XOR U3874 ( .A(in[831]), .B(n3921), .Z(n2607) );
  NANDN U3875 ( .A(n2402), .B(n2271), .Z(n2272) );
  XOR U3876 ( .A(n2607), .B(n2272), .Z(out[1450]) );
  XOR U3877 ( .A(in[768]), .B(n3925), .Z(n2611) );
  NANDN U3878 ( .A(n2403), .B(n2273), .Z(n2274) );
  XOR U3879 ( .A(n2611), .B(n2274), .Z(out[1451]) );
  XOR U3880 ( .A(in[769]), .B(n3929), .Z(n2617) );
  NANDN U3881 ( .A(n2404), .B(n2275), .Z(n2276) );
  XOR U3882 ( .A(n2617), .B(n2276), .Z(out[1452]) );
  XNOR U3883 ( .A(n3934), .B(in[770]), .Z(n2621) );
  NANDN U3884 ( .A(n2405), .B(n2277), .Z(n2278) );
  XNOR U3885 ( .A(n2621), .B(n2278), .Z(out[1453]) );
  IV U3886 ( .A(n3177), .Z(n3938) );
  XOR U3887 ( .A(n3938), .B(in[771]), .Z(n2625) );
  NANDN U3888 ( .A(n2406), .B(n2279), .Z(n2280) );
  XOR U3889 ( .A(n2625), .B(n2280), .Z(out[1454]) );
  IV U3890 ( .A(n3179), .Z(n3945) );
  XOR U3891 ( .A(n3945), .B(in[772]), .Z(n2629) );
  NANDN U3892 ( .A(n2407), .B(n2281), .Z(n2282) );
  XOR U3893 ( .A(n2629), .B(n2282), .Z(out[1455]) );
  IV U3894 ( .A(n3181), .Z(n3949) );
  XOR U3895 ( .A(n3949), .B(in[773]), .Z(n2633) );
  NANDN U3896 ( .A(n2409), .B(n2283), .Z(n2284) );
  XOR U3897 ( .A(n2633), .B(n2284), .Z(out[1456]) );
  IV U3898 ( .A(n3183), .Z(n3953) );
  XOR U3899 ( .A(n3953), .B(in[774]), .Z(n2637) );
  NANDN U3900 ( .A(n2410), .B(n2285), .Z(n2286) );
  XOR U3901 ( .A(n2637), .B(n2286), .Z(out[1457]) );
  IV U3902 ( .A(n3185), .Z(n3957) );
  XOR U3903 ( .A(n3957), .B(in[775]), .Z(n2641) );
  NANDN U3904 ( .A(n2411), .B(n2287), .Z(n2288) );
  XOR U3905 ( .A(n2641), .B(n2288), .Z(out[1458]) );
  IV U3906 ( .A(n3187), .Z(n3961) );
  XOR U3907 ( .A(n3961), .B(in[776]), .Z(n2645) );
  NAND U3908 ( .A(n2289), .B(n2412), .Z(n2290) );
  XOR U3909 ( .A(n2645), .B(n2290), .Z(out[1459]) );
  XOR U3910 ( .A(in[682]), .B(n4298), .Z(n2774) );
  XOR U3911 ( .A(in[616]), .B(n4150), .Z(n4516) );
  XNOR U3912 ( .A(in[207]), .B(n3968), .Z(n4513) );
  NANDN U3913 ( .A(n4516), .B(n4513), .Z(n2291) );
  XNOR U3914 ( .A(n2774), .B(n2291), .Z(out[145]) );
  IV U3915 ( .A(n3189), .Z(n3965) );
  XOR U3916 ( .A(in[777]), .B(n3965), .Z(n2649) );
  NAND U3917 ( .A(n2292), .B(n2414), .Z(n2293) );
  XOR U3918 ( .A(n2649), .B(n2293), .Z(out[1460]) );
  IV U3919 ( .A(n3191), .Z(n3969) );
  XOR U3920 ( .A(n3969), .B(in[778]), .Z(n2653) );
  NAND U3921 ( .A(n2294), .B(n2416), .Z(n2295) );
  XOR U3922 ( .A(n2653), .B(n2295), .Z(out[1461]) );
  IV U3923 ( .A(n2296), .Z(n3973) );
  XOR U3924 ( .A(n3973), .B(in[779]), .Z(n2659) );
  NANDN U3925 ( .A(n2418), .B(n2297), .Z(n2298) );
  XOR U3926 ( .A(n2659), .B(n2298), .Z(out[1462]) );
  IV U3927 ( .A(n3198), .Z(n3977) );
  XOR U3928 ( .A(in[780]), .B(n3977), .Z(n2663) );
  NANDN U3929 ( .A(n2419), .B(n2299), .Z(n2300) );
  XOR U3930 ( .A(n2663), .B(n2300), .Z(out[1463]) );
  IV U3931 ( .A(n3200), .Z(n3981) );
  XOR U3932 ( .A(in[781]), .B(n3981), .Z(n2667) );
  NANDN U3933 ( .A(n2420), .B(n2301), .Z(n2302) );
  XOR U3934 ( .A(n2667), .B(n2302), .Z(out[1464]) );
  IV U3935 ( .A(n3203), .Z(n3988) );
  XOR U3936 ( .A(in[782]), .B(n3988), .Z(n2671) );
  NAND U3937 ( .A(n2303), .B(n2421), .Z(n2304) );
  XOR U3938 ( .A(n2671), .B(n2304), .Z(out[1465]) );
  IV U3939 ( .A(n3206), .Z(n3992) );
  XOR U3940 ( .A(in[783]), .B(n3992), .Z(n2675) );
  NAND U3941 ( .A(n2305), .B(n2424), .Z(n2306) );
  XOR U3942 ( .A(n2675), .B(n2306), .Z(out[1466]) );
  IV U3943 ( .A(n3209), .Z(n3996) );
  XOR U3944 ( .A(in[784]), .B(n3996), .Z(n2679) );
  NAND U3945 ( .A(n2307), .B(n2426), .Z(n2308) );
  XOR U3946 ( .A(n2679), .B(n2308), .Z(out[1467]) );
  IV U3947 ( .A(n3212), .Z(n4000) );
  XOR U3948 ( .A(in[785]), .B(n4000), .Z(n2683) );
  NAND U3949 ( .A(n2309), .B(n2428), .Z(n2310) );
  XOR U3950 ( .A(n2683), .B(n2310), .Z(out[1468]) );
  XOR U3951 ( .A(in[786]), .B(n4004), .Z(n2430) );
  NAND U3952 ( .A(n2311), .B(n2431), .Z(n2312) );
  XNOR U3953 ( .A(n2430), .B(n2312), .Z(out[1469]) );
  XOR U3954 ( .A(in[683]), .B(n4300), .Z(n2778) );
  XOR U3955 ( .A(in[617]), .B(n4154), .Z(n4555) );
  XNOR U3956 ( .A(in[208]), .B(n3972), .Z(n4552) );
  NANDN U3957 ( .A(n4555), .B(n4552), .Z(n2313) );
  XNOR U3958 ( .A(n2778), .B(n2313), .Z(out[146]) );
  XOR U3959 ( .A(in[787]), .B(n4008), .Z(n2691) );
  NAND U3960 ( .A(n2314), .B(n2433), .Z(n2315) );
  XOR U3961 ( .A(n2691), .B(n2315), .Z(out[1470]) );
  XOR U3962 ( .A(in[788]), .B(n4012), .Z(n2695) );
  NAND U3963 ( .A(n2316), .B(n2435), .Z(n2317) );
  XOR U3964 ( .A(n2695), .B(n2317), .Z(out[1471]) );
  NANDN U3965 ( .A(n2318), .B(n2437), .Z(n2319) );
  XOR U3966 ( .A(n2438), .B(n2319), .Z(out[1472]) );
  NANDN U3967 ( .A(n2320), .B(n2440), .Z(n2321) );
  XOR U3968 ( .A(n2441), .B(n2321), .Z(out[1473]) );
  NANDN U3969 ( .A(n2322), .B(n2443), .Z(n2323) );
  XOR U3970 ( .A(n2444), .B(n2323), .Z(out[1474]) );
  NANDN U3971 ( .A(n2324), .B(n2447), .Z(n2325) );
  XOR U3972 ( .A(n2448), .B(n2325), .Z(out[1475]) );
  NANDN U3973 ( .A(n2326), .B(n2453), .Z(n2327) );
  XOR U3974 ( .A(n2454), .B(n2327), .Z(out[1476]) );
  NANDN U3975 ( .A(n2328), .B(n2457), .Z(n2329) );
  XOR U3976 ( .A(n2458), .B(n2329), .Z(out[1477]) );
  NANDN U3977 ( .A(n2330), .B(n2461), .Z(n2331) );
  XOR U3978 ( .A(n2462), .B(n2331), .Z(out[1478]) );
  NANDN U3979 ( .A(n2332), .B(n2465), .Z(n2333) );
  XOR U3980 ( .A(n2466), .B(n2333), .Z(out[1479]) );
  XNOR U3981 ( .A(in[684]), .B(n4302), .Z(n2909) );
  XOR U3982 ( .A(in[618]), .B(n4164), .Z(n4584) );
  XNOR U3983 ( .A(in[209]), .B(n3976), .Z(n4581) );
  NANDN U3984 ( .A(n4584), .B(n4581), .Z(n2334) );
  XOR U3985 ( .A(n2909), .B(n2334), .Z(out[147]) );
  NANDN U3986 ( .A(n2335), .B(n2470), .Z(n2336) );
  XOR U3987 ( .A(n2471), .B(n2336), .Z(out[1480]) );
  IV U3988 ( .A(n2337), .Z(n2473) );
  NANDN U3989 ( .A(n2338), .B(n2473), .Z(n2339) );
  XOR U3990 ( .A(n2474), .B(n2339), .Z(out[1481]) );
  IV U3991 ( .A(n2340), .Z(n2476) );
  NANDN U3992 ( .A(n2341), .B(n2476), .Z(n2342) );
  XOR U3993 ( .A(n2477), .B(n2342), .Z(out[1482]) );
  IV U3994 ( .A(n2343), .Z(n2478) );
  NANDN U3995 ( .A(n2344), .B(n2478), .Z(n2345) );
  XOR U3996 ( .A(n2479), .B(n2345), .Z(out[1483]) );
  IV U3997 ( .A(n2346), .Z(n2482) );
  NANDN U3998 ( .A(n2347), .B(n2482), .Z(n2348) );
  XOR U3999 ( .A(n2483), .B(n2348), .Z(out[1484]) );
  IV U4000 ( .A(n2349), .Z(n2487) );
  NANDN U4001 ( .A(n2350), .B(n2487), .Z(n2351) );
  XOR U4002 ( .A(n2488), .B(n2351), .Z(out[1485]) );
  IV U4003 ( .A(n2352), .Z(n2491) );
  NANDN U4004 ( .A(n2353), .B(n2491), .Z(n2354) );
  XNOR U4005 ( .A(n2490), .B(n2354), .Z(out[1486]) );
  IV U4006 ( .A(n2356), .Z(n2495) );
  OR U4007 ( .A(n2503), .B(n2358), .Z(n2359) );
  XOR U4008 ( .A(n2504), .B(n2359), .Z(out[1489]) );
  XNOR U4009 ( .A(in[685]), .B(n4304), .Z(n2912) );
  XOR U4010 ( .A(in[619]), .B(n4168), .Z(n4609) );
  XNOR U4011 ( .A(in[210]), .B(n3980), .Z(n4606) );
  NANDN U4012 ( .A(n4609), .B(n4606), .Z(n2360) );
  XOR U4013 ( .A(n2912), .B(n2360), .Z(out[148]) );
  OR U4014 ( .A(n2507), .B(n2361), .Z(n2362) );
  XOR U4015 ( .A(n2508), .B(n2362), .Z(out[1490]) );
  OR U4016 ( .A(n2511), .B(n2363), .Z(n2364) );
  XOR U4017 ( .A(n2512), .B(n2364), .Z(out[1491]) );
  OR U4018 ( .A(n2515), .B(n2365), .Z(n2366) );
  XOR U4019 ( .A(n2516), .B(n2366), .Z(out[1492]) );
  OR U4020 ( .A(n2519), .B(n2367), .Z(n2368) );
  XOR U4021 ( .A(n2520), .B(n2368), .Z(out[1493]) );
  NANDN U4022 ( .A(n2369), .B(n2523), .Z(n2370) );
  XOR U4023 ( .A(n2524), .B(n2370), .Z(out[1494]) );
  NANDN U4024 ( .A(n2371), .B(n2527), .Z(n2372) );
  XNOR U4025 ( .A(n2528), .B(n2372), .Z(out[1495]) );
  NANDN U4026 ( .A(n2373), .B(n2532), .Z(n2374) );
  XNOR U4027 ( .A(n2533), .B(n2374), .Z(out[1496]) );
  NANDN U4028 ( .A(n2375), .B(n2536), .Z(n2376) );
  XNOR U4029 ( .A(n2537), .B(n2376), .Z(out[1497]) );
  NANDN U4030 ( .A(n2377), .B(n2540), .Z(n2378) );
  XNOR U4031 ( .A(n2541), .B(n2378), .Z(out[1498]) );
  XOR U4032 ( .A(in[686]), .B(n4306), .Z(n2915) );
  XOR U4033 ( .A(in[620]), .B(n4172), .Z(n4638) );
  XOR U4034 ( .A(in[211]), .B(n3987), .Z(n4635) );
  NANDN U4035 ( .A(n4638), .B(n4635), .Z(n2380) );
  XNOR U4036 ( .A(n2915), .B(n2380), .Z(out[149]) );
  XOR U4037 ( .A(in[1424]), .B(n3209), .Z(n4408) );
  XNOR U4038 ( .A(in[1047]), .B(n4501), .Z(n2893) );
  NANDN U4039 ( .A(n4408), .B(n2893), .Z(n2381) );
  XNOR U4040 ( .A(n4407), .B(n2381), .Z(out[14]) );
  NANDN U4041 ( .A(n2382), .B(n2548), .Z(n2383) );
  XNOR U4042 ( .A(n2549), .B(n2383), .Z(out[1500]) );
  NANDN U4043 ( .A(n2384), .B(n2552), .Z(n2385) );
  XNOR U4044 ( .A(n2553), .B(n2385), .Z(out[1501]) );
  NANDN U4045 ( .A(n2386), .B(n2556), .Z(n2387) );
  XNOR U4046 ( .A(n2557), .B(n2387), .Z(out[1502]) );
  NANDN U4047 ( .A(n2388), .B(n2560), .Z(n2389) );
  XNOR U4048 ( .A(n2561), .B(n2389), .Z(out[1503]) );
  NANDN U4049 ( .A(n2390), .B(n2565), .Z(n2391) );
  XNOR U4050 ( .A(n2566), .B(n2391), .Z(out[1504]) );
  XOR U4051 ( .A(in[687]), .B(n4308), .Z(n2918) );
  XOR U4052 ( .A(in[621]), .B(n4176), .Z(n4668) );
  XOR U4053 ( .A(in[212]), .B(n3991), .Z(n4665) );
  NANDN U4054 ( .A(n4668), .B(n4665), .Z(n2397) );
  XNOR U4055 ( .A(n2918), .B(n2397), .Z(out[150]) );
  XOR U4056 ( .A(in[688]), .B(n4315), .Z(n2921) );
  XOR U4057 ( .A(in[622]), .B(n3900), .Z(n4683) );
  XOR U4058 ( .A(in[213]), .B(n3995), .Z(n4680) );
  NANDN U4059 ( .A(n4683), .B(n4680), .Z(n2408) );
  XNOR U4060 ( .A(n2921), .B(n2408), .Z(out[151]) );
  NANDN U4061 ( .A(n2412), .B(n2645), .Z(n2413) );
  XOR U4062 ( .A(n2646), .B(n2413), .Z(out[1523]) );
  NANDN U4063 ( .A(n2414), .B(n2649), .Z(n2415) );
  XOR U4064 ( .A(n2650), .B(n2415), .Z(out[1524]) );
  NANDN U4065 ( .A(n2416), .B(n2653), .Z(n2417) );
  XOR U4066 ( .A(n2654), .B(n2417), .Z(out[1525]) );
  NANDN U4067 ( .A(n2421), .B(n2671), .Z(n2422) );
  XOR U4068 ( .A(n2672), .B(n2422), .Z(out[1529]) );
  XOR U4069 ( .A(in[689]), .B(n4318), .Z(n2927) );
  XOR U4070 ( .A(in[214]), .B(n3999), .Z(n4697) );
  XNOR U4071 ( .A(in[623]), .B(n3904), .Z(n4699) );
  NANDN U4072 ( .A(n4697), .B(n4699), .Z(n2423) );
  XNOR U4073 ( .A(n2927), .B(n2423), .Z(out[152]) );
  NANDN U4074 ( .A(n2424), .B(n2675), .Z(n2425) );
  XOR U4075 ( .A(n2676), .B(n2425), .Z(out[1530]) );
  NANDN U4076 ( .A(n2426), .B(n2679), .Z(n2427) );
  XOR U4077 ( .A(n2680), .B(n2427), .Z(out[1531]) );
  NANDN U4078 ( .A(n2428), .B(n2683), .Z(n2429) );
  XOR U4079 ( .A(n2684), .B(n2429), .Z(out[1532]) );
  IV U4080 ( .A(n2430), .Z(n2687) );
  NANDN U4081 ( .A(n2431), .B(n2687), .Z(n2432) );
  XOR U4082 ( .A(n2688), .B(n2432), .Z(out[1533]) );
  NANDN U4083 ( .A(n2433), .B(n2691), .Z(n2434) );
  XOR U4084 ( .A(n2692), .B(n2434), .Z(out[1534]) );
  NANDN U4085 ( .A(n2435), .B(n2695), .Z(n2436) );
  XOR U4086 ( .A(n2696), .B(n2436), .Z(out[1535]) );
  ANDN U4087 ( .B(n2444), .A(n2443), .Z(n2445) );
  XOR U4088 ( .A(n2446), .B(n2445), .Z(out[1538]) );
  ANDN U4089 ( .B(n2448), .A(n2447), .Z(n2451) );
  XOR U4090 ( .A(n2449), .B(round_const_3), .Z(n2450) );
  XNOR U4091 ( .A(n2451), .B(n2450), .Z(out[1539]) );
  XOR U4092 ( .A(in[690]), .B(n4321), .Z(n2930) );
  XOR U4093 ( .A(in[624]), .B(n3908), .Z(n4734) );
  XOR U4094 ( .A(in[215]), .B(n4003), .Z(n4731) );
  NANDN U4095 ( .A(n4734), .B(n4731), .Z(n2452) );
  XNOR U4096 ( .A(n2930), .B(n2452), .Z(out[153]) );
  ANDN U4097 ( .B(n2454), .A(n2453), .Z(n2455) );
  XOR U4098 ( .A(n2456), .B(n2455), .Z(out[1540]) );
  ANDN U4099 ( .B(n2458), .A(n2457), .Z(n2459) );
  XOR U4100 ( .A(n2460), .B(n2459), .Z(out[1541]) );
  ANDN U4101 ( .B(n2462), .A(n2461), .Z(n2463) );
  XOR U4102 ( .A(n2464), .B(n2463), .Z(out[1542]) );
  ANDN U4103 ( .B(n2466), .A(n2465), .Z(n2467) );
  XOR U4104 ( .A(n2468), .B(n2467), .Z(out[1543]) );
  ANDN U4105 ( .B(n2479), .A(n2478), .Z(n2480) );
  XNOR U4106 ( .A(n2481), .B(n2480), .Z(out[1547]) );
  ANDN U4107 ( .B(n2483), .A(n2482), .Z(n2484) );
  XNOR U4108 ( .A(n2485), .B(n2484), .Z(out[1548]) );
  XOR U4109 ( .A(in[691]), .B(n4324), .Z(n2933) );
  XOR U4110 ( .A(in[216]), .B(n4007), .Z(n4779) );
  XNOR U4111 ( .A(in[625]), .B(n3912), .Z(n4781) );
  NANDN U4112 ( .A(n4779), .B(n4781), .Z(n2489) );
  XNOR U4113 ( .A(n2933), .B(n2489), .Z(out[154]) );
  NOR U4114 ( .A(n2491), .B(n2490), .Z(n2492) );
  XOR U4115 ( .A(n2493), .B(n2492), .Z(out[1550]) );
  NOR U4116 ( .A(n2495), .B(n2494), .Z(n2498) );
  XNOR U4117 ( .A(n2496), .B(round_const_15), .Z(n2497) );
  XNOR U4118 ( .A(n2498), .B(n2497), .Z(out[1551]) );
  NOR U4119 ( .A(n2500), .B(n2499), .Z(n2501) );
  XOR U4120 ( .A(n2502), .B(n2501), .Z(out[1552]) );
  AND U4121 ( .A(n2504), .B(n2503), .Z(n2505) );
  XOR U4122 ( .A(n2506), .B(n2505), .Z(out[1553]) );
  AND U4123 ( .A(n2508), .B(n2507), .Z(n2509) );
  XOR U4124 ( .A(n2510), .B(n2509), .Z(out[1554]) );
  AND U4125 ( .A(n2512), .B(n2511), .Z(n2513) );
  XOR U4126 ( .A(n2514), .B(n2513), .Z(out[1555]) );
  AND U4127 ( .A(n2516), .B(n2515), .Z(n2517) );
  XOR U4128 ( .A(n2518), .B(n2517), .Z(out[1556]) );
  AND U4129 ( .A(n2520), .B(n2519), .Z(n2521) );
  XOR U4130 ( .A(n2522), .B(n2521), .Z(out[1557]) );
  ANDN U4131 ( .B(n2524), .A(n2523), .Z(n2525) );
  XOR U4132 ( .A(n2526), .B(n2525), .Z(out[1558]) );
  NOR U4133 ( .A(n2528), .B(n2527), .Z(n2529) );
  XOR U4134 ( .A(n2530), .B(n2529), .Z(out[1559]) );
  XOR U4135 ( .A(in[692]), .B(n4327), .Z(n2936) );
  XOR U4136 ( .A(in[217]), .B(n4011), .Z(n4822) );
  XNOR U4137 ( .A(in[626]), .B(n3916), .Z(n4824) );
  NANDN U4138 ( .A(n4822), .B(n4824), .Z(n2531) );
  XNOR U4139 ( .A(n2936), .B(n2531), .Z(out[155]) );
  NOR U4140 ( .A(n2533), .B(n2532), .Z(n2534) );
  XOR U4141 ( .A(n2535), .B(n2534), .Z(out[1560]) );
  NOR U4142 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U4143 ( .A(n2539), .B(n2538), .Z(out[1561]) );
  NOR U4144 ( .A(n2541), .B(n2540), .Z(n2542) );
  XOR U4145 ( .A(n2543), .B(n2542), .Z(out[1562]) );
  NOR U4146 ( .A(n2545), .B(n2544), .Z(n2546) );
  XOR U4147 ( .A(n2547), .B(n2546), .Z(out[1563]) );
  NOR U4148 ( .A(n2549), .B(n2548), .Z(n2550) );
  XOR U4149 ( .A(n2551), .B(n2550), .Z(out[1564]) );
  NOR U4150 ( .A(n2553), .B(n2552), .Z(n2554) );
  XOR U4151 ( .A(n2555), .B(n2554), .Z(out[1565]) );
  NOR U4152 ( .A(n2557), .B(n2556), .Z(n2558) );
  XOR U4153 ( .A(n2559), .B(n2558), .Z(out[1566]) );
  NOR U4154 ( .A(n2561), .B(n2560), .Z(n2564) );
  XNOR U4155 ( .A(n2562), .B(round_const_31), .Z(n2563) );
  XNOR U4156 ( .A(n2564), .B(n2563), .Z(out[1567]) );
  NOR U4157 ( .A(n2566), .B(n2565), .Z(n2567) );
  XOR U4158 ( .A(n2568), .B(n2567), .Z(out[1568]) );
  NOR U4159 ( .A(n2570), .B(n2569), .Z(n2571) );
  XOR U4160 ( .A(n2572), .B(n2571), .Z(out[1569]) );
  XOR U4161 ( .A(in[693]), .B(n4330), .Z(n2938) );
  XOR U4162 ( .A(in[218]), .B(n4015), .Z(n4866) );
  XNOR U4163 ( .A(in[627]), .B(n2573), .Z(n4868) );
  NANDN U4164 ( .A(n4866), .B(n4868), .Z(n2574) );
  XNOR U4165 ( .A(n2938), .B(n2574), .Z(out[156]) );
  NOR U4166 ( .A(n2576), .B(n2575), .Z(n2577) );
  XOR U4167 ( .A(n2578), .B(n2577), .Z(out[1570]) );
  NOR U4168 ( .A(n2580), .B(n2579), .Z(n2581) );
  XOR U4169 ( .A(n2582), .B(n2581), .Z(out[1571]) );
  NOR U4170 ( .A(n2584), .B(n2583), .Z(n2585) );
  XOR U4171 ( .A(n2586), .B(n2585), .Z(out[1572]) );
  NOR U4172 ( .A(n2588), .B(n2587), .Z(n2589) );
  XOR U4173 ( .A(n2590), .B(n2589), .Z(out[1573]) );
  NOR U4174 ( .A(n2592), .B(n2591), .Z(n2593) );
  XNOR U4175 ( .A(n2594), .B(n2593), .Z(out[1574]) );
  ANDN U4176 ( .B(n2596), .A(n2595), .Z(n2597) );
  XOR U4177 ( .A(n2598), .B(n2597), .Z(out[1575]) );
  ANDN U4178 ( .B(n2600), .A(n2599), .Z(n2601) );
  XOR U4179 ( .A(n2602), .B(n2601), .Z(out[1576]) );
  ANDN U4180 ( .B(n2604), .A(n2603), .Z(n2605) );
  XOR U4181 ( .A(n2606), .B(n2605), .Z(out[1577]) );
  NOR U4182 ( .A(n2608), .B(n2607), .Z(n2609) );
  XOR U4183 ( .A(n2610), .B(n2609), .Z(out[1578]) );
  ANDN U4184 ( .B(n2612), .A(n2611), .Z(n2613) );
  XOR U4185 ( .A(n2614), .B(n2613), .Z(out[1579]) );
  XOR U4186 ( .A(in[694]), .B(n4333), .Z(n2940) );
  XOR U4187 ( .A(in[219]), .B(n4019), .Z(n4910) );
  XNOR U4188 ( .A(in[628]), .B(n2615), .Z(n4912) );
  NANDN U4189 ( .A(n4910), .B(n4912), .Z(n2616) );
  XNOR U4190 ( .A(n2940), .B(n2616), .Z(out[157]) );
  ANDN U4191 ( .B(n2618), .A(n2617), .Z(n2619) );
  XOR U4192 ( .A(n2620), .B(n2619), .Z(out[1580]) );
  AND U4193 ( .A(n2622), .B(n2621), .Z(n2623) );
  XOR U4194 ( .A(n2624), .B(n2623), .Z(out[1581]) );
  ANDN U4195 ( .B(n2626), .A(n2625), .Z(n2627) );
  XOR U4196 ( .A(n2628), .B(n2627), .Z(out[1582]) );
  ANDN U4197 ( .B(n2630), .A(n2629), .Z(n2631) );
  XOR U4198 ( .A(n2632), .B(n2631), .Z(out[1583]) );
  ANDN U4199 ( .B(n2634), .A(n2633), .Z(n2635) );
  XOR U4200 ( .A(n2636), .B(n2635), .Z(out[1584]) );
  ANDN U4201 ( .B(n2638), .A(n2637), .Z(n2639) );
  XOR U4202 ( .A(n2640), .B(n2639), .Z(out[1585]) );
  ANDN U4203 ( .B(n2642), .A(n2641), .Z(n2643) );
  XOR U4204 ( .A(n2644), .B(n2643), .Z(out[1586]) );
  ANDN U4205 ( .B(n2646), .A(n2645), .Z(n2647) );
  XOR U4206 ( .A(n2648), .B(n2647), .Z(out[1587]) );
  ANDN U4207 ( .B(n2650), .A(n2649), .Z(n2651) );
  XOR U4208 ( .A(n2652), .B(n2651), .Z(out[1588]) );
  ANDN U4209 ( .B(n2654), .A(n2653), .Z(n2655) );
  XOR U4210 ( .A(n2656), .B(n2655), .Z(out[1589]) );
  XOR U4211 ( .A(in[695]), .B(n4336), .Z(n2942) );
  XNOR U4212 ( .A(in[220]), .B(n4023), .Z(n4954) );
  XNOR U4213 ( .A(in[629]), .B(n2657), .Z(n4956) );
  NANDN U4214 ( .A(n4954), .B(n4956), .Z(n2658) );
  XNOR U4215 ( .A(n2942), .B(n2658), .Z(out[158]) );
  ANDN U4216 ( .B(n2660), .A(n2659), .Z(n2661) );
  XNOR U4217 ( .A(n2662), .B(n2661), .Z(out[1590]) );
  ANDN U4218 ( .B(n2664), .A(n2663), .Z(n2665) );
  XNOR U4219 ( .A(n2666), .B(n2665), .Z(out[1591]) );
  ANDN U4220 ( .B(n2668), .A(n2667), .Z(n2669) );
  XNOR U4221 ( .A(n2670), .B(n2669), .Z(out[1592]) );
  ANDN U4222 ( .B(n2672), .A(n2671), .Z(n2673) );
  XOR U4223 ( .A(n2674), .B(n2673), .Z(out[1593]) );
  ANDN U4224 ( .B(n2676), .A(n2675), .Z(n2677) );
  XOR U4225 ( .A(n2678), .B(n2677), .Z(out[1594]) );
  ANDN U4226 ( .B(n2680), .A(n2679), .Z(n2681) );
  XOR U4227 ( .A(n2682), .B(n2681), .Z(out[1595]) );
  ANDN U4228 ( .B(n2684), .A(n2683), .Z(n2685) );
  XOR U4229 ( .A(n2686), .B(n2685), .Z(out[1596]) );
  ANDN U4230 ( .B(n2688), .A(n2687), .Z(n2689) );
  XOR U4231 ( .A(n2690), .B(n2689), .Z(out[1597]) );
  ANDN U4232 ( .B(n2692), .A(n2691), .Z(n2693) );
  XOR U4233 ( .A(n2694), .B(n2693), .Z(out[1598]) );
  XOR U4234 ( .A(in[696]), .B(n4180), .Z(n2944) );
  XNOR U4235 ( .A(in[221]), .B(n4031), .Z(n4998) );
  XNOR U4236 ( .A(in[630]), .B(n3069), .Z(n5000) );
  NANDN U4237 ( .A(n4998), .B(n5000), .Z(n2698) );
  XNOR U4238 ( .A(n2944), .B(n2698), .Z(out[159]) );
  XOR U4239 ( .A(in[1425]), .B(n3212), .Z(n4442) );
  XNOR U4240 ( .A(in[1048]), .B(n4504), .Z(n2896) );
  NANDN U4241 ( .A(n4442), .B(n2896), .Z(n2699) );
  XNOR U4242 ( .A(n4441), .B(n2699), .Z(out[15]) );
  XOR U4243 ( .A(in[697]), .B(n4183), .Z(n2946) );
  XNOR U4244 ( .A(in[222]), .B(n4035), .Z(n5042) );
  XNOR U4245 ( .A(in[631]), .B(n3071), .Z(n5044) );
  NANDN U4246 ( .A(n5042), .B(n5044), .Z(n2700) );
  XNOR U4247 ( .A(n2946), .B(n2700), .Z(out[160]) );
  XOR U4248 ( .A(in[698]), .B(n4186), .Z(n2948) );
  XNOR U4249 ( .A(in[223]), .B(n4039), .Z(n5083) );
  XNOR U4250 ( .A(in[632]), .B(n3074), .Z(n5085) );
  NANDN U4251 ( .A(n5083), .B(n5085), .Z(n2701) );
  XNOR U4252 ( .A(n2948), .B(n2701), .Z(out[161]) );
  XOR U4253 ( .A(in[699]), .B(n4189), .Z(n2952) );
  XNOR U4254 ( .A(in[633]), .B(n2702), .Z(n5120) );
  XOR U4255 ( .A(in[224]), .B(n4043), .Z(n5117) );
  NAND U4256 ( .A(n5120), .B(n5117), .Z(n2703) );
  XNOR U4257 ( .A(n2952), .B(n2703), .Z(out[162]) );
  XOR U4258 ( .A(in[700]), .B(n4192), .Z(n2954) );
  XNOR U4259 ( .A(in[634]), .B(n2704), .Z(n5163) );
  XOR U4260 ( .A(in[225]), .B(n4047), .Z(n5160) );
  NAND U4261 ( .A(n5163), .B(n5160), .Z(n2705) );
  XOR U4262 ( .A(n2954), .B(n2705), .Z(out[163]) );
  XOR U4263 ( .A(in[701]), .B(n4195), .Z(n2956) );
  ANDN U4264 ( .B(n3117), .A(n2706), .Z(n2707) );
  XNOR U4265 ( .A(n2956), .B(n2707), .Z(out[164]) );
  XOR U4266 ( .A(in[702]), .B(n4200), .Z(n2958) );
  ANDN U4267 ( .B(n3141), .A(n2708), .Z(n2709) );
  XNOR U4268 ( .A(n2958), .B(n2709), .Z(out[165]) );
  XNOR U4269 ( .A(in[703]), .B(n4201), .Z(n2960) );
  ANDN U4270 ( .B(n3160), .A(n2710), .Z(n2711) );
  XNOR U4271 ( .A(n2960), .B(n2711), .Z(out[166]) );
  XOR U4272 ( .A(in[640]), .B(n4202), .Z(n2962) );
  ANDN U4273 ( .B(n3171), .A(n2712), .Z(n2713) );
  XNOR U4274 ( .A(n2962), .B(n2713), .Z(out[167]) );
  XOR U4275 ( .A(in[641]), .B(n4203), .Z(n2964) );
  NOR U4276 ( .A(n2714), .B(n3196), .Z(n2715) );
  XNOR U4277 ( .A(n2964), .B(n2715), .Z(out[168]) );
  XOR U4278 ( .A(in[642]), .B(n4204), .Z(n2966) );
  NOR U4279 ( .A(n2716), .B(n3226), .Z(n2717) );
  XNOR U4280 ( .A(n2966), .B(n2717), .Z(out[169]) );
  XOR U4281 ( .A(in[1426]), .B(n4004), .Z(n4480) );
  XNOR U4282 ( .A(in[1049]), .B(n4507), .Z(n2899) );
  NANDN U4283 ( .A(n4480), .B(n2899), .Z(n2718) );
  XNOR U4284 ( .A(n4479), .B(n2718), .Z(out[16]) );
  XOR U4285 ( .A(in[643]), .B(n4205), .Z(n2968) );
  NOR U4286 ( .A(n2719), .B(n3250), .Z(n2720) );
  XNOR U4287 ( .A(n2968), .B(n2720), .Z(out[170]) );
  XOR U4288 ( .A(in[644]), .B(n4206), .Z(n2970) );
  NOR U4289 ( .A(n2721), .B(n3262), .Z(n2722) );
  XNOR U4290 ( .A(n2970), .B(n2722), .Z(out[171]) );
  XOR U4291 ( .A(in[645]), .B(n4207), .Z(n2976) );
  NOR U4292 ( .A(n2723), .B(n3272), .Z(n2724) );
  XNOR U4293 ( .A(n2976), .B(n2724), .Z(out[172]) );
  XOR U4294 ( .A(in[646]), .B(n4210), .Z(n2978) );
  NOR U4295 ( .A(n3306), .B(n2813), .Z(n2725) );
  XNOR U4296 ( .A(n2978), .B(n2725), .Z(out[173]) );
  XOR U4297 ( .A(in[647]), .B(n4213), .Z(n2980) );
  NOR U4298 ( .A(n3336), .B(n2815), .Z(n2726) );
  XNOR U4299 ( .A(n2980), .B(n2726), .Z(out[174]) );
  XNOR U4300 ( .A(in[648]), .B(n4218), .Z(n2982) );
  NOR U4301 ( .A(n3364), .B(n2817), .Z(n2727) );
  XNOR U4302 ( .A(n2982), .B(n2727), .Z(out[175]) );
  XOR U4303 ( .A(in[649]), .B(n4221), .Z(n2984) );
  NOR U4304 ( .A(n3392), .B(n2822), .Z(n2728) );
  XNOR U4305 ( .A(n2984), .B(n2728), .Z(out[176]) );
  XOR U4306 ( .A(in[650]), .B(n4224), .Z(n2986) );
  NOR U4307 ( .A(n3427), .B(n2824), .Z(n2729) );
  XNOR U4308 ( .A(n2986), .B(n2729), .Z(out[177]) );
  IV U4309 ( .A(n3096), .Z(n4227) );
  XOR U4310 ( .A(in[651]), .B(n4227), .Z(n2988) );
  NOR U4311 ( .A(n3462), .B(n2826), .Z(n2730) );
  XNOR U4312 ( .A(n2988), .B(n2730), .Z(out[178]) );
  IV U4313 ( .A(n3098), .Z(n4230) );
  XOR U4314 ( .A(in[652]), .B(n4230), .Z(n2990) );
  NOR U4315 ( .A(n3484), .B(n2828), .Z(n2731) );
  XNOR U4316 ( .A(n2990), .B(n2731), .Z(out[179]) );
  XOR U4317 ( .A(in[1427]), .B(n3217), .Z(n4514) );
  XNOR U4318 ( .A(in[1050]), .B(n4510), .Z(n2902) );
  NANDN U4319 ( .A(n4514), .B(n2902), .Z(n2732) );
  XNOR U4320 ( .A(n4513), .B(n2732), .Z(out[17]) );
  IV U4321 ( .A(n3102), .Z(n4233) );
  XOR U4322 ( .A(in[653]), .B(n4233), .Z(n2992) );
  NOR U4323 ( .A(n3506), .B(n2830), .Z(n2733) );
  XNOR U4324 ( .A(n2992), .B(n2733), .Z(out[180]) );
  IV U4325 ( .A(n3104), .Z(n4236) );
  XOR U4326 ( .A(in[654]), .B(n4236), .Z(n2994) );
  NOR U4327 ( .A(n3521), .B(n2832), .Z(n2734) );
  XNOR U4328 ( .A(n2994), .B(n2734), .Z(out[181]) );
  XNOR U4329 ( .A(in[655]), .B(n4237), .Z(n2999) );
  NOR U4330 ( .A(n3549), .B(n2834), .Z(n2735) );
  XNOR U4331 ( .A(n2999), .B(n2735), .Z(out[182]) );
  XNOR U4332 ( .A(in[656]), .B(n4240), .Z(n3002) );
  NOR U4333 ( .A(n3579), .B(n2836), .Z(n2736) );
  XNOR U4334 ( .A(n3002), .B(n2736), .Z(out[183]) );
  XNOR U4335 ( .A(in[657]), .B(n4241), .Z(n3005) );
  NOR U4336 ( .A(n3603), .B(n2838), .Z(n2737) );
  XNOR U4337 ( .A(n3005), .B(n2737), .Z(out[184]) );
  XNOR U4338 ( .A(in[658]), .B(n4246), .Z(n3008) );
  NOR U4339 ( .A(n3633), .B(n2840), .Z(n2738) );
  XNOR U4340 ( .A(n3008), .B(n2738), .Z(out[185]) );
  XNOR U4341 ( .A(in[659]), .B(n4249), .Z(n3011) );
  NOR U4342 ( .A(n3677), .B(n2845), .Z(n2739) );
  XNOR U4343 ( .A(n3011), .B(n2739), .Z(out[186]) );
  XOR U4344 ( .A(in[660]), .B(n4252), .Z(n3013) );
  NOR U4345 ( .A(n3721), .B(n2847), .Z(n2740) );
  XOR U4346 ( .A(n3013), .B(n2740), .Z(out[187]) );
  XOR U4347 ( .A(in[661]), .B(n4255), .Z(n3016) );
  NOR U4348 ( .A(n3767), .B(n2849), .Z(n2741) );
  XOR U4349 ( .A(n3016), .B(n2741), .Z(out[188]) );
  XOR U4350 ( .A(in[662]), .B(n4256), .Z(n3019) );
  XOR U4351 ( .A(in[1428]), .B(n3220), .Z(n4553) );
  XNOR U4352 ( .A(in[1051]), .B(n2742), .Z(n2905) );
  NANDN U4353 ( .A(n4553), .B(n2905), .Z(n2743) );
  XNOR U4354 ( .A(n4552), .B(n2743), .Z(out[18]) );
  XOR U4355 ( .A(in[663]), .B(n4257), .Z(n3020) );
  XOR U4356 ( .A(in[664]), .B(n4258), .Z(n3023) );
  NANDN U4357 ( .A(n2857), .B(n3942), .Z(n2744) );
  XOR U4358 ( .A(n2858), .B(n2744), .Z(out[192]) );
  XNOR U4359 ( .A(in[1034]), .B(n4458), .Z(n2761) );
  ANDN U4360 ( .B(n3985), .A(n2860), .Z(n2745) );
  XNOR U4361 ( .A(n2761), .B(n2745), .Z(out[193]) );
  XNOR U4362 ( .A(in[1035]), .B(n4461), .Z(n2974) );
  ANDN U4363 ( .B(n4029), .A(n2746), .Z(n2747) );
  XNOR U4364 ( .A(n2974), .B(n2747), .Z(out[194]) );
  XOR U4365 ( .A(n4464), .B(in[1036]), .Z(n3172) );
  ANDN U4366 ( .B(n4073), .A(n2748), .Z(n2749) );
  XNOR U4367 ( .A(n3172), .B(n2749), .Z(out[195]) );
  XOR U4368 ( .A(n4467), .B(in[1037]), .Z(n3428) );
  ANDN U4369 ( .B(n4117), .A(n2750), .Z(n2751) );
  XNOR U4370 ( .A(n3428), .B(n2751), .Z(out[196]) );
  XOR U4371 ( .A(n4470), .B(in[1038]), .Z(n3722) );
  ANDN U4372 ( .B(n4161), .A(n2752), .Z(n2753) );
  XNOR U4373 ( .A(n3722), .B(n2753), .Z(out[197]) );
  XOR U4374 ( .A(n4473), .B(in[1039]), .Z(n4162) );
  ANDN U4375 ( .B(n4199), .A(n2754), .Z(n2755) );
  XNOR U4376 ( .A(n4162), .B(n2755), .Z(out[198]) );
  XOR U4377 ( .A(n4476), .B(in[1040]), .Z(n4445) );
  ANDN U4378 ( .B(n4217), .A(n2756), .Z(n2757) );
  XNOR U4379 ( .A(n4445), .B(n2757), .Z(out[199]) );
  XOR U4380 ( .A(in[1429]), .B(n2758), .Z(n4582) );
  XNOR U4381 ( .A(in[1052]), .B(n2759), .Z(n2908) );
  NANDN U4382 ( .A(n4582), .B(n2908), .Z(n2760) );
  XNOR U4383 ( .A(n4581), .B(n2760), .Z(out[19]) );
  XOR U4384 ( .A(n3177), .B(in[1411]), .Z(n3983) );
  IV U4385 ( .A(n2761), .Z(n2859) );
  NANDN U4386 ( .A(n3983), .B(n2859), .Z(n2762) );
  XNOR U4387 ( .A(n3984), .B(n2762), .Z(out[1]) );
  XOR U4388 ( .A(n4483), .B(in[1041]), .Z(n4735) );
  ANDN U4389 ( .B(n4245), .A(n2763), .Z(n2764) );
  XNOR U4390 ( .A(n4735), .B(n2764), .Z(out[200]) );
  XOR U4391 ( .A(n4486), .B(in[1042]), .Z(n5164) );
  ANDN U4392 ( .B(n4263), .A(n2765), .Z(n2766) );
  XNOR U4393 ( .A(n5164), .B(n2766), .Z(out[201]) );
  NAND U4394 ( .A(n4289), .B(n2882), .Z(n2767) );
  XNOR U4395 ( .A(n2881), .B(n2767), .Z(out[202]) );
  NANDN U4396 ( .A(n2884), .B(n4314), .Z(n2768) );
  XNOR U4397 ( .A(n2885), .B(n2768), .Z(out[203]) );
  NANDN U4398 ( .A(n2886), .B(n4346), .Z(n2769) );
  XNOR U4399 ( .A(n2887), .B(n2769), .Z(out[204]) );
  NANDN U4400 ( .A(n2888), .B(n4377), .Z(n2770) );
  XNOR U4401 ( .A(n2889), .B(n2770), .Z(out[205]) );
  IV U4402 ( .A(n2771), .Z(n2894) );
  IV U4403 ( .A(n2772), .Z(n2897) );
  IV U4404 ( .A(n2773), .Z(n2900) );
  IV U4405 ( .A(n2774), .Z(n2903) );
  XOR U4406 ( .A(in[1430]), .B(n2775), .Z(n4607) );
  XNOR U4407 ( .A(in[1053]), .B(n2776), .Z(n2911) );
  NANDN U4408 ( .A(n4607), .B(n2911), .Z(n2777) );
  XNOR U4409 ( .A(n4606), .B(n2777), .Z(out[20]) );
  IV U4410 ( .A(n2778), .Z(n2906) );
  XOR U4411 ( .A(in[1054]), .B(n4526), .Z(n2783) );
  IV U4412 ( .A(n2783), .Z(n2914) );
  XOR U4413 ( .A(in[1055]), .B(n4530), .Z(n2797) );
  IV U4414 ( .A(n2797), .Z(n2917) );
  XOR U4415 ( .A(in[1056]), .B(n4534), .Z(n2820) );
  IV U4416 ( .A(n2820), .Z(n2920) );
  XOR U4417 ( .A(in[1057]), .B(n4538), .Z(n2843) );
  IV U4418 ( .A(n2843), .Z(n2926) );
  NOR U4419 ( .A(n4699), .B(n2927), .Z(n2779) );
  XOR U4420 ( .A(n2926), .B(n2779), .Z(out[216]) );
  XOR U4421 ( .A(in[1058]), .B(n4542), .Z(n2867) );
  IV U4422 ( .A(n2867), .Z(n2929) );
  XOR U4423 ( .A(in[1059]), .B(n4546), .Z(n2891) );
  IV U4424 ( .A(n2891), .Z(n2932) );
  NOR U4425 ( .A(n4781), .B(n2933), .Z(n2780) );
  XOR U4426 ( .A(n2932), .B(n2780), .Z(out[218]) );
  XNOR U4427 ( .A(in[1060]), .B(n4550), .Z(n2924) );
  IV U4428 ( .A(n2924), .Z(n2935) );
  NOR U4429 ( .A(n4824), .B(n2936), .Z(n2781) );
  XOR U4430 ( .A(n2935), .B(n2781), .Z(out[219]) );
  XOR U4431 ( .A(in[1431]), .B(n2782), .Z(n4636) );
  OR U4432 ( .A(n4636), .B(n2783), .Z(n2784) );
  XNOR U4433 ( .A(n4635), .B(n2784), .Z(out[21]) );
  XNOR U4434 ( .A(in[1061]), .B(n4556), .Z(n2950) );
  NOR U4435 ( .A(n4868), .B(n2938), .Z(n2785) );
  XNOR U4436 ( .A(n2950), .B(n2785), .Z(out[220]) );
  XNOR U4437 ( .A(in[1062]), .B(n4558), .Z(n2972) );
  NOR U4438 ( .A(n4912), .B(n2940), .Z(n2786) );
  XNOR U4439 ( .A(n2972), .B(n2786), .Z(out[221]) );
  XNOR U4440 ( .A(in[1063]), .B(n4339), .Z(n2996) );
  NOR U4441 ( .A(n4956), .B(n2942), .Z(n2787) );
  XNOR U4442 ( .A(n2996), .B(n2787), .Z(out[222]) );
  XNOR U4443 ( .A(in[1064]), .B(n4341), .Z(n3026) );
  NOR U4444 ( .A(n5000), .B(n2944), .Z(n2788) );
  XNOR U4445 ( .A(n3026), .B(n2788), .Z(out[223]) );
  XNOR U4446 ( .A(in[1065]), .B(n4347), .Z(n3046) );
  NOR U4447 ( .A(n5044), .B(n2946), .Z(n2789) );
  XNOR U4448 ( .A(n3046), .B(n2789), .Z(out[224]) );
  XNOR U4449 ( .A(in[1066]), .B(n4349), .Z(n3058) );
  NOR U4450 ( .A(n5085), .B(n2948), .Z(n2790) );
  XNOR U4451 ( .A(n3058), .B(n2790), .Z(out[225]) );
  XNOR U4452 ( .A(in[1067]), .B(n4351), .Z(n3079) );
  NOR U4453 ( .A(n5120), .B(n2952), .Z(n2791) );
  XNOR U4454 ( .A(n3079), .B(n2791), .Z(out[226]) );
  XNOR U4455 ( .A(in[1068]), .B(n4354), .Z(n3100) );
  XOR U4456 ( .A(in[1069]), .B(n4357), .Z(n3115) );
  NANDN U4457 ( .A(n2792), .B(n2956), .Z(n2793) );
  XNOR U4458 ( .A(n3115), .B(n2793), .Z(out[228]) );
  XOR U4459 ( .A(in[1070]), .B(n4360), .Z(n3139) );
  NANDN U4460 ( .A(n2794), .B(n2958), .Z(n2795) );
  XNOR U4461 ( .A(n3139), .B(n2795), .Z(out[229]) );
  XOR U4462 ( .A(in[1432]), .B(n2796), .Z(n4666) );
  OR U4463 ( .A(n4666), .B(n2797), .Z(n2798) );
  XNOR U4464 ( .A(n4665), .B(n2798), .Z(out[22]) );
  XNOR U4465 ( .A(in[1071]), .B(n4362), .Z(n3157) );
  NANDN U4466 ( .A(n2799), .B(n2960), .Z(n2800) );
  XOR U4467 ( .A(n3157), .B(n2800), .Z(out[230]) );
  XOR U4468 ( .A(in[1072]), .B(n4365), .Z(n3169) );
  NANDN U4469 ( .A(n2801), .B(n2962), .Z(n2802) );
  XNOR U4470 ( .A(n3169), .B(n2802), .Z(out[231]) );
  XOR U4471 ( .A(in[1073]), .B(n4368), .Z(n3194) );
  NANDN U4472 ( .A(n2803), .B(n2964), .Z(n2804) );
  XNOR U4473 ( .A(n3194), .B(n2804), .Z(out[232]) );
  XOR U4474 ( .A(in[1074]), .B(n4371), .Z(n3223) );
  NANDN U4475 ( .A(n2805), .B(n2966), .Z(n2806) );
  XNOR U4476 ( .A(n3223), .B(n2806), .Z(out[233]) );
  XOR U4477 ( .A(in[1075]), .B(n4378), .Z(n3247) );
  NANDN U4478 ( .A(n2807), .B(n2968), .Z(n2808) );
  XNOR U4479 ( .A(n3247), .B(n2808), .Z(out[234]) );
  XOR U4480 ( .A(in[1076]), .B(n4381), .Z(n3259) );
  NANDN U4481 ( .A(n2809), .B(n2970), .Z(n2810) );
  XNOR U4482 ( .A(n3259), .B(n2810), .Z(out[235]) );
  XOR U4483 ( .A(in[1077]), .B(n4384), .Z(n3269) );
  NANDN U4484 ( .A(n2811), .B(n2976), .Z(n2812) );
  XNOR U4485 ( .A(n3269), .B(n2812), .Z(out[236]) );
  XOR U4486 ( .A(in[1078]), .B(n4387), .Z(n3303) );
  NAND U4487 ( .A(n2813), .B(n2978), .Z(n2814) );
  XNOR U4488 ( .A(n3303), .B(n2814), .Z(out[237]) );
  XOR U4489 ( .A(in[1079]), .B(n4390), .Z(n3333) );
  NAND U4490 ( .A(n2815), .B(n2980), .Z(n2816) );
  XNOR U4491 ( .A(n3333), .B(n2816), .Z(out[238]) );
  XNOR U4492 ( .A(in[1080]), .B(n4392), .Z(n3361) );
  NAND U4493 ( .A(n2817), .B(n2982), .Z(n2818) );
  XOR U4494 ( .A(n3361), .B(n2818), .Z(out[239]) );
  XOR U4495 ( .A(in[1433]), .B(n2819), .Z(n4681) );
  OR U4496 ( .A(n4681), .B(n2820), .Z(n2821) );
  XNOR U4497 ( .A(n4680), .B(n2821), .Z(out[23]) );
  XOR U4498 ( .A(in[1081]), .B(n4395), .Z(n3389) );
  NAND U4499 ( .A(n2822), .B(n2984), .Z(n2823) );
  XNOR U4500 ( .A(n3389), .B(n2823), .Z(out[240]) );
  XOR U4501 ( .A(in[1082]), .B(n4398), .Z(n3424) );
  NAND U4502 ( .A(n2824), .B(n2986), .Z(n2825) );
  XOR U4503 ( .A(n3424), .B(n2825), .Z(out[241]) );
  XOR U4504 ( .A(in[1083]), .B(n4401), .Z(n3459) );
  NAND U4505 ( .A(n2826), .B(n2988), .Z(n2827) );
  XOR U4506 ( .A(n3459), .B(n2827), .Z(out[242]) );
  XNOR U4507 ( .A(in[1084]), .B(n4404), .Z(n3481) );
  NAND U4508 ( .A(n2828), .B(n2990), .Z(n2829) );
  XOR U4509 ( .A(n3481), .B(n2829), .Z(out[243]) );
  XNOR U4510 ( .A(in[1085]), .B(n4411), .Z(n3503) );
  NAND U4511 ( .A(n2830), .B(n2992), .Z(n2831) );
  XOR U4512 ( .A(n3503), .B(n2831), .Z(out[244]) );
  XNOR U4513 ( .A(in[1086]), .B(n4414), .Z(n3518) );
  NAND U4514 ( .A(n2832), .B(n2994), .Z(n2833) );
  XOR U4515 ( .A(n3518), .B(n2833), .Z(out[245]) );
  XOR U4516 ( .A(in[1087]), .B(n4417), .Z(n2998) );
  NAND U4517 ( .A(n2834), .B(n2999), .Z(n2835) );
  XNOR U4518 ( .A(n2998), .B(n2835), .Z(out[246]) );
  XOR U4519 ( .A(in[1024]), .B(n4420), .Z(n3001) );
  NAND U4520 ( .A(n2836), .B(n3002), .Z(n2837) );
  XNOR U4521 ( .A(n3001), .B(n2837), .Z(out[247]) );
  XOR U4522 ( .A(in[1025]), .B(n4423), .Z(n3004) );
  NAND U4523 ( .A(n2838), .B(n3005), .Z(n2839) );
  XNOR U4524 ( .A(n3004), .B(n2839), .Z(out[248]) );
  XOR U4525 ( .A(in[1026]), .B(n4426), .Z(n3007) );
  NAND U4526 ( .A(n2840), .B(n3008), .Z(n2841) );
  XNOR U4527 ( .A(n3007), .B(n2841), .Z(out[249]) );
  XOR U4528 ( .A(in[1434]), .B(n2842), .Z(n4698) );
  OR U4529 ( .A(n4698), .B(n2843), .Z(n2844) );
  XOR U4530 ( .A(n4697), .B(n2844), .Z(out[24]) );
  XOR U4531 ( .A(in[1027]), .B(n4429), .Z(n3010) );
  NAND U4532 ( .A(n2845), .B(n3011), .Z(n2846) );
  XNOR U4533 ( .A(n3010), .B(n2846), .Z(out[250]) );
  XOR U4534 ( .A(in[1028]), .B(n4432), .Z(n3014) );
  IV U4535 ( .A(n3014), .Z(n3718) );
  NANDN U4536 ( .A(n3013), .B(n2847), .Z(n2848) );
  XOR U4537 ( .A(n3718), .B(n2848), .Z(out[251]) );
  XOR U4538 ( .A(in[1029]), .B(n4435), .Z(n3017) );
  IV U4539 ( .A(n3017), .Z(n3764) );
  NANDN U4540 ( .A(n3016), .B(n2849), .Z(n2850) );
  XOR U4541 ( .A(n3764), .B(n2850), .Z(out[252]) );
  XOR U4542 ( .A(in[1030]), .B(n4438), .Z(n3808) );
  NANDN U4543 ( .A(n3019), .B(n2851), .Z(n2852) );
  XOR U4544 ( .A(n3808), .B(n2852), .Z(out[253]) );
  XOR U4545 ( .A(in[1031]), .B(n4449), .Z(n3021) );
  IV U4546 ( .A(n3021), .Z(n3852) );
  NANDN U4547 ( .A(n3020), .B(n2853), .Z(n2854) );
  XOR U4548 ( .A(n3852), .B(n2854), .Z(out[254]) );
  XOR U4549 ( .A(in[1032]), .B(n4452), .Z(n3024) );
  IV U4550 ( .A(n3024), .Z(n3896) );
  NANDN U4551 ( .A(n3023), .B(n2855), .Z(n2856) );
  XOR U4552 ( .A(n3896), .B(n2856), .Z(out[255]) );
  ANDN U4553 ( .B(n2860), .A(n2859), .Z(n2861) );
  XOR U4554 ( .A(n3983), .B(n2861), .Z(out[257]) );
  XNOR U4555 ( .A(n3945), .B(in[1412]), .Z(n4027) );
  NANDN U4556 ( .A(n2862), .B(n2974), .Z(n2863) );
  XNOR U4557 ( .A(n4027), .B(n2863), .Z(out[258]) );
  XNOR U4558 ( .A(n3949), .B(in[1413]), .Z(n4071) );
  NANDN U4559 ( .A(n2864), .B(n3172), .Z(n2865) );
  XNOR U4560 ( .A(n4071), .B(n2865), .Z(out[259]) );
  XOR U4561 ( .A(in[1435]), .B(n2866), .Z(n4732) );
  OR U4562 ( .A(n4732), .B(n2867), .Z(n2868) );
  XNOR U4563 ( .A(n4731), .B(n2868), .Z(out[25]) );
  XNOR U4564 ( .A(n3953), .B(in[1414]), .Z(n4115) );
  NANDN U4565 ( .A(n2869), .B(n3428), .Z(n2870) );
  XNOR U4566 ( .A(n4115), .B(n2870), .Z(out[260]) );
  XNOR U4567 ( .A(n3957), .B(in[1415]), .Z(n4159) );
  NANDN U4568 ( .A(n2871), .B(n3722), .Z(n2872) );
  XNOR U4569 ( .A(n4159), .B(n2872), .Z(out[261]) );
  XNOR U4570 ( .A(n3961), .B(in[1416]), .Z(n4197) );
  NANDN U4571 ( .A(n2873), .B(n4162), .Z(n2874) );
  XNOR U4572 ( .A(n4197), .B(n2874), .Z(out[262]) );
  XNOR U4573 ( .A(in[1417]), .B(n3965), .Z(n4446) );
  NANDN U4574 ( .A(n2875), .B(n4445), .Z(n2876) );
  XNOR U4575 ( .A(n4446), .B(n2876), .Z(out[263]) );
  XNOR U4576 ( .A(n3969), .B(in[1418]), .Z(n4736) );
  NANDN U4577 ( .A(n2877), .B(n4735), .Z(n2878) );
  XNOR U4578 ( .A(n4736), .B(n2878), .Z(out[264]) );
  XNOR U4579 ( .A(n3973), .B(in[1419]), .Z(n5165) );
  NANDN U4580 ( .A(n2879), .B(n5164), .Z(n2880) );
  XNOR U4581 ( .A(n5165), .B(n2880), .Z(out[265]) );
  NOR U4582 ( .A(n2882), .B(n2881), .Z(n2883) );
  XOR U4583 ( .A(n4287), .B(n2883), .Z(out[266]) );
  XOR U4584 ( .A(in[1436]), .B(n2890), .Z(n4780) );
  OR U4585 ( .A(n4780), .B(n2891), .Z(n2892) );
  XOR U4586 ( .A(n4779), .B(n2892), .Z(out[26]) );
  NOR U4587 ( .A(n2894), .B(n2893), .Z(n2895) );
  XOR U4588 ( .A(n4408), .B(n2895), .Z(out[270]) );
  NOR U4589 ( .A(n2897), .B(n2896), .Z(n2898) );
  XOR U4590 ( .A(n4442), .B(n2898), .Z(out[271]) );
  NOR U4591 ( .A(n2900), .B(n2899), .Z(n2901) );
  XOR U4592 ( .A(n4480), .B(n2901), .Z(out[272]) );
  NOR U4593 ( .A(n2903), .B(n2902), .Z(n2904) );
  XOR U4594 ( .A(n4514), .B(n2904), .Z(out[273]) );
  NOR U4595 ( .A(n2906), .B(n2905), .Z(n2907) );
  XOR U4596 ( .A(n4553), .B(n2907), .Z(out[274]) );
  NOR U4597 ( .A(n2909), .B(n2908), .Z(n2910) );
  XOR U4598 ( .A(n4582), .B(n2910), .Z(out[275]) );
  NOR U4599 ( .A(n2912), .B(n2911), .Z(n2913) );
  XOR U4600 ( .A(n4607), .B(n2913), .Z(out[276]) );
  ANDN U4601 ( .B(n2915), .A(n2914), .Z(n2916) );
  XOR U4602 ( .A(n4636), .B(n2916), .Z(out[277]) );
  ANDN U4603 ( .B(n2918), .A(n2917), .Z(n2919) );
  XOR U4604 ( .A(n4666), .B(n2919), .Z(out[278]) );
  ANDN U4605 ( .B(n2921), .A(n2920), .Z(n2922) );
  XOR U4606 ( .A(n4681), .B(n2922), .Z(out[279]) );
  XOR U4607 ( .A(in[1437]), .B(n2923), .Z(n4823) );
  OR U4608 ( .A(n4823), .B(n2924), .Z(n2925) );
  XOR U4609 ( .A(n4822), .B(n2925), .Z(out[27]) );
  ANDN U4610 ( .B(n2927), .A(n2926), .Z(n2928) );
  XOR U4611 ( .A(n4698), .B(n2928), .Z(out[280]) );
  ANDN U4612 ( .B(n2930), .A(n2929), .Z(n2931) );
  XOR U4613 ( .A(n4732), .B(n2931), .Z(out[281]) );
  ANDN U4614 ( .B(n2933), .A(n2932), .Z(n2934) );
  XOR U4615 ( .A(n4780), .B(n2934), .Z(out[282]) );
  ANDN U4616 ( .B(n2936), .A(n2935), .Z(n2937) );
  XOR U4617 ( .A(n4823), .B(n2937), .Z(out[283]) );
  XOR U4618 ( .A(in[1438]), .B(n4056), .Z(n4865) );
  NAND U4619 ( .A(n2938), .B(n2950), .Z(n2939) );
  XNOR U4620 ( .A(n4865), .B(n2939), .Z(out[284]) );
  XOR U4621 ( .A(in[1439]), .B(n4060), .Z(n4909) );
  NAND U4622 ( .A(n2940), .B(n2972), .Z(n2941) );
  XNOR U4623 ( .A(n4909), .B(n2941), .Z(out[285]) );
  XOR U4624 ( .A(in[1440]), .B(n4064), .Z(n4953) );
  NAND U4625 ( .A(n2942), .B(n2996), .Z(n2943) );
  XNOR U4626 ( .A(n4953), .B(n2943), .Z(out[286]) );
  XOR U4627 ( .A(in[1441]), .B(n4068), .Z(n4997) );
  NAND U4628 ( .A(n2944), .B(n3026), .Z(n2945) );
  XNOR U4629 ( .A(n4997), .B(n2945), .Z(out[287]) );
  XOR U4630 ( .A(in[1442]), .B(n4076), .Z(n5041) );
  NAND U4631 ( .A(n2946), .B(n3046), .Z(n2947) );
  XNOR U4632 ( .A(n5041), .B(n2947), .Z(out[288]) );
  XOR U4633 ( .A(in[1443]), .B(n4080), .Z(n5082) );
  NAND U4634 ( .A(n2948), .B(n3058), .Z(n2949) );
  XNOR U4635 ( .A(n5082), .B(n2949), .Z(out[289]) );
  OR U4636 ( .A(n4865), .B(n2950), .Z(n2951) );
  XOR U4637 ( .A(n4866), .B(n2951), .Z(out[28]) );
  XOR U4638 ( .A(in[1444]), .B(n4084), .Z(n5118) );
  NAND U4639 ( .A(n2952), .B(n3079), .Z(n2953) );
  XNOR U4640 ( .A(n5118), .B(n2953), .Z(out[290]) );
  XNOR U4641 ( .A(in[1445]), .B(n4088), .Z(n5161) );
  NANDN U4642 ( .A(n2954), .B(n3100), .Z(n2955) );
  XNOR U4643 ( .A(n5161), .B(n2955), .Z(out[291]) );
  OR U4644 ( .A(n3115), .B(n2956), .Z(n2957) );
  XNOR U4645 ( .A(n3114), .B(n2957), .Z(out[292]) );
  OR U4646 ( .A(n3139), .B(n2958), .Z(n2959) );
  XNOR U4647 ( .A(n3138), .B(n2959), .Z(out[293]) );
  NANDN U4648 ( .A(n2960), .B(n3157), .Z(n2961) );
  XNOR U4649 ( .A(n3158), .B(n2961), .Z(out[294]) );
  OR U4650 ( .A(n3169), .B(n2962), .Z(n2963) );
  XNOR U4651 ( .A(n3168), .B(n2963), .Z(out[295]) );
  OR U4652 ( .A(n3194), .B(n2964), .Z(n2965) );
  XNOR U4653 ( .A(n3193), .B(n2965), .Z(out[296]) );
  OR U4654 ( .A(n3223), .B(n2966), .Z(n2967) );
  XOR U4655 ( .A(n3224), .B(n2967), .Z(out[297]) );
  OR U4656 ( .A(n3247), .B(n2968), .Z(n2969) );
  XOR U4657 ( .A(n3248), .B(n2969), .Z(out[298]) );
  OR U4658 ( .A(n3259), .B(n2970), .Z(n2971) );
  XOR U4659 ( .A(n3260), .B(n2971), .Z(out[299]) );
  OR U4660 ( .A(n4909), .B(n2972), .Z(n2973) );
  XOR U4661 ( .A(n4910), .B(n2973), .Z(out[29]) );
  OR U4662 ( .A(n4027), .B(n2974), .Z(n2975) );
  XNOR U4663 ( .A(n4026), .B(n2975), .Z(out[2]) );
  OR U4664 ( .A(n3269), .B(n2976), .Z(n2977) );
  XOR U4665 ( .A(n3270), .B(n2977), .Z(out[300]) );
  OR U4666 ( .A(n3303), .B(n2978), .Z(n2979) );
  XOR U4667 ( .A(n3304), .B(n2979), .Z(out[301]) );
  OR U4668 ( .A(n3333), .B(n2980), .Z(n2981) );
  XOR U4669 ( .A(n3334), .B(n2981), .Z(out[302]) );
  NANDN U4670 ( .A(n2982), .B(n3361), .Z(n2983) );
  XOR U4671 ( .A(n3362), .B(n2983), .Z(out[303]) );
  OR U4672 ( .A(n3389), .B(n2984), .Z(n2985) );
  XOR U4673 ( .A(n3390), .B(n2985), .Z(out[304]) );
  NANDN U4674 ( .A(n2986), .B(n3424), .Z(n2987) );
  XOR U4675 ( .A(n3425), .B(n2987), .Z(out[305]) );
  NANDN U4676 ( .A(n2988), .B(n3459), .Z(n2989) );
  XOR U4677 ( .A(n3460), .B(n2989), .Z(out[306]) );
  NANDN U4678 ( .A(n2990), .B(n3481), .Z(n2991) );
  XOR U4679 ( .A(n3482), .B(n2991), .Z(out[307]) );
  NANDN U4680 ( .A(n2992), .B(n3503), .Z(n2993) );
  XOR U4681 ( .A(n3504), .B(n2993), .Z(out[308]) );
  NANDN U4682 ( .A(n2994), .B(n3518), .Z(n2995) );
  XOR U4683 ( .A(n3519), .B(n2995), .Z(out[309]) );
  OR U4684 ( .A(n4953), .B(n2996), .Z(n2997) );
  XOR U4685 ( .A(n4954), .B(n2997), .Z(out[30]) );
  IV U4686 ( .A(n2998), .Z(n3546) );
  NANDN U4687 ( .A(n2999), .B(n3546), .Z(n3000) );
  XOR U4688 ( .A(n3547), .B(n3000), .Z(out[310]) );
  IV U4689 ( .A(n3001), .Z(n3576) );
  NANDN U4690 ( .A(n3002), .B(n3576), .Z(n3003) );
  XOR U4691 ( .A(n3577), .B(n3003), .Z(out[311]) );
  IV U4692 ( .A(n3004), .Z(n3600) );
  NANDN U4693 ( .A(n3005), .B(n3600), .Z(n3006) );
  XOR U4694 ( .A(n3601), .B(n3006), .Z(out[312]) );
  IV U4695 ( .A(n3007), .Z(n3630) );
  NANDN U4696 ( .A(n3008), .B(n3630), .Z(n3009) );
  XOR U4697 ( .A(n3631), .B(n3009), .Z(out[313]) );
  IV U4698 ( .A(n3010), .Z(n3674) );
  NANDN U4699 ( .A(n3011), .B(n3674), .Z(n3012) );
  XOR U4700 ( .A(n3675), .B(n3012), .Z(out[314]) );
  NANDN U4701 ( .A(n3014), .B(n3013), .Z(n3015) );
  XOR U4702 ( .A(n3719), .B(n3015), .Z(out[315]) );
  NANDN U4703 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U4704 ( .A(n3765), .B(n3018), .Z(out[316]) );
  NANDN U4705 ( .A(n3021), .B(n3020), .Z(n3022) );
  XOR U4706 ( .A(n3853), .B(n3022), .Z(out[318]) );
  NANDN U4707 ( .A(n3024), .B(n3023), .Z(n3025) );
  XOR U4708 ( .A(n3897), .B(n3025), .Z(out[319]) );
  OR U4709 ( .A(n4997), .B(n3026), .Z(n3027) );
  XOR U4710 ( .A(n4998), .B(n3027), .Z(out[31]) );
  XOR U4711 ( .A(in[72]), .B(n4452), .Z(n3264) );
  XOR U4712 ( .A(in[1317]), .B(n4284), .Z(n3617) );
  XNOR U4713 ( .A(in[1244]), .B(n3028), .Z(n3614) );
  NANDN U4714 ( .A(n3617), .B(n3614), .Z(n3029) );
  XNOR U4715 ( .A(n3264), .B(n3029), .Z(out[320]) );
  XOR U4716 ( .A(in[73]), .B(n4455), .Z(n3151) );
  IV U4717 ( .A(n3151), .Z(n3267) );
  XOR U4718 ( .A(in[1318]), .B(n4290), .Z(n3621) );
  XNOR U4719 ( .A(in[1245]), .B(n3030), .Z(n3618) );
  NANDN U4720 ( .A(n3621), .B(n3618), .Z(n3031) );
  XOR U4721 ( .A(n3267), .B(n3031), .Z(out[321]) );
  XOR U4722 ( .A(in[74]), .B(n4458), .Z(n3153) );
  IV U4723 ( .A(n3153), .Z(n3274) );
  XOR U4724 ( .A(in[1319]), .B(n4292), .Z(n3625) );
  XNOR U4725 ( .A(in[1246]), .B(n3032), .Z(n3622) );
  NANDN U4726 ( .A(n3625), .B(n3622), .Z(n3033) );
  XOR U4727 ( .A(n3274), .B(n3033), .Z(out[322]) );
  XOR U4728 ( .A(in[75]), .B(n4461), .Z(n3155) );
  IV U4729 ( .A(n3155), .Z(n3277) );
  XOR U4730 ( .A(in[1320]), .B(n4294), .Z(n3629) );
  XNOR U4731 ( .A(in[1247]), .B(n3034), .Z(n3626) );
  NANDN U4732 ( .A(n3629), .B(n3626), .Z(n3035) );
  XOR U4733 ( .A(n3277), .B(n3035), .Z(out[323]) );
  XNOR U4734 ( .A(n4464), .B(in[76]), .Z(n3280) );
  XOR U4735 ( .A(in[1321]), .B(n4296), .Z(n3637) );
  XNOR U4736 ( .A(in[1248]), .B(n3036), .Z(n3634) );
  NANDN U4737 ( .A(n3637), .B(n3634), .Z(n3037) );
  XNOR U4738 ( .A(n3280), .B(n3037), .Z(out[324]) );
  XNOR U4739 ( .A(n4467), .B(in[77]), .Z(n3283) );
  XOR U4740 ( .A(in[1322]), .B(n4298), .Z(n3641) );
  XNOR U4741 ( .A(in[1249]), .B(n3038), .Z(n3638) );
  NANDN U4742 ( .A(n3641), .B(n3638), .Z(n3039) );
  XNOR U4743 ( .A(n3283), .B(n3039), .Z(out[325]) );
  XNOR U4744 ( .A(n4470), .B(in[78]), .Z(n3286) );
  XOR U4745 ( .A(in[1323]), .B(n4300), .Z(n3645) );
  XOR U4746 ( .A(in[1250]), .B(n4126), .Z(n3642) );
  NANDN U4747 ( .A(n3645), .B(n3642), .Z(n3040) );
  XNOR U4748 ( .A(n3286), .B(n3040), .Z(out[326]) );
  XNOR U4749 ( .A(n4473), .B(in[79]), .Z(n3289) );
  XOR U4750 ( .A(in[1324]), .B(n4302), .Z(n3649) );
  XNOR U4751 ( .A(in[1251]), .B(n3041), .Z(n3646) );
  NANDN U4752 ( .A(n3649), .B(n3646), .Z(n3042) );
  XNOR U4753 ( .A(n3289), .B(n3042), .Z(out[327]) );
  XNOR U4754 ( .A(n4476), .B(in[80]), .Z(n3292) );
  XOR U4755 ( .A(in[1325]), .B(n4304), .Z(n3653) );
  XNOR U4756 ( .A(in[1252]), .B(n3043), .Z(n3650) );
  NANDN U4757 ( .A(n3653), .B(n3650), .Z(n3044) );
  XNOR U4758 ( .A(n3292), .B(n3044), .Z(out[328]) );
  XNOR U4759 ( .A(n4483), .B(in[81]), .Z(n3295) );
  XNOR U4760 ( .A(in[1253]), .B(n4138), .Z(n3655) );
  XNOR U4761 ( .A(in[1326]), .B(n4306), .Z(n3657) );
  NANDN U4762 ( .A(n3655), .B(n3657), .Z(n3045) );
  XNOR U4763 ( .A(n3295), .B(n3045), .Z(out[329]) );
  OR U4764 ( .A(n5041), .B(n3046), .Z(n3047) );
  XOR U4765 ( .A(n5042), .B(n3047), .Z(out[32]) );
  XNOR U4766 ( .A(n4486), .B(in[82]), .Z(n3298) );
  XNOR U4767 ( .A(in[1254]), .B(n4142), .Z(n3659) );
  XNOR U4768 ( .A(in[1327]), .B(n4308), .Z(n3661) );
  NANDN U4769 ( .A(n3659), .B(n3661), .Z(n3048) );
  XNOR U4770 ( .A(n3298), .B(n3048), .Z(out[330]) );
  XNOR U4771 ( .A(n4489), .B(in[83]), .Z(n3301) );
  XNOR U4772 ( .A(in[1255]), .B(n4146), .Z(n3663) );
  XNOR U4773 ( .A(in[1328]), .B(n4315), .Z(n3665) );
  NANDN U4774 ( .A(n3663), .B(n3665), .Z(n3049) );
  XNOR U4775 ( .A(n3301), .B(n3049), .Z(out[331]) );
  XNOR U4776 ( .A(in[84]), .B(n4492), .Z(n3308) );
  XNOR U4777 ( .A(in[1256]), .B(n4150), .Z(n3667) );
  XNOR U4778 ( .A(in[1329]), .B(n4318), .Z(n3669) );
  NANDN U4779 ( .A(n3667), .B(n3669), .Z(n3050) );
  XNOR U4780 ( .A(n3308), .B(n3050), .Z(out[332]) );
  XNOR U4781 ( .A(in[85]), .B(n4495), .Z(n3311) );
  XNOR U4782 ( .A(in[1257]), .B(n4154), .Z(n3671) );
  XNOR U4783 ( .A(in[1330]), .B(n4321), .Z(n3673) );
  NANDN U4784 ( .A(n3671), .B(n3673), .Z(n3051) );
  XNOR U4785 ( .A(n3311), .B(n3051), .Z(out[333]) );
  XNOR U4786 ( .A(in[86]), .B(n4498), .Z(n3314) );
  XNOR U4787 ( .A(in[1258]), .B(n4164), .Z(n3679) );
  XNOR U4788 ( .A(in[1331]), .B(n4324), .Z(n3681) );
  NANDN U4789 ( .A(n3679), .B(n3681), .Z(n3052) );
  XNOR U4790 ( .A(n3314), .B(n3052), .Z(out[334]) );
  XNOR U4791 ( .A(in[87]), .B(n4501), .Z(n3317) );
  XNOR U4792 ( .A(in[1259]), .B(n4168), .Z(n3683) );
  XNOR U4793 ( .A(in[1332]), .B(n4327), .Z(n3685) );
  NANDN U4794 ( .A(n3683), .B(n3685), .Z(n3053) );
  XNOR U4795 ( .A(n3317), .B(n3053), .Z(out[335]) );
  XNOR U4796 ( .A(in[88]), .B(n4504), .Z(n3320) );
  XNOR U4797 ( .A(in[1260]), .B(n4172), .Z(n3687) );
  XNOR U4798 ( .A(in[1333]), .B(n4330), .Z(n3689) );
  NANDN U4799 ( .A(n3687), .B(n3689), .Z(n3054) );
  XNOR U4800 ( .A(n3320), .B(n3054), .Z(out[336]) );
  XNOR U4801 ( .A(in[89]), .B(n4507), .Z(n3323) );
  XNOR U4802 ( .A(in[1261]), .B(n4176), .Z(n3691) );
  XNOR U4803 ( .A(in[1334]), .B(n4333), .Z(n3693) );
  NANDN U4804 ( .A(n3691), .B(n3693), .Z(n3055) );
  XNOR U4805 ( .A(n3323), .B(n3055), .Z(out[337]) );
  XNOR U4806 ( .A(in[90]), .B(n4510), .Z(n3325) );
  XNOR U4807 ( .A(in[1262]), .B(n3900), .Z(n3695) );
  XNOR U4808 ( .A(in[1335]), .B(n4336), .Z(n3697) );
  NANDN U4809 ( .A(n3695), .B(n3697), .Z(n3056) );
  XNOR U4810 ( .A(n3325), .B(n3056), .Z(out[338]) );
  XOR U4811 ( .A(in[91]), .B(n4517), .Z(n3327) );
  XNOR U4812 ( .A(in[1263]), .B(n3904), .Z(n3699) );
  XNOR U4813 ( .A(in[1336]), .B(n4180), .Z(n3701) );
  NANDN U4814 ( .A(n3699), .B(n3701), .Z(n3057) );
  XNOR U4815 ( .A(n3327), .B(n3057), .Z(out[339]) );
  OR U4816 ( .A(n5082), .B(n3058), .Z(n3059) );
  XOR U4817 ( .A(n5083), .B(n3059), .Z(out[33]) );
  XOR U4818 ( .A(in[92]), .B(n4520), .Z(n3329) );
  XNOR U4819 ( .A(in[1264]), .B(n3908), .Z(n3703) );
  XNOR U4820 ( .A(in[1337]), .B(n4183), .Z(n3705) );
  NANDN U4821 ( .A(n3703), .B(n3705), .Z(n3060) );
  XNOR U4822 ( .A(n3329), .B(n3060), .Z(out[340]) );
  XOR U4823 ( .A(in[93]), .B(n4523), .Z(n3331) );
  XNOR U4824 ( .A(in[1265]), .B(n3912), .Z(n3707) );
  XNOR U4825 ( .A(in[1338]), .B(n4186), .Z(n3709) );
  NANDN U4826 ( .A(n3707), .B(n3709), .Z(n3061) );
  XNOR U4827 ( .A(n3331), .B(n3061), .Z(out[341]) );
  XNOR U4828 ( .A(in[94]), .B(n4526), .Z(n3337) );
  XNOR U4829 ( .A(in[1266]), .B(n3916), .Z(n3711) );
  XNOR U4830 ( .A(in[1339]), .B(n4189), .Z(n3713) );
  NANDN U4831 ( .A(n3711), .B(n3713), .Z(n3062) );
  XNOR U4832 ( .A(n3337), .B(n3062), .Z(out[342]) );
  XNOR U4833 ( .A(in[95]), .B(n4530), .Z(n3339) );
  XOR U4834 ( .A(in[1267]), .B(n3920), .Z(n3715) );
  XNOR U4835 ( .A(in[1340]), .B(n3063), .Z(n3717) );
  NANDN U4836 ( .A(n3715), .B(n3717), .Z(n3064) );
  XNOR U4837 ( .A(n3339), .B(n3064), .Z(out[343]) );
  XNOR U4838 ( .A(in[96]), .B(n4534), .Z(n3341) );
  XOR U4839 ( .A(in[1268]), .B(n3924), .Z(n3725) );
  XNOR U4840 ( .A(in[1341]), .B(n3065), .Z(n3727) );
  NANDN U4841 ( .A(n3725), .B(n3727), .Z(n3066) );
  XNOR U4842 ( .A(n3341), .B(n3066), .Z(out[344]) );
  XNOR U4843 ( .A(in[97]), .B(n4538), .Z(n3343) );
  XOR U4844 ( .A(in[1269]), .B(n3928), .Z(n3729) );
  XNOR U4845 ( .A(in[1342]), .B(n3067), .Z(n3731) );
  NANDN U4846 ( .A(n3729), .B(n3731), .Z(n3068) );
  XNOR U4847 ( .A(n3343), .B(n3068), .Z(out[345]) );
  XNOR U4848 ( .A(in[98]), .B(n4542), .Z(n3345) );
  IV U4849 ( .A(n3069), .Z(n3932) );
  XOR U4850 ( .A(in[1270]), .B(n3932), .Z(n3733) );
  XNOR U4851 ( .A(in[1343]), .B(n4201), .Z(n3735) );
  NANDN U4852 ( .A(n3733), .B(n3735), .Z(n3070) );
  XNOR U4853 ( .A(n3345), .B(n3070), .Z(out[346]) );
  XNOR U4854 ( .A(in[99]), .B(n4546), .Z(n3347) );
  IV U4855 ( .A(n3071), .Z(n3936) );
  XOR U4856 ( .A(in[1271]), .B(n3936), .Z(n3737) );
  XNOR U4857 ( .A(in[1280]), .B(n3072), .Z(n3739) );
  NANDN U4858 ( .A(n3737), .B(n3739), .Z(n3073) );
  XNOR U4859 ( .A(n3347), .B(n3073), .Z(out[347]) );
  XOR U4860 ( .A(in[100]), .B(n4550), .Z(n3201) );
  IV U4861 ( .A(n3201), .Z(n3350) );
  IV U4862 ( .A(n3074), .Z(n3943) );
  XOR U4863 ( .A(in[1272]), .B(n3943), .Z(n3741) );
  XNOR U4864 ( .A(in[1281]), .B(n3075), .Z(n3743) );
  NANDN U4865 ( .A(n3741), .B(n3743), .Z(n3076) );
  XOR U4866 ( .A(n3350), .B(n3076), .Z(out[348]) );
  XOR U4867 ( .A(in[101]), .B(n4556), .Z(n3204) );
  IV U4868 ( .A(n3204), .Z(n3353) );
  XOR U4869 ( .A(in[1273]), .B(n3947), .Z(n3745) );
  XNOR U4870 ( .A(in[1282]), .B(n3077), .Z(n3747) );
  NANDN U4871 ( .A(n3745), .B(n3747), .Z(n3078) );
  XOR U4872 ( .A(n3353), .B(n3078), .Z(out[349]) );
  OR U4873 ( .A(n5118), .B(n3079), .Z(n3080) );
  XNOR U4874 ( .A(n5117), .B(n3080), .Z(out[34]) );
  XOR U4875 ( .A(in[102]), .B(n4558), .Z(n3207) );
  IV U4876 ( .A(n3207), .Z(n3356) );
  XOR U4877 ( .A(in[1274]), .B(n3951), .Z(n3749) );
  XNOR U4878 ( .A(in[1283]), .B(n3081), .Z(n3751) );
  NANDN U4879 ( .A(n3749), .B(n3751), .Z(n3082) );
  XOR U4880 ( .A(n3356), .B(n3082), .Z(out[350]) );
  XOR U4881 ( .A(in[103]), .B(n4339), .Z(n3210) );
  IV U4882 ( .A(n3210), .Z(n3359) );
  XNOR U4883 ( .A(in[1275]), .B(n3955), .Z(n3753) );
  XNOR U4884 ( .A(in[1284]), .B(n3083), .Z(n3755) );
  NANDN U4885 ( .A(n3753), .B(n3755), .Z(n3084) );
  XOR U4886 ( .A(n3359), .B(n3084), .Z(out[351]) );
  XOR U4887 ( .A(in[104]), .B(n4341), .Z(n3213) );
  IV U4888 ( .A(n3213), .Z(n3366) );
  XNOR U4889 ( .A(in[1276]), .B(n3959), .Z(n3757) );
  XNOR U4890 ( .A(in[1285]), .B(n3085), .Z(n3759) );
  NANDN U4891 ( .A(n3757), .B(n3759), .Z(n3086) );
  XOR U4892 ( .A(n3366), .B(n3086), .Z(out[352]) );
  XOR U4893 ( .A(in[105]), .B(n4347), .Z(n3215) );
  IV U4894 ( .A(n3215), .Z(n3369) );
  XNOR U4895 ( .A(in[1277]), .B(n3963), .Z(n3761) );
  XNOR U4896 ( .A(in[1286]), .B(n3087), .Z(n3763) );
  NANDN U4897 ( .A(n3761), .B(n3763), .Z(n3088) );
  XOR U4898 ( .A(n3369), .B(n3088), .Z(out[353]) );
  XOR U4899 ( .A(in[106]), .B(n4349), .Z(n3218) );
  IV U4900 ( .A(n3218), .Z(n3372) );
  XNOR U4901 ( .A(in[1278]), .B(n3967), .Z(n3769) );
  XNOR U4902 ( .A(in[1287]), .B(n3089), .Z(n3771) );
  NANDN U4903 ( .A(n3769), .B(n3771), .Z(n3090) );
  XOR U4904 ( .A(n3372), .B(n3090), .Z(out[354]) );
  XOR U4905 ( .A(in[107]), .B(n4351), .Z(n3221) );
  IV U4906 ( .A(n3221), .Z(n3375) );
  XNOR U4907 ( .A(in[1279]), .B(n3971), .Z(n3773) );
  XNOR U4908 ( .A(in[1288]), .B(n4218), .Z(n3775) );
  NANDN U4909 ( .A(n3773), .B(n3775), .Z(n3091) );
  XOR U4910 ( .A(n3375), .B(n3091), .Z(out[355]) );
  XOR U4911 ( .A(in[108]), .B(n4354), .Z(n3227) );
  IV U4912 ( .A(n3227), .Z(n3377) );
  XNOR U4913 ( .A(in[1216]), .B(n3975), .Z(n3777) );
  XNOR U4914 ( .A(in[1289]), .B(n3092), .Z(n3779) );
  NANDN U4915 ( .A(n3777), .B(n3779), .Z(n3093) );
  XOR U4916 ( .A(n3377), .B(n3093), .Z(out[356]) );
  XOR U4917 ( .A(in[109]), .B(n4357), .Z(n3229) );
  IV U4918 ( .A(n3229), .Z(n3379) );
  XNOR U4919 ( .A(in[1217]), .B(n3979), .Z(n3781) );
  XNOR U4920 ( .A(in[1290]), .B(n3094), .Z(n3783) );
  NANDN U4921 ( .A(n3781), .B(n3783), .Z(n3095) );
  XOR U4922 ( .A(n3379), .B(n3095), .Z(out[357]) );
  XOR U4923 ( .A(in[110]), .B(n4360), .Z(n3231) );
  IV U4924 ( .A(n3231), .Z(n3381) );
  XNOR U4925 ( .A(in[1218]), .B(n3986), .Z(n3785) );
  XNOR U4926 ( .A(in[1291]), .B(n3096), .Z(n3787) );
  NANDN U4927 ( .A(n3785), .B(n3787), .Z(n3097) );
  XOR U4928 ( .A(n3381), .B(n3097), .Z(out[358]) );
  XOR U4929 ( .A(in[111]), .B(n4362), .Z(n3233) );
  IV U4930 ( .A(n3233), .Z(n3383) );
  XNOR U4931 ( .A(in[1219]), .B(n3990), .Z(n3789) );
  XNOR U4932 ( .A(in[1292]), .B(n3098), .Z(n3791) );
  NANDN U4933 ( .A(n3789), .B(n3791), .Z(n3099) );
  XOR U4934 ( .A(n3383), .B(n3099), .Z(out[359]) );
  OR U4935 ( .A(n5161), .B(n3100), .Z(n3101) );
  XNOR U4936 ( .A(n5160), .B(n3101), .Z(out[35]) );
  XOR U4937 ( .A(in[112]), .B(n4365), .Z(n3235) );
  IV U4938 ( .A(n3235), .Z(n3385) );
  XOR U4939 ( .A(in[1293]), .B(n3102), .Z(n3795) );
  XOR U4940 ( .A(in[1220]), .B(n3994), .Z(n3792) );
  NANDN U4941 ( .A(n3795), .B(n3792), .Z(n3103) );
  XOR U4942 ( .A(n3385), .B(n3103), .Z(out[360]) );
  XOR U4943 ( .A(in[113]), .B(n4368), .Z(n3237) );
  IV U4944 ( .A(n3237), .Z(n3387) );
  XOR U4945 ( .A(in[1294]), .B(n3104), .Z(n3799) );
  XOR U4946 ( .A(in[1221]), .B(n3998), .Z(n3796) );
  NANDN U4947 ( .A(n3799), .B(n3796), .Z(n3105) );
  XOR U4948 ( .A(n3387), .B(n3105), .Z(out[361]) );
  XOR U4949 ( .A(in[114]), .B(n4371), .Z(n3239) );
  IV U4950 ( .A(n3239), .Z(n3393) );
  XOR U4951 ( .A(in[1295]), .B(n4237), .Z(n3803) );
  XOR U4952 ( .A(in[1222]), .B(n4002), .Z(n3800) );
  NANDN U4953 ( .A(n3803), .B(n3800), .Z(n3106) );
  XOR U4954 ( .A(n3393), .B(n3106), .Z(out[362]) );
  XOR U4955 ( .A(in[115]), .B(n4378), .Z(n3241) );
  IV U4956 ( .A(n3241), .Z(n3395) );
  XOR U4957 ( .A(in[1296]), .B(n4240), .Z(n3807) );
  XOR U4958 ( .A(in[1223]), .B(n4006), .Z(n3804) );
  NANDN U4959 ( .A(n3807), .B(n3804), .Z(n3107) );
  XOR U4960 ( .A(n3395), .B(n3107), .Z(out[363]) );
  XOR U4961 ( .A(in[116]), .B(n4381), .Z(n3243) );
  IV U4962 ( .A(n3243), .Z(n3398) );
  XOR U4963 ( .A(in[1297]), .B(n4241), .Z(n3815) );
  XOR U4964 ( .A(in[1224]), .B(n4010), .Z(n3812) );
  NANDN U4965 ( .A(n3815), .B(n3812), .Z(n3108) );
  XOR U4966 ( .A(n3398), .B(n3108), .Z(out[364]) );
  XOR U4967 ( .A(in[117]), .B(n4384), .Z(n3245) );
  IV U4968 ( .A(n3245), .Z(n3402) );
  XOR U4969 ( .A(in[1298]), .B(n4246), .Z(n3819) );
  XOR U4970 ( .A(in[1225]), .B(n4014), .Z(n3816) );
  NANDN U4971 ( .A(n3819), .B(n3816), .Z(n3109) );
  XOR U4972 ( .A(n3402), .B(n3109), .Z(out[365]) );
  XOR U4973 ( .A(in[118]), .B(n4387), .Z(n3251) );
  IV U4974 ( .A(n3251), .Z(n3406) );
  XOR U4975 ( .A(in[1299]), .B(n4249), .Z(n3823) );
  XOR U4976 ( .A(in[1226]), .B(n4018), .Z(n3820) );
  NANDN U4977 ( .A(n3823), .B(n3820), .Z(n3110) );
  XOR U4978 ( .A(n3406), .B(n3110), .Z(out[366]) );
  XOR U4979 ( .A(in[119]), .B(n4390), .Z(n3253) );
  IV U4980 ( .A(n3253), .Z(n3410) );
  XOR U4981 ( .A(in[1300]), .B(n4252), .Z(n3827) );
  XNOR U4982 ( .A(in[1227]), .B(n4022), .Z(n3824) );
  NANDN U4983 ( .A(n3827), .B(n3824), .Z(n3111) );
  XOR U4984 ( .A(n3410), .B(n3111), .Z(out[367]) );
  XOR U4985 ( .A(in[120]), .B(n4392), .Z(n3255) );
  IV U4986 ( .A(n3255), .Z(n3413) );
  XOR U4987 ( .A(in[1301]), .B(n4255), .Z(n3831) );
  XOR U4988 ( .A(in[1228]), .B(n4030), .Z(n3828) );
  NANDN U4989 ( .A(n3831), .B(n3828), .Z(n3112) );
  XOR U4990 ( .A(n3413), .B(n3112), .Z(out[368]) );
  XOR U4991 ( .A(in[121]), .B(n4395), .Z(n3257) );
  IV U4992 ( .A(n3257), .Z(n3416) );
  XOR U4993 ( .A(in[1302]), .B(n4256), .Z(n3835) );
  XOR U4994 ( .A(in[1229]), .B(n4034), .Z(n3832) );
  NANDN U4995 ( .A(n3835), .B(n3832), .Z(n3113) );
  XOR U4996 ( .A(n3416), .B(n3113), .Z(out[369]) );
  ANDN U4997 ( .B(n3115), .A(n3114), .Z(n3116) );
  XOR U4998 ( .A(n3117), .B(n3116), .Z(out[36]) );
  XOR U4999 ( .A(in[122]), .B(n4398), .Z(n3419) );
  XOR U5000 ( .A(in[1303]), .B(n4257), .Z(n3839) );
  XNOR U5001 ( .A(in[1230]), .B(n3118), .Z(n3836) );
  NANDN U5002 ( .A(n3839), .B(n3836), .Z(n3119) );
  XOR U5003 ( .A(n3419), .B(n3119), .Z(out[370]) );
  XOR U5004 ( .A(in[123]), .B(n4401), .Z(n3422) );
  XOR U5005 ( .A(in[1304]), .B(n4258), .Z(n3843) );
  XNOR U5006 ( .A(in[1231]), .B(n3120), .Z(n3840) );
  NANDN U5007 ( .A(n3843), .B(n3840), .Z(n3121) );
  XOR U5008 ( .A(n3422), .B(n3121), .Z(out[371]) );
  XOR U5009 ( .A(in[124]), .B(n4404), .Z(n3430) );
  XOR U5010 ( .A(in[1305]), .B(n4259), .Z(n3847) );
  XNOR U5011 ( .A(in[1232]), .B(n3122), .Z(n3844) );
  NANDN U5012 ( .A(n3847), .B(n3844), .Z(n3123) );
  XNOR U5013 ( .A(n3430), .B(n3123), .Z(out[372]) );
  XOR U5014 ( .A(in[125]), .B(n4411), .Z(n3433) );
  XOR U5015 ( .A(in[1306]), .B(n4260), .Z(n3851) );
  XNOR U5016 ( .A(in[1233]), .B(n3124), .Z(n3848) );
  NANDN U5017 ( .A(n3851), .B(n3848), .Z(n3125) );
  XNOR U5018 ( .A(n3433), .B(n3125), .Z(out[373]) );
  XOR U5019 ( .A(in[126]), .B(n4414), .Z(n3436) );
  XOR U5020 ( .A(in[1307]), .B(n4261), .Z(n3859) );
  XNOR U5021 ( .A(in[1234]), .B(n3126), .Z(n3856) );
  NANDN U5022 ( .A(n3859), .B(n3856), .Z(n3127) );
  XNOR U5023 ( .A(n3436), .B(n3127), .Z(out[374]) );
  XOR U5024 ( .A(in[127]), .B(n4417), .Z(n3439) );
  XOR U5025 ( .A(in[1308]), .B(n4264), .Z(n3863) );
  XNOR U5026 ( .A(in[1235]), .B(n3128), .Z(n3860) );
  NANDN U5027 ( .A(n3863), .B(n3860), .Z(n3129) );
  XNOR U5028 ( .A(n3439), .B(n3129), .Z(out[375]) );
  XOR U5029 ( .A(in[64]), .B(n4420), .Z(n3442) );
  XOR U5030 ( .A(in[1309]), .B(n4265), .Z(n3867) );
  XNOR U5031 ( .A(in[1236]), .B(n3130), .Z(n3864) );
  NANDN U5032 ( .A(n3867), .B(n3864), .Z(n3131) );
  XNOR U5033 ( .A(n3442), .B(n3131), .Z(out[376]) );
  XOR U5034 ( .A(in[65]), .B(n4423), .Z(n3445) );
  XOR U5035 ( .A(in[1310]), .B(n4266), .Z(n3871) );
  XNOR U5036 ( .A(in[1237]), .B(n3132), .Z(n3868) );
  NANDN U5037 ( .A(n3871), .B(n3868), .Z(n3133) );
  XNOR U5038 ( .A(n3445), .B(n3133), .Z(out[377]) );
  XOR U5039 ( .A(in[66]), .B(n4426), .Z(n3448) );
  XOR U5040 ( .A(in[1311]), .B(n4267), .Z(n3875) );
  XNOR U5041 ( .A(in[1238]), .B(n3134), .Z(n3872) );
  NANDN U5042 ( .A(n3875), .B(n3872), .Z(n3135) );
  XNOR U5043 ( .A(n3448), .B(n3135), .Z(out[378]) );
  XOR U5044 ( .A(in[67]), .B(n4429), .Z(n3451) );
  XOR U5045 ( .A(in[1312]), .B(n4270), .Z(n3879) );
  XNOR U5046 ( .A(in[1239]), .B(n3136), .Z(n3876) );
  NANDN U5047 ( .A(n3879), .B(n3876), .Z(n3137) );
  XNOR U5048 ( .A(n3451), .B(n3137), .Z(out[379]) );
  ANDN U5049 ( .B(n3139), .A(n3138), .Z(n3140) );
  XOR U5050 ( .A(n3141), .B(n3140), .Z(out[37]) );
  XOR U5051 ( .A(in[68]), .B(n4432), .Z(n3454) );
  XOR U5052 ( .A(in[1313]), .B(n4273), .Z(n3883) );
  XNOR U5053 ( .A(in[1240]), .B(n3142), .Z(n3880) );
  NANDN U5054 ( .A(n3883), .B(n3880), .Z(n3143) );
  XNOR U5055 ( .A(n3454), .B(n3143), .Z(out[380]) );
  XOR U5056 ( .A(in[69]), .B(n4435), .Z(n3457) );
  XOR U5057 ( .A(in[1314]), .B(n4276), .Z(n3887) );
  XNOR U5058 ( .A(in[1241]), .B(n3144), .Z(n3884) );
  NANDN U5059 ( .A(n3887), .B(n3884), .Z(n3145) );
  XNOR U5060 ( .A(n3457), .B(n3145), .Z(out[381]) );
  XOR U5061 ( .A(in[70]), .B(n4438), .Z(n3464) );
  XOR U5062 ( .A(in[1315]), .B(n3146), .Z(n3891) );
  XNOR U5063 ( .A(in[1242]), .B(n3147), .Z(n3888) );
  NANDN U5064 ( .A(n3891), .B(n3888), .Z(n3148) );
  XOR U5065 ( .A(n3464), .B(n3148), .Z(out[382]) );
  XOR U5066 ( .A(in[71]), .B(n4449), .Z(n3467) );
  XOR U5067 ( .A(in[1316]), .B(n4282), .Z(n3895) );
  XNOR U5068 ( .A(in[1243]), .B(n3149), .Z(n3892) );
  NANDN U5069 ( .A(n3895), .B(n3892), .Z(n3150) );
  XNOR U5070 ( .A(n3467), .B(n3150), .Z(out[383]) );
  XOR U5071 ( .A(in[497]), .B(n4139), .Z(n3469) );
  XOR U5072 ( .A(in[498]), .B(n4143), .Z(n3471) );
  ANDN U5073 ( .B(n3621), .A(n3151), .Z(n3152) );
  XNOR U5074 ( .A(n3471), .B(n3152), .Z(out[385]) );
  XOR U5075 ( .A(in[499]), .B(n4147), .Z(n3473) );
  ANDN U5076 ( .B(n3625), .A(n3153), .Z(n3154) );
  XNOR U5077 ( .A(n3473), .B(n3154), .Z(out[386]) );
  XOR U5078 ( .A(in[500]), .B(n4151), .Z(n3475) );
  ANDN U5079 ( .B(n3629), .A(n3155), .Z(n3156) );
  XNOR U5080 ( .A(n3475), .B(n3156), .Z(out[387]) );
  XOR U5081 ( .A(in[501]), .B(n4155), .Z(n3477) );
  XOR U5082 ( .A(in[502]), .B(n4165), .Z(n3478) );
  NOR U5083 ( .A(n3158), .B(n3157), .Z(n3159) );
  XOR U5084 ( .A(n3160), .B(n3159), .Z(out[38]) );
  XOR U5085 ( .A(in[503]), .B(n4169), .Z(n3479) );
  XOR U5086 ( .A(in[504]), .B(n4173), .Z(n3480) );
  XOR U5087 ( .A(in[505]), .B(n4177), .Z(n3485) );
  XOR U5088 ( .A(in[506]), .B(n3901), .Z(n3486) );
  NOR U5089 ( .A(n3657), .B(n3295), .Z(n3161) );
  XNOR U5090 ( .A(n3486), .B(n3161), .Z(out[393]) );
  XOR U5091 ( .A(in[507]), .B(n3905), .Z(n3488) );
  NOR U5092 ( .A(n3661), .B(n3298), .Z(n3162) );
  XNOR U5093 ( .A(n3488), .B(n3162), .Z(out[394]) );
  XOR U5094 ( .A(in[508]), .B(n3909), .Z(n3490) );
  NOR U5095 ( .A(n3665), .B(n3301), .Z(n3163) );
  XNOR U5096 ( .A(n3490), .B(n3163), .Z(out[395]) );
  XOR U5097 ( .A(in[509]), .B(n3913), .Z(n3492) );
  NOR U5098 ( .A(n3669), .B(n3308), .Z(n3164) );
  XNOR U5099 ( .A(n3492), .B(n3164), .Z(out[396]) );
  XOR U5100 ( .A(in[510]), .B(n3917), .Z(n3494) );
  NOR U5101 ( .A(n3673), .B(n3311), .Z(n3165) );
  XNOR U5102 ( .A(n3494), .B(n3165), .Z(out[397]) );
  XOR U5103 ( .A(in[511]), .B(n3921), .Z(n3496) );
  NOR U5104 ( .A(n3681), .B(n3314), .Z(n3166) );
  XNOR U5105 ( .A(n3496), .B(n3166), .Z(out[398]) );
  XOR U5106 ( .A(in[448]), .B(n3925), .Z(n3498) );
  NOR U5107 ( .A(n3685), .B(n3317), .Z(n3167) );
  XNOR U5108 ( .A(n3498), .B(n3167), .Z(out[399]) );
  ANDN U5109 ( .B(n3169), .A(n3168), .Z(n3170) );
  XOR U5110 ( .A(n3171), .B(n3170), .Z(out[39]) );
  OR U5111 ( .A(n4071), .B(n3172), .Z(n3173) );
  XNOR U5112 ( .A(n4070), .B(n3173), .Z(out[3]) );
  XOR U5113 ( .A(in[449]), .B(n3929), .Z(n3500) );
  NOR U5114 ( .A(n3689), .B(n3320), .Z(n3174) );
  XNOR U5115 ( .A(n3500), .B(n3174), .Z(out[400]) );
  XOR U5116 ( .A(n3175), .B(in[450]), .Z(n3502) );
  NOR U5117 ( .A(n3693), .B(n3323), .Z(n3176) );
  XOR U5118 ( .A(n3502), .B(n3176), .Z(out[401]) );
  XOR U5119 ( .A(n3177), .B(in[451]), .Z(n3507) );
  NOR U5120 ( .A(n3697), .B(n3325), .Z(n3178) );
  XOR U5121 ( .A(n3507), .B(n3178), .Z(out[402]) );
  XOR U5122 ( .A(n3179), .B(in[452]), .Z(n3508) );
  NOR U5123 ( .A(n3701), .B(n3327), .Z(n3180) );
  XOR U5124 ( .A(n3508), .B(n3180), .Z(out[403]) );
  XOR U5125 ( .A(n3181), .B(in[453]), .Z(n3509) );
  NOR U5126 ( .A(n3705), .B(n3329), .Z(n3182) );
  XOR U5127 ( .A(n3509), .B(n3182), .Z(out[404]) );
  XOR U5128 ( .A(n3183), .B(in[454]), .Z(n3510) );
  NOR U5129 ( .A(n3709), .B(n3331), .Z(n3184) );
  XOR U5130 ( .A(n3510), .B(n3184), .Z(out[405]) );
  XOR U5131 ( .A(n3185), .B(in[455]), .Z(n3511) );
  NOR U5132 ( .A(n3713), .B(n3337), .Z(n3186) );
  XOR U5133 ( .A(n3511), .B(n3186), .Z(out[406]) );
  XOR U5134 ( .A(n3187), .B(in[456]), .Z(n3512) );
  NOR U5135 ( .A(n3717), .B(n3339), .Z(n3188) );
  XOR U5136 ( .A(n3512), .B(n3188), .Z(out[407]) );
  XOR U5137 ( .A(in[457]), .B(n3189), .Z(n3513) );
  NOR U5138 ( .A(n3727), .B(n3341), .Z(n3190) );
  XOR U5139 ( .A(n3513), .B(n3190), .Z(out[408]) );
  XOR U5140 ( .A(n3191), .B(in[458]), .Z(n3514) );
  NOR U5141 ( .A(n3731), .B(n3343), .Z(n3192) );
  XOR U5142 ( .A(n3514), .B(n3192), .Z(out[409]) );
  ANDN U5143 ( .B(n3194), .A(n3193), .Z(n3195) );
  XNOR U5144 ( .A(n3196), .B(n3195), .Z(out[40]) );
  XOR U5145 ( .A(n3973), .B(in[459]), .Z(n3515) );
  NOR U5146 ( .A(n3735), .B(n3345), .Z(n3197) );
  XNOR U5147 ( .A(n3515), .B(n3197), .Z(out[410]) );
  XOR U5148 ( .A(in[460]), .B(n3198), .Z(n3517) );
  NOR U5149 ( .A(n3739), .B(n3347), .Z(n3199) );
  XOR U5150 ( .A(n3517), .B(n3199), .Z(out[411]) );
  XOR U5151 ( .A(in[461]), .B(n3200), .Z(n3349) );
  NOR U5152 ( .A(n3201), .B(n3743), .Z(n3202) );
  XOR U5153 ( .A(n3349), .B(n3202), .Z(out[412]) );
  XOR U5154 ( .A(in[462]), .B(n3203), .Z(n3352) );
  NOR U5155 ( .A(n3204), .B(n3747), .Z(n3205) );
  XOR U5156 ( .A(n3352), .B(n3205), .Z(out[413]) );
  XOR U5157 ( .A(in[463]), .B(n3206), .Z(n3355) );
  NOR U5158 ( .A(n3207), .B(n3751), .Z(n3208) );
  XOR U5159 ( .A(n3355), .B(n3208), .Z(out[414]) );
  XOR U5160 ( .A(in[464]), .B(n3209), .Z(n3358) );
  NOR U5161 ( .A(n3210), .B(n3755), .Z(n3211) );
  XOR U5162 ( .A(n3358), .B(n3211), .Z(out[415]) );
  XOR U5163 ( .A(in[465]), .B(n3212), .Z(n3365) );
  NOR U5164 ( .A(n3213), .B(n3759), .Z(n3214) );
  XOR U5165 ( .A(n3365), .B(n3214), .Z(out[416]) );
  XOR U5166 ( .A(in[466]), .B(n4004), .Z(n3368) );
  NOR U5167 ( .A(n3215), .B(n3763), .Z(n3216) );
  XOR U5168 ( .A(n3368), .B(n3216), .Z(out[417]) );
  XOR U5169 ( .A(in[467]), .B(n3217), .Z(n3371) );
  NOR U5170 ( .A(n3218), .B(n3771), .Z(n3219) );
  XOR U5171 ( .A(n3371), .B(n3219), .Z(out[418]) );
  XOR U5172 ( .A(in[468]), .B(n3220), .Z(n3374) );
  NOR U5173 ( .A(n3221), .B(n3775), .Z(n3222) );
  XOR U5174 ( .A(n3374), .B(n3222), .Z(out[419]) );
  AND U5175 ( .A(n3224), .B(n3223), .Z(n3225) );
  XNOR U5176 ( .A(n3226), .B(n3225), .Z(out[41]) );
  XOR U5177 ( .A(in[469]), .B(n4016), .Z(n3542) );
  NOR U5178 ( .A(n3227), .B(n3779), .Z(n3228) );
  XNOR U5179 ( .A(n3542), .B(n3228), .Z(out[420]) );
  XOR U5180 ( .A(in[470]), .B(n4020), .Z(n3544) );
  NOR U5181 ( .A(n3229), .B(n3783), .Z(n3230) );
  XNOR U5182 ( .A(n3544), .B(n3230), .Z(out[421]) );
  XOR U5183 ( .A(in[471]), .B(n4024), .Z(n3551) );
  NOR U5184 ( .A(n3231), .B(n3787), .Z(n3232) );
  XNOR U5185 ( .A(n3551), .B(n3232), .Z(out[422]) );
  XOR U5186 ( .A(in[472]), .B(n4032), .Z(n3554) );
  NOR U5187 ( .A(n3233), .B(n3791), .Z(n3234) );
  XNOR U5188 ( .A(n3554), .B(n3234), .Z(out[423]) );
  XOR U5189 ( .A(in[473]), .B(n4036), .Z(n3557) );
  ANDN U5190 ( .B(n3795), .A(n3235), .Z(n3236) );
  XNOR U5191 ( .A(n3557), .B(n3236), .Z(out[424]) );
  XOR U5192 ( .A(in[474]), .B(n4040), .Z(n3560) );
  ANDN U5193 ( .B(n3799), .A(n3237), .Z(n3238) );
  XNOR U5194 ( .A(n3560), .B(n3238), .Z(out[425]) );
  XOR U5195 ( .A(in[475]), .B(n4044), .Z(n3563) );
  ANDN U5196 ( .B(n3803), .A(n3239), .Z(n3240) );
  XNOR U5197 ( .A(n3563), .B(n3240), .Z(out[426]) );
  XOR U5198 ( .A(in[476]), .B(n4048), .Z(n3566) );
  ANDN U5199 ( .B(n3807), .A(n3241), .Z(n3242) );
  XNOR U5200 ( .A(n3566), .B(n3242), .Z(out[427]) );
  XOR U5201 ( .A(in[477]), .B(n4052), .Z(n3568) );
  ANDN U5202 ( .B(n3815), .A(n3243), .Z(n3244) );
  XNOR U5203 ( .A(n3568), .B(n3244), .Z(out[428]) );
  XOR U5204 ( .A(in[478]), .B(n4056), .Z(n3401) );
  ANDN U5205 ( .B(n3819), .A(n3245), .Z(n3246) );
  XOR U5206 ( .A(n3401), .B(n3246), .Z(out[429]) );
  AND U5207 ( .A(n3248), .B(n3247), .Z(n3249) );
  XNOR U5208 ( .A(n3250), .B(n3249), .Z(out[42]) );
  XOR U5209 ( .A(in[479]), .B(n4060), .Z(n3405) );
  ANDN U5210 ( .B(n3823), .A(n3251), .Z(n3252) );
  XOR U5211 ( .A(n3405), .B(n3252), .Z(out[430]) );
  XOR U5212 ( .A(in[480]), .B(n4064), .Z(n3409) );
  ANDN U5213 ( .B(n3827), .A(n3253), .Z(n3254) );
  XOR U5214 ( .A(n3409), .B(n3254), .Z(out[431]) );
  XOR U5215 ( .A(in[481]), .B(n4068), .Z(n3412) );
  ANDN U5216 ( .B(n3831), .A(n3255), .Z(n3256) );
  XOR U5217 ( .A(n3412), .B(n3256), .Z(out[432]) );
  XOR U5218 ( .A(in[482]), .B(n4076), .Z(n3415) );
  ANDN U5219 ( .B(n3835), .A(n3257), .Z(n3258) );
  XOR U5220 ( .A(n3415), .B(n3258), .Z(out[433]) );
  XOR U5221 ( .A(in[483]), .B(n4080), .Z(n3418) );
  XOR U5222 ( .A(in[484]), .B(n4084), .Z(n3421) );
  XOR U5223 ( .A(in[485]), .B(n4088), .Z(n3588) );
  XOR U5224 ( .A(in[486]), .B(n4091), .Z(n3590) );
  XOR U5225 ( .A(in[487]), .B(n4095), .Z(n3592) );
  XOR U5226 ( .A(in[488]), .B(n4099), .Z(n3594) );
  AND U5227 ( .A(n3260), .B(n3259), .Z(n3261) );
  XNOR U5228 ( .A(n3262), .B(n3261), .Z(out[43]) );
  XOR U5229 ( .A(in[489]), .B(n4103), .Z(n3596) );
  XOR U5230 ( .A(in[490]), .B(n4107), .Z(n3598) );
  XOR U5231 ( .A(in[491]), .B(n4111), .Z(n3604) );
  XOR U5232 ( .A(in[492]), .B(n4119), .Z(n3605) );
  XOR U5233 ( .A(in[493]), .B(n4123), .Z(n3606) );
  XOR U5234 ( .A(in[494]), .B(n4127), .Z(n3608) );
  XOR U5235 ( .A(in[495]), .B(n4131), .Z(n3610) );
  XOR U5236 ( .A(in[496]), .B(n4135), .Z(n3612) );
  XOR U5237 ( .A(in[886]), .B(n3263), .Z(n3615) );
  NAND U5238 ( .A(n3264), .B(n3469), .Z(n3265) );
  XOR U5239 ( .A(n3615), .B(n3265), .Z(out[448]) );
  XOR U5240 ( .A(in[887]), .B(n3266), .Z(n3619) );
  NANDN U5241 ( .A(n3267), .B(n3471), .Z(n3268) );
  XOR U5242 ( .A(n3619), .B(n3268), .Z(out[449]) );
  AND U5243 ( .A(n3270), .B(n3269), .Z(n3271) );
  XNOR U5244 ( .A(n3272), .B(n3271), .Z(out[44]) );
  XOR U5245 ( .A(in[888]), .B(n3273), .Z(n3623) );
  NANDN U5246 ( .A(n3274), .B(n3473), .Z(n3275) );
  XOR U5247 ( .A(n3623), .B(n3275), .Z(out[450]) );
  XOR U5248 ( .A(in[889]), .B(n3276), .Z(n3627) );
  NANDN U5249 ( .A(n3277), .B(n3475), .Z(n3278) );
  XOR U5250 ( .A(n3627), .B(n3278), .Z(out[451]) );
  XOR U5251 ( .A(in[890]), .B(n3279), .Z(n3635) );
  NANDN U5252 ( .A(n3477), .B(n3280), .Z(n3281) );
  XOR U5253 ( .A(n3635), .B(n3281), .Z(out[452]) );
  XOR U5254 ( .A(in[891]), .B(n3282), .Z(n3639) );
  NANDN U5255 ( .A(n3478), .B(n3283), .Z(n3284) );
  XNOR U5256 ( .A(n3639), .B(n3284), .Z(out[453]) );
  XOR U5257 ( .A(in[892]), .B(n3285), .Z(n3643) );
  NANDN U5258 ( .A(n3479), .B(n3286), .Z(n3287) );
  XNOR U5259 ( .A(n3643), .B(n3287), .Z(out[454]) );
  XOR U5260 ( .A(in[893]), .B(n3288), .Z(n3647) );
  NANDN U5261 ( .A(n3480), .B(n3289), .Z(n3290) );
  XNOR U5262 ( .A(n3647), .B(n3290), .Z(out[455]) );
  XOR U5263 ( .A(in[894]), .B(n3291), .Z(n3651) );
  NANDN U5264 ( .A(n3485), .B(n3292), .Z(n3293) );
  XOR U5265 ( .A(n3651), .B(n3293), .Z(out[456]) );
  IV U5266 ( .A(n3294), .Z(n3902) );
  XOR U5267 ( .A(in[895]), .B(n3902), .Z(n3654) );
  NAND U5268 ( .A(n3295), .B(n3486), .Z(n3296) );
  XNOR U5269 ( .A(n3654), .B(n3296), .Z(out[457]) );
  IV U5270 ( .A(n3297), .Z(n3906) );
  XOR U5271 ( .A(in[832]), .B(n3906), .Z(n3658) );
  NAND U5272 ( .A(n3298), .B(n3488), .Z(n3299) );
  XNOR U5273 ( .A(n3658), .B(n3299), .Z(out[458]) );
  IV U5274 ( .A(n3300), .Z(n3910) );
  XOR U5275 ( .A(in[833]), .B(n3910), .Z(n3662) );
  NAND U5276 ( .A(n3301), .B(n3490), .Z(n3302) );
  XNOR U5277 ( .A(n3662), .B(n3302), .Z(out[459]) );
  AND U5278 ( .A(n3304), .B(n3303), .Z(n3305) );
  XNOR U5279 ( .A(n3306), .B(n3305), .Z(out[45]) );
  IV U5280 ( .A(n3307), .Z(n3914) );
  XOR U5281 ( .A(in[834]), .B(n3914), .Z(n3666) );
  NAND U5282 ( .A(n3308), .B(n3492), .Z(n3309) );
  XNOR U5283 ( .A(n3666), .B(n3309), .Z(out[460]) );
  IV U5284 ( .A(n3310), .Z(n3918) );
  XOR U5285 ( .A(in[835]), .B(n3918), .Z(n3670) );
  NAND U5286 ( .A(n3311), .B(n3494), .Z(n3312) );
  XNOR U5287 ( .A(n3670), .B(n3312), .Z(out[461]) );
  IV U5288 ( .A(n3313), .Z(n3922) );
  XOR U5289 ( .A(in[836]), .B(n3922), .Z(n3678) );
  NAND U5290 ( .A(n3314), .B(n3496), .Z(n3315) );
  XNOR U5291 ( .A(n3678), .B(n3315), .Z(out[462]) );
  IV U5292 ( .A(n3316), .Z(n3926) );
  XOR U5293 ( .A(in[837]), .B(n3926), .Z(n3682) );
  NAND U5294 ( .A(n3317), .B(n3498), .Z(n3318) );
  XNOR U5295 ( .A(n3682), .B(n3318), .Z(out[463]) );
  IV U5296 ( .A(n3319), .Z(n3930) );
  XOR U5297 ( .A(in[838]), .B(n3930), .Z(n3686) );
  NAND U5298 ( .A(n3320), .B(n3500), .Z(n3321) );
  XNOR U5299 ( .A(n3686), .B(n3321), .Z(out[464]) );
  XNOR U5300 ( .A(in[839]), .B(n3322), .Z(n3690) );
  NANDN U5301 ( .A(n3502), .B(n3323), .Z(n3324) );
  XNOR U5302 ( .A(n3690), .B(n3324), .Z(out[465]) );
  XNOR U5303 ( .A(in[840]), .B(n3937), .Z(n3694) );
  NANDN U5304 ( .A(n3507), .B(n3325), .Z(n3326) );
  XNOR U5305 ( .A(n3694), .B(n3326), .Z(out[466]) );
  XNOR U5306 ( .A(in[841]), .B(n3944), .Z(n3698) );
  NANDN U5307 ( .A(n3508), .B(n3327), .Z(n3328) );
  XNOR U5308 ( .A(n3698), .B(n3328), .Z(out[467]) );
  XNOR U5309 ( .A(in[842]), .B(n3948), .Z(n3702) );
  NANDN U5310 ( .A(n3509), .B(n3329), .Z(n3330) );
  XNOR U5311 ( .A(n3702), .B(n3330), .Z(out[468]) );
  XNOR U5312 ( .A(in[843]), .B(n3952), .Z(n3706) );
  NANDN U5313 ( .A(n3510), .B(n3331), .Z(n3332) );
  XNOR U5314 ( .A(n3706), .B(n3332), .Z(out[469]) );
  AND U5315 ( .A(n3334), .B(n3333), .Z(n3335) );
  XNOR U5316 ( .A(n3336), .B(n3335), .Z(out[46]) );
  XNOR U5317 ( .A(in[844]), .B(n3956), .Z(n3710) );
  NANDN U5318 ( .A(n3511), .B(n3337), .Z(n3338) );
  XNOR U5319 ( .A(n3710), .B(n3338), .Z(out[470]) );
  XNOR U5320 ( .A(in[845]), .B(n3960), .Z(n3714) );
  NANDN U5321 ( .A(n3512), .B(n3339), .Z(n3340) );
  XNOR U5322 ( .A(n3714), .B(n3340), .Z(out[471]) );
  XNOR U5323 ( .A(in[846]), .B(n3964), .Z(n3724) );
  NANDN U5324 ( .A(n3513), .B(n3341), .Z(n3342) );
  XNOR U5325 ( .A(n3724), .B(n3342), .Z(out[472]) );
  XNOR U5326 ( .A(in[847]), .B(n3968), .Z(n3728) );
  NANDN U5327 ( .A(n3514), .B(n3343), .Z(n3344) );
  XNOR U5328 ( .A(n3728), .B(n3344), .Z(out[473]) );
  XNOR U5329 ( .A(in[848]), .B(n3972), .Z(n3732) );
  NAND U5330 ( .A(n3345), .B(n3515), .Z(n3346) );
  XNOR U5331 ( .A(n3732), .B(n3346), .Z(out[474]) );
  XNOR U5332 ( .A(in[849]), .B(n3976), .Z(n3736) );
  NANDN U5333 ( .A(n3517), .B(n3347), .Z(n3348) );
  XNOR U5334 ( .A(n3736), .B(n3348), .Z(out[475]) );
  XNOR U5335 ( .A(in[850]), .B(n3980), .Z(n3740) );
  IV U5336 ( .A(n3349), .Z(n3522) );
  NANDN U5337 ( .A(n3350), .B(n3522), .Z(n3351) );
  XNOR U5338 ( .A(n3740), .B(n3351), .Z(out[476]) );
  XOR U5339 ( .A(in[851]), .B(n3987), .Z(n3524) );
  IV U5340 ( .A(n3352), .Z(n3525) );
  NANDN U5341 ( .A(n3353), .B(n3525), .Z(n3354) );
  XNOR U5342 ( .A(n3524), .B(n3354), .Z(out[477]) );
  XOR U5343 ( .A(in[852]), .B(n3991), .Z(n3527) );
  IV U5344 ( .A(n3355), .Z(n3528) );
  NANDN U5345 ( .A(n3356), .B(n3528), .Z(n3357) );
  XNOR U5346 ( .A(n3527), .B(n3357), .Z(out[478]) );
  XOR U5347 ( .A(in[853]), .B(n3995), .Z(n3530) );
  IV U5348 ( .A(n3358), .Z(n3531) );
  NANDN U5349 ( .A(n3359), .B(n3531), .Z(n3360) );
  XNOR U5350 ( .A(n3530), .B(n3360), .Z(out[479]) );
  ANDN U5351 ( .B(n3362), .A(n3361), .Z(n3363) );
  XNOR U5352 ( .A(n3364), .B(n3363), .Z(out[47]) );
  XOR U5353 ( .A(in[854]), .B(n3999), .Z(n3756) );
  IV U5354 ( .A(n3365), .Z(n3533) );
  NANDN U5355 ( .A(n3366), .B(n3533), .Z(n3367) );
  XOR U5356 ( .A(n3756), .B(n3367), .Z(out[480]) );
  XOR U5357 ( .A(in[855]), .B(n4003), .Z(n3535) );
  IV U5358 ( .A(n3368), .Z(n3536) );
  NANDN U5359 ( .A(n3369), .B(n3536), .Z(n3370) );
  XNOR U5360 ( .A(n3535), .B(n3370), .Z(out[481]) );
  XOR U5361 ( .A(in[856]), .B(n4007), .Z(n3768) );
  IV U5362 ( .A(n3371), .Z(n3538) );
  NANDN U5363 ( .A(n3372), .B(n3538), .Z(n3373) );
  XOR U5364 ( .A(n3768), .B(n3373), .Z(out[482]) );
  XOR U5365 ( .A(in[857]), .B(n4011), .Z(n3772) );
  IV U5366 ( .A(n3374), .Z(n3540) );
  NANDN U5367 ( .A(n3375), .B(n3540), .Z(n3376) );
  XOR U5368 ( .A(n3772), .B(n3376), .Z(out[483]) );
  XOR U5369 ( .A(in[858]), .B(n4015), .Z(n3776) );
  NANDN U5370 ( .A(n3377), .B(n3542), .Z(n3378) );
  XOR U5371 ( .A(n3776), .B(n3378), .Z(out[484]) );
  XOR U5372 ( .A(in[859]), .B(n4019), .Z(n3780) );
  NANDN U5373 ( .A(n3379), .B(n3544), .Z(n3380) );
  XOR U5374 ( .A(n3780), .B(n3380), .Z(out[485]) );
  XOR U5375 ( .A(in[860]), .B(n4023), .Z(n3550) );
  NANDN U5376 ( .A(n3381), .B(n3551), .Z(n3382) );
  XNOR U5377 ( .A(n3550), .B(n3382), .Z(out[486]) );
  XOR U5378 ( .A(in[861]), .B(n4031), .Z(n3553) );
  NANDN U5379 ( .A(n3383), .B(n3554), .Z(n3384) );
  XNOR U5380 ( .A(n3553), .B(n3384), .Z(out[487]) );
  XOR U5381 ( .A(in[862]), .B(n4035), .Z(n3556) );
  NANDN U5382 ( .A(n3385), .B(n3557), .Z(n3386) );
  XNOR U5383 ( .A(n3556), .B(n3386), .Z(out[488]) );
  XOR U5384 ( .A(in[863]), .B(n4039), .Z(n3559) );
  NANDN U5385 ( .A(n3387), .B(n3560), .Z(n3388) );
  XNOR U5386 ( .A(n3559), .B(n3388), .Z(out[489]) );
  AND U5387 ( .A(n3390), .B(n3389), .Z(n3391) );
  XNOR U5388 ( .A(n3392), .B(n3391), .Z(out[48]) );
  XOR U5389 ( .A(in[864]), .B(n4043), .Z(n3562) );
  NANDN U5390 ( .A(n3393), .B(n3563), .Z(n3394) );
  XNOR U5391 ( .A(n3562), .B(n3394), .Z(out[490]) );
  XOR U5392 ( .A(in[865]), .B(n4047), .Z(n3565) );
  NANDN U5393 ( .A(n3395), .B(n3566), .Z(n3396) );
  XNOR U5394 ( .A(n3565), .B(n3396), .Z(out[491]) );
  XNOR U5395 ( .A(n3397), .B(in[866]), .Z(n3813) );
  NANDN U5396 ( .A(n3398), .B(n3568), .Z(n3399) );
  XNOR U5397 ( .A(n3813), .B(n3399), .Z(out[492]) );
  XNOR U5398 ( .A(n3400), .B(in[867]), .Z(n3817) );
  IV U5399 ( .A(n3401), .Z(n3570) );
  NANDN U5400 ( .A(n3402), .B(n3570), .Z(n3403) );
  XNOR U5401 ( .A(n3817), .B(n3403), .Z(out[493]) );
  XNOR U5402 ( .A(n3404), .B(in[868]), .Z(n3821) );
  IV U5403 ( .A(n3405), .Z(n3572) );
  NANDN U5404 ( .A(n3406), .B(n3572), .Z(n3407) );
  XNOR U5405 ( .A(n3821), .B(n3407), .Z(out[494]) );
  XNOR U5406 ( .A(n3408), .B(in[869]), .Z(n3825) );
  IV U5407 ( .A(n3409), .Z(n3574) );
  NANDN U5408 ( .A(n3410), .B(n3574), .Z(n3411) );
  XNOR U5409 ( .A(n3825), .B(n3411), .Z(out[495]) );
  XOR U5410 ( .A(in[870]), .B(n4067), .Z(n3829) );
  IV U5411 ( .A(n3412), .Z(n3580) );
  NANDN U5412 ( .A(n3413), .B(n3580), .Z(n3414) );
  XOR U5413 ( .A(n3829), .B(n3414), .Z(out[496]) );
  XOR U5414 ( .A(in[871]), .B(n4075), .Z(n3833) );
  IV U5415 ( .A(n3415), .Z(n3582) );
  NANDN U5416 ( .A(n3416), .B(n3582), .Z(n3417) );
  XOR U5417 ( .A(n3833), .B(n3417), .Z(out[497]) );
  XOR U5418 ( .A(in[872]), .B(n4079), .Z(n3837) );
  IV U5419 ( .A(n3418), .Z(n3584) );
  NANDN U5420 ( .A(n3419), .B(n3584), .Z(n3420) );
  XOR U5421 ( .A(n3837), .B(n3420), .Z(out[498]) );
  XOR U5422 ( .A(in[873]), .B(n4083), .Z(n3841) );
  IV U5423 ( .A(n3421), .Z(n3586) );
  NANDN U5424 ( .A(n3422), .B(n3586), .Z(n3423) );
  XOR U5425 ( .A(n3841), .B(n3423), .Z(out[499]) );
  ANDN U5426 ( .B(n3425), .A(n3424), .Z(n3426) );
  XNOR U5427 ( .A(n3427), .B(n3426), .Z(out[49]) );
  OR U5428 ( .A(n4115), .B(n3428), .Z(n3429) );
  XNOR U5429 ( .A(n4114), .B(n3429), .Z(out[4]) );
  XOR U5430 ( .A(in[874]), .B(n4087), .Z(n3845) );
  NAND U5431 ( .A(n3430), .B(n3588), .Z(n3431) );
  XOR U5432 ( .A(n3845), .B(n3431), .Z(out[500]) );
  XOR U5433 ( .A(in[875]), .B(n3432), .Z(n3849) );
  NAND U5434 ( .A(n3433), .B(n3590), .Z(n3434) );
  XOR U5435 ( .A(n3849), .B(n3434), .Z(out[501]) );
  XOR U5436 ( .A(in[876]), .B(n3435), .Z(n3857) );
  NAND U5437 ( .A(n3436), .B(n3592), .Z(n3437) );
  XOR U5438 ( .A(n3857), .B(n3437), .Z(out[502]) );
  XOR U5439 ( .A(in[877]), .B(n3438), .Z(n3861) );
  NAND U5440 ( .A(n3439), .B(n3594), .Z(n3440) );
  XOR U5441 ( .A(n3861), .B(n3440), .Z(out[503]) );
  XOR U5442 ( .A(in[878]), .B(n3441), .Z(n3865) );
  NAND U5443 ( .A(n3442), .B(n3596), .Z(n3443) );
  XOR U5444 ( .A(n3865), .B(n3443), .Z(out[504]) );
  XOR U5445 ( .A(in[879]), .B(n3444), .Z(n3869) );
  NAND U5446 ( .A(n3445), .B(n3598), .Z(n3446) );
  XOR U5447 ( .A(n3869), .B(n3446), .Z(out[505]) );
  XOR U5448 ( .A(in[880]), .B(n3447), .Z(n3873) );
  NANDN U5449 ( .A(n3604), .B(n3448), .Z(n3449) );
  XOR U5450 ( .A(n3873), .B(n3449), .Z(out[506]) );
  XOR U5451 ( .A(in[881]), .B(n3450), .Z(n3877) );
  NANDN U5452 ( .A(n3605), .B(n3451), .Z(n3452) );
  XOR U5453 ( .A(n3877), .B(n3452), .Z(out[507]) );
  XOR U5454 ( .A(in[882]), .B(n3453), .Z(n3881) );
  NAND U5455 ( .A(n3454), .B(n3606), .Z(n3455) );
  XOR U5456 ( .A(n3881), .B(n3455), .Z(out[508]) );
  XOR U5457 ( .A(in[883]), .B(n3456), .Z(n3885) );
  NAND U5458 ( .A(n3457), .B(n3608), .Z(n3458) );
  XOR U5459 ( .A(n3885), .B(n3458), .Z(out[509]) );
  ANDN U5460 ( .B(n3460), .A(n3459), .Z(n3461) );
  XNOR U5461 ( .A(n3462), .B(n3461), .Z(out[50]) );
  XOR U5462 ( .A(in[884]), .B(n3463), .Z(n3889) );
  NANDN U5463 ( .A(n3464), .B(n3610), .Z(n3465) );
  XOR U5464 ( .A(n3889), .B(n3465), .Z(out[510]) );
  XOR U5465 ( .A(in[885]), .B(n3466), .Z(n3893) );
  NAND U5466 ( .A(n3467), .B(n3612), .Z(n3468) );
  XOR U5467 ( .A(n3893), .B(n3468), .Z(out[511]) );
  NANDN U5468 ( .A(n3469), .B(n3615), .Z(n3470) );
  XNOR U5469 ( .A(n3614), .B(n3470), .Z(out[512]) );
  NANDN U5470 ( .A(n3471), .B(n3619), .Z(n3472) );
  XNOR U5471 ( .A(n3618), .B(n3472), .Z(out[513]) );
  NANDN U5472 ( .A(n3473), .B(n3623), .Z(n3474) );
  XNOR U5473 ( .A(n3622), .B(n3474), .Z(out[514]) );
  NANDN U5474 ( .A(n3475), .B(n3627), .Z(n3476) );
  XNOR U5475 ( .A(n3626), .B(n3476), .Z(out[515]) );
  ANDN U5476 ( .B(n3482), .A(n3481), .Z(n3483) );
  XNOR U5477 ( .A(n3484), .B(n3483), .Z(out[51]) );
  OR U5478 ( .A(n3654), .B(n3486), .Z(n3487) );
  XOR U5479 ( .A(n3655), .B(n3487), .Z(out[521]) );
  OR U5480 ( .A(n3658), .B(n3488), .Z(n3489) );
  XOR U5481 ( .A(n3659), .B(n3489), .Z(out[522]) );
  OR U5482 ( .A(n3662), .B(n3490), .Z(n3491) );
  XOR U5483 ( .A(n3663), .B(n3491), .Z(out[523]) );
  OR U5484 ( .A(n3666), .B(n3492), .Z(n3493) );
  XOR U5485 ( .A(n3667), .B(n3493), .Z(out[524]) );
  OR U5486 ( .A(n3670), .B(n3494), .Z(n3495) );
  XOR U5487 ( .A(n3671), .B(n3495), .Z(out[525]) );
  OR U5488 ( .A(n3678), .B(n3496), .Z(n3497) );
  XOR U5489 ( .A(n3679), .B(n3497), .Z(out[526]) );
  OR U5490 ( .A(n3682), .B(n3498), .Z(n3499) );
  XOR U5491 ( .A(n3683), .B(n3499), .Z(out[527]) );
  OR U5492 ( .A(n3686), .B(n3500), .Z(n3501) );
  XOR U5493 ( .A(n3687), .B(n3501), .Z(out[528]) );
  ANDN U5494 ( .B(n3504), .A(n3503), .Z(n3505) );
  XNOR U5495 ( .A(n3506), .B(n3505), .Z(out[52]) );
  OR U5496 ( .A(n3732), .B(n3515), .Z(n3516) );
  XOR U5497 ( .A(n3733), .B(n3516), .Z(out[538]) );
  ANDN U5498 ( .B(n3519), .A(n3518), .Z(n3520) );
  XNOR U5499 ( .A(n3521), .B(n3520), .Z(out[53]) );
  OR U5500 ( .A(n3740), .B(n3522), .Z(n3523) );
  XOR U5501 ( .A(n3741), .B(n3523), .Z(out[540]) );
  IV U5502 ( .A(n3524), .Z(n3744) );
  NANDN U5503 ( .A(n3525), .B(n3744), .Z(n3526) );
  XOR U5504 ( .A(n3745), .B(n3526), .Z(out[541]) );
  IV U5505 ( .A(n3527), .Z(n3748) );
  NANDN U5506 ( .A(n3528), .B(n3748), .Z(n3529) );
  XOR U5507 ( .A(n3749), .B(n3529), .Z(out[542]) );
  IV U5508 ( .A(n3530), .Z(n3752) );
  NANDN U5509 ( .A(n3531), .B(n3752), .Z(n3532) );
  XOR U5510 ( .A(n3753), .B(n3532), .Z(out[543]) );
  NANDN U5511 ( .A(n3533), .B(n3756), .Z(n3534) );
  XOR U5512 ( .A(n3757), .B(n3534), .Z(out[544]) );
  IV U5513 ( .A(n3535), .Z(n3760) );
  NANDN U5514 ( .A(n3536), .B(n3760), .Z(n3537) );
  XOR U5515 ( .A(n3761), .B(n3537), .Z(out[545]) );
  NANDN U5516 ( .A(n3538), .B(n3768), .Z(n3539) );
  XOR U5517 ( .A(n3769), .B(n3539), .Z(out[546]) );
  NANDN U5518 ( .A(n3540), .B(n3772), .Z(n3541) );
  XOR U5519 ( .A(n3773), .B(n3541), .Z(out[547]) );
  NANDN U5520 ( .A(n3542), .B(n3776), .Z(n3543) );
  XOR U5521 ( .A(n3777), .B(n3543), .Z(out[548]) );
  NANDN U5522 ( .A(n3544), .B(n3780), .Z(n3545) );
  XOR U5523 ( .A(n3781), .B(n3545), .Z(out[549]) );
  ANDN U5524 ( .B(n3547), .A(n3546), .Z(n3548) );
  XNOR U5525 ( .A(n3549), .B(n3548), .Z(out[54]) );
  IV U5526 ( .A(n3550), .Z(n3784) );
  NANDN U5527 ( .A(n3551), .B(n3784), .Z(n3552) );
  XOR U5528 ( .A(n3785), .B(n3552), .Z(out[550]) );
  IV U5529 ( .A(n3553), .Z(n3788) );
  NANDN U5530 ( .A(n3554), .B(n3788), .Z(n3555) );
  XOR U5531 ( .A(n3789), .B(n3555), .Z(out[551]) );
  IV U5532 ( .A(n3556), .Z(n3793) );
  NANDN U5533 ( .A(n3557), .B(n3793), .Z(n3558) );
  XNOR U5534 ( .A(n3792), .B(n3558), .Z(out[552]) );
  IV U5535 ( .A(n3559), .Z(n3797) );
  NANDN U5536 ( .A(n3560), .B(n3797), .Z(n3561) );
  XNOR U5537 ( .A(n3796), .B(n3561), .Z(out[553]) );
  IV U5538 ( .A(n3562), .Z(n3801) );
  NANDN U5539 ( .A(n3563), .B(n3801), .Z(n3564) );
  XNOR U5540 ( .A(n3800), .B(n3564), .Z(out[554]) );
  IV U5541 ( .A(n3565), .Z(n3805) );
  NANDN U5542 ( .A(n3566), .B(n3805), .Z(n3567) );
  XNOR U5543 ( .A(n3804), .B(n3567), .Z(out[555]) );
  OR U5544 ( .A(n3813), .B(n3568), .Z(n3569) );
  XNOR U5545 ( .A(n3812), .B(n3569), .Z(out[556]) );
  OR U5546 ( .A(n3817), .B(n3570), .Z(n3571) );
  XNOR U5547 ( .A(n3816), .B(n3571), .Z(out[557]) );
  OR U5548 ( .A(n3821), .B(n3572), .Z(n3573) );
  XNOR U5549 ( .A(n3820), .B(n3573), .Z(out[558]) );
  OR U5550 ( .A(n3825), .B(n3574), .Z(n3575) );
  XNOR U5551 ( .A(n3824), .B(n3575), .Z(out[559]) );
  ANDN U5552 ( .B(n3577), .A(n3576), .Z(n3578) );
  XNOR U5553 ( .A(n3579), .B(n3578), .Z(out[55]) );
  NANDN U5554 ( .A(n3580), .B(n3829), .Z(n3581) );
  XNOR U5555 ( .A(n3828), .B(n3581), .Z(out[560]) );
  NANDN U5556 ( .A(n3582), .B(n3833), .Z(n3583) );
  XNOR U5557 ( .A(n3832), .B(n3583), .Z(out[561]) );
  NANDN U5558 ( .A(n3584), .B(n3837), .Z(n3585) );
  XNOR U5559 ( .A(n3836), .B(n3585), .Z(out[562]) );
  NANDN U5560 ( .A(n3586), .B(n3841), .Z(n3587) );
  XNOR U5561 ( .A(n3840), .B(n3587), .Z(out[563]) );
  NANDN U5562 ( .A(n3588), .B(n3845), .Z(n3589) );
  XNOR U5563 ( .A(n3844), .B(n3589), .Z(out[564]) );
  NANDN U5564 ( .A(n3590), .B(n3849), .Z(n3591) );
  XNOR U5565 ( .A(n3848), .B(n3591), .Z(out[565]) );
  NANDN U5566 ( .A(n3592), .B(n3857), .Z(n3593) );
  XNOR U5567 ( .A(n3856), .B(n3593), .Z(out[566]) );
  NANDN U5568 ( .A(n3594), .B(n3861), .Z(n3595) );
  XNOR U5569 ( .A(n3860), .B(n3595), .Z(out[567]) );
  NANDN U5570 ( .A(n3596), .B(n3865), .Z(n3597) );
  XNOR U5571 ( .A(n3864), .B(n3597), .Z(out[568]) );
  NANDN U5572 ( .A(n3598), .B(n3869), .Z(n3599) );
  XNOR U5573 ( .A(n3868), .B(n3599), .Z(out[569]) );
  ANDN U5574 ( .B(n3601), .A(n3600), .Z(n3602) );
  XNOR U5575 ( .A(n3603), .B(n3602), .Z(out[56]) );
  NANDN U5576 ( .A(n3606), .B(n3881), .Z(n3607) );
  XNOR U5577 ( .A(n3880), .B(n3607), .Z(out[572]) );
  NANDN U5578 ( .A(n3608), .B(n3885), .Z(n3609) );
  XNOR U5579 ( .A(n3884), .B(n3609), .Z(out[573]) );
  NANDN U5580 ( .A(n3610), .B(n3889), .Z(n3611) );
  XNOR U5581 ( .A(n3888), .B(n3611), .Z(out[574]) );
  NANDN U5582 ( .A(n3612), .B(n3893), .Z(n3613) );
  XNOR U5583 ( .A(n3892), .B(n3613), .Z(out[575]) );
  NOR U5584 ( .A(n3615), .B(n3614), .Z(n3616) );
  XOR U5585 ( .A(n3617), .B(n3616), .Z(out[576]) );
  NOR U5586 ( .A(n3619), .B(n3618), .Z(n3620) );
  XOR U5587 ( .A(n3621), .B(n3620), .Z(out[577]) );
  NOR U5588 ( .A(n3623), .B(n3622), .Z(n3624) );
  XOR U5589 ( .A(n3625), .B(n3624), .Z(out[578]) );
  NOR U5590 ( .A(n3627), .B(n3626), .Z(n3628) );
  XOR U5591 ( .A(n3629), .B(n3628), .Z(out[579]) );
  ANDN U5592 ( .B(n3631), .A(n3630), .Z(n3632) );
  XNOR U5593 ( .A(n3633), .B(n3632), .Z(out[57]) );
  NOR U5594 ( .A(n3635), .B(n3634), .Z(n3636) );
  XOR U5595 ( .A(n3637), .B(n3636), .Z(out[580]) );
  ANDN U5596 ( .B(n3639), .A(n3638), .Z(n3640) );
  XOR U5597 ( .A(n3641), .B(n3640), .Z(out[581]) );
  ANDN U5598 ( .B(n3643), .A(n3642), .Z(n3644) );
  XOR U5599 ( .A(n3645), .B(n3644), .Z(out[582]) );
  ANDN U5600 ( .B(n3647), .A(n3646), .Z(n3648) );
  XOR U5601 ( .A(n3649), .B(n3648), .Z(out[583]) );
  NOR U5602 ( .A(n3651), .B(n3650), .Z(n3652) );
  XOR U5603 ( .A(n3653), .B(n3652), .Z(out[584]) );
  AND U5604 ( .A(n3655), .B(n3654), .Z(n3656) );
  XNOR U5605 ( .A(n3657), .B(n3656), .Z(out[585]) );
  AND U5606 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U5607 ( .A(n3661), .B(n3660), .Z(out[586]) );
  AND U5608 ( .A(n3663), .B(n3662), .Z(n3664) );
  XNOR U5609 ( .A(n3665), .B(n3664), .Z(out[587]) );
  AND U5610 ( .A(n3667), .B(n3666), .Z(n3668) );
  XNOR U5611 ( .A(n3669), .B(n3668), .Z(out[588]) );
  AND U5612 ( .A(n3671), .B(n3670), .Z(n3672) );
  XNOR U5613 ( .A(n3673), .B(n3672), .Z(out[589]) );
  ANDN U5614 ( .B(n3675), .A(n3674), .Z(n3676) );
  XNOR U5615 ( .A(n3677), .B(n3676), .Z(out[58]) );
  AND U5616 ( .A(n3679), .B(n3678), .Z(n3680) );
  XNOR U5617 ( .A(n3681), .B(n3680), .Z(out[590]) );
  AND U5618 ( .A(n3683), .B(n3682), .Z(n3684) );
  XNOR U5619 ( .A(n3685), .B(n3684), .Z(out[591]) );
  AND U5620 ( .A(n3687), .B(n3686), .Z(n3688) );
  XNOR U5621 ( .A(n3689), .B(n3688), .Z(out[592]) );
  AND U5622 ( .A(n3691), .B(n3690), .Z(n3692) );
  XNOR U5623 ( .A(n3693), .B(n3692), .Z(out[593]) );
  AND U5624 ( .A(n3695), .B(n3694), .Z(n3696) );
  XNOR U5625 ( .A(n3697), .B(n3696), .Z(out[594]) );
  AND U5626 ( .A(n3699), .B(n3698), .Z(n3700) );
  XNOR U5627 ( .A(n3701), .B(n3700), .Z(out[595]) );
  AND U5628 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR U5629 ( .A(n3705), .B(n3704), .Z(out[596]) );
  AND U5630 ( .A(n3707), .B(n3706), .Z(n3708) );
  XNOR U5631 ( .A(n3709), .B(n3708), .Z(out[597]) );
  AND U5632 ( .A(n3711), .B(n3710), .Z(n3712) );
  XNOR U5633 ( .A(n3713), .B(n3712), .Z(out[598]) );
  AND U5634 ( .A(n3715), .B(n3714), .Z(n3716) );
  XNOR U5635 ( .A(n3717), .B(n3716), .Z(out[599]) );
  ANDN U5636 ( .B(n3719), .A(n3718), .Z(n3720) );
  XNOR U5637 ( .A(n3721), .B(n3720), .Z(out[59]) );
  OR U5638 ( .A(n4159), .B(n3722), .Z(n3723) );
  XNOR U5639 ( .A(n4158), .B(n3723), .Z(out[5]) );
  AND U5640 ( .A(n3725), .B(n3724), .Z(n3726) );
  XNOR U5641 ( .A(n3727), .B(n3726), .Z(out[600]) );
  AND U5642 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U5643 ( .A(n3731), .B(n3730), .Z(out[601]) );
  AND U5644 ( .A(n3733), .B(n3732), .Z(n3734) );
  XNOR U5645 ( .A(n3735), .B(n3734), .Z(out[602]) );
  AND U5646 ( .A(n3737), .B(n3736), .Z(n3738) );
  XNOR U5647 ( .A(n3739), .B(n3738), .Z(out[603]) );
  AND U5648 ( .A(n3741), .B(n3740), .Z(n3742) );
  XNOR U5649 ( .A(n3743), .B(n3742), .Z(out[604]) );
  ANDN U5650 ( .B(n3745), .A(n3744), .Z(n3746) );
  XNOR U5651 ( .A(n3747), .B(n3746), .Z(out[605]) );
  ANDN U5652 ( .B(n3749), .A(n3748), .Z(n3750) );
  XNOR U5653 ( .A(n3751), .B(n3750), .Z(out[606]) );
  ANDN U5654 ( .B(n3753), .A(n3752), .Z(n3754) );
  XNOR U5655 ( .A(n3755), .B(n3754), .Z(out[607]) );
  ANDN U5656 ( .B(n3757), .A(n3756), .Z(n3758) );
  XNOR U5657 ( .A(n3759), .B(n3758), .Z(out[608]) );
  ANDN U5658 ( .B(n3761), .A(n3760), .Z(n3762) );
  XNOR U5659 ( .A(n3763), .B(n3762), .Z(out[609]) );
  ANDN U5660 ( .B(n3765), .A(n3764), .Z(n3766) );
  XNOR U5661 ( .A(n3767), .B(n3766), .Z(out[60]) );
  ANDN U5662 ( .B(n3769), .A(n3768), .Z(n3770) );
  XNOR U5663 ( .A(n3771), .B(n3770), .Z(out[610]) );
  ANDN U5664 ( .B(n3773), .A(n3772), .Z(n3774) );
  XNOR U5665 ( .A(n3775), .B(n3774), .Z(out[611]) );
  ANDN U5666 ( .B(n3777), .A(n3776), .Z(n3778) );
  XNOR U5667 ( .A(n3779), .B(n3778), .Z(out[612]) );
  ANDN U5668 ( .B(n3781), .A(n3780), .Z(n3782) );
  XNOR U5669 ( .A(n3783), .B(n3782), .Z(out[613]) );
  ANDN U5670 ( .B(n3785), .A(n3784), .Z(n3786) );
  XNOR U5671 ( .A(n3787), .B(n3786), .Z(out[614]) );
  ANDN U5672 ( .B(n3789), .A(n3788), .Z(n3790) );
  XNOR U5673 ( .A(n3791), .B(n3790), .Z(out[615]) );
  NOR U5674 ( .A(n3793), .B(n3792), .Z(n3794) );
  XOR U5675 ( .A(n3795), .B(n3794), .Z(out[616]) );
  NOR U5676 ( .A(n3797), .B(n3796), .Z(n3798) );
  XOR U5677 ( .A(n3799), .B(n3798), .Z(out[617]) );
  NOR U5678 ( .A(n3801), .B(n3800), .Z(n3802) );
  XOR U5679 ( .A(n3803), .B(n3802), .Z(out[618]) );
  NOR U5680 ( .A(n3805), .B(n3804), .Z(n3806) );
  XOR U5681 ( .A(n3807), .B(n3806), .Z(out[619]) );
  ANDN U5682 ( .B(n3809), .A(n3808), .Z(n3810) );
  XOR U5683 ( .A(n3811), .B(n3810), .Z(out[61]) );
  ANDN U5684 ( .B(n3813), .A(n3812), .Z(n3814) );
  XOR U5685 ( .A(n3815), .B(n3814), .Z(out[620]) );
  ANDN U5686 ( .B(n3817), .A(n3816), .Z(n3818) );
  XOR U5687 ( .A(n3819), .B(n3818), .Z(out[621]) );
  ANDN U5688 ( .B(n3821), .A(n3820), .Z(n3822) );
  XOR U5689 ( .A(n3823), .B(n3822), .Z(out[622]) );
  ANDN U5690 ( .B(n3825), .A(n3824), .Z(n3826) );
  XOR U5691 ( .A(n3827), .B(n3826), .Z(out[623]) );
  NOR U5692 ( .A(n3829), .B(n3828), .Z(n3830) );
  XOR U5693 ( .A(n3831), .B(n3830), .Z(out[624]) );
  NOR U5694 ( .A(n3833), .B(n3832), .Z(n3834) );
  XOR U5695 ( .A(n3835), .B(n3834), .Z(out[625]) );
  NOR U5696 ( .A(n3837), .B(n3836), .Z(n3838) );
  XOR U5697 ( .A(n3839), .B(n3838), .Z(out[626]) );
  NOR U5698 ( .A(n3841), .B(n3840), .Z(n3842) );
  XOR U5699 ( .A(n3843), .B(n3842), .Z(out[627]) );
  NOR U5700 ( .A(n3845), .B(n3844), .Z(n3846) );
  XOR U5701 ( .A(n3847), .B(n3846), .Z(out[628]) );
  NOR U5702 ( .A(n3849), .B(n3848), .Z(n3850) );
  XOR U5703 ( .A(n3851), .B(n3850), .Z(out[629]) );
  ANDN U5704 ( .B(n3853), .A(n3852), .Z(n3854) );
  XOR U5705 ( .A(n3855), .B(n3854), .Z(out[62]) );
  NOR U5706 ( .A(n3857), .B(n3856), .Z(n3858) );
  XOR U5707 ( .A(n3859), .B(n3858), .Z(out[630]) );
  NOR U5708 ( .A(n3861), .B(n3860), .Z(n3862) );
  XOR U5709 ( .A(n3863), .B(n3862), .Z(out[631]) );
  NOR U5710 ( .A(n3865), .B(n3864), .Z(n3866) );
  XOR U5711 ( .A(n3867), .B(n3866), .Z(out[632]) );
  NOR U5712 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U5713 ( .A(n3871), .B(n3870), .Z(out[633]) );
  NOR U5714 ( .A(n3873), .B(n3872), .Z(n3874) );
  XOR U5715 ( .A(n3875), .B(n3874), .Z(out[634]) );
  NOR U5716 ( .A(n3877), .B(n3876), .Z(n3878) );
  XOR U5717 ( .A(n3879), .B(n3878), .Z(out[635]) );
  NOR U5718 ( .A(n3881), .B(n3880), .Z(n3882) );
  XOR U5719 ( .A(n3883), .B(n3882), .Z(out[636]) );
  NOR U5720 ( .A(n3885), .B(n3884), .Z(n3886) );
  XOR U5721 ( .A(n3887), .B(n3886), .Z(out[637]) );
  NOR U5722 ( .A(n3889), .B(n3888), .Z(n3890) );
  XOR U5723 ( .A(n3891), .B(n3890), .Z(out[638]) );
  NOR U5724 ( .A(n3893), .B(n3892), .Z(n3894) );
  XOR U5725 ( .A(n3895), .B(n3894), .Z(out[639]) );
  ANDN U5726 ( .B(n3897), .A(n3896), .Z(n3898) );
  XOR U5727 ( .A(n3899), .B(n3898), .Z(out[63]) );
  XOR U5728 ( .A(in[302]), .B(n3900), .Z(n4181) );
  IV U5729 ( .A(n4181), .Z(n4340) );
  XOR U5730 ( .A(in[1146]), .B(n3901), .Z(n4716) );
  XOR U5731 ( .A(in[1535]), .B(n3902), .Z(n4718) );
  OR U5732 ( .A(n4716), .B(n4718), .Z(n3903) );
  XOR U5733 ( .A(n4340), .B(n3903), .Z(out[640]) );
  XOR U5734 ( .A(in[303]), .B(n3904), .Z(n4184) );
  IV U5735 ( .A(n4184), .Z(n4342) );
  XOR U5736 ( .A(in[1147]), .B(n3905), .Z(n4720) );
  XOR U5737 ( .A(in[1472]), .B(n3906), .Z(n4722) );
  OR U5738 ( .A(n4720), .B(n4722), .Z(n3907) );
  XOR U5739 ( .A(n4342), .B(n3907), .Z(out[641]) );
  XOR U5740 ( .A(in[304]), .B(n3908), .Z(n4187) );
  IV U5741 ( .A(n4187), .Z(n4348) );
  XOR U5742 ( .A(in[1148]), .B(n3909), .Z(n4724) );
  XOR U5743 ( .A(in[1473]), .B(n3910), .Z(n4726) );
  OR U5744 ( .A(n4724), .B(n4726), .Z(n3911) );
  XOR U5745 ( .A(n4348), .B(n3911), .Z(out[642]) );
  XOR U5746 ( .A(in[305]), .B(n3912), .Z(n4190) );
  IV U5747 ( .A(n4190), .Z(n4350) );
  XOR U5748 ( .A(in[1149]), .B(n3913), .Z(n4728) );
  XOR U5749 ( .A(in[1474]), .B(n3914), .Z(n4730) );
  OR U5750 ( .A(n4728), .B(n4730), .Z(n3915) );
  XOR U5751 ( .A(n4350), .B(n3915), .Z(out[643]) );
  XOR U5752 ( .A(in[306]), .B(n3916), .Z(n4193) );
  IV U5753 ( .A(n4193), .Z(n4352) );
  XOR U5754 ( .A(in[1150]), .B(n3917), .Z(n4740) );
  XOR U5755 ( .A(in[1475]), .B(n3918), .Z(n4742) );
  OR U5756 ( .A(n4740), .B(n4742), .Z(n3919) );
  XOR U5757 ( .A(n4352), .B(n3919), .Z(out[644]) );
  XOR U5758 ( .A(in[307]), .B(n3920), .Z(n4355) );
  XOR U5759 ( .A(in[1151]), .B(n3921), .Z(n4744) );
  XOR U5760 ( .A(in[1476]), .B(n3922), .Z(n4746) );
  OR U5761 ( .A(n4744), .B(n4746), .Z(n3923) );
  XOR U5762 ( .A(n4355), .B(n3923), .Z(out[645]) );
  XOR U5763 ( .A(in[308]), .B(n3924), .Z(n4358) );
  XOR U5764 ( .A(in[1088]), .B(n3925), .Z(n4748) );
  XOR U5765 ( .A(in[1477]), .B(n3926), .Z(n4750) );
  OR U5766 ( .A(n4748), .B(n4750), .Z(n3927) );
  XOR U5767 ( .A(n4358), .B(n3927), .Z(out[646]) );
  XOR U5768 ( .A(in[309]), .B(n3928), .Z(n4361) );
  XOR U5769 ( .A(in[1089]), .B(n3929), .Z(n4752) );
  XOR U5770 ( .A(in[1478]), .B(n3930), .Z(n4754) );
  OR U5771 ( .A(n4752), .B(n4754), .Z(n3931) );
  XOR U5772 ( .A(n4361), .B(n3931), .Z(out[647]) );
  XOR U5773 ( .A(in[310]), .B(n3932), .Z(n4363) );
  XOR U5774 ( .A(in[1479]), .B(n3933), .Z(n4758) );
  XNOR U5775 ( .A(n3934), .B(in[1090]), .Z(n4755) );
  NANDN U5776 ( .A(n4758), .B(n4755), .Z(n3935) );
  XOR U5777 ( .A(n4363), .B(n3935), .Z(out[648]) );
  XOR U5778 ( .A(in[311]), .B(n3936), .Z(n4366) );
  XNOR U5779 ( .A(n3938), .B(in[1091]), .Z(n4759) );
  NANDN U5780 ( .A(n4762), .B(n4759), .Z(n3939) );
  XOR U5781 ( .A(n4366), .B(n3939), .Z(out[649]) );
  XOR U5782 ( .A(in[312]), .B(n3943), .Z(n4369) );
  XNOR U5783 ( .A(n3945), .B(in[1092]), .Z(n4763) );
  NANDN U5784 ( .A(n4766), .B(n4763), .Z(n3946) );
  XOR U5785 ( .A(n4369), .B(n3946), .Z(out[650]) );
  XOR U5786 ( .A(in[313]), .B(n3947), .Z(n4372) );
  XNOR U5787 ( .A(n3949), .B(in[1093]), .Z(n4767) );
  NANDN U5788 ( .A(n4770), .B(n4767), .Z(n3950) );
  XOR U5789 ( .A(n4372), .B(n3950), .Z(out[651]) );
  XOR U5790 ( .A(in[314]), .B(n3951), .Z(n4379) );
  XNOR U5791 ( .A(n3953), .B(in[1094]), .Z(n4771) );
  NANDN U5792 ( .A(n4774), .B(n4771), .Z(n3954) );
  XOR U5793 ( .A(n4379), .B(n3954), .Z(out[652]) );
  XOR U5794 ( .A(in[315]), .B(n3955), .Z(n4208) );
  IV U5795 ( .A(n4208), .Z(n4382) );
  XNOR U5796 ( .A(n3957), .B(in[1095]), .Z(n4775) );
  NANDN U5797 ( .A(n4778), .B(n4775), .Z(n3958) );
  XOR U5798 ( .A(n4382), .B(n3958), .Z(out[653]) );
  XOR U5799 ( .A(in[316]), .B(n3959), .Z(n4211) );
  IV U5800 ( .A(n4211), .Z(n4385) );
  XNOR U5801 ( .A(n3961), .B(in[1096]), .Z(n4782) );
  NANDN U5802 ( .A(n4785), .B(n4782), .Z(n3962) );
  XOR U5803 ( .A(n4385), .B(n3962), .Z(out[654]) );
  XOR U5804 ( .A(in[317]), .B(n3963), .Z(n4214) );
  IV U5805 ( .A(n4214), .Z(n4388) );
  XNOR U5806 ( .A(in[1097]), .B(n3965), .Z(n4786) );
  NANDN U5807 ( .A(n4789), .B(n4786), .Z(n3966) );
  XOR U5808 ( .A(n4388), .B(n3966), .Z(out[655]) );
  XOR U5809 ( .A(in[318]), .B(n3967), .Z(n4219) );
  IV U5810 ( .A(n4219), .Z(n4391) );
  XNOR U5811 ( .A(n3969), .B(in[1098]), .Z(n4790) );
  NANDN U5812 ( .A(n4793), .B(n4790), .Z(n3970) );
  XOR U5813 ( .A(n4391), .B(n3970), .Z(out[656]) );
  XOR U5814 ( .A(in[319]), .B(n3971), .Z(n4222) );
  IV U5815 ( .A(n4222), .Z(n4393) );
  XNOR U5816 ( .A(n3973), .B(in[1099]), .Z(n4794) );
  NANDN U5817 ( .A(n4797), .B(n4794), .Z(n3974) );
  XOR U5818 ( .A(n4393), .B(n3974), .Z(out[657]) );
  XOR U5819 ( .A(in[256]), .B(n3975), .Z(n4225) );
  IV U5820 ( .A(n4225), .Z(n4396) );
  XNOR U5821 ( .A(in[1100]), .B(n3977), .Z(n4798) );
  NANDN U5822 ( .A(n4801), .B(n4798), .Z(n3978) );
  XOR U5823 ( .A(n4396), .B(n3978), .Z(out[658]) );
  XOR U5824 ( .A(in[257]), .B(n3979), .Z(n4228) );
  IV U5825 ( .A(n4228), .Z(n4399) );
  XNOR U5826 ( .A(in[1101]), .B(n3981), .Z(n4802) );
  NANDN U5827 ( .A(n4805), .B(n4802), .Z(n3982) );
  XOR U5828 ( .A(n4399), .B(n3982), .Z(out[659]) );
  XOR U5829 ( .A(in[258]), .B(n3986), .Z(n4231) );
  IV U5830 ( .A(n4231), .Z(n4402) );
  XOR U5831 ( .A(in[1491]), .B(n3987), .Z(n4809) );
  XNOR U5832 ( .A(in[1102]), .B(n3988), .Z(n4806) );
  NANDN U5833 ( .A(n4809), .B(n4806), .Z(n3989) );
  XOR U5834 ( .A(n4402), .B(n3989), .Z(out[660]) );
  XOR U5835 ( .A(in[259]), .B(n3990), .Z(n4234) );
  IV U5836 ( .A(n4234), .Z(n4405) );
  XOR U5837 ( .A(in[1492]), .B(n3991), .Z(n4813) );
  XNOR U5838 ( .A(in[1103]), .B(n3992), .Z(n4810) );
  NANDN U5839 ( .A(n4813), .B(n4810), .Z(n3993) );
  XOR U5840 ( .A(n4405), .B(n3993), .Z(out[661]) );
  XOR U5841 ( .A(in[260]), .B(n3994), .Z(n4412) );
  XOR U5842 ( .A(in[1493]), .B(n3995), .Z(n4817) );
  XNOR U5843 ( .A(in[1104]), .B(n3996), .Z(n4814) );
  NANDN U5844 ( .A(n4817), .B(n4814), .Z(n3997) );
  XNOR U5845 ( .A(n4412), .B(n3997), .Z(out[662]) );
  XOR U5846 ( .A(in[261]), .B(n3998), .Z(n4415) );
  XOR U5847 ( .A(in[1494]), .B(n3999), .Z(n4238) );
  IV U5848 ( .A(n4238), .Z(n4821) );
  XNOR U5849 ( .A(in[1105]), .B(n4000), .Z(n4818) );
  NANDN U5850 ( .A(n4821), .B(n4818), .Z(n4001) );
  XNOR U5851 ( .A(n4415), .B(n4001), .Z(out[663]) );
  XOR U5852 ( .A(in[262]), .B(n4002), .Z(n4418) );
  XOR U5853 ( .A(in[1495]), .B(n4003), .Z(n4828) );
  XOR U5854 ( .A(in[1106]), .B(n4004), .Z(n4825) );
  NANDN U5855 ( .A(n4828), .B(n4825), .Z(n4005) );
  XNOR U5856 ( .A(n4418), .B(n4005), .Z(out[664]) );
  XOR U5857 ( .A(in[263]), .B(n4006), .Z(n4421) );
  XOR U5858 ( .A(in[1496]), .B(n4007), .Z(n4242) );
  IV U5859 ( .A(n4242), .Z(n4832) );
  XNOR U5860 ( .A(in[1107]), .B(n4008), .Z(n4829) );
  NANDN U5861 ( .A(n4832), .B(n4829), .Z(n4009) );
  XNOR U5862 ( .A(n4421), .B(n4009), .Z(out[665]) );
  XOR U5863 ( .A(in[264]), .B(n4010), .Z(n4424) );
  XOR U5864 ( .A(in[1497]), .B(n4011), .Z(n4247) );
  IV U5865 ( .A(n4247), .Z(n4836) );
  XNOR U5866 ( .A(in[1108]), .B(n4012), .Z(n4833) );
  NANDN U5867 ( .A(n4836), .B(n4833), .Z(n4013) );
  XNOR U5868 ( .A(n4424), .B(n4013), .Z(out[666]) );
  XOR U5869 ( .A(in[265]), .B(n4014), .Z(n4427) );
  XOR U5870 ( .A(in[1498]), .B(n4015), .Z(n4250) );
  IV U5871 ( .A(n4250), .Z(n4840) );
  XNOR U5872 ( .A(in[1109]), .B(n4016), .Z(n4837) );
  NANDN U5873 ( .A(n4840), .B(n4837), .Z(n4017) );
  XNOR U5874 ( .A(n4427), .B(n4017), .Z(out[667]) );
  XOR U5875 ( .A(in[266]), .B(n4018), .Z(n4430) );
  XOR U5876 ( .A(in[1499]), .B(n4019), .Z(n4253) );
  IV U5877 ( .A(n4253), .Z(n4844) );
  XNOR U5878 ( .A(in[1110]), .B(n4020), .Z(n4841) );
  NANDN U5879 ( .A(n4844), .B(n4841), .Z(n4021) );
  XNOR U5880 ( .A(n4430), .B(n4021), .Z(out[668]) );
  XNOR U5881 ( .A(in[267]), .B(n4022), .Z(n4433) );
  XOR U5882 ( .A(in[1500]), .B(n4023), .Z(n4848) );
  XNOR U5883 ( .A(in[1111]), .B(n4024), .Z(n4845) );
  NANDN U5884 ( .A(n4848), .B(n4845), .Z(n4025) );
  XNOR U5885 ( .A(n4433), .B(n4025), .Z(out[669]) );
  ANDN U5886 ( .B(n4027), .A(n4026), .Z(n4028) );
  XOR U5887 ( .A(n4029), .B(n4028), .Z(out[66]) );
  XOR U5888 ( .A(in[268]), .B(n4030), .Z(n4436) );
  XOR U5889 ( .A(in[1501]), .B(n4031), .Z(n4852) );
  XNOR U5890 ( .A(in[1112]), .B(n4032), .Z(n4849) );
  NANDN U5891 ( .A(n4852), .B(n4849), .Z(n4033) );
  XNOR U5892 ( .A(n4436), .B(n4033), .Z(out[670]) );
  XOR U5893 ( .A(in[269]), .B(n4034), .Z(n4439) );
  XOR U5894 ( .A(in[1502]), .B(n4035), .Z(n4856) );
  XNOR U5895 ( .A(in[1113]), .B(n4036), .Z(n4853) );
  NANDN U5896 ( .A(n4856), .B(n4853), .Z(n4037) );
  XNOR U5897 ( .A(n4439), .B(n4037), .Z(out[671]) );
  XOR U5898 ( .A(in[270]), .B(n4038), .Z(n4450) );
  XOR U5899 ( .A(in[1503]), .B(n4039), .Z(n4860) );
  XNOR U5900 ( .A(in[1114]), .B(n4040), .Z(n4857) );
  NANDN U5901 ( .A(n4860), .B(n4857), .Z(n4041) );
  XNOR U5902 ( .A(n4450), .B(n4041), .Z(out[672]) );
  XOR U5903 ( .A(in[271]), .B(n4042), .Z(n4453) );
  XOR U5904 ( .A(in[1504]), .B(n4043), .Z(n4864) );
  XNOR U5905 ( .A(in[1115]), .B(n4044), .Z(n4861) );
  NANDN U5906 ( .A(n4864), .B(n4861), .Z(n4045) );
  XNOR U5907 ( .A(n4453), .B(n4045), .Z(out[673]) );
  XOR U5908 ( .A(in[272]), .B(n4046), .Z(n4456) );
  XOR U5909 ( .A(in[1505]), .B(n4047), .Z(n4872) );
  XNOR U5910 ( .A(in[1116]), .B(n4048), .Z(n4869) );
  NANDN U5911 ( .A(n4872), .B(n4869), .Z(n4049) );
  XNOR U5912 ( .A(n4456), .B(n4049), .Z(out[674]) );
  XOR U5913 ( .A(in[273]), .B(n4050), .Z(n4459) );
  XOR U5914 ( .A(n4051), .B(in[1506]), .Z(n4876) );
  XNOR U5915 ( .A(in[1117]), .B(n4052), .Z(n4873) );
  NANDN U5916 ( .A(n4876), .B(n4873), .Z(n4053) );
  XNOR U5917 ( .A(n4459), .B(n4053), .Z(out[675]) );
  XOR U5918 ( .A(in[274]), .B(n4054), .Z(n4462) );
  XOR U5919 ( .A(n4055), .B(in[1507]), .Z(n4880) );
  XOR U5920 ( .A(in[1118]), .B(n4056), .Z(n4877) );
  NANDN U5921 ( .A(n4880), .B(n4877), .Z(n4057) );
  XNOR U5922 ( .A(n4462), .B(n4057), .Z(out[676]) );
  XOR U5923 ( .A(in[275]), .B(n4058), .Z(n4465) );
  XOR U5924 ( .A(n4059), .B(in[1508]), .Z(n4884) );
  XOR U5925 ( .A(in[1119]), .B(n4060), .Z(n4881) );
  NANDN U5926 ( .A(n4884), .B(n4881), .Z(n4061) );
  XNOR U5927 ( .A(n4465), .B(n4061), .Z(out[677]) );
  XOR U5928 ( .A(in[276]), .B(n4062), .Z(n4468) );
  XOR U5929 ( .A(n4063), .B(in[1509]), .Z(n4888) );
  XOR U5930 ( .A(in[1120]), .B(n4064), .Z(n4885) );
  NANDN U5931 ( .A(n4888), .B(n4885), .Z(n4065) );
  XNOR U5932 ( .A(n4468), .B(n4065), .Z(out[678]) );
  XOR U5933 ( .A(in[277]), .B(n4066), .Z(n4471) );
  XOR U5934 ( .A(in[1510]), .B(n4067), .Z(n4268) );
  IV U5935 ( .A(n4268), .Z(n4892) );
  XOR U5936 ( .A(in[1121]), .B(n4068), .Z(n4889) );
  NANDN U5937 ( .A(n4892), .B(n4889), .Z(n4069) );
  XNOR U5938 ( .A(n4471), .B(n4069), .Z(out[679]) );
  ANDN U5939 ( .B(n4071), .A(n4070), .Z(n4072) );
  XOR U5940 ( .A(n4073), .B(n4072), .Z(out[67]) );
  XOR U5941 ( .A(in[278]), .B(n4074), .Z(n4474) );
  XOR U5942 ( .A(in[1511]), .B(n4075), .Z(n4271) );
  IV U5943 ( .A(n4271), .Z(n4896) );
  XOR U5944 ( .A(in[1122]), .B(n4076), .Z(n4893) );
  NANDN U5945 ( .A(n4896), .B(n4893), .Z(n4077) );
  XNOR U5946 ( .A(n4474), .B(n4077), .Z(out[680]) );
  XOR U5947 ( .A(in[279]), .B(n4078), .Z(n4477) );
  XOR U5948 ( .A(in[1512]), .B(n4079), .Z(n4274) );
  IV U5949 ( .A(n4274), .Z(n4900) );
  XOR U5950 ( .A(in[1123]), .B(n4080), .Z(n4897) );
  NANDN U5951 ( .A(n4900), .B(n4897), .Z(n4081) );
  XNOR U5952 ( .A(n4477), .B(n4081), .Z(out[681]) );
  XOR U5953 ( .A(in[280]), .B(n4082), .Z(n4484) );
  XOR U5954 ( .A(in[1513]), .B(n4083), .Z(n4277) );
  IV U5955 ( .A(n4277), .Z(n4904) );
  XOR U5956 ( .A(in[1124]), .B(n4084), .Z(n4901) );
  NANDN U5957 ( .A(n4904), .B(n4901), .Z(n4085) );
  XNOR U5958 ( .A(n4484), .B(n4085), .Z(out[682]) );
  XOR U5959 ( .A(in[281]), .B(n4086), .Z(n4487) );
  XOR U5960 ( .A(in[1514]), .B(n4087), .Z(n4280) );
  IV U5961 ( .A(n4280), .Z(n4908) );
  XNOR U5962 ( .A(in[1125]), .B(n4088), .Z(n4905) );
  NANDN U5963 ( .A(n4908), .B(n4905), .Z(n4089) );
  XNOR U5964 ( .A(n4487), .B(n4089), .Z(out[683]) );
  XOR U5965 ( .A(in[282]), .B(n4090), .Z(n4490) );
  XOR U5966 ( .A(in[1126]), .B(n4091), .Z(n4914) );
  XNOR U5967 ( .A(in[1515]), .B(n4092), .Z(n4916) );
  NANDN U5968 ( .A(n4914), .B(n4916), .Z(n4093) );
  XNOR U5969 ( .A(n4490), .B(n4093), .Z(out[684]) );
  XOR U5970 ( .A(in[283]), .B(n4094), .Z(n4493) );
  XOR U5971 ( .A(in[1127]), .B(n4095), .Z(n4918) );
  XNOR U5972 ( .A(in[1516]), .B(n4096), .Z(n4920) );
  NANDN U5973 ( .A(n4918), .B(n4920), .Z(n4097) );
  XNOR U5974 ( .A(n4493), .B(n4097), .Z(out[685]) );
  XOR U5975 ( .A(in[284]), .B(n4098), .Z(n4496) );
  XOR U5976 ( .A(in[1128]), .B(n4099), .Z(n4922) );
  XNOR U5977 ( .A(in[1517]), .B(n4100), .Z(n4924) );
  NANDN U5978 ( .A(n4922), .B(n4924), .Z(n4101) );
  XNOR U5979 ( .A(n4496), .B(n4101), .Z(out[686]) );
  XOR U5980 ( .A(in[285]), .B(n4102), .Z(n4499) );
  XOR U5981 ( .A(in[1129]), .B(n4103), .Z(n4926) );
  XNOR U5982 ( .A(in[1518]), .B(n4104), .Z(n4928) );
  NANDN U5983 ( .A(n4926), .B(n4928), .Z(n4105) );
  XNOR U5984 ( .A(n4499), .B(n4105), .Z(out[687]) );
  XOR U5985 ( .A(in[286]), .B(n4106), .Z(n4502) );
  XOR U5986 ( .A(in[1130]), .B(n4107), .Z(n4930) );
  XNOR U5987 ( .A(in[1519]), .B(n4108), .Z(n4932) );
  NANDN U5988 ( .A(n4930), .B(n4932), .Z(n4109) );
  XNOR U5989 ( .A(n4502), .B(n4109), .Z(out[688]) );
  XOR U5990 ( .A(in[287]), .B(n4110), .Z(n4505) );
  XNOR U5991 ( .A(in[1131]), .B(n4111), .Z(n4934) );
  XNOR U5992 ( .A(in[1520]), .B(n4112), .Z(n4936) );
  NANDN U5993 ( .A(n4934), .B(n4936), .Z(n4113) );
  XNOR U5994 ( .A(n4505), .B(n4113), .Z(out[689]) );
  ANDN U5995 ( .B(n4115), .A(n4114), .Z(n4116) );
  XOR U5996 ( .A(n4117), .B(n4116), .Z(out[68]) );
  XOR U5997 ( .A(in[288]), .B(n4118), .Z(n4508) );
  XNOR U5998 ( .A(in[1132]), .B(n4119), .Z(n4938) );
  XNOR U5999 ( .A(in[1521]), .B(n4120), .Z(n4940) );
  NANDN U6000 ( .A(n4938), .B(n4940), .Z(n4121) );
  XNOR U6001 ( .A(n4508), .B(n4121), .Z(out[690]) );
  XOR U6002 ( .A(in[289]), .B(n4122), .Z(n4511) );
  XOR U6003 ( .A(in[1133]), .B(n4123), .Z(n4942) );
  XNOR U6004 ( .A(in[1522]), .B(n4124), .Z(n4944) );
  NANDN U6005 ( .A(n4942), .B(n4944), .Z(n4125) );
  XNOR U6006 ( .A(n4511), .B(n4125), .Z(out[691]) );
  XOR U6007 ( .A(in[290]), .B(n4126), .Z(n4518) );
  XOR U6008 ( .A(in[1134]), .B(n4127), .Z(n4946) );
  XNOR U6009 ( .A(in[1523]), .B(n4128), .Z(n4948) );
  NANDN U6010 ( .A(n4946), .B(n4948), .Z(n4129) );
  XNOR U6011 ( .A(n4518), .B(n4129), .Z(out[692]) );
  XOR U6012 ( .A(in[291]), .B(n4130), .Z(n4521) );
  XOR U6013 ( .A(in[1135]), .B(n4131), .Z(n4950) );
  XNOR U6014 ( .A(in[1524]), .B(n4132), .Z(n4952) );
  NANDN U6015 ( .A(n4950), .B(n4952), .Z(n4133) );
  XNOR U6016 ( .A(n4521), .B(n4133), .Z(out[693]) );
  XOR U6017 ( .A(in[292]), .B(n4134), .Z(n4524) );
  XOR U6018 ( .A(in[1136]), .B(n4135), .Z(n4958) );
  XNOR U6019 ( .A(in[1525]), .B(n4136), .Z(n4960) );
  NANDN U6020 ( .A(n4958), .B(n4960), .Z(n4137) );
  XNOR U6021 ( .A(n4524), .B(n4137), .Z(out[694]) );
  XOR U6022 ( .A(in[293]), .B(n4138), .Z(n4309) );
  IV U6023 ( .A(n4309), .Z(n4528) );
  XOR U6024 ( .A(in[1137]), .B(n4139), .Z(n4962) );
  XNOR U6025 ( .A(in[1526]), .B(n4140), .Z(n4964) );
  NANDN U6026 ( .A(n4962), .B(n4964), .Z(n4141) );
  XOR U6027 ( .A(n4528), .B(n4141), .Z(out[695]) );
  XOR U6028 ( .A(in[294]), .B(n4142), .Z(n4316) );
  IV U6029 ( .A(n4316), .Z(n4532) );
  XOR U6030 ( .A(in[1138]), .B(n4143), .Z(n4966) );
  XNOR U6031 ( .A(in[1527]), .B(n4144), .Z(n4968) );
  NANDN U6032 ( .A(n4966), .B(n4968), .Z(n4145) );
  XOR U6033 ( .A(n4532), .B(n4145), .Z(out[696]) );
  XOR U6034 ( .A(in[295]), .B(n4146), .Z(n4319) );
  IV U6035 ( .A(n4319), .Z(n4536) );
  XOR U6036 ( .A(in[1139]), .B(n4147), .Z(n4970) );
  XNOR U6037 ( .A(in[1528]), .B(n4148), .Z(n4972) );
  NANDN U6038 ( .A(n4970), .B(n4972), .Z(n4149) );
  XOR U6039 ( .A(n4536), .B(n4149), .Z(out[697]) );
  XOR U6040 ( .A(in[296]), .B(n4150), .Z(n4322) );
  IV U6041 ( .A(n4322), .Z(n4540) );
  XOR U6042 ( .A(in[1140]), .B(n4151), .Z(n4974) );
  XNOR U6043 ( .A(in[1529]), .B(n4152), .Z(n4976) );
  NANDN U6044 ( .A(n4974), .B(n4976), .Z(n4153) );
  XOR U6045 ( .A(n4540), .B(n4153), .Z(out[698]) );
  XOR U6046 ( .A(in[297]), .B(n4154), .Z(n4325) );
  IV U6047 ( .A(n4325), .Z(n4544) );
  XNOR U6048 ( .A(in[1141]), .B(n4155), .Z(n4978) );
  XNOR U6049 ( .A(in[1530]), .B(n4156), .Z(n4980) );
  NANDN U6050 ( .A(n4978), .B(n4980), .Z(n4157) );
  XOR U6051 ( .A(n4544), .B(n4157), .Z(out[699]) );
  ANDN U6052 ( .B(n4159), .A(n4158), .Z(n4160) );
  XOR U6053 ( .A(n4161), .B(n4160), .Z(out[69]) );
  OR U6054 ( .A(n4197), .B(n4162), .Z(n4163) );
  XNOR U6055 ( .A(n4196), .B(n4163), .Z(out[6]) );
  XOR U6056 ( .A(in[298]), .B(n4164), .Z(n4328) );
  IV U6057 ( .A(n4328), .Z(n4548) );
  XNOR U6058 ( .A(in[1142]), .B(n4165), .Z(n4982) );
  XNOR U6059 ( .A(in[1531]), .B(n4166), .Z(n4984) );
  OR U6060 ( .A(n4982), .B(n4984), .Z(n4167) );
  XOR U6061 ( .A(n4548), .B(n4167), .Z(out[700]) );
  XOR U6062 ( .A(in[299]), .B(n4168), .Z(n4331) );
  IV U6063 ( .A(n4331), .Z(n4551) );
  XNOR U6064 ( .A(in[1143]), .B(n4169), .Z(n4986) );
  XNOR U6065 ( .A(in[1532]), .B(n4170), .Z(n4988) );
  OR U6066 ( .A(n4986), .B(n4988), .Z(n4171) );
  XOR U6067 ( .A(n4551), .B(n4171), .Z(out[701]) );
  XOR U6068 ( .A(in[300]), .B(n4172), .Z(n4334) );
  IV U6069 ( .A(n4334), .Z(n4557) );
  XNOR U6070 ( .A(in[1144]), .B(n4173), .Z(n4990) );
  XNOR U6071 ( .A(in[1533]), .B(n4174), .Z(n4992) );
  OR U6072 ( .A(n4990), .B(n4992), .Z(n4175) );
  XOR U6073 ( .A(n4557), .B(n4175), .Z(out[702]) );
  XOR U6074 ( .A(in[301]), .B(n4176), .Z(n4337) );
  IV U6075 ( .A(n4337), .Z(n4559) );
  XNOR U6076 ( .A(in[1145]), .B(n4177), .Z(n4994) );
  XNOR U6077 ( .A(in[1534]), .B(n4178), .Z(n4996) );
  NANDN U6078 ( .A(n4994), .B(n4996), .Z(n4179) );
  XOR U6079 ( .A(n4559), .B(n4179), .Z(out[703]) );
  XOR U6080 ( .A(in[376]), .B(n4180), .Z(n4560) );
  ANDN U6081 ( .B(n4718), .A(n4181), .Z(n4182) );
  XOR U6082 ( .A(n4560), .B(n4182), .Z(out[704]) );
  XOR U6083 ( .A(in[377]), .B(n4183), .Z(n4563) );
  ANDN U6084 ( .B(n4722), .A(n4184), .Z(n4185) );
  XOR U6085 ( .A(n4563), .B(n4185), .Z(out[705]) );
  XOR U6086 ( .A(in[378]), .B(n4186), .Z(n4566) );
  ANDN U6087 ( .B(n4726), .A(n4187), .Z(n4188) );
  XOR U6088 ( .A(n4566), .B(n4188), .Z(out[706]) );
  XOR U6089 ( .A(in[379]), .B(n4189), .Z(n4569) );
  ANDN U6090 ( .B(n4730), .A(n4190), .Z(n4191) );
  XOR U6091 ( .A(n4569), .B(n4191), .Z(out[707]) );
  XOR U6092 ( .A(in[380]), .B(n4192), .Z(n4572) );
  ANDN U6093 ( .B(n4742), .A(n4193), .Z(n4194) );
  XNOR U6094 ( .A(n4572), .B(n4194), .Z(out[708]) );
  XOR U6095 ( .A(in[381]), .B(n4195), .Z(n4574) );
  ANDN U6096 ( .B(n4197), .A(n4196), .Z(n4198) );
  XOR U6097 ( .A(n4199), .B(n4198), .Z(out[70]) );
  XOR U6098 ( .A(in[382]), .B(n4200), .Z(n4576) );
  XOR U6099 ( .A(in[383]), .B(n4201), .Z(n4578) );
  XOR U6100 ( .A(in[320]), .B(n4202), .Z(n4585) );
  XOR U6101 ( .A(in[321]), .B(n4203), .Z(n4587) );
  XOR U6102 ( .A(in[322]), .B(n4204), .Z(n4589) );
  XOR U6103 ( .A(in[323]), .B(n4205), .Z(n4591) );
  XOR U6104 ( .A(in[324]), .B(n4206), .Z(n4593) );
  XOR U6105 ( .A(in[325]), .B(n4207), .Z(n4595) );
  ANDN U6106 ( .B(n4778), .A(n4208), .Z(n4209) );
  XNOR U6107 ( .A(n4595), .B(n4209), .Z(out[717]) );
  XOR U6108 ( .A(in[326]), .B(n4210), .Z(n4597) );
  ANDN U6109 ( .B(n4785), .A(n4211), .Z(n4212) );
  XNOR U6110 ( .A(n4597), .B(n4212), .Z(out[718]) );
  XOR U6111 ( .A(in[327]), .B(n4213), .Z(n4599) );
  ANDN U6112 ( .B(n4789), .A(n4214), .Z(n4215) );
  XNOR U6113 ( .A(n4599), .B(n4215), .Z(out[719]) );
  ANDN U6114 ( .B(n4446), .A(n4448), .Z(n4216) );
  XOR U6115 ( .A(n4217), .B(n4216), .Z(out[71]) );
  XOR U6116 ( .A(in[328]), .B(n4218), .Z(n4601) );
  ANDN U6117 ( .B(n4793), .A(n4219), .Z(n4220) );
  XOR U6118 ( .A(n4601), .B(n4220), .Z(out[720]) );
  XOR U6119 ( .A(in[329]), .B(n4221), .Z(n4604) );
  ANDN U6120 ( .B(n4797), .A(n4222), .Z(n4223) );
  XNOR U6121 ( .A(n4604), .B(n4223), .Z(out[721]) );
  XOR U6122 ( .A(in[330]), .B(n4224), .Z(n4610) );
  ANDN U6123 ( .B(n4801), .A(n4225), .Z(n4226) );
  XNOR U6124 ( .A(n4610), .B(n4226), .Z(out[722]) );
  XOR U6125 ( .A(in[331]), .B(n4227), .Z(n4612) );
  ANDN U6126 ( .B(n4805), .A(n4228), .Z(n4229) );
  XNOR U6127 ( .A(n4612), .B(n4229), .Z(out[723]) );
  XOR U6128 ( .A(in[332]), .B(n4230), .Z(n4614) );
  ANDN U6129 ( .B(n4809), .A(n4231), .Z(n4232) );
  XNOR U6130 ( .A(n4614), .B(n4232), .Z(out[724]) );
  XOR U6131 ( .A(in[333]), .B(n4233), .Z(n4616) );
  ANDN U6132 ( .B(n4813), .A(n4234), .Z(n4235) );
  XNOR U6133 ( .A(n4616), .B(n4235), .Z(out[725]) );
  XOR U6134 ( .A(in[334]), .B(n4236), .Z(n4618) );
  XOR U6135 ( .A(in[335]), .B(n4237), .Z(n4620) );
  NOR U6136 ( .A(n4238), .B(n4415), .Z(n4239) );
  XOR U6137 ( .A(n4620), .B(n4239), .Z(out[727]) );
  XOR U6138 ( .A(in[336]), .B(n4240), .Z(n4623) );
  XOR U6139 ( .A(in[337]), .B(n4241), .Z(n4626) );
  NOR U6140 ( .A(n4242), .B(n4421), .Z(n4243) );
  XOR U6141 ( .A(n4626), .B(n4243), .Z(out[729]) );
  ANDN U6142 ( .B(n4736), .A(n4738), .Z(n4244) );
  XOR U6143 ( .A(n4245), .B(n4244), .Z(out[72]) );
  XOR U6144 ( .A(in[338]), .B(n4246), .Z(n4629) );
  NOR U6145 ( .A(n4247), .B(n4424), .Z(n4248) );
  XOR U6146 ( .A(n4629), .B(n4248), .Z(out[730]) );
  XOR U6147 ( .A(in[339]), .B(n4249), .Z(n4632) );
  NOR U6148 ( .A(n4250), .B(n4427), .Z(n4251) );
  XOR U6149 ( .A(n4632), .B(n4251), .Z(out[731]) );
  XOR U6150 ( .A(in[340]), .B(n4252), .Z(n4639) );
  NOR U6151 ( .A(n4253), .B(n4430), .Z(n4254) );
  XOR U6152 ( .A(n4639), .B(n4254), .Z(out[732]) );
  XOR U6153 ( .A(in[341]), .B(n4255), .Z(n4642) );
  XOR U6154 ( .A(in[342]), .B(n4256), .Z(n4645) );
  XOR U6155 ( .A(in[343]), .B(n4257), .Z(n4648) );
  XOR U6156 ( .A(in[344]), .B(n4258), .Z(n4649) );
  XOR U6157 ( .A(in[345]), .B(n4259), .Z(n4652) );
  XOR U6158 ( .A(in[346]), .B(n4260), .Z(n4655) );
  XOR U6159 ( .A(in[347]), .B(n4261), .Z(n4658) );
  ANDN U6160 ( .B(n5165), .A(n5167), .Z(n4262) );
  XOR U6161 ( .A(n4263), .B(n4262), .Z(out[73]) );
  XOR U6162 ( .A(in[348]), .B(n4264), .Z(n4661) );
  XOR U6163 ( .A(in[349]), .B(n4265), .Z(n4664) );
  XOR U6164 ( .A(in[350]), .B(n4266), .Z(n4669) );
  XOR U6165 ( .A(in[351]), .B(n4267), .Z(n4670) );
  NOR U6166 ( .A(n4268), .B(n4471), .Z(n4269) );
  XOR U6167 ( .A(n4670), .B(n4269), .Z(out[743]) );
  XOR U6168 ( .A(in[352]), .B(n4270), .Z(n4671) );
  NOR U6169 ( .A(n4271), .B(n4474), .Z(n4272) );
  XOR U6170 ( .A(n4671), .B(n4272), .Z(out[744]) );
  XOR U6171 ( .A(in[353]), .B(n4273), .Z(n4672) );
  NOR U6172 ( .A(n4274), .B(n4477), .Z(n4275) );
  XOR U6173 ( .A(n4672), .B(n4275), .Z(out[745]) );
  XOR U6174 ( .A(in[354]), .B(n4276), .Z(n4673) );
  NOR U6175 ( .A(n4277), .B(n4484), .Z(n4278) );
  XOR U6176 ( .A(n4673), .B(n4278), .Z(out[746]) );
  XOR U6177 ( .A(in[355]), .B(n4279), .Z(n4674) );
  NOR U6178 ( .A(n4280), .B(n4487), .Z(n4281) );
  XNOR U6179 ( .A(n4674), .B(n4281), .Z(out[747]) );
  XOR U6180 ( .A(in[356]), .B(n4282), .Z(n4676) );
  NOR U6181 ( .A(n4916), .B(n4490), .Z(n4283) );
  XOR U6182 ( .A(n4676), .B(n4283), .Z(out[748]) );
  XOR U6183 ( .A(in[357]), .B(n4284), .Z(n4677) );
  NOR U6184 ( .A(n4920), .B(n4493), .Z(n4285) );
  XOR U6185 ( .A(n4677), .B(n4285), .Z(out[749]) );
  ANDN U6186 ( .B(n4287), .A(n4286), .Z(n4288) );
  XOR U6187 ( .A(n4289), .B(n4288), .Z(out[74]) );
  XOR U6188 ( .A(in[358]), .B(n4290), .Z(n4678) );
  NOR U6189 ( .A(n4924), .B(n4496), .Z(n4291) );
  XOR U6190 ( .A(n4678), .B(n4291), .Z(out[750]) );
  XOR U6191 ( .A(in[359]), .B(n4292), .Z(n4679) );
  NOR U6192 ( .A(n4928), .B(n4499), .Z(n4293) );
  XOR U6193 ( .A(n4679), .B(n4293), .Z(out[751]) );
  XOR U6194 ( .A(in[360]), .B(n4294), .Z(n4684) );
  NOR U6195 ( .A(n4932), .B(n4502), .Z(n4295) );
  XOR U6196 ( .A(n4684), .B(n4295), .Z(out[752]) );
  XOR U6197 ( .A(in[361]), .B(n4296), .Z(n4685) );
  NOR U6198 ( .A(n4936), .B(n4505), .Z(n4297) );
  XOR U6199 ( .A(n4685), .B(n4297), .Z(out[753]) );
  XOR U6200 ( .A(in[362]), .B(n4298), .Z(n4686) );
  NOR U6201 ( .A(n4940), .B(n4508), .Z(n4299) );
  XOR U6202 ( .A(n4686), .B(n4299), .Z(out[754]) );
  XOR U6203 ( .A(in[363]), .B(n4300), .Z(n4687) );
  NOR U6204 ( .A(n4944), .B(n4511), .Z(n4301) );
  XOR U6205 ( .A(n4687), .B(n4301), .Z(out[755]) );
  XOR U6206 ( .A(in[364]), .B(n4302), .Z(n4688) );
  NOR U6207 ( .A(n4948), .B(n4518), .Z(n4303) );
  XOR U6208 ( .A(n4688), .B(n4303), .Z(out[756]) );
  XOR U6209 ( .A(in[365]), .B(n4304), .Z(n4689) );
  NOR U6210 ( .A(n4952), .B(n4521), .Z(n4305) );
  XOR U6211 ( .A(n4689), .B(n4305), .Z(out[757]) );
  XOR U6212 ( .A(in[366]), .B(n4306), .Z(n4690) );
  NOR U6213 ( .A(n4960), .B(n4524), .Z(n4307) );
  XOR U6214 ( .A(n4690), .B(n4307), .Z(out[758]) );
  XOR U6215 ( .A(in[367]), .B(n4308), .Z(n4527) );
  NOR U6216 ( .A(n4309), .B(n4964), .Z(n4310) );
  XOR U6217 ( .A(n4527), .B(n4310), .Z(out[759]) );
  ANDN U6218 ( .B(n4312), .A(n4311), .Z(n4313) );
  XOR U6219 ( .A(n4314), .B(n4313), .Z(out[75]) );
  XOR U6220 ( .A(in[368]), .B(n4315), .Z(n4531) );
  NOR U6221 ( .A(n4316), .B(n4968), .Z(n4317) );
  XOR U6222 ( .A(n4531), .B(n4317), .Z(out[760]) );
  XOR U6223 ( .A(in[369]), .B(n4318), .Z(n4535) );
  NOR U6224 ( .A(n4319), .B(n4972), .Z(n4320) );
  XOR U6225 ( .A(n4535), .B(n4320), .Z(out[761]) );
  XOR U6226 ( .A(in[370]), .B(n4321), .Z(n4539) );
  NOR U6227 ( .A(n4322), .B(n4976), .Z(n4323) );
  XOR U6228 ( .A(n4539), .B(n4323), .Z(out[762]) );
  XOR U6229 ( .A(in[371]), .B(n4324), .Z(n4543) );
  NOR U6230 ( .A(n4325), .B(n4980), .Z(n4326) );
  XOR U6231 ( .A(n4543), .B(n4326), .Z(out[763]) );
  XOR U6232 ( .A(in[372]), .B(n4327), .Z(n4547) );
  ANDN U6233 ( .B(n4984), .A(n4328), .Z(n4329) );
  XOR U6234 ( .A(n4547), .B(n4329), .Z(out[764]) );
  XOR U6235 ( .A(in[373]), .B(n4330), .Z(n4706) );
  ANDN U6236 ( .B(n4988), .A(n4331), .Z(n4332) );
  XOR U6237 ( .A(n4706), .B(n4332), .Z(out[765]) );
  XOR U6238 ( .A(in[374]), .B(n4333), .Z(n4709) );
  ANDN U6239 ( .B(n4992), .A(n4334), .Z(n4335) );
  XOR U6240 ( .A(n4709), .B(n4335), .Z(out[766]) );
  XOR U6241 ( .A(in[375]), .B(n4336), .Z(n4712) );
  NOR U6242 ( .A(n4337), .B(n4996), .Z(n4338) );
  XOR U6243 ( .A(n4712), .B(n4338), .Z(out[767]) );
  XOR U6244 ( .A(in[743]), .B(n4339), .Z(n4561) );
  IV U6245 ( .A(n4561), .Z(n4715) );
  XOR U6246 ( .A(in[744]), .B(n4341), .Z(n4564) );
  IV U6247 ( .A(n4564), .Z(n4719) );
  ANDN U6248 ( .B(n4344), .A(n4343), .Z(n4345) );
  XOR U6249 ( .A(n4346), .B(n4345), .Z(out[76]) );
  XOR U6250 ( .A(in[745]), .B(n4347), .Z(n4567) );
  IV U6251 ( .A(n4567), .Z(n4723) );
  XOR U6252 ( .A(in[746]), .B(n4349), .Z(n4570) );
  IV U6253 ( .A(n4570), .Z(n4727) );
  XNOR U6254 ( .A(in[747]), .B(n4351), .Z(n4739) );
  NANDN U6255 ( .A(n4352), .B(n4572), .Z(n4353) );
  XOR U6256 ( .A(n4739), .B(n4353), .Z(out[772]) );
  XNOR U6257 ( .A(in[748]), .B(n4354), .Z(n4743) );
  NANDN U6258 ( .A(n4355), .B(n4574), .Z(n4356) );
  XOR U6259 ( .A(n4743), .B(n4356), .Z(out[773]) );
  XNOR U6260 ( .A(in[749]), .B(n4357), .Z(n4747) );
  NANDN U6261 ( .A(n4358), .B(n4576), .Z(n4359) );
  XOR U6262 ( .A(n4747), .B(n4359), .Z(out[774]) );
  XOR U6263 ( .A(in[750]), .B(n4360), .Z(n4579) );
  IV U6264 ( .A(n4579), .Z(n4751) );
  XNOR U6265 ( .A(in[751]), .B(n4362), .Z(n4756) );
  NANDN U6266 ( .A(n4363), .B(n4585), .Z(n4364) );
  XOR U6267 ( .A(n4756), .B(n4364), .Z(out[776]) );
  XNOR U6268 ( .A(in[752]), .B(n4365), .Z(n4760) );
  NANDN U6269 ( .A(n4366), .B(n4587), .Z(n4367) );
  XOR U6270 ( .A(n4760), .B(n4367), .Z(out[777]) );
  XNOR U6271 ( .A(in[753]), .B(n4368), .Z(n4764) );
  NANDN U6272 ( .A(n4369), .B(n4589), .Z(n4370) );
  XOR U6273 ( .A(n4764), .B(n4370), .Z(out[778]) );
  XNOR U6274 ( .A(in[754]), .B(n4371), .Z(n4768) );
  NANDN U6275 ( .A(n4372), .B(n4591), .Z(n4373) );
  XOR U6276 ( .A(n4768), .B(n4373), .Z(out[779]) );
  ANDN U6277 ( .B(n4375), .A(n4374), .Z(n4376) );
  XOR U6278 ( .A(n4377), .B(n4376), .Z(out[77]) );
  XNOR U6279 ( .A(in[755]), .B(n4378), .Z(n4772) );
  NANDN U6280 ( .A(n4379), .B(n4593), .Z(n4380) );
  XOR U6281 ( .A(n4772), .B(n4380), .Z(out[780]) );
  XNOR U6282 ( .A(in[756]), .B(n4381), .Z(n4776) );
  NANDN U6283 ( .A(n4382), .B(n4595), .Z(n4383) );
  XOR U6284 ( .A(n4776), .B(n4383), .Z(out[781]) );
  XNOR U6285 ( .A(in[757]), .B(n4384), .Z(n4783) );
  NANDN U6286 ( .A(n4385), .B(n4597), .Z(n4386) );
  XOR U6287 ( .A(n4783), .B(n4386), .Z(out[782]) );
  XNOR U6288 ( .A(in[758]), .B(n4387), .Z(n4787) );
  NANDN U6289 ( .A(n4388), .B(n4599), .Z(n4389) );
  XOR U6290 ( .A(n4787), .B(n4389), .Z(out[783]) );
  XOR U6291 ( .A(in[759]), .B(n4390), .Z(n4602) );
  IV U6292 ( .A(n4602), .Z(n4791) );
  XNOR U6293 ( .A(in[760]), .B(n4392), .Z(n4795) );
  NANDN U6294 ( .A(n4393), .B(n4604), .Z(n4394) );
  XOR U6295 ( .A(n4795), .B(n4394), .Z(out[785]) );
  XNOR U6296 ( .A(in[761]), .B(n4395), .Z(n4799) );
  NANDN U6297 ( .A(n4396), .B(n4610), .Z(n4397) );
  XOR U6298 ( .A(n4799), .B(n4397), .Z(out[786]) );
  XOR U6299 ( .A(in[762]), .B(n4398), .Z(n4803) );
  NANDN U6300 ( .A(n4399), .B(n4612), .Z(n4400) );
  XOR U6301 ( .A(n4803), .B(n4400), .Z(out[787]) );
  XOR U6302 ( .A(in[763]), .B(n4401), .Z(n4807) );
  NANDN U6303 ( .A(n4402), .B(n4614), .Z(n4403) );
  XOR U6304 ( .A(n4807), .B(n4403), .Z(out[788]) );
  XNOR U6305 ( .A(in[764]), .B(n4404), .Z(n4811) );
  NANDN U6306 ( .A(n4405), .B(n4616), .Z(n4406) );
  XOR U6307 ( .A(n4811), .B(n4406), .Z(out[789]) );
  ANDN U6308 ( .B(n4408), .A(n4407), .Z(n4409) );
  XOR U6309 ( .A(n4410), .B(n4409), .Z(out[78]) );
  XNOR U6310 ( .A(in[765]), .B(n4411), .Z(n4815) );
  NAND U6311 ( .A(n4412), .B(n4618), .Z(n4413) );
  XOR U6312 ( .A(n4815), .B(n4413), .Z(out[790]) );
  XOR U6313 ( .A(in[766]), .B(n4414), .Z(n4621) );
  IV U6314 ( .A(n4621), .Z(n4819) );
  NANDN U6315 ( .A(n4620), .B(n4415), .Z(n4416) );
  XOR U6316 ( .A(n4819), .B(n4416), .Z(out[791]) );
  XOR U6317 ( .A(in[767]), .B(n4417), .Z(n4624) );
  IV U6318 ( .A(n4624), .Z(n4826) );
  NANDN U6319 ( .A(n4623), .B(n4418), .Z(n4419) );
  XOR U6320 ( .A(n4826), .B(n4419), .Z(out[792]) );
  XOR U6321 ( .A(in[704]), .B(n4420), .Z(n4627) );
  IV U6322 ( .A(n4627), .Z(n4830) );
  NANDN U6323 ( .A(n4626), .B(n4421), .Z(n4422) );
  XOR U6324 ( .A(n4830), .B(n4422), .Z(out[793]) );
  XOR U6325 ( .A(in[705]), .B(n4423), .Z(n4630) );
  IV U6326 ( .A(n4630), .Z(n4834) );
  NANDN U6327 ( .A(n4629), .B(n4424), .Z(n4425) );
  XOR U6328 ( .A(n4834), .B(n4425), .Z(out[794]) );
  XOR U6329 ( .A(in[706]), .B(n4426), .Z(n4633) );
  IV U6330 ( .A(n4633), .Z(n4838) );
  NANDN U6331 ( .A(n4632), .B(n4427), .Z(n4428) );
  XOR U6332 ( .A(n4838), .B(n4428), .Z(out[795]) );
  XOR U6333 ( .A(in[707]), .B(n4429), .Z(n4640) );
  IV U6334 ( .A(n4640), .Z(n4842) );
  NANDN U6335 ( .A(n4639), .B(n4430), .Z(n4431) );
  XOR U6336 ( .A(n4842), .B(n4431), .Z(out[796]) );
  XOR U6337 ( .A(in[708]), .B(n4432), .Z(n4643) );
  IV U6338 ( .A(n4643), .Z(n4846) );
  NANDN U6339 ( .A(n4642), .B(n4433), .Z(n4434) );
  XOR U6340 ( .A(n4846), .B(n4434), .Z(out[797]) );
  XOR U6341 ( .A(in[709]), .B(n4435), .Z(n4646) );
  IV U6342 ( .A(n4646), .Z(n4850) );
  NANDN U6343 ( .A(n4645), .B(n4436), .Z(n4437) );
  XOR U6344 ( .A(n4850), .B(n4437), .Z(out[798]) );
  XOR U6345 ( .A(in[710]), .B(n4438), .Z(n4854) );
  NANDN U6346 ( .A(n4648), .B(n4439), .Z(n4440) );
  XOR U6347 ( .A(n4854), .B(n4440), .Z(out[799]) );
  ANDN U6348 ( .B(n4442), .A(n4441), .Z(n4443) );
  XOR U6349 ( .A(n4444), .B(n4443), .Z(out[79]) );
  OR U6350 ( .A(n4446), .B(n4445), .Z(n4447) );
  XNOR U6351 ( .A(n4448), .B(n4447), .Z(out[7]) );
  XOR U6352 ( .A(in[711]), .B(n4449), .Z(n4650) );
  IV U6353 ( .A(n4650), .Z(n4858) );
  NANDN U6354 ( .A(n4649), .B(n4450), .Z(n4451) );
  XOR U6355 ( .A(n4858), .B(n4451), .Z(out[800]) );
  XOR U6356 ( .A(in[712]), .B(n4452), .Z(n4653) );
  IV U6357 ( .A(n4653), .Z(n4862) );
  NANDN U6358 ( .A(n4652), .B(n4453), .Z(n4454) );
  XOR U6359 ( .A(n4862), .B(n4454), .Z(out[801]) );
  XOR U6360 ( .A(in[713]), .B(n4455), .Z(n4656) );
  IV U6361 ( .A(n4656), .Z(n4870) );
  NANDN U6362 ( .A(n4655), .B(n4456), .Z(n4457) );
  XOR U6363 ( .A(n4870), .B(n4457), .Z(out[802]) );
  XOR U6364 ( .A(in[714]), .B(n4458), .Z(n4659) );
  IV U6365 ( .A(n4659), .Z(n4874) );
  NANDN U6366 ( .A(n4658), .B(n4459), .Z(n4460) );
  XOR U6367 ( .A(n4874), .B(n4460), .Z(out[803]) );
  XOR U6368 ( .A(in[715]), .B(n4461), .Z(n4662) );
  IV U6369 ( .A(n4662), .Z(n4878) );
  NANDN U6370 ( .A(n4661), .B(n4462), .Z(n4463) );
  XOR U6371 ( .A(n4878), .B(n4463), .Z(out[804]) );
  XNOR U6372 ( .A(n4464), .B(in[716]), .Z(n4882) );
  NANDN U6373 ( .A(n4664), .B(n4465), .Z(n4466) );
  XNOR U6374 ( .A(n4882), .B(n4466), .Z(out[805]) );
  XNOR U6375 ( .A(n4467), .B(in[717]), .Z(n4886) );
  NANDN U6376 ( .A(n4669), .B(n4468), .Z(n4469) );
  XNOR U6377 ( .A(n4886), .B(n4469), .Z(out[806]) );
  XNOR U6378 ( .A(n4470), .B(in[718]), .Z(n4890) );
  NANDN U6379 ( .A(n4670), .B(n4471), .Z(n4472) );
  XNOR U6380 ( .A(n4890), .B(n4472), .Z(out[807]) );
  XNOR U6381 ( .A(n4473), .B(in[719]), .Z(n4894) );
  NANDN U6382 ( .A(n4671), .B(n4474), .Z(n4475) );
  XNOR U6383 ( .A(n4894), .B(n4475), .Z(out[808]) );
  XNOR U6384 ( .A(n4476), .B(in[720]), .Z(n4898) );
  NANDN U6385 ( .A(n4672), .B(n4477), .Z(n4478) );
  XNOR U6386 ( .A(n4898), .B(n4478), .Z(out[809]) );
  ANDN U6387 ( .B(n4480), .A(n4479), .Z(n4481) );
  XOR U6388 ( .A(n4482), .B(n4481), .Z(out[80]) );
  XNOR U6389 ( .A(n4483), .B(in[721]), .Z(n4902) );
  NANDN U6390 ( .A(n4673), .B(n4484), .Z(n4485) );
  XNOR U6391 ( .A(n4902), .B(n4485), .Z(out[810]) );
  XNOR U6392 ( .A(n4486), .B(in[722]), .Z(n4906) );
  NAND U6393 ( .A(n4487), .B(n4674), .Z(n4488) );
  XNOR U6394 ( .A(n4906), .B(n4488), .Z(out[811]) );
  XNOR U6395 ( .A(n4489), .B(in[723]), .Z(n4913) );
  NANDN U6396 ( .A(n4676), .B(n4490), .Z(n4491) );
  XNOR U6397 ( .A(n4913), .B(n4491), .Z(out[812]) );
  XNOR U6398 ( .A(in[724]), .B(n4492), .Z(n4917) );
  NANDN U6399 ( .A(n4677), .B(n4493), .Z(n4494) );
  XNOR U6400 ( .A(n4917), .B(n4494), .Z(out[813]) );
  XNOR U6401 ( .A(in[725]), .B(n4495), .Z(n4921) );
  NANDN U6402 ( .A(n4678), .B(n4496), .Z(n4497) );
  XNOR U6403 ( .A(n4921), .B(n4497), .Z(out[814]) );
  XNOR U6404 ( .A(in[726]), .B(n4498), .Z(n4925) );
  NANDN U6405 ( .A(n4679), .B(n4499), .Z(n4500) );
  XNOR U6406 ( .A(n4925), .B(n4500), .Z(out[815]) );
  XNOR U6407 ( .A(in[727]), .B(n4501), .Z(n4929) );
  NANDN U6408 ( .A(n4684), .B(n4502), .Z(n4503) );
  XNOR U6409 ( .A(n4929), .B(n4503), .Z(out[816]) );
  XNOR U6410 ( .A(in[728]), .B(n4504), .Z(n4933) );
  NANDN U6411 ( .A(n4685), .B(n4505), .Z(n4506) );
  XNOR U6412 ( .A(n4933), .B(n4506), .Z(out[817]) );
  XNOR U6413 ( .A(in[729]), .B(n4507), .Z(n4937) );
  NANDN U6414 ( .A(n4686), .B(n4508), .Z(n4509) );
  XNOR U6415 ( .A(n4937), .B(n4509), .Z(out[818]) );
  XNOR U6416 ( .A(in[730]), .B(n4510), .Z(n4941) );
  NANDN U6417 ( .A(n4687), .B(n4511), .Z(n4512) );
  XNOR U6418 ( .A(n4941), .B(n4512), .Z(out[819]) );
  ANDN U6419 ( .B(n4514), .A(n4513), .Z(n4515) );
  XOR U6420 ( .A(n4516), .B(n4515), .Z(out[81]) );
  XOR U6421 ( .A(in[731]), .B(n4517), .Z(n4945) );
  NANDN U6422 ( .A(n4688), .B(n4518), .Z(n4519) );
  XNOR U6423 ( .A(n4945), .B(n4519), .Z(out[820]) );
  XOR U6424 ( .A(in[732]), .B(n4520), .Z(n4949) );
  NANDN U6425 ( .A(n4689), .B(n4521), .Z(n4522) );
  XNOR U6426 ( .A(n4949), .B(n4522), .Z(out[821]) );
  XOR U6427 ( .A(in[733]), .B(n4523), .Z(n4957) );
  NANDN U6428 ( .A(n4690), .B(n4524), .Z(n4525) );
  XNOR U6429 ( .A(n4957), .B(n4525), .Z(out[822]) );
  XNOR U6430 ( .A(in[734]), .B(n4526), .Z(n4961) );
  IV U6431 ( .A(n4527), .Z(n4691) );
  NANDN U6432 ( .A(n4528), .B(n4691), .Z(n4529) );
  XNOR U6433 ( .A(n4961), .B(n4529), .Z(out[823]) );
  XNOR U6434 ( .A(in[735]), .B(n4530), .Z(n4965) );
  IV U6435 ( .A(n4531), .Z(n4693) );
  NANDN U6436 ( .A(n4532), .B(n4693), .Z(n4533) );
  XNOR U6437 ( .A(n4965), .B(n4533), .Z(out[824]) );
  XNOR U6438 ( .A(in[736]), .B(n4534), .Z(n4969) );
  IV U6439 ( .A(n4535), .Z(n4695) );
  NANDN U6440 ( .A(n4536), .B(n4695), .Z(n4537) );
  XNOR U6441 ( .A(n4969), .B(n4537), .Z(out[825]) );
  XNOR U6442 ( .A(in[737]), .B(n4538), .Z(n4973) );
  IV U6443 ( .A(n4539), .Z(n4700) );
  NANDN U6444 ( .A(n4540), .B(n4700), .Z(n4541) );
  XNOR U6445 ( .A(n4973), .B(n4541), .Z(out[826]) );
  XNOR U6446 ( .A(in[738]), .B(n4542), .Z(n4977) );
  IV U6447 ( .A(n4543), .Z(n4702) );
  NANDN U6448 ( .A(n4544), .B(n4702), .Z(n4545) );
  XNOR U6449 ( .A(n4977), .B(n4545), .Z(out[827]) );
  XNOR U6450 ( .A(in[739]), .B(n4546), .Z(n4981) );
  IV U6451 ( .A(n4547), .Z(n4704) );
  NANDN U6452 ( .A(n4548), .B(n4704), .Z(n4549) );
  XNOR U6453 ( .A(n4981), .B(n4549), .Z(out[828]) );
  XOR U6454 ( .A(in[740]), .B(n4550), .Z(n4707) );
  IV U6455 ( .A(n4707), .Z(n4985) );
  ANDN U6456 ( .B(n4553), .A(n4552), .Z(n4554) );
  XOR U6457 ( .A(n4555), .B(n4554), .Z(out[82]) );
  XOR U6458 ( .A(in[741]), .B(n4556), .Z(n4710) );
  IV U6459 ( .A(n4710), .Z(n4989) );
  XOR U6460 ( .A(in[742]), .B(n4558), .Z(n4713) );
  IV U6461 ( .A(n4713), .Z(n4993) );
  NANDN U6462 ( .A(n4561), .B(n4560), .Z(n4562) );
  XOR U6463 ( .A(n4716), .B(n4562), .Z(out[832]) );
  NANDN U6464 ( .A(n4564), .B(n4563), .Z(n4565) );
  XOR U6465 ( .A(n4720), .B(n4565), .Z(out[833]) );
  NANDN U6466 ( .A(n4567), .B(n4566), .Z(n4568) );
  XOR U6467 ( .A(n4724), .B(n4568), .Z(out[834]) );
  NANDN U6468 ( .A(n4570), .B(n4569), .Z(n4571) );
  XOR U6469 ( .A(n4728), .B(n4571), .Z(out[835]) );
  NANDN U6470 ( .A(n4572), .B(n4739), .Z(n4573) );
  XOR U6471 ( .A(n4740), .B(n4573), .Z(out[836]) );
  NANDN U6472 ( .A(n4574), .B(n4743), .Z(n4575) );
  XOR U6473 ( .A(n4744), .B(n4575), .Z(out[837]) );
  NANDN U6474 ( .A(n4576), .B(n4747), .Z(n4577) );
  XOR U6475 ( .A(n4748), .B(n4577), .Z(out[838]) );
  NANDN U6476 ( .A(n4579), .B(n4578), .Z(n4580) );
  XOR U6477 ( .A(n4752), .B(n4580), .Z(out[839]) );
  ANDN U6478 ( .B(n4582), .A(n4581), .Z(n4583) );
  XOR U6479 ( .A(n4584), .B(n4583), .Z(out[83]) );
  NANDN U6480 ( .A(n4585), .B(n4756), .Z(n4586) );
  XNOR U6481 ( .A(n4755), .B(n4586), .Z(out[840]) );
  NANDN U6482 ( .A(n4587), .B(n4760), .Z(n4588) );
  XNOR U6483 ( .A(n4759), .B(n4588), .Z(out[841]) );
  NANDN U6484 ( .A(n4589), .B(n4764), .Z(n4590) );
  XNOR U6485 ( .A(n4763), .B(n4590), .Z(out[842]) );
  NANDN U6486 ( .A(n4591), .B(n4768), .Z(n4592) );
  XNOR U6487 ( .A(n4767), .B(n4592), .Z(out[843]) );
  NANDN U6488 ( .A(n4593), .B(n4772), .Z(n4594) );
  XNOR U6489 ( .A(n4771), .B(n4594), .Z(out[844]) );
  NANDN U6490 ( .A(n4595), .B(n4776), .Z(n4596) );
  XNOR U6491 ( .A(n4775), .B(n4596), .Z(out[845]) );
  NANDN U6492 ( .A(n4597), .B(n4783), .Z(n4598) );
  XNOR U6493 ( .A(n4782), .B(n4598), .Z(out[846]) );
  NANDN U6494 ( .A(n4599), .B(n4787), .Z(n4600) );
  XNOR U6495 ( .A(n4786), .B(n4600), .Z(out[847]) );
  NANDN U6496 ( .A(n4602), .B(n4601), .Z(n4603) );
  XNOR U6497 ( .A(n4790), .B(n4603), .Z(out[848]) );
  NANDN U6498 ( .A(n4604), .B(n4795), .Z(n4605) );
  XNOR U6499 ( .A(n4794), .B(n4605), .Z(out[849]) );
  ANDN U6500 ( .B(n4607), .A(n4606), .Z(n4608) );
  XOR U6501 ( .A(n4609), .B(n4608), .Z(out[84]) );
  NANDN U6502 ( .A(n4610), .B(n4799), .Z(n4611) );
  XNOR U6503 ( .A(n4798), .B(n4611), .Z(out[850]) );
  NANDN U6504 ( .A(n4612), .B(n4803), .Z(n4613) );
  XNOR U6505 ( .A(n4802), .B(n4613), .Z(out[851]) );
  NANDN U6506 ( .A(n4614), .B(n4807), .Z(n4615) );
  XNOR U6507 ( .A(n4806), .B(n4615), .Z(out[852]) );
  NANDN U6508 ( .A(n4616), .B(n4811), .Z(n4617) );
  XNOR U6509 ( .A(n4810), .B(n4617), .Z(out[853]) );
  NANDN U6510 ( .A(n4618), .B(n4815), .Z(n4619) );
  XNOR U6511 ( .A(n4814), .B(n4619), .Z(out[854]) );
  NANDN U6512 ( .A(n4621), .B(n4620), .Z(n4622) );
  XNOR U6513 ( .A(n4818), .B(n4622), .Z(out[855]) );
  NANDN U6514 ( .A(n4624), .B(n4623), .Z(n4625) );
  XNOR U6515 ( .A(n4825), .B(n4625), .Z(out[856]) );
  NANDN U6516 ( .A(n4627), .B(n4626), .Z(n4628) );
  XNOR U6517 ( .A(n4829), .B(n4628), .Z(out[857]) );
  NANDN U6518 ( .A(n4630), .B(n4629), .Z(n4631) );
  XNOR U6519 ( .A(n4833), .B(n4631), .Z(out[858]) );
  NANDN U6520 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U6521 ( .A(n4837), .B(n4634), .Z(out[859]) );
  ANDN U6522 ( .B(n4636), .A(n4635), .Z(n4637) );
  XOR U6523 ( .A(n4638), .B(n4637), .Z(out[85]) );
  NANDN U6524 ( .A(n4640), .B(n4639), .Z(n4641) );
  XNOR U6525 ( .A(n4841), .B(n4641), .Z(out[860]) );
  NANDN U6526 ( .A(n4643), .B(n4642), .Z(n4644) );
  XNOR U6527 ( .A(n4845), .B(n4644), .Z(out[861]) );
  NANDN U6528 ( .A(n4646), .B(n4645), .Z(n4647) );
  XNOR U6529 ( .A(n4849), .B(n4647), .Z(out[862]) );
  NANDN U6530 ( .A(n4650), .B(n4649), .Z(n4651) );
  XNOR U6531 ( .A(n4857), .B(n4651), .Z(out[864]) );
  NANDN U6532 ( .A(n4653), .B(n4652), .Z(n4654) );
  XNOR U6533 ( .A(n4861), .B(n4654), .Z(out[865]) );
  NANDN U6534 ( .A(n4656), .B(n4655), .Z(n4657) );
  XNOR U6535 ( .A(n4869), .B(n4657), .Z(out[866]) );
  NANDN U6536 ( .A(n4659), .B(n4658), .Z(n4660) );
  XNOR U6537 ( .A(n4873), .B(n4660), .Z(out[867]) );
  NANDN U6538 ( .A(n4662), .B(n4661), .Z(n4663) );
  XNOR U6539 ( .A(n4877), .B(n4663), .Z(out[868]) );
  ANDN U6540 ( .B(n4666), .A(n4665), .Z(n4667) );
  XOR U6541 ( .A(n4668), .B(n4667), .Z(out[86]) );
  OR U6542 ( .A(n4906), .B(n4674), .Z(n4675) );
  XNOR U6543 ( .A(n4905), .B(n4675), .Z(out[875]) );
  ANDN U6544 ( .B(n4681), .A(n4680), .Z(n4682) );
  XOR U6545 ( .A(n4683), .B(n4682), .Z(out[87]) );
  OR U6546 ( .A(n4961), .B(n4691), .Z(n4692) );
  XOR U6547 ( .A(n4962), .B(n4692), .Z(out[887]) );
  OR U6548 ( .A(n4965), .B(n4693), .Z(n4694) );
  XOR U6549 ( .A(n4966), .B(n4694), .Z(out[888]) );
  OR U6550 ( .A(n4969), .B(n4695), .Z(n4696) );
  XOR U6551 ( .A(n4970), .B(n4696), .Z(out[889]) );
  OR U6552 ( .A(n4973), .B(n4700), .Z(n4701) );
  XOR U6553 ( .A(n4974), .B(n4701), .Z(out[890]) );
  OR U6554 ( .A(n4977), .B(n4702), .Z(n4703) );
  XOR U6555 ( .A(n4978), .B(n4703), .Z(out[891]) );
  OR U6556 ( .A(n4981), .B(n4704), .Z(n4705) );
  XOR U6557 ( .A(n4982), .B(n4705), .Z(out[892]) );
  NANDN U6558 ( .A(n4707), .B(n4706), .Z(n4708) );
  XOR U6559 ( .A(n4986), .B(n4708), .Z(out[893]) );
  NANDN U6560 ( .A(n4710), .B(n4709), .Z(n4711) );
  XOR U6561 ( .A(n4990), .B(n4711), .Z(out[894]) );
  NANDN U6562 ( .A(n4713), .B(n4712), .Z(n4714) );
  XOR U6563 ( .A(n4994), .B(n4714), .Z(out[895]) );
  ANDN U6564 ( .B(n4716), .A(n4715), .Z(n4717) );
  XOR U6565 ( .A(n4718), .B(n4717), .Z(out[896]) );
  ANDN U6566 ( .B(n4720), .A(n4719), .Z(n4721) );
  XOR U6567 ( .A(n4722), .B(n4721), .Z(out[897]) );
  ANDN U6568 ( .B(n4724), .A(n4723), .Z(n4725) );
  XOR U6569 ( .A(n4726), .B(n4725), .Z(out[898]) );
  ANDN U6570 ( .B(n4728), .A(n4727), .Z(n4729) );
  XOR U6571 ( .A(n4730), .B(n4729), .Z(out[899]) );
  ANDN U6572 ( .B(n4732), .A(n4731), .Z(n4733) );
  XOR U6573 ( .A(n4734), .B(n4733), .Z(out[89]) );
  OR U6574 ( .A(n4736), .B(n4735), .Z(n4737) );
  XNOR U6575 ( .A(n4738), .B(n4737), .Z(out[8]) );
  ANDN U6576 ( .B(n4740), .A(n4739), .Z(n4741) );
  XOR U6577 ( .A(n4742), .B(n4741), .Z(out[900]) );
  ANDN U6578 ( .B(n4744), .A(n4743), .Z(n4745) );
  XOR U6579 ( .A(n4746), .B(n4745), .Z(out[901]) );
  ANDN U6580 ( .B(n4748), .A(n4747), .Z(n4749) );
  XOR U6581 ( .A(n4750), .B(n4749), .Z(out[902]) );
  ANDN U6582 ( .B(n4752), .A(n4751), .Z(n4753) );
  XOR U6583 ( .A(n4754), .B(n4753), .Z(out[903]) );
  NOR U6584 ( .A(n4756), .B(n4755), .Z(n4757) );
  XOR U6585 ( .A(n4758), .B(n4757), .Z(out[904]) );
  NOR U6586 ( .A(n4760), .B(n4759), .Z(n4761) );
  XOR U6587 ( .A(n4762), .B(n4761), .Z(out[905]) );
  NOR U6588 ( .A(n4764), .B(n4763), .Z(n4765) );
  XOR U6589 ( .A(n4766), .B(n4765), .Z(out[906]) );
  NOR U6590 ( .A(n4768), .B(n4767), .Z(n4769) );
  XOR U6591 ( .A(n4770), .B(n4769), .Z(out[907]) );
  NOR U6592 ( .A(n4772), .B(n4771), .Z(n4773) );
  XOR U6593 ( .A(n4774), .B(n4773), .Z(out[908]) );
  NOR U6594 ( .A(n4776), .B(n4775), .Z(n4777) );
  XOR U6595 ( .A(n4778), .B(n4777), .Z(out[909]) );
  NOR U6596 ( .A(n4783), .B(n4782), .Z(n4784) );
  XOR U6597 ( .A(n4785), .B(n4784), .Z(out[910]) );
  NOR U6598 ( .A(n4787), .B(n4786), .Z(n4788) );
  XOR U6599 ( .A(n4789), .B(n4788), .Z(out[911]) );
  NOR U6600 ( .A(n4791), .B(n4790), .Z(n4792) );
  XOR U6601 ( .A(n4793), .B(n4792), .Z(out[912]) );
  NOR U6602 ( .A(n4795), .B(n4794), .Z(n4796) );
  XOR U6603 ( .A(n4797), .B(n4796), .Z(out[913]) );
  NOR U6604 ( .A(n4799), .B(n4798), .Z(n4800) );
  XOR U6605 ( .A(n4801), .B(n4800), .Z(out[914]) );
  NOR U6606 ( .A(n4803), .B(n4802), .Z(n4804) );
  XOR U6607 ( .A(n4805), .B(n4804), .Z(out[915]) );
  NOR U6608 ( .A(n4807), .B(n4806), .Z(n4808) );
  XOR U6609 ( .A(n4809), .B(n4808), .Z(out[916]) );
  NOR U6610 ( .A(n4811), .B(n4810), .Z(n4812) );
  XOR U6611 ( .A(n4813), .B(n4812), .Z(out[917]) );
  NOR U6612 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U6613 ( .A(n4817), .B(n4816), .Z(out[918]) );
  NOR U6614 ( .A(n4819), .B(n4818), .Z(n4820) );
  XOR U6615 ( .A(n4821), .B(n4820), .Z(out[919]) );
  NOR U6616 ( .A(n4826), .B(n4825), .Z(n4827) );
  XOR U6617 ( .A(n4828), .B(n4827), .Z(out[920]) );
  NOR U6618 ( .A(n4830), .B(n4829), .Z(n4831) );
  XOR U6619 ( .A(n4832), .B(n4831), .Z(out[921]) );
  NOR U6620 ( .A(n4834), .B(n4833), .Z(n4835) );
  XOR U6621 ( .A(n4836), .B(n4835), .Z(out[922]) );
  NOR U6622 ( .A(n4838), .B(n4837), .Z(n4839) );
  XOR U6623 ( .A(n4840), .B(n4839), .Z(out[923]) );
  NOR U6624 ( .A(n4842), .B(n4841), .Z(n4843) );
  XOR U6625 ( .A(n4844), .B(n4843), .Z(out[924]) );
  NOR U6626 ( .A(n4846), .B(n4845), .Z(n4847) );
  XOR U6627 ( .A(n4848), .B(n4847), .Z(out[925]) );
  NOR U6628 ( .A(n4850), .B(n4849), .Z(n4851) );
  XOR U6629 ( .A(n4852), .B(n4851), .Z(out[926]) );
  NOR U6630 ( .A(n4854), .B(n4853), .Z(n4855) );
  XOR U6631 ( .A(n4856), .B(n4855), .Z(out[927]) );
  NOR U6632 ( .A(n4858), .B(n4857), .Z(n4859) );
  XOR U6633 ( .A(n4860), .B(n4859), .Z(out[928]) );
  NOR U6634 ( .A(n4862), .B(n4861), .Z(n4863) );
  XOR U6635 ( .A(n4864), .B(n4863), .Z(out[929]) );
  AND U6636 ( .A(n4866), .B(n4865), .Z(n4867) );
  XNOR U6637 ( .A(n4868), .B(n4867), .Z(out[92]) );
  NOR U6638 ( .A(n4870), .B(n4869), .Z(n4871) );
  XOR U6639 ( .A(n4872), .B(n4871), .Z(out[930]) );
  NOR U6640 ( .A(n4874), .B(n4873), .Z(n4875) );
  XOR U6641 ( .A(n4876), .B(n4875), .Z(out[931]) );
  NOR U6642 ( .A(n4878), .B(n4877), .Z(n4879) );
  XOR U6643 ( .A(n4880), .B(n4879), .Z(out[932]) );
  ANDN U6644 ( .B(n4882), .A(n4881), .Z(n4883) );
  XOR U6645 ( .A(n4884), .B(n4883), .Z(out[933]) );
  ANDN U6646 ( .B(n4886), .A(n4885), .Z(n4887) );
  XOR U6647 ( .A(n4888), .B(n4887), .Z(out[934]) );
  ANDN U6648 ( .B(n4890), .A(n4889), .Z(n4891) );
  XOR U6649 ( .A(n4892), .B(n4891), .Z(out[935]) );
  ANDN U6650 ( .B(n4894), .A(n4893), .Z(n4895) );
  XOR U6651 ( .A(n4896), .B(n4895), .Z(out[936]) );
  ANDN U6652 ( .B(n4898), .A(n4897), .Z(n4899) );
  XOR U6653 ( .A(n4900), .B(n4899), .Z(out[937]) );
  ANDN U6654 ( .B(n4902), .A(n4901), .Z(n4903) );
  XOR U6655 ( .A(n4904), .B(n4903), .Z(out[938]) );
  ANDN U6656 ( .B(n4906), .A(n4905), .Z(n4907) );
  XOR U6657 ( .A(n4908), .B(n4907), .Z(out[939]) );
  AND U6658 ( .A(n4910), .B(n4909), .Z(n4911) );
  XNOR U6659 ( .A(n4912), .B(n4911), .Z(out[93]) );
  AND U6660 ( .A(n4914), .B(n4913), .Z(n4915) );
  XNOR U6661 ( .A(n4916), .B(n4915), .Z(out[940]) );
  AND U6662 ( .A(n4918), .B(n4917), .Z(n4919) );
  XNOR U6663 ( .A(n4920), .B(n4919), .Z(out[941]) );
  AND U6664 ( .A(n4922), .B(n4921), .Z(n4923) );
  XNOR U6665 ( .A(n4924), .B(n4923), .Z(out[942]) );
  AND U6666 ( .A(n4926), .B(n4925), .Z(n4927) );
  XNOR U6667 ( .A(n4928), .B(n4927), .Z(out[943]) );
  AND U6668 ( .A(n4930), .B(n4929), .Z(n4931) );
  XNOR U6669 ( .A(n4932), .B(n4931), .Z(out[944]) );
  AND U6670 ( .A(n4934), .B(n4933), .Z(n4935) );
  XNOR U6671 ( .A(n4936), .B(n4935), .Z(out[945]) );
  AND U6672 ( .A(n4938), .B(n4937), .Z(n4939) );
  XNOR U6673 ( .A(n4940), .B(n4939), .Z(out[946]) );
  AND U6674 ( .A(n4942), .B(n4941), .Z(n4943) );
  XNOR U6675 ( .A(n4944), .B(n4943), .Z(out[947]) );
  AND U6676 ( .A(n4946), .B(n4945), .Z(n4947) );
  XNOR U6677 ( .A(n4948), .B(n4947), .Z(out[948]) );
  AND U6678 ( .A(n4950), .B(n4949), .Z(n4951) );
  XNOR U6679 ( .A(n4952), .B(n4951), .Z(out[949]) );
  AND U6680 ( .A(n4954), .B(n4953), .Z(n4955) );
  XNOR U6681 ( .A(n4956), .B(n4955), .Z(out[94]) );
  AND U6682 ( .A(n4958), .B(n4957), .Z(n4959) );
  XNOR U6683 ( .A(n4960), .B(n4959), .Z(out[950]) );
  AND U6684 ( .A(n4962), .B(n4961), .Z(n4963) );
  XNOR U6685 ( .A(n4964), .B(n4963), .Z(out[951]) );
  AND U6686 ( .A(n4966), .B(n4965), .Z(n4967) );
  XNOR U6687 ( .A(n4968), .B(n4967), .Z(out[952]) );
  AND U6688 ( .A(n4970), .B(n4969), .Z(n4971) );
  XNOR U6689 ( .A(n4972), .B(n4971), .Z(out[953]) );
  AND U6690 ( .A(n4974), .B(n4973), .Z(n4975) );
  XNOR U6691 ( .A(n4976), .B(n4975), .Z(out[954]) );
  AND U6692 ( .A(n4978), .B(n4977), .Z(n4979) );
  XNOR U6693 ( .A(n4980), .B(n4979), .Z(out[955]) );
  AND U6694 ( .A(n4982), .B(n4981), .Z(n4983) );
  XOR U6695 ( .A(n4984), .B(n4983), .Z(out[956]) );
  ANDN U6696 ( .B(n4986), .A(n4985), .Z(n4987) );
  XOR U6697 ( .A(n4988), .B(n4987), .Z(out[957]) );
  ANDN U6698 ( .B(n4990), .A(n4989), .Z(n4991) );
  XOR U6699 ( .A(n4992), .B(n4991), .Z(out[958]) );
  ANDN U6700 ( .B(n4994), .A(n4993), .Z(n4995) );
  XNOR U6701 ( .A(n4996), .B(n4995), .Z(out[959]) );
  AND U6702 ( .A(n4998), .B(n4997), .Z(n4999) );
  XNOR U6703 ( .A(n5000), .B(n4999), .Z(out[95]) );
  ANDN U6704 ( .B(n5002), .A(n5001), .Z(n5003) );
  XOR U6705 ( .A(n5004), .B(n5003), .Z(out[960]) );
  ANDN U6706 ( .B(n5006), .A(n5005), .Z(n5007) );
  XOR U6707 ( .A(n5008), .B(n5007), .Z(out[961]) );
  ANDN U6708 ( .B(n5010), .A(n5009), .Z(n5011) );
  XOR U6709 ( .A(n5012), .B(n5011), .Z(out[962]) );
  ANDN U6710 ( .B(n5014), .A(n5013), .Z(n5015) );
  XOR U6711 ( .A(n5016), .B(n5015), .Z(out[963]) );
  ANDN U6712 ( .B(n5018), .A(n5017), .Z(n5019) );
  XOR U6713 ( .A(n5020), .B(n5019), .Z(out[964]) );
  ANDN U6714 ( .B(n5022), .A(n5021), .Z(n5023) );
  XOR U6715 ( .A(n5024), .B(n5023), .Z(out[965]) );
  ANDN U6716 ( .B(n5026), .A(n5025), .Z(n5027) );
  XOR U6717 ( .A(n5028), .B(n5027), .Z(out[966]) );
  ANDN U6718 ( .B(n5030), .A(n5029), .Z(n5031) );
  XOR U6719 ( .A(n5032), .B(n5031), .Z(out[967]) );
  ANDN U6720 ( .B(n5034), .A(n5033), .Z(n5035) );
  XOR U6721 ( .A(n5036), .B(n5035), .Z(out[968]) );
  ANDN U6722 ( .B(n5038), .A(n5037), .Z(n5039) );
  XOR U6723 ( .A(n5040), .B(n5039), .Z(out[969]) );
  AND U6724 ( .A(n5042), .B(n5041), .Z(n5043) );
  XNOR U6725 ( .A(n5044), .B(n5043), .Z(out[96]) );
  ANDN U6726 ( .B(n5046), .A(n5045), .Z(n5047) );
  XOR U6727 ( .A(n5048), .B(n5047), .Z(out[970]) );
  ANDN U6728 ( .B(n5050), .A(n5049), .Z(n5051) );
  XOR U6729 ( .A(n5052), .B(n5051), .Z(out[971]) );
  ANDN U6730 ( .B(n5054), .A(n5053), .Z(n5055) );
  XOR U6731 ( .A(n5056), .B(n5055), .Z(out[972]) );
  ANDN U6732 ( .B(n5058), .A(n5057), .Z(n5059) );
  XOR U6733 ( .A(n5060), .B(n5059), .Z(out[973]) );
  ANDN U6734 ( .B(n5062), .A(n5061), .Z(n5063) );
  XOR U6735 ( .A(n5064), .B(n5063), .Z(out[974]) );
  ANDN U6736 ( .B(n5066), .A(n5065), .Z(n5067) );
  XOR U6737 ( .A(n5068), .B(n5067), .Z(out[975]) );
  ANDN U6738 ( .B(n5079), .A(n5078), .Z(n5080) );
  XOR U6739 ( .A(n5081), .B(n5080), .Z(out[979]) );
  AND U6740 ( .A(n5083), .B(n5082), .Z(n5084) );
  XNOR U6741 ( .A(n5085), .B(n5084), .Z(out[97]) );
  ANDN U6742 ( .B(n5111), .A(n5110), .Z(n5112) );
  XOR U6743 ( .A(n5113), .B(n5112), .Z(out[988]) );
  ANDN U6744 ( .B(n5118), .A(n5117), .Z(n5119) );
  XNOR U6745 ( .A(n5120), .B(n5119), .Z(out[98]) );
  ANDN U6746 ( .B(n5125), .A(n5124), .Z(n5126) );
  XOR U6747 ( .A(n5127), .B(n5126), .Z(out[991]) );
  ANDN U6748 ( .B(n5129), .A(n5128), .Z(n5130) );
  XOR U6749 ( .A(n5131), .B(n5130), .Z(out[992]) );
  ANDN U6750 ( .B(n5133), .A(n5132), .Z(n5134) );
  XOR U6751 ( .A(n5135), .B(n5134), .Z(out[993]) );
  ANDN U6752 ( .B(n5137), .A(n5136), .Z(n5138) );
  XOR U6753 ( .A(n5139), .B(n5138), .Z(out[994]) );
  ANDN U6754 ( .B(n5141), .A(n5140), .Z(n5142) );
  XNOR U6755 ( .A(n5143), .B(n5142), .Z(out[995]) );
  ANDN U6756 ( .B(n5145), .A(n5144), .Z(n5146) );
  XNOR U6757 ( .A(n5147), .B(n5146), .Z(out[996]) );
  ANDN U6758 ( .B(n5149), .A(n5148), .Z(n5150) );
  XNOR U6759 ( .A(n5151), .B(n5150), .Z(out[997]) );
  AND U6760 ( .A(n5153), .B(n5152), .Z(n5154) );
  XNOR U6761 ( .A(n5155), .B(n5154), .Z(out[998]) );
  ANDN U6762 ( .B(n5157), .A(n5156), .Z(n5158) );
  XNOR U6763 ( .A(n5159), .B(n5158), .Z(out[999]) );
  ANDN U6764 ( .B(n5161), .A(n5160), .Z(n5162) );
  XNOR U6765 ( .A(n5163), .B(n5162), .Z(out[99]) );
  OR U6766 ( .A(n5165), .B(n5164), .Z(n5166) );
  XNOR U6767 ( .A(n5167), .B(n5166), .Z(out[9]) );
endmodule


module round_4 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_31, round_const_15, round_const_7, round_const_3, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156;
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XNOR U1 ( .A(n1716), .B(n1717), .Z(n3088) );
  XOR U2 ( .A(n1432), .B(n1390), .Z(n4458) );
  XOR U3 ( .A(n1394), .B(n1434), .Z(n4461) );
  XOR U4 ( .A(n1435), .B(n1398), .Z(n4464) );
  XOR U5 ( .A(n1438), .B(n1406), .Z(n4470) );
  NAND U6 ( .A(n2901), .B(n4476), .Z(n1) );
  XNOR U7 ( .A(n2900), .B(n1), .Z(out[208]) );
  AND U8 ( .A(n4671), .B(n4670), .Z(n2) );
  XNOR U9 ( .A(n4672), .B(n2), .Z(out[87]) );
  AND U10 ( .A(n4813), .B(n4812), .Z(n3) );
  XNOR U11 ( .A(n4814), .B(n3), .Z(out[91]) );
  NAND U12 ( .A(n4638), .B(n4844), .Z(n4) );
  XNOR U13 ( .A(n4843), .B(n4), .Z(out[863]) );
  AND U14 ( .A(n4740), .B(n4352), .Z(n5) );
  XNOR U15 ( .A(n4570), .B(n5), .Z(out[710]) );
  XNOR U16 ( .A(n1452), .B(n1014), .Z(n2759) );
  XNOR U17 ( .A(n1456), .B(n1040), .Z(n2783) );
  XNOR U18 ( .A(n1460), .B(n1053), .Z(n2797) );
  XNOR U19 ( .A(n1462), .B(n1066), .Z(n2820) );
  XNOR U20 ( .A(n1474), .B(n1107), .Z(n2891) );
  XNOR U21 ( .A(n1450), .B(n1758), .Z(n3216) );
  XOR U22 ( .A(n1447), .B(n755), .Z(n4486) );
  XOR U23 ( .A(n1453), .B(n800), .Z(n4495) );
  XNOR U24 ( .A(n3974), .B(in[1489]), .Z(n4791) );
  NANDN U25 ( .A(n2919), .B(n4658), .Z(n6) );
  XNOR U26 ( .A(n2918), .B(n6), .Z(out[214]) );
  ANDN U27 ( .B(n1908), .A(n1501), .Z(n7) );
  XNOR U28 ( .A(n1761), .B(n7), .Z(out[1064]) );
  ANDN U29 ( .B(n1912), .A(n1505), .Z(n8) );
  XNOR U30 ( .A(n1763), .B(n8), .Z(out[1065]) );
  NANDN U31 ( .A(n1515), .B(n1920), .Z(n9) );
  XNOR U32 ( .A(n1767), .B(n9), .Z(out[1067]) );
  ANDN U33 ( .B(n1950), .A(n1543), .Z(n10) );
  XNOR U34 ( .A(n1782), .B(n10), .Z(out[1074]) );
  ANDN U35 ( .B(n1958), .A(n1553), .Z(n11) );
  XNOR U36 ( .A(n1786), .B(n11), .Z(out[1076]) );
  ANDN U37 ( .B(n1962), .A(n1557), .Z(n12) );
  XNOR U38 ( .A(n1788), .B(n12), .Z(out[1077]) );
  ANDN U39 ( .B(n1968), .A(n1561), .Z(n13) );
  XNOR U40 ( .A(n1790), .B(n13), .Z(out[1078]) );
  NANDN U41 ( .A(n3982), .B(n3981), .Z(n14) );
  XNOR U42 ( .A(n3983), .B(n14), .Z(out[65]) );
  NANDN U43 ( .A(n4880), .B(n4660), .Z(n15) );
  XNOR U44 ( .A(n4879), .B(n15), .Z(out[871]) );
  NAND U45 ( .A(n2859), .B(n2858), .Z(n16) );
  XNOR U46 ( .A(n3939), .B(n16), .Z(out[256]) );
  NANDN U47 ( .A(n2888), .B(n2887), .Z(n17) );
  XNOR U48 ( .A(n4338), .B(n17), .Z(out[268]) );
  ANDN U49 ( .B(n5006), .A(n1611), .Z(n18) );
  XNOR U50 ( .A(n1822), .B(n18), .Z(out[1091]) );
  ANDN U51 ( .B(n4830), .A(n4421), .Z(n19) );
  XNOR U52 ( .A(n4623), .B(n19), .Z(out[731]) );
  NANDN U53 ( .A(n4430), .B(n4842), .Z(n20) );
  XNOR U54 ( .A(n4635), .B(n20), .Z(out[734]) );
  NANDN U55 ( .A(n4433), .B(n4846), .Z(n21) );
  XNOR U56 ( .A(n4638), .B(n21), .Z(out[735]) );
  XNOR U57 ( .A(n1454), .B(n1027), .Z(n2776) );
  XNOR U58 ( .A(n1748), .B(n1749), .Z(n3105) );
  XNOR U59 ( .A(n1484), .B(n1153), .Z(n4058) );
  XNOR U60 ( .A(n1487), .B(n1166), .Z(n4062) );
  XNOR U61 ( .A(n1490), .B(n1181), .Z(n4066) );
  XNOR U62 ( .A(n1226), .B(n1499), .Z(n4082) );
  XNOR U63 ( .A(n1415), .B(n1688), .Z(n3173) );
  XNOR U64 ( .A(n1419), .B(n1696), .Z(n3177) );
  XNOR U65 ( .A(n1423), .B(n1704), .Z(n3181) );
  XNOR U66 ( .A(n1428), .B(n1708), .Z(n3183) );
  XNOR U67 ( .A(n1448), .B(n1754), .Z(n3213) );
  XOR U68 ( .A(n1439), .B(n1410), .Z(n4477) );
  XOR U69 ( .A(n740), .B(n1443), .Z(n4483) );
  XNOR U70 ( .A(n1463), .B(n871), .Z(n4511) );
  XOR U71 ( .A(n1479), .B(n931), .Z(n4524) );
  XOR U72 ( .A(n819), .B(n1491), .Z(n4540) );
  XNOR U73 ( .A(n3950), .B(in[1483]), .Z(n4764) );
  XNOR U74 ( .A(n3954), .B(in[1484]), .Z(n4768) );
  NAND U75 ( .A(n2895), .B(n4404), .Z(n22) );
  XNOR U76 ( .A(n2894), .B(n22), .Z(out[206]) );
  NAND U77 ( .A(n2898), .B(n4438), .Z(n23) );
  XNOR U78 ( .A(n2897), .B(n23), .Z(out[207]) );
  NAND U79 ( .A(n2904), .B(n4510), .Z(n24) );
  XNOR U80 ( .A(n2903), .B(n24), .Z(out[209]) );
  NAND U81 ( .A(n2910), .B(n4578), .Z(n25) );
  XNOR U82 ( .A(n2909), .B(n25), .Z(out[211]) );
  NANDN U83 ( .A(n2928), .B(n4689), .Z(n26) );
  XNOR U84 ( .A(n2927), .B(n26), .Z(out[216]) );
  NANDN U85 ( .A(n2931), .B(n4724), .Z(n27) );
  XNOR U86 ( .A(n2930), .B(n27), .Z(out[217]) );
  ANDN U87 ( .B(n1926), .A(n1519), .Z(n28) );
  XNOR U88 ( .A(n1768), .B(n28), .Z(out[1068]) );
  ANDN U89 ( .B(n1942), .A(n1535), .Z(n29) );
  XNOR U90 ( .A(n1778), .B(n29), .Z(out[1072]) );
  ANDN U91 ( .B(n1946), .A(n1539), .Z(n30) );
  XNOR U92 ( .A(n1780), .B(n30), .Z(out[1073]) );
  ANDN U93 ( .B(n1992), .A(n1585), .Z(n31) );
  XNOR U94 ( .A(n1804), .B(n31), .Z(out[1084]) );
  AND U95 ( .A(n4770), .B(n4769), .Z(n32) );
  XNOR U96 ( .A(n4771), .B(n32), .Z(out[90]) );
  NAND U97 ( .A(n3939), .B(n3938), .Z(n33) );
  XNOR U98 ( .A(n3940), .B(n33), .Z(out[64]) );
  ANDN U99 ( .B(n4679), .A(n4947), .Z(n34) );
  XNOR U100 ( .A(n4948), .B(n34), .Z(out[886]) );
  NANDN U101 ( .A(n4884), .B(n4661), .Z(n35) );
  XNOR U102 ( .A(n4883), .B(n35), .Z(out[872]) );
  AND U103 ( .A(n3015), .B(n3806), .Z(n36) );
  XNOR U104 ( .A(n3807), .B(n36), .Z(out[317]) );
  NANDN U105 ( .A(n2890), .B(n2889), .Z(n37) );
  XNOR U106 ( .A(n4369), .B(n37), .Z(out[269]) );
  AND U107 ( .A(n4736), .B(n4349), .Z(n38) );
  XNOR U108 ( .A(n4568), .B(n38), .Z(out[709]) );
  AND U109 ( .A(n4756), .B(n4363), .Z(n39) );
  XNOR U110 ( .A(n4583), .B(n39), .Z(out[714]) );
  ANDN U111 ( .B(n4998), .A(n1603), .Z(n40) );
  XNOR U112 ( .A(n1816), .B(n40), .Z(out[1089]) );
  ANDN U113 ( .B(n5022), .A(n1627), .Z(n41) );
  XNOR U114 ( .A(n1833), .B(n41), .Z(out[1095]) );
  ANDN U115 ( .B(n5030), .A(n1636), .Z(n42) );
  XNOR U116 ( .A(n1837), .B(n42), .Z(out[1097]) );
  ANDN U117 ( .B(n5038), .A(n1640), .Z(n43) );
  XNOR U118 ( .A(n1839), .B(n43), .Z(out[1098]) );
  AND U119 ( .A(n5067), .B(n1673), .Z(n44) );
  XNOR U120 ( .A(n1857), .B(n44), .Z(out[1106]) );
  NAND U121 ( .A(n2570), .B(n2394), .Z(n45) );
  XNOR U122 ( .A(n2571), .B(n45), .Z(out[1505]) );
  NAND U123 ( .A(n2576), .B(n2395), .Z(n46) );
  XNOR U124 ( .A(n2577), .B(n46), .Z(out[1506]) );
  NAND U125 ( .A(n2580), .B(n2396), .Z(n47) );
  XNOR U126 ( .A(n2581), .B(n47), .Z(out[1507]) );
  NANDN U127 ( .A(n4409), .B(n4811), .Z(n48) );
  XNOR U128 ( .A(n4614), .B(n48), .Z(out[727]) );
  NANDN U129 ( .A(n4453), .B(n4866), .Z(n49) );
  XNOR U130 ( .A(n4648), .B(n49), .Z(out[739]) );
  NANDN U131 ( .A(n2856), .B(n3897), .Z(n50) );
  XNOR U132 ( .A(n3019), .B(n50), .Z(out[191]) );
  ANDN U133 ( .B(n2675), .A(n2305), .Z(n51) );
  XNOR U134 ( .A(n2423), .B(n51), .Z(out[1401]) );
  XNOR U135 ( .A(n1433), .B(n1721), .Z(n2298) );
  XNOR U136 ( .A(n1503), .B(n1241), .Z(n2217) );
  XNOR U137 ( .A(n1468), .B(n1094), .Z(n2867) );
  XNOR U138 ( .A(n574), .B(n691), .Z(n4049) );
  XNOR U139 ( .A(n1482), .B(n1140), .Z(n4054) );
  XNOR U140 ( .A(n1417), .B(n1692), .Z(n3175) );
  XNOR U141 ( .A(n1662), .B(n1663), .Z(n3059) );
  XNOR U142 ( .A(n1430), .B(n1713), .Z(n3185) );
  XNOR U143 ( .A(n1683), .B(n1684), .Z(n3071) );
  XNOR U144 ( .A(n1436), .B(n1729), .Z(n3196) );
  XNOR U145 ( .A(n1695), .B(n1696), .Z(n3079) );
  XNOR U146 ( .A(n1446), .B(n1749), .Z(n4002) );
  XNOR U147 ( .A(n1744), .B(n1745), .Z(n3103) );
  XOR U148 ( .A(n725), .B(n1441), .Z(n4480) );
  XOR U149 ( .A(n856), .B(n1461), .Z(n4504) );
  XNOR U150 ( .A(n3935), .B(in[1480]), .Z(n4752) );
  XNOR U151 ( .A(n3942), .B(in[1481]), .Z(n4756) );
  XNOR U152 ( .A(n3946), .B(in[1482]), .Z(n4760) );
  XNOR U153 ( .A(n3962), .B(in[1486]), .Z(n4779) );
  AND U154 ( .A(n2004), .B(n1595), .Z(n52) );
  XNOR U155 ( .A(n1810), .B(n52), .Z(out[1087]) );
  ANDN U156 ( .B(n1954), .A(n1547), .Z(n53) );
  XNOR U157 ( .A(n1784), .B(n53), .Z(out[1075]) );
  ANDN U158 ( .B(n1984), .A(n1577), .Z(n54) );
  XNOR U159 ( .A(n1800), .B(n54), .Z(out[1082]) );
  ANDN U160 ( .B(n1996), .A(n1589), .Z(n55) );
  XNOR U161 ( .A(n1806), .B(n55), .Z(out[1085]) );
  ANDN U162 ( .B(n2000), .A(n1593), .Z(n56) );
  XNOR U163 ( .A(n1808), .B(n56), .Z(out[1086]) );
  OR U164 ( .A(n5016), .B(n1832), .Z(n57) );
  XNOR U165 ( .A(n5015), .B(n57), .Z(out[1222]) );
  NANDN U166 ( .A(n4872), .B(n4654), .Z(n58) );
  XNOR U167 ( .A(n4871), .B(n58), .Z(out[869]) );
  NANDN U168 ( .A(n4876), .B(n4659), .Z(n59) );
  XNOR U169 ( .A(n4875), .B(n59), .Z(out[870]) );
  NANDN U170 ( .A(n4888), .B(n4662), .Z(n60) );
  XNOR U171 ( .A(n4887), .B(n60), .Z(out[873]) );
  NANDN U172 ( .A(n4892), .B(n4663), .Z(n61) );
  XNOR U173 ( .A(n4891), .B(n61), .Z(out[874]) );
  ANDN U174 ( .B(n4666), .A(n4903), .Z(n62) );
  XNOR U175 ( .A(n4904), .B(n62), .Z(out[876]) );
  ANDN U176 ( .B(n4667), .A(n4907), .Z(n63) );
  XNOR U177 ( .A(n4908), .B(n63), .Z(out[877]) );
  ANDN U178 ( .B(n4668), .A(n4911), .Z(n64) );
  XNOR U179 ( .A(n4912), .B(n64), .Z(out[878]) );
  ANDN U180 ( .B(n4669), .A(n4915), .Z(n65) );
  XNOR U181 ( .A(n4916), .B(n65), .Z(out[879]) );
  ANDN U182 ( .B(n4674), .A(n4923), .Z(n66) );
  XNOR U183 ( .A(n4924), .B(n66), .Z(out[881]) );
  ANDN U184 ( .B(n4675), .A(n4927), .Z(n67) );
  XNOR U185 ( .A(n4928), .B(n67), .Z(out[882]) );
  ANDN U186 ( .B(n4677), .A(n4935), .Z(n68) );
  XNOR U187 ( .A(n4936), .B(n68), .Z(out[884]) );
  ANDN U188 ( .B(n4678), .A(n4939), .Z(n69) );
  XNOR U189 ( .A(n4940), .B(n69), .Z(out[885]) );
  AND U190 ( .A(n3420), .B(n2987), .Z(n70) );
  XNOR U191 ( .A(n3421), .B(n70), .Z(out[305]) );
  NAND U192 ( .A(n2545), .B(n2381), .Z(n71) );
  XNOR U193 ( .A(n2546), .B(n71), .Z(out[1499]) );
  NAND U194 ( .A(n4744), .B(n4355), .Z(n72) );
  XNOR U195 ( .A(n4572), .B(n72), .Z(out[711]) );
  AND U196 ( .A(n4748), .B(n4357), .Z(n73) );
  XNOR U197 ( .A(n4579), .B(n73), .Z(out[712]) );
  ANDN U198 ( .B(n4994), .A(n1599), .Z(n74) );
  XNOR U199 ( .A(n1813), .B(n74), .Z(out[1088]) );
  ANDN U200 ( .B(n5010), .A(n1615), .Z(n75) );
  XNOR U201 ( .A(n1827), .B(n75), .Z(out[1092]) );
  ANDN U202 ( .B(n5014), .A(n1619), .Z(n76) );
  XNOR U203 ( .A(n1830), .B(n76), .Z(out[1093]) );
  ANDN U204 ( .B(n5046), .A(n1648), .Z(n77) );
  XNOR U205 ( .A(n1843), .B(n77), .Z(out[1100]) );
  ANDN U206 ( .B(n5050), .A(n1652), .Z(n78) );
  XNOR U207 ( .A(n1845), .B(n78), .Z(out[1101]) );
  ANDN U208 ( .B(n5054), .A(n1656), .Z(n79) );
  XNOR U209 ( .A(n1849), .B(n79), .Z(out[1102]) );
  AND U210 ( .A(n5061), .B(n1664), .Z(n80) );
  XNOR U211 ( .A(n1853), .B(n80), .Z(out[1104]) );
  AND U212 ( .A(n5064), .B(n1668), .Z(n81) );
  XNOR U213 ( .A(n1855), .B(n81), .Z(out[1105]) );
  ANDN U214 ( .B(n5071), .A(n1677), .Z(n82) );
  XNOR U215 ( .A(n1859), .B(n82), .Z(out[1107]) );
  ANDN U216 ( .B(n5093), .A(n1701), .Z(n83) );
  XNOR U217 ( .A(n1873), .B(n83), .Z(out[1113]) );
  ANDN U218 ( .B(n5096), .A(n1705), .Z(n84) );
  XNOR U219 ( .A(n1875), .B(n84), .Z(out[1114]) );
  NAND U220 ( .A(n2584), .B(n2397), .Z(n85) );
  XNOR U221 ( .A(n2585), .B(n85), .Z(out[1508]) );
  NANDN U222 ( .A(n4424), .B(n4834), .Z(n86) );
  XNOR U223 ( .A(n4629), .B(n86), .Z(out[732]) );
  NANDN U224 ( .A(n2852), .B(n3809), .Z(n87) );
  XNOR U225 ( .A(n3015), .B(n87), .Z(out[189]) );
  NANDN U226 ( .A(n2854), .B(n3853), .Z(n88) );
  XNOR U227 ( .A(n3016), .B(n88), .Z(out[190]) );
  OR U228 ( .A(n5085), .B(n5086), .Z(n89) );
  XNOR U229 ( .A(n5087), .B(n89), .Z(out[983]) );
  ANDN U230 ( .B(n2515), .A(n2224), .Z(n90) );
  XNOR U231 ( .A(n2365), .B(n90), .Z(out[1363]) );
  ANDN U232 ( .B(n2527), .A(n2231), .Z(n91) );
  XNOR U233 ( .A(n2371), .B(n91), .Z(out[1366]) );
  OR U234 ( .A(n5111), .B(n5112), .Z(n92) );
  XNOR U235 ( .A(n5113), .B(n92), .Z(out[990]) );
  ANDN U236 ( .B(n2544), .A(n2239), .Z(n93) );
  XNOR U237 ( .A(n2379), .B(n93), .Z(out[1370]) );
  ANDN U238 ( .B(n2569), .A(n2252), .Z(n94) );
  XNOR U239 ( .A(n2392), .B(n94), .Z(out[1376]) );
  NANDN U240 ( .A(n3282), .B(n3643), .Z(n95) );
  XNOR U241 ( .A(n3475), .B(n95), .Z(out[390]) );
  ANDN U242 ( .B(n2440), .A(n2439), .Z(n96) );
  XNOR U243 ( .A(n2441), .B(round_const[0]), .Z(n97) );
  XOR U244 ( .A(n96), .B(n97), .Z(out[1536]) );
  XNOR U245 ( .A(n1712), .B(n1356), .Z(n3931) );
  XNOR U246 ( .A(n1464), .B(n1079), .Z(n2843) );
  XNOR U247 ( .A(n1493), .B(n1196), .Z(n4074) );
  XNOR U248 ( .A(n1411), .B(n1684), .Z(n3171) );
  XNOR U249 ( .A(n1421), .B(n1700), .Z(n3179) );
  XNOR U250 ( .A(n1666), .B(n1667), .Z(n3061) );
  XNOR U251 ( .A(n1671), .B(n1672), .Z(n3063) );
  XNOR U252 ( .A(n1679), .B(n1680), .Z(n3068) );
  XNOR U253 ( .A(n1687), .B(n1688), .Z(n3073) );
  XNOR U254 ( .A(n1691), .B(n1692), .Z(n3077) );
  XNOR U255 ( .A(n1442), .B(n1745), .Z(n3208) );
  XNOR U256 ( .A(n1720), .B(n1721), .Z(n3090) );
  XNOR U257 ( .A(n1732), .B(n1733), .Z(n3098) );
  XNOR U258 ( .A(n1736), .B(n1737), .Z(n3100) );
  XOR U259 ( .A(n1455), .B(n826), .Z(n4498) );
  XOR U260 ( .A(n841), .B(n1457), .Z(n4501) );
  XNOR U261 ( .A(n1465), .B(n886), .Z(n4514) );
  XNOR U262 ( .A(n1469), .B(n901), .Z(n4517) );
  XOR U263 ( .A(n1485), .B(n691), .Z(n4532) );
  XNOR U264 ( .A(n3966), .B(in[1487]), .Z(n4783) );
  XNOR U265 ( .A(n3970), .B(in[1488]), .Z(n4787) );
  XNOR U266 ( .A(n3978), .B(in[1490]), .Z(n4795) );
  NAND U267 ( .A(n2907), .B(n4549), .Z(n98) );
  XNOR U268 ( .A(n2906), .B(n98), .Z(out[210]) );
  NANDN U269 ( .A(n2916), .B(n4628), .Z(n99) );
  XNOR U270 ( .A(n2915), .B(n99), .Z(out[213]) );
  ANDN U271 ( .B(n2955), .A(n5152), .Z(n100) );
  XNOR U272 ( .A(n3096), .B(n100), .Z(out[227]) );
  ANDN U273 ( .B(n1930), .A(n1523), .Z(n101) );
  XNOR U274 ( .A(n1770), .B(n101), .Z(out[1069]) );
  ANDN U275 ( .B(n1934), .A(n1527), .Z(n102) );
  XNOR U276 ( .A(n1772), .B(n102), .Z(out[1070]) );
  ANDN U277 ( .B(n1938), .A(n1531), .Z(n103) );
  XNOR U278 ( .A(n1774), .B(n103), .Z(out[1071]) );
  ANDN U279 ( .B(n4673), .A(n4919), .Z(n104) );
  XNOR U280 ( .A(n4920), .B(n104), .Z(out[880]) );
  ANDN U281 ( .B(n4676), .A(n4931), .Z(n105) );
  XNOR U282 ( .A(n4932), .B(n105), .Z(out[883]) );
  AND U283 ( .A(n2604), .B(n2403), .Z(n106) );
  XNOR U284 ( .A(n2605), .B(n106), .Z(out[1513]) );
  NAND U285 ( .A(n2608), .B(n2404), .Z(n107) );
  XNOR U286 ( .A(n2609), .B(n107), .Z(out[1514]) );
  NANDN U287 ( .A(n4456), .B(n4870), .Z(n108) );
  XNOR U288 ( .A(n4651), .B(n108), .Z(out[740]) );
  NANDN U289 ( .A(n4459), .B(n4874), .Z(n109) );
  XNOR U290 ( .A(n4654), .B(n109), .Z(out[741]) );
  NANDN U291 ( .A(n4462), .B(n4878), .Z(n110) );
  XNOR U292 ( .A(n4659), .B(n110), .Z(out[742]) );
  ANDN U293 ( .B(n5026), .A(n1632), .Z(n111) );
  XNOR U294 ( .A(n1835), .B(n111), .Z(out[1096]) );
  NAND U295 ( .A(n2496), .B(n2357), .Z(n112) );
  XNOR U296 ( .A(n2495), .B(n112), .Z(out[1487]) );
  NAND U297 ( .A(n2501), .B(n2359), .Z(n113) );
  XNOR U298 ( .A(n2500), .B(n113), .Z(out[1488]) );
  AND U299 ( .A(n5058), .B(n1660), .Z(n114) );
  XNOR U300 ( .A(n1851), .B(n114), .Z(out[1103]) );
  ANDN U301 ( .B(n5078), .A(n1681), .Z(n115) );
  XNOR U302 ( .A(n1861), .B(n115), .Z(out[1108]) );
  ANDN U303 ( .B(n5084), .A(n1689), .Z(n116) );
  XNOR U304 ( .A(n1865), .B(n116), .Z(out[1110]) );
  AND U305 ( .A(n2612), .B(n2405), .Z(n117) );
  XNOR U306 ( .A(n2613), .B(n117), .Z(out[1515]) );
  AND U307 ( .A(n2664), .B(n2421), .Z(n118) );
  XNOR U308 ( .A(n2665), .B(n118), .Z(out[1527]) );
  NANDN U309 ( .A(n4444), .B(n4850), .Z(n119) );
  XNOR U310 ( .A(n4639), .B(n119), .Z(out[736]) );
  NANDN U311 ( .A(n4447), .B(n4854), .Z(n120) );
  XNOR U312 ( .A(n4642), .B(n120), .Z(out[737]) );
  NANDN U313 ( .A(n4450), .B(n4862), .Z(n121) );
  XNOR U314 ( .A(n4645), .B(n121), .Z(out[738]) );
  ANDN U315 ( .B(n2556), .A(n2245), .Z(n122) );
  XNOR U316 ( .A(n2386), .B(n122), .Z(out[1373]) );
  ANDN U317 ( .B(n3505), .A(n3700), .Z(n123) );
  XNOR U318 ( .A(n3701), .B(n123), .Z(out[532]) );
  ANDN U319 ( .B(n3507), .A(n3708), .Z(n124) );
  XNOR U320 ( .A(n3709), .B(n124), .Z(out[534]) );
  ANDN U321 ( .B(n3508), .A(n3712), .Z(n125) );
  XNOR U322 ( .A(n3713), .B(n125), .Z(out[535]) );
  ANDN U323 ( .B(n3509), .A(n3722), .Z(n126) );
  XNOR U324 ( .A(n3723), .B(n126), .Z(out[536]) );
  ANDN U325 ( .B(n3513), .A(n3734), .Z(n127) );
  XNOR U326 ( .A(n3735), .B(n127), .Z(out[539]) );
  ANDN U327 ( .B(n2649), .A(n2291), .Z(n128) );
  XNOR U328 ( .A(n2414), .B(n128), .Z(out[1395]) );
  ANDN U329 ( .B(n2653), .A(n2294), .Z(n129) );
  XNOR U330 ( .A(n2416), .B(n129), .Z(out[1396]) );
  ANDN U331 ( .B(n2657), .A(n2296), .Z(n130) );
  XNOR U332 ( .A(n2418), .B(n130), .Z(out[1397]) );
  OR U333 ( .A(n5079), .B(n5080), .Z(n131) );
  XNOR U334 ( .A(n5081), .B(n131), .Z(out[981]) );
  OR U335 ( .A(n5088), .B(n5089), .Z(n132) );
  XNOR U336 ( .A(n5090), .B(n132), .Z(out[984]) );
  OR U337 ( .A(n5091), .B(n5092), .Z(n133) );
  XNOR U338 ( .A(n5093), .B(n133), .Z(out[985]) );
  OR U339 ( .A(n5094), .B(n5095), .Z(n134) );
  XNOR U340 ( .A(n5096), .B(n134), .Z(out[986]) );
  OR U341 ( .A(n5097), .B(n5098), .Z(n135) );
  XNOR U342 ( .A(n5099), .B(n135), .Z(out[987]) );
  OR U343 ( .A(n5104), .B(n5105), .Z(n136) );
  XNOR U344 ( .A(n5106), .B(n136), .Z(out[989]) );
  NOR U345 ( .A(n5138), .B(n5139), .Z(n137) );
  XNOR U346 ( .A(n5140), .B(n137), .Z(out[997]) );
  ANDN U347 ( .B(n2466), .A(n2465), .Z(n138) );
  XNOR U348 ( .A(n2464), .B(n138), .Z(out[1542]) );
  NAND U349 ( .A(n3837), .B(n3415), .Z(n139) );
  XNOR U350 ( .A(n3414), .B(n139), .Z(out[434]) );
  NANDN U351 ( .A(n3444), .B(n3873), .Z(n140) );
  XNOR U352 ( .A(n3602), .B(n140), .Z(out[442]) );
  NANDN U353 ( .A(n3447), .B(n3877), .Z(n141) );
  XNOR U354 ( .A(n3603), .B(n141), .Z(out[443]) );
  ANDN U355 ( .B(n3893), .A(n3463), .Z(n142) );
  XNOR U356 ( .A(n3610), .B(n142), .Z(out[447]) );
  NANDN U357 ( .A(n3276), .B(n3635), .Z(n143) );
  XNOR U358 ( .A(n3473), .B(n143), .Z(out[388]) );
  NANDN U359 ( .A(n3279), .B(n3639), .Z(n144) );
  XNOR U360 ( .A(n3474), .B(n144), .Z(out[389]) );
  NANDN U361 ( .A(n3285), .B(n3647), .Z(n145) );
  XNOR U362 ( .A(n3476), .B(n145), .Z(out[391]) );
  NANDN U363 ( .A(n3288), .B(n3651), .Z(n146) );
  XNOR U364 ( .A(n3481), .B(n146), .Z(out[392]) );
  ANDN U365 ( .B(n2472), .A(n2471), .Z(n147) );
  XNOR U366 ( .A(n2470), .B(n147), .Z(out[1544]) );
  ANDN U367 ( .B(n2475), .A(n2474), .Z(n148) );
  XNOR U368 ( .A(n2473), .B(n148), .Z(out[1545]) );
  ANDN U369 ( .B(n2478), .A(n2477), .Z(n149) );
  XNOR U370 ( .A(n2476), .B(n149), .Z(out[1546]) );
  NOR U371 ( .A(n4696), .B(n4545), .Z(n150) );
  XNOR U372 ( .A(n4975), .B(n150), .Z(out[829]) );
  NOR U373 ( .A(n4699), .B(n4551), .Z(n151) );
  XNOR U374 ( .A(n4979), .B(n151), .Z(out[830]) );
  NOR U375 ( .A(n4702), .B(n4553), .Z(n152) );
  XNOR U376 ( .A(n4983), .B(n152), .Z(out[831]) );
  NOR U377 ( .A(n4554), .B(n4334), .Z(n153) );
  XNOR U378 ( .A(n4705), .B(n153), .Z(out[768]) );
  NOR U379 ( .A(n4557), .B(n4336), .Z(n154) );
  XNOR U380 ( .A(n4709), .B(n154), .Z(out[769]) );
  NOR U381 ( .A(n4560), .B(n4342), .Z(n155) );
  XNOR U382 ( .A(n4713), .B(n155), .Z(out[770]) );
  NOR U383 ( .A(n4563), .B(n4344), .Z(n156) );
  XNOR U384 ( .A(n4717), .B(n156), .Z(out[771]) );
  NOR U385 ( .A(n4572), .B(n4355), .Z(n157) );
  XNOR U386 ( .A(n4741), .B(n157), .Z(out[775]) );
  NOR U387 ( .A(n4595), .B(n4385), .Z(n158) );
  XNOR U388 ( .A(n4781), .B(n158), .Z(out[784]) );
  ANDN U389 ( .B(n2697), .A(n2696), .Z(n159) );
  XNOR U390 ( .A(n2698), .B(round_const_7), .Z(n160) );
  XOR U391 ( .A(n159), .B(n160), .Z(out[1599]) );
  XNOR U392 ( .A(n1478), .B(n1127), .Z(n2924) );
  XNOR U393 ( .A(n1496), .B(n1211), .Z(n4078) );
  XNOR U394 ( .A(n1440), .B(n1741), .Z(n3205) );
  XNOR U395 ( .A(n1699), .B(n1700), .Z(n3081) );
  XNOR U396 ( .A(n1703), .B(n1704), .Z(n3083) );
  XNOR U397 ( .A(n1707), .B(n1708), .Z(n3085) );
  XNOR U398 ( .A(n1724), .B(n1725), .Z(n3092) );
  XNOR U399 ( .A(n1728), .B(n1729), .Z(n3094) );
  XNOR U400 ( .A(n1753), .B(n1754), .Z(n3107) );
  XNOR U401 ( .A(n1757), .B(n1758), .Z(n3109) );
  XOR U402 ( .A(n1437), .B(n1402), .Z(n4467) );
  XOR U403 ( .A(n770), .B(n1449), .Z(n4489) );
  XOR U404 ( .A(n785), .B(n1451), .Z(n4492) );
  XOR U405 ( .A(n1475), .B(n916), .Z(n4520) );
  XOR U406 ( .A(n1483), .B(n946), .Z(n4528) );
  XOR U407 ( .A(n708), .B(n1488), .Z(n4536) );
  XNOR U408 ( .A(n3958), .B(in[1485]), .Z(n4775) );
  NAND U409 ( .A(n2913), .B(n4603), .Z(n161) );
  XNOR U410 ( .A(n2912), .B(n161), .Z(out[212]) );
  ANDN U411 ( .B(n1916), .A(n1511), .Z(n162) );
  XNOR U412 ( .A(n1765), .B(n162), .Z(out[1066]) );
  ANDN U413 ( .B(n1988), .A(n1581), .Z(n163) );
  XNOR U414 ( .A(n1802), .B(n163), .Z(out[1083]) );
  NAND U415 ( .A(n2592), .B(n2400), .Z(n164) );
  XNOR U416 ( .A(n2593), .B(n164), .Z(out[1510]) );
  AND U417 ( .A(n2596), .B(n2401), .Z(n165) );
  XNOR U418 ( .A(n2597), .B(n165), .Z(out[1511]) );
  AND U419 ( .A(n2600), .B(n2402), .Z(n166) );
  XNOR U420 ( .A(n2601), .B(n166), .Z(out[1512]) );
  NANDN U421 ( .A(n2886), .B(n2885), .Z(n167) );
  XNOR U422 ( .A(n4306), .B(n167), .Z(out[267]) );
  AND U423 ( .A(n4752), .B(n4360), .Z(n168) );
  XNOR U424 ( .A(n4581), .B(n168), .Z(out[713]) );
  AND U425 ( .A(n4760), .B(n4366), .Z(n169) );
  XNOR U426 ( .A(n4585), .B(n169), .Z(out[715]) );
  ANDN U427 ( .B(n5002), .A(n1607), .Z(n170) );
  XNOR U428 ( .A(n1819), .B(n170), .Z(out[1090]) );
  ANDN U429 ( .B(n5018), .A(n1623), .Z(n171) );
  XNOR U430 ( .A(n1832), .B(n171), .Z(out[1094]) );
  ANDN U431 ( .B(n5042), .A(n1644), .Z(n172) );
  XNOR U432 ( .A(n1841), .B(n172), .Z(out[1099]) );
  ANDN U433 ( .B(n5081), .A(n1685), .Z(n173) );
  XNOR U434 ( .A(n1863), .B(n173), .Z(out[1109]) );
  ANDN U435 ( .B(n5087), .A(n1693), .Z(n174) );
  XNOR U436 ( .A(n1867), .B(n174), .Z(out[1111]) );
  ANDN U437 ( .B(n5090), .A(n1697), .Z(n175) );
  XNOR U438 ( .A(n1871), .B(n175), .Z(out[1112]) );
  ANDN U439 ( .B(n5103), .A(n1714), .Z(n176) );
  XNOR U440 ( .A(n1879), .B(n176), .Z(out[1116]) );
  ANDN U441 ( .B(n5106), .A(n1718), .Z(n177) );
  XNOR U442 ( .A(n1881), .B(n177), .Z(out[1117]) );
  AND U443 ( .A(n4764), .B(n4373), .Z(n178) );
  XNOR U444 ( .A(n4587), .B(n178), .Z(out[716]) );
  NAND U445 ( .A(n2588), .B(n2398), .Z(n179) );
  XNOR U446 ( .A(n2589), .B(n179), .Z(out[1509]) );
  ANDN U447 ( .B(n5129), .A(n1738), .Z(n180) );
  XNOR U448 ( .A(n1893), .B(n180), .Z(out[1122]) );
  AND U449 ( .A(n2618), .B(n2406), .Z(n181) );
  XNOR U450 ( .A(n2619), .B(n181), .Z(out[1516]) );
  ANDN U451 ( .B(n2407), .A(n2622), .Z(n182) );
  XNOR U452 ( .A(n2623), .B(n182), .Z(out[1517]) );
  AND U453 ( .A(n2626), .B(n2408), .Z(n183) );
  XNOR U454 ( .A(n2627), .B(n183), .Z(out[1518]) );
  AND U455 ( .A(n2630), .B(n2409), .Z(n184) );
  XNOR U456 ( .A(n2631), .B(n184), .Z(out[1519]) );
  AND U457 ( .A(n2634), .B(n2411), .Z(n185) );
  XNOR U458 ( .A(n2635), .B(n185), .Z(out[1520]) );
  ANDN U459 ( .B(n4818), .A(n4412), .Z(n186) );
  XNOR U460 ( .A(n4617), .B(n186), .Z(out[728]) );
  AND U461 ( .A(n2638), .B(n2412), .Z(n187) );
  XNOR U462 ( .A(n2639), .B(n187), .Z(out[1521]) );
  AND U463 ( .A(n2642), .B(n2413), .Z(n188) );
  XNOR U464 ( .A(n2643), .B(n188), .Z(out[1522]) );
  NANDN U465 ( .A(n4427), .B(n4838), .Z(n189) );
  XNOR U466 ( .A(n4632), .B(n189), .Z(out[733]) );
  AND U467 ( .A(n2660), .B(n2420), .Z(n190) );
  XNOR U468 ( .A(n2661), .B(n190), .Z(out[1526]) );
  AND U469 ( .A(n2668), .B(n2422), .Z(n191) );
  XNOR U470 ( .A(n2669), .B(n191), .Z(out[1528]) );
  NANDN U471 ( .A(n2241), .B(n2548), .Z(n192) );
  XNOR U472 ( .A(n2381), .B(n192), .Z(out[1371]) );
  ANDN U473 ( .B(n2552), .A(n2243), .Z(n193) );
  XNOR U474 ( .A(n2384), .B(n193), .Z(out[1372]) );
  ANDN U475 ( .B(n3504), .A(n3696), .Z(n194) );
  XNOR U476 ( .A(n3697), .B(n194), .Z(out[531]) );
  ANDN U477 ( .B(n3506), .A(n3704), .Z(n195) );
  XNOR U478 ( .A(n3705), .B(n195), .Z(out[533]) );
  ANDN U479 ( .B(n3510), .A(n3726), .Z(n196) );
  XNOR U480 ( .A(n3727), .B(n196), .Z(out[537]) );
  NAND U481 ( .A(n3602), .B(n3871), .Z(n197) );
  XNOR U482 ( .A(n3870), .B(n197), .Z(out[570]) );
  NAND U483 ( .A(n3603), .B(n3875), .Z(n198) );
  XNOR U484 ( .A(n3874), .B(n198), .Z(out[571]) );
  NAND U485 ( .A(n3473), .B(n3633), .Z(n199) );
  XNOR U486 ( .A(n3632), .B(n199), .Z(out[516]) );
  NANDN U487 ( .A(n3637), .B(n3474), .Z(n200) );
  XNOR U488 ( .A(n3636), .B(n200), .Z(out[517]) );
  NANDN U489 ( .A(n3641), .B(n3475), .Z(n201) );
  XNOR U490 ( .A(n3640), .B(n201), .Z(out[518]) );
  NANDN U491 ( .A(n3645), .B(n3476), .Z(n202) );
  XNOR U492 ( .A(n3644), .B(n202), .Z(out[519]) );
  NAND U493 ( .A(n3481), .B(n3649), .Z(n203) );
  XNOR U494 ( .A(n3648), .B(n203), .Z(out[520]) );
  ANDN U495 ( .B(n3498), .A(n3688), .Z(n204) );
  XNOR U496 ( .A(n3689), .B(n204), .Z(out[529]) );
  ANDN U497 ( .B(n3503), .A(n3692), .Z(n205) );
  XNOR U498 ( .A(n3693), .B(n205), .Z(out[530]) );
  ANDN U499 ( .B(n2679), .A(n2307), .Z(n206) );
  XNOR U500 ( .A(n2426), .B(n206), .Z(out[1402]) );
  OR U501 ( .A(n5059), .B(n5060), .Z(n207) );
  XNOR U502 ( .A(n5061), .B(n207), .Z(out[976]) );
  OR U503 ( .A(n5062), .B(n5063), .Z(n208) );
  XNOR U504 ( .A(n5064), .B(n208), .Z(out[977]) );
  OR U505 ( .A(n5065), .B(n5066), .Z(n209) );
  XNOR U506 ( .A(n5067), .B(n209), .Z(out[978]) );
  OR U507 ( .A(n5076), .B(n5077), .Z(n210) );
  XNOR U508 ( .A(n5078), .B(n210), .Z(out[980]) );
  ANDN U509 ( .B(n2494), .A(n2213), .Z(n211) );
  XNOR U510 ( .A(n2355), .B(n211), .Z(out[1358]) );
  OR U511 ( .A(n5082), .B(n5083), .Z(n212) );
  XNOR U512 ( .A(n5084), .B(n212), .Z(out[982]) );
  NANDN U513 ( .A(n2215), .B(n2497), .Z(n213) );
  XNOR U514 ( .A(n2357), .B(n213), .Z(out[1359]) );
  NANDN U515 ( .A(n2218), .B(n2503), .Z(n214) );
  XNOR U516 ( .A(n2359), .B(n214), .Z(out[1360]) );
  ANDN U517 ( .B(n2531), .A(n2233), .Z(n215) );
  XNOR U518 ( .A(n2373), .B(n215), .Z(out[1367]) );
  ANDN U519 ( .B(n2560), .A(n2247), .Z(n216) );
  XNOR U520 ( .A(n2388), .B(n216), .Z(out[1374]) );
  ANDN U521 ( .B(n2563), .A(n2249), .Z(n217) );
  XNOR U522 ( .A(n2390), .B(n217), .Z(out[1375]) );
  ANDN U523 ( .B(n2449), .A(n2448), .Z(n218) );
  XNOR U524 ( .A(n2447), .B(n218), .Z(out[1538]) );
  ANDN U525 ( .B(n2468), .A(n2467), .Z(n219) );
  XNOR U526 ( .A(n2469), .B(round_const_7), .Z(n220) );
  XOR U527 ( .A(n219), .B(n220), .Z(out[1543]) );
  NAND U528 ( .A(n3841), .B(n3418), .Z(n221) );
  XNOR U529 ( .A(n3417), .B(n221), .Z(out[435]) );
  ANDN U530 ( .B(n3845), .A(n3426), .Z(n222) );
  XNOR U531 ( .A(n3586), .B(n222), .Z(out[436]) );
  ANDN U532 ( .B(n3849), .A(n3429), .Z(n223) );
  XNOR U533 ( .A(n3588), .B(n223), .Z(out[437]) );
  ANDN U534 ( .B(n3857), .A(n3432), .Z(n224) );
  XNOR U535 ( .A(n3590), .B(n224), .Z(out[438]) );
  ANDN U536 ( .B(n3861), .A(n3435), .Z(n225) );
  XNOR U537 ( .A(n3592), .B(n225), .Z(out[439]) );
  ANDN U538 ( .B(n3865), .A(n3438), .Z(n226) );
  XNOR U539 ( .A(n3594), .B(n226), .Z(out[440]) );
  ANDN U540 ( .B(n3869), .A(n3441), .Z(n227) );
  XNOR U541 ( .A(n3596), .B(n227), .Z(out[441]) );
  ANDN U542 ( .B(n3881), .A(n3450), .Z(n228) );
  XNOR U543 ( .A(n3604), .B(n228), .Z(out[444]) );
  ANDN U544 ( .B(n3885), .A(n3453), .Z(n229) );
  XNOR U545 ( .A(n3606), .B(n229), .Z(out[445]) );
  AND U546 ( .A(n3889), .B(n3460), .Z(n230) );
  XNOR U547 ( .A(n3608), .B(n230), .Z(out[446]) );
  ANDN U548 ( .B(n3615), .A(n3260), .Z(n231) );
  XNOR U549 ( .A(n3465), .B(n231), .Z(out[384]) );
  ANDN U550 ( .B(n2485), .A(n2484), .Z(n232) );
  XNOR U551 ( .A(n2483), .B(n232), .Z(out[1548]) );
  NANDN U552 ( .A(n1918), .B(n1767), .Z(n233) );
  XNOR U553 ( .A(n1917), .B(n233), .Z(out[1195]) );
  XNOR U554 ( .A(in[1162]), .B(n848), .Z(n234) );
  XNOR U555 ( .A(in[1164]), .B(n878), .Z(n235) );
  XNOR U556 ( .A(in[1166]), .B(n908), .Z(n236) );
  XNOR U557 ( .A(in[1167]), .B(n923), .Z(n237) );
  XOR U558 ( .A(in[1469]), .B(in[509]), .Z(n239) );
  XNOR U559 ( .A(in[829]), .B(in[189]), .Z(n238) );
  XNOR U560 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U561 ( .A(in[1149]), .B(n240), .Z(n1109) );
  XOR U562 ( .A(in[1598]), .B(in[638]), .Z(n242) );
  XNOR U563 ( .A(in[958]), .B(in[318]), .Z(n241) );
  XNOR U564 ( .A(n242), .B(n241), .Z(n243) );
  XNOR U565 ( .A(in[1278]), .B(n243), .Z(n1676) );
  XNOR U566 ( .A(n1109), .B(n1676), .Z(n3287) );
  XOR U567 ( .A(in[254]), .B(n3287), .Z(n3938) );
  XOR U568 ( .A(in[1345]), .B(in[65]), .Z(n245) );
  XNOR U569 ( .A(in[1025]), .B(in[385]), .Z(n244) );
  XNOR U570 ( .A(n245), .B(n244), .Z(n246) );
  XNOR U571 ( .A(in[705]), .B(n246), .Z(n1684) );
  XOR U572 ( .A(in[1474]), .B(in[514]), .Z(n248) );
  XNOR U573 ( .A(in[834]), .B(in[194]), .Z(n247) );
  XNOR U574 ( .A(n248), .B(n247), .Z(n249) );
  XOR U575 ( .A(in[1154]), .B(n249), .Z(n1411) );
  XOR U576 ( .A(in[1410]), .B(n3171), .Z(n3939) );
  XOR U577 ( .A(in[137]), .B(in[457]), .Z(n251) );
  XNOR U578 ( .A(in[777]), .B(in[1417]), .Z(n250) );
  XNOR U579 ( .A(n251), .B(n250), .Z(n252) );
  XNOR U580 ( .A(in[1097]), .B(n252), .Z(n1368) );
  XOR U581 ( .A(in[328]), .B(in[8]), .Z(n254) );
  XNOR U582 ( .A(in[968]), .B(in[648]), .Z(n253) );
  XNOR U583 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U584 ( .A(in[1288]), .B(n255), .Z(n1424) );
  XOR U585 ( .A(n1368), .B(n1424), .Z(n4449) );
  XNOR U586 ( .A(in[1033]), .B(n4449), .Z(n2859) );
  OR U587 ( .A(n3939), .B(n2859), .Z(n256) );
  XOR U588 ( .A(n3938), .B(n256), .Z(out[0]) );
  XOR U589 ( .A(in[1515]), .B(in[555]), .Z(n258) );
  XNOR U590 ( .A(in[875]), .B(in[235]), .Z(n257) );
  XNOR U591 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U592 ( .A(in[1195]), .B(n259), .Z(n1530) );
  XOR U593 ( .A(in[1386]), .B(in[106]), .Z(n261) );
  XNOR U594 ( .A(in[1066]), .B(in[746]), .Z(n260) );
  XNOR U595 ( .A(n261), .B(n260), .Z(n262) );
  XNOR U596 ( .A(in[426]), .B(n262), .Z(n712) );
  XOR U597 ( .A(n1530), .B(n712), .Z(n4109) );
  XOR U598 ( .A(in[171]), .B(n4109), .Z(n1501) );
  XOR U599 ( .A(in[140]), .B(in[460]), .Z(n264) );
  XNOR U600 ( .A(in[1100]), .B(in[1420]), .Z(n263) );
  XNOR U601 ( .A(n264), .B(n263), .Z(n265) );
  XNOR U602 ( .A(in[780]), .B(n265), .Z(n1390) );
  XOR U603 ( .A(in[971]), .B(in[1291]), .Z(n267) );
  XNOR U604 ( .A(in[11]), .B(in[331]), .Z(n266) );
  XNOR U605 ( .A(n267), .B(n266), .Z(n268) );
  XOR U606 ( .A(in[651]), .B(n268), .Z(n1432) );
  XNOR U607 ( .A(in[1356]), .B(n4458), .Z(n1908) );
  XOR U608 ( .A(in[1364]), .B(in[724]), .Z(n270) );
  XNOR U609 ( .A(in[84]), .B(in[404]), .Z(n269) );
  XNOR U610 ( .A(n270), .B(n269), .Z(n271) );
  XNOR U611 ( .A(in[1044]), .B(n271), .Z(n1014) );
  XOR U612 ( .A(in[1555]), .B(in[595]), .Z(n273) );
  XNOR U613 ( .A(in[915]), .B(in[275]), .Z(n272) );
  XNOR U614 ( .A(n273), .B(n272), .Z(n274) );
  XNOR U615 ( .A(in[1235]), .B(n274), .Z(n726) );
  XOR U616 ( .A(n1014), .B(n726), .Z(n4248) );
  XOR U617 ( .A(in[980]), .B(n4248), .Z(n1905) );
  NANDN U618 ( .A(n1908), .B(n1905), .Z(n275) );
  XNOR U619 ( .A(n1501), .B(n275), .Z(out[1000]) );
  XOR U620 ( .A(in[1516]), .B(in[556]), .Z(n277) );
  XNOR U621 ( .A(in[876]), .B(in[236]), .Z(n276) );
  XNOR U622 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U623 ( .A(in[1196]), .B(n278), .Z(n1534) );
  XOR U624 ( .A(in[1387]), .B(in[107]), .Z(n280) );
  XNOR U625 ( .A(in[1067]), .B(in[747]), .Z(n279) );
  XNOR U626 ( .A(n280), .B(n279), .Z(n281) );
  XNOR U627 ( .A(in[427]), .B(n281), .Z(n723) );
  XOR U628 ( .A(n1534), .B(n723), .Z(n4117) );
  XOR U629 ( .A(in[172]), .B(n4117), .Z(n1505) );
  XOR U630 ( .A(in[972]), .B(in[12]), .Z(n283) );
  XNOR U631 ( .A(in[1292]), .B(in[332]), .Z(n282) );
  XNOR U632 ( .A(n283), .B(n282), .Z(n284) );
  XNOR U633 ( .A(in[652]), .B(n284), .Z(n1434) );
  XOR U634 ( .A(in[141]), .B(in[461]), .Z(n286) );
  XNOR U635 ( .A(in[1101]), .B(in[1421]), .Z(n285) );
  XNOR U636 ( .A(n286), .B(n285), .Z(n287) );
  XOR U637 ( .A(in[781]), .B(n287), .Z(n1394) );
  XNOR U638 ( .A(in[1357]), .B(n4461), .Z(n1912) );
  XOR U639 ( .A(in[1365]), .B(in[725]), .Z(n289) );
  XNOR U640 ( .A(in[85]), .B(in[405]), .Z(n288) );
  XNOR U641 ( .A(n289), .B(n288), .Z(n290) );
  XNOR U642 ( .A(in[1045]), .B(n290), .Z(n1027) );
  XOR U643 ( .A(in[1556]), .B(in[596]), .Z(n292) );
  XNOR U644 ( .A(in[916]), .B(in[276]), .Z(n291) );
  XNOR U645 ( .A(n292), .B(n291), .Z(n293) );
  XNOR U646 ( .A(in[1236]), .B(n293), .Z(n741) );
  XOR U647 ( .A(n1027), .B(n741), .Z(n4249) );
  XOR U648 ( .A(in[981]), .B(n4249), .Z(n1909) );
  NANDN U649 ( .A(n1912), .B(n1909), .Z(n294) );
  XNOR U650 ( .A(n1505), .B(n294), .Z(out[1001]) );
  XOR U651 ( .A(in[1388]), .B(in[108]), .Z(n296) );
  XNOR U652 ( .A(in[1068]), .B(in[748]), .Z(n295) );
  XNOR U653 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U654 ( .A(in[428]), .B(n297), .Z(n1598) );
  XOR U655 ( .A(in[1517]), .B(in[557]), .Z(n299) );
  XNOR U656 ( .A(in[877]), .B(in[237]), .Z(n298) );
  XNOR U657 ( .A(n299), .B(n298), .Z(n300) );
  XNOR U658 ( .A(in[1197]), .B(n300), .Z(n1538) );
  XOR U659 ( .A(n1598), .B(n1538), .Z(n1373) );
  XOR U660 ( .A(in[173]), .B(n1373), .Z(n1511) );
  XOR U661 ( .A(in[142]), .B(in[1422]), .Z(n302) );
  XNOR U662 ( .A(in[1102]), .B(in[782]), .Z(n301) );
  XNOR U663 ( .A(n302), .B(n301), .Z(n303) );
  XNOR U664 ( .A(in[462]), .B(n303), .Z(n1398) );
  XOR U665 ( .A(in[973]), .B(in[13]), .Z(n305) );
  XNOR U666 ( .A(in[1293]), .B(in[333]), .Z(n304) );
  XNOR U667 ( .A(n305), .B(n304), .Z(n306) );
  XOR U668 ( .A(in[653]), .B(n306), .Z(n1435) );
  XNOR U669 ( .A(in[1358]), .B(n4464), .Z(n1916) );
  XOR U670 ( .A(in[1366]), .B(in[726]), .Z(n308) );
  XNOR U671 ( .A(in[86]), .B(in[406]), .Z(n307) );
  XNOR U672 ( .A(n308), .B(n307), .Z(n309) );
  XNOR U673 ( .A(in[1046]), .B(n309), .Z(n1040) );
  XOR U674 ( .A(in[1557]), .B(in[597]), .Z(n311) );
  XNOR U675 ( .A(in[917]), .B(in[277]), .Z(n310) );
  XNOR U676 ( .A(n311), .B(n310), .Z(n312) );
  XNOR U677 ( .A(in[1237]), .B(n312), .Z(n756) );
  XOR U678 ( .A(n1040), .B(n756), .Z(n4250) );
  XOR U679 ( .A(in[982]), .B(n4250), .Z(n1913) );
  NANDN U680 ( .A(n1916), .B(n1913), .Z(n313) );
  XNOR U681 ( .A(n1511), .B(n313), .Z(out[1002]) );
  XOR U682 ( .A(in[1389]), .B(in[109]), .Z(n315) );
  XNOR U683 ( .A(in[1069]), .B(in[749]), .Z(n314) );
  XNOR U684 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U685 ( .A(in[429]), .B(n316), .Z(n1602) );
  XOR U686 ( .A(in[1518]), .B(in[558]), .Z(n318) );
  XNOR U687 ( .A(in[878]), .B(in[238]), .Z(n317) );
  XNOR U688 ( .A(n318), .B(n317), .Z(n319) );
  XNOR U689 ( .A(in[1198]), .B(n319), .Z(n1542) );
  XOR U690 ( .A(n1602), .B(n1542), .Z(n1413) );
  XOR U691 ( .A(in[174]), .B(n1413), .Z(n1515) );
  XOR U692 ( .A(in[143]), .B(in[1423]), .Z(n321) );
  XNOR U693 ( .A(in[1103]), .B(in[783]), .Z(n320) );
  XNOR U694 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U695 ( .A(in[463]), .B(n322), .Z(n1402) );
  XOR U696 ( .A(in[974]), .B(in[14]), .Z(n324) );
  XNOR U697 ( .A(in[1294]), .B(in[334]), .Z(n323) );
  XNOR U698 ( .A(n324), .B(n323), .Z(n325) );
  XOR U699 ( .A(in[654]), .B(n325), .Z(n1437) );
  XNOR U700 ( .A(in[1359]), .B(n4467), .Z(n1920) );
  XOR U701 ( .A(in[1367]), .B(in[727]), .Z(n327) );
  XNOR U702 ( .A(in[87]), .B(in[407]), .Z(n326) );
  XNOR U703 ( .A(n327), .B(n326), .Z(n328) );
  XNOR U704 ( .A(in[1047]), .B(n328), .Z(n1053) );
  XOR U705 ( .A(in[1558]), .B(in[598]), .Z(n330) );
  XNOR U706 ( .A(in[918]), .B(in[278]), .Z(n329) );
  XNOR U707 ( .A(n330), .B(n329), .Z(n331) );
  XNOR U708 ( .A(in[1238]), .B(n331), .Z(n771) );
  XOR U709 ( .A(n1053), .B(n771), .Z(n4251) );
  XOR U710 ( .A(in[983]), .B(n4251), .Z(n1917) );
  NANDN U711 ( .A(n1920), .B(n1917), .Z(n332) );
  XNOR U712 ( .A(n1515), .B(n332), .Z(out[1003]) );
  XOR U713 ( .A(in[1390]), .B(in[110]), .Z(n334) );
  XNOR U714 ( .A(in[1070]), .B(in[750]), .Z(n333) );
  XNOR U715 ( .A(n334), .B(n333), .Z(n335) );
  XNOR U716 ( .A(in[430]), .B(n335), .Z(n1606) );
  XOR U717 ( .A(in[1519]), .B(in[559]), .Z(n337) );
  XNOR U718 ( .A(in[879]), .B(in[239]), .Z(n336) );
  XNOR U719 ( .A(n337), .B(n336), .Z(n338) );
  XNOR U720 ( .A(in[1199]), .B(n338), .Z(n1546) );
  XOR U721 ( .A(n1606), .B(n1546), .Z(n1425) );
  XOR U722 ( .A(in[175]), .B(n1425), .Z(n1519) );
  XOR U723 ( .A(in[144]), .B(in[1424]), .Z(n340) );
  XNOR U724 ( .A(in[1104]), .B(in[784]), .Z(n339) );
  XNOR U725 ( .A(n340), .B(n339), .Z(n341) );
  XNOR U726 ( .A(in[464]), .B(n341), .Z(n1406) );
  XOR U727 ( .A(in[975]), .B(in[15]), .Z(n343) );
  XNOR U728 ( .A(in[1295]), .B(in[335]), .Z(n342) );
  XNOR U729 ( .A(n343), .B(n342), .Z(n344) );
  XOR U730 ( .A(in[655]), .B(n344), .Z(n1438) );
  XNOR U731 ( .A(in[1360]), .B(n4470), .Z(n1926) );
  XOR U732 ( .A(in[1368]), .B(in[728]), .Z(n346) );
  XNOR U733 ( .A(in[88]), .B(in[408]), .Z(n345) );
  XNOR U734 ( .A(n346), .B(n345), .Z(n347) );
  XNOR U735 ( .A(in[1048]), .B(n347), .Z(n1066) );
  XOR U736 ( .A(in[1559]), .B(in[599]), .Z(n349) );
  XNOR U737 ( .A(in[919]), .B(in[279]), .Z(n348) );
  XNOR U738 ( .A(n349), .B(n348), .Z(n350) );
  XNOR U739 ( .A(in[1239]), .B(n350), .Z(n786) );
  XOR U740 ( .A(n1066), .B(n786), .Z(n4252) );
  XOR U741 ( .A(in[984]), .B(n4252), .Z(n1923) );
  NANDN U742 ( .A(n1926), .B(n1923), .Z(n351) );
  XNOR U743 ( .A(n1519), .B(n351), .Z(out[1004]) );
  XOR U744 ( .A(in[1391]), .B(in[111]), .Z(n353) );
  XNOR U745 ( .A(in[1071]), .B(in[751]), .Z(n352) );
  XNOR U746 ( .A(n353), .B(n352), .Z(n354) );
  XNOR U747 ( .A(in[431]), .B(n354), .Z(n1610) );
  XOR U748 ( .A(in[1520]), .B(in[560]), .Z(n356) );
  XNOR U749 ( .A(in[880]), .B(in[240]), .Z(n355) );
  XNOR U750 ( .A(n356), .B(n355), .Z(n357) );
  XNOR U751 ( .A(in[1200]), .B(n357), .Z(n1552) );
  XOR U752 ( .A(n1610), .B(n1552), .Z(n1444) );
  XOR U753 ( .A(in[176]), .B(n1444), .Z(n1523) );
  XOR U754 ( .A(in[145]), .B(in[1425]), .Z(n359) );
  XNOR U755 ( .A(in[1105]), .B(in[785]), .Z(n358) );
  XNOR U756 ( .A(n359), .B(n358), .Z(n360) );
  XNOR U757 ( .A(in[465]), .B(n360), .Z(n1410) );
  XOR U758 ( .A(in[976]), .B(in[16]), .Z(n362) );
  XNOR U759 ( .A(in[1296]), .B(in[336]), .Z(n361) );
  XNOR U760 ( .A(n362), .B(n361), .Z(n363) );
  XOR U761 ( .A(in[656]), .B(n363), .Z(n1439) );
  XNOR U762 ( .A(in[1361]), .B(n4477), .Z(n1930) );
  XOR U763 ( .A(in[1369]), .B(in[729]), .Z(n365) );
  XNOR U764 ( .A(in[89]), .B(in[409]), .Z(n364) );
  XNOR U765 ( .A(n365), .B(n364), .Z(n366) );
  XNOR U766 ( .A(in[1049]), .B(n366), .Z(n1079) );
  XOR U767 ( .A(in[1560]), .B(in[600]), .Z(n368) );
  XNOR U768 ( .A(in[920]), .B(in[280]), .Z(n367) );
  XNOR U769 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U770 ( .A(in[1240]), .B(n369), .Z(n801) );
  XOR U771 ( .A(n1079), .B(n801), .Z(n4253) );
  XOR U772 ( .A(in[985]), .B(n4253), .Z(n1927) );
  NANDN U773 ( .A(n1930), .B(n1927), .Z(n370) );
  XNOR U774 ( .A(n1523), .B(n370), .Z(out[1005]) );
  XOR U775 ( .A(in[1392]), .B(in[112]), .Z(n372) );
  XNOR U776 ( .A(in[1072]), .B(in[752]), .Z(n371) );
  XNOR U777 ( .A(n372), .B(n371), .Z(n373) );
  XNOR U778 ( .A(in[432]), .B(n373), .Z(n1614) );
  XOR U779 ( .A(in[1521]), .B(in[561]), .Z(n375) );
  XNOR U780 ( .A(in[881]), .B(in[241]), .Z(n374) );
  XNOR U781 ( .A(n375), .B(n374), .Z(n376) );
  XNOR U782 ( .A(in[1201]), .B(n376), .Z(n1556) );
  XOR U783 ( .A(n1614), .B(n1556), .Z(n1472) );
  XOR U784 ( .A(in[177]), .B(n1472), .Z(n1527) );
  XOR U785 ( .A(in[17]), .B(in[657]), .Z(n378) );
  XNOR U786 ( .A(in[977]), .B(in[337]), .Z(n377) );
  XNOR U787 ( .A(n378), .B(n377), .Z(n379) );
  XNOR U788 ( .A(in[1297]), .B(n379), .Z(n1441) );
  XOR U789 ( .A(in[1426]), .B(in[466]), .Z(n381) );
  XNOR U790 ( .A(in[786]), .B(in[146]), .Z(n380) );
  XNOR U791 ( .A(n381), .B(n380), .Z(n382) );
  XOR U792 ( .A(in[1106]), .B(n382), .Z(n725) );
  XNOR U793 ( .A(n4480), .B(in[1362]), .Z(n1934) );
  XOR U794 ( .A(in[1370]), .B(in[730]), .Z(n384) );
  XNOR U795 ( .A(in[90]), .B(in[410]), .Z(n383) );
  XNOR U796 ( .A(n384), .B(n383), .Z(n385) );
  XNOR U797 ( .A(in[1050]), .B(n385), .Z(n1094) );
  XOR U798 ( .A(in[1561]), .B(in[601]), .Z(n387) );
  XNOR U799 ( .A(in[921]), .B(in[281]), .Z(n386) );
  XNOR U800 ( .A(n387), .B(n386), .Z(n388) );
  XNOR U801 ( .A(in[1241]), .B(n388), .Z(n827) );
  XOR U802 ( .A(n1094), .B(n827), .Z(n4254) );
  XOR U803 ( .A(in[986]), .B(n4254), .Z(n1931) );
  NANDN U804 ( .A(n1934), .B(n1931), .Z(n389) );
  XNOR U805 ( .A(n1527), .B(n389), .Z(out[1006]) );
  XOR U806 ( .A(in[1393]), .B(in[113]), .Z(n391) );
  XNOR U807 ( .A(in[1073]), .B(in[753]), .Z(n390) );
  XNOR U808 ( .A(n391), .B(n390), .Z(n392) );
  XNOR U809 ( .A(in[433]), .B(n392), .Z(n1618) );
  XOR U810 ( .A(in[1522]), .B(in[562]), .Z(n394) );
  XNOR U811 ( .A(in[882]), .B(in[242]), .Z(n393) );
  XNOR U812 ( .A(n394), .B(n393), .Z(n395) );
  XNOR U813 ( .A(in[1202]), .B(n395), .Z(n1560) );
  XOR U814 ( .A(n1618), .B(n1560), .Z(n1507) );
  XOR U815 ( .A(in[178]), .B(n1507), .Z(n1531) );
  XOR U816 ( .A(in[978]), .B(in[18]), .Z(n397) );
  XNOR U817 ( .A(in[1298]), .B(in[338]), .Z(n396) );
  XNOR U818 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U819 ( .A(in[658]), .B(n398), .Z(n1443) );
  XOR U820 ( .A(in[147]), .B(in[1427]), .Z(n400) );
  XNOR U821 ( .A(in[1107]), .B(in[787]), .Z(n399) );
  XNOR U822 ( .A(n400), .B(n399), .Z(n401) );
  XOR U823 ( .A(in[467]), .B(n401), .Z(n740) );
  XNOR U824 ( .A(in[1363]), .B(n4483), .Z(n1938) );
  XOR U825 ( .A(in[1371]), .B(in[731]), .Z(n403) );
  XNOR U826 ( .A(in[91]), .B(in[411]), .Z(n402) );
  XNOR U827 ( .A(n403), .B(n402), .Z(n404) );
  XNOR U828 ( .A(in[1051]), .B(n404), .Z(n1107) );
  XOR U829 ( .A(in[1562]), .B(in[602]), .Z(n406) );
  XNOR U830 ( .A(in[922]), .B(in[282]), .Z(n405) );
  XNOR U831 ( .A(n406), .B(n405), .Z(n407) );
  XNOR U832 ( .A(in[1242]), .B(n407), .Z(n842) );
  XOR U833 ( .A(n1107), .B(n842), .Z(n4255) );
  XOR U834 ( .A(in[987]), .B(n4255), .Z(n1935) );
  NANDN U835 ( .A(n1938), .B(n1935), .Z(n408) );
  XNOR U836 ( .A(n1531), .B(n408), .Z(out[1007]) );
  XOR U837 ( .A(in[1394]), .B(in[114]), .Z(n410) );
  XNOR U838 ( .A(in[1074]), .B(in[754]), .Z(n409) );
  XNOR U839 ( .A(n410), .B(n409), .Z(n411) );
  XNOR U840 ( .A(in[434]), .B(n411), .Z(n1622) );
  XOR U841 ( .A(in[1523]), .B(in[563]), .Z(n413) );
  XNOR U842 ( .A(in[883]), .B(in[243]), .Z(n412) );
  XNOR U843 ( .A(n413), .B(n412), .Z(n414) );
  XNOR U844 ( .A(in[1203]), .B(n414), .Z(n1564) );
  XOR U845 ( .A(n1622), .B(n1564), .Z(n1549) );
  XOR U846 ( .A(in[179]), .B(n1549), .Z(n1535) );
  XOR U847 ( .A(in[148]), .B(in[1428]), .Z(n416) );
  XNOR U848 ( .A(in[1108]), .B(in[788]), .Z(n415) );
  XNOR U849 ( .A(n416), .B(n415), .Z(n417) );
  XNOR U850 ( .A(in[468]), .B(n417), .Z(n755) );
  XOR U851 ( .A(in[979]), .B(in[19]), .Z(n419) );
  XNOR U852 ( .A(in[1299]), .B(in[339]), .Z(n418) );
  XNOR U853 ( .A(n419), .B(n418), .Z(n420) );
  XOR U854 ( .A(in[659]), .B(n420), .Z(n1447) );
  XNOR U855 ( .A(in[1364]), .B(n4486), .Z(n1942) );
  XOR U856 ( .A(in[1372]), .B(in[732]), .Z(n422) );
  XNOR U857 ( .A(in[92]), .B(in[412]), .Z(n421) );
  XNOR U858 ( .A(n422), .B(n421), .Z(n423) );
  XNOR U859 ( .A(in[1052]), .B(n423), .Z(n1127) );
  XOR U860 ( .A(in[1563]), .B(in[603]), .Z(n425) );
  XNOR U861 ( .A(in[923]), .B(in[283]), .Z(n424) );
  XNOR U862 ( .A(n425), .B(n424), .Z(n426) );
  XNOR U863 ( .A(in[1243]), .B(n426), .Z(n857) );
  XOR U864 ( .A(n1127), .B(n857), .Z(n4258) );
  XOR U865 ( .A(in[988]), .B(n4258), .Z(n1939) );
  NANDN U866 ( .A(n1942), .B(n1939), .Z(n427) );
  XNOR U867 ( .A(n1535), .B(n427), .Z(out[1008]) );
  XOR U868 ( .A(in[1395]), .B(in[115]), .Z(n429) );
  XNOR U869 ( .A(in[1075]), .B(in[755]), .Z(n428) );
  XNOR U870 ( .A(n429), .B(n428), .Z(n430) );
  XNOR U871 ( .A(in[435]), .B(n430), .Z(n1626) );
  XOR U872 ( .A(in[1524]), .B(in[564]), .Z(n432) );
  XNOR U873 ( .A(in[884]), .B(in[244]), .Z(n431) );
  XNOR U874 ( .A(n432), .B(n431), .Z(n433) );
  XNOR U875 ( .A(in[1204]), .B(n433), .Z(n1568) );
  XOR U876 ( .A(n1626), .B(n1568), .Z(n1591) );
  XOR U877 ( .A(in[180]), .B(n1591), .Z(n1539) );
  XOR U878 ( .A(in[340]), .B(in[660]), .Z(n435) );
  XNOR U879 ( .A(in[20]), .B(in[1300]), .Z(n434) );
  XNOR U880 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U881 ( .A(in[980]), .B(n436), .Z(n1449) );
  XOR U882 ( .A(in[149]), .B(in[1429]), .Z(n438) );
  XNOR U883 ( .A(in[1109]), .B(in[789]), .Z(n437) );
  XNOR U884 ( .A(n438), .B(n437), .Z(n439) );
  XOR U885 ( .A(in[469]), .B(n439), .Z(n770) );
  XNOR U886 ( .A(in[1365]), .B(n4489), .Z(n1946) );
  XOR U887 ( .A(in[1373]), .B(in[733]), .Z(n441) );
  XNOR U888 ( .A(in[93]), .B(in[413]), .Z(n440) );
  XNOR U889 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U890 ( .A(in[1053]), .B(n442), .Z(n1140) );
  XOR U891 ( .A(in[1564]), .B(in[604]), .Z(n444) );
  XNOR U892 ( .A(in[924]), .B(in[284]), .Z(n443) );
  XNOR U893 ( .A(n444), .B(n443), .Z(n445) );
  XNOR U894 ( .A(in[1244]), .B(n445), .Z(n872) );
  XOR U895 ( .A(n1140), .B(n872), .Z(n4259) );
  XOR U896 ( .A(in[989]), .B(n4259), .Z(n1943) );
  NANDN U897 ( .A(n1946), .B(n1943), .Z(n446) );
  XNOR U898 ( .A(n1539), .B(n446), .Z(out[1009]) );
  XOR U899 ( .A(in[1339]), .B(in[59]), .Z(n448) );
  XNOR U900 ( .A(in[699]), .B(in[379]), .Z(n447) );
  XNOR U901 ( .A(n448), .B(n447), .Z(n449) );
  XNOR U902 ( .A(in[1019]), .B(n449), .Z(n1098) );
  XOR U903 ( .A(in[1530]), .B(in[570]), .Z(n451) );
  XNOR U904 ( .A(in[1210]), .B(in[250]), .Z(n450) );
  XNOR U905 ( .A(n451), .B(n450), .Z(n452) );
  XNOR U906 ( .A(in[890]), .B(n452), .Z(n564) );
  XOR U907 ( .A(n1098), .B(n564), .Z(n3953) );
  XOR U908 ( .A(in[635]), .B(n3953), .Z(n2707) );
  IV U909 ( .A(n2707), .Z(n2793) );
  XOR U910 ( .A(in[161]), .B(in[1441]), .Z(n454) );
  XNOR U911 ( .A(in[801]), .B(in[1121]), .Z(n453) );
  XNOR U912 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U913 ( .A(in[481]), .B(n455), .Z(n691) );
  XOR U914 ( .A(in[1570]), .B(in[610]), .Z(n457) );
  XNOR U915 ( .A(in[930]), .B(in[290]), .Z(n456) );
  XNOR U916 ( .A(n457), .B(n456), .Z(n458) );
  XOR U917 ( .A(in[1250]), .B(n458), .Z(n574) );
  XOR U918 ( .A(in[226]), .B(n4049), .Z(n3117) );
  XOR U919 ( .A(in[1510]), .B(in[550]), .Z(n460) );
  XNOR U920 ( .A(in[870]), .B(in[230]), .Z(n459) );
  XNOR U921 ( .A(n460), .B(n459), .Z(n461) );
  XNOR U922 ( .A(in[1190]), .B(n461), .Z(n1510) );
  XOR U923 ( .A(in[1061]), .B(in[421]), .Z(n463) );
  XNOR U924 ( .A(in[741]), .B(in[1381]), .Z(n462) );
  XNOR U925 ( .A(n463), .B(n462), .Z(n464) );
  XNOR U926 ( .A(in[101]), .B(n464), .Z(n610) );
  XNOR U927 ( .A(n1510), .B(n610), .Z(n4089) );
  IV U928 ( .A(n4089), .Z(n1253) );
  XOR U929 ( .A(in[1446]), .B(n1253), .Z(n3114) );
  NANDN U930 ( .A(n3117), .B(n3114), .Z(n465) );
  XOR U931 ( .A(n2793), .B(n465), .Z(out[100]) );
  XOR U932 ( .A(in[1396]), .B(in[116]), .Z(n467) );
  XNOR U933 ( .A(in[1076]), .B(in[756]), .Z(n466) );
  XNOR U934 ( .A(n467), .B(n466), .Z(n468) );
  XNOR U935 ( .A(in[436]), .B(n468), .Z(n1631) );
  XOR U936 ( .A(in[1525]), .B(in[565]), .Z(n470) );
  XNOR U937 ( .A(in[885]), .B(in[245]), .Z(n469) );
  XNOR U938 ( .A(n470), .B(n469), .Z(n471) );
  XNOR U939 ( .A(in[1205]), .B(n471), .Z(n1572) );
  XOR U940 ( .A(n1631), .B(n1572), .Z(n4153) );
  XOR U941 ( .A(in[181]), .B(n4153), .Z(n1543) );
  XOR U942 ( .A(in[341]), .B(in[661]), .Z(n473) );
  XNOR U943 ( .A(in[21]), .B(in[1301]), .Z(n472) );
  XNOR U944 ( .A(n473), .B(n472), .Z(n474) );
  XNOR U945 ( .A(in[981]), .B(n474), .Z(n1451) );
  XOR U946 ( .A(in[150]), .B(in[1430]), .Z(n476) );
  XNOR U947 ( .A(in[1110]), .B(in[790]), .Z(n475) );
  XNOR U948 ( .A(n476), .B(n475), .Z(n477) );
  XOR U949 ( .A(in[470]), .B(n477), .Z(n785) );
  XNOR U950 ( .A(in[1366]), .B(n4492), .Z(n1950) );
  XOR U951 ( .A(in[1374]), .B(in[734]), .Z(n479) );
  XNOR U952 ( .A(in[94]), .B(in[414]), .Z(n478) );
  XNOR U953 ( .A(n479), .B(n478), .Z(n480) );
  XNOR U954 ( .A(in[1054]), .B(n480), .Z(n1153) );
  XOR U955 ( .A(in[1565]), .B(in[605]), .Z(n482) );
  XNOR U956 ( .A(in[925]), .B(in[285]), .Z(n481) );
  XNOR U957 ( .A(n482), .B(n481), .Z(n483) );
  XNOR U958 ( .A(in[1245]), .B(n483), .Z(n887) );
  XOR U959 ( .A(n1153), .B(n887), .Z(n4260) );
  XOR U960 ( .A(in[990]), .B(n4260), .Z(n1947) );
  NANDN U961 ( .A(n1950), .B(n1947), .Z(n484) );
  XNOR U962 ( .A(n1543), .B(n484), .Z(out[1010]) );
  XOR U963 ( .A(in[1526]), .B(in[566]), .Z(n486) );
  XNOR U964 ( .A(in[886]), .B(in[246]), .Z(n485) );
  XNOR U965 ( .A(n486), .B(n485), .Z(n487) );
  XNOR U966 ( .A(in[1206]), .B(n487), .Z(n1576) );
  XOR U967 ( .A(in[1397]), .B(in[117]), .Z(n489) );
  XNOR U968 ( .A(in[1077]), .B(in[757]), .Z(n488) );
  XNOR U969 ( .A(n489), .B(n488), .Z(n490) );
  XNOR U970 ( .A(in[437]), .B(n490), .Z(n1635) );
  XOR U971 ( .A(n1576), .B(n1635), .Z(n4163) );
  XOR U972 ( .A(in[182]), .B(n4163), .Z(n1547) );
  XOR U973 ( .A(in[151]), .B(in[1431]), .Z(n492) );
  XNOR U974 ( .A(in[1111]), .B(in[791]), .Z(n491) );
  XNOR U975 ( .A(n492), .B(n491), .Z(n493) );
  XNOR U976 ( .A(in[471]), .B(n493), .Z(n800) );
  XOR U977 ( .A(in[342]), .B(in[662]), .Z(n495) );
  XNOR U978 ( .A(in[22]), .B(in[1302]), .Z(n494) );
  XNOR U979 ( .A(n495), .B(n494), .Z(n496) );
  XOR U980 ( .A(in[982]), .B(n496), .Z(n1453) );
  XNOR U981 ( .A(in[1367]), .B(n4495), .Z(n1954) );
  XOR U982 ( .A(in[1375]), .B(in[735]), .Z(n498) );
  XNOR U983 ( .A(in[95]), .B(in[415]), .Z(n497) );
  XNOR U984 ( .A(n498), .B(n497), .Z(n499) );
  XNOR U985 ( .A(in[1055]), .B(n499), .Z(n1166) );
  XOR U986 ( .A(in[1566]), .B(in[606]), .Z(n501) );
  XNOR U987 ( .A(in[926]), .B(in[286]), .Z(n500) );
  XNOR U988 ( .A(n501), .B(n500), .Z(n502) );
  XNOR U989 ( .A(in[1246]), .B(n502), .Z(n902) );
  XOR U990 ( .A(n1166), .B(n902), .Z(n4261) );
  XOR U991 ( .A(in[991]), .B(n4261), .Z(n1951) );
  NANDN U992 ( .A(n1954), .B(n1951), .Z(n503) );
  XNOR U993 ( .A(n1547), .B(n503), .Z(out[1011]) );
  XOR U994 ( .A(in[1527]), .B(in[567]), .Z(n505) );
  XNOR U995 ( .A(in[887]), .B(in[247]), .Z(n504) );
  XNOR U996 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U997 ( .A(in[1207]), .B(n506), .Z(n1580) );
  XOR U998 ( .A(in[1398]), .B(in[118]), .Z(n508) );
  XNOR U999 ( .A(in[1078]), .B(in[758]), .Z(n507) );
  XNOR U1000 ( .A(n508), .B(n507), .Z(n509) );
  XNOR U1001 ( .A(in[438]), .B(n509), .Z(n1639) );
  XOR U1002 ( .A(n1580), .B(n1639), .Z(n4167) );
  XOR U1003 ( .A(in[183]), .B(n4167), .Z(n1553) );
  XOR U1004 ( .A(in[152]), .B(in[1432]), .Z(n511) );
  XNOR U1005 ( .A(in[1112]), .B(in[792]), .Z(n510) );
  XNOR U1006 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U1007 ( .A(in[472]), .B(n512), .Z(n826) );
  XOR U1008 ( .A(in[343]), .B(in[663]), .Z(n514) );
  XNOR U1009 ( .A(in[23]), .B(in[1303]), .Z(n513) );
  XNOR U1010 ( .A(n514), .B(n513), .Z(n515) );
  XOR U1011 ( .A(in[983]), .B(n515), .Z(n1455) );
  XNOR U1012 ( .A(in[1368]), .B(n4498), .Z(n1958) );
  XOR U1013 ( .A(in[1376]), .B(in[736]), .Z(n517) );
  XNOR U1014 ( .A(in[96]), .B(in[416]), .Z(n516) );
  XNOR U1015 ( .A(n517), .B(n516), .Z(n518) );
  XNOR U1016 ( .A(in[1056]), .B(n518), .Z(n1181) );
  XOR U1017 ( .A(in[1567]), .B(in[607]), .Z(n520) );
  XNOR U1018 ( .A(in[927]), .B(in[287]), .Z(n519) );
  XNOR U1019 ( .A(n520), .B(n519), .Z(n521) );
  XNOR U1020 ( .A(in[1247]), .B(n521), .Z(n917) );
  XOR U1021 ( .A(n1181), .B(n917), .Z(n4264) );
  XOR U1022 ( .A(in[992]), .B(n4264), .Z(n1955) );
  NANDN U1023 ( .A(n1958), .B(n1955), .Z(n522) );
  XNOR U1024 ( .A(n1553), .B(n522), .Z(out[1012]) );
  XOR U1025 ( .A(in[1528]), .B(in[568]), .Z(n524) );
  XNOR U1026 ( .A(in[888]), .B(in[248]), .Z(n523) );
  XNOR U1027 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U1028 ( .A(in[1208]), .B(n525), .Z(n1584) );
  XOR U1029 ( .A(in[1399]), .B(in[119]), .Z(n527) );
  XNOR U1030 ( .A(in[1079]), .B(in[759]), .Z(n526) );
  XNOR U1031 ( .A(n527), .B(n526), .Z(n528) );
  XNOR U1032 ( .A(in[439]), .B(n528), .Z(n1643) );
  XOR U1033 ( .A(n1584), .B(n1643), .Z(n4171) );
  XOR U1034 ( .A(in[184]), .B(n4171), .Z(n1557) );
  XOR U1035 ( .A(in[344]), .B(in[664]), .Z(n530) );
  XNOR U1036 ( .A(in[24]), .B(in[1304]), .Z(n529) );
  XNOR U1037 ( .A(n530), .B(n529), .Z(n531) );
  XNOR U1038 ( .A(in[984]), .B(n531), .Z(n1457) );
  XOR U1039 ( .A(in[153]), .B(in[1433]), .Z(n533) );
  XNOR U1040 ( .A(in[1113]), .B(in[793]), .Z(n532) );
  XNOR U1041 ( .A(n533), .B(n532), .Z(n534) );
  XOR U1042 ( .A(in[473]), .B(n534), .Z(n841) );
  XNOR U1043 ( .A(in[1369]), .B(n4501), .Z(n1962) );
  XOR U1044 ( .A(in[1377]), .B(in[737]), .Z(n536) );
  XNOR U1045 ( .A(in[97]), .B(in[417]), .Z(n535) );
  XNOR U1046 ( .A(n536), .B(n535), .Z(n537) );
  XNOR U1047 ( .A(in[1057]), .B(n537), .Z(n1196) );
  XOR U1048 ( .A(in[1568]), .B(in[608]), .Z(n539) );
  XNOR U1049 ( .A(in[928]), .B(in[288]), .Z(n538) );
  XNOR U1050 ( .A(n539), .B(n538), .Z(n540) );
  XNOR U1051 ( .A(in[1248]), .B(n540), .Z(n932) );
  XOR U1052 ( .A(n1196), .B(n932), .Z(n4267) );
  XOR U1053 ( .A(in[993]), .B(n4267), .Z(n1959) );
  NANDN U1054 ( .A(n1962), .B(n1959), .Z(n541) );
  XNOR U1055 ( .A(n1557), .B(n541), .Z(out[1013]) );
  XOR U1056 ( .A(in[1529]), .B(in[569]), .Z(n543) );
  XNOR U1057 ( .A(in[889]), .B(in[249]), .Z(n542) );
  XNOR U1058 ( .A(n543), .B(n542), .Z(n544) );
  XNOR U1059 ( .A(in[1209]), .B(n544), .Z(n1588) );
  XOR U1060 ( .A(in[1400]), .B(in[120]), .Z(n546) );
  XNOR U1061 ( .A(in[1080]), .B(in[760]), .Z(n545) );
  XNOR U1062 ( .A(n546), .B(n545), .Z(n547) );
  XNOR U1063 ( .A(in[440]), .B(n547), .Z(n1647) );
  XOR U1064 ( .A(n1588), .B(n1647), .Z(n4175) );
  XOR U1065 ( .A(in[185]), .B(n4175), .Z(n1561) );
  XOR U1066 ( .A(in[345]), .B(in[665]), .Z(n549) );
  XNOR U1067 ( .A(in[25]), .B(in[1305]), .Z(n548) );
  XNOR U1068 ( .A(n549), .B(n548), .Z(n550) );
  XNOR U1069 ( .A(in[985]), .B(n550), .Z(n1461) );
  XOR U1070 ( .A(in[154]), .B(in[1434]), .Z(n552) );
  XNOR U1071 ( .A(in[1114]), .B(in[794]), .Z(n551) );
  XNOR U1072 ( .A(n552), .B(n551), .Z(n553) );
  XOR U1073 ( .A(in[474]), .B(n553), .Z(n856) );
  XNOR U1074 ( .A(in[1370]), .B(n4504), .Z(n1968) );
  XOR U1075 ( .A(in[1569]), .B(in[609]), .Z(n555) );
  XNOR U1076 ( .A(in[929]), .B(in[289]), .Z(n554) );
  XNOR U1077 ( .A(n555), .B(n554), .Z(n556) );
  XNOR U1078 ( .A(in[1249]), .B(n556), .Z(n947) );
  XOR U1079 ( .A(in[1378]), .B(in[738]), .Z(n558) );
  XNOR U1080 ( .A(in[98]), .B(in[418]), .Z(n557) );
  XNOR U1081 ( .A(n558), .B(n557), .Z(n559) );
  XNOR U1082 ( .A(in[1058]), .B(n559), .Z(n1211) );
  XOR U1083 ( .A(n947), .B(n1211), .Z(n4270) );
  XOR U1084 ( .A(in[994]), .B(n4270), .Z(n1965) );
  NANDN U1085 ( .A(n1968), .B(n1965), .Z(n560) );
  XNOR U1086 ( .A(n1561), .B(n560), .Z(out[1014]) );
  XOR U1087 ( .A(in[1401]), .B(in[121]), .Z(n562) );
  XNOR U1088 ( .A(in[1081]), .B(in[761]), .Z(n561) );
  XNOR U1089 ( .A(n562), .B(n561), .Z(n563) );
  XNOR U1090 ( .A(in[441]), .B(n563), .Z(n1651) );
  XOR U1091 ( .A(n564), .B(n1651), .Z(n1798) );
  XOR U1092 ( .A(in[186]), .B(n1798), .Z(n1565) );
  XOR U1093 ( .A(in[155]), .B(in[1435]), .Z(n566) );
  XNOR U1094 ( .A(in[1115]), .B(in[795]), .Z(n565) );
  XNOR U1095 ( .A(n566), .B(n565), .Z(n567) );
  XNOR U1096 ( .A(in[475]), .B(n567), .Z(n871) );
  XOR U1097 ( .A(in[346]), .B(in[666]), .Z(n569) );
  XNOR U1098 ( .A(in[26]), .B(in[1306]), .Z(n568) );
  XNOR U1099 ( .A(n569), .B(n568), .Z(n570) );
  XOR U1100 ( .A(in[986]), .B(n570), .Z(n1463) );
  IV U1101 ( .A(n4511), .Z(n2743) );
  XOR U1102 ( .A(in[1371]), .B(n2743), .Z(n1369) );
  IV U1103 ( .A(n1369), .Z(n1972) );
  XOR U1104 ( .A(in[1379]), .B(in[739]), .Z(n572) );
  XNOR U1105 ( .A(in[99]), .B(in[419]), .Z(n571) );
  XNOR U1106 ( .A(n572), .B(n571), .Z(n573) );
  XOR U1107 ( .A(in[1059]), .B(n573), .Z(n1226) );
  XNOR U1108 ( .A(n574), .B(n1226), .Z(n4273) );
  XNOR U1109 ( .A(in[995]), .B(n4273), .Z(n1969) );
  NANDN U1110 ( .A(n1972), .B(n1969), .Z(n575) );
  XNOR U1111 ( .A(n1565), .B(n575), .Z(out[1015]) );
  XOR U1112 ( .A(in[1402]), .B(in[122]), .Z(n577) );
  XNOR U1113 ( .A(in[1082]), .B(in[762]), .Z(n576) );
  XNOR U1114 ( .A(n577), .B(n576), .Z(n578) );
  XNOR U1115 ( .A(in[442]), .B(n578), .Z(n1655) );
  XOR U1116 ( .A(in[1531]), .B(in[571]), .Z(n580) );
  XNOR U1117 ( .A(in[1211]), .B(in[251]), .Z(n579) );
  XNOR U1118 ( .A(n580), .B(n579), .Z(n581) );
  XNOR U1119 ( .A(in[891]), .B(n581), .Z(n653) );
  XOR U1120 ( .A(n1655), .B(n653), .Z(n1824) );
  XOR U1121 ( .A(in[187]), .B(n1824), .Z(n1569) );
  XOR U1122 ( .A(in[156]), .B(in[1436]), .Z(n583) );
  XNOR U1123 ( .A(in[1116]), .B(in[796]), .Z(n582) );
  XNOR U1124 ( .A(n583), .B(n582), .Z(n584) );
  XNOR U1125 ( .A(in[476]), .B(n584), .Z(n886) );
  XOR U1126 ( .A(in[347]), .B(in[667]), .Z(n586) );
  XNOR U1127 ( .A(in[27]), .B(in[1307]), .Z(n585) );
  XNOR U1128 ( .A(n586), .B(n585), .Z(n587) );
  XOR U1129 ( .A(in[987]), .B(n587), .Z(n1465) );
  IV U1130 ( .A(n4514), .Z(n2760) );
  XOR U1131 ( .A(in[1372]), .B(n2760), .Z(n1379) );
  IV U1132 ( .A(n1379), .Z(n1976) );
  XOR U1133 ( .A(in[1060]), .B(in[420]), .Z(n589) );
  XNOR U1134 ( .A(in[740]), .B(in[1380]), .Z(n588) );
  XNOR U1135 ( .A(n589), .B(n588), .Z(n590) );
  XNOR U1136 ( .A(in[100]), .B(n590), .Z(n1241) );
  XOR U1137 ( .A(in[1571]), .B(in[611]), .Z(n592) );
  XNOR U1138 ( .A(in[931]), .B(in[291]), .Z(n591) );
  XNOR U1139 ( .A(n592), .B(n591), .Z(n593) );
  XNOR U1140 ( .A(in[1251]), .B(n593), .Z(n657) );
  XOR U1141 ( .A(n1241), .B(n657), .Z(n4276) );
  XOR U1142 ( .A(in[996]), .B(n4276), .Z(n1973) );
  NANDN U1143 ( .A(n1976), .B(n1973), .Z(n594) );
  XNOR U1144 ( .A(n1569), .B(n594), .Z(out[1016]) );
  XOR U1145 ( .A(in[1403]), .B(in[123]), .Z(n596) );
  XNOR U1146 ( .A(in[1083]), .B(in[763]), .Z(n595) );
  XNOR U1147 ( .A(n596), .B(n595), .Z(n597) );
  XNOR U1148 ( .A(in[443]), .B(n597), .Z(n1659) );
  XOR U1149 ( .A(in[1532]), .B(in[572]), .Z(n599) );
  XNOR U1150 ( .A(in[1212]), .B(in[252]), .Z(n598) );
  XNOR U1151 ( .A(n599), .B(n598), .Z(n600) );
  XNOR U1152 ( .A(in[892]), .B(n600), .Z(n818) );
  XOR U1153 ( .A(n1659), .B(n818), .Z(n1847) );
  XOR U1154 ( .A(in[188]), .B(n1847), .Z(n1573) );
  XOR U1155 ( .A(in[157]), .B(in[1437]), .Z(n602) );
  XNOR U1156 ( .A(in[1117]), .B(in[797]), .Z(n601) );
  XNOR U1157 ( .A(n602), .B(n601), .Z(n603) );
  XNOR U1158 ( .A(in[477]), .B(n603), .Z(n901) );
  XOR U1159 ( .A(in[348]), .B(in[668]), .Z(n605) );
  XNOR U1160 ( .A(in[28]), .B(in[1308]), .Z(n604) );
  XNOR U1161 ( .A(n605), .B(n604), .Z(n606) );
  XOR U1162 ( .A(in[988]), .B(n606), .Z(n1469) );
  IV U1163 ( .A(n4517), .Z(n2777) );
  XOR U1164 ( .A(in[1373]), .B(n2777), .Z(n1385) );
  IV U1165 ( .A(n1385), .Z(n1980) );
  XOR U1166 ( .A(in[1572]), .B(in[612]), .Z(n608) );
  XNOR U1167 ( .A(in[932]), .B(in[292]), .Z(n607) );
  XNOR U1168 ( .A(n608), .B(n607), .Z(n609) );
  XNOR U1169 ( .A(in[1252]), .B(n609), .Z(n820) );
  XOR U1170 ( .A(n610), .B(n820), .Z(n4278) );
  XOR U1171 ( .A(in[997]), .B(n4278), .Z(n1977) );
  NANDN U1172 ( .A(n1980), .B(n1977), .Z(n611) );
  XNOR U1173 ( .A(n1573), .B(n611), .Z(out[1017]) );
  XOR U1174 ( .A(in[1404]), .B(in[124]), .Z(n613) );
  XNOR U1175 ( .A(in[1084]), .B(in[764]), .Z(n612) );
  XNOR U1176 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U1177 ( .A(in[444]), .B(n614), .Z(n1663) );
  XOR U1178 ( .A(in[1533]), .B(in[573]), .Z(n616) );
  XNOR U1179 ( .A(in[1213]), .B(in[253]), .Z(n615) );
  XNOR U1180 ( .A(n616), .B(n615), .Z(n617) );
  XNOR U1181 ( .A(in[893]), .B(n617), .Z(n977) );
  XOR U1182 ( .A(n1663), .B(n977), .Z(n1869) );
  XOR U1183 ( .A(in[189]), .B(n1869), .Z(n1577) );
  XOR U1184 ( .A(in[158]), .B(in[1438]), .Z(n619) );
  XNOR U1185 ( .A(in[1118]), .B(in[798]), .Z(n618) );
  XNOR U1186 ( .A(n619), .B(n618), .Z(n620) );
  XNOR U1187 ( .A(in[478]), .B(n620), .Z(n916) );
  XOR U1188 ( .A(in[349]), .B(in[669]), .Z(n622) );
  XNOR U1189 ( .A(in[29]), .B(in[1309]), .Z(n621) );
  XNOR U1190 ( .A(n622), .B(n621), .Z(n623) );
  XOR U1191 ( .A(in[989]), .B(n623), .Z(n1475) );
  XNOR U1192 ( .A(in[1374]), .B(n4520), .Z(n1984) );
  XOR U1193 ( .A(in[1062]), .B(in[422]), .Z(n625) );
  XNOR U1194 ( .A(in[742]), .B(in[1382]), .Z(n624) );
  XNOR U1195 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U1196 ( .A(in[102]), .B(n626), .Z(n661) );
  XOR U1197 ( .A(in[1573]), .B(in[613]), .Z(n628) );
  XNOR U1198 ( .A(in[933]), .B(in[293]), .Z(n627) );
  XNOR U1199 ( .A(n628), .B(n627), .Z(n629) );
  XNOR U1200 ( .A(in[1253]), .B(n629), .Z(n979) );
  XOR U1201 ( .A(n661), .B(n979), .Z(n4284) );
  XOR U1202 ( .A(in[998]), .B(n4284), .Z(n1981) );
  NANDN U1203 ( .A(n1984), .B(n1981), .Z(n630) );
  XNOR U1204 ( .A(n1577), .B(n630), .Z(out[1018]) );
  XOR U1205 ( .A(in[1405]), .B(in[125]), .Z(n632) );
  XNOR U1206 ( .A(in[1085]), .B(in[765]), .Z(n631) );
  XNOR U1207 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U1208 ( .A(in[445]), .B(n633), .Z(n1667) );
  XOR U1209 ( .A(in[1534]), .B(in[894]), .Z(n635) );
  XNOR U1210 ( .A(in[574]), .B(in[1214]), .Z(n634) );
  XNOR U1211 ( .A(n635), .B(n634), .Z(n636) );
  XNOR U1212 ( .A(in[254]), .B(n636), .Z(n1114) );
  XOR U1213 ( .A(n1667), .B(n1114), .Z(n1891) );
  XOR U1214 ( .A(in[190]), .B(n1891), .Z(n1581) );
  XOR U1215 ( .A(in[1439]), .B(in[479]), .Z(n638) );
  XNOR U1216 ( .A(in[799]), .B(in[159]), .Z(n637) );
  XNOR U1217 ( .A(n638), .B(n637), .Z(n639) );
  XNOR U1218 ( .A(in[1119]), .B(n639), .Z(n931) );
  XOR U1219 ( .A(in[350]), .B(in[670]), .Z(n641) );
  XNOR U1220 ( .A(in[30]), .B(in[1310]), .Z(n640) );
  XNOR U1221 ( .A(n641), .B(n640), .Z(n642) );
  XOR U1222 ( .A(in[990]), .B(n642), .Z(n1479) );
  XNOR U1223 ( .A(in[1375]), .B(n4524), .Z(n1988) );
  XOR U1224 ( .A(in[1063]), .B(in[423]), .Z(n644) );
  XNOR U1225 ( .A(in[743]), .B(in[1383]), .Z(n643) );
  XNOR U1226 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U1227 ( .A(in[103]), .B(n645), .Z(n824) );
  XOR U1228 ( .A(in[1574]), .B(in[614]), .Z(n647) );
  XNOR U1229 ( .A(in[934]), .B(in[294]), .Z(n646) );
  XNOR U1230 ( .A(n647), .B(n646), .Z(n648) );
  XNOR U1231 ( .A(in[1254]), .B(n648), .Z(n1023) );
  XOR U1232 ( .A(n824), .B(n1023), .Z(n4286) );
  XOR U1233 ( .A(in[999]), .B(n4286), .Z(n1985) );
  NANDN U1234 ( .A(n1988), .B(n1985), .Z(n649) );
  XNOR U1235 ( .A(n1581), .B(n649), .Z(out[1019]) );
  XOR U1236 ( .A(in[1340]), .B(in[60]), .Z(n651) );
  XNOR U1237 ( .A(in[700]), .B(in[380]), .Z(n650) );
  XNOR U1238 ( .A(n651), .B(n650), .Z(n652) );
  XNOR U1239 ( .A(in[1020]), .B(n652), .Z(n1108) );
  XOR U1240 ( .A(n653), .B(n1108), .Z(n3957) );
  XOR U1241 ( .A(in[636]), .B(n3957), .Z(n2709) );
  IV U1242 ( .A(n2709), .Z(n2795) );
  XOR U1243 ( .A(in[162]), .B(in[1442]), .Z(n655) );
  XNOR U1244 ( .A(in[802]), .B(in[1122]), .Z(n654) );
  XNOR U1245 ( .A(n655), .B(n654), .Z(n656) );
  XOR U1246 ( .A(in[482]), .B(n656), .Z(n708) );
  XOR U1247 ( .A(n657), .B(n708), .Z(n3396) );
  IV U1248 ( .A(n3396), .Z(n4053) );
  XOR U1249 ( .A(in[227]), .B(n4053), .Z(n3137) );
  XOR U1250 ( .A(in[1511]), .B(in[551]), .Z(n659) );
  XNOR U1251 ( .A(in[871]), .B(in[231]), .Z(n658) );
  XNOR U1252 ( .A(n659), .B(n658), .Z(n660) );
  XNOR U1253 ( .A(in[1191]), .B(n660), .Z(n1514) );
  XNOR U1254 ( .A(n661), .B(n1514), .Z(n4093) );
  IV U1255 ( .A(n4093), .Z(n1268) );
  XOR U1256 ( .A(in[1447]), .B(n1268), .Z(n3134) );
  NANDN U1257 ( .A(n3137), .B(n3134), .Z(n662) );
  XOR U1258 ( .A(n2795), .B(n662), .Z(out[101]) );
  XOR U1259 ( .A(in[1406]), .B(in[126]), .Z(n664) );
  XNOR U1260 ( .A(in[1086]), .B(in[766]), .Z(n663) );
  XNOR U1261 ( .A(n664), .B(n663), .Z(n665) );
  XNOR U1262 ( .A(in[446]), .B(n665), .Z(n1672) );
  XOR U1263 ( .A(in[1535]), .B(in[575]), .Z(n667) );
  XNOR U1264 ( .A(in[895]), .B(in[255]), .Z(n666) );
  XNOR U1265 ( .A(n667), .B(n666), .Z(n668) );
  XNOR U1266 ( .A(in[1215]), .B(n668), .Z(n1262) );
  XOR U1267 ( .A(n1672), .B(n1262), .Z(n1921) );
  XOR U1268 ( .A(in[191]), .B(n1921), .Z(n1585) );
  XOR U1269 ( .A(in[1440]), .B(in[480]), .Z(n670) );
  XNOR U1270 ( .A(in[800]), .B(in[160]), .Z(n669) );
  XNOR U1271 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1272 ( .A(in[1120]), .B(n671), .Z(n946) );
  XOR U1273 ( .A(in[351]), .B(in[671]), .Z(n673) );
  XNOR U1274 ( .A(in[31]), .B(in[1311]), .Z(n672) );
  XNOR U1275 ( .A(n673), .B(n672), .Z(n674) );
  XOR U1276 ( .A(in[991]), .B(n674), .Z(n1483) );
  XNOR U1277 ( .A(in[1376]), .B(n4528), .Z(n1992) );
  XOR U1278 ( .A(in[1064]), .B(in[424]), .Z(n676) );
  XNOR U1279 ( .A(in[744]), .B(in[1384]), .Z(n675) );
  XNOR U1280 ( .A(n676), .B(n675), .Z(n677) );
  XNOR U1281 ( .A(in[104]), .B(n677), .Z(n983) );
  XOR U1282 ( .A(in[1575]), .B(in[615]), .Z(n679) );
  XNOR U1283 ( .A(in[935]), .B(in[295]), .Z(n678) );
  XNOR U1284 ( .A(n679), .B(n678), .Z(n680) );
  XNOR U1285 ( .A(in[1255]), .B(n680), .Z(n1036) );
  XOR U1286 ( .A(n983), .B(n1036), .Z(n4288) );
  XOR U1287 ( .A(in[1000]), .B(n4288), .Z(n1989) );
  NANDN U1288 ( .A(n1992), .B(n1989), .Z(n681) );
  XNOR U1289 ( .A(n1585), .B(n681), .Z(out[1020]) );
  XOR U1290 ( .A(in[1407]), .B(in[127]), .Z(n683) );
  XNOR U1291 ( .A(in[1087]), .B(in[767]), .Z(n682) );
  XNOR U1292 ( .A(n683), .B(n682), .Z(n684) );
  XNOR U1293 ( .A(in[447]), .B(n684), .Z(n1675) );
  XOR U1294 ( .A(in[1472]), .B(in[512]), .Z(n686) );
  XNOR U1295 ( .A(in[832]), .B(in[192]), .Z(n685) );
  XNOR U1296 ( .A(n686), .B(n685), .Z(n687) );
  XNOR U1297 ( .A(in[1152]), .B(n687), .Z(n1327) );
  XOR U1298 ( .A(n1675), .B(n1327), .Z(n1963) );
  XOR U1299 ( .A(in[128]), .B(n1963), .Z(n1589) );
  XOR U1300 ( .A(in[352]), .B(in[672]), .Z(n689) );
  XNOR U1301 ( .A(in[32]), .B(in[1312]), .Z(n688) );
  XNOR U1302 ( .A(n689), .B(n688), .Z(n690) );
  XOR U1303 ( .A(in[992]), .B(n690), .Z(n1485) );
  XNOR U1304 ( .A(in[1377]), .B(n4532), .Z(n1996) );
  XOR U1305 ( .A(in[1065]), .B(in[425]), .Z(n693) );
  XNOR U1306 ( .A(in[745]), .B(in[1385]), .Z(n692) );
  XNOR U1307 ( .A(n693), .B(n692), .Z(n694) );
  XNOR U1308 ( .A(in[105]), .B(n694), .Z(n1118) );
  XOR U1309 ( .A(in[1576]), .B(in[616]), .Z(n696) );
  XNOR U1310 ( .A(in[936]), .B(in[296]), .Z(n695) );
  XNOR U1311 ( .A(n696), .B(n695), .Z(n697) );
  XNOR U1312 ( .A(in[1256]), .B(n697), .Z(n1049) );
  XOR U1313 ( .A(n1118), .B(n1049), .Z(n4290) );
  XOR U1314 ( .A(in[1001]), .B(n4290), .Z(n1993) );
  NANDN U1315 ( .A(n1996), .B(n1993), .Z(n698) );
  XNOR U1316 ( .A(n1589), .B(n698), .Z(out[1021]) );
  XOR U1317 ( .A(in[1344]), .B(in[64]), .Z(n700) );
  XNOR U1318 ( .A(in[1024]), .B(in[384]), .Z(n699) );
  XNOR U1319 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1320 ( .A(in[704]), .B(n701), .Z(n1680) );
  XOR U1321 ( .A(in[1473]), .B(in[513]), .Z(n703) );
  XNOR U1322 ( .A(in[833]), .B(in[193]), .Z(n702) );
  XNOR U1323 ( .A(n703), .B(n702), .Z(n704) );
  XNOR U1324 ( .A(in[1153]), .B(n704), .Z(n1372) );
  XOR U1325 ( .A(n1680), .B(n1372), .Z(n2005) );
  XOR U1326 ( .A(in[129]), .B(n2005), .Z(n1593) );
  XOR U1327 ( .A(in[353]), .B(in[673]), .Z(n706) );
  XNOR U1328 ( .A(in[33]), .B(in[1313]), .Z(n705) );
  XNOR U1329 ( .A(n706), .B(n705), .Z(n707) );
  XNOR U1330 ( .A(in[993]), .B(n707), .Z(n1488) );
  XNOR U1331 ( .A(in[1378]), .B(n4536), .Z(n2000) );
  XOR U1332 ( .A(in[1577]), .B(in[617]), .Z(n710) );
  XNOR U1333 ( .A(in[937]), .B(in[297]), .Z(n709) );
  XNOR U1334 ( .A(n710), .B(n709), .Z(n711) );
  XNOR U1335 ( .A(in[1257]), .B(n711), .Z(n1062) );
  XOR U1336 ( .A(n712), .B(n1062), .Z(n4292) );
  XOR U1337 ( .A(in[1002]), .B(n4292), .Z(n1997) );
  NANDN U1338 ( .A(n2000), .B(n1997), .Z(n713) );
  XNOR U1339 ( .A(n1593), .B(n713), .Z(out[1022]) );
  IV U1340 ( .A(n3171), .Z(n3932) );
  XOR U1341 ( .A(n3932), .B(in[130]), .Z(n1595) );
  XOR U1342 ( .A(in[354]), .B(in[674]), .Z(n715) );
  XNOR U1343 ( .A(in[34]), .B(in[1314]), .Z(n714) );
  XNOR U1344 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1345 ( .A(in[994]), .B(n716), .Z(n1491) );
  XOR U1346 ( .A(in[163]), .B(in[1443]), .Z(n718) );
  XNOR U1347 ( .A(in[803]), .B(in[1123]), .Z(n717) );
  XNOR U1348 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1349 ( .A(in[483]), .B(n719), .Z(n819) );
  XNOR U1350 ( .A(in[1379]), .B(n4540), .Z(n2004) );
  XOR U1351 ( .A(in[1578]), .B(in[618]), .Z(n721) );
  XNOR U1352 ( .A(in[938]), .B(in[298]), .Z(n720) );
  XNOR U1353 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U1354 ( .A(in[1258]), .B(n722), .Z(n1075) );
  XOR U1355 ( .A(n723), .B(n1075), .Z(n4294) );
  XOR U1356 ( .A(in[1003]), .B(n4294), .Z(n2001) );
  NANDN U1357 ( .A(n2004), .B(n2001), .Z(n724) );
  XOR U1358 ( .A(n1595), .B(n724), .Z(out[1023]) );
  XNOR U1359 ( .A(n726), .B(n725), .Z(n3985) );
  XOR U1360 ( .A(in[531]), .B(n3985), .Z(n1599) );
  XOR U1361 ( .A(in[35]), .B(in[675]), .Z(n728) );
  XNOR U1362 ( .A(in[355]), .B(in[1315]), .Z(n727) );
  XNOR U1363 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1364 ( .A(in[995]), .B(n729), .Z(n1494) );
  XOR U1365 ( .A(in[164]), .B(in[1444]), .Z(n731) );
  XNOR U1366 ( .A(in[804]), .B(in[1124]), .Z(n730) );
  XNOR U1367 ( .A(n731), .B(n730), .Z(n732) );
  XNOR U1368 ( .A(in[484]), .B(n732), .Z(n978) );
  XOR U1369 ( .A(n1494), .B(n978), .Z(n4544) );
  XNOR U1370 ( .A(in[1380]), .B(n4544), .Z(n4992) );
  XOR U1371 ( .A(in[1346]), .B(in[66]), .Z(n734) );
  XNOR U1372 ( .A(in[1026]), .B(in[386]), .Z(n733) );
  XNOR U1373 ( .A(n734), .B(n733), .Z(n735) );
  XNOR U1374 ( .A(in[706]), .B(n735), .Z(n1688) );
  XOR U1375 ( .A(in[1475]), .B(in[515]), .Z(n737) );
  XNOR U1376 ( .A(in[835]), .B(in[195]), .Z(n736) );
  XNOR U1377 ( .A(n737), .B(n736), .Z(n738) );
  XOR U1378 ( .A(in[1155]), .B(n738), .Z(n1415) );
  XOR U1379 ( .A(in[131]), .B(n3173), .Z(n4994) );
  OR U1380 ( .A(n4992), .B(n4994), .Z(n739) );
  XNOR U1381 ( .A(n1599), .B(n739), .Z(out[1024]) );
  XNOR U1382 ( .A(n741), .B(n740), .Z(n3989) );
  XOR U1383 ( .A(in[532]), .B(n3989), .Z(n1603) );
  XOR U1384 ( .A(in[1445]), .B(in[165]), .Z(n743) );
  XNOR U1385 ( .A(in[805]), .B(in[1125]), .Z(n742) );
  XNOR U1386 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U1387 ( .A(in[485]), .B(n744), .Z(n1022) );
  XOR U1388 ( .A(in[36]), .B(in[676]), .Z(n746) );
  XNOR U1389 ( .A(in[356]), .B(in[1316]), .Z(n745) );
  XNOR U1390 ( .A(n746), .B(n745), .Z(n747) );
  XNOR U1391 ( .A(in[996]), .B(n747), .Z(n1497) );
  XOR U1392 ( .A(n1022), .B(n1497), .Z(n4550) );
  XNOR U1393 ( .A(in[1381]), .B(n4550), .Z(n4996) );
  XOR U1394 ( .A(in[1347]), .B(in[67]), .Z(n749) );
  XNOR U1395 ( .A(in[1027]), .B(in[387]), .Z(n748) );
  XNOR U1396 ( .A(n749), .B(n748), .Z(n750) );
  XNOR U1397 ( .A(in[707]), .B(n750), .Z(n1692) );
  XOR U1398 ( .A(in[1476]), .B(in[516]), .Z(n752) );
  XNOR U1399 ( .A(in[836]), .B(in[196]), .Z(n751) );
  XNOR U1400 ( .A(n752), .B(n751), .Z(n753) );
  XOR U1401 ( .A(in[1156]), .B(n753), .Z(n1417) );
  XOR U1402 ( .A(in[132]), .B(n3175), .Z(n4998) );
  OR U1403 ( .A(n4996), .B(n4998), .Z(n754) );
  XNOR U1404 ( .A(n1603), .B(n754), .Z(out[1025]) );
  XOR U1405 ( .A(n756), .B(n755), .Z(n2008) );
  XOR U1406 ( .A(in[533]), .B(n2008), .Z(n1607) );
  XOR U1407 ( .A(in[166]), .B(in[806]), .Z(n758) );
  XNOR U1408 ( .A(in[1126]), .B(in[486]), .Z(n757) );
  XNOR U1409 ( .A(n758), .B(n757), .Z(n759) );
  XNOR U1410 ( .A(in[1446]), .B(n759), .Z(n1035) );
  XOR U1411 ( .A(in[37]), .B(in[677]), .Z(n761) );
  XNOR U1412 ( .A(in[357]), .B(in[1317]), .Z(n760) );
  XNOR U1413 ( .A(n761), .B(n760), .Z(n762) );
  XNOR U1414 ( .A(in[997]), .B(n762), .Z(n1500) );
  XOR U1415 ( .A(n1035), .B(n1500), .Z(n4552) );
  XNOR U1416 ( .A(in[1382]), .B(n4552), .Z(n5000) );
  XOR U1417 ( .A(in[1348]), .B(in[68]), .Z(n764) );
  XNOR U1418 ( .A(in[1028]), .B(in[388]), .Z(n763) );
  XNOR U1419 ( .A(n764), .B(n763), .Z(n765) );
  XNOR U1420 ( .A(in[708]), .B(n765), .Z(n1696) );
  XOR U1421 ( .A(in[1477]), .B(in[517]), .Z(n767) );
  XNOR U1422 ( .A(in[837]), .B(in[197]), .Z(n766) );
  XNOR U1423 ( .A(n767), .B(n766), .Z(n768) );
  XOR U1424 ( .A(in[1157]), .B(n768), .Z(n1419) );
  XOR U1425 ( .A(in[133]), .B(n3177), .Z(n5002) );
  OR U1426 ( .A(n5000), .B(n5002), .Z(n769) );
  XNOR U1427 ( .A(n1607), .B(n769), .Z(out[1026]) );
  XNOR U1428 ( .A(n771), .B(n770), .Z(n3997) );
  XOR U1429 ( .A(in[534]), .B(n3997), .Z(n1611) );
  XOR U1430 ( .A(in[167]), .B(in[807]), .Z(n773) );
  XNOR U1431 ( .A(in[1127]), .B(in[487]), .Z(n772) );
  XNOR U1432 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U1433 ( .A(in[1447]), .B(n774), .Z(n1048) );
  XOR U1434 ( .A(in[38]), .B(in[678]), .Z(n776) );
  XNOR U1435 ( .A(in[358]), .B(in[1318]), .Z(n775) );
  XNOR U1436 ( .A(n776), .B(n775), .Z(n777) );
  XNOR U1437 ( .A(in[998]), .B(n777), .Z(n1504) );
  XOR U1438 ( .A(n1048), .B(n1504), .Z(n4333) );
  XNOR U1439 ( .A(in[1383]), .B(n4333), .Z(n5004) );
  XOR U1440 ( .A(in[1349]), .B(in[69]), .Z(n779) );
  XNOR U1441 ( .A(in[1029]), .B(in[389]), .Z(n778) );
  XNOR U1442 ( .A(n779), .B(n778), .Z(n780) );
  XNOR U1443 ( .A(in[709]), .B(n780), .Z(n1700) );
  XOR U1444 ( .A(in[1478]), .B(in[518]), .Z(n782) );
  XNOR U1445 ( .A(in[838]), .B(in[198]), .Z(n781) );
  XNOR U1446 ( .A(n782), .B(n781), .Z(n783) );
  XOR U1447 ( .A(in[1158]), .B(n783), .Z(n1421) );
  XOR U1448 ( .A(in[134]), .B(n3179), .Z(n5006) );
  OR U1449 ( .A(n5004), .B(n5006), .Z(n784) );
  XNOR U1450 ( .A(n1611), .B(n784), .Z(out[1027]) );
  XNOR U1451 ( .A(n786), .B(n785), .Z(n4001) );
  XOR U1452 ( .A(in[535]), .B(n4001), .Z(n1615) );
  XOR U1453 ( .A(in[39]), .B(in[679]), .Z(n788) );
  XNOR U1454 ( .A(in[359]), .B(in[1319]), .Z(n787) );
  XNOR U1455 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1456 ( .A(in[999]), .B(n789), .Z(n1509) );
  XOR U1457 ( .A(in[168]), .B(in[1448]), .Z(n791) );
  XNOR U1458 ( .A(in[1128]), .B(in[808]), .Z(n790) );
  XNOR U1459 ( .A(n791), .B(n790), .Z(n792) );
  XNOR U1460 ( .A(in[488]), .B(n792), .Z(n1061) );
  XOR U1461 ( .A(n1509), .B(n1061), .Z(n4335) );
  XNOR U1462 ( .A(in[1384]), .B(n4335), .Z(n5008) );
  XOR U1463 ( .A(in[1350]), .B(in[70]), .Z(n794) );
  XNOR U1464 ( .A(in[1030]), .B(in[390]), .Z(n793) );
  XNOR U1465 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U1466 ( .A(in[710]), .B(n795), .Z(n1704) );
  XOR U1467 ( .A(in[199]), .B(in[1479]), .Z(n797) );
  XNOR U1468 ( .A(in[1159]), .B(in[839]), .Z(n796) );
  XNOR U1469 ( .A(n797), .B(n796), .Z(n798) );
  XOR U1470 ( .A(in[519]), .B(n798), .Z(n1423) );
  XOR U1471 ( .A(in[135]), .B(n3181), .Z(n5010) );
  OR U1472 ( .A(n5008), .B(n5010), .Z(n799) );
  XNOR U1473 ( .A(n1615), .B(n799), .Z(out[1028]) );
  XOR U1474 ( .A(n801), .B(n800), .Z(n2012) );
  XOR U1475 ( .A(in[536]), .B(n2012), .Z(n1619) );
  XOR U1476 ( .A(in[680]), .B(in[1320]), .Z(n803) );
  XNOR U1477 ( .A(in[40]), .B(in[360]), .Z(n802) );
  XNOR U1478 ( .A(n803), .B(n802), .Z(n804) );
  XNOR U1479 ( .A(in[1000]), .B(n804), .Z(n1513) );
  XOR U1480 ( .A(in[169]), .B(in[1449]), .Z(n806) );
  XNOR U1481 ( .A(in[1129]), .B(in[809]), .Z(n805) );
  XNOR U1482 ( .A(n806), .B(n805), .Z(n807) );
  XNOR U1483 ( .A(in[489]), .B(n807), .Z(n1074) );
  XOR U1484 ( .A(n1513), .B(n1074), .Z(n4341) );
  XNOR U1485 ( .A(in[1385]), .B(n4341), .Z(n5012) );
  XOR U1486 ( .A(in[1351]), .B(in[711]), .Z(n809) );
  XNOR U1487 ( .A(in[1031]), .B(in[391]), .Z(n808) );
  XNOR U1488 ( .A(n809), .B(n808), .Z(n810) );
  XNOR U1489 ( .A(in[71]), .B(n810), .Z(n1708) );
  XOR U1490 ( .A(in[1480]), .B(in[520]), .Z(n812) );
  XNOR U1491 ( .A(in[840]), .B(in[200]), .Z(n811) );
  XNOR U1492 ( .A(n812), .B(n811), .Z(n813) );
  XOR U1493 ( .A(in[1160]), .B(n813), .Z(n1428) );
  XOR U1494 ( .A(in[136]), .B(n3183), .Z(n5014) );
  OR U1495 ( .A(n5012), .B(n5014), .Z(n814) );
  XNOR U1496 ( .A(n1619), .B(n814), .Z(out[1029]) );
  XOR U1497 ( .A(in[1341]), .B(in[61]), .Z(n816) );
  XNOR U1498 ( .A(in[701]), .B(in[381]), .Z(n815) );
  XNOR U1499 ( .A(n816), .B(n815), .Z(n817) );
  XNOR U1500 ( .A(in[1021]), .B(n817), .Z(n1131) );
  XOR U1501 ( .A(n818), .B(n1131), .Z(n3961) );
  XOR U1502 ( .A(in[637]), .B(n3961), .Z(n2711) );
  IV U1503 ( .A(n2711), .Z(n2800) );
  XOR U1504 ( .A(n820), .B(n819), .Z(n3400) );
  IV U1505 ( .A(n3400), .Z(n4057) );
  XOR U1506 ( .A(in[228]), .B(n4057), .Z(n3156) );
  XOR U1507 ( .A(in[1512]), .B(in[552]), .Z(n822) );
  XNOR U1508 ( .A(in[872]), .B(in[232]), .Z(n821) );
  XNOR U1509 ( .A(n822), .B(n821), .Z(n823) );
  XNOR U1510 ( .A(in[1192]), .B(n823), .Z(n1518) );
  XNOR U1511 ( .A(n824), .B(n1518), .Z(n4097) );
  IV U1512 ( .A(n4097), .Z(n1280) );
  XOR U1513 ( .A(in[1448]), .B(n1280), .Z(n3154) );
  NANDN U1514 ( .A(n3156), .B(n3154), .Z(n825) );
  XOR U1515 ( .A(n2800), .B(n825), .Z(out[102]) );
  XOR U1516 ( .A(n827), .B(n826), .Z(n2015) );
  XOR U1517 ( .A(in[537]), .B(n2015), .Z(n1623) );
  XOR U1518 ( .A(in[1352]), .B(in[712]), .Z(n829) );
  XNOR U1519 ( .A(in[1032]), .B(in[392]), .Z(n828) );
  XNOR U1520 ( .A(n829), .B(n828), .Z(n830) );
  XNOR U1521 ( .A(in[72]), .B(n830), .Z(n1713) );
  XOR U1522 ( .A(in[1481]), .B(in[521]), .Z(n832) );
  XNOR U1523 ( .A(in[841]), .B(in[201]), .Z(n831) );
  XNOR U1524 ( .A(n832), .B(n831), .Z(n833) );
  XOR U1525 ( .A(in[1161]), .B(n833), .Z(n1430) );
  XOR U1526 ( .A(in[137]), .B(n3185), .Z(n5018) );
  XOR U1527 ( .A(in[170]), .B(in[1450]), .Z(n835) );
  XNOR U1528 ( .A(in[1130]), .B(in[810]), .Z(n834) );
  XNOR U1529 ( .A(n835), .B(n834), .Z(n836) );
  XNOR U1530 ( .A(in[490]), .B(n836), .Z(n1090) );
  XOR U1531 ( .A(in[681]), .B(in[1321]), .Z(n838) );
  XNOR U1532 ( .A(in[41]), .B(in[361]), .Z(n837) );
  XNOR U1533 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U1534 ( .A(in[1001]), .B(n839), .Z(n1517) );
  XOR U1535 ( .A(n1090), .B(n1517), .Z(n4343) );
  XOR U1536 ( .A(in[1386]), .B(n4343), .Z(n5015) );
  NANDN U1537 ( .A(n5018), .B(n5015), .Z(n840) );
  XNOR U1538 ( .A(n1623), .B(n840), .Z(out[1030]) );
  XNOR U1539 ( .A(n842), .B(n841), .Z(n4013) );
  XOR U1540 ( .A(in[538]), .B(n4013), .Z(n1627) );
  XOR U1541 ( .A(in[1353]), .B(in[393]), .Z(n844) );
  XNOR U1542 ( .A(in[713]), .B(in[73]), .Z(n843) );
  XNOR U1543 ( .A(n844), .B(n843), .Z(n845) );
  XNOR U1544 ( .A(in[1033]), .B(n845), .Z(n1717) );
  XOR U1545 ( .A(in[1482]), .B(in[522]), .Z(n847) );
  XNOR U1546 ( .A(in[842]), .B(in[202]), .Z(n846) );
  XNOR U1547 ( .A(n847), .B(n846), .Z(n848) );
  XOR U1548 ( .A(n1717), .B(n234), .Z(n3187) );
  XOR U1549 ( .A(in[138]), .B(n3187), .Z(n5022) );
  XOR U1550 ( .A(in[811]), .B(in[491]), .Z(n850) );
  XNOR U1551 ( .A(in[1451]), .B(in[1131]), .Z(n849) );
  XNOR U1552 ( .A(n850), .B(n849), .Z(n851) );
  XNOR U1553 ( .A(in[171]), .B(n851), .Z(n1103) );
  XOR U1554 ( .A(in[682]), .B(in[1322]), .Z(n853) );
  XNOR U1555 ( .A(in[42]), .B(in[362]), .Z(n852) );
  XNOR U1556 ( .A(n853), .B(n852), .Z(n854) );
  XNOR U1557 ( .A(in[1002]), .B(n854), .Z(n1522) );
  XOR U1558 ( .A(n1103), .B(n1522), .Z(n4345) );
  XOR U1559 ( .A(in[1387]), .B(n4345), .Z(n5019) );
  NANDN U1560 ( .A(n5022), .B(n5019), .Z(n855) );
  XNOR U1561 ( .A(n1627), .B(n855), .Z(out[1031]) );
  XNOR U1562 ( .A(n857), .B(n856), .Z(n4017) );
  XOR U1563 ( .A(in[539]), .B(n4017), .Z(n1632) );
  XOR U1564 ( .A(in[1354]), .B(in[714]), .Z(n859) );
  XNOR U1565 ( .A(in[74]), .B(in[394]), .Z(n858) );
  XNOR U1566 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U1567 ( .A(in[1034]), .B(n860), .Z(n1721) );
  XOR U1568 ( .A(in[1483]), .B(in[523]), .Z(n862) );
  XNOR U1569 ( .A(in[843]), .B(in[203]), .Z(n861) );
  XNOR U1570 ( .A(n862), .B(n861), .Z(n863) );
  XOR U1571 ( .A(in[1163]), .B(n863), .Z(n1433) );
  XOR U1572 ( .A(n2298), .B(in[139]), .Z(n5026) );
  XOR U1573 ( .A(in[683]), .B(in[1323]), .Z(n865) );
  XNOR U1574 ( .A(in[43]), .B(in[363]), .Z(n864) );
  XNOR U1575 ( .A(n865), .B(n864), .Z(n866) );
  XNOR U1576 ( .A(in[1003]), .B(n866), .Z(n1526) );
  XOR U1577 ( .A(in[812]), .B(in[492]), .Z(n868) );
  XNOR U1578 ( .A(in[1452]), .B(in[1132]), .Z(n867) );
  XNOR U1579 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1580 ( .A(in[172]), .B(n869), .Z(n1123) );
  XOR U1581 ( .A(n1526), .B(n1123), .Z(n4348) );
  XOR U1582 ( .A(in[1388]), .B(n4348), .Z(n5023) );
  NANDN U1583 ( .A(n5026), .B(n5023), .Z(n870) );
  XNOR U1584 ( .A(n1632), .B(n870), .Z(out[1032]) );
  XOR U1585 ( .A(n872), .B(n871), .Z(n4021) );
  XOR U1586 ( .A(in[540]), .B(n4021), .Z(n1636) );
  XOR U1587 ( .A(in[1355]), .B(in[715]), .Z(n874) );
  XNOR U1588 ( .A(in[1035]), .B(in[395]), .Z(n873) );
  XNOR U1589 ( .A(n874), .B(n873), .Z(n875) );
  XNOR U1590 ( .A(in[75]), .B(n875), .Z(n1725) );
  XOR U1591 ( .A(in[1484]), .B(in[524]), .Z(n877) );
  XNOR U1592 ( .A(in[844]), .B(in[204]), .Z(n876) );
  XNOR U1593 ( .A(n877), .B(n876), .Z(n878) );
  XOR U1594 ( .A(n1725), .B(n235), .Z(n3194) );
  XOR U1595 ( .A(in[140]), .B(n3194), .Z(n5030) );
  XOR U1596 ( .A(in[1324]), .B(in[44]), .Z(n880) );
  XNOR U1597 ( .A(in[684]), .B(in[364]), .Z(n879) );
  XNOR U1598 ( .A(n880), .B(n879), .Z(n881) );
  XNOR U1599 ( .A(in[1004]), .B(n881), .Z(n1529) );
  XOR U1600 ( .A(in[813]), .B(in[493]), .Z(n883) );
  XNOR U1601 ( .A(in[1453]), .B(in[1133]), .Z(n882) );
  XNOR U1602 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U1603 ( .A(in[173]), .B(n884), .Z(n1136) );
  XOR U1604 ( .A(n1529), .B(n1136), .Z(n4351) );
  XOR U1605 ( .A(in[1389]), .B(n4351), .Z(n5027) );
  NANDN U1606 ( .A(n5030), .B(n5027), .Z(n885) );
  XNOR U1607 ( .A(n1636), .B(n885), .Z(out[1033]) );
  XOR U1608 ( .A(n887), .B(n886), .Z(n4029) );
  XOR U1609 ( .A(in[541]), .B(n4029), .Z(n1640) );
  XOR U1610 ( .A(in[76]), .B(in[1036]), .Z(n889) );
  XNOR U1611 ( .A(in[716]), .B(in[396]), .Z(n888) );
  XNOR U1612 ( .A(n889), .B(n888), .Z(n890) );
  XNOR U1613 ( .A(in[1356]), .B(n890), .Z(n1729) );
  XOR U1614 ( .A(in[1485]), .B(in[525]), .Z(n892) );
  XNOR U1615 ( .A(in[845]), .B(in[205]), .Z(n891) );
  XNOR U1616 ( .A(n892), .B(n891), .Z(n893) );
  XOR U1617 ( .A(in[1165]), .B(n893), .Z(n1436) );
  XOR U1618 ( .A(in[141]), .B(n3196), .Z(n5038) );
  XOR U1619 ( .A(in[814]), .B(in[494]), .Z(n895) );
  XNOR U1620 ( .A(in[1454]), .B(in[1134]), .Z(n894) );
  XNOR U1621 ( .A(n895), .B(n894), .Z(n896) );
  XNOR U1622 ( .A(in[174]), .B(n896), .Z(n1149) );
  XOR U1623 ( .A(in[1325]), .B(in[45]), .Z(n898) );
  XNOR U1624 ( .A(in[685]), .B(in[365]), .Z(n897) );
  XNOR U1625 ( .A(n898), .B(n897), .Z(n899) );
  XNOR U1626 ( .A(in[1005]), .B(n899), .Z(n1533) );
  XOR U1627 ( .A(n1149), .B(n1533), .Z(n4354) );
  XOR U1628 ( .A(in[1390]), .B(n4354), .Z(n5035) );
  NANDN U1629 ( .A(n5038), .B(n5035), .Z(n900) );
  XNOR U1630 ( .A(n1640), .B(n900), .Z(out[1034]) );
  XOR U1631 ( .A(n902), .B(n901), .Z(n4033) );
  XOR U1632 ( .A(in[542]), .B(n4033), .Z(n1644) );
  XOR U1633 ( .A(in[77]), .B(in[1037]), .Z(n904) );
  XNOR U1634 ( .A(in[717]), .B(in[397]), .Z(n903) );
  XNOR U1635 ( .A(n904), .B(n903), .Z(n905) );
  XNOR U1636 ( .A(in[1357]), .B(n905), .Z(n1733) );
  XOR U1637 ( .A(in[1486]), .B(in[526]), .Z(n907) );
  XNOR U1638 ( .A(in[846]), .B(in[206]), .Z(n906) );
  XNOR U1639 ( .A(n907), .B(n906), .Z(n908) );
  XOR U1640 ( .A(n1733), .B(n236), .Z(n3199) );
  XOR U1641 ( .A(in[142]), .B(n3199), .Z(n5042) );
  XOR U1642 ( .A(in[1326]), .B(in[46]), .Z(n910) );
  XNOR U1643 ( .A(in[686]), .B(in[366]), .Z(n909) );
  XNOR U1644 ( .A(n910), .B(n909), .Z(n911) );
  XNOR U1645 ( .A(in[1006]), .B(n911), .Z(n1537) );
  XOR U1646 ( .A(in[815]), .B(in[495]), .Z(n913) );
  XNOR U1647 ( .A(in[1455]), .B(in[1135]), .Z(n912) );
  XNOR U1648 ( .A(n913), .B(n912), .Z(n914) );
  XNOR U1649 ( .A(in[175]), .B(n914), .Z(n1162) );
  XOR U1650 ( .A(n1537), .B(n1162), .Z(n4356) );
  XOR U1651 ( .A(in[1391]), .B(n4356), .Z(n5039) );
  NANDN U1652 ( .A(n5042), .B(n5039), .Z(n915) );
  XNOR U1653 ( .A(n1644), .B(n915), .Z(out[1035]) );
  XOR U1654 ( .A(n917), .B(n916), .Z(n4037) );
  XOR U1655 ( .A(in[543]), .B(n4037), .Z(n1648) );
  XOR U1656 ( .A(in[78]), .B(in[1038]), .Z(n919) );
  XNOR U1657 ( .A(in[718]), .B(in[398]), .Z(n918) );
  XNOR U1658 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U1659 ( .A(in[1358]), .B(n920), .Z(n1737) );
  XOR U1660 ( .A(in[1487]), .B(in[527]), .Z(n922) );
  XNOR U1661 ( .A(in[847]), .B(in[207]), .Z(n921) );
  XNOR U1662 ( .A(n922), .B(n921), .Z(n923) );
  XOR U1663 ( .A(n1737), .B(n237), .Z(n3202) );
  XOR U1664 ( .A(in[143]), .B(n3202), .Z(n5046) );
  XOR U1665 ( .A(in[816]), .B(in[496]), .Z(n925) );
  XNOR U1666 ( .A(in[1456]), .B(in[1136]), .Z(n924) );
  XNOR U1667 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U1668 ( .A(in[176]), .B(n926), .Z(n1177) );
  XOR U1669 ( .A(in[1327]), .B(in[47]), .Z(n928) );
  XNOR U1670 ( .A(in[687]), .B(in[367]), .Z(n927) );
  XNOR U1671 ( .A(n928), .B(n927), .Z(n929) );
  XNOR U1672 ( .A(in[1007]), .B(n929), .Z(n1541) );
  XOR U1673 ( .A(n1177), .B(n1541), .Z(n4359) );
  XOR U1674 ( .A(in[1392]), .B(n4359), .Z(n5043) );
  NANDN U1675 ( .A(n5046), .B(n5043), .Z(n930) );
  XNOR U1676 ( .A(n1648), .B(n930), .Z(out[1036]) );
  XOR U1677 ( .A(n932), .B(n931), .Z(n4041) );
  XOR U1678 ( .A(in[544]), .B(n4041), .Z(n1652) );
  XOR U1679 ( .A(in[79]), .B(in[1039]), .Z(n934) );
  XNOR U1680 ( .A(in[719]), .B(in[399]), .Z(n933) );
  XNOR U1681 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U1682 ( .A(in[1359]), .B(n935), .Z(n1741) );
  XOR U1683 ( .A(in[1488]), .B(in[528]), .Z(n937) );
  XNOR U1684 ( .A(in[848]), .B(in[208]), .Z(n936) );
  XNOR U1685 ( .A(n937), .B(n936), .Z(n938) );
  XOR U1686 ( .A(in[1168]), .B(n938), .Z(n1440) );
  XOR U1687 ( .A(in[144]), .B(n3205), .Z(n5050) );
  XOR U1688 ( .A(in[1328]), .B(in[48]), .Z(n940) );
  XNOR U1689 ( .A(in[688]), .B(in[368]), .Z(n939) );
  XNOR U1690 ( .A(n940), .B(n939), .Z(n941) );
  XNOR U1691 ( .A(in[1008]), .B(n941), .Z(n1545) );
  XOR U1692 ( .A(in[817]), .B(in[497]), .Z(n943) );
  XNOR U1693 ( .A(in[1457]), .B(in[1137]), .Z(n942) );
  XNOR U1694 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U1695 ( .A(in[177]), .B(n944), .Z(n1192) );
  XOR U1696 ( .A(n1545), .B(n1192), .Z(n4362) );
  XOR U1697 ( .A(in[1393]), .B(n4362), .Z(n5047) );
  NANDN U1698 ( .A(n5050), .B(n5047), .Z(n945) );
  XNOR U1699 ( .A(n1652), .B(n945), .Z(out[1037]) );
  XOR U1700 ( .A(n947), .B(n946), .Z(n4045) );
  XOR U1701 ( .A(in[545]), .B(n4045), .Z(n1656) );
  XOR U1702 ( .A(in[80]), .B(in[1040]), .Z(n949) );
  XNOR U1703 ( .A(in[720]), .B(in[400]), .Z(n948) );
  XNOR U1704 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1705 ( .A(in[1360]), .B(n950), .Z(n1745) );
  XOR U1706 ( .A(in[1489]), .B(in[529]), .Z(n952) );
  XNOR U1707 ( .A(in[849]), .B(in[209]), .Z(n951) );
  XNOR U1708 ( .A(n952), .B(n951), .Z(n953) );
  XOR U1709 ( .A(in[1169]), .B(n953), .Z(n1442) );
  XOR U1710 ( .A(in[145]), .B(n3208), .Z(n5054) );
  XOR U1711 ( .A(in[1329]), .B(in[49]), .Z(n955) );
  XNOR U1712 ( .A(in[689]), .B(in[369]), .Z(n954) );
  XNOR U1713 ( .A(n955), .B(n954), .Z(n956) );
  XNOR U1714 ( .A(in[1009]), .B(n956), .Z(n1551) );
  XOR U1715 ( .A(in[818]), .B(in[498]), .Z(n958) );
  XNOR U1716 ( .A(in[1458]), .B(in[1138]), .Z(n957) );
  XNOR U1717 ( .A(n958), .B(n957), .Z(n959) );
  XNOR U1718 ( .A(in[178]), .B(n959), .Z(n1207) );
  XOR U1719 ( .A(n1551), .B(n1207), .Z(n4365) );
  XOR U1720 ( .A(in[1394]), .B(n4365), .Z(n5051) );
  NANDN U1721 ( .A(n5054), .B(n5051), .Z(n960) );
  XNOR U1722 ( .A(n1656), .B(n960), .Z(out[1038]) );
  IV U1723 ( .A(n4049), .Z(n3393) );
  XOR U1724 ( .A(n3393), .B(in[546]), .Z(n1660) );
  XOR U1725 ( .A(in[81]), .B(in[1041]), .Z(n962) );
  XNOR U1726 ( .A(in[721]), .B(in[401]), .Z(n961) );
  XNOR U1727 ( .A(n962), .B(n961), .Z(n963) );
  XNOR U1728 ( .A(in[1361]), .B(n963), .Z(n1749) );
  XOR U1729 ( .A(in[1490]), .B(in[530]), .Z(n965) );
  XNOR U1730 ( .A(in[850]), .B(in[210]), .Z(n964) );
  XNOR U1731 ( .A(n965), .B(n964), .Z(n966) );
  XOR U1732 ( .A(in[1170]), .B(n966), .Z(n1446) );
  XOR U1733 ( .A(in[146]), .B(n4002), .Z(n5058) );
  XOR U1734 ( .A(in[1330]), .B(in[50]), .Z(n968) );
  XNOR U1735 ( .A(in[690]), .B(in[370]), .Z(n967) );
  XNOR U1736 ( .A(n968), .B(n967), .Z(n969) );
  XNOR U1737 ( .A(in[1010]), .B(n969), .Z(n1555) );
  XOR U1738 ( .A(in[819]), .B(in[499]), .Z(n971) );
  XNOR U1739 ( .A(in[1459]), .B(in[1139]), .Z(n970) );
  XNOR U1740 ( .A(n971), .B(n970), .Z(n972) );
  XNOR U1741 ( .A(in[179]), .B(n972), .Z(n1222) );
  XOR U1742 ( .A(n1555), .B(n1222), .Z(n4372) );
  XOR U1743 ( .A(in[1395]), .B(n4372), .Z(n5055) );
  NANDN U1744 ( .A(n5058), .B(n5055), .Z(n973) );
  XOR U1745 ( .A(n1660), .B(n973), .Z(out[1039]) );
  XOR U1746 ( .A(in[1342]), .B(in[62]), .Z(n975) );
  XNOR U1747 ( .A(in[702]), .B(in[382]), .Z(n974) );
  XNOR U1748 ( .A(n975), .B(n974), .Z(n976) );
  XNOR U1749 ( .A(in[1022]), .B(n976), .Z(n1144) );
  XOR U1750 ( .A(n977), .B(n1144), .Z(n3965) );
  XOR U1751 ( .A(in[638]), .B(n3965), .Z(n2713) );
  IV U1752 ( .A(n2713), .Z(n2802) );
  XOR U1753 ( .A(n979), .B(n978), .Z(n4061) );
  XOR U1754 ( .A(in[229]), .B(n4061), .Z(n3167) );
  XOR U1755 ( .A(in[1513]), .B(in[553]), .Z(n981) );
  XNOR U1756 ( .A(in[873]), .B(in[233]), .Z(n980) );
  XNOR U1757 ( .A(n981), .B(n980), .Z(n982) );
  XNOR U1758 ( .A(in[1193]), .B(n982), .Z(n1521) );
  XNOR U1759 ( .A(n983), .B(n1521), .Z(n4101) );
  IV U1760 ( .A(n4101), .Z(n1292) );
  XOR U1761 ( .A(in[1449]), .B(n1292), .Z(n3164) );
  NANDN U1762 ( .A(n3167), .B(n3164), .Z(n984) );
  XOR U1763 ( .A(n2802), .B(n984), .Z(out[103]) );
  XOR U1764 ( .A(n3396), .B(in[547]), .Z(n1664) );
  XOR U1765 ( .A(in[1042]), .B(in[402]), .Z(n986) );
  XNOR U1766 ( .A(in[722]), .B(in[82]), .Z(n985) );
  XNOR U1767 ( .A(n986), .B(n985), .Z(n987) );
  XNOR U1768 ( .A(in[1362]), .B(n987), .Z(n1754) );
  XOR U1769 ( .A(in[851]), .B(in[1171]), .Z(n989) );
  XNOR U1770 ( .A(in[1491]), .B(in[211]), .Z(n988) );
  XNOR U1771 ( .A(n989), .B(n988), .Z(n990) );
  XOR U1772 ( .A(in[531]), .B(n990), .Z(n1448) );
  IV U1773 ( .A(n3213), .Z(n4006) );
  XNOR U1774 ( .A(in[147]), .B(n4006), .Z(n5061) );
  XOR U1775 ( .A(in[1331]), .B(in[51]), .Z(n992) );
  XNOR U1776 ( .A(in[691]), .B(in[371]), .Z(n991) );
  XNOR U1777 ( .A(n992), .B(n991), .Z(n993) );
  XNOR U1778 ( .A(in[1011]), .B(n993), .Z(n1559) );
  XOR U1779 ( .A(in[820]), .B(in[500]), .Z(n995) );
  XNOR U1780 ( .A(in[1460]), .B(in[1140]), .Z(n994) );
  XNOR U1781 ( .A(n995), .B(n994), .Z(n996) );
  XNOR U1782 ( .A(in[180]), .B(n996), .Z(n1237) );
  XOR U1783 ( .A(n1559), .B(n1237), .Z(n4375) );
  XOR U1784 ( .A(in[1396]), .B(n4375), .Z(n5060) );
  NANDN U1785 ( .A(n5061), .B(n5060), .Z(n997) );
  XOR U1786 ( .A(n1664), .B(n997), .Z(out[1040]) );
  XOR U1787 ( .A(n3400), .B(in[548]), .Z(n1668) );
  XOR U1788 ( .A(in[83]), .B(in[1043]), .Z(n999) );
  XNOR U1789 ( .A(in[723]), .B(in[403]), .Z(n998) );
  XNOR U1790 ( .A(n999), .B(n998), .Z(n1000) );
  XNOR U1791 ( .A(in[1363]), .B(n1000), .Z(n1758) );
  XOR U1792 ( .A(in[852]), .B(in[1172]), .Z(n1002) );
  XNOR U1793 ( .A(in[1492]), .B(in[212]), .Z(n1001) );
  XNOR U1794 ( .A(n1002), .B(n1001), .Z(n1003) );
  XOR U1795 ( .A(in[532]), .B(n1003), .Z(n1450) );
  IV U1796 ( .A(n3216), .Z(n4010) );
  XNOR U1797 ( .A(in[148]), .B(n4010), .Z(n5064) );
  XOR U1798 ( .A(in[1332]), .B(in[52]), .Z(n1005) );
  XNOR U1799 ( .A(in[692]), .B(in[372]), .Z(n1004) );
  XNOR U1800 ( .A(n1005), .B(n1004), .Z(n1006) );
  XNOR U1801 ( .A(in[1012]), .B(n1006), .Z(n1563) );
  XOR U1802 ( .A(in[821]), .B(in[501]), .Z(n1008) );
  XNOR U1803 ( .A(in[1461]), .B(in[1141]), .Z(n1007) );
  XNOR U1804 ( .A(n1008), .B(n1007), .Z(n1009) );
  XNOR U1805 ( .A(in[181]), .B(n1009), .Z(n1252) );
  XOR U1806 ( .A(n1563), .B(n1252), .Z(n4378) );
  XOR U1807 ( .A(in[1397]), .B(n4378), .Z(n5063) );
  NANDN U1808 ( .A(n5064), .B(n5063), .Z(n1010) );
  XOR U1809 ( .A(n1668), .B(n1010), .Z(out[1041]) );
  IV U1810 ( .A(n4061), .Z(n3404) );
  XOR U1811 ( .A(n3404), .B(in[549]), .Z(n1673) );
  XOR U1812 ( .A(in[853]), .B(in[1173]), .Z(n1012) );
  XNOR U1813 ( .A(in[1493]), .B(in[213]), .Z(n1011) );
  XNOR U1814 ( .A(n1012), .B(n1011), .Z(n1013) );
  XOR U1815 ( .A(in[533]), .B(n1013), .Z(n1452) );
  IV U1816 ( .A(n2759), .Z(n4014) );
  XNOR U1817 ( .A(in[149]), .B(n4014), .Z(n5067) );
  XOR U1818 ( .A(in[822]), .B(in[502]), .Z(n1016) );
  XNOR U1819 ( .A(in[1462]), .B(in[1142]), .Z(n1015) );
  XNOR U1820 ( .A(n1016), .B(n1015), .Z(n1017) );
  XNOR U1821 ( .A(in[182]), .B(n1017), .Z(n1267) );
  XOR U1822 ( .A(in[1333]), .B(in[53]), .Z(n1019) );
  XNOR U1823 ( .A(in[693]), .B(in[373]), .Z(n1018) );
  XNOR U1824 ( .A(n1019), .B(n1018), .Z(n1020) );
  XNOR U1825 ( .A(in[1013]), .B(n1020), .Z(n1567) );
  XOR U1826 ( .A(n1267), .B(n1567), .Z(n4381) );
  XOR U1827 ( .A(in[1398]), .B(n4381), .Z(n5066) );
  NANDN U1828 ( .A(n5067), .B(n5066), .Z(n1021) );
  XOR U1829 ( .A(n1673), .B(n1021), .Z(out[1042]) );
  XOR U1830 ( .A(n1023), .B(n1022), .Z(n2038) );
  XOR U1831 ( .A(in[550]), .B(n2038), .Z(n1677) );
  XOR U1832 ( .A(in[854]), .B(in[1174]), .Z(n1025) );
  XNOR U1833 ( .A(in[1494]), .B(in[214]), .Z(n1024) );
  XNOR U1834 ( .A(n1025), .B(n1024), .Z(n1026) );
  XOR U1835 ( .A(in[534]), .B(n1026), .Z(n1454) );
  XOR U1836 ( .A(in[150]), .B(n2776), .Z(n5071) );
  XOR U1837 ( .A(in[1334]), .B(in[54]), .Z(n1029) );
  XNOR U1838 ( .A(in[694]), .B(in[374]), .Z(n1028) );
  XNOR U1839 ( .A(n1029), .B(n1028), .Z(n1030) );
  XNOR U1840 ( .A(in[1014]), .B(n1030), .Z(n1571) );
  XOR U1841 ( .A(in[823]), .B(in[503]), .Z(n1032) );
  XNOR U1842 ( .A(in[1463]), .B(in[1143]), .Z(n1031) );
  XNOR U1843 ( .A(n1032), .B(n1031), .Z(n1033) );
  XNOR U1844 ( .A(in[183]), .B(n1033), .Z(n1279) );
  XOR U1845 ( .A(n1571), .B(n1279), .Z(n4384) );
  XOR U1846 ( .A(in[1399]), .B(n4384), .Z(n5068) );
  NANDN U1847 ( .A(n5071), .B(n5068), .Z(n1034) );
  XNOR U1848 ( .A(n1677), .B(n1034), .Z(out[1043]) );
  XOR U1849 ( .A(n1036), .B(n1035), .Z(n2041) );
  XOR U1850 ( .A(in[551]), .B(n2041), .Z(n1681) );
  XOR U1851 ( .A(in[855]), .B(in[1175]), .Z(n1038) );
  XNOR U1852 ( .A(in[1495]), .B(in[215]), .Z(n1037) );
  XNOR U1853 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1854 ( .A(in[535]), .B(n1039), .Z(n1456) );
  XOR U1855 ( .A(in[151]), .B(n2783), .Z(n5078) );
  XOR U1856 ( .A(in[824]), .B(in[504]), .Z(n1042) );
  XNOR U1857 ( .A(in[1464]), .B(in[1144]), .Z(n1041) );
  XNOR U1858 ( .A(n1042), .B(n1041), .Z(n1043) );
  XNOR U1859 ( .A(in[184]), .B(n1043), .Z(n1285) );
  XOR U1860 ( .A(in[1335]), .B(in[55]), .Z(n1045) );
  XNOR U1861 ( .A(in[695]), .B(in[375]), .Z(n1044) );
  XNOR U1862 ( .A(n1045), .B(n1044), .Z(n1046) );
  XNOR U1863 ( .A(in[1015]), .B(n1046), .Z(n1575) );
  XOR U1864 ( .A(n1285), .B(n1575), .Z(n4386) );
  XOR U1865 ( .A(in[1400]), .B(n4386), .Z(n5077) );
  NANDN U1866 ( .A(n5078), .B(n5077), .Z(n1047) );
  XNOR U1867 ( .A(n1681), .B(n1047), .Z(out[1044]) );
  XOR U1868 ( .A(n1049), .B(n1048), .Z(n2045) );
  XOR U1869 ( .A(in[552]), .B(n2045), .Z(n1685) );
  XOR U1870 ( .A(in[856]), .B(in[1176]), .Z(n1051) );
  XNOR U1871 ( .A(in[1496]), .B(in[216]), .Z(n1050) );
  XNOR U1872 ( .A(n1051), .B(n1050), .Z(n1052) );
  XOR U1873 ( .A(in[536]), .B(n1052), .Z(n1460) );
  XOR U1874 ( .A(in[152]), .B(n2797), .Z(n5081) );
  XOR U1875 ( .A(in[825]), .B(in[505]), .Z(n1055) );
  XNOR U1876 ( .A(in[1465]), .B(in[1145]), .Z(n1054) );
  XNOR U1877 ( .A(n1055), .B(n1054), .Z(n1056) );
  XNOR U1878 ( .A(in[185]), .B(n1056), .Z(n1297) );
  XOR U1879 ( .A(in[1336]), .B(in[56]), .Z(n1058) );
  XNOR U1880 ( .A(in[696]), .B(in[376]), .Z(n1057) );
  XNOR U1881 ( .A(n1058), .B(n1057), .Z(n1059) );
  XNOR U1882 ( .A(in[1016]), .B(n1059), .Z(n1579) );
  XOR U1883 ( .A(n1297), .B(n1579), .Z(n4389) );
  XOR U1884 ( .A(in[1401]), .B(n4389), .Z(n5080) );
  NANDN U1885 ( .A(n5081), .B(n5080), .Z(n1060) );
  XNOR U1886 ( .A(n1685), .B(n1060), .Z(out[1045]) );
  XOR U1887 ( .A(n1062), .B(n1061), .Z(n2047) );
  XOR U1888 ( .A(in[553]), .B(n2047), .Z(n1689) );
  XOR U1889 ( .A(in[857]), .B(in[1177]), .Z(n1064) );
  XNOR U1890 ( .A(in[1497]), .B(in[217]), .Z(n1063) );
  XNOR U1891 ( .A(n1064), .B(n1063), .Z(n1065) );
  XOR U1892 ( .A(in[537]), .B(n1065), .Z(n1462) );
  XOR U1893 ( .A(in[153]), .B(n2820), .Z(n5084) );
  XOR U1894 ( .A(in[1337]), .B(in[57]), .Z(n1068) );
  XNOR U1895 ( .A(in[697]), .B(in[377]), .Z(n1067) );
  XNOR U1896 ( .A(n1068), .B(n1067), .Z(n1069) );
  XNOR U1897 ( .A(in[1017]), .B(n1069), .Z(n1583) );
  XOR U1898 ( .A(in[826]), .B(in[506]), .Z(n1071) );
  XNOR U1899 ( .A(in[1466]), .B(in[1146]), .Z(n1070) );
  XNOR U1900 ( .A(n1071), .B(n1070), .Z(n1072) );
  XNOR U1901 ( .A(in[186]), .B(n1072), .Z(n1309) );
  XOR U1902 ( .A(n1583), .B(n1309), .Z(n2114) );
  IV U1903 ( .A(n2114), .Z(n4392) );
  XNOR U1904 ( .A(in[1402]), .B(n4392), .Z(n5083) );
  NANDN U1905 ( .A(n5084), .B(n5083), .Z(n1073) );
  XNOR U1906 ( .A(n1689), .B(n1073), .Z(out[1046]) );
  XOR U1907 ( .A(n1075), .B(n1074), .Z(n2049) );
  XOR U1908 ( .A(in[554]), .B(n2049), .Z(n1693) );
  XOR U1909 ( .A(in[858]), .B(in[1178]), .Z(n1077) );
  XNOR U1910 ( .A(in[1498]), .B(in[218]), .Z(n1076) );
  XNOR U1911 ( .A(n1077), .B(n1076), .Z(n1078) );
  XOR U1912 ( .A(in[538]), .B(n1078), .Z(n1464) );
  XOR U1913 ( .A(in[154]), .B(n2843), .Z(n5087) );
  XOR U1914 ( .A(in[1338]), .B(in[58]), .Z(n1081) );
  XNOR U1915 ( .A(in[698]), .B(in[378]), .Z(n1080) );
  XNOR U1916 ( .A(n1081), .B(n1080), .Z(n1082) );
  XNOR U1917 ( .A(in[1018]), .B(n1082), .Z(n1587) );
  XOR U1918 ( .A(in[827]), .B(in[507]), .Z(n1084) );
  XNOR U1919 ( .A(in[1467]), .B(in[1147]), .Z(n1083) );
  XNOR U1920 ( .A(n1084), .B(n1083), .Z(n1085) );
  XNOR U1921 ( .A(in[187]), .B(n1085), .Z(n1313) );
  XOR U1922 ( .A(n1587), .B(n1313), .Z(n2116) );
  IV U1923 ( .A(n2116), .Z(n4395) );
  XNOR U1924 ( .A(in[1403]), .B(n4395), .Z(n5086) );
  NANDN U1925 ( .A(n5087), .B(n5086), .Z(n1086) );
  XNOR U1926 ( .A(n1693), .B(n1086), .Z(out[1047]) );
  XOR U1927 ( .A(in[1579]), .B(in[619]), .Z(n1088) );
  XNOR U1928 ( .A(in[939]), .B(in[299]), .Z(n1087) );
  XNOR U1929 ( .A(n1088), .B(n1087), .Z(n1089) );
  XNOR U1930 ( .A(in[1259]), .B(n1089), .Z(n1597) );
  XNOR U1931 ( .A(n1090), .B(n1597), .Z(n3428) );
  IV U1932 ( .A(n3428), .Z(n4090) );
  XOR U1933 ( .A(in[555]), .B(n4090), .Z(n1697) );
  XOR U1934 ( .A(in[859]), .B(in[1179]), .Z(n1092) );
  XNOR U1935 ( .A(in[1499]), .B(in[219]), .Z(n1091) );
  XNOR U1936 ( .A(n1092), .B(n1091), .Z(n1093) );
  XOR U1937 ( .A(in[539]), .B(n1093), .Z(n1468) );
  XOR U1938 ( .A(in[155]), .B(n2867), .Z(n5090) );
  XOR U1939 ( .A(in[828]), .B(in[508]), .Z(n1096) );
  XNOR U1940 ( .A(in[1468]), .B(in[1148]), .Z(n1095) );
  XNOR U1941 ( .A(n1096), .B(n1095), .Z(n1097) );
  XNOR U1942 ( .A(in[188]), .B(n1097), .Z(n1317) );
  XOR U1943 ( .A(n1098), .B(n1317), .Z(n4398) );
  XOR U1944 ( .A(in[1404]), .B(n4398), .Z(n5089) );
  NANDN U1945 ( .A(n5090), .B(n5089), .Z(n1099) );
  XNOR U1946 ( .A(n1697), .B(n1099), .Z(out[1048]) );
  XOR U1947 ( .A(in[1580]), .B(in[620]), .Z(n1101) );
  XNOR U1948 ( .A(in[940]), .B(in[300]), .Z(n1100) );
  XNOR U1949 ( .A(n1101), .B(n1100), .Z(n1102) );
  XNOR U1950 ( .A(in[1260]), .B(n1102), .Z(n1601) );
  XNOR U1951 ( .A(n1103), .B(n1601), .Z(n3431) );
  IV U1952 ( .A(n3431), .Z(n4094) );
  XOR U1953 ( .A(in[556]), .B(n4094), .Z(n1701) );
  XOR U1954 ( .A(in[860]), .B(in[1180]), .Z(n1105) );
  XNOR U1955 ( .A(in[1500]), .B(in[220]), .Z(n1104) );
  XNOR U1956 ( .A(n1105), .B(n1104), .Z(n1106) );
  XOR U1957 ( .A(in[540]), .B(n1106), .Z(n1474) );
  XOR U1958 ( .A(in[156]), .B(n2891), .Z(n5093) );
  XOR U1959 ( .A(n1109), .B(n1108), .Z(n4405) );
  XOR U1960 ( .A(in[1405]), .B(n4405), .Z(n5092) );
  NANDN U1961 ( .A(n5093), .B(n5092), .Z(n1110) );
  XNOR U1962 ( .A(n1701), .B(n1110), .Z(out[1049]) );
  XOR U1963 ( .A(in[1343]), .B(in[63]), .Z(n1112) );
  XNOR U1964 ( .A(in[703]), .B(in[383]), .Z(n1111) );
  XNOR U1965 ( .A(n1112), .B(n1111), .Z(n1113) );
  XNOR U1966 ( .A(in[1023]), .B(n1113), .Z(n1157) );
  XOR U1967 ( .A(n1114), .B(n1157), .Z(n3969) );
  XOR U1968 ( .A(in[639]), .B(n3969), .Z(n2715) );
  IV U1969 ( .A(n2715), .Z(n2804) );
  XNOR U1970 ( .A(in[230]), .B(n2038), .Z(n3192) );
  XOR U1971 ( .A(in[874]), .B(in[1194]), .Z(n1116) );
  XNOR U1972 ( .A(in[1514]), .B(in[234]), .Z(n1115) );
  XNOR U1973 ( .A(n1116), .B(n1115), .Z(n1117) );
  XNOR U1974 ( .A(in[554]), .B(n1117), .Z(n1525) );
  XNOR U1975 ( .A(n1118), .B(n1525), .Z(n4105) );
  IV U1976 ( .A(n4105), .Z(n1298) );
  XOR U1977 ( .A(in[1450]), .B(n1298), .Z(n3189) );
  NAND U1978 ( .A(n3192), .B(n3189), .Z(n1119) );
  XOR U1979 ( .A(n2804), .B(n1119), .Z(out[104]) );
  XOR U1980 ( .A(in[1581]), .B(in[621]), .Z(n1121) );
  XNOR U1981 ( .A(in[941]), .B(in[301]), .Z(n1120) );
  XNOR U1982 ( .A(n1121), .B(n1120), .Z(n1122) );
  XNOR U1983 ( .A(in[1261]), .B(n1122), .Z(n1605) );
  XNOR U1984 ( .A(n1123), .B(n1605), .Z(n3434) );
  IV U1985 ( .A(n3434), .Z(n4098) );
  XOR U1986 ( .A(in[557]), .B(n4098), .Z(n1705) );
  XOR U1987 ( .A(in[861]), .B(in[1181]), .Z(n1125) );
  XNOR U1988 ( .A(in[1501]), .B(in[221]), .Z(n1124) );
  XNOR U1989 ( .A(n1125), .B(n1124), .Z(n1126) );
  XOR U1990 ( .A(in[541]), .B(n1126), .Z(n1478) );
  XOR U1991 ( .A(in[157]), .B(n2924), .Z(n5096) );
  XOR U1992 ( .A(in[830]), .B(in[510]), .Z(n1129) );
  XNOR U1993 ( .A(in[1470]), .B(in[1150]), .Z(n1128) );
  XNOR U1994 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1995 ( .A(in[190]), .B(n1130), .Z(n1321) );
  XOR U1996 ( .A(n1131), .B(n1321), .Z(n4408) );
  XOR U1997 ( .A(in[1406]), .B(n4408), .Z(n5095) );
  NANDN U1998 ( .A(n5096), .B(n5095), .Z(n1132) );
  XNOR U1999 ( .A(n1705), .B(n1132), .Z(out[1050]) );
  XOR U2000 ( .A(in[1582]), .B(in[622]), .Z(n1134) );
  XNOR U2001 ( .A(in[942]), .B(in[302]), .Z(n1133) );
  XNOR U2002 ( .A(n1134), .B(n1133), .Z(n1135) );
  XNOR U2003 ( .A(in[1262]), .B(n1135), .Z(n1609) );
  XNOR U2004 ( .A(n1136), .B(n1609), .Z(n3437) );
  IV U2005 ( .A(n3437), .Z(n4102) );
  XOR U2006 ( .A(in[558]), .B(n4102), .Z(n1709) );
  XOR U2007 ( .A(in[862]), .B(in[1182]), .Z(n1138) );
  XNOR U2008 ( .A(in[1502]), .B(in[222]), .Z(n1137) );
  XNOR U2009 ( .A(n1138), .B(n1137), .Z(n1139) );
  XOR U2010 ( .A(in[542]), .B(n1139), .Z(n1482) );
  XNOR U2011 ( .A(in[158]), .B(n4054), .Z(n1458) );
  IV U2012 ( .A(n1458), .Z(n5099) );
  XOR U2013 ( .A(in[831]), .B(in[511]), .Z(n1142) );
  XNOR U2014 ( .A(in[1471]), .B(in[1151]), .Z(n1141) );
  XNOR U2015 ( .A(n1142), .B(n1141), .Z(n1143) );
  XNOR U2016 ( .A(in[191]), .B(n1143), .Z(n1325) );
  XOR U2017 ( .A(n1144), .B(n1325), .Z(n4411) );
  XOR U2018 ( .A(in[1407]), .B(n4411), .Z(n5098) );
  NANDN U2019 ( .A(n5099), .B(n5098), .Z(n1145) );
  XNOR U2020 ( .A(n1709), .B(n1145), .Z(out[1051]) );
  XOR U2021 ( .A(in[1583]), .B(in[623]), .Z(n1147) );
  XNOR U2022 ( .A(in[943]), .B(in[303]), .Z(n1146) );
  XNOR U2023 ( .A(n1147), .B(n1146), .Z(n1148) );
  XNOR U2024 ( .A(in[1263]), .B(n1148), .Z(n1613) );
  XNOR U2025 ( .A(n1149), .B(n1613), .Z(n3440) );
  IV U2026 ( .A(n3440), .Z(n4106) );
  XOR U2027 ( .A(in[559]), .B(n4106), .Z(n1714) );
  XOR U2028 ( .A(in[863]), .B(in[1183]), .Z(n1151) );
  XNOR U2029 ( .A(in[1503]), .B(in[223]), .Z(n1150) );
  XNOR U2030 ( .A(n1151), .B(n1150), .Z(n1152) );
  XOR U2031 ( .A(in[543]), .B(n1152), .Z(n1484) );
  XOR U2032 ( .A(in[159]), .B(n4058), .Z(n5103) );
  XOR U2033 ( .A(in[768]), .B(in[1088]), .Z(n1155) );
  XNOR U2034 ( .A(in[448]), .B(in[1408]), .Z(n1154) );
  XNOR U2035 ( .A(n1155), .B(n1154), .Z(n1156) );
  XNOR U2036 ( .A(in[128]), .B(n1156), .Z(n1332) );
  XOR U2037 ( .A(n1157), .B(n1332), .Z(n4414) );
  XOR U2038 ( .A(in[1344]), .B(n4414), .Z(n5100) );
  NANDN U2039 ( .A(n5103), .B(n5100), .Z(n1158) );
  XNOR U2040 ( .A(n1714), .B(n1158), .Z(out[1052]) );
  XOR U2041 ( .A(in[1584]), .B(in[624]), .Z(n1160) );
  XNOR U2042 ( .A(in[944]), .B(in[304]), .Z(n1159) );
  XNOR U2043 ( .A(n1160), .B(n1159), .Z(n1161) );
  XNOR U2044 ( .A(in[1264]), .B(n1161), .Z(n1617) );
  XNOR U2045 ( .A(n1162), .B(n1617), .Z(n3443) );
  IV U2046 ( .A(n3443), .Z(n4110) );
  XOR U2047 ( .A(in[560]), .B(n4110), .Z(n1718) );
  XOR U2048 ( .A(in[224]), .B(in[864]), .Z(n1164) );
  XNOR U2049 ( .A(in[1184]), .B(in[1504]), .Z(n1163) );
  XNOR U2050 ( .A(n1164), .B(n1163), .Z(n1165) );
  XOR U2051 ( .A(in[544]), .B(n1165), .Z(n1487) );
  XOR U2052 ( .A(in[160]), .B(n4062), .Z(n5106) );
  XOR U2053 ( .A(in[1280]), .B(in[640]), .Z(n1168) );
  XNOR U2054 ( .A(in[960]), .B(in[320]), .Z(n1167) );
  XNOR U2055 ( .A(n1168), .B(n1167), .Z(n1169) );
  XNOR U2056 ( .A(in[0]), .B(n1169), .Z(n1261) );
  XOR U2057 ( .A(in[769]), .B(in[1089]), .Z(n1171) );
  XNOR U2058 ( .A(in[449]), .B(in[1409]), .Z(n1170) );
  XNOR U2059 ( .A(n1171), .B(n1170), .Z(n1172) );
  XNOR U2060 ( .A(in[129]), .B(n1172), .Z(n1336) );
  XOR U2061 ( .A(n1261), .B(n1336), .Z(n4417) );
  XOR U2062 ( .A(in[1345]), .B(n4417), .Z(n5105) );
  NANDN U2063 ( .A(n5106), .B(n5105), .Z(n1173) );
  XNOR U2064 ( .A(n1718), .B(n1173), .Z(out[1053]) );
  XOR U2065 ( .A(in[1585]), .B(in[625]), .Z(n1175) );
  XNOR U2066 ( .A(in[945]), .B(in[305]), .Z(n1174) );
  XNOR U2067 ( .A(n1175), .B(n1174), .Z(n1176) );
  XNOR U2068 ( .A(in[1265]), .B(n1176), .Z(n1621) );
  XNOR U2069 ( .A(n1177), .B(n1621), .Z(n3446) );
  IV U2070 ( .A(n3446), .Z(n4118) );
  XOR U2071 ( .A(in[561]), .B(n4118), .Z(n1722) );
  XOR U2072 ( .A(in[225]), .B(in[865]), .Z(n1179) );
  XNOR U2073 ( .A(in[1185]), .B(in[1505]), .Z(n1178) );
  XNOR U2074 ( .A(n1179), .B(n1178), .Z(n1180) );
  XOR U2075 ( .A(in[545]), .B(n1180), .Z(n1490) );
  XNOR U2076 ( .A(in[161]), .B(n4066), .Z(n1466) );
  IV U2077 ( .A(n1466), .Z(n5113) );
  XOR U2078 ( .A(in[1]), .B(in[641]), .Z(n1183) );
  XNOR U2079 ( .A(in[961]), .B(in[321]), .Z(n1182) );
  XNOR U2080 ( .A(n1183), .B(n1182), .Z(n1184) );
  XNOR U2081 ( .A(in[1281]), .B(n1184), .Z(n1326) );
  XOR U2082 ( .A(in[1090]), .B(in[450]), .Z(n1186) );
  XNOR U2083 ( .A(in[130]), .B(in[770]), .Z(n1185) );
  XNOR U2084 ( .A(n1186), .B(n1185), .Z(n1187) );
  XNOR U2085 ( .A(in[1410]), .B(n1187), .Z(n1340) );
  XOR U2086 ( .A(n1326), .B(n1340), .Z(n4420) );
  XOR U2087 ( .A(in[1346]), .B(n4420), .Z(n5112) );
  NANDN U2088 ( .A(n5113), .B(n5112), .Z(n1188) );
  XNOR U2089 ( .A(n1722), .B(n1188), .Z(out[1054]) );
  XOR U2090 ( .A(in[1586]), .B(in[626]), .Z(n1190) );
  XNOR U2091 ( .A(in[946]), .B(in[306]), .Z(n1189) );
  XNOR U2092 ( .A(n1190), .B(n1189), .Z(n1191) );
  XNOR U2093 ( .A(in[1266]), .B(n1191), .Z(n1625) );
  XNOR U2094 ( .A(n1192), .B(n1625), .Z(n3449) );
  IV U2095 ( .A(n3449), .Z(n4122) );
  XOR U2096 ( .A(in[562]), .B(n4122), .Z(n1726) );
  XOR U2097 ( .A(in[1186]), .B(in[1506]), .Z(n1194) );
  XNOR U2098 ( .A(in[546]), .B(in[866]), .Z(n1193) );
  XNOR U2099 ( .A(n1194), .B(n1193), .Z(n1195) );
  XOR U2100 ( .A(in[226]), .B(n1195), .Z(n1493) );
  XNOR U2101 ( .A(in[162]), .B(n4074), .Z(n1470) );
  IV U2102 ( .A(n1470), .Z(n5117) );
  XOR U2103 ( .A(in[2]), .B(in[642]), .Z(n1198) );
  XNOR U2104 ( .A(in[962]), .B(in[322]), .Z(n1197) );
  XNOR U2105 ( .A(n1198), .B(n1197), .Z(n1199) );
  XNOR U2106 ( .A(in[1282]), .B(n1199), .Z(n1371) );
  XOR U2107 ( .A(in[771]), .B(in[1091]), .Z(n1201) );
  XNOR U2108 ( .A(in[451]), .B(in[1411]), .Z(n1200) );
  XNOR U2109 ( .A(n1201), .B(n1200), .Z(n1202) );
  XNOR U2110 ( .A(in[131]), .B(n1202), .Z(n1344) );
  XOR U2111 ( .A(n1371), .B(n1344), .Z(n4423) );
  XOR U2112 ( .A(in[1347]), .B(n4423), .Z(n5114) );
  NANDN U2113 ( .A(n5117), .B(n5114), .Z(n1203) );
  XNOR U2114 ( .A(n1726), .B(n1203), .Z(out[1055]) );
  XOR U2115 ( .A(in[1587]), .B(in[627]), .Z(n1205) );
  XNOR U2116 ( .A(in[947]), .B(in[307]), .Z(n1204) );
  XNOR U2117 ( .A(n1205), .B(n1204), .Z(n1206) );
  XNOR U2118 ( .A(in[1267]), .B(n1206), .Z(n1630) );
  XNOR U2119 ( .A(n1207), .B(n1630), .Z(n3452) );
  IV U2120 ( .A(n3452), .Z(n4126) );
  XOR U2121 ( .A(in[563]), .B(n4126), .Z(n1730) );
  XOR U2122 ( .A(in[1187]), .B(in[1507]), .Z(n1209) );
  XNOR U2123 ( .A(in[547]), .B(in[867]), .Z(n1208) );
  XNOR U2124 ( .A(n1209), .B(n1208), .Z(n1210) );
  XOR U2125 ( .A(in[227]), .B(n1210), .Z(n1496) );
  XNOR U2126 ( .A(in[163]), .B(n4078), .Z(n1476) );
  IV U2127 ( .A(n1476), .Z(n5121) );
  XOR U2128 ( .A(in[772]), .B(in[1092]), .Z(n1213) );
  XNOR U2129 ( .A(in[452]), .B(in[1412]), .Z(n1212) );
  XNOR U2130 ( .A(n1213), .B(n1212), .Z(n1214) );
  XNOR U2131 ( .A(in[132]), .B(n1214), .Z(n1348) );
  XOR U2132 ( .A(in[323]), .B(in[643]), .Z(n1216) );
  XNOR U2133 ( .A(in[963]), .B(in[3]), .Z(n1215) );
  XNOR U2134 ( .A(n1216), .B(n1215), .Z(n1217) );
  XNOR U2135 ( .A(in[1283]), .B(n1217), .Z(n1412) );
  XOR U2136 ( .A(n1348), .B(n1412), .Z(n4426) );
  XOR U2137 ( .A(in[1348]), .B(n4426), .Z(n5118) );
  NANDN U2138 ( .A(n5121), .B(n5118), .Z(n1218) );
  XNOR U2139 ( .A(n1730), .B(n1218), .Z(out[1056]) );
  XOR U2140 ( .A(in[1588]), .B(in[628]), .Z(n1220) );
  XNOR U2141 ( .A(in[948]), .B(in[308]), .Z(n1219) );
  XNOR U2142 ( .A(n1220), .B(n1219), .Z(n1221) );
  XNOR U2143 ( .A(in[1268]), .B(n1221), .Z(n1634) );
  XNOR U2144 ( .A(n1222), .B(n1634), .Z(n3459) );
  IV U2145 ( .A(n3459), .Z(n4130) );
  XOR U2146 ( .A(in[564]), .B(n4130), .Z(n1734) );
  XOR U2147 ( .A(in[1188]), .B(in[1508]), .Z(n1224) );
  XNOR U2148 ( .A(in[548]), .B(in[868]), .Z(n1223) );
  XNOR U2149 ( .A(n1224), .B(n1223), .Z(n1225) );
  XNOR U2150 ( .A(in[228]), .B(n1225), .Z(n1499) );
  XNOR U2151 ( .A(in[164]), .B(n4082), .Z(n1480) );
  IV U2152 ( .A(n1480), .Z(n5125) );
  XOR U2153 ( .A(in[773]), .B(in[1093]), .Z(n1228) );
  XNOR U2154 ( .A(in[453]), .B(in[1413]), .Z(n1227) );
  XNOR U2155 ( .A(n1228), .B(n1227), .Z(n1229) );
  XNOR U2156 ( .A(in[133]), .B(n1229), .Z(n1352) );
  XOR U2157 ( .A(in[324]), .B(in[644]), .Z(n1231) );
  XNOR U2158 ( .A(in[964]), .B(in[4]), .Z(n1230) );
  XNOR U2159 ( .A(n1231), .B(n1230), .Z(n1232) );
  XNOR U2160 ( .A(in[1284]), .B(n1232), .Z(n1416) );
  XOR U2161 ( .A(n1352), .B(n1416), .Z(n4429) );
  XOR U2162 ( .A(in[1349]), .B(n4429), .Z(n5122) );
  NANDN U2163 ( .A(n5125), .B(n5122), .Z(n1233) );
  XNOR U2164 ( .A(n1734), .B(n1233), .Z(out[1057]) );
  XOR U2165 ( .A(in[1589]), .B(in[629]), .Z(n1235) );
  XNOR U2166 ( .A(in[949]), .B(in[309]), .Z(n1234) );
  XNOR U2167 ( .A(n1235), .B(n1234), .Z(n1236) );
  XNOR U2168 ( .A(in[1269]), .B(n1236), .Z(n1638) );
  XNOR U2169 ( .A(n1237), .B(n1638), .Z(n3462) );
  IV U2170 ( .A(n3462), .Z(n4134) );
  XOR U2171 ( .A(in[565]), .B(n4134), .Z(n1738) );
  XOR U2172 ( .A(in[1189]), .B(in[1509]), .Z(n1239) );
  XNOR U2173 ( .A(in[549]), .B(in[869]), .Z(n1238) );
  XNOR U2174 ( .A(n1239), .B(n1238), .Z(n1240) );
  XOR U2175 ( .A(in[229]), .B(n1240), .Z(n1503) );
  XOR U2176 ( .A(in[165]), .B(n2217), .Z(n5129) );
  XOR U2177 ( .A(in[774]), .B(in[1094]), .Z(n1243) );
  XNOR U2178 ( .A(in[454]), .B(in[1414]), .Z(n1242) );
  XNOR U2179 ( .A(n1243), .B(n1242), .Z(n1244) );
  XNOR U2180 ( .A(in[134]), .B(n1244), .Z(n1356) );
  XOR U2181 ( .A(in[325]), .B(in[645]), .Z(n1246) );
  XNOR U2182 ( .A(in[965]), .B(in[5]), .Z(n1245) );
  XNOR U2183 ( .A(n1246), .B(n1245), .Z(n1247) );
  XNOR U2184 ( .A(in[1285]), .B(n1247), .Z(n1418) );
  XOR U2185 ( .A(n1356), .B(n1418), .Z(n2130) );
  IV U2186 ( .A(n2130), .Z(n4432) );
  XNOR U2187 ( .A(in[1350]), .B(n4432), .Z(n5126) );
  NANDN U2188 ( .A(n5129), .B(n5126), .Z(n1248) );
  XNOR U2189 ( .A(n1738), .B(n1248), .Z(out[1058]) );
  XOR U2190 ( .A(in[1590]), .B(in[630]), .Z(n1250) );
  XNOR U2191 ( .A(in[950]), .B(in[310]), .Z(n1249) );
  XNOR U2192 ( .A(n1250), .B(n1249), .Z(n1251) );
  XNOR U2193 ( .A(in[1270]), .B(n1251), .Z(n1642) );
  XNOR U2194 ( .A(n1252), .B(n1642), .Z(n3259) );
  IV U2195 ( .A(n3259), .Z(n4138) );
  XOR U2196 ( .A(in[566]), .B(n4138), .Z(n1742) );
  XNOR U2197 ( .A(in[166]), .B(n1253), .Z(n5133) );
  XOR U2198 ( .A(in[775]), .B(in[1095]), .Z(n1255) );
  XNOR U2199 ( .A(in[455]), .B(in[1415]), .Z(n1254) );
  XNOR U2200 ( .A(n1255), .B(n1254), .Z(n1256) );
  XNOR U2201 ( .A(in[135]), .B(n1256), .Z(n1360) );
  XOR U2202 ( .A(in[326]), .B(in[6]), .Z(n1258) );
  XNOR U2203 ( .A(in[966]), .B(in[646]), .Z(n1257) );
  XNOR U2204 ( .A(n1258), .B(n1257), .Z(n1259) );
  XNOR U2205 ( .A(in[1286]), .B(n1259), .Z(n1420) );
  XOR U2206 ( .A(n1360), .B(n1420), .Z(n4443) );
  XOR U2207 ( .A(in[1351]), .B(n4443), .Z(n5130) );
  NAND U2208 ( .A(n5133), .B(n5130), .Z(n1260) );
  XNOR U2209 ( .A(n1742), .B(n1260), .Z(out[1059]) );
  XOR U2210 ( .A(n1262), .B(n1261), .Z(n3973) );
  XOR U2211 ( .A(in[576]), .B(n3973), .Z(n2717) );
  IV U2212 ( .A(n2717), .Z(n2806) );
  XNOR U2213 ( .A(in[1451]), .B(n4109), .Z(n3220) );
  XNOR U2214 ( .A(in[231]), .B(n2041), .Z(n3222) );
  NANDN U2215 ( .A(n3220), .B(n3222), .Z(n1263) );
  XOR U2216 ( .A(n2806), .B(n1263), .Z(out[105]) );
  XOR U2217 ( .A(in[1591]), .B(in[631]), .Z(n1265) );
  XNOR U2218 ( .A(in[951]), .B(in[311]), .Z(n1264) );
  XNOR U2219 ( .A(n1265), .B(n1264), .Z(n1266) );
  XNOR U2220 ( .A(in[1271]), .B(n1266), .Z(n1646) );
  XNOR U2221 ( .A(n1267), .B(n1646), .Z(n3262) );
  IV U2222 ( .A(n3262), .Z(n4142) );
  XOR U2223 ( .A(in[567]), .B(n4142), .Z(n1746) );
  XNOR U2224 ( .A(in[167]), .B(n1268), .Z(n5137) );
  XOR U2225 ( .A(in[776]), .B(in[1096]), .Z(n1270) );
  XNOR U2226 ( .A(in[456]), .B(in[1416]), .Z(n1269) );
  XNOR U2227 ( .A(n1270), .B(n1269), .Z(n1271) );
  XNOR U2228 ( .A(in[136]), .B(n1271), .Z(n1364) );
  XOR U2229 ( .A(in[327]), .B(in[7]), .Z(n1273) );
  XNOR U2230 ( .A(in[967]), .B(in[647]), .Z(n1272) );
  XNOR U2231 ( .A(n1273), .B(n1272), .Z(n1274) );
  XNOR U2232 ( .A(in[1287]), .B(n1274), .Z(n1422) );
  XOR U2233 ( .A(n1364), .B(n1422), .Z(n4446) );
  XOR U2234 ( .A(in[1352]), .B(n4446), .Z(n5134) );
  NAND U2235 ( .A(n5137), .B(n5134), .Z(n1275) );
  XNOR U2236 ( .A(n1746), .B(n1275), .Z(out[1060]) );
  XOR U2237 ( .A(in[632]), .B(in[1592]), .Z(n1277) );
  XNOR U2238 ( .A(in[1272]), .B(in[312]), .Z(n1276) );
  XNOR U2239 ( .A(n1277), .B(n1276), .Z(n1278) );
  XNOR U2240 ( .A(in[952]), .B(n1278), .Z(n1650) );
  XNOR U2241 ( .A(n1279), .B(n1650), .Z(n3269) );
  IV U2242 ( .A(n3269), .Z(n4146) );
  XOR U2243 ( .A(in[568]), .B(n4146), .Z(n1750) );
  XNOR U2244 ( .A(in[168]), .B(n1280), .Z(n5140) );
  XOR U2245 ( .A(in[1353]), .B(n4449), .Z(n5139) );
  NAND U2246 ( .A(n5140), .B(n5139), .Z(n1281) );
  XNOR U2247 ( .A(n1750), .B(n1281), .Z(out[1061]) );
  XOR U2248 ( .A(in[633]), .B(in[1593]), .Z(n1283) );
  XNOR U2249 ( .A(in[1273]), .B(in[313]), .Z(n1282) );
  XNOR U2250 ( .A(n1283), .B(n1282), .Z(n1284) );
  XNOR U2251 ( .A(in[953]), .B(n1284), .Z(n1654) );
  XNOR U2252 ( .A(n1285), .B(n1654), .Z(n3272) );
  IV U2253 ( .A(n3272), .Z(n4150) );
  XOR U2254 ( .A(in[569]), .B(n4150), .Z(n1755) );
  XOR U2255 ( .A(in[778]), .B(in[1098]), .Z(n1287) );
  XNOR U2256 ( .A(in[458]), .B(in[1418]), .Z(n1286) );
  XNOR U2257 ( .A(n1287), .B(n1286), .Z(n1288) );
  XNOR U2258 ( .A(in[138]), .B(n1288), .Z(n1378) );
  XOR U2259 ( .A(in[329]), .B(in[969]), .Z(n1290) );
  XNOR U2260 ( .A(in[9]), .B(in[649]), .Z(n1289) );
  XNOR U2261 ( .A(n1290), .B(n1289), .Z(n1291) );
  XNOR U2262 ( .A(in[1289]), .B(n1291), .Z(n1429) );
  XOR U2263 ( .A(n1378), .B(n1429), .Z(n4452) );
  XNOR U2264 ( .A(in[1354]), .B(n4452), .Z(n5142) );
  XNOR U2265 ( .A(in[169]), .B(n1292), .Z(n5144) );
  NANDN U2266 ( .A(n5142), .B(n5144), .Z(n1293) );
  XNOR U2267 ( .A(n1755), .B(n1293), .Z(out[1062]) );
  XOR U2268 ( .A(in[634]), .B(in[1594]), .Z(n1295) );
  XNOR U2269 ( .A(in[1274]), .B(in[314]), .Z(n1294) );
  XNOR U2270 ( .A(n1295), .B(n1294), .Z(n1296) );
  XNOR U2271 ( .A(in[954]), .B(n1296), .Z(n1658) );
  XNOR U2272 ( .A(n1297), .B(n1658), .Z(n3275) );
  IV U2273 ( .A(n3275), .Z(n4154) );
  XOR U2274 ( .A(in[570]), .B(n4154), .Z(n1759) );
  XNOR U2275 ( .A(in[170]), .B(n1298), .Z(n5148) );
  XOR U2276 ( .A(in[1419]), .B(in[779]), .Z(n1300) );
  XNOR U2277 ( .A(in[1099]), .B(in[459]), .Z(n1299) );
  XNOR U2278 ( .A(n1300), .B(n1299), .Z(n1301) );
  XNOR U2279 ( .A(in[139]), .B(n1301), .Z(n1384) );
  XOR U2280 ( .A(in[1290]), .B(in[650]), .Z(n1303) );
  XNOR U2281 ( .A(in[970]), .B(in[330]), .Z(n1302) );
  XNOR U2282 ( .A(n1303), .B(n1302), .Z(n1304) );
  XNOR U2283 ( .A(in[10]), .B(n1304), .Z(n1431) );
  XOR U2284 ( .A(n1384), .B(n1431), .Z(n4455) );
  XOR U2285 ( .A(in[1355]), .B(n4455), .Z(n5145) );
  NAND U2286 ( .A(n5148), .B(n5145), .Z(n1305) );
  XNOR U2287 ( .A(n1759), .B(n1305), .Z(out[1063]) );
  XOR U2288 ( .A(in[955]), .B(in[1275]), .Z(n1307) );
  XNOR U2289 ( .A(in[1595]), .B(in[315]), .Z(n1306) );
  XNOR U2290 ( .A(n1307), .B(n1306), .Z(n1308) );
  XOR U2291 ( .A(in[635]), .B(n1308), .Z(n1662) );
  XOR U2292 ( .A(n1309), .B(n1662), .Z(n4164) );
  XOR U2293 ( .A(in[571]), .B(n4164), .Z(n1761) );
  XOR U2294 ( .A(in[956]), .B(in[1276]), .Z(n1311) );
  XNOR U2295 ( .A(in[1596]), .B(in[316]), .Z(n1310) );
  XNOR U2296 ( .A(n1311), .B(n1310), .Z(n1312) );
  XOR U2297 ( .A(in[636]), .B(n1312), .Z(n1666) );
  XOR U2298 ( .A(n1313), .B(n1666), .Z(n4168) );
  XOR U2299 ( .A(in[572]), .B(n4168), .Z(n1763) );
  XOR U2300 ( .A(in[957]), .B(in[1277]), .Z(n1315) );
  XNOR U2301 ( .A(in[1597]), .B(in[317]), .Z(n1314) );
  XNOR U2302 ( .A(n1315), .B(n1314), .Z(n1316) );
  XOR U2303 ( .A(in[637]), .B(n1316), .Z(n1671) );
  XOR U2304 ( .A(n1317), .B(n1671), .Z(n4172) );
  XOR U2305 ( .A(in[573]), .B(n4172), .Z(n1765) );
  IV U2306 ( .A(n3287), .Z(n4176) );
  XOR U2307 ( .A(in[574]), .B(n4176), .Z(n1767) );
  XOR U2308 ( .A(in[959]), .B(in[1279]), .Z(n1319) );
  XNOR U2309 ( .A(in[1599]), .B(in[319]), .Z(n1318) );
  XNOR U2310 ( .A(n1319), .B(n1318), .Z(n1320) );
  XOR U2311 ( .A(in[639]), .B(n1320), .Z(n1679) );
  XOR U2312 ( .A(n1321), .B(n1679), .Z(n3290) );
  XOR U2313 ( .A(in[575]), .B(n3290), .Z(n1768) );
  XOR U2314 ( .A(in[896]), .B(in[1216]), .Z(n1323) );
  XNOR U2315 ( .A(in[1536]), .B(in[256]), .Z(n1322) );
  XNOR U2316 ( .A(n1323), .B(n1322), .Z(n1324) );
  XOR U2317 ( .A(in[576]), .B(n1324), .Z(n1683) );
  XOR U2318 ( .A(n1325), .B(n1683), .Z(n3293) );
  XOR U2319 ( .A(in[512]), .B(n3293), .Z(n1770) );
  XOR U2320 ( .A(n1327), .B(n1326), .Z(n3977) );
  XOR U2321 ( .A(in[577]), .B(n3977), .Z(n2720) );
  IV U2322 ( .A(n2720), .Z(n2808) );
  XNOR U2323 ( .A(in[1452]), .B(n4117), .Z(n3244) );
  XNOR U2324 ( .A(in[232]), .B(n2045), .Z(n3246) );
  NANDN U2325 ( .A(n3244), .B(n3246), .Z(n1328) );
  XOR U2326 ( .A(n2808), .B(n1328), .Z(out[106]) );
  XOR U2327 ( .A(in[897]), .B(in[1217]), .Z(n1330) );
  XNOR U2328 ( .A(in[1537]), .B(in[257]), .Z(n1329) );
  XNOR U2329 ( .A(n1330), .B(n1329), .Z(n1331) );
  XOR U2330 ( .A(in[577]), .B(n1331), .Z(n1687) );
  XOR U2331 ( .A(n1332), .B(n1687), .Z(n3296) );
  XOR U2332 ( .A(in[513]), .B(n3296), .Z(n1772) );
  XOR U2333 ( .A(in[1538]), .B(in[578]), .Z(n1334) );
  XNOR U2334 ( .A(in[898]), .B(in[258]), .Z(n1333) );
  XNOR U2335 ( .A(n1334), .B(n1333), .Z(n1335) );
  XOR U2336 ( .A(in[1218]), .B(n1335), .Z(n1691) );
  XOR U2337 ( .A(n1336), .B(n1691), .Z(n3303) );
  XOR U2338 ( .A(in[514]), .B(n3303), .Z(n1774) );
  XOR U2339 ( .A(in[1539]), .B(in[579]), .Z(n1338) );
  XNOR U2340 ( .A(in[899]), .B(in[259]), .Z(n1337) );
  XNOR U2341 ( .A(n1338), .B(n1337), .Z(n1339) );
  XOR U2342 ( .A(in[1219]), .B(n1339), .Z(n1695) );
  XOR U2343 ( .A(n1340), .B(n1695), .Z(n3306) );
  XOR U2344 ( .A(in[515]), .B(n3306), .Z(n1778) );
  XOR U2345 ( .A(in[1540]), .B(in[580]), .Z(n1342) );
  XNOR U2346 ( .A(in[900]), .B(in[260]), .Z(n1341) );
  XNOR U2347 ( .A(n1342), .B(n1341), .Z(n1343) );
  XOR U2348 ( .A(in[1220]), .B(n1343), .Z(n1699) );
  XOR U2349 ( .A(n1344), .B(n1699), .Z(n3309) );
  XOR U2350 ( .A(in[516]), .B(n3309), .Z(n1780) );
  XOR U2351 ( .A(in[1541]), .B(in[581]), .Z(n1346) );
  XNOR U2352 ( .A(in[901]), .B(in[261]), .Z(n1345) );
  XNOR U2353 ( .A(n1346), .B(n1345), .Z(n1347) );
  XOR U2354 ( .A(in[1221]), .B(n1347), .Z(n1703) );
  XOR U2355 ( .A(n1348), .B(n1703), .Z(n3312) );
  XOR U2356 ( .A(in[517]), .B(n3312), .Z(n1782) );
  XOR U2357 ( .A(in[1542]), .B(in[582]), .Z(n1350) );
  XNOR U2358 ( .A(in[902]), .B(in[262]), .Z(n1349) );
  XNOR U2359 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U2360 ( .A(in[1222]), .B(n1351), .Z(n1707) );
  XOR U2361 ( .A(n1352), .B(n1707), .Z(n3315) );
  XOR U2362 ( .A(in[518]), .B(n3315), .Z(n1784) );
  XOR U2363 ( .A(in[1543]), .B(in[583]), .Z(n1354) );
  XNOR U2364 ( .A(in[903]), .B(in[263]), .Z(n1353) );
  XNOR U2365 ( .A(n1354), .B(n1353), .Z(n1355) );
  XOR U2366 ( .A(in[1223]), .B(n1355), .Z(n1712) );
  IV U2367 ( .A(n3931), .Z(n3318) );
  XOR U2368 ( .A(in[519]), .B(n3318), .Z(n1786) );
  XOR U2369 ( .A(in[1544]), .B(in[584]), .Z(n1358) );
  XNOR U2370 ( .A(in[904]), .B(in[264]), .Z(n1357) );
  XNOR U2371 ( .A(n1358), .B(n1357), .Z(n1359) );
  XOR U2372 ( .A(in[1224]), .B(n1359), .Z(n1716) );
  XOR U2373 ( .A(n1360), .B(n1716), .Z(n3935) );
  XOR U2374 ( .A(in[520]), .B(n3935), .Z(n1788) );
  XOR U2375 ( .A(in[1545]), .B(in[585]), .Z(n1362) );
  XNOR U2376 ( .A(in[905]), .B(in[265]), .Z(n1361) );
  XNOR U2377 ( .A(n1362), .B(n1361), .Z(n1363) );
  XOR U2378 ( .A(in[1225]), .B(n1363), .Z(n1720) );
  XOR U2379 ( .A(n1364), .B(n1720), .Z(n3942) );
  XOR U2380 ( .A(in[521]), .B(n3942), .Z(n1790) );
  XOR U2381 ( .A(in[1546]), .B(in[586]), .Z(n1366) );
  XNOR U2382 ( .A(in[906]), .B(in[266]), .Z(n1365) );
  XNOR U2383 ( .A(n1366), .B(n1365), .Z(n1367) );
  XOR U2384 ( .A(in[1226]), .B(n1367), .Z(n1724) );
  XOR U2385 ( .A(n1368), .B(n1724), .Z(n3946) );
  XOR U2386 ( .A(in[522]), .B(n3946), .Z(n1792) );
  NOR U2387 ( .A(n1369), .B(n1565), .Z(n1370) );
  XNOR U2388 ( .A(n1792), .B(n1370), .Z(out[1079]) );
  XOR U2389 ( .A(n1372), .B(n1371), .Z(n3984) );
  XOR U2390 ( .A(in[578]), .B(n3984), .Z(n2722) );
  IV U2391 ( .A(n2722), .Z(n2810) );
  IV U2392 ( .A(n1373), .Z(n4121) );
  XOR U2393 ( .A(in[1453]), .B(n4121), .Z(n3256) );
  XNOR U2394 ( .A(in[233]), .B(n2047), .Z(n3258) );
  NANDN U2395 ( .A(n3256), .B(n3258), .Z(n1374) );
  XOR U2396 ( .A(n2810), .B(n1374), .Z(out[107]) );
  XOR U2397 ( .A(in[1547]), .B(in[587]), .Z(n1376) );
  XNOR U2398 ( .A(in[907]), .B(in[267]), .Z(n1375) );
  XNOR U2399 ( .A(n1376), .B(n1375), .Z(n1377) );
  XOR U2400 ( .A(in[1227]), .B(n1377), .Z(n1728) );
  XOR U2401 ( .A(n1378), .B(n1728), .Z(n3950) );
  XOR U2402 ( .A(in[523]), .B(n3950), .Z(n1794) );
  NOR U2403 ( .A(n1379), .B(n1569), .Z(n1380) );
  XNOR U2404 ( .A(n1794), .B(n1380), .Z(out[1080]) );
  XOR U2405 ( .A(in[1548]), .B(in[588]), .Z(n1382) );
  XNOR U2406 ( .A(in[908]), .B(in[268]), .Z(n1381) );
  XNOR U2407 ( .A(n1382), .B(n1381), .Z(n1383) );
  XOR U2408 ( .A(in[1228]), .B(n1383), .Z(n1732) );
  XOR U2409 ( .A(n1384), .B(n1732), .Z(n3954) );
  XOR U2410 ( .A(in[524]), .B(n3954), .Z(n1796) );
  NOR U2411 ( .A(n1385), .B(n1573), .Z(n1386) );
  XNOR U2412 ( .A(n1796), .B(n1386), .Z(out[1081]) );
  XOR U2413 ( .A(in[1549]), .B(in[589]), .Z(n1388) );
  XNOR U2414 ( .A(in[909]), .B(in[269]), .Z(n1387) );
  XNOR U2415 ( .A(n1388), .B(n1387), .Z(n1389) );
  XOR U2416 ( .A(in[1229]), .B(n1389), .Z(n1736) );
  XOR U2417 ( .A(n1390), .B(n1736), .Z(n3958) );
  XOR U2418 ( .A(in[525]), .B(n3958), .Z(n1800) );
  XOR U2419 ( .A(in[1550]), .B(in[590]), .Z(n1392) );
  XNOR U2420 ( .A(in[910]), .B(in[270]), .Z(n1391) );
  XNOR U2421 ( .A(n1392), .B(n1391), .Z(n1393) );
  XNOR U2422 ( .A(in[1230]), .B(n1393), .Z(n1740) );
  XOR U2423 ( .A(n1740), .B(n1394), .Z(n3962) );
  XOR U2424 ( .A(in[526]), .B(n3962), .Z(n1802) );
  XOR U2425 ( .A(in[1551]), .B(in[591]), .Z(n1396) );
  XNOR U2426 ( .A(in[911]), .B(in[271]), .Z(n1395) );
  XNOR U2427 ( .A(n1396), .B(n1395), .Z(n1397) );
  XOR U2428 ( .A(in[1231]), .B(n1397), .Z(n1744) );
  XOR U2429 ( .A(n1398), .B(n1744), .Z(n3966) );
  XOR U2430 ( .A(in[527]), .B(n3966), .Z(n1804) );
  XOR U2431 ( .A(in[1552]), .B(in[592]), .Z(n1400) );
  XNOR U2432 ( .A(in[912]), .B(in[272]), .Z(n1399) );
  XNOR U2433 ( .A(n1400), .B(n1399), .Z(n1401) );
  XOR U2434 ( .A(in[1232]), .B(n1401), .Z(n1748) );
  XOR U2435 ( .A(n1402), .B(n1748), .Z(n3970) );
  XOR U2436 ( .A(in[528]), .B(n3970), .Z(n1806) );
  XOR U2437 ( .A(in[1553]), .B(in[593]), .Z(n1404) );
  XNOR U2438 ( .A(in[913]), .B(in[273]), .Z(n1403) );
  XNOR U2439 ( .A(n1404), .B(n1403), .Z(n1405) );
  XOR U2440 ( .A(in[1233]), .B(n1405), .Z(n1753) );
  XOR U2441 ( .A(n1406), .B(n1753), .Z(n3974) );
  XOR U2442 ( .A(in[529]), .B(n3974), .Z(n1808) );
  XOR U2443 ( .A(in[1554]), .B(in[594]), .Z(n1408) );
  XNOR U2444 ( .A(in[914]), .B(in[274]), .Z(n1407) );
  XNOR U2445 ( .A(n1408), .B(n1407), .Z(n1409) );
  XOR U2446 ( .A(in[1234]), .B(n1409), .Z(n1757) );
  XOR U2447 ( .A(n1410), .B(n1757), .Z(n3978) );
  XOR U2448 ( .A(in[530]), .B(n3978), .Z(n1810) );
  XNOR U2449 ( .A(in[957]), .B(n3961), .Z(n1813) );
  XNOR U2450 ( .A(in[958]), .B(n3965), .Z(n1816) );
  XNOR U2451 ( .A(n1412), .B(n1411), .Z(n3988) );
  XOR U2452 ( .A(in[579]), .B(n3988), .Z(n2724) );
  IV U2453 ( .A(n2724), .Z(n2812) );
  IV U2454 ( .A(n1413), .Z(n4125) );
  XOR U2455 ( .A(in[1454]), .B(n4125), .Z(n3266) );
  XNOR U2456 ( .A(in[234]), .B(n2049), .Z(n3268) );
  NANDN U2457 ( .A(n3266), .B(n3268), .Z(n1414) );
  XOR U2458 ( .A(n2812), .B(n1414), .Z(out[108]) );
  XNOR U2459 ( .A(in[959]), .B(n3969), .Z(n1819) );
  XNOR U2460 ( .A(in[896]), .B(n3973), .Z(n1822) );
  XNOR U2461 ( .A(in[897]), .B(n3977), .Z(n1827) );
  XNOR U2462 ( .A(in[898]), .B(n3984), .Z(n1830) );
  XNOR U2463 ( .A(in[899]), .B(n3988), .Z(n1832) );
  XOR U2464 ( .A(n1416), .B(n1415), .Z(n2013) );
  XOR U2465 ( .A(in[900]), .B(n2013), .Z(n1833) );
  XOR U2466 ( .A(n1418), .B(n1417), .Z(n2016) );
  XOR U2467 ( .A(in[901]), .B(n2016), .Z(n1835) );
  XOR U2468 ( .A(n1420), .B(n1419), .Z(n2018) );
  XOR U2469 ( .A(in[902]), .B(n2018), .Z(n1837) );
  XOR U2470 ( .A(n1422), .B(n1421), .Z(n2020) );
  XOR U2471 ( .A(in[903]), .B(n2020), .Z(n1839) );
  XOR U2472 ( .A(n1424), .B(n1423), .Z(n2022) );
  XOR U2473 ( .A(in[904]), .B(n2022), .Z(n1841) );
  IV U2474 ( .A(n2013), .Z(n3992) );
  XOR U2475 ( .A(in[580]), .B(n3992), .Z(n2814) );
  IV U2476 ( .A(n1425), .Z(n4129) );
  XOR U2477 ( .A(in[1455]), .B(n4129), .Z(n3300) );
  XNOR U2478 ( .A(in[235]), .B(n4090), .Z(n3302) );
  NANDN U2479 ( .A(n3300), .B(n3302), .Z(n1426) );
  XNOR U2480 ( .A(n2814), .B(n1426), .Z(out[109]) );
  XNOR U2481 ( .A(in[200]), .B(n3935), .Z(n4280) );
  XOR U2482 ( .A(in[1420]), .B(n3194), .Z(n4281) );
  XNOR U2483 ( .A(n4483), .B(in[1043]), .Z(n2882) );
  NANDN U2484 ( .A(n4281), .B(n2882), .Z(n1427) );
  XNOR U2485 ( .A(n4280), .B(n1427), .Z(out[10]) );
  XOR U2486 ( .A(n1429), .B(n1428), .Z(n2024) );
  XOR U2487 ( .A(in[905]), .B(n2024), .Z(n1843) );
  XOR U2488 ( .A(n1431), .B(n1430), .Z(n2027) );
  XOR U2489 ( .A(in[906]), .B(n2027), .Z(n1845) );
  XOR U2490 ( .A(n1432), .B(n234), .Z(n4020) );
  XOR U2491 ( .A(in[907]), .B(n4020), .Z(n1849) );
  XOR U2492 ( .A(n1434), .B(n1433), .Z(n2030) );
  XOR U2493 ( .A(in[908]), .B(n2030), .Z(n1851) );
  XOR U2494 ( .A(n1435), .B(n235), .Z(n4032) );
  XOR U2495 ( .A(in[909]), .B(n4032), .Z(n1853) );
  XNOR U2496 ( .A(n1437), .B(n1436), .Z(n3118) );
  XOR U2497 ( .A(in[910]), .B(n3118), .Z(n1855) );
  XOR U2498 ( .A(n1438), .B(n236), .Z(n4040) );
  XOR U2499 ( .A(in[911]), .B(n4040), .Z(n1857) );
  XOR U2500 ( .A(n1439), .B(n237), .Z(n4044) );
  XOR U2501 ( .A(in[912]), .B(n4044), .Z(n1859) );
  XOR U2502 ( .A(n1441), .B(n1440), .Z(n2036) );
  XOR U2503 ( .A(in[913]), .B(n2036), .Z(n1861) );
  XOR U2504 ( .A(n1443), .B(n1442), .Z(n2039) );
  XOR U2505 ( .A(in[914]), .B(n2039), .Z(n1863) );
  IV U2506 ( .A(n2016), .Z(n3996) );
  XOR U2507 ( .A(in[581]), .B(n3996), .Z(n2816) );
  IV U2508 ( .A(n1444), .Z(n4133) );
  XOR U2509 ( .A(in[1456]), .B(n4133), .Z(n3330) );
  XNOR U2510 ( .A(in[236]), .B(n4094), .Z(n3332) );
  NANDN U2511 ( .A(n3330), .B(n3332), .Z(n1445) );
  XNOR U2512 ( .A(n2816), .B(n1445), .Z(out[110]) );
  XNOR U2513 ( .A(n1447), .B(n1446), .Z(n3124) );
  XOR U2514 ( .A(in[915]), .B(n3124), .Z(n1865) );
  XOR U2515 ( .A(n1449), .B(n1448), .Z(n3126) );
  XOR U2516 ( .A(in[916]), .B(n3126), .Z(n1867) );
  XOR U2517 ( .A(n1451), .B(n1450), .Z(n3128) );
  XOR U2518 ( .A(in[917]), .B(n3128), .Z(n1871) );
  XNOR U2519 ( .A(n1453), .B(n1452), .Z(n3130) );
  XOR U2520 ( .A(in[918]), .B(n3130), .Z(n1873) );
  XNOR U2521 ( .A(n1455), .B(n1454), .Z(n3132) );
  XOR U2522 ( .A(in[919]), .B(n3132), .Z(n1875) );
  XOR U2523 ( .A(n1457), .B(n1456), .Z(n3138) );
  XOR U2524 ( .A(in[920]), .B(n3138), .Z(n1877) );
  NOR U2525 ( .A(n1458), .B(n1709), .Z(n1459) );
  XNOR U2526 ( .A(n1877), .B(n1459), .Z(out[1115]) );
  XOR U2527 ( .A(n1461), .B(n1460), .Z(n3140) );
  XOR U2528 ( .A(in[921]), .B(n3140), .Z(n1879) );
  XNOR U2529 ( .A(n1463), .B(n1462), .Z(n3143) );
  XOR U2530 ( .A(in[922]), .B(n3143), .Z(n1881) );
  XNOR U2531 ( .A(n1465), .B(n1464), .Z(n3145) );
  XOR U2532 ( .A(in[923]), .B(n3145), .Z(n1883) );
  NOR U2533 ( .A(n1466), .B(n1722), .Z(n1467) );
  XNOR U2534 ( .A(n1883), .B(n1467), .Z(out[1118]) );
  XNOR U2535 ( .A(n1469), .B(n1468), .Z(n3024) );
  XOR U2536 ( .A(in[924]), .B(n3024), .Z(n1885) );
  NOR U2537 ( .A(n1470), .B(n1726), .Z(n1471) );
  XNOR U2538 ( .A(n1885), .B(n1471), .Z(out[1119]) );
  IV U2539 ( .A(n2018), .Z(n4000) );
  XOR U2540 ( .A(in[582]), .B(n4000), .Z(n2818) );
  IV U2541 ( .A(n1472), .Z(n4137) );
  XOR U2542 ( .A(in[1457]), .B(n4137), .Z(n3358) );
  XNOR U2543 ( .A(in[237]), .B(n4098), .Z(n3360) );
  NANDN U2544 ( .A(n3358), .B(n3360), .Z(n1473) );
  XNOR U2545 ( .A(n2818), .B(n1473), .Z(out[111]) );
  XNOR U2546 ( .A(n1475), .B(n1474), .Z(n3026) );
  XOR U2547 ( .A(in[925]), .B(n3026), .Z(n1887) );
  NOR U2548 ( .A(n1476), .B(n1730), .Z(n1477) );
  XNOR U2549 ( .A(n1887), .B(n1477), .Z(out[1120]) );
  XNOR U2550 ( .A(n1479), .B(n1478), .Z(n3028) );
  XOR U2551 ( .A(in[926]), .B(n3028), .Z(n1889) );
  NOR U2552 ( .A(n1480), .B(n1734), .Z(n1481) );
  XNOR U2553 ( .A(n1889), .B(n1481), .Z(out[1121]) );
  XNOR U2554 ( .A(n1483), .B(n1482), .Z(n3030) );
  XOR U2555 ( .A(in[927]), .B(n3030), .Z(n1893) );
  XNOR U2556 ( .A(n1485), .B(n1484), .Z(n3032) );
  XOR U2557 ( .A(in[928]), .B(n3032), .Z(n1895) );
  NOR U2558 ( .A(n5133), .B(n1742), .Z(n1486) );
  XNOR U2559 ( .A(n1895), .B(n1486), .Z(out[1123]) );
  XOR U2560 ( .A(n1488), .B(n1487), .Z(n3034) );
  XOR U2561 ( .A(in[929]), .B(n3034), .Z(n1897) );
  NOR U2562 ( .A(n5137), .B(n1746), .Z(n1489) );
  XNOR U2563 ( .A(n1897), .B(n1489), .Z(out[1124]) );
  XOR U2564 ( .A(n1491), .B(n1490), .Z(n2170) );
  XOR U2565 ( .A(in[930]), .B(n2170), .Z(n1899) );
  NOR U2566 ( .A(n5140), .B(n1750), .Z(n1492) );
  XNOR U2567 ( .A(n1899), .B(n1492), .Z(out[1125]) );
  XOR U2568 ( .A(n1494), .B(n1493), .Z(n3037) );
  XOR U2569 ( .A(in[931]), .B(n3037), .Z(n1901) );
  NOR U2570 ( .A(n5144), .B(n1755), .Z(n1495) );
  XNOR U2571 ( .A(n1901), .B(n1495), .Z(out[1126]) );
  XOR U2572 ( .A(n1497), .B(n1496), .Z(n3039) );
  XOR U2573 ( .A(in[932]), .B(n3039), .Z(n1903) );
  NOR U2574 ( .A(n5148), .B(n1759), .Z(n1498) );
  XNOR U2575 ( .A(n1903), .B(n1498), .Z(out[1127]) );
  XOR U2576 ( .A(n1500), .B(n1499), .Z(n4136) );
  XOR U2577 ( .A(in[933]), .B(n4136), .Z(n1906) );
  NAND U2578 ( .A(n1501), .B(n1761), .Z(n1502) );
  XNOR U2579 ( .A(n1906), .B(n1502), .Z(out[1128]) );
  XNOR U2580 ( .A(n1504), .B(n1503), .Z(n4140) );
  XOR U2581 ( .A(in[934]), .B(n4140), .Z(n1910) );
  NAND U2582 ( .A(n1505), .B(n1763), .Z(n1506) );
  XNOR U2583 ( .A(n1910), .B(n1506), .Z(out[1129]) );
  IV U2584 ( .A(n2020), .Z(n4004) );
  XOR U2585 ( .A(in[583]), .B(n4004), .Z(n2823) );
  IV U2586 ( .A(n1507), .Z(n4141) );
  XOR U2587 ( .A(in[1458]), .B(n4141), .Z(n3386) );
  XNOR U2588 ( .A(in[238]), .B(n4102), .Z(n3388) );
  NANDN U2589 ( .A(n3386), .B(n3388), .Z(n1508) );
  XNOR U2590 ( .A(n2823), .B(n1508), .Z(out[112]) );
  XOR U2591 ( .A(n1510), .B(n1509), .Z(n4144) );
  XOR U2592 ( .A(in[935]), .B(n4144), .Z(n1914) );
  NAND U2593 ( .A(n1511), .B(n1765), .Z(n1512) );
  XNOR U2594 ( .A(n1914), .B(n1512), .Z(out[1130]) );
  XOR U2595 ( .A(n1514), .B(n1513), .Z(n4148) );
  XOR U2596 ( .A(in[936]), .B(n4148), .Z(n1918) );
  NANDN U2597 ( .A(n1767), .B(n1515), .Z(n1516) );
  XNOR U2598 ( .A(n1918), .B(n1516), .Z(out[1131]) );
  XOR U2599 ( .A(n1518), .B(n1517), .Z(n4152) );
  XOR U2600 ( .A(in[937]), .B(n4152), .Z(n1924) );
  NAND U2601 ( .A(n1519), .B(n1768), .Z(n1520) );
  XNOR U2602 ( .A(n1924), .B(n1520), .Z(out[1132]) );
  XOR U2603 ( .A(n1522), .B(n1521), .Z(n4162) );
  XOR U2604 ( .A(in[938]), .B(n4162), .Z(n1928) );
  NAND U2605 ( .A(n1523), .B(n1770), .Z(n1524) );
  XNOR U2606 ( .A(n1928), .B(n1524), .Z(out[1133]) );
  XOR U2607 ( .A(n1526), .B(n1525), .Z(n4166) );
  XOR U2608 ( .A(in[939]), .B(n4166), .Z(n1932) );
  NAND U2609 ( .A(n1527), .B(n1772), .Z(n1528) );
  XNOR U2610 ( .A(n1932), .B(n1528), .Z(out[1134]) );
  XOR U2611 ( .A(n1530), .B(n1529), .Z(n4170) );
  XOR U2612 ( .A(in[940]), .B(n4170), .Z(n1936) );
  NAND U2613 ( .A(n1531), .B(n1774), .Z(n1532) );
  XNOR U2614 ( .A(n1936), .B(n1532), .Z(out[1135]) );
  XOR U2615 ( .A(n1534), .B(n1533), .Z(n4174) );
  XOR U2616 ( .A(in[941]), .B(n4174), .Z(n1940) );
  NAND U2617 ( .A(n1535), .B(n1778), .Z(n1536) );
  XNOR U2618 ( .A(n1940), .B(n1536), .Z(out[1136]) );
  XOR U2619 ( .A(n1538), .B(n1537), .Z(n3898) );
  XOR U2620 ( .A(in[942]), .B(n3898), .Z(n1944) );
  NAND U2621 ( .A(n1539), .B(n1780), .Z(n1540) );
  XNOR U2622 ( .A(n1944), .B(n1540), .Z(out[1137]) );
  XOR U2623 ( .A(n1542), .B(n1541), .Z(n3902) );
  XOR U2624 ( .A(in[943]), .B(n3902), .Z(n1948) );
  NAND U2625 ( .A(n1543), .B(n1782), .Z(n1544) );
  XNOR U2626 ( .A(n1948), .B(n1544), .Z(out[1138]) );
  XOR U2627 ( .A(n1546), .B(n1545), .Z(n3906) );
  XOR U2628 ( .A(in[944]), .B(n3906), .Z(n1952) );
  NAND U2629 ( .A(n1547), .B(n1784), .Z(n1548) );
  XNOR U2630 ( .A(n1952), .B(n1548), .Z(out[1139]) );
  IV U2631 ( .A(n2022), .Z(n4008) );
  XOR U2632 ( .A(in[584]), .B(n4008), .Z(n2825) );
  IV U2633 ( .A(n1549), .Z(n4145) );
  XOR U2634 ( .A(in[1459]), .B(n4145), .Z(n3421) );
  XNOR U2635 ( .A(in[239]), .B(n4106), .Z(n3423) );
  NANDN U2636 ( .A(n3421), .B(n3423), .Z(n1550) );
  XNOR U2637 ( .A(n2825), .B(n1550), .Z(out[113]) );
  XOR U2638 ( .A(n1552), .B(n1551), .Z(n3910) );
  XOR U2639 ( .A(in[945]), .B(n3910), .Z(n1956) );
  NAND U2640 ( .A(n1553), .B(n1786), .Z(n1554) );
  XNOR U2641 ( .A(n1956), .B(n1554), .Z(out[1140]) );
  XOR U2642 ( .A(n1556), .B(n1555), .Z(n3914) );
  XOR U2643 ( .A(in[946]), .B(n3914), .Z(n1960) );
  NAND U2644 ( .A(n1557), .B(n1788), .Z(n1558) );
  XNOR U2645 ( .A(n1960), .B(n1558), .Z(out[1141]) );
  XNOR U2646 ( .A(n1560), .B(n1559), .Z(n3918) );
  IV U2647 ( .A(n3918), .Z(n2574) );
  XOR U2648 ( .A(in[947]), .B(n2574), .Z(n1966) );
  NAND U2649 ( .A(n1561), .B(n1790), .Z(n1562) );
  XNOR U2650 ( .A(n1966), .B(n1562), .Z(out[1142]) );
  XNOR U2651 ( .A(n1564), .B(n1563), .Z(n3922) );
  IV U2652 ( .A(n3922), .Z(n2616) );
  XOR U2653 ( .A(in[948]), .B(n2616), .Z(n1970) );
  NAND U2654 ( .A(n1565), .B(n1792), .Z(n1566) );
  XNOR U2655 ( .A(n1970), .B(n1566), .Z(out[1143]) );
  XNOR U2656 ( .A(n1568), .B(n1567), .Z(n3926) );
  IV U2657 ( .A(n3926), .Z(n2658) );
  XOR U2658 ( .A(in[949]), .B(n2658), .Z(n1974) );
  NAND U2659 ( .A(n1569), .B(n1794), .Z(n1570) );
  XNOR U2660 ( .A(n1974), .B(n1570), .Z(out[1144]) );
  XOR U2661 ( .A(n1572), .B(n1571), .Z(n3065) );
  XOR U2662 ( .A(in[950]), .B(n3065), .Z(n1978) );
  NAND U2663 ( .A(n1573), .B(n1796), .Z(n1574) );
  XNOR U2664 ( .A(n1978), .B(n1574), .Z(out[1145]) );
  XOR U2665 ( .A(n1576), .B(n1575), .Z(n3067) );
  XOR U2666 ( .A(in[951]), .B(n3067), .Z(n1982) );
  NAND U2667 ( .A(n1577), .B(n1800), .Z(n1578) );
  XNOR U2668 ( .A(n1982), .B(n1578), .Z(out[1146]) );
  XOR U2669 ( .A(n1580), .B(n1579), .Z(n3070) );
  XOR U2670 ( .A(in[952]), .B(n3070), .Z(n1986) );
  NAND U2671 ( .A(n1581), .B(n1802), .Z(n1582) );
  XNOR U2672 ( .A(n1986), .B(n1582), .Z(out[1147]) );
  XNOR U2673 ( .A(n1584), .B(n1583), .Z(n3945) );
  IV U2674 ( .A(n3945), .Z(n2703) );
  XOR U2675 ( .A(in[953]), .B(n2703), .Z(n1990) );
  NAND U2676 ( .A(n1585), .B(n1804), .Z(n1586) );
  XNOR U2677 ( .A(n1990), .B(n1586), .Z(out[1148]) );
  XNOR U2678 ( .A(n1588), .B(n1587), .Z(n3949) );
  IV U2679 ( .A(n3949), .Z(n2705) );
  XOR U2680 ( .A(in[954]), .B(n2705), .Z(n1994) );
  NAND U2681 ( .A(n1589), .B(n1806), .Z(n1590) );
  XNOR U2682 ( .A(n1994), .B(n1590), .Z(out[1149]) );
  IV U2683 ( .A(n2024), .Z(n4012) );
  XOR U2684 ( .A(in[585]), .B(n4012), .Z(n2827) );
  IV U2685 ( .A(n1591), .Z(n4149) );
  XOR U2686 ( .A(in[1460]), .B(n4149), .Z(n3456) );
  XNOR U2687 ( .A(in[240]), .B(n4110), .Z(n3458) );
  NANDN U2688 ( .A(n3456), .B(n3458), .Z(n1592) );
  XNOR U2689 ( .A(n2827), .B(n1592), .Z(out[114]) );
  XOR U2690 ( .A(in[955]), .B(n3953), .Z(n1998) );
  NAND U2691 ( .A(n1593), .B(n1808), .Z(n1594) );
  XNOR U2692 ( .A(n1998), .B(n1594), .Z(out[1150]) );
  XOR U2693 ( .A(in[956]), .B(n3957), .Z(n2002) );
  NANDN U2694 ( .A(n1595), .B(n1810), .Z(n1596) );
  XNOR U2695 ( .A(n2002), .B(n1596), .Z(out[1151]) );
  XOR U2696 ( .A(n1598), .B(n1597), .Z(n4296) );
  XOR U2697 ( .A(in[1004]), .B(n4296), .Z(n1812) );
  NAND U2698 ( .A(n1599), .B(n1813), .Z(n1600) );
  XNOR U2699 ( .A(n1812), .B(n1600), .Z(out[1152]) );
  XOR U2700 ( .A(n1602), .B(n1601), .Z(n4298) );
  XOR U2701 ( .A(in[1005]), .B(n4298), .Z(n1815) );
  NAND U2702 ( .A(n1603), .B(n1816), .Z(n1604) );
  XNOR U2703 ( .A(n1815), .B(n1604), .Z(out[1153]) );
  XOR U2704 ( .A(n1606), .B(n1605), .Z(n4300) );
  XOR U2705 ( .A(in[1006]), .B(n4300), .Z(n1818) );
  NAND U2706 ( .A(n1607), .B(n1819), .Z(n1608) );
  XNOR U2707 ( .A(n1818), .B(n1608), .Z(out[1154]) );
  XOR U2708 ( .A(n1610), .B(n1609), .Z(n4302) );
  XOR U2709 ( .A(in[1007]), .B(n4302), .Z(n1821) );
  NAND U2710 ( .A(n1611), .B(n1822), .Z(n1612) );
  XNOR U2711 ( .A(n1821), .B(n1612), .Z(out[1155]) );
  XOR U2712 ( .A(n1614), .B(n1613), .Z(n4309) );
  XOR U2713 ( .A(in[1008]), .B(n4309), .Z(n1826) );
  NAND U2714 ( .A(n1615), .B(n1827), .Z(n1616) );
  XNOR U2715 ( .A(n1826), .B(n1616), .Z(out[1156]) );
  XOR U2716 ( .A(n1618), .B(n1617), .Z(n4312) );
  XOR U2717 ( .A(in[1009]), .B(n4312), .Z(n1829) );
  NAND U2718 ( .A(n1619), .B(n1830), .Z(n1620) );
  XNOR U2719 ( .A(n1829), .B(n1620), .Z(out[1157]) );
  XOR U2720 ( .A(n1622), .B(n1621), .Z(n4315) );
  XOR U2721 ( .A(in[1010]), .B(n4315), .Z(n5016) );
  NAND U2722 ( .A(n1623), .B(n1832), .Z(n1624) );
  XNOR U2723 ( .A(n5016), .B(n1624), .Z(out[1158]) );
  XOR U2724 ( .A(n1626), .B(n1625), .Z(n4318) );
  XOR U2725 ( .A(in[1011]), .B(n4318), .Z(n5020) );
  NAND U2726 ( .A(n1627), .B(n1833), .Z(n1628) );
  XNOR U2727 ( .A(n5020), .B(n1628), .Z(out[1159]) );
  IV U2728 ( .A(n2027), .Z(n4016) );
  XOR U2729 ( .A(in[586]), .B(n4016), .Z(n2829) );
  XNOR U2730 ( .A(in[1461]), .B(n4153), .Z(n3478) );
  XNOR U2731 ( .A(in[241]), .B(n4118), .Z(n3480) );
  NANDN U2732 ( .A(n3478), .B(n3480), .Z(n1629) );
  XNOR U2733 ( .A(n2829), .B(n1629), .Z(out[115]) );
  XOR U2734 ( .A(n1631), .B(n1630), .Z(n4321) );
  XOR U2735 ( .A(in[1012]), .B(n4321), .Z(n5024) );
  NAND U2736 ( .A(n1632), .B(n1835), .Z(n1633) );
  XNOR U2737 ( .A(n5024), .B(n1633), .Z(out[1160]) );
  XOR U2738 ( .A(n1635), .B(n1634), .Z(n4324) );
  XOR U2739 ( .A(in[1013]), .B(n4324), .Z(n5028) );
  NAND U2740 ( .A(n1636), .B(n1837), .Z(n1637) );
  XNOR U2741 ( .A(n5028), .B(n1637), .Z(out[1161]) );
  XOR U2742 ( .A(n1639), .B(n1638), .Z(n4327) );
  XOR U2743 ( .A(in[1014]), .B(n4327), .Z(n5036) );
  NAND U2744 ( .A(n1640), .B(n1839), .Z(n1641) );
  XNOR U2745 ( .A(n5036), .B(n1641), .Z(out[1162]) );
  XOR U2746 ( .A(n1643), .B(n1642), .Z(n4330) );
  XOR U2747 ( .A(in[1015]), .B(n4330), .Z(n5040) );
  NAND U2748 ( .A(n1644), .B(n1841), .Z(n1645) );
  XNOR U2749 ( .A(n5040), .B(n1645), .Z(out[1163]) );
  XOR U2750 ( .A(n1647), .B(n1646), .Z(n4178) );
  XOR U2751 ( .A(in[1016]), .B(n4178), .Z(n5044) );
  NAND U2752 ( .A(n1648), .B(n1843), .Z(n1649) );
  XNOR U2753 ( .A(n5044), .B(n1649), .Z(out[1164]) );
  XOR U2754 ( .A(n1651), .B(n1650), .Z(n4181) );
  XOR U2755 ( .A(in[1017]), .B(n4181), .Z(n5048) );
  NAND U2756 ( .A(n1652), .B(n1845), .Z(n1653) );
  XNOR U2757 ( .A(n5048), .B(n1653), .Z(out[1165]) );
  XOR U2758 ( .A(n1655), .B(n1654), .Z(n4184) );
  XOR U2759 ( .A(in[1018]), .B(n4184), .Z(n5052) );
  NAND U2760 ( .A(n1656), .B(n1849), .Z(n1657) );
  XNOR U2761 ( .A(n5052), .B(n1657), .Z(out[1166]) );
  XOR U2762 ( .A(n1659), .B(n1658), .Z(n4187) );
  XOR U2763 ( .A(in[1019]), .B(n4187), .Z(n5056) );
  NANDN U2764 ( .A(n1660), .B(n1851), .Z(n1661) );
  XNOR U2765 ( .A(n5056), .B(n1661), .Z(out[1167]) );
  IV U2766 ( .A(n3059), .Z(n4190) );
  XOR U2767 ( .A(in[1020]), .B(n4190), .Z(n5059) );
  NANDN U2768 ( .A(n1664), .B(n1853), .Z(n1665) );
  XOR U2769 ( .A(n5059), .B(n1665), .Z(out[1168]) );
  IV U2770 ( .A(n3061), .Z(n4193) );
  XOR U2771 ( .A(in[1021]), .B(n4193), .Z(n5062) );
  NANDN U2772 ( .A(n1668), .B(n1855), .Z(n1669) );
  XOR U2773 ( .A(n5062), .B(n1669), .Z(out[1169]) );
  XNOR U2774 ( .A(in[587]), .B(n4020), .Z(n2831) );
  XNOR U2775 ( .A(in[1462]), .B(n4163), .Z(n3500) );
  XNOR U2776 ( .A(in[242]), .B(n4122), .Z(n3502) );
  NANDN U2777 ( .A(n3500), .B(n3502), .Z(n1670) );
  XNOR U2778 ( .A(n2831), .B(n1670), .Z(out[116]) );
  IV U2779 ( .A(n3063), .Z(n4198) );
  XOR U2780 ( .A(in[1022]), .B(n4198), .Z(n5065) );
  NANDN U2781 ( .A(n1673), .B(n1857), .Z(n1674) );
  XOR U2782 ( .A(n5065), .B(n1674), .Z(out[1170]) );
  XOR U2783 ( .A(n1676), .B(n1675), .Z(n4199) );
  XOR U2784 ( .A(in[1023]), .B(n4199), .Z(n5069) );
  NAND U2785 ( .A(n1677), .B(n1859), .Z(n1678) );
  XNOR U2786 ( .A(n5069), .B(n1678), .Z(out[1171]) );
  IV U2787 ( .A(n3068), .Z(n4200) );
  XOR U2788 ( .A(in[960]), .B(n4200), .Z(n5076) );
  NAND U2789 ( .A(n1681), .B(n1861), .Z(n1682) );
  XOR U2790 ( .A(n5076), .B(n1682), .Z(out[1172]) );
  IV U2791 ( .A(n3071), .Z(n4201) );
  XOR U2792 ( .A(in[961]), .B(n4201), .Z(n5079) );
  NAND U2793 ( .A(n1685), .B(n1863), .Z(n1686) );
  XOR U2794 ( .A(n5079), .B(n1686), .Z(out[1173]) );
  IV U2795 ( .A(n3073), .Z(n4202) );
  XOR U2796 ( .A(in[962]), .B(n4202), .Z(n5082) );
  NAND U2797 ( .A(n1689), .B(n1865), .Z(n1690) );
  XOR U2798 ( .A(n5082), .B(n1690), .Z(out[1174]) );
  IV U2799 ( .A(n3077), .Z(n4203) );
  XOR U2800 ( .A(in[963]), .B(n4203), .Z(n5085) );
  NAND U2801 ( .A(n1693), .B(n1867), .Z(n1694) );
  XOR U2802 ( .A(n5085), .B(n1694), .Z(out[1175]) );
  IV U2803 ( .A(n3079), .Z(n4204) );
  XOR U2804 ( .A(in[964]), .B(n4204), .Z(n5088) );
  NAND U2805 ( .A(n1697), .B(n1871), .Z(n1698) );
  XOR U2806 ( .A(n5088), .B(n1698), .Z(out[1176]) );
  IV U2807 ( .A(n3081), .Z(n4205) );
  XOR U2808 ( .A(in[965]), .B(n4205), .Z(n5091) );
  NAND U2809 ( .A(n1701), .B(n1873), .Z(n1702) );
  XOR U2810 ( .A(n5091), .B(n1702), .Z(out[1177]) );
  IV U2811 ( .A(n3083), .Z(n4208) );
  XOR U2812 ( .A(in[966]), .B(n4208), .Z(n5094) );
  NAND U2813 ( .A(n1705), .B(n1875), .Z(n1706) );
  XOR U2814 ( .A(n5094), .B(n1706), .Z(out[1178]) );
  IV U2815 ( .A(n3085), .Z(n4211) );
  XOR U2816 ( .A(in[967]), .B(n4211), .Z(n5097) );
  NAND U2817 ( .A(n1709), .B(n1877), .Z(n1710) );
  XOR U2818 ( .A(n5097), .B(n1710), .Z(out[1179]) );
  IV U2819 ( .A(n2030), .Z(n4028) );
  XOR U2820 ( .A(in[588]), .B(n4028), .Z(n2833) );
  XNOR U2821 ( .A(in[1463]), .B(n4167), .Z(n3515) );
  XNOR U2822 ( .A(in[243]), .B(n4126), .Z(n3517) );
  NANDN U2823 ( .A(n3515), .B(n3517), .Z(n1711) );
  XNOR U2824 ( .A(n2833), .B(n1711), .Z(out[117]) );
  XNOR U2825 ( .A(n1713), .B(n1712), .Z(n4216) );
  XOR U2826 ( .A(in[968]), .B(n4216), .Z(n5101) );
  NAND U2827 ( .A(n1714), .B(n1879), .Z(n1715) );
  XNOR U2828 ( .A(n5101), .B(n1715), .Z(out[1180]) );
  IV U2829 ( .A(n3088), .Z(n4219) );
  XOR U2830 ( .A(in[969]), .B(n4219), .Z(n5104) );
  NAND U2831 ( .A(n1718), .B(n1881), .Z(n1719) );
  XOR U2832 ( .A(n5104), .B(n1719), .Z(out[1181]) );
  IV U2833 ( .A(n3090), .Z(n4222) );
  XOR U2834 ( .A(in[970]), .B(n4222), .Z(n5111) );
  NAND U2835 ( .A(n1722), .B(n1883), .Z(n1723) );
  XOR U2836 ( .A(n5111), .B(n1723), .Z(out[1182]) );
  XOR U2837 ( .A(in[971]), .B(n3092), .Z(n5115) );
  NAND U2838 ( .A(n1726), .B(n1885), .Z(n1727) );
  XNOR U2839 ( .A(n5115), .B(n1727), .Z(out[1183]) );
  XOR U2840 ( .A(in[972]), .B(n3094), .Z(n5119) );
  NAND U2841 ( .A(n1730), .B(n1887), .Z(n1731) );
  XNOR U2842 ( .A(n5119), .B(n1731), .Z(out[1184]) );
  XOR U2843 ( .A(in[973]), .B(n3098), .Z(n5123) );
  NAND U2844 ( .A(n1734), .B(n1889), .Z(n1735) );
  XNOR U2845 ( .A(n5123), .B(n1735), .Z(out[1185]) );
  XOR U2846 ( .A(in[974]), .B(n3100), .Z(n5127) );
  NAND U2847 ( .A(n1738), .B(n1893), .Z(n1739) );
  XNOR U2848 ( .A(n5127), .B(n1739), .Z(out[1186]) );
  XOR U2849 ( .A(n1741), .B(n1740), .Z(n4237) );
  XOR U2850 ( .A(in[975]), .B(n4237), .Z(n5131) );
  NAND U2851 ( .A(n1742), .B(n1895), .Z(n1743) );
  XNOR U2852 ( .A(n5131), .B(n1743), .Z(out[1187]) );
  XOR U2853 ( .A(in[976]), .B(n3103), .Z(n5135) );
  NAND U2854 ( .A(n1746), .B(n1897), .Z(n1747) );
  XNOR U2855 ( .A(n5135), .B(n1747), .Z(out[1188]) );
  IV U2856 ( .A(n3105), .Z(n4239) );
  XOR U2857 ( .A(in[977]), .B(n4239), .Z(n5138) );
  NAND U2858 ( .A(n1750), .B(n1899), .Z(n1751) );
  XOR U2859 ( .A(n5138), .B(n1751), .Z(out[1189]) );
  XNOR U2860 ( .A(in[589]), .B(n4032), .Z(n2835) );
  XNOR U2861 ( .A(in[1464]), .B(n4171), .Z(n3545) );
  XNOR U2862 ( .A(in[244]), .B(n4130), .Z(n3547) );
  NANDN U2863 ( .A(n3545), .B(n3547), .Z(n1752) );
  XNOR U2864 ( .A(n2835), .B(n1752), .Z(out[118]) );
  XOR U2865 ( .A(in[978]), .B(n3107), .Z(n5141) );
  NAND U2866 ( .A(n1755), .B(n1901), .Z(n1756) );
  XNOR U2867 ( .A(n5141), .B(n1756), .Z(out[1190]) );
  XOR U2868 ( .A(in[979]), .B(n3109), .Z(n5146) );
  NAND U2869 ( .A(n1759), .B(n1903), .Z(n1760) );
  XNOR U2870 ( .A(n5146), .B(n1760), .Z(out[1191]) );
  OR U2871 ( .A(n1906), .B(n1761), .Z(n1762) );
  XNOR U2872 ( .A(n1905), .B(n1762), .Z(out[1192]) );
  OR U2873 ( .A(n1910), .B(n1763), .Z(n1764) );
  XNOR U2874 ( .A(n1909), .B(n1764), .Z(out[1193]) );
  OR U2875 ( .A(n1914), .B(n1765), .Z(n1766) );
  XNOR U2876 ( .A(n1913), .B(n1766), .Z(out[1194]) );
  OR U2877 ( .A(n1924), .B(n1768), .Z(n1769) );
  XNOR U2878 ( .A(n1923), .B(n1769), .Z(out[1196]) );
  OR U2879 ( .A(n1928), .B(n1770), .Z(n1771) );
  XNOR U2880 ( .A(n1927), .B(n1771), .Z(out[1197]) );
  OR U2881 ( .A(n1932), .B(n1772), .Z(n1773) );
  XNOR U2882 ( .A(n1931), .B(n1773), .Z(out[1198]) );
  OR U2883 ( .A(n1936), .B(n1774), .Z(n1775) );
  XNOR U2884 ( .A(n1935), .B(n1775), .Z(out[1199]) );
  IV U2885 ( .A(n3118), .Z(n4036) );
  XOR U2886 ( .A(in[590]), .B(n4036), .Z(n2837) );
  XNOR U2887 ( .A(in[1465]), .B(n4175), .Z(n3575) );
  XNOR U2888 ( .A(in[245]), .B(n4134), .Z(n3577) );
  NANDN U2889 ( .A(n3575), .B(n3577), .Z(n1776) );
  XNOR U2890 ( .A(n2837), .B(n1776), .Z(out[119]) );
  XNOR U2891 ( .A(in[201]), .B(n3942), .Z(n4305) );
  XOR U2892 ( .A(in[1421]), .B(n3196), .Z(n4306) );
  XNOR U2893 ( .A(in[1044]), .B(n4486), .Z(n2886) );
  NANDN U2894 ( .A(n4306), .B(n2886), .Z(n1777) );
  XNOR U2895 ( .A(n4305), .B(n1777), .Z(out[11]) );
  OR U2896 ( .A(n1940), .B(n1778), .Z(n1779) );
  XNOR U2897 ( .A(n1939), .B(n1779), .Z(out[1200]) );
  OR U2898 ( .A(n1944), .B(n1780), .Z(n1781) );
  XNOR U2899 ( .A(n1943), .B(n1781), .Z(out[1201]) );
  OR U2900 ( .A(n1948), .B(n1782), .Z(n1783) );
  XNOR U2901 ( .A(n1947), .B(n1783), .Z(out[1202]) );
  OR U2902 ( .A(n1952), .B(n1784), .Z(n1785) );
  XNOR U2903 ( .A(n1951), .B(n1785), .Z(out[1203]) );
  OR U2904 ( .A(n1956), .B(n1786), .Z(n1787) );
  XNOR U2905 ( .A(n1955), .B(n1787), .Z(out[1204]) );
  OR U2906 ( .A(n1960), .B(n1788), .Z(n1789) );
  XNOR U2907 ( .A(n1959), .B(n1789), .Z(out[1205]) );
  OR U2908 ( .A(n1966), .B(n1790), .Z(n1791) );
  XNOR U2909 ( .A(n1965), .B(n1791), .Z(out[1206]) );
  OR U2910 ( .A(n1970), .B(n1792), .Z(n1793) );
  XNOR U2911 ( .A(n1969), .B(n1793), .Z(out[1207]) );
  OR U2912 ( .A(n1974), .B(n1794), .Z(n1795) );
  XNOR U2913 ( .A(n1973), .B(n1795), .Z(out[1208]) );
  OR U2914 ( .A(n1978), .B(n1796), .Z(n1797) );
  XNOR U2915 ( .A(n1977), .B(n1797), .Z(out[1209]) );
  XNOR U2916 ( .A(in[591]), .B(n4040), .Z(n2839) );
  IV U2917 ( .A(n1798), .Z(n3899) );
  XOR U2918 ( .A(in[1466]), .B(n3899), .Z(n3599) );
  XNOR U2919 ( .A(in[246]), .B(n4138), .Z(n3601) );
  NANDN U2920 ( .A(n3599), .B(n3601), .Z(n1799) );
  XNOR U2921 ( .A(n2839), .B(n1799), .Z(out[120]) );
  OR U2922 ( .A(n1982), .B(n1800), .Z(n1801) );
  XNOR U2923 ( .A(n1981), .B(n1801), .Z(out[1210]) );
  OR U2924 ( .A(n1986), .B(n1802), .Z(n1803) );
  XNOR U2925 ( .A(n1985), .B(n1803), .Z(out[1211]) );
  OR U2926 ( .A(n1990), .B(n1804), .Z(n1805) );
  XNOR U2927 ( .A(n1989), .B(n1805), .Z(out[1212]) );
  OR U2928 ( .A(n1994), .B(n1806), .Z(n1807) );
  XNOR U2929 ( .A(n1993), .B(n1807), .Z(out[1213]) );
  OR U2930 ( .A(n1998), .B(n1808), .Z(n1809) );
  XNOR U2931 ( .A(n1997), .B(n1809), .Z(out[1214]) );
  OR U2932 ( .A(n2002), .B(n1810), .Z(n1811) );
  XNOR U2933 ( .A(n2001), .B(n1811), .Z(out[1215]) );
  IV U2934 ( .A(n1812), .Z(n4991) );
  NANDN U2935 ( .A(n1813), .B(n4991), .Z(n1814) );
  XOR U2936 ( .A(n4992), .B(n1814), .Z(out[1216]) );
  IV U2937 ( .A(n1815), .Z(n4995) );
  NANDN U2938 ( .A(n1816), .B(n4995), .Z(n1817) );
  XOR U2939 ( .A(n4996), .B(n1817), .Z(out[1217]) );
  IV U2940 ( .A(n1818), .Z(n4999) );
  NANDN U2941 ( .A(n1819), .B(n4999), .Z(n1820) );
  XOR U2942 ( .A(n5000), .B(n1820), .Z(out[1218]) );
  IV U2943 ( .A(n1821), .Z(n5003) );
  NANDN U2944 ( .A(n1822), .B(n5003), .Z(n1823) );
  XOR U2945 ( .A(n5004), .B(n1823), .Z(out[1219]) );
  XNOR U2946 ( .A(in[592]), .B(n4044), .Z(n2841) );
  IV U2947 ( .A(n1824), .Z(n3903) );
  XOR U2948 ( .A(in[1467]), .B(n3903), .Z(n3629) );
  XNOR U2949 ( .A(in[247]), .B(n4142), .Z(n3631) );
  NANDN U2950 ( .A(n3629), .B(n3631), .Z(n1825) );
  XNOR U2951 ( .A(n2841), .B(n1825), .Z(out[121]) );
  IV U2952 ( .A(n1826), .Z(n5007) );
  NANDN U2953 ( .A(n1827), .B(n5007), .Z(n1828) );
  XOR U2954 ( .A(n5008), .B(n1828), .Z(out[1220]) );
  IV U2955 ( .A(n1829), .Z(n5011) );
  NANDN U2956 ( .A(n1830), .B(n5011), .Z(n1831) );
  XOR U2957 ( .A(n5012), .B(n1831), .Z(out[1221]) );
  OR U2958 ( .A(n5020), .B(n1833), .Z(n1834) );
  XNOR U2959 ( .A(n5019), .B(n1834), .Z(out[1223]) );
  OR U2960 ( .A(n5024), .B(n1835), .Z(n1836) );
  XNOR U2961 ( .A(n5023), .B(n1836), .Z(out[1224]) );
  OR U2962 ( .A(n5028), .B(n1837), .Z(n1838) );
  XNOR U2963 ( .A(n5027), .B(n1838), .Z(out[1225]) );
  OR U2964 ( .A(n5036), .B(n1839), .Z(n1840) );
  XNOR U2965 ( .A(n5035), .B(n1840), .Z(out[1226]) );
  OR U2966 ( .A(n5040), .B(n1841), .Z(n1842) );
  XNOR U2967 ( .A(n5039), .B(n1842), .Z(out[1227]) );
  OR U2968 ( .A(n5044), .B(n1843), .Z(n1844) );
  XNOR U2969 ( .A(n5043), .B(n1844), .Z(out[1228]) );
  OR U2970 ( .A(n5048), .B(n1845), .Z(n1846) );
  XNOR U2971 ( .A(n5047), .B(n1846), .Z(out[1229]) );
  IV U2972 ( .A(n2036), .Z(n4048) );
  XOR U2973 ( .A(in[593]), .B(n4048), .Z(n2846) );
  IV U2974 ( .A(n1847), .Z(n3907) );
  XOR U2975 ( .A(in[1468]), .B(n3907), .Z(n3673) );
  XNOR U2976 ( .A(in[248]), .B(n4146), .Z(n3675) );
  NANDN U2977 ( .A(n3673), .B(n3675), .Z(n1848) );
  XNOR U2978 ( .A(n2846), .B(n1848), .Z(out[122]) );
  OR U2979 ( .A(n5052), .B(n1849), .Z(n1850) );
  XNOR U2980 ( .A(n5051), .B(n1850), .Z(out[1230]) );
  OR U2981 ( .A(n5056), .B(n1851), .Z(n1852) );
  XNOR U2982 ( .A(n5055), .B(n1852), .Z(out[1231]) );
  NANDN U2983 ( .A(n1853), .B(n5059), .Z(n1854) );
  XNOR U2984 ( .A(n5060), .B(n1854), .Z(out[1232]) );
  NANDN U2985 ( .A(n1855), .B(n5062), .Z(n1856) );
  XNOR U2986 ( .A(n5063), .B(n1856), .Z(out[1233]) );
  NANDN U2987 ( .A(n1857), .B(n5065), .Z(n1858) );
  XNOR U2988 ( .A(n5066), .B(n1858), .Z(out[1234]) );
  OR U2989 ( .A(n5069), .B(n1859), .Z(n1860) );
  XNOR U2990 ( .A(n5068), .B(n1860), .Z(out[1235]) );
  NANDN U2991 ( .A(n1861), .B(n5076), .Z(n1862) );
  XNOR U2992 ( .A(n5077), .B(n1862), .Z(out[1236]) );
  NANDN U2993 ( .A(n1863), .B(n5079), .Z(n1864) );
  XNOR U2994 ( .A(n5080), .B(n1864), .Z(out[1237]) );
  NANDN U2995 ( .A(n1865), .B(n5082), .Z(n1866) );
  XNOR U2996 ( .A(n5083), .B(n1866), .Z(out[1238]) );
  NANDN U2997 ( .A(n1867), .B(n5085), .Z(n1868) );
  XNOR U2998 ( .A(n5086), .B(n1868), .Z(out[1239]) );
  IV U2999 ( .A(n2039), .Z(n4052) );
  XOR U3000 ( .A(in[594]), .B(n4052), .Z(n2848) );
  IV U3001 ( .A(n1869), .Z(n3911) );
  XOR U3002 ( .A(in[1469]), .B(n3911), .Z(n3717) );
  XNOR U3003 ( .A(in[249]), .B(n4150), .Z(n3719) );
  NANDN U3004 ( .A(n3717), .B(n3719), .Z(n1870) );
  XNOR U3005 ( .A(n2848), .B(n1870), .Z(out[123]) );
  NANDN U3006 ( .A(n1871), .B(n5088), .Z(n1872) );
  XNOR U3007 ( .A(n5089), .B(n1872), .Z(out[1240]) );
  NANDN U3008 ( .A(n1873), .B(n5091), .Z(n1874) );
  XNOR U3009 ( .A(n5092), .B(n1874), .Z(out[1241]) );
  NANDN U3010 ( .A(n1875), .B(n5094), .Z(n1876) );
  XNOR U3011 ( .A(n5095), .B(n1876), .Z(out[1242]) );
  NANDN U3012 ( .A(n1877), .B(n5097), .Z(n1878) );
  XNOR U3013 ( .A(n5098), .B(n1878), .Z(out[1243]) );
  OR U3014 ( .A(n5101), .B(n1879), .Z(n1880) );
  XNOR U3015 ( .A(n5100), .B(n1880), .Z(out[1244]) );
  NANDN U3016 ( .A(n1881), .B(n5104), .Z(n1882) );
  XNOR U3017 ( .A(n5105), .B(n1882), .Z(out[1245]) );
  NANDN U3018 ( .A(n1883), .B(n5111), .Z(n1884) );
  XNOR U3019 ( .A(n5112), .B(n1884), .Z(out[1246]) );
  OR U3020 ( .A(n5115), .B(n1885), .Z(n1886) );
  XNOR U3021 ( .A(n5114), .B(n1886), .Z(out[1247]) );
  OR U3022 ( .A(n5119), .B(n1887), .Z(n1888) );
  XNOR U3023 ( .A(n5118), .B(n1888), .Z(out[1248]) );
  OR U3024 ( .A(n5123), .B(n1889), .Z(n1890) );
  XNOR U3025 ( .A(n5122), .B(n1890), .Z(out[1249]) );
  IV U3026 ( .A(n3124), .Z(n4056) );
  XOR U3027 ( .A(in[595]), .B(n4056), .Z(n2850) );
  IV U3028 ( .A(n1891), .Z(n3915) );
  XOR U3029 ( .A(in[1470]), .B(n3915), .Z(n3763) );
  XNOR U3030 ( .A(in[250]), .B(n4154), .Z(n3765) );
  NANDN U3031 ( .A(n3763), .B(n3765), .Z(n1892) );
  XNOR U3032 ( .A(n2850), .B(n1892), .Z(out[124]) );
  OR U3033 ( .A(n5127), .B(n1893), .Z(n1894) );
  XNOR U3034 ( .A(n5126), .B(n1894), .Z(out[1250]) );
  OR U3035 ( .A(n5131), .B(n1895), .Z(n1896) );
  XNOR U3036 ( .A(n5130), .B(n1896), .Z(out[1251]) );
  OR U3037 ( .A(n5135), .B(n1897), .Z(n1898) );
  XNOR U3038 ( .A(n5134), .B(n1898), .Z(out[1252]) );
  NANDN U3039 ( .A(n1899), .B(n5138), .Z(n1900) );
  XNOR U3040 ( .A(n5139), .B(n1900), .Z(out[1253]) );
  OR U3041 ( .A(n5141), .B(n1901), .Z(n1902) );
  XOR U3042 ( .A(n5142), .B(n1902), .Z(out[1254]) );
  OR U3043 ( .A(n5146), .B(n1903), .Z(n1904) );
  XNOR U3044 ( .A(n5145), .B(n1904), .Z(out[1255]) );
  ANDN U3045 ( .B(n1906), .A(n1905), .Z(n1907) );
  XOR U3046 ( .A(n1908), .B(n1907), .Z(out[1256]) );
  ANDN U3047 ( .B(n1910), .A(n1909), .Z(n1911) );
  XOR U3048 ( .A(n1912), .B(n1911), .Z(out[1257]) );
  ANDN U3049 ( .B(n1914), .A(n1913), .Z(n1915) );
  XOR U3050 ( .A(n1916), .B(n1915), .Z(out[1258]) );
  ANDN U3051 ( .B(n1918), .A(n1917), .Z(n1919) );
  XOR U3052 ( .A(n1920), .B(n1919), .Z(out[1259]) );
  IV U3053 ( .A(n3126), .Z(n4060) );
  XOR U3054 ( .A(in[596]), .B(n4060), .Z(n2852) );
  IV U3055 ( .A(n1921), .Z(n3919) );
  XOR U3056 ( .A(in[1471]), .B(n3919), .Z(n3807) );
  IV U3057 ( .A(n4164), .Z(n3278) );
  XOR U3058 ( .A(in[251]), .B(n3278), .Z(n3809) );
  OR U3059 ( .A(n3807), .B(n3809), .Z(n1922) );
  XNOR U3060 ( .A(n2852), .B(n1922), .Z(out[125]) );
  ANDN U3061 ( .B(n1924), .A(n1923), .Z(n1925) );
  XOR U3062 ( .A(n1926), .B(n1925), .Z(out[1260]) );
  ANDN U3063 ( .B(n1928), .A(n1927), .Z(n1929) );
  XOR U3064 ( .A(n1930), .B(n1929), .Z(out[1261]) );
  ANDN U3065 ( .B(n1932), .A(n1931), .Z(n1933) );
  XOR U3066 ( .A(n1934), .B(n1933), .Z(out[1262]) );
  ANDN U3067 ( .B(n1936), .A(n1935), .Z(n1937) );
  XOR U3068 ( .A(n1938), .B(n1937), .Z(out[1263]) );
  ANDN U3069 ( .B(n1940), .A(n1939), .Z(n1941) );
  XOR U3070 ( .A(n1942), .B(n1941), .Z(out[1264]) );
  ANDN U3071 ( .B(n1944), .A(n1943), .Z(n1945) );
  XOR U3072 ( .A(n1946), .B(n1945), .Z(out[1265]) );
  ANDN U3073 ( .B(n1948), .A(n1947), .Z(n1949) );
  XOR U3074 ( .A(n1950), .B(n1949), .Z(out[1266]) );
  ANDN U3075 ( .B(n1952), .A(n1951), .Z(n1953) );
  XOR U3076 ( .A(n1954), .B(n1953), .Z(out[1267]) );
  ANDN U3077 ( .B(n1956), .A(n1955), .Z(n1957) );
  XOR U3078 ( .A(n1958), .B(n1957), .Z(out[1268]) );
  ANDN U3079 ( .B(n1960), .A(n1959), .Z(n1961) );
  XOR U3080 ( .A(n1962), .B(n1961), .Z(out[1269]) );
  IV U3081 ( .A(n3128), .Z(n4064) );
  XOR U3082 ( .A(in[597]), .B(n4064), .Z(n2854) );
  IV U3083 ( .A(n1963), .Z(n3923) );
  XOR U3084 ( .A(in[1408]), .B(n3923), .Z(n3851) );
  IV U3085 ( .A(n4168), .Z(n3281) );
  XOR U3086 ( .A(in[252]), .B(n3281), .Z(n3853) );
  OR U3087 ( .A(n3851), .B(n3853), .Z(n1964) );
  XNOR U3088 ( .A(n2854), .B(n1964), .Z(out[126]) );
  ANDN U3089 ( .B(n1966), .A(n1965), .Z(n1967) );
  XOR U3090 ( .A(n1968), .B(n1967), .Z(out[1270]) );
  ANDN U3091 ( .B(n1970), .A(n1969), .Z(n1971) );
  XOR U3092 ( .A(n1972), .B(n1971), .Z(out[1271]) );
  ANDN U3093 ( .B(n1974), .A(n1973), .Z(n1975) );
  XOR U3094 ( .A(n1976), .B(n1975), .Z(out[1272]) );
  ANDN U3095 ( .B(n1978), .A(n1977), .Z(n1979) );
  XOR U3096 ( .A(n1980), .B(n1979), .Z(out[1273]) );
  ANDN U3097 ( .B(n1982), .A(n1981), .Z(n1983) );
  XOR U3098 ( .A(n1984), .B(n1983), .Z(out[1274]) );
  ANDN U3099 ( .B(n1986), .A(n1985), .Z(n1987) );
  XOR U3100 ( .A(n1988), .B(n1987), .Z(out[1275]) );
  ANDN U3101 ( .B(n1990), .A(n1989), .Z(n1991) );
  XOR U3102 ( .A(n1992), .B(n1991), .Z(out[1276]) );
  ANDN U3103 ( .B(n1994), .A(n1993), .Z(n1995) );
  XOR U3104 ( .A(n1996), .B(n1995), .Z(out[1277]) );
  ANDN U3105 ( .B(n1998), .A(n1997), .Z(n1999) );
  XOR U3106 ( .A(n2000), .B(n1999), .Z(out[1278]) );
  ANDN U3107 ( .B(n2002), .A(n2001), .Z(n2003) );
  XOR U3108 ( .A(n2004), .B(n2003), .Z(out[1279]) );
  IV U3109 ( .A(n3130), .Z(n4072) );
  XOR U3110 ( .A(in[598]), .B(n4072), .Z(n2856) );
  IV U3111 ( .A(n2005), .Z(n3927) );
  XOR U3112 ( .A(in[1409]), .B(n3927), .Z(n3895) );
  IV U3113 ( .A(n4172), .Z(n3284) );
  XOR U3114 ( .A(in[253]), .B(n3284), .Z(n3897) );
  OR U3115 ( .A(n3895), .B(n3897), .Z(n2006) );
  XNOR U3116 ( .A(n2856), .B(n2006), .Z(out[127]) );
  XOR U3117 ( .A(in[50]), .B(n4315), .Z(n2183) );
  XNOR U3118 ( .A(in[1172]), .B(n3989), .Z(n2440) );
  XNOR U3119 ( .A(in[1536]), .B(n3973), .Z(n2441) );
  NANDN U3120 ( .A(n2440), .B(n2441), .Z(n2007) );
  XNOR U3121 ( .A(n2183), .B(n2007), .Z(out[1280]) );
  XOR U3122 ( .A(in[51]), .B(n4318), .Z(n2185) );
  IV U3123 ( .A(n2008), .Z(n3993) );
  XOR U3124 ( .A(in[1173]), .B(n3993), .Z(n2443) );
  XNOR U3125 ( .A(in[1537]), .B(n3977), .Z(n2097) );
  IV U3126 ( .A(n2097), .Z(n2444) );
  OR U3127 ( .A(n2443), .B(n2444), .Z(n2009) );
  XNOR U3128 ( .A(n2185), .B(n2009), .Z(out[1281]) );
  XOR U3129 ( .A(in[52]), .B(n4321), .Z(n2188) );
  XNOR U3130 ( .A(in[1174]), .B(n3997), .Z(n2449) );
  XNOR U3131 ( .A(in[1538]), .B(n3984), .Z(n2447) );
  NANDN U3132 ( .A(n2449), .B(n2447), .Z(n2010) );
  XNOR U3133 ( .A(n2188), .B(n2010), .Z(out[1282]) );
  XOR U3134 ( .A(in[53]), .B(n4324), .Z(n2190) );
  XNOR U3135 ( .A(in[1175]), .B(n4001), .Z(n2451) );
  XNOR U3136 ( .A(in[1539]), .B(n3988), .Z(n2452) );
  NANDN U3137 ( .A(n2451), .B(n2452), .Z(n2011) );
  XNOR U3138 ( .A(n2190), .B(n2011), .Z(out[1283]) );
  XOR U3139 ( .A(in[54]), .B(n4327), .Z(n2192) );
  IV U3140 ( .A(n2012), .Z(n4005) );
  XOR U3141 ( .A(in[1176]), .B(n4005), .Z(n2457) );
  XOR U3142 ( .A(in[1540]), .B(n2013), .Z(n2101) );
  IV U3143 ( .A(n2101), .Z(n2459) );
  OR U3144 ( .A(n2457), .B(n2459), .Z(n2014) );
  XNOR U3145 ( .A(n2192), .B(n2014), .Z(out[1284]) );
  XOR U3146 ( .A(in[55]), .B(n4330), .Z(n2194) );
  IV U3147 ( .A(n2015), .Z(n4009) );
  XOR U3148 ( .A(in[1177]), .B(n4009), .Z(n2461) );
  XOR U3149 ( .A(in[1541]), .B(n2016), .Z(n2103) );
  IV U3150 ( .A(n2103), .Z(n2463) );
  OR U3151 ( .A(n2461), .B(n2463), .Z(n2017) );
  XNOR U3152 ( .A(n2194), .B(n2017), .Z(out[1285]) );
  XOR U3153 ( .A(in[56]), .B(n4178), .Z(n2196) );
  XNOR U3154 ( .A(in[1178]), .B(n4013), .Z(n2466) );
  XOR U3155 ( .A(in[1542]), .B(n2018), .Z(n2464) );
  NANDN U3156 ( .A(n2466), .B(n2464), .Z(n2019) );
  XNOR U3157 ( .A(n2196), .B(n2019), .Z(out[1286]) );
  XOR U3158 ( .A(in[57]), .B(n4181), .Z(n2198) );
  XNOR U3159 ( .A(in[1179]), .B(n4017), .Z(n2468) );
  XOR U3160 ( .A(in[1543]), .B(n2020), .Z(n2469) );
  NANDN U3161 ( .A(n2468), .B(n2469), .Z(n2021) );
  XNOR U3162 ( .A(n2198), .B(n2021), .Z(out[1287]) );
  XOR U3163 ( .A(in[58]), .B(n4184), .Z(n2200) );
  XNOR U3164 ( .A(in[1180]), .B(n4021), .Z(n2472) );
  XOR U3165 ( .A(in[1544]), .B(n2022), .Z(n2470) );
  NANDN U3166 ( .A(n2472), .B(n2470), .Z(n2023) );
  XNOR U3167 ( .A(n2200), .B(n2023), .Z(out[1288]) );
  XOR U3168 ( .A(in[59]), .B(n4187), .Z(n2202) );
  XNOR U3169 ( .A(in[1181]), .B(n4029), .Z(n2475) );
  XOR U3170 ( .A(in[1545]), .B(n2024), .Z(n2473) );
  NANDN U3171 ( .A(n2475), .B(n2473), .Z(n2025) );
  XNOR U3172 ( .A(n2202), .B(n2025), .Z(out[1289]) );
  XOR U3173 ( .A(in[665]), .B(n4253), .Z(n2858) );
  IV U3174 ( .A(n3132), .Z(n4076) );
  XOR U3175 ( .A(in[599]), .B(n4076), .Z(n3940) );
  OR U3176 ( .A(n3940), .B(n3938), .Z(n2026) );
  XNOR U3177 ( .A(n2858), .B(n2026), .Z(out[128]) );
  XOR U3178 ( .A(in[60]), .B(n3059), .Z(n2204) );
  XNOR U3179 ( .A(in[1182]), .B(n4033), .Z(n2478) );
  XOR U3180 ( .A(in[1546]), .B(n2027), .Z(n2476) );
  NANDN U3181 ( .A(n2478), .B(n2476), .Z(n2028) );
  XNOR U3182 ( .A(n2204), .B(n2028), .Z(out[1290]) );
  XOR U3183 ( .A(in[61]), .B(n3061), .Z(n2206) );
  XNOR U3184 ( .A(in[1183]), .B(n4037), .Z(n2480) );
  XOR U3185 ( .A(in[1547]), .B(n4020), .Z(n2482) );
  NANDN U3186 ( .A(n2480), .B(n2482), .Z(n2029) );
  XNOR U3187 ( .A(n2206), .B(n2029), .Z(out[1291]) );
  XOR U3188 ( .A(in[62]), .B(n3063), .Z(n2209) );
  XNOR U3189 ( .A(in[1184]), .B(n4041), .Z(n2485) );
  XOR U3190 ( .A(in[1548]), .B(n2030), .Z(n2483) );
  NANDN U3191 ( .A(n2485), .B(n2483), .Z(n2031) );
  XNOR U3192 ( .A(n2209), .B(n2031), .Z(out[1292]) );
  XOR U3193 ( .A(in[63]), .B(n4199), .Z(n2211) );
  XNOR U3194 ( .A(in[1185]), .B(n4045), .Z(n2487) );
  XOR U3195 ( .A(in[1549]), .B(n4032), .Z(n2489) );
  NANDN U3196 ( .A(n2487), .B(n2489), .Z(n2032) );
  XNOR U3197 ( .A(n2211), .B(n2032), .Z(out[1293]) );
  XOR U3198 ( .A(in[0]), .B(n3068), .Z(n2213) );
  XOR U3199 ( .A(in[1550]), .B(n4036), .Z(n2494) );
  XNOR U3200 ( .A(n3393), .B(in[1186]), .Z(n2491) );
  NANDN U3201 ( .A(n2494), .B(n2491), .Z(n2033) );
  XNOR U3202 ( .A(n2213), .B(n2033), .Z(out[1294]) );
  XOR U3203 ( .A(in[1]), .B(n3071), .Z(n2215) );
  XNOR U3204 ( .A(in[1551]), .B(n4040), .Z(n2497) );
  XNOR U3205 ( .A(n3396), .B(in[1187]), .Z(n2495) );
  NANDN U3206 ( .A(n2497), .B(n2495), .Z(n2034) );
  XNOR U3207 ( .A(n2215), .B(n2034), .Z(out[1295]) );
  XOR U3208 ( .A(in[2]), .B(n3073), .Z(n2218) );
  XNOR U3209 ( .A(in[1552]), .B(n4044), .Z(n2503) );
  XNOR U3210 ( .A(n3400), .B(in[1188]), .Z(n2500) );
  NANDN U3211 ( .A(n2503), .B(n2500), .Z(n2035) );
  XNOR U3212 ( .A(n2218), .B(n2035), .Z(out[1296]) );
  XOR U3213 ( .A(in[3]), .B(n3077), .Z(n2220) );
  XOR U3214 ( .A(n3404), .B(in[1189]), .Z(n2505) );
  XOR U3215 ( .A(in[1553]), .B(n2036), .Z(n2117) );
  IV U3216 ( .A(n2117), .Z(n2507) );
  OR U3217 ( .A(n2505), .B(n2507), .Z(n2037) );
  XNOR U3218 ( .A(n2220), .B(n2037), .Z(out[1297]) );
  XOR U3219 ( .A(in[4]), .B(n3079), .Z(n2222) );
  IV U3220 ( .A(n2038), .Z(n4065) );
  XOR U3221 ( .A(in[1190]), .B(n4065), .Z(n2509) );
  XOR U3222 ( .A(in[1554]), .B(n2039), .Z(n2119) );
  IV U3223 ( .A(n2119), .Z(n2511) );
  OR U3224 ( .A(n2509), .B(n2511), .Z(n2040) );
  XNOR U3225 ( .A(n2222), .B(n2040), .Z(out[1298]) );
  XOR U3226 ( .A(in[5]), .B(n3081), .Z(n2224) );
  IV U3227 ( .A(n2041), .Z(n4073) );
  XOR U3228 ( .A(in[1191]), .B(n4073), .Z(n2513) );
  XOR U3229 ( .A(in[1555]), .B(n4056), .Z(n2515) );
  OR U3230 ( .A(n2513), .B(n2515), .Z(n2042) );
  XNOR U3231 ( .A(n2224), .B(n2042), .Z(out[1299]) );
  XOR U3232 ( .A(in[666]), .B(n4254), .Z(n2861) );
  IV U3233 ( .A(n3138), .Z(n4080) );
  XOR U3234 ( .A(in[600]), .B(n4080), .Z(n3983) );
  XNOR U3235 ( .A(in[255]), .B(n3290), .Z(n3982) );
  NANDN U3236 ( .A(n3983), .B(n3982), .Z(n2043) );
  XNOR U3237 ( .A(n2861), .B(n2043), .Z(out[129]) );
  XNOR U3238 ( .A(in[202]), .B(n3946), .Z(n4337) );
  XOR U3239 ( .A(in[1422]), .B(n3199), .Z(n4338) );
  XNOR U3240 ( .A(in[1045]), .B(n4489), .Z(n2888) );
  NANDN U3241 ( .A(n4338), .B(n2888), .Z(n2044) );
  XNOR U3242 ( .A(n4337), .B(n2044), .Z(out[12]) );
  XOR U3243 ( .A(in[6]), .B(n3083), .Z(n2226) );
  IV U3244 ( .A(n2045), .Z(n4077) );
  XOR U3245 ( .A(in[1192]), .B(n4077), .Z(n2517) );
  XOR U3246 ( .A(in[1556]), .B(n3126), .Z(n2121) );
  IV U3247 ( .A(n2121), .Z(n2519) );
  OR U3248 ( .A(n2517), .B(n2519), .Z(n2046) );
  XNOR U3249 ( .A(n2226), .B(n2046), .Z(out[1300]) );
  XOR U3250 ( .A(in[7]), .B(n3085), .Z(n2228) );
  IV U3251 ( .A(n2047), .Z(n4081) );
  XOR U3252 ( .A(in[1193]), .B(n4081), .Z(n2521) );
  XOR U3253 ( .A(in[1557]), .B(n3128), .Z(n2123) );
  IV U3254 ( .A(n2123), .Z(n2523) );
  OR U3255 ( .A(n2521), .B(n2523), .Z(n2048) );
  XNOR U3256 ( .A(n2228), .B(n2048), .Z(out[1301]) );
  XOR U3257 ( .A(in[8]), .B(n4216), .Z(n2231) );
  IV U3258 ( .A(n2049), .Z(n4085) );
  XOR U3259 ( .A(in[1194]), .B(n4085), .Z(n2525) );
  XOR U3260 ( .A(in[1558]), .B(n4072), .Z(n2527) );
  OR U3261 ( .A(n2525), .B(n2527), .Z(n2050) );
  XNOR U3262 ( .A(n2231), .B(n2050), .Z(out[1302]) );
  XOR U3263 ( .A(in[9]), .B(n3088), .Z(n2233) );
  XOR U3264 ( .A(in[1559]), .B(n4076), .Z(n2531) );
  XOR U3265 ( .A(in[1195]), .B(n4090), .Z(n2529) );
  NANDN U3266 ( .A(n2531), .B(n2529), .Z(n2051) );
  XNOR U3267 ( .A(n2233), .B(n2051), .Z(out[1303]) );
  XOR U3268 ( .A(in[10]), .B(n3090), .Z(n2235) );
  XOR U3269 ( .A(in[1560]), .B(n3138), .Z(n2125) );
  IV U3270 ( .A(n2125), .Z(n2536) );
  XOR U3271 ( .A(in[1196]), .B(n4094), .Z(n2534) );
  NANDN U3272 ( .A(n2536), .B(n2534), .Z(n2052) );
  XNOR U3273 ( .A(n2235), .B(n2052), .Z(out[1304]) );
  XOR U3274 ( .A(in[11]), .B(n3092), .Z(n2237) );
  XOR U3275 ( .A(in[1561]), .B(n3140), .Z(n2127) );
  IV U3276 ( .A(n2127), .Z(n2540) );
  XOR U3277 ( .A(in[1197]), .B(n4098), .Z(n2538) );
  NANDN U3278 ( .A(n2540), .B(n2538), .Z(n2053) );
  XNOR U3279 ( .A(n2237), .B(n2053), .Z(out[1305]) );
  XOR U3280 ( .A(in[12]), .B(n3094), .Z(n2239) );
  IV U3281 ( .A(n3143), .Z(n4088) );
  XOR U3282 ( .A(in[1562]), .B(n4088), .Z(n2544) );
  XOR U3283 ( .A(in[1198]), .B(n4102), .Z(n2542) );
  NANDN U3284 ( .A(n2544), .B(n2542), .Z(n2054) );
  XNOR U3285 ( .A(n2239), .B(n2054), .Z(out[1306]) );
  XOR U3286 ( .A(in[13]), .B(n3098), .Z(n2241) );
  IV U3287 ( .A(n3145), .Z(n4092) );
  XOR U3288 ( .A(in[1563]), .B(n4092), .Z(n2548) );
  XOR U3289 ( .A(in[1199]), .B(n4106), .Z(n2546) );
  NANDN U3290 ( .A(n2548), .B(n2546), .Z(n2055) );
  XNOR U3291 ( .A(n2241), .B(n2055), .Z(out[1307]) );
  XOR U3292 ( .A(in[14]), .B(n3100), .Z(n2243) );
  IV U3293 ( .A(n3024), .Z(n4096) );
  XOR U3294 ( .A(in[1564]), .B(n4096), .Z(n2552) );
  XOR U3295 ( .A(in[1200]), .B(n4110), .Z(n2550) );
  NANDN U3296 ( .A(n2552), .B(n2550), .Z(n2056) );
  XNOR U3297 ( .A(n2243), .B(n2056), .Z(out[1308]) );
  XOR U3298 ( .A(in[15]), .B(n4237), .Z(n2245) );
  IV U3299 ( .A(n3026), .Z(n4100) );
  XOR U3300 ( .A(in[1565]), .B(n4100), .Z(n2556) );
  XOR U3301 ( .A(in[1201]), .B(n4118), .Z(n2554) );
  NANDN U3302 ( .A(n2556), .B(n2554), .Z(n2057) );
  XNOR U3303 ( .A(n2245), .B(n2057), .Z(out[1309]) );
  XOR U3304 ( .A(in[667]), .B(n4255), .Z(n2747) );
  IV U3305 ( .A(n2747), .Z(n2863) );
  IV U3306 ( .A(n3140), .Z(n4084) );
  XOR U3307 ( .A(in[601]), .B(n4084), .Z(n4027) );
  XNOR U3308 ( .A(in[192]), .B(n3293), .Z(n4024) );
  NANDN U3309 ( .A(n4027), .B(n4024), .Z(n2058) );
  XOR U3310 ( .A(n2863), .B(n2058), .Z(out[130]) );
  XOR U3311 ( .A(in[16]), .B(n3103), .Z(n2247) );
  IV U3312 ( .A(n3028), .Z(n4104) );
  XOR U3313 ( .A(in[1566]), .B(n4104), .Z(n2560) );
  XOR U3314 ( .A(in[1202]), .B(n4122), .Z(n2558) );
  NANDN U3315 ( .A(n2560), .B(n2558), .Z(n2059) );
  XNOR U3316 ( .A(n2247), .B(n2059), .Z(out[1310]) );
  XOR U3317 ( .A(in[17]), .B(n3105), .Z(n2249) );
  IV U3318 ( .A(n3030), .Z(n4108) );
  XOR U3319 ( .A(in[1567]), .B(n4108), .Z(n2563) );
  XOR U3320 ( .A(in[1203]), .B(n4126), .Z(n2562) );
  NANDN U3321 ( .A(n2563), .B(n2562), .Z(n2060) );
  XNOR U3322 ( .A(n2249), .B(n2060), .Z(out[1311]) );
  XOR U3323 ( .A(in[18]), .B(n3107), .Z(n2252) );
  IV U3324 ( .A(n3032), .Z(n4116) );
  XOR U3325 ( .A(in[1568]), .B(n4116), .Z(n2569) );
  XOR U3326 ( .A(in[1204]), .B(n4130), .Z(n2567) );
  NANDN U3327 ( .A(n2569), .B(n2567), .Z(n2061) );
  XNOR U3328 ( .A(n2252), .B(n2061), .Z(out[1312]) );
  XOR U3329 ( .A(in[19]), .B(n3109), .Z(n2254) );
  XOR U3330 ( .A(in[1569]), .B(n3034), .Z(n2131) );
  IV U3331 ( .A(n2131), .Z(n2573) );
  XOR U3332 ( .A(in[1205]), .B(n4134), .Z(n2571) );
  NANDN U3333 ( .A(n2573), .B(n2571), .Z(n2062) );
  XNOR U3334 ( .A(n2254), .B(n2062), .Z(out[1313]) );
  XOR U3335 ( .A(in[20]), .B(n4248), .Z(n2256) );
  XOR U3336 ( .A(in[1570]), .B(n2170), .Z(n2133) );
  IV U3337 ( .A(n2133), .Z(n2579) );
  XOR U3338 ( .A(in[1206]), .B(n4138), .Z(n2577) );
  NANDN U3339 ( .A(n2579), .B(n2577), .Z(n2063) );
  XNOR U3340 ( .A(n2256), .B(n2063), .Z(out[1314]) );
  XOR U3341 ( .A(in[21]), .B(n4249), .Z(n2258) );
  XOR U3342 ( .A(in[1571]), .B(n3037), .Z(n2135) );
  IV U3343 ( .A(n2135), .Z(n2583) );
  XOR U3344 ( .A(in[1207]), .B(n4142), .Z(n2581) );
  NANDN U3345 ( .A(n2583), .B(n2581), .Z(n2064) );
  XNOR U3346 ( .A(n2258), .B(n2064), .Z(out[1315]) );
  XOR U3347 ( .A(in[22]), .B(n4250), .Z(n2260) );
  XOR U3348 ( .A(in[1572]), .B(n3039), .Z(n2138) );
  IV U3349 ( .A(n2138), .Z(n2587) );
  XOR U3350 ( .A(in[1208]), .B(n4146), .Z(n2585) );
  NANDN U3351 ( .A(n2587), .B(n2585), .Z(n2065) );
  XNOR U3352 ( .A(n2260), .B(n2065), .Z(out[1316]) );
  XOR U3353 ( .A(in[23]), .B(n4251), .Z(n2262) );
  XNOR U3354 ( .A(in[1573]), .B(n4136), .Z(n2140) );
  IV U3355 ( .A(n2140), .Z(n2591) );
  XOR U3356 ( .A(in[1209]), .B(n4150), .Z(n2589) );
  NANDN U3357 ( .A(n2591), .B(n2589), .Z(n2066) );
  XNOR U3358 ( .A(n2262), .B(n2066), .Z(out[1317]) );
  XOR U3359 ( .A(in[24]), .B(n4252), .Z(n2264) );
  XNOR U3360 ( .A(in[1574]), .B(n4140), .Z(n2595) );
  XOR U3361 ( .A(in[1210]), .B(n4154), .Z(n2593) );
  NAND U3362 ( .A(n2595), .B(n2593), .Z(n2067) );
  XNOR U3363 ( .A(n2264), .B(n2067), .Z(out[1318]) );
  XOR U3364 ( .A(in[25]), .B(n4253), .Z(n2266) );
  XOR U3365 ( .A(in[1211]), .B(n4164), .Z(n2597) );
  XNOR U3366 ( .A(in[1575]), .B(n4144), .Z(n2143) );
  IV U3367 ( .A(n2143), .Z(n2599) );
  OR U3368 ( .A(n2597), .B(n2599), .Z(n2068) );
  XNOR U3369 ( .A(n2266), .B(n2068), .Z(out[1319]) );
  XOR U3370 ( .A(in[668]), .B(n4258), .Z(n2749) );
  IV U3371 ( .A(n2749), .Z(n2865) );
  XOR U3372 ( .A(in[602]), .B(n4088), .Z(n4071) );
  XNOR U3373 ( .A(in[193]), .B(n3296), .Z(n4068) );
  NANDN U3374 ( .A(n4071), .B(n4068), .Z(n2069) );
  XOR U3375 ( .A(n2865), .B(n2069), .Z(out[131]) );
  XOR U3376 ( .A(in[26]), .B(n4254), .Z(n2268) );
  XOR U3377 ( .A(in[1212]), .B(n4168), .Z(n2601) );
  XNOR U3378 ( .A(in[1576]), .B(n4148), .Z(n2145) );
  IV U3379 ( .A(n2145), .Z(n2603) );
  OR U3380 ( .A(n2601), .B(n2603), .Z(n2070) );
  XNOR U3381 ( .A(n2268), .B(n2070), .Z(out[1320]) );
  XOR U3382 ( .A(in[27]), .B(n4255), .Z(n2270) );
  XOR U3383 ( .A(in[1213]), .B(n4172), .Z(n2605) );
  XNOR U3384 ( .A(in[1577]), .B(n4152), .Z(n2147) );
  IV U3385 ( .A(n2147), .Z(n2607) );
  OR U3386 ( .A(n2605), .B(n2607), .Z(n2071) );
  XNOR U3387 ( .A(n2270), .B(n2071), .Z(out[1321]) );
  XOR U3388 ( .A(in[28]), .B(n4258), .Z(n2273) );
  XNOR U3389 ( .A(in[1578]), .B(n4162), .Z(n2149) );
  IV U3390 ( .A(n2149), .Z(n2611) );
  XOR U3391 ( .A(in[1214]), .B(n4176), .Z(n2609) );
  NANDN U3392 ( .A(n2611), .B(n2609), .Z(n2072) );
  XNOR U3393 ( .A(n2273), .B(n2072), .Z(out[1322]) );
  XOR U3394 ( .A(in[29]), .B(n4259), .Z(n2275) );
  XOR U3395 ( .A(in[1215]), .B(n3290), .Z(n2613) );
  XNOR U3396 ( .A(in[1579]), .B(n4166), .Z(n2151) );
  IV U3397 ( .A(n2151), .Z(n2615) );
  OR U3398 ( .A(n2613), .B(n2615), .Z(n2073) );
  XNOR U3399 ( .A(n2275), .B(n2073), .Z(out[1323]) );
  XOR U3400 ( .A(in[30]), .B(n4260), .Z(n2277) );
  XOR U3401 ( .A(in[1152]), .B(n3293), .Z(n2619) );
  XNOR U3402 ( .A(in[1580]), .B(n4170), .Z(n2153) );
  IV U3403 ( .A(n2153), .Z(n2621) );
  OR U3404 ( .A(n2619), .B(n2621), .Z(n2074) );
  XNOR U3405 ( .A(n2277), .B(n2074), .Z(out[1324]) );
  XOR U3406 ( .A(in[31]), .B(n4261), .Z(n2279) );
  XOR U3407 ( .A(in[1153]), .B(n3296), .Z(n2623) );
  XNOR U3408 ( .A(in[1581]), .B(n4174), .Z(n2155) );
  IV U3409 ( .A(n2155), .Z(n2625) );
  OR U3410 ( .A(n2623), .B(n2625), .Z(n2075) );
  XNOR U3411 ( .A(n2279), .B(n2075), .Z(out[1325]) );
  XOR U3412 ( .A(in[32]), .B(n4264), .Z(n2281) );
  XOR U3413 ( .A(in[1154]), .B(n3303), .Z(n2627) );
  XNOR U3414 ( .A(in[1582]), .B(n3898), .Z(n2158) );
  IV U3415 ( .A(n2158), .Z(n2629) );
  OR U3416 ( .A(n2627), .B(n2629), .Z(n2076) );
  XNOR U3417 ( .A(n2281), .B(n2076), .Z(out[1326]) );
  XOR U3418 ( .A(in[33]), .B(n4267), .Z(n2283) );
  XOR U3419 ( .A(in[1155]), .B(n3306), .Z(n2631) );
  XNOR U3420 ( .A(in[1583]), .B(n3902), .Z(n2160) );
  IV U3421 ( .A(n2160), .Z(n2633) );
  OR U3422 ( .A(n2631), .B(n2633), .Z(n2077) );
  XNOR U3423 ( .A(n2283), .B(n2077), .Z(out[1327]) );
  XOR U3424 ( .A(in[34]), .B(n4270), .Z(n2285) );
  XOR U3425 ( .A(in[1156]), .B(n3309), .Z(n2635) );
  XNOR U3426 ( .A(in[1584]), .B(n3906), .Z(n2162) );
  IV U3427 ( .A(n2162), .Z(n2637) );
  OR U3428 ( .A(n2635), .B(n2637), .Z(n2078) );
  XNOR U3429 ( .A(n2285), .B(n2078), .Z(out[1328]) );
  IV U3430 ( .A(n4273), .Z(n3142) );
  XOR U3431 ( .A(in[35]), .B(n3142), .Z(n2287) );
  XOR U3432 ( .A(in[1157]), .B(n3312), .Z(n2639) );
  XNOR U3433 ( .A(in[1585]), .B(n3910), .Z(n2164) );
  IV U3434 ( .A(n2164), .Z(n2641) );
  OR U3435 ( .A(n2639), .B(n2641), .Z(n2079) );
  XNOR U3436 ( .A(n2287), .B(n2079), .Z(out[1329]) );
  XOR U3437 ( .A(in[669]), .B(n4259), .Z(n2751) );
  IV U3438 ( .A(n2751), .Z(n2870) );
  XOR U3439 ( .A(in[603]), .B(n4092), .Z(n4115) );
  XNOR U3440 ( .A(in[194]), .B(n3303), .Z(n4112) );
  NANDN U3441 ( .A(n4115), .B(n4112), .Z(n2080) );
  XOR U3442 ( .A(n2870), .B(n2080), .Z(out[132]) );
  XOR U3443 ( .A(in[36]), .B(n4276), .Z(n2289) );
  XOR U3444 ( .A(in[1158]), .B(n3315), .Z(n2643) );
  XNOR U3445 ( .A(in[1586]), .B(n3914), .Z(n2166) );
  IV U3446 ( .A(n2166), .Z(n2645) );
  OR U3447 ( .A(n2643), .B(n2645), .Z(n2081) );
  XNOR U3448 ( .A(n2289), .B(n2081), .Z(out[1330]) );
  XOR U3449 ( .A(in[37]), .B(n4278), .Z(n2291) );
  XOR U3450 ( .A(in[1159]), .B(n3318), .Z(n2647) );
  XOR U3451 ( .A(in[1587]), .B(n2574), .Z(n2649) );
  OR U3452 ( .A(n2647), .B(n2649), .Z(n2082) );
  XNOR U3453 ( .A(n2291), .B(n2082), .Z(out[1331]) );
  XOR U3454 ( .A(in[38]), .B(n4284), .Z(n2294) );
  XOR U3455 ( .A(in[1160]), .B(n3935), .Z(n2651) );
  XOR U3456 ( .A(in[1588]), .B(n2616), .Z(n2653) );
  OR U3457 ( .A(n2651), .B(n2653), .Z(n2083) );
  XNOR U3458 ( .A(n2294), .B(n2083), .Z(out[1332]) );
  XOR U3459 ( .A(in[39]), .B(n4286), .Z(n2296) );
  XOR U3460 ( .A(in[1161]), .B(n3942), .Z(n2655) );
  XOR U3461 ( .A(in[1589]), .B(n2658), .Z(n2657) );
  OR U3462 ( .A(n2655), .B(n2657), .Z(n2084) );
  XNOR U3463 ( .A(n2296), .B(n2084), .Z(out[1333]) );
  XOR U3464 ( .A(in[40]), .B(n4288), .Z(n2299) );
  XOR U3465 ( .A(in[1162]), .B(n3946), .Z(n2661) );
  XNOR U3466 ( .A(in[1590]), .B(n3065), .Z(n2663) );
  NANDN U3467 ( .A(n2661), .B(n2663), .Z(n2085) );
  XNOR U3468 ( .A(n2299), .B(n2085), .Z(out[1334]) );
  XOR U3469 ( .A(in[41]), .B(n4290), .Z(n2301) );
  XOR U3470 ( .A(in[1163]), .B(n3950), .Z(n2665) );
  XNOR U3471 ( .A(in[1591]), .B(n3067), .Z(n2667) );
  NANDN U3472 ( .A(n2665), .B(n2667), .Z(n2086) );
  XNOR U3473 ( .A(n2301), .B(n2086), .Z(out[1335]) );
  XOR U3474 ( .A(in[42]), .B(n4292), .Z(n2303) );
  XOR U3475 ( .A(in[1164]), .B(n3954), .Z(n2669) );
  XNOR U3476 ( .A(in[1592]), .B(n3070), .Z(n2671) );
  NANDN U3477 ( .A(n2669), .B(n2671), .Z(n2087) );
  XNOR U3478 ( .A(n2303), .B(n2087), .Z(out[1336]) );
  XOR U3479 ( .A(in[43]), .B(n4294), .Z(n2305) );
  XOR U3480 ( .A(in[1165]), .B(n3958), .Z(n2673) );
  XOR U3481 ( .A(in[1593]), .B(n2703), .Z(n2675) );
  OR U3482 ( .A(n2673), .B(n2675), .Z(n2088) );
  XNOR U3483 ( .A(n2305), .B(n2088), .Z(out[1337]) );
  XOR U3484 ( .A(in[44]), .B(n4296), .Z(n2307) );
  XOR U3485 ( .A(in[1166]), .B(n3962), .Z(n2677) );
  XOR U3486 ( .A(in[1594]), .B(n2705), .Z(n2679) );
  OR U3487 ( .A(n2677), .B(n2679), .Z(n2089) );
  XNOR U3488 ( .A(n2307), .B(n2089), .Z(out[1338]) );
  XOR U3489 ( .A(in[45]), .B(n4298), .Z(n2309) );
  XOR U3490 ( .A(in[1167]), .B(n3966), .Z(n2681) );
  XNOR U3491 ( .A(in[1595]), .B(n3953), .Z(n2174) );
  IV U3492 ( .A(n2174), .Z(n2683) );
  OR U3493 ( .A(n2681), .B(n2683), .Z(n2090) );
  XNOR U3494 ( .A(n2309), .B(n2090), .Z(out[1339]) );
  XOR U3495 ( .A(in[670]), .B(n4260), .Z(n2753) );
  IV U3496 ( .A(n2753), .Z(n2872) );
  XOR U3497 ( .A(in[604]), .B(n4096), .Z(n4159) );
  XNOR U3498 ( .A(in[195]), .B(n3306), .Z(n4156) );
  NANDN U3499 ( .A(n4159), .B(n4156), .Z(n2091) );
  XOR U3500 ( .A(n2872), .B(n2091), .Z(out[133]) );
  XOR U3501 ( .A(in[46]), .B(n4300), .Z(n2311) );
  XOR U3502 ( .A(in[1168]), .B(n3970), .Z(n2685) );
  XNOR U3503 ( .A(in[1596]), .B(n3957), .Z(n2176) );
  IV U3504 ( .A(n2176), .Z(n2687) );
  OR U3505 ( .A(n2685), .B(n2687), .Z(n2092) );
  XNOR U3506 ( .A(n2311), .B(n2092), .Z(out[1340]) );
  XOR U3507 ( .A(in[47]), .B(n4302), .Z(n2313) );
  XOR U3508 ( .A(in[1169]), .B(n3974), .Z(n2689) );
  XNOR U3509 ( .A(in[1597]), .B(n3961), .Z(n2178) );
  IV U3510 ( .A(n2178), .Z(n2691) );
  OR U3511 ( .A(n2689), .B(n2691), .Z(n2093) );
  XNOR U3512 ( .A(n2313), .B(n2093), .Z(out[1341]) );
  XOR U3513 ( .A(in[48]), .B(n4309), .Z(n2316) );
  XOR U3514 ( .A(in[1170]), .B(n3978), .Z(n2693) );
  XNOR U3515 ( .A(in[1598]), .B(n3965), .Z(n2180) );
  IV U3516 ( .A(n2180), .Z(n2695) );
  OR U3517 ( .A(n2693), .B(n2695), .Z(n2094) );
  XNOR U3518 ( .A(n2316), .B(n2094), .Z(out[1342]) );
  XOR U3519 ( .A(in[49]), .B(n4312), .Z(n2318) );
  XNOR U3520 ( .A(in[1171]), .B(n3985), .Z(n2697) );
  XNOR U3521 ( .A(in[1599]), .B(n3969), .Z(n2698) );
  NANDN U3522 ( .A(n2697), .B(n2698), .Z(n2095) );
  XNOR U3523 ( .A(n2318), .B(n2095), .Z(out[1343]) );
  XNOR U3524 ( .A(in[427]), .B(n4345), .Z(n2320) );
  NOR U3525 ( .A(n2441), .B(n2183), .Z(n2096) );
  XNOR U3526 ( .A(n2320), .B(n2096), .Z(out[1344]) );
  XNOR U3527 ( .A(in[428]), .B(n4348), .Z(n2322) );
  NOR U3528 ( .A(n2097), .B(n2185), .Z(n2098) );
  XNOR U3529 ( .A(n2322), .B(n2098), .Z(out[1345]) );
  XNOR U3530 ( .A(in[429]), .B(n4351), .Z(n2324) );
  NOR U3531 ( .A(n2447), .B(n2188), .Z(n2099) );
  XNOR U3532 ( .A(n2324), .B(n2099), .Z(out[1346]) );
  XNOR U3533 ( .A(in[430]), .B(n4354), .Z(n2326) );
  NOR U3534 ( .A(n2452), .B(n2190), .Z(n2100) );
  XNOR U3535 ( .A(n2326), .B(n2100), .Z(out[1347]) );
  XNOR U3536 ( .A(in[431]), .B(n4356), .Z(n2328) );
  NOR U3537 ( .A(n2101), .B(n2192), .Z(n2102) );
  XNOR U3538 ( .A(n2328), .B(n2102), .Z(out[1348]) );
  XNOR U3539 ( .A(in[432]), .B(n4359), .Z(n2330) );
  NOR U3540 ( .A(n2103), .B(n2194), .Z(n2104) );
  XNOR U3541 ( .A(n2330), .B(n2104), .Z(out[1349]) );
  XOR U3542 ( .A(in[671]), .B(n4261), .Z(n2755) );
  IV U3543 ( .A(n2755), .Z(n2874) );
  XOR U3544 ( .A(in[605]), .B(n4100), .Z(n4197) );
  XNOR U3545 ( .A(in[196]), .B(n3309), .Z(n4194) );
  NANDN U3546 ( .A(n4197), .B(n4194), .Z(n2105) );
  XOR U3547 ( .A(n2874), .B(n2105), .Z(out[134]) );
  XNOR U3548 ( .A(in[433]), .B(n4362), .Z(n2332) );
  NOR U3549 ( .A(n2464), .B(n2196), .Z(n2106) );
  XNOR U3550 ( .A(n2332), .B(n2106), .Z(out[1350]) );
  XNOR U3551 ( .A(in[434]), .B(n4365), .Z(n2334) );
  NOR U3552 ( .A(n2469), .B(n2198), .Z(n2107) );
  XNOR U3553 ( .A(n2334), .B(n2107), .Z(out[1351]) );
  XNOR U3554 ( .A(in[435]), .B(n4372), .Z(n2337) );
  NOR U3555 ( .A(n2470), .B(n2200), .Z(n2108) );
  XNOR U3556 ( .A(n2337), .B(n2108), .Z(out[1352]) );
  XNOR U3557 ( .A(in[436]), .B(n4375), .Z(n2340) );
  NOR U3558 ( .A(n2473), .B(n2202), .Z(n2109) );
  XNOR U3559 ( .A(n2340), .B(n2109), .Z(out[1353]) );
  XNOR U3560 ( .A(in[437]), .B(n4378), .Z(n2343) );
  NOR U3561 ( .A(n2476), .B(n2204), .Z(n2110) );
  XNOR U3562 ( .A(n2343), .B(n2110), .Z(out[1354]) );
  XNOR U3563 ( .A(in[438]), .B(n4381), .Z(n2346) );
  NOR U3564 ( .A(n2482), .B(n2206), .Z(n2111) );
  XNOR U3565 ( .A(n2346), .B(n2111), .Z(out[1355]) );
  XNOR U3566 ( .A(in[439]), .B(n4384), .Z(n2349) );
  NOR U3567 ( .A(n2483), .B(n2209), .Z(n2112) );
  XNOR U3568 ( .A(n2349), .B(n2112), .Z(out[1356]) );
  XNOR U3569 ( .A(in[440]), .B(n4386), .Z(n2352) );
  NOR U3570 ( .A(n2489), .B(n2211), .Z(n2113) );
  XNOR U3571 ( .A(n2352), .B(n2113), .Z(out[1357]) );
  XNOR U3572 ( .A(in[441]), .B(n4389), .Z(n2355) );
  XOR U3573 ( .A(in[442]), .B(n2114), .Z(n2357) );
  XOR U3574 ( .A(in[672]), .B(n4264), .Z(n2757) );
  IV U3575 ( .A(n2757), .Z(n2876) );
  XOR U3576 ( .A(in[606]), .B(n4104), .Z(n4215) );
  XNOR U3577 ( .A(in[197]), .B(n3312), .Z(n4442) );
  NANDN U3578 ( .A(n4215), .B(n4442), .Z(n2115) );
  XOR U3579 ( .A(n2876), .B(n2115), .Z(out[135]) );
  XOR U3580 ( .A(in[443]), .B(n2116), .Z(n2359) );
  XNOR U3581 ( .A(in[444]), .B(n4398), .Z(n2360) );
  NOR U3582 ( .A(n2117), .B(n2220), .Z(n2118) );
  XNOR U3583 ( .A(n2360), .B(n2118), .Z(out[1361]) );
  XNOR U3584 ( .A(in[445]), .B(n4405), .Z(n2363) );
  NOR U3585 ( .A(n2119), .B(n2222), .Z(n2120) );
  XNOR U3586 ( .A(n2363), .B(n2120), .Z(out[1362]) );
  XNOR U3587 ( .A(in[446]), .B(n4408), .Z(n2365) );
  XNOR U3588 ( .A(in[447]), .B(n4411), .Z(n2367) );
  NOR U3589 ( .A(n2121), .B(n2226), .Z(n2122) );
  XNOR U3590 ( .A(n2367), .B(n2122), .Z(out[1364]) );
  XNOR U3591 ( .A(in[384]), .B(n4414), .Z(n2369) );
  NOR U3592 ( .A(n2123), .B(n2228), .Z(n2124) );
  XNOR U3593 ( .A(n2369), .B(n2124), .Z(out[1365]) );
  XNOR U3594 ( .A(in[385]), .B(n4417), .Z(n2371) );
  XNOR U3595 ( .A(in[386]), .B(n4420), .Z(n2373) );
  XNOR U3596 ( .A(in[387]), .B(n4423), .Z(n2375) );
  NOR U3597 ( .A(n2125), .B(n2235), .Z(n2126) );
  XNOR U3598 ( .A(n2375), .B(n2126), .Z(out[1368]) );
  XNOR U3599 ( .A(in[388]), .B(n4426), .Z(n2377) );
  NOR U3600 ( .A(n2127), .B(n2237), .Z(n2128) );
  XNOR U3601 ( .A(n2377), .B(n2128), .Z(out[1369]) );
  XOR U3602 ( .A(in[673]), .B(n4267), .Z(n2764) );
  IV U3603 ( .A(n2764), .Z(n2878) );
  XOR U3604 ( .A(in[607]), .B(n4108), .Z(n4243) );
  XNOR U3605 ( .A(in[198]), .B(n3315), .Z(n4728) );
  NANDN U3606 ( .A(n4243), .B(n4728), .Z(n2129) );
  XOR U3607 ( .A(n2878), .B(n2129), .Z(out[136]) );
  XNOR U3608 ( .A(in[389]), .B(n4429), .Z(n2379) );
  XOR U3609 ( .A(in[390]), .B(n2130), .Z(n2381) );
  XNOR U3610 ( .A(in[391]), .B(n4443), .Z(n2384) );
  XNOR U3611 ( .A(in[392]), .B(n4446), .Z(n2386) );
  XNOR U3612 ( .A(in[393]), .B(n4449), .Z(n2388) );
  XNOR U3613 ( .A(in[394]), .B(n4452), .Z(n2390) );
  XNOR U3614 ( .A(in[395]), .B(n4455), .Z(n2392) );
  XNOR U3615 ( .A(n4458), .B(in[396]), .Z(n2394) );
  NOR U3616 ( .A(n2131), .B(n2254), .Z(n2132) );
  XOR U3617 ( .A(n2394), .B(n2132), .Z(out[1377]) );
  XNOR U3618 ( .A(n4461), .B(in[397]), .Z(n2395) );
  NOR U3619 ( .A(n2133), .B(n2256), .Z(n2134) );
  XOR U3620 ( .A(n2395), .B(n2134), .Z(out[1378]) );
  XNOR U3621 ( .A(n4464), .B(in[398]), .Z(n2396) );
  NOR U3622 ( .A(n2135), .B(n2258), .Z(n2136) );
  XOR U3623 ( .A(n2396), .B(n2136), .Z(out[1379]) );
  XOR U3624 ( .A(in[674]), .B(n4270), .Z(n2766) );
  IV U3625 ( .A(n2766), .Z(n2880) );
  XOR U3626 ( .A(in[608]), .B(n4116), .Z(n4257) );
  XNOR U3627 ( .A(in[199]), .B(n3318), .Z(n5156) );
  NANDN U3628 ( .A(n4257), .B(n5156), .Z(n2137) );
  XOR U3629 ( .A(n2880), .B(n2137), .Z(out[137]) );
  XNOR U3630 ( .A(n4467), .B(in[399]), .Z(n2397) );
  NOR U3631 ( .A(n2138), .B(n2260), .Z(n2139) );
  XOR U3632 ( .A(n2397), .B(n2139), .Z(out[1380]) );
  XNOR U3633 ( .A(n4470), .B(in[400]), .Z(n2398) );
  NOR U3634 ( .A(n2140), .B(n2262), .Z(n2141) );
  XOR U3635 ( .A(n2398), .B(n2141), .Z(out[1381]) );
  XNOR U3636 ( .A(n4477), .B(in[401]), .Z(n2400) );
  NOR U3637 ( .A(n2595), .B(n2264), .Z(n2142) );
  XOR U3638 ( .A(n2400), .B(n2142), .Z(out[1382]) );
  XNOR U3639 ( .A(n4480), .B(in[402]), .Z(n2401) );
  NOR U3640 ( .A(n2143), .B(n2266), .Z(n2144) );
  XOR U3641 ( .A(n2401), .B(n2144), .Z(out[1383]) );
  XNOR U3642 ( .A(n4483), .B(in[403]), .Z(n2402) );
  NOR U3643 ( .A(n2145), .B(n2268), .Z(n2146) );
  XOR U3644 ( .A(n2402), .B(n2146), .Z(out[1384]) );
  XNOR U3645 ( .A(in[404]), .B(n4486), .Z(n2403) );
  NOR U3646 ( .A(n2147), .B(n2270), .Z(n2148) );
  XOR U3647 ( .A(n2403), .B(n2148), .Z(out[1385]) );
  XNOR U3648 ( .A(in[405]), .B(n4489), .Z(n2404) );
  NOR U3649 ( .A(n2149), .B(n2273), .Z(n2150) );
  XOR U3650 ( .A(n2404), .B(n2150), .Z(out[1386]) );
  XNOR U3651 ( .A(in[406]), .B(n4492), .Z(n2405) );
  NOR U3652 ( .A(n2151), .B(n2275), .Z(n2152) );
  XOR U3653 ( .A(n2405), .B(n2152), .Z(out[1387]) );
  XNOR U3654 ( .A(in[407]), .B(n4495), .Z(n2406) );
  NOR U3655 ( .A(n2153), .B(n2277), .Z(n2154) );
  XOR U3656 ( .A(n2406), .B(n2154), .Z(out[1388]) );
  XNOR U3657 ( .A(in[408]), .B(n4498), .Z(n2407) );
  NOR U3658 ( .A(n2155), .B(n2279), .Z(n2156) );
  XOR U3659 ( .A(n2407), .B(n2156), .Z(out[1389]) );
  XOR U3660 ( .A(in[675]), .B(n4273), .Z(n2883) );
  IV U3661 ( .A(n3034), .Z(n4120) );
  XOR U3662 ( .A(in[609]), .B(n4120), .Z(n4283) );
  NANDN U3663 ( .A(n4283), .B(n4280), .Z(n2157) );
  XOR U3664 ( .A(n2883), .B(n2157), .Z(out[138]) );
  XNOR U3665 ( .A(in[409]), .B(n4501), .Z(n2408) );
  NOR U3666 ( .A(n2158), .B(n2281), .Z(n2159) );
  XOR U3667 ( .A(n2408), .B(n2159), .Z(out[1390]) );
  XNOR U3668 ( .A(in[410]), .B(n4504), .Z(n2409) );
  NOR U3669 ( .A(n2160), .B(n2283), .Z(n2161) );
  XOR U3670 ( .A(n2409), .B(n2161), .Z(out[1391]) );
  XOR U3671 ( .A(in[411]), .B(n4511), .Z(n2411) );
  NOR U3672 ( .A(n2162), .B(n2285), .Z(n2163) );
  XOR U3673 ( .A(n2411), .B(n2163), .Z(out[1392]) );
  XOR U3674 ( .A(in[412]), .B(n4514), .Z(n2412) );
  NOR U3675 ( .A(n2164), .B(n2287), .Z(n2165) );
  XOR U3676 ( .A(n2412), .B(n2165), .Z(out[1393]) );
  XOR U3677 ( .A(in[413]), .B(n4517), .Z(n2413) );
  NOR U3678 ( .A(n2166), .B(n2289), .Z(n2167) );
  XOR U3679 ( .A(n2413), .B(n2167), .Z(out[1394]) );
  XOR U3680 ( .A(in[414]), .B(n4520), .Z(n2414) );
  XOR U3681 ( .A(in[415]), .B(n4524), .Z(n2416) );
  XOR U3682 ( .A(in[416]), .B(n4528), .Z(n2418) );
  XNOR U3683 ( .A(in[417]), .B(n4532), .Z(n2420) );
  NOR U3684 ( .A(n2663), .B(n2299), .Z(n2168) );
  XOR U3685 ( .A(n2420), .B(n2168), .Z(out[1398]) );
  XNOR U3686 ( .A(in[418]), .B(n4536), .Z(n2421) );
  NOR U3687 ( .A(n2667), .B(n2301), .Z(n2169) );
  XOR U3688 ( .A(n2421), .B(n2169), .Z(out[1399]) );
  XOR U3689 ( .A(in[676]), .B(n4276), .Z(n2885) );
  IV U3690 ( .A(n2170), .Z(n4124) );
  XOR U3691 ( .A(in[610]), .B(n4124), .Z(n4308) );
  NANDN U3692 ( .A(n4308), .B(n4305), .Z(n2171) );
  XNOR U3693 ( .A(n2885), .B(n2171), .Z(out[139]) );
  XNOR U3694 ( .A(in[203]), .B(n3950), .Z(n4368) );
  XOR U3695 ( .A(in[1423]), .B(n3202), .Z(n4369) );
  XNOR U3696 ( .A(in[1046]), .B(n4492), .Z(n2890) );
  NANDN U3697 ( .A(n4369), .B(n2890), .Z(n2172) );
  XNOR U3698 ( .A(n4368), .B(n2172), .Z(out[13]) );
  XNOR U3699 ( .A(in[419]), .B(n4540), .Z(n2422) );
  NOR U3700 ( .A(n2671), .B(n2303), .Z(n2173) );
  XOR U3701 ( .A(n2422), .B(n2173), .Z(out[1400]) );
  XNOR U3702 ( .A(in[420]), .B(n4544), .Z(n2423) );
  XNOR U3703 ( .A(in[421]), .B(n4550), .Z(n2426) );
  XNOR U3704 ( .A(in[422]), .B(n4552), .Z(n2428) );
  NOR U3705 ( .A(n2174), .B(n2309), .Z(n2175) );
  XNOR U3706 ( .A(n2428), .B(n2175), .Z(out[1403]) );
  XNOR U3707 ( .A(in[423]), .B(n4333), .Z(n2430) );
  NOR U3708 ( .A(n2176), .B(n2311), .Z(n2177) );
  XNOR U3709 ( .A(n2430), .B(n2177), .Z(out[1404]) );
  XNOR U3710 ( .A(in[424]), .B(n4335), .Z(n2433) );
  NOR U3711 ( .A(n2178), .B(n2313), .Z(n2179) );
  XNOR U3712 ( .A(n2433), .B(n2179), .Z(out[1405]) );
  XNOR U3713 ( .A(in[425]), .B(n4341), .Z(n2435) );
  NOR U3714 ( .A(n2180), .B(n2316), .Z(n2181) );
  XNOR U3715 ( .A(n2435), .B(n2181), .Z(out[1406]) );
  XNOR U3716 ( .A(in[426]), .B(n4343), .Z(n2437) );
  NOR U3717 ( .A(n2698), .B(n2318), .Z(n2182) );
  XNOR U3718 ( .A(n2437), .B(n2182), .Z(out[1407]) );
  XOR U3719 ( .A(in[789]), .B(n4014), .Z(n2439) );
  NAND U3720 ( .A(n2183), .B(n2320), .Z(n2184) );
  XOR U3721 ( .A(n2439), .B(n2184), .Z(out[1408]) );
  IV U3722 ( .A(n2776), .Z(n4018) );
  XOR U3723 ( .A(in[790]), .B(n4018), .Z(n2442) );
  NAND U3724 ( .A(n2185), .B(n2322), .Z(n2186) );
  XOR U3725 ( .A(n2442), .B(n2186), .Z(out[1409]) );
  XOR U3726 ( .A(in[677]), .B(n4278), .Z(n2887) );
  IV U3727 ( .A(n3037), .Z(n4128) );
  XOR U3728 ( .A(in[611]), .B(n4128), .Z(n4340) );
  NANDN U3729 ( .A(n4340), .B(n4337), .Z(n2187) );
  XNOR U3730 ( .A(n2887), .B(n2187), .Z(out[140]) );
  IV U3731 ( .A(n2783), .Z(n4022) );
  XOR U3732 ( .A(in[791]), .B(n4022), .Z(n2448) );
  NAND U3733 ( .A(n2188), .B(n2324), .Z(n2189) );
  XOR U3734 ( .A(n2448), .B(n2189), .Z(out[1410]) );
  IV U3735 ( .A(n2797), .Z(n4030) );
  XOR U3736 ( .A(in[792]), .B(n4030), .Z(n2450) );
  NAND U3737 ( .A(n2190), .B(n2326), .Z(n2191) );
  XOR U3738 ( .A(n2450), .B(n2191), .Z(out[1411]) );
  IV U3739 ( .A(n2820), .Z(n4034) );
  XOR U3740 ( .A(in[793]), .B(n4034), .Z(n2456) );
  NAND U3741 ( .A(n2192), .B(n2328), .Z(n2193) );
  XOR U3742 ( .A(n2456), .B(n2193), .Z(out[1412]) );
  IV U3743 ( .A(n2843), .Z(n4038) );
  XOR U3744 ( .A(in[794]), .B(n4038), .Z(n2460) );
  NAND U3745 ( .A(n2194), .B(n2330), .Z(n2195) );
  XOR U3746 ( .A(n2460), .B(n2195), .Z(out[1413]) );
  IV U3747 ( .A(n2867), .Z(n4042) );
  XOR U3748 ( .A(in[795]), .B(n4042), .Z(n2465) );
  NAND U3749 ( .A(n2196), .B(n2332), .Z(n2197) );
  XOR U3750 ( .A(n2465), .B(n2197), .Z(out[1414]) );
  IV U3751 ( .A(n2891), .Z(n4046) );
  XOR U3752 ( .A(in[796]), .B(n4046), .Z(n2467) );
  NAND U3753 ( .A(n2198), .B(n2334), .Z(n2199) );
  XOR U3754 ( .A(n2467), .B(n2199), .Z(out[1415]) );
  IV U3755 ( .A(n2924), .Z(n4050) );
  XOR U3756 ( .A(in[797]), .B(n4050), .Z(n2471) );
  NAND U3757 ( .A(n2200), .B(n2337), .Z(n2201) );
  XOR U3758 ( .A(n2471), .B(n2201), .Z(out[1416]) );
  XOR U3759 ( .A(in[798]), .B(n4054), .Z(n2339) );
  NAND U3760 ( .A(n2202), .B(n2340), .Z(n2203) );
  XNOR U3761 ( .A(n2339), .B(n2203), .Z(out[1417]) );
  XOR U3762 ( .A(in[799]), .B(n4058), .Z(n2342) );
  NAND U3763 ( .A(n2204), .B(n2343), .Z(n2205) );
  XNOR U3764 ( .A(n2342), .B(n2205), .Z(out[1418]) );
  XOR U3765 ( .A(in[800]), .B(n4062), .Z(n2345) );
  NAND U3766 ( .A(n2206), .B(n2346), .Z(n2207) );
  XNOR U3767 ( .A(n2345), .B(n2207), .Z(out[1419]) );
  XOR U3768 ( .A(in[678]), .B(n4284), .Z(n2889) );
  IV U3769 ( .A(n3039), .Z(n4132) );
  XOR U3770 ( .A(in[612]), .B(n4132), .Z(n4371) );
  NANDN U3771 ( .A(n4371), .B(n4368), .Z(n2208) );
  XNOR U3772 ( .A(n2889), .B(n2208), .Z(out[141]) );
  XOR U3773 ( .A(in[801]), .B(n4066), .Z(n2348) );
  NAND U3774 ( .A(n2209), .B(n2349), .Z(n2210) );
  XNOR U3775 ( .A(n2348), .B(n2210), .Z(out[1420]) );
  XOR U3776 ( .A(in[802]), .B(n4074), .Z(n2351) );
  NAND U3777 ( .A(n2211), .B(n2352), .Z(n2212) );
  XNOR U3778 ( .A(n2351), .B(n2212), .Z(out[1421]) );
  XOR U3779 ( .A(in[803]), .B(n4078), .Z(n2354) );
  NAND U3780 ( .A(n2213), .B(n2355), .Z(n2214) );
  XNOR U3781 ( .A(n2354), .B(n2214), .Z(out[1422]) );
  XOR U3782 ( .A(in[804]), .B(n4082), .Z(n2358) );
  NANDN U3783 ( .A(n2357), .B(n2215), .Z(n2216) );
  XNOR U3784 ( .A(n2358), .B(n2216), .Z(out[1423]) );
  IV U3785 ( .A(n2217), .Z(n4086) );
  XOR U3786 ( .A(in[805]), .B(n4086), .Z(n2501) );
  NANDN U3787 ( .A(n2359), .B(n2218), .Z(n2219) );
  XOR U3788 ( .A(n2501), .B(n2219), .Z(out[1424]) );
  XNOR U3789 ( .A(in[806]), .B(n4089), .Z(n2504) );
  NAND U3790 ( .A(n2220), .B(n2360), .Z(n2221) );
  XNOR U3791 ( .A(n2504), .B(n2221), .Z(out[1425]) );
  XNOR U3792 ( .A(in[807]), .B(n4093), .Z(n2508) );
  NAND U3793 ( .A(n2222), .B(n2363), .Z(n2223) );
  XNOR U3794 ( .A(n2508), .B(n2223), .Z(out[1426]) );
  XNOR U3795 ( .A(in[808]), .B(n4097), .Z(n2512) );
  NAND U3796 ( .A(n2224), .B(n2365), .Z(n2225) );
  XNOR U3797 ( .A(n2512), .B(n2225), .Z(out[1427]) );
  XNOR U3798 ( .A(in[809]), .B(n4101), .Z(n2516) );
  NAND U3799 ( .A(n2226), .B(n2367), .Z(n2227) );
  XNOR U3800 ( .A(n2516), .B(n2227), .Z(out[1428]) );
  XNOR U3801 ( .A(in[810]), .B(n4105), .Z(n2520) );
  NAND U3802 ( .A(n2228), .B(n2369), .Z(n2229) );
  XNOR U3803 ( .A(n2520), .B(n2229), .Z(out[1429]) );
  XOR U3804 ( .A(in[679]), .B(n4286), .Z(n2772) );
  XOR U3805 ( .A(in[613]), .B(n4136), .Z(n4404) );
  XNOR U3806 ( .A(in[204]), .B(n3954), .Z(n4401) );
  NANDN U3807 ( .A(n4404), .B(n4401), .Z(n2230) );
  XNOR U3808 ( .A(n2772), .B(n2230), .Z(out[142]) );
  XNOR U3809 ( .A(in[811]), .B(n4109), .Z(n2524) );
  NAND U3810 ( .A(n2231), .B(n2371), .Z(n2232) );
  XOR U3811 ( .A(n2524), .B(n2232), .Z(out[1430]) );
  XNOR U3812 ( .A(in[812]), .B(n4117), .Z(n2528) );
  NAND U3813 ( .A(n2233), .B(n2373), .Z(n2234) );
  XOR U3814 ( .A(n2528), .B(n2234), .Z(out[1431]) );
  XOR U3815 ( .A(in[813]), .B(n4121), .Z(n2533) );
  NAND U3816 ( .A(n2235), .B(n2375), .Z(n2236) );
  XOR U3817 ( .A(n2533), .B(n2236), .Z(out[1432]) );
  XOR U3818 ( .A(in[814]), .B(n4125), .Z(n2537) );
  NAND U3819 ( .A(n2237), .B(n2377), .Z(n2238) );
  XOR U3820 ( .A(n2537), .B(n2238), .Z(out[1433]) );
  XOR U3821 ( .A(in[815]), .B(n4129), .Z(n2541) );
  NAND U3822 ( .A(n2239), .B(n2379), .Z(n2240) );
  XOR U3823 ( .A(n2541), .B(n2240), .Z(out[1434]) );
  XOR U3824 ( .A(in[816]), .B(n4133), .Z(n2545) );
  NANDN U3825 ( .A(n2381), .B(n2241), .Z(n2242) );
  XOR U3826 ( .A(n2545), .B(n2242), .Z(out[1435]) );
  XOR U3827 ( .A(in[817]), .B(n4137), .Z(n2549) );
  NAND U3828 ( .A(n2243), .B(n2384), .Z(n2244) );
  XOR U3829 ( .A(n2549), .B(n2244), .Z(out[1436]) );
  XOR U3830 ( .A(in[818]), .B(n4141), .Z(n2553) );
  NAND U3831 ( .A(n2245), .B(n2386), .Z(n2246) );
  XOR U3832 ( .A(n2553), .B(n2246), .Z(out[1437]) );
  XOR U3833 ( .A(in[819]), .B(n4145), .Z(n2557) );
  NAND U3834 ( .A(n2247), .B(n2388), .Z(n2248) );
  XOR U3835 ( .A(n2557), .B(n2248), .Z(out[1438]) );
  XOR U3836 ( .A(in[820]), .B(n4149), .Z(n2561) );
  NAND U3837 ( .A(n2249), .B(n2390), .Z(n2250) );
  XOR U3838 ( .A(n2561), .B(n2250), .Z(out[1439]) );
  XOR U3839 ( .A(in[680]), .B(n4288), .Z(n2773) );
  XOR U3840 ( .A(in[614]), .B(n4140), .Z(n4438) );
  XNOR U3841 ( .A(in[205]), .B(n3958), .Z(n4435) );
  NANDN U3842 ( .A(n4438), .B(n4435), .Z(n2251) );
  XNOR U3843 ( .A(n2773), .B(n2251), .Z(out[143]) );
  XNOR U3844 ( .A(in[821]), .B(n4153), .Z(n2566) );
  NAND U3845 ( .A(n2252), .B(n2392), .Z(n2253) );
  XOR U3846 ( .A(n2566), .B(n2253), .Z(out[1440]) );
  XNOR U3847 ( .A(in[822]), .B(n4163), .Z(n2570) );
  NANDN U3848 ( .A(n2394), .B(n2254), .Z(n2255) );
  XOR U3849 ( .A(n2570), .B(n2255), .Z(out[1441]) );
  XNOR U3850 ( .A(in[823]), .B(n4167), .Z(n2576) );
  NANDN U3851 ( .A(n2395), .B(n2256), .Z(n2257) );
  XOR U3852 ( .A(n2576), .B(n2257), .Z(out[1442]) );
  XNOR U3853 ( .A(in[824]), .B(n4171), .Z(n2580) );
  NANDN U3854 ( .A(n2396), .B(n2258), .Z(n2259) );
  XOR U3855 ( .A(n2580), .B(n2259), .Z(out[1443]) );
  XNOR U3856 ( .A(in[825]), .B(n4175), .Z(n2584) );
  NANDN U3857 ( .A(n2397), .B(n2260), .Z(n2261) );
  XOR U3858 ( .A(n2584), .B(n2261), .Z(out[1444]) );
  XOR U3859 ( .A(in[826]), .B(n3899), .Z(n2588) );
  NANDN U3860 ( .A(n2398), .B(n2262), .Z(n2263) );
  XOR U3861 ( .A(n2588), .B(n2263), .Z(out[1445]) );
  XOR U3862 ( .A(in[827]), .B(n3903), .Z(n2592) );
  NANDN U3863 ( .A(n2400), .B(n2264), .Z(n2265) );
  XOR U3864 ( .A(n2592), .B(n2265), .Z(out[1446]) );
  XOR U3865 ( .A(in[828]), .B(n3907), .Z(n2596) );
  NANDN U3866 ( .A(n2401), .B(n2266), .Z(n2267) );
  XOR U3867 ( .A(n2596), .B(n2267), .Z(out[1447]) );
  XOR U3868 ( .A(in[829]), .B(n3911), .Z(n2600) );
  NANDN U3869 ( .A(n2402), .B(n2268), .Z(n2269) );
  XOR U3870 ( .A(n2600), .B(n2269), .Z(out[1448]) );
  XOR U3871 ( .A(in[830]), .B(n3915), .Z(n2604) );
  NANDN U3872 ( .A(n2403), .B(n2270), .Z(n2271) );
  XOR U3873 ( .A(n2604), .B(n2271), .Z(out[1449]) );
  XOR U3874 ( .A(in[681]), .B(n4290), .Z(n2774) );
  XOR U3875 ( .A(in[615]), .B(n4144), .Z(n4476) );
  XNOR U3876 ( .A(in[206]), .B(n3962), .Z(n4473) );
  NANDN U3877 ( .A(n4476), .B(n4473), .Z(n2272) );
  XNOR U3878 ( .A(n2774), .B(n2272), .Z(out[144]) );
  XOR U3879 ( .A(in[831]), .B(n3919), .Z(n2608) );
  NANDN U3880 ( .A(n2404), .B(n2273), .Z(n2274) );
  XOR U3881 ( .A(n2608), .B(n2274), .Z(out[1450]) );
  XOR U3882 ( .A(in[768]), .B(n3923), .Z(n2612) );
  NANDN U3883 ( .A(n2405), .B(n2275), .Z(n2276) );
  XOR U3884 ( .A(n2612), .B(n2276), .Z(out[1451]) );
  XOR U3885 ( .A(in[769]), .B(n3927), .Z(n2618) );
  NANDN U3886 ( .A(n2406), .B(n2277), .Z(n2278) );
  XOR U3887 ( .A(n2618), .B(n2278), .Z(out[1452]) );
  XNOR U3888 ( .A(n3932), .B(in[770]), .Z(n2622) );
  NANDN U3889 ( .A(n2407), .B(n2279), .Z(n2280) );
  XNOR U3890 ( .A(n2622), .B(n2280), .Z(out[1453]) );
  IV U3891 ( .A(n3173), .Z(n3936) );
  XOR U3892 ( .A(n3936), .B(in[771]), .Z(n2626) );
  NANDN U3893 ( .A(n2408), .B(n2281), .Z(n2282) );
  XOR U3894 ( .A(n2626), .B(n2282), .Z(out[1454]) );
  IV U3895 ( .A(n3175), .Z(n3943) );
  XOR U3896 ( .A(n3943), .B(in[772]), .Z(n2630) );
  NANDN U3897 ( .A(n2409), .B(n2283), .Z(n2284) );
  XOR U3898 ( .A(n2630), .B(n2284), .Z(out[1455]) );
  IV U3899 ( .A(n3177), .Z(n3947) );
  XOR U3900 ( .A(n3947), .B(in[773]), .Z(n2634) );
  NANDN U3901 ( .A(n2411), .B(n2285), .Z(n2286) );
  XOR U3902 ( .A(n2634), .B(n2286), .Z(out[1456]) );
  IV U3903 ( .A(n3179), .Z(n3951) );
  XOR U3904 ( .A(n3951), .B(in[774]), .Z(n2638) );
  NANDN U3905 ( .A(n2412), .B(n2287), .Z(n2288) );
  XOR U3906 ( .A(n2638), .B(n2288), .Z(out[1457]) );
  IV U3907 ( .A(n3181), .Z(n3955) );
  XOR U3908 ( .A(n3955), .B(in[775]), .Z(n2642) );
  NANDN U3909 ( .A(n2413), .B(n2289), .Z(n2290) );
  XOR U3910 ( .A(n2642), .B(n2290), .Z(out[1458]) );
  IV U3911 ( .A(n3183), .Z(n3959) );
  XOR U3912 ( .A(n3959), .B(in[776]), .Z(n2646) );
  NAND U3913 ( .A(n2291), .B(n2414), .Z(n2292) );
  XOR U3914 ( .A(n2646), .B(n2292), .Z(out[1459]) );
  XOR U3915 ( .A(in[682]), .B(n4292), .Z(n2775) );
  XOR U3916 ( .A(in[616]), .B(n4148), .Z(n4510) );
  XNOR U3917 ( .A(in[207]), .B(n3966), .Z(n4507) );
  NANDN U3918 ( .A(n4510), .B(n4507), .Z(n2293) );
  XNOR U3919 ( .A(n2775), .B(n2293), .Z(out[145]) );
  IV U3920 ( .A(n3185), .Z(n3963) );
  XOR U3921 ( .A(in[777]), .B(n3963), .Z(n2650) );
  NAND U3922 ( .A(n2294), .B(n2416), .Z(n2295) );
  XOR U3923 ( .A(n2650), .B(n2295), .Z(out[1460]) );
  IV U3924 ( .A(n3187), .Z(n3967) );
  XOR U3925 ( .A(n3967), .B(in[778]), .Z(n2654) );
  NAND U3926 ( .A(n2296), .B(n2418), .Z(n2297) );
  XOR U3927 ( .A(n2654), .B(n2297), .Z(out[1461]) );
  IV U3928 ( .A(n2298), .Z(n3971) );
  XOR U3929 ( .A(n3971), .B(in[779]), .Z(n2660) );
  NANDN U3930 ( .A(n2420), .B(n2299), .Z(n2300) );
  XOR U3931 ( .A(n2660), .B(n2300), .Z(out[1462]) );
  IV U3932 ( .A(n3194), .Z(n3975) );
  XOR U3933 ( .A(in[780]), .B(n3975), .Z(n2664) );
  NANDN U3934 ( .A(n2421), .B(n2301), .Z(n2302) );
  XOR U3935 ( .A(n2664), .B(n2302), .Z(out[1463]) );
  IV U3936 ( .A(n3196), .Z(n3979) );
  XOR U3937 ( .A(in[781]), .B(n3979), .Z(n2668) );
  NANDN U3938 ( .A(n2422), .B(n2303), .Z(n2304) );
  XOR U3939 ( .A(n2668), .B(n2304), .Z(out[1464]) );
  IV U3940 ( .A(n3199), .Z(n3986) );
  XOR U3941 ( .A(in[782]), .B(n3986), .Z(n2672) );
  NAND U3942 ( .A(n2305), .B(n2423), .Z(n2306) );
  XOR U3943 ( .A(n2672), .B(n2306), .Z(out[1465]) );
  IV U3944 ( .A(n3202), .Z(n3990) );
  XOR U3945 ( .A(in[783]), .B(n3990), .Z(n2676) );
  NAND U3946 ( .A(n2307), .B(n2426), .Z(n2308) );
  XOR U3947 ( .A(n2676), .B(n2308), .Z(out[1466]) );
  IV U3948 ( .A(n3205), .Z(n3994) );
  XOR U3949 ( .A(in[784]), .B(n3994), .Z(n2680) );
  NAND U3950 ( .A(n2309), .B(n2428), .Z(n2310) );
  XOR U3951 ( .A(n2680), .B(n2310), .Z(out[1467]) );
  IV U3952 ( .A(n3208), .Z(n3998) );
  XOR U3953 ( .A(in[785]), .B(n3998), .Z(n2684) );
  NAND U3954 ( .A(n2311), .B(n2430), .Z(n2312) );
  XOR U3955 ( .A(n2684), .B(n2312), .Z(out[1468]) );
  XOR U3956 ( .A(in[786]), .B(n4002), .Z(n2432) );
  NAND U3957 ( .A(n2313), .B(n2433), .Z(n2314) );
  XNOR U3958 ( .A(n2432), .B(n2314), .Z(out[1469]) );
  XOR U3959 ( .A(in[683]), .B(n4294), .Z(n2779) );
  XOR U3960 ( .A(in[617]), .B(n4152), .Z(n4549) );
  XNOR U3961 ( .A(in[208]), .B(n3970), .Z(n4546) );
  NANDN U3962 ( .A(n4549), .B(n4546), .Z(n2315) );
  XNOR U3963 ( .A(n2779), .B(n2315), .Z(out[146]) );
  XOR U3964 ( .A(in[787]), .B(n4006), .Z(n2692) );
  NAND U3965 ( .A(n2316), .B(n2435), .Z(n2317) );
  XOR U3966 ( .A(n2692), .B(n2317), .Z(out[1470]) );
  XOR U3967 ( .A(in[788]), .B(n4010), .Z(n2696) );
  NAND U3968 ( .A(n2318), .B(n2437), .Z(n2319) );
  XOR U3969 ( .A(n2696), .B(n2319), .Z(out[1471]) );
  NANDN U3970 ( .A(n2320), .B(n2439), .Z(n2321) );
  XOR U3971 ( .A(n2440), .B(n2321), .Z(out[1472]) );
  NANDN U3972 ( .A(n2322), .B(n2442), .Z(n2323) );
  XOR U3973 ( .A(n2443), .B(n2323), .Z(out[1473]) );
  NANDN U3974 ( .A(n2324), .B(n2448), .Z(n2325) );
  XOR U3975 ( .A(n2449), .B(n2325), .Z(out[1474]) );
  NANDN U3976 ( .A(n2326), .B(n2450), .Z(n2327) );
  XOR U3977 ( .A(n2451), .B(n2327), .Z(out[1475]) );
  NANDN U3978 ( .A(n2328), .B(n2456), .Z(n2329) );
  XOR U3979 ( .A(n2457), .B(n2329), .Z(out[1476]) );
  NANDN U3980 ( .A(n2330), .B(n2460), .Z(n2331) );
  XOR U3981 ( .A(n2461), .B(n2331), .Z(out[1477]) );
  NANDN U3982 ( .A(n2332), .B(n2465), .Z(n2333) );
  XOR U3983 ( .A(n2466), .B(n2333), .Z(out[1478]) );
  NANDN U3984 ( .A(n2334), .B(n2467), .Z(n2335) );
  XOR U3985 ( .A(n2468), .B(n2335), .Z(out[1479]) );
  XNOR U3986 ( .A(in[684]), .B(n4296), .Z(n2910) );
  XOR U3987 ( .A(in[618]), .B(n4162), .Z(n4578) );
  XNOR U3988 ( .A(in[209]), .B(n3974), .Z(n4575) );
  NANDN U3989 ( .A(n4578), .B(n4575), .Z(n2336) );
  XOR U3990 ( .A(n2910), .B(n2336), .Z(out[147]) );
  NANDN U3991 ( .A(n2337), .B(n2471), .Z(n2338) );
  XOR U3992 ( .A(n2472), .B(n2338), .Z(out[1480]) );
  IV U3993 ( .A(n2339), .Z(n2474) );
  NANDN U3994 ( .A(n2340), .B(n2474), .Z(n2341) );
  XOR U3995 ( .A(n2475), .B(n2341), .Z(out[1481]) );
  IV U3996 ( .A(n2342), .Z(n2477) );
  NANDN U3997 ( .A(n2343), .B(n2477), .Z(n2344) );
  XOR U3998 ( .A(n2478), .B(n2344), .Z(out[1482]) );
  IV U3999 ( .A(n2345), .Z(n2479) );
  NANDN U4000 ( .A(n2346), .B(n2479), .Z(n2347) );
  XOR U4001 ( .A(n2480), .B(n2347), .Z(out[1483]) );
  IV U4002 ( .A(n2348), .Z(n2484) );
  NANDN U4003 ( .A(n2349), .B(n2484), .Z(n2350) );
  XOR U4004 ( .A(n2485), .B(n2350), .Z(out[1484]) );
  IV U4005 ( .A(n2351), .Z(n2486) );
  NANDN U4006 ( .A(n2352), .B(n2486), .Z(n2353) );
  XOR U4007 ( .A(n2487), .B(n2353), .Z(out[1485]) );
  IV U4008 ( .A(n2354), .Z(n2492) );
  NANDN U4009 ( .A(n2355), .B(n2492), .Z(n2356) );
  XNOR U4010 ( .A(n2491), .B(n2356), .Z(out[1486]) );
  IV U4011 ( .A(n2358), .Z(n2496) );
  OR U4012 ( .A(n2504), .B(n2360), .Z(n2361) );
  XOR U4013 ( .A(n2505), .B(n2361), .Z(out[1489]) );
  XNOR U4014 ( .A(in[685]), .B(n4298), .Z(n2913) );
  XOR U4015 ( .A(in[619]), .B(n4166), .Z(n4603) );
  XNOR U4016 ( .A(in[210]), .B(n3978), .Z(n4600) );
  NANDN U4017 ( .A(n4603), .B(n4600), .Z(n2362) );
  XOR U4018 ( .A(n2913), .B(n2362), .Z(out[148]) );
  OR U4019 ( .A(n2508), .B(n2363), .Z(n2364) );
  XOR U4020 ( .A(n2509), .B(n2364), .Z(out[1490]) );
  OR U4021 ( .A(n2512), .B(n2365), .Z(n2366) );
  XOR U4022 ( .A(n2513), .B(n2366), .Z(out[1491]) );
  OR U4023 ( .A(n2516), .B(n2367), .Z(n2368) );
  XOR U4024 ( .A(n2517), .B(n2368), .Z(out[1492]) );
  OR U4025 ( .A(n2520), .B(n2369), .Z(n2370) );
  XOR U4026 ( .A(n2521), .B(n2370), .Z(out[1493]) );
  NANDN U4027 ( .A(n2371), .B(n2524), .Z(n2372) );
  XOR U4028 ( .A(n2525), .B(n2372), .Z(out[1494]) );
  NANDN U4029 ( .A(n2373), .B(n2528), .Z(n2374) );
  XNOR U4030 ( .A(n2529), .B(n2374), .Z(out[1495]) );
  NANDN U4031 ( .A(n2375), .B(n2533), .Z(n2376) );
  XNOR U4032 ( .A(n2534), .B(n2376), .Z(out[1496]) );
  NANDN U4033 ( .A(n2377), .B(n2537), .Z(n2378) );
  XNOR U4034 ( .A(n2538), .B(n2378), .Z(out[1497]) );
  NANDN U4035 ( .A(n2379), .B(n2541), .Z(n2380) );
  XNOR U4036 ( .A(n2542), .B(n2380), .Z(out[1498]) );
  XOR U4037 ( .A(in[686]), .B(n4300), .Z(n2916) );
  XOR U4038 ( .A(in[620]), .B(n4170), .Z(n4628) );
  XOR U4039 ( .A(in[211]), .B(n3985), .Z(n4625) );
  NANDN U4040 ( .A(n4628), .B(n4625), .Z(n2382) );
  XNOR U4041 ( .A(n2916), .B(n2382), .Z(out[149]) );
  XOR U4042 ( .A(in[1424]), .B(n3205), .Z(n4402) );
  XNOR U4043 ( .A(in[1047]), .B(n4495), .Z(n2894) );
  NANDN U4044 ( .A(n4402), .B(n2894), .Z(n2383) );
  XNOR U4045 ( .A(n4401), .B(n2383), .Z(out[14]) );
  NANDN U4046 ( .A(n2384), .B(n2549), .Z(n2385) );
  XNOR U4047 ( .A(n2550), .B(n2385), .Z(out[1500]) );
  NANDN U4048 ( .A(n2386), .B(n2553), .Z(n2387) );
  XNOR U4049 ( .A(n2554), .B(n2387), .Z(out[1501]) );
  NANDN U4050 ( .A(n2388), .B(n2557), .Z(n2389) );
  XNOR U4051 ( .A(n2558), .B(n2389), .Z(out[1502]) );
  NANDN U4052 ( .A(n2390), .B(n2561), .Z(n2391) );
  XNOR U4053 ( .A(n2562), .B(n2391), .Z(out[1503]) );
  NANDN U4054 ( .A(n2392), .B(n2566), .Z(n2393) );
  XNOR U4055 ( .A(n2567), .B(n2393), .Z(out[1504]) );
  XOR U4056 ( .A(in[687]), .B(n4302), .Z(n2919) );
  XOR U4057 ( .A(in[621]), .B(n4174), .Z(n4658) );
  XOR U4058 ( .A(in[212]), .B(n3989), .Z(n4655) );
  NANDN U4059 ( .A(n4658), .B(n4655), .Z(n2399) );
  XNOR U4060 ( .A(n2919), .B(n2399), .Z(out[150]) );
  XOR U4061 ( .A(in[688]), .B(n4309), .Z(n2922) );
  XOR U4062 ( .A(in[213]), .B(n3993), .Z(n4670) );
  XNOR U4063 ( .A(in[622]), .B(n3898), .Z(n4672) );
  NANDN U4064 ( .A(n4670), .B(n4672), .Z(n2410) );
  XNOR U4065 ( .A(n2922), .B(n2410), .Z(out[151]) );
  NANDN U4066 ( .A(n2414), .B(n2646), .Z(n2415) );
  XOR U4067 ( .A(n2647), .B(n2415), .Z(out[1523]) );
  NANDN U4068 ( .A(n2416), .B(n2650), .Z(n2417) );
  XOR U4069 ( .A(n2651), .B(n2417), .Z(out[1524]) );
  NANDN U4070 ( .A(n2418), .B(n2654), .Z(n2419) );
  XOR U4071 ( .A(n2655), .B(n2419), .Z(out[1525]) );
  NANDN U4072 ( .A(n2423), .B(n2672), .Z(n2424) );
  XOR U4073 ( .A(n2673), .B(n2424), .Z(out[1529]) );
  XOR U4074 ( .A(in[689]), .B(n4312), .Z(n2928) );
  XOR U4075 ( .A(in[623]), .B(n3902), .Z(n4689) );
  XOR U4076 ( .A(in[214]), .B(n3997), .Z(n4686) );
  NANDN U4077 ( .A(n4689), .B(n4686), .Z(n2425) );
  XNOR U4078 ( .A(n2928), .B(n2425), .Z(out[152]) );
  NANDN U4079 ( .A(n2426), .B(n2676), .Z(n2427) );
  XOR U4080 ( .A(n2677), .B(n2427), .Z(out[1530]) );
  NANDN U4081 ( .A(n2428), .B(n2680), .Z(n2429) );
  XOR U4082 ( .A(n2681), .B(n2429), .Z(out[1531]) );
  NANDN U4083 ( .A(n2430), .B(n2684), .Z(n2431) );
  XOR U4084 ( .A(n2685), .B(n2431), .Z(out[1532]) );
  IV U4085 ( .A(n2432), .Z(n2688) );
  NANDN U4086 ( .A(n2433), .B(n2688), .Z(n2434) );
  XOR U4087 ( .A(n2689), .B(n2434), .Z(out[1533]) );
  NANDN U4088 ( .A(n2435), .B(n2692), .Z(n2436) );
  XOR U4089 ( .A(n2693), .B(n2436), .Z(out[1534]) );
  NANDN U4090 ( .A(n2437), .B(n2696), .Z(n2438) );
  XOR U4091 ( .A(n2697), .B(n2438), .Z(out[1535]) );
  ANDN U4092 ( .B(n2443), .A(n2442), .Z(n2446) );
  XNOR U4093 ( .A(n2444), .B(round_const[1]), .Z(n2445) );
  XNOR U4094 ( .A(n2446), .B(n2445), .Z(out[1537]) );
  ANDN U4095 ( .B(n2451), .A(n2450), .Z(n2454) );
  XOR U4096 ( .A(n2452), .B(round_const_3), .Z(n2453) );
  XNOR U4097 ( .A(n2454), .B(n2453), .Z(out[1539]) );
  XOR U4098 ( .A(in[690]), .B(n4315), .Z(n2931) );
  XOR U4099 ( .A(in[624]), .B(n3906), .Z(n4724) );
  XOR U4100 ( .A(in[215]), .B(n4001), .Z(n4721) );
  NANDN U4101 ( .A(n4724), .B(n4721), .Z(n2455) );
  XNOR U4102 ( .A(n2931), .B(n2455), .Z(out[153]) );
  ANDN U4103 ( .B(n2457), .A(n2456), .Z(n2458) );
  XOR U4104 ( .A(n2459), .B(n2458), .Z(out[1540]) );
  ANDN U4105 ( .B(n2461), .A(n2460), .Z(n2462) );
  XOR U4106 ( .A(n2463), .B(n2462), .Z(out[1541]) );
  ANDN U4107 ( .B(n2480), .A(n2479), .Z(n2481) );
  XNOR U4108 ( .A(n2482), .B(n2481), .Z(out[1547]) );
  ANDN U4109 ( .B(n2487), .A(n2486), .Z(n2488) );
  XNOR U4110 ( .A(n2489), .B(n2488), .Z(out[1549]) );
  XOR U4111 ( .A(in[691]), .B(n4318), .Z(n2934) );
  XOR U4112 ( .A(in[216]), .B(n4005), .Z(n4769) );
  XNOR U4113 ( .A(in[625]), .B(n3910), .Z(n4771) );
  NANDN U4114 ( .A(n4769), .B(n4771), .Z(n2490) );
  XNOR U4115 ( .A(n2934), .B(n2490), .Z(out[154]) );
  NOR U4116 ( .A(n2492), .B(n2491), .Z(n2493) );
  XOR U4117 ( .A(n2494), .B(n2493), .Z(out[1550]) );
  NOR U4118 ( .A(n2496), .B(n2495), .Z(n2499) );
  XNOR U4119 ( .A(n2497), .B(round_const_15), .Z(n2498) );
  XNOR U4120 ( .A(n2499), .B(n2498), .Z(out[1551]) );
  NOR U4121 ( .A(n2501), .B(n2500), .Z(n2502) );
  XOR U4122 ( .A(n2503), .B(n2502), .Z(out[1552]) );
  AND U4123 ( .A(n2505), .B(n2504), .Z(n2506) );
  XOR U4124 ( .A(n2507), .B(n2506), .Z(out[1553]) );
  AND U4125 ( .A(n2509), .B(n2508), .Z(n2510) );
  XOR U4126 ( .A(n2511), .B(n2510), .Z(out[1554]) );
  AND U4127 ( .A(n2513), .B(n2512), .Z(n2514) );
  XOR U4128 ( .A(n2515), .B(n2514), .Z(out[1555]) );
  AND U4129 ( .A(n2517), .B(n2516), .Z(n2518) );
  XOR U4130 ( .A(n2519), .B(n2518), .Z(out[1556]) );
  AND U4131 ( .A(n2521), .B(n2520), .Z(n2522) );
  XOR U4132 ( .A(n2523), .B(n2522), .Z(out[1557]) );
  ANDN U4133 ( .B(n2525), .A(n2524), .Z(n2526) );
  XOR U4134 ( .A(n2527), .B(n2526), .Z(out[1558]) );
  NOR U4135 ( .A(n2529), .B(n2528), .Z(n2530) );
  XOR U4136 ( .A(n2531), .B(n2530), .Z(out[1559]) );
  XOR U4137 ( .A(in[692]), .B(n4321), .Z(n2937) );
  XOR U4138 ( .A(in[217]), .B(n4009), .Z(n4812) );
  XNOR U4139 ( .A(in[626]), .B(n3914), .Z(n4814) );
  NANDN U4140 ( .A(n4812), .B(n4814), .Z(n2532) );
  XNOR U4141 ( .A(n2937), .B(n2532), .Z(out[155]) );
  NOR U4142 ( .A(n2534), .B(n2533), .Z(n2535) );
  XOR U4143 ( .A(n2536), .B(n2535), .Z(out[1560]) );
  NOR U4144 ( .A(n2538), .B(n2537), .Z(n2539) );
  XOR U4145 ( .A(n2540), .B(n2539), .Z(out[1561]) );
  NOR U4146 ( .A(n2542), .B(n2541), .Z(n2543) );
  XOR U4147 ( .A(n2544), .B(n2543), .Z(out[1562]) );
  NOR U4148 ( .A(n2546), .B(n2545), .Z(n2547) );
  XOR U4149 ( .A(n2548), .B(n2547), .Z(out[1563]) );
  NOR U4150 ( .A(n2550), .B(n2549), .Z(n2551) );
  XOR U4151 ( .A(n2552), .B(n2551), .Z(out[1564]) );
  NOR U4152 ( .A(n2554), .B(n2553), .Z(n2555) );
  XOR U4153 ( .A(n2556), .B(n2555), .Z(out[1565]) );
  NOR U4154 ( .A(n2558), .B(n2557), .Z(n2559) );
  XOR U4155 ( .A(n2560), .B(n2559), .Z(out[1566]) );
  NOR U4156 ( .A(n2562), .B(n2561), .Z(n2565) );
  XNOR U4157 ( .A(n2563), .B(round_const_31), .Z(n2564) );
  XNOR U4158 ( .A(n2565), .B(n2564), .Z(out[1567]) );
  NOR U4159 ( .A(n2567), .B(n2566), .Z(n2568) );
  XOR U4160 ( .A(n2569), .B(n2568), .Z(out[1568]) );
  NOR U4161 ( .A(n2571), .B(n2570), .Z(n2572) );
  XOR U4162 ( .A(n2573), .B(n2572), .Z(out[1569]) );
  XOR U4163 ( .A(in[693]), .B(n4324), .Z(n2939) );
  XNOR U4164 ( .A(in[218]), .B(n4013), .Z(n4856) );
  XNOR U4165 ( .A(in[627]), .B(n2574), .Z(n4858) );
  NANDN U4166 ( .A(n4856), .B(n4858), .Z(n2575) );
  XNOR U4167 ( .A(n2939), .B(n2575), .Z(out[156]) );
  NOR U4168 ( .A(n2577), .B(n2576), .Z(n2578) );
  XOR U4169 ( .A(n2579), .B(n2578), .Z(out[1570]) );
  NOR U4170 ( .A(n2581), .B(n2580), .Z(n2582) );
  XOR U4171 ( .A(n2583), .B(n2582), .Z(out[1571]) );
  NOR U4172 ( .A(n2585), .B(n2584), .Z(n2586) );
  XOR U4173 ( .A(n2587), .B(n2586), .Z(out[1572]) );
  NOR U4174 ( .A(n2589), .B(n2588), .Z(n2590) );
  XOR U4175 ( .A(n2591), .B(n2590), .Z(out[1573]) );
  NOR U4176 ( .A(n2593), .B(n2592), .Z(n2594) );
  XNOR U4177 ( .A(n2595), .B(n2594), .Z(out[1574]) );
  ANDN U4178 ( .B(n2597), .A(n2596), .Z(n2598) );
  XOR U4179 ( .A(n2599), .B(n2598), .Z(out[1575]) );
  ANDN U4180 ( .B(n2601), .A(n2600), .Z(n2602) );
  XOR U4181 ( .A(n2603), .B(n2602), .Z(out[1576]) );
  ANDN U4182 ( .B(n2605), .A(n2604), .Z(n2606) );
  XOR U4183 ( .A(n2607), .B(n2606), .Z(out[1577]) );
  NOR U4184 ( .A(n2609), .B(n2608), .Z(n2610) );
  XOR U4185 ( .A(n2611), .B(n2610), .Z(out[1578]) );
  ANDN U4186 ( .B(n2613), .A(n2612), .Z(n2614) );
  XOR U4187 ( .A(n2615), .B(n2614), .Z(out[1579]) );
  XOR U4188 ( .A(in[694]), .B(n4327), .Z(n2941) );
  XNOR U4189 ( .A(in[219]), .B(n4017), .Z(n4900) );
  XNOR U4190 ( .A(in[628]), .B(n2616), .Z(n4902) );
  NANDN U4191 ( .A(n4900), .B(n4902), .Z(n2617) );
  XNOR U4192 ( .A(n2941), .B(n2617), .Z(out[157]) );
  ANDN U4193 ( .B(n2619), .A(n2618), .Z(n2620) );
  XOR U4194 ( .A(n2621), .B(n2620), .Z(out[1580]) );
  AND U4195 ( .A(n2623), .B(n2622), .Z(n2624) );
  XOR U4196 ( .A(n2625), .B(n2624), .Z(out[1581]) );
  ANDN U4197 ( .B(n2627), .A(n2626), .Z(n2628) );
  XOR U4198 ( .A(n2629), .B(n2628), .Z(out[1582]) );
  ANDN U4199 ( .B(n2631), .A(n2630), .Z(n2632) );
  XOR U4200 ( .A(n2633), .B(n2632), .Z(out[1583]) );
  ANDN U4201 ( .B(n2635), .A(n2634), .Z(n2636) );
  XOR U4202 ( .A(n2637), .B(n2636), .Z(out[1584]) );
  ANDN U4203 ( .B(n2639), .A(n2638), .Z(n2640) );
  XOR U4204 ( .A(n2641), .B(n2640), .Z(out[1585]) );
  ANDN U4205 ( .B(n2643), .A(n2642), .Z(n2644) );
  XOR U4206 ( .A(n2645), .B(n2644), .Z(out[1586]) );
  ANDN U4207 ( .B(n2647), .A(n2646), .Z(n2648) );
  XOR U4208 ( .A(n2649), .B(n2648), .Z(out[1587]) );
  ANDN U4209 ( .B(n2651), .A(n2650), .Z(n2652) );
  XOR U4210 ( .A(n2653), .B(n2652), .Z(out[1588]) );
  ANDN U4211 ( .B(n2655), .A(n2654), .Z(n2656) );
  XOR U4212 ( .A(n2657), .B(n2656), .Z(out[1589]) );
  XOR U4213 ( .A(in[695]), .B(n4330), .Z(n2943) );
  XNOR U4214 ( .A(in[220]), .B(n4021), .Z(n4944) );
  XNOR U4215 ( .A(in[629]), .B(n2658), .Z(n4946) );
  NANDN U4216 ( .A(n4944), .B(n4946), .Z(n2659) );
  XNOR U4217 ( .A(n2943), .B(n2659), .Z(out[158]) );
  ANDN U4218 ( .B(n2661), .A(n2660), .Z(n2662) );
  XNOR U4219 ( .A(n2663), .B(n2662), .Z(out[1590]) );
  ANDN U4220 ( .B(n2665), .A(n2664), .Z(n2666) );
  XNOR U4221 ( .A(n2667), .B(n2666), .Z(out[1591]) );
  ANDN U4222 ( .B(n2669), .A(n2668), .Z(n2670) );
  XNOR U4223 ( .A(n2671), .B(n2670), .Z(out[1592]) );
  ANDN U4224 ( .B(n2673), .A(n2672), .Z(n2674) );
  XOR U4225 ( .A(n2675), .B(n2674), .Z(out[1593]) );
  ANDN U4226 ( .B(n2677), .A(n2676), .Z(n2678) );
  XOR U4227 ( .A(n2679), .B(n2678), .Z(out[1594]) );
  ANDN U4228 ( .B(n2681), .A(n2680), .Z(n2682) );
  XOR U4229 ( .A(n2683), .B(n2682), .Z(out[1595]) );
  ANDN U4230 ( .B(n2685), .A(n2684), .Z(n2686) );
  XOR U4231 ( .A(n2687), .B(n2686), .Z(out[1596]) );
  ANDN U4232 ( .B(n2689), .A(n2688), .Z(n2690) );
  XOR U4233 ( .A(n2691), .B(n2690), .Z(out[1597]) );
  ANDN U4234 ( .B(n2693), .A(n2692), .Z(n2694) );
  XOR U4235 ( .A(n2695), .B(n2694), .Z(out[1598]) );
  XOR U4236 ( .A(in[696]), .B(n4178), .Z(n2945) );
  XNOR U4237 ( .A(in[221]), .B(n4029), .Z(n4988) );
  XNOR U4238 ( .A(in[630]), .B(n3065), .Z(n4990) );
  NANDN U4239 ( .A(n4988), .B(n4990), .Z(n2699) );
  XNOR U4240 ( .A(n2945), .B(n2699), .Z(out[159]) );
  XOR U4241 ( .A(in[1425]), .B(n3208), .Z(n4436) );
  XNOR U4242 ( .A(in[1048]), .B(n4498), .Z(n2897) );
  NANDN U4243 ( .A(n4436), .B(n2897), .Z(n2700) );
  XNOR U4244 ( .A(n4435), .B(n2700), .Z(out[15]) );
  XOR U4245 ( .A(in[697]), .B(n4181), .Z(n2947) );
  XNOR U4246 ( .A(in[222]), .B(n4033), .Z(n5032) );
  XNOR U4247 ( .A(in[631]), .B(n3067), .Z(n5034) );
  NANDN U4248 ( .A(n5032), .B(n5034), .Z(n2701) );
  XNOR U4249 ( .A(n2947), .B(n2701), .Z(out[160]) );
  XOR U4250 ( .A(in[698]), .B(n4184), .Z(n2949) );
  XNOR U4251 ( .A(in[223]), .B(n4037), .Z(n5073) );
  XNOR U4252 ( .A(in[632]), .B(n3070), .Z(n5075) );
  NANDN U4253 ( .A(n5073), .B(n5075), .Z(n2702) );
  XNOR U4254 ( .A(n2949), .B(n2702), .Z(out[161]) );
  XOR U4255 ( .A(in[699]), .B(n4187), .Z(n2953) );
  XNOR U4256 ( .A(in[633]), .B(n2703), .Z(n5110) );
  XOR U4257 ( .A(in[224]), .B(n4041), .Z(n5107) );
  NAND U4258 ( .A(n5110), .B(n5107), .Z(n2704) );
  XNOR U4259 ( .A(n2953), .B(n2704), .Z(out[162]) );
  XOR U4260 ( .A(in[700]), .B(n4190), .Z(n2955) );
  XNOR U4261 ( .A(in[634]), .B(n2705), .Z(n5152) );
  XOR U4262 ( .A(in[225]), .B(n4045), .Z(n5149) );
  NAND U4263 ( .A(n5152), .B(n5149), .Z(n2706) );
  XOR U4264 ( .A(n2955), .B(n2706), .Z(out[163]) );
  XOR U4265 ( .A(in[701]), .B(n4193), .Z(n2957) );
  ANDN U4266 ( .B(n3117), .A(n2707), .Z(n2708) );
  XNOR U4267 ( .A(n2957), .B(n2708), .Z(out[164]) );
  XOR U4268 ( .A(in[702]), .B(n4198), .Z(n2959) );
  ANDN U4269 ( .B(n3137), .A(n2709), .Z(n2710) );
  XNOR U4270 ( .A(n2959), .B(n2710), .Z(out[165]) );
  XNOR U4271 ( .A(in[703]), .B(n4199), .Z(n2961) );
  ANDN U4272 ( .B(n3156), .A(n2711), .Z(n2712) );
  XNOR U4273 ( .A(n2961), .B(n2712), .Z(out[166]) );
  XOR U4274 ( .A(in[640]), .B(n4200), .Z(n2963) );
  ANDN U4275 ( .B(n3167), .A(n2713), .Z(n2714) );
  XNOR U4276 ( .A(n2963), .B(n2714), .Z(out[167]) );
  XOR U4277 ( .A(in[641]), .B(n4201), .Z(n2965) );
  NOR U4278 ( .A(n2715), .B(n3192), .Z(n2716) );
  XNOR U4279 ( .A(n2965), .B(n2716), .Z(out[168]) );
  XOR U4280 ( .A(in[642]), .B(n4202), .Z(n2967) );
  NOR U4281 ( .A(n2717), .B(n3222), .Z(n2718) );
  XNOR U4282 ( .A(n2967), .B(n2718), .Z(out[169]) );
  XOR U4283 ( .A(in[1426]), .B(n4002), .Z(n4474) );
  XNOR U4284 ( .A(in[1049]), .B(n4501), .Z(n2900) );
  NANDN U4285 ( .A(n4474), .B(n2900), .Z(n2719) );
  XNOR U4286 ( .A(n4473), .B(n2719), .Z(out[16]) );
  XOR U4287 ( .A(in[643]), .B(n4203), .Z(n2969) );
  NOR U4288 ( .A(n2720), .B(n3246), .Z(n2721) );
  XNOR U4289 ( .A(n2969), .B(n2721), .Z(out[170]) );
  XOR U4290 ( .A(in[644]), .B(n4204), .Z(n2971) );
  NOR U4291 ( .A(n2722), .B(n3258), .Z(n2723) );
  XNOR U4292 ( .A(n2971), .B(n2723), .Z(out[171]) );
  XOR U4293 ( .A(in[645]), .B(n4205), .Z(n2977) );
  NOR U4294 ( .A(n2724), .B(n3268), .Z(n2725) );
  XNOR U4295 ( .A(n2977), .B(n2725), .Z(out[172]) );
  XOR U4296 ( .A(in[646]), .B(n4208), .Z(n2979) );
  NOR U4297 ( .A(n3302), .B(n2814), .Z(n2726) );
  XNOR U4298 ( .A(n2979), .B(n2726), .Z(out[173]) );
  XOR U4299 ( .A(in[647]), .B(n4211), .Z(n2981) );
  NOR U4300 ( .A(n3332), .B(n2816), .Z(n2727) );
  XNOR U4301 ( .A(n2981), .B(n2727), .Z(out[174]) );
  XNOR U4302 ( .A(in[648]), .B(n4216), .Z(n2983) );
  NOR U4303 ( .A(n3360), .B(n2818), .Z(n2728) );
  XNOR U4304 ( .A(n2983), .B(n2728), .Z(out[175]) );
  XOR U4305 ( .A(in[649]), .B(n4219), .Z(n2985) );
  NOR U4306 ( .A(n3388), .B(n2823), .Z(n2729) );
  XNOR U4307 ( .A(n2985), .B(n2729), .Z(out[176]) );
  XOR U4308 ( .A(in[650]), .B(n3090), .Z(n2987) );
  NOR U4309 ( .A(n3423), .B(n2825), .Z(n2730) );
  XOR U4310 ( .A(n2987), .B(n2730), .Z(out[177]) );
  IV U4311 ( .A(n3092), .Z(n4225) );
  XOR U4312 ( .A(in[651]), .B(n4225), .Z(n2988) );
  NOR U4313 ( .A(n3458), .B(n2827), .Z(n2731) );
  XNOR U4314 ( .A(n2988), .B(n2731), .Z(out[178]) );
  IV U4315 ( .A(n3094), .Z(n4228) );
  XOR U4316 ( .A(in[652]), .B(n4228), .Z(n2990) );
  NOR U4317 ( .A(n3480), .B(n2829), .Z(n2732) );
  XNOR U4318 ( .A(n2990), .B(n2732), .Z(out[179]) );
  XOR U4319 ( .A(in[1427]), .B(n3213), .Z(n4508) );
  XNOR U4320 ( .A(in[1050]), .B(n4504), .Z(n2903) );
  NANDN U4321 ( .A(n4508), .B(n2903), .Z(n2733) );
  XNOR U4322 ( .A(n4507), .B(n2733), .Z(out[17]) );
  IV U4323 ( .A(n3098), .Z(n4231) );
  XOR U4324 ( .A(in[653]), .B(n4231), .Z(n2992) );
  NOR U4325 ( .A(n3502), .B(n2831), .Z(n2734) );
  XNOR U4326 ( .A(n2992), .B(n2734), .Z(out[180]) );
  IV U4327 ( .A(n3100), .Z(n4234) );
  XOR U4328 ( .A(in[654]), .B(n4234), .Z(n2994) );
  NOR U4329 ( .A(n3517), .B(n2833), .Z(n2735) );
  XNOR U4330 ( .A(n2994), .B(n2735), .Z(out[181]) );
  XNOR U4331 ( .A(in[655]), .B(n4237), .Z(n2999) );
  NOR U4332 ( .A(n3547), .B(n2835), .Z(n2736) );
  XNOR U4333 ( .A(n2999), .B(n2736), .Z(out[182]) );
  IV U4334 ( .A(n3103), .Z(n4238) );
  XOR U4335 ( .A(in[656]), .B(n4238), .Z(n3001) );
  NOR U4336 ( .A(n3577), .B(n2837), .Z(n2737) );
  XNOR U4337 ( .A(n3001), .B(n2737), .Z(out[183]) );
  XOR U4338 ( .A(in[657]), .B(n4239), .Z(n3003) );
  NOR U4339 ( .A(n3601), .B(n2839), .Z(n2738) );
  XNOR U4340 ( .A(n3003), .B(n2738), .Z(out[184]) );
  IV U4341 ( .A(n3107), .Z(n4244) );
  XOR U4342 ( .A(in[658]), .B(n4244), .Z(n3005) );
  NOR U4343 ( .A(n3631), .B(n2841), .Z(n2739) );
  XNOR U4344 ( .A(n3005), .B(n2739), .Z(out[185]) );
  IV U4345 ( .A(n3109), .Z(n4247) );
  XOR U4346 ( .A(in[659]), .B(n4247), .Z(n3007) );
  NOR U4347 ( .A(n3675), .B(n2846), .Z(n2740) );
  XNOR U4348 ( .A(n3007), .B(n2740), .Z(out[186]) );
  XOR U4349 ( .A(in[660]), .B(n4248), .Z(n3009) );
  NOR U4350 ( .A(n3719), .B(n2848), .Z(n2741) );
  XOR U4351 ( .A(n3009), .B(n2741), .Z(out[187]) );
  XOR U4352 ( .A(in[661]), .B(n4249), .Z(n3012) );
  NOR U4353 ( .A(n3765), .B(n2850), .Z(n2742) );
  XOR U4354 ( .A(n3012), .B(n2742), .Z(out[188]) );
  XOR U4355 ( .A(in[662]), .B(n4250), .Z(n3015) );
  XOR U4356 ( .A(in[1428]), .B(n3216), .Z(n4547) );
  XNOR U4357 ( .A(in[1051]), .B(n2743), .Z(n2906) );
  NANDN U4358 ( .A(n4547), .B(n2906), .Z(n2744) );
  XNOR U4359 ( .A(n4546), .B(n2744), .Z(out[18]) );
  XOR U4360 ( .A(in[663]), .B(n4251), .Z(n3016) );
  XOR U4361 ( .A(in[664]), .B(n4252), .Z(n3019) );
  NANDN U4362 ( .A(n2858), .B(n3940), .Z(n2745) );
  XOR U4363 ( .A(n2859), .B(n2745), .Z(out[192]) );
  XNOR U4364 ( .A(in[1034]), .B(n4452), .Z(n2762) );
  ANDN U4365 ( .B(n3983), .A(n2861), .Z(n2746) );
  XNOR U4366 ( .A(n2762), .B(n2746), .Z(out[193]) );
  XNOR U4367 ( .A(in[1035]), .B(n4455), .Z(n2975) );
  ANDN U4368 ( .B(n4027), .A(n2747), .Z(n2748) );
  XNOR U4369 ( .A(n2975), .B(n2748), .Z(out[194]) );
  XOR U4370 ( .A(n4458), .B(in[1036]), .Z(n3168) );
  ANDN U4371 ( .B(n4071), .A(n2749), .Z(n2750) );
  XNOR U4372 ( .A(n3168), .B(n2750), .Z(out[195]) );
  XOR U4373 ( .A(n4461), .B(in[1037]), .Z(n3424) );
  ANDN U4374 ( .B(n4115), .A(n2751), .Z(n2752) );
  XNOR U4375 ( .A(n3424), .B(n2752), .Z(out[196]) );
  XOR U4376 ( .A(n4464), .B(in[1038]), .Z(n3720) );
  ANDN U4377 ( .B(n4159), .A(n2753), .Z(n2754) );
  XNOR U4378 ( .A(n3720), .B(n2754), .Z(out[197]) );
  XOR U4379 ( .A(n4467), .B(in[1039]), .Z(n4160) );
  ANDN U4380 ( .B(n4197), .A(n2755), .Z(n2756) );
  XNOR U4381 ( .A(n4160), .B(n2756), .Z(out[198]) );
  XOR U4382 ( .A(n4470), .B(in[1040]), .Z(n4439) );
  ANDN U4383 ( .B(n4215), .A(n2757), .Z(n2758) );
  XNOR U4384 ( .A(n4439), .B(n2758), .Z(out[199]) );
  XOR U4385 ( .A(in[1429]), .B(n2759), .Z(n4576) );
  XNOR U4386 ( .A(in[1052]), .B(n2760), .Z(n2909) );
  NANDN U4387 ( .A(n4576), .B(n2909), .Z(n2761) );
  XNOR U4388 ( .A(n4575), .B(n2761), .Z(out[19]) );
  XOR U4389 ( .A(n3173), .B(in[1411]), .Z(n3981) );
  IV U4390 ( .A(n2762), .Z(n2860) );
  NANDN U4391 ( .A(n3981), .B(n2860), .Z(n2763) );
  XNOR U4392 ( .A(n3982), .B(n2763), .Z(out[1]) );
  XOR U4393 ( .A(n4477), .B(in[1041]), .Z(n4725) );
  ANDN U4394 ( .B(n4243), .A(n2764), .Z(n2765) );
  XNOR U4395 ( .A(n4725), .B(n2765), .Z(out[200]) );
  XOR U4396 ( .A(n4480), .B(in[1042]), .Z(n5153) );
  ANDN U4397 ( .B(n4257), .A(n2766), .Z(n2767) );
  XNOR U4398 ( .A(n5153), .B(n2767), .Z(out[201]) );
  NAND U4399 ( .A(n4283), .B(n2883), .Z(n2768) );
  XNOR U4400 ( .A(n2882), .B(n2768), .Z(out[202]) );
  NANDN U4401 ( .A(n2885), .B(n4308), .Z(n2769) );
  XNOR U4402 ( .A(n2886), .B(n2769), .Z(out[203]) );
  NANDN U4403 ( .A(n2887), .B(n4340), .Z(n2770) );
  XNOR U4404 ( .A(n2888), .B(n2770), .Z(out[204]) );
  NANDN U4405 ( .A(n2889), .B(n4371), .Z(n2771) );
  XNOR U4406 ( .A(n2890), .B(n2771), .Z(out[205]) );
  IV U4407 ( .A(n2772), .Z(n2895) );
  IV U4408 ( .A(n2773), .Z(n2898) );
  IV U4409 ( .A(n2774), .Z(n2901) );
  IV U4410 ( .A(n2775), .Z(n2904) );
  XOR U4411 ( .A(in[1430]), .B(n2776), .Z(n4601) );
  XNOR U4412 ( .A(in[1053]), .B(n2777), .Z(n2912) );
  NANDN U4413 ( .A(n4601), .B(n2912), .Z(n2778) );
  XNOR U4414 ( .A(n4600), .B(n2778), .Z(out[20]) );
  IV U4415 ( .A(n2779), .Z(n2907) );
  XOR U4416 ( .A(in[1054]), .B(n4520), .Z(n2784) );
  IV U4417 ( .A(n2784), .Z(n2915) );
  XOR U4418 ( .A(in[1055]), .B(n4524), .Z(n2798) );
  IV U4419 ( .A(n2798), .Z(n2918) );
  XOR U4420 ( .A(in[1056]), .B(n4528), .Z(n2821) );
  IV U4421 ( .A(n2821), .Z(n2921) );
  NOR U4422 ( .A(n4672), .B(n2922), .Z(n2780) );
  XOR U4423 ( .A(n2921), .B(n2780), .Z(out[215]) );
  XOR U4424 ( .A(in[1057]), .B(n4532), .Z(n2844) );
  IV U4425 ( .A(n2844), .Z(n2927) );
  XOR U4426 ( .A(in[1058]), .B(n4536), .Z(n2868) );
  IV U4427 ( .A(n2868), .Z(n2930) );
  XOR U4428 ( .A(in[1059]), .B(n4540), .Z(n2892) );
  IV U4429 ( .A(n2892), .Z(n2933) );
  NOR U4430 ( .A(n4771), .B(n2934), .Z(n2781) );
  XOR U4431 ( .A(n2933), .B(n2781), .Z(out[218]) );
  XNOR U4432 ( .A(in[1060]), .B(n4544), .Z(n2925) );
  IV U4433 ( .A(n2925), .Z(n2936) );
  NOR U4434 ( .A(n4814), .B(n2937), .Z(n2782) );
  XOR U4435 ( .A(n2936), .B(n2782), .Z(out[219]) );
  XOR U4436 ( .A(in[1431]), .B(n2783), .Z(n4626) );
  OR U4437 ( .A(n4626), .B(n2784), .Z(n2785) );
  XNOR U4438 ( .A(n4625), .B(n2785), .Z(out[21]) );
  XNOR U4439 ( .A(in[1061]), .B(n4550), .Z(n2951) );
  NOR U4440 ( .A(n4858), .B(n2939), .Z(n2786) );
  XNOR U4441 ( .A(n2951), .B(n2786), .Z(out[220]) );
  XNOR U4442 ( .A(in[1062]), .B(n4552), .Z(n2973) );
  NOR U4443 ( .A(n4902), .B(n2941), .Z(n2787) );
  XNOR U4444 ( .A(n2973), .B(n2787), .Z(out[221]) );
  XNOR U4445 ( .A(in[1063]), .B(n4333), .Z(n2996) );
  NOR U4446 ( .A(n4946), .B(n2943), .Z(n2788) );
  XNOR U4447 ( .A(n2996), .B(n2788), .Z(out[222]) );
  XNOR U4448 ( .A(in[1064]), .B(n4335), .Z(n3022) );
  NOR U4449 ( .A(n4990), .B(n2945), .Z(n2789) );
  XNOR U4450 ( .A(n3022), .B(n2789), .Z(out[223]) );
  XNOR U4451 ( .A(in[1065]), .B(n4341), .Z(n3042) );
  NOR U4452 ( .A(n5034), .B(n2947), .Z(n2790) );
  XNOR U4453 ( .A(n3042), .B(n2790), .Z(out[224]) );
  XNOR U4454 ( .A(in[1066]), .B(n4343), .Z(n3054) );
  NOR U4455 ( .A(n5075), .B(n2949), .Z(n2791) );
  XNOR U4456 ( .A(n3054), .B(n2791), .Z(out[225]) );
  XNOR U4457 ( .A(in[1067]), .B(n4345), .Z(n3075) );
  NOR U4458 ( .A(n5110), .B(n2953), .Z(n2792) );
  XNOR U4459 ( .A(n3075), .B(n2792), .Z(out[226]) );
  XNOR U4460 ( .A(in[1068]), .B(n4348), .Z(n3096) );
  XOR U4461 ( .A(in[1069]), .B(n4351), .Z(n3115) );
  NANDN U4462 ( .A(n2793), .B(n2957), .Z(n2794) );
  XNOR U4463 ( .A(n3115), .B(n2794), .Z(out[228]) );
  XOR U4464 ( .A(in[1070]), .B(n4354), .Z(n3135) );
  NANDN U4465 ( .A(n2795), .B(n2959), .Z(n2796) );
  XNOR U4466 ( .A(n3135), .B(n2796), .Z(out[229]) );
  XOR U4467 ( .A(in[1432]), .B(n2797), .Z(n4656) );
  OR U4468 ( .A(n4656), .B(n2798), .Z(n2799) );
  XNOR U4469 ( .A(n4655), .B(n2799), .Z(out[22]) );
  XNOR U4470 ( .A(in[1071]), .B(n4356), .Z(n3153) );
  NANDN U4471 ( .A(n2800), .B(n2961), .Z(n2801) );
  XOR U4472 ( .A(n3153), .B(n2801), .Z(out[230]) );
  XOR U4473 ( .A(in[1072]), .B(n4359), .Z(n3165) );
  NANDN U4474 ( .A(n2802), .B(n2963), .Z(n2803) );
  XNOR U4475 ( .A(n3165), .B(n2803), .Z(out[231]) );
  XOR U4476 ( .A(in[1073]), .B(n4362), .Z(n3190) );
  NANDN U4477 ( .A(n2804), .B(n2965), .Z(n2805) );
  XNOR U4478 ( .A(n3190), .B(n2805), .Z(out[232]) );
  XOR U4479 ( .A(in[1074]), .B(n4365), .Z(n3219) );
  NANDN U4480 ( .A(n2806), .B(n2967), .Z(n2807) );
  XNOR U4481 ( .A(n3219), .B(n2807), .Z(out[233]) );
  XOR U4482 ( .A(in[1075]), .B(n4372), .Z(n3243) );
  NANDN U4483 ( .A(n2808), .B(n2969), .Z(n2809) );
  XNOR U4484 ( .A(n3243), .B(n2809), .Z(out[234]) );
  XOR U4485 ( .A(in[1076]), .B(n4375), .Z(n3255) );
  NANDN U4486 ( .A(n2810), .B(n2971), .Z(n2811) );
  XNOR U4487 ( .A(n3255), .B(n2811), .Z(out[235]) );
  XOR U4488 ( .A(in[1077]), .B(n4378), .Z(n3265) );
  NANDN U4489 ( .A(n2812), .B(n2977), .Z(n2813) );
  XNOR U4490 ( .A(n3265), .B(n2813), .Z(out[236]) );
  XOR U4491 ( .A(in[1078]), .B(n4381), .Z(n3299) );
  NAND U4492 ( .A(n2814), .B(n2979), .Z(n2815) );
  XNOR U4493 ( .A(n3299), .B(n2815), .Z(out[237]) );
  XOR U4494 ( .A(in[1079]), .B(n4384), .Z(n3329) );
  NAND U4495 ( .A(n2816), .B(n2981), .Z(n2817) );
  XNOR U4496 ( .A(n3329), .B(n2817), .Z(out[238]) );
  XNOR U4497 ( .A(in[1080]), .B(n4386), .Z(n3357) );
  NAND U4498 ( .A(n2818), .B(n2983), .Z(n2819) );
  XOR U4499 ( .A(n3357), .B(n2819), .Z(out[239]) );
  XOR U4500 ( .A(in[1433]), .B(n2820), .Z(n4671) );
  OR U4501 ( .A(n4671), .B(n2821), .Z(n2822) );
  XOR U4502 ( .A(n4670), .B(n2822), .Z(out[23]) );
  XOR U4503 ( .A(in[1081]), .B(n4389), .Z(n3385) );
  NAND U4504 ( .A(n2823), .B(n2985), .Z(n2824) );
  XNOR U4505 ( .A(n3385), .B(n2824), .Z(out[240]) );
  XOR U4506 ( .A(in[1082]), .B(n4392), .Z(n3420) );
  NANDN U4507 ( .A(n2987), .B(n2825), .Z(n2826) );
  XOR U4508 ( .A(n3420), .B(n2826), .Z(out[241]) );
  XOR U4509 ( .A(in[1083]), .B(n4395), .Z(n3455) );
  NAND U4510 ( .A(n2827), .B(n2988), .Z(n2828) );
  XOR U4511 ( .A(n3455), .B(n2828), .Z(out[242]) );
  XNOR U4512 ( .A(in[1084]), .B(n4398), .Z(n3477) );
  NAND U4513 ( .A(n2829), .B(n2990), .Z(n2830) );
  XOR U4514 ( .A(n3477), .B(n2830), .Z(out[243]) );
  XNOR U4515 ( .A(in[1085]), .B(n4405), .Z(n3499) );
  NAND U4516 ( .A(n2831), .B(n2992), .Z(n2832) );
  XOR U4517 ( .A(n3499), .B(n2832), .Z(out[244]) );
  XNOR U4518 ( .A(in[1086]), .B(n4408), .Z(n3514) );
  NAND U4519 ( .A(n2833), .B(n2994), .Z(n2834) );
  XOR U4520 ( .A(n3514), .B(n2834), .Z(out[245]) );
  XOR U4521 ( .A(in[1087]), .B(n4411), .Z(n2998) );
  NAND U4522 ( .A(n2835), .B(n2999), .Z(n2836) );
  XNOR U4523 ( .A(n2998), .B(n2836), .Z(out[246]) );
  XNOR U4524 ( .A(in[1024]), .B(n4414), .Z(n3574) );
  NAND U4525 ( .A(n2837), .B(n3001), .Z(n2838) );
  XOR U4526 ( .A(n3574), .B(n2838), .Z(out[247]) );
  XNOR U4527 ( .A(in[1025]), .B(n4417), .Z(n3598) );
  NAND U4528 ( .A(n2839), .B(n3003), .Z(n2840) );
  XOR U4529 ( .A(n3598), .B(n2840), .Z(out[248]) );
  XNOR U4530 ( .A(in[1026]), .B(n4420), .Z(n3628) );
  NAND U4531 ( .A(n2841), .B(n3005), .Z(n2842) );
  XOR U4532 ( .A(n3628), .B(n2842), .Z(out[249]) );
  XOR U4533 ( .A(in[1434]), .B(n2843), .Z(n4687) );
  OR U4534 ( .A(n4687), .B(n2844), .Z(n2845) );
  XNOR U4535 ( .A(n4686), .B(n2845), .Z(out[24]) );
  XNOR U4536 ( .A(in[1027]), .B(n4423), .Z(n3672) );
  NAND U4537 ( .A(n2846), .B(n3007), .Z(n2847) );
  XOR U4538 ( .A(n3672), .B(n2847), .Z(out[250]) );
  XOR U4539 ( .A(in[1028]), .B(n4426), .Z(n3010) );
  IV U4540 ( .A(n3010), .Z(n3716) );
  NANDN U4541 ( .A(n3009), .B(n2848), .Z(n2849) );
  XOR U4542 ( .A(n3716), .B(n2849), .Z(out[251]) );
  XOR U4543 ( .A(in[1029]), .B(n4429), .Z(n3013) );
  IV U4544 ( .A(n3013), .Z(n3762) );
  NANDN U4545 ( .A(n3012), .B(n2850), .Z(n2851) );
  XOR U4546 ( .A(n3762), .B(n2851), .Z(out[252]) );
  XOR U4547 ( .A(in[1030]), .B(n4432), .Z(n3806) );
  NANDN U4548 ( .A(n3015), .B(n2852), .Z(n2853) );
  XOR U4549 ( .A(n3806), .B(n2853), .Z(out[253]) );
  XOR U4550 ( .A(in[1031]), .B(n4443), .Z(n3017) );
  IV U4551 ( .A(n3017), .Z(n3850) );
  NANDN U4552 ( .A(n3016), .B(n2854), .Z(n2855) );
  XOR U4553 ( .A(n3850), .B(n2855), .Z(out[254]) );
  XOR U4554 ( .A(in[1032]), .B(n4446), .Z(n3020) );
  IV U4555 ( .A(n3020), .Z(n3894) );
  NANDN U4556 ( .A(n3019), .B(n2856), .Z(n2857) );
  XOR U4557 ( .A(n3894), .B(n2857), .Z(out[255]) );
  ANDN U4558 ( .B(n2861), .A(n2860), .Z(n2862) );
  XOR U4559 ( .A(n3981), .B(n2862), .Z(out[257]) );
  XNOR U4560 ( .A(n3943), .B(in[1412]), .Z(n4025) );
  NANDN U4561 ( .A(n2863), .B(n2975), .Z(n2864) );
  XNOR U4562 ( .A(n4025), .B(n2864), .Z(out[258]) );
  XNOR U4563 ( .A(n3947), .B(in[1413]), .Z(n4069) );
  NANDN U4564 ( .A(n2865), .B(n3168), .Z(n2866) );
  XNOR U4565 ( .A(n4069), .B(n2866), .Z(out[259]) );
  XOR U4566 ( .A(in[1435]), .B(n2867), .Z(n4722) );
  OR U4567 ( .A(n4722), .B(n2868), .Z(n2869) );
  XNOR U4568 ( .A(n4721), .B(n2869), .Z(out[25]) );
  XNOR U4569 ( .A(n3951), .B(in[1414]), .Z(n4113) );
  NANDN U4570 ( .A(n2870), .B(n3424), .Z(n2871) );
  XNOR U4571 ( .A(n4113), .B(n2871), .Z(out[260]) );
  XNOR U4572 ( .A(n3955), .B(in[1415]), .Z(n4157) );
  NANDN U4573 ( .A(n2872), .B(n3720), .Z(n2873) );
  XNOR U4574 ( .A(n4157), .B(n2873), .Z(out[261]) );
  XNOR U4575 ( .A(n3959), .B(in[1416]), .Z(n4195) );
  NANDN U4576 ( .A(n2874), .B(n4160), .Z(n2875) );
  XNOR U4577 ( .A(n4195), .B(n2875), .Z(out[262]) );
  XNOR U4578 ( .A(in[1417]), .B(n3963), .Z(n4440) );
  NANDN U4579 ( .A(n2876), .B(n4439), .Z(n2877) );
  XNOR U4580 ( .A(n4440), .B(n2877), .Z(out[263]) );
  XNOR U4581 ( .A(n3967), .B(in[1418]), .Z(n4726) );
  NANDN U4582 ( .A(n2878), .B(n4725), .Z(n2879) );
  XNOR U4583 ( .A(n4726), .B(n2879), .Z(out[264]) );
  XNOR U4584 ( .A(n3971), .B(in[1419]), .Z(n5154) );
  NANDN U4585 ( .A(n2880), .B(n5153), .Z(n2881) );
  XNOR U4586 ( .A(n5154), .B(n2881), .Z(out[265]) );
  NOR U4587 ( .A(n2883), .B(n2882), .Z(n2884) );
  XOR U4588 ( .A(n4281), .B(n2884), .Z(out[266]) );
  XOR U4589 ( .A(in[1436]), .B(n2891), .Z(n4770) );
  OR U4590 ( .A(n4770), .B(n2892), .Z(n2893) );
  XOR U4591 ( .A(n4769), .B(n2893), .Z(out[26]) );
  NOR U4592 ( .A(n2895), .B(n2894), .Z(n2896) );
  XOR U4593 ( .A(n4402), .B(n2896), .Z(out[270]) );
  NOR U4594 ( .A(n2898), .B(n2897), .Z(n2899) );
  XOR U4595 ( .A(n4436), .B(n2899), .Z(out[271]) );
  NOR U4596 ( .A(n2901), .B(n2900), .Z(n2902) );
  XOR U4597 ( .A(n4474), .B(n2902), .Z(out[272]) );
  NOR U4598 ( .A(n2904), .B(n2903), .Z(n2905) );
  XOR U4599 ( .A(n4508), .B(n2905), .Z(out[273]) );
  NOR U4600 ( .A(n2907), .B(n2906), .Z(n2908) );
  XOR U4601 ( .A(n4547), .B(n2908), .Z(out[274]) );
  NOR U4602 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U4603 ( .A(n4576), .B(n2911), .Z(out[275]) );
  NOR U4604 ( .A(n2913), .B(n2912), .Z(n2914) );
  XOR U4605 ( .A(n4601), .B(n2914), .Z(out[276]) );
  ANDN U4606 ( .B(n2916), .A(n2915), .Z(n2917) );
  XOR U4607 ( .A(n4626), .B(n2917), .Z(out[277]) );
  ANDN U4608 ( .B(n2919), .A(n2918), .Z(n2920) );
  XOR U4609 ( .A(n4656), .B(n2920), .Z(out[278]) );
  ANDN U4610 ( .B(n2922), .A(n2921), .Z(n2923) );
  XOR U4611 ( .A(n4671), .B(n2923), .Z(out[279]) );
  XOR U4612 ( .A(in[1437]), .B(n2924), .Z(n4813) );
  OR U4613 ( .A(n4813), .B(n2925), .Z(n2926) );
  XOR U4614 ( .A(n4812), .B(n2926), .Z(out[27]) );
  ANDN U4615 ( .B(n2928), .A(n2927), .Z(n2929) );
  XOR U4616 ( .A(n4687), .B(n2929), .Z(out[280]) );
  ANDN U4617 ( .B(n2931), .A(n2930), .Z(n2932) );
  XOR U4618 ( .A(n4722), .B(n2932), .Z(out[281]) );
  ANDN U4619 ( .B(n2934), .A(n2933), .Z(n2935) );
  XOR U4620 ( .A(n4770), .B(n2935), .Z(out[282]) );
  ANDN U4621 ( .B(n2937), .A(n2936), .Z(n2938) );
  XOR U4622 ( .A(n4813), .B(n2938), .Z(out[283]) );
  XOR U4623 ( .A(in[1438]), .B(n4054), .Z(n4855) );
  NAND U4624 ( .A(n2939), .B(n2951), .Z(n2940) );
  XNOR U4625 ( .A(n4855), .B(n2940), .Z(out[284]) );
  XOR U4626 ( .A(in[1439]), .B(n4058), .Z(n4899) );
  NAND U4627 ( .A(n2941), .B(n2973), .Z(n2942) );
  XNOR U4628 ( .A(n4899), .B(n2942), .Z(out[285]) );
  XOR U4629 ( .A(in[1440]), .B(n4062), .Z(n4943) );
  NAND U4630 ( .A(n2943), .B(n2996), .Z(n2944) );
  XNOR U4631 ( .A(n4943), .B(n2944), .Z(out[286]) );
  XOR U4632 ( .A(in[1441]), .B(n4066), .Z(n4987) );
  NAND U4633 ( .A(n2945), .B(n3022), .Z(n2946) );
  XNOR U4634 ( .A(n4987), .B(n2946), .Z(out[287]) );
  XOR U4635 ( .A(in[1442]), .B(n4074), .Z(n5031) );
  NAND U4636 ( .A(n2947), .B(n3042), .Z(n2948) );
  XNOR U4637 ( .A(n5031), .B(n2948), .Z(out[288]) );
  XOR U4638 ( .A(in[1443]), .B(n4078), .Z(n5072) );
  NAND U4639 ( .A(n2949), .B(n3054), .Z(n2950) );
  XNOR U4640 ( .A(n5072), .B(n2950), .Z(out[289]) );
  OR U4641 ( .A(n4855), .B(n2951), .Z(n2952) );
  XOR U4642 ( .A(n4856), .B(n2952), .Z(out[28]) );
  XOR U4643 ( .A(in[1444]), .B(n4082), .Z(n5108) );
  NAND U4644 ( .A(n2953), .B(n3075), .Z(n2954) );
  XNOR U4645 ( .A(n5108), .B(n2954), .Z(out[290]) );
  XNOR U4646 ( .A(in[1445]), .B(n4086), .Z(n5150) );
  NANDN U4647 ( .A(n2955), .B(n3096), .Z(n2956) );
  XNOR U4648 ( .A(n5150), .B(n2956), .Z(out[291]) );
  OR U4649 ( .A(n3115), .B(n2957), .Z(n2958) );
  XNOR U4650 ( .A(n3114), .B(n2958), .Z(out[292]) );
  OR U4651 ( .A(n3135), .B(n2959), .Z(n2960) );
  XNOR U4652 ( .A(n3134), .B(n2960), .Z(out[293]) );
  NANDN U4653 ( .A(n2961), .B(n3153), .Z(n2962) );
  XNOR U4654 ( .A(n3154), .B(n2962), .Z(out[294]) );
  OR U4655 ( .A(n3165), .B(n2963), .Z(n2964) );
  XNOR U4656 ( .A(n3164), .B(n2964), .Z(out[295]) );
  OR U4657 ( .A(n3190), .B(n2965), .Z(n2966) );
  XNOR U4658 ( .A(n3189), .B(n2966), .Z(out[296]) );
  OR U4659 ( .A(n3219), .B(n2967), .Z(n2968) );
  XOR U4660 ( .A(n3220), .B(n2968), .Z(out[297]) );
  OR U4661 ( .A(n3243), .B(n2969), .Z(n2970) );
  XOR U4662 ( .A(n3244), .B(n2970), .Z(out[298]) );
  OR U4663 ( .A(n3255), .B(n2971), .Z(n2972) );
  XOR U4664 ( .A(n3256), .B(n2972), .Z(out[299]) );
  OR U4665 ( .A(n4899), .B(n2973), .Z(n2974) );
  XOR U4666 ( .A(n4900), .B(n2974), .Z(out[29]) );
  OR U4667 ( .A(n4025), .B(n2975), .Z(n2976) );
  XNOR U4668 ( .A(n4024), .B(n2976), .Z(out[2]) );
  OR U4669 ( .A(n3265), .B(n2977), .Z(n2978) );
  XOR U4670 ( .A(n3266), .B(n2978), .Z(out[300]) );
  OR U4671 ( .A(n3299), .B(n2979), .Z(n2980) );
  XOR U4672 ( .A(n3300), .B(n2980), .Z(out[301]) );
  OR U4673 ( .A(n3329), .B(n2981), .Z(n2982) );
  XOR U4674 ( .A(n3330), .B(n2982), .Z(out[302]) );
  NANDN U4675 ( .A(n2983), .B(n3357), .Z(n2984) );
  XOR U4676 ( .A(n3358), .B(n2984), .Z(out[303]) );
  OR U4677 ( .A(n3385), .B(n2985), .Z(n2986) );
  XOR U4678 ( .A(n3386), .B(n2986), .Z(out[304]) );
  NANDN U4679 ( .A(n2988), .B(n3455), .Z(n2989) );
  XOR U4680 ( .A(n3456), .B(n2989), .Z(out[306]) );
  NANDN U4681 ( .A(n2990), .B(n3477), .Z(n2991) );
  XOR U4682 ( .A(n3478), .B(n2991), .Z(out[307]) );
  NANDN U4683 ( .A(n2992), .B(n3499), .Z(n2993) );
  XOR U4684 ( .A(n3500), .B(n2993), .Z(out[308]) );
  NANDN U4685 ( .A(n2994), .B(n3514), .Z(n2995) );
  XOR U4686 ( .A(n3515), .B(n2995), .Z(out[309]) );
  OR U4687 ( .A(n4943), .B(n2996), .Z(n2997) );
  XOR U4688 ( .A(n4944), .B(n2997), .Z(out[30]) );
  IV U4689 ( .A(n2998), .Z(n3544) );
  NANDN U4690 ( .A(n2999), .B(n3544), .Z(n3000) );
  XOR U4691 ( .A(n3545), .B(n3000), .Z(out[310]) );
  NANDN U4692 ( .A(n3001), .B(n3574), .Z(n3002) );
  XOR U4693 ( .A(n3575), .B(n3002), .Z(out[311]) );
  NANDN U4694 ( .A(n3003), .B(n3598), .Z(n3004) );
  XOR U4695 ( .A(n3599), .B(n3004), .Z(out[312]) );
  NANDN U4696 ( .A(n3005), .B(n3628), .Z(n3006) );
  XOR U4697 ( .A(n3629), .B(n3006), .Z(out[313]) );
  NANDN U4698 ( .A(n3007), .B(n3672), .Z(n3008) );
  XOR U4699 ( .A(n3673), .B(n3008), .Z(out[314]) );
  NANDN U4700 ( .A(n3010), .B(n3009), .Z(n3011) );
  XOR U4701 ( .A(n3717), .B(n3011), .Z(out[315]) );
  NANDN U4702 ( .A(n3013), .B(n3012), .Z(n3014) );
  XOR U4703 ( .A(n3763), .B(n3014), .Z(out[316]) );
  NANDN U4704 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U4705 ( .A(n3851), .B(n3018), .Z(out[318]) );
  NANDN U4706 ( .A(n3020), .B(n3019), .Z(n3021) );
  XOR U4707 ( .A(n3895), .B(n3021), .Z(out[319]) );
  OR U4708 ( .A(n4987), .B(n3022), .Z(n3023) );
  XOR U4709 ( .A(n4988), .B(n3023), .Z(out[31]) );
  XOR U4710 ( .A(in[72]), .B(n4446), .Z(n3260) );
  XOR U4711 ( .A(in[1317]), .B(n4278), .Z(n3615) );
  XNOR U4712 ( .A(in[1244]), .B(n3024), .Z(n3612) );
  NANDN U4713 ( .A(n3615), .B(n3612), .Z(n3025) );
  XNOR U4714 ( .A(n3260), .B(n3025), .Z(out[320]) );
  XOR U4715 ( .A(in[73]), .B(n4449), .Z(n3147) );
  IV U4716 ( .A(n3147), .Z(n3263) );
  XOR U4717 ( .A(in[1318]), .B(n4284), .Z(n3619) );
  XNOR U4718 ( .A(in[1245]), .B(n3026), .Z(n3616) );
  NANDN U4719 ( .A(n3619), .B(n3616), .Z(n3027) );
  XOR U4720 ( .A(n3263), .B(n3027), .Z(out[321]) );
  XOR U4721 ( .A(in[74]), .B(n4452), .Z(n3149) );
  IV U4722 ( .A(n3149), .Z(n3270) );
  XOR U4723 ( .A(in[1319]), .B(n4286), .Z(n3623) );
  XNOR U4724 ( .A(in[1246]), .B(n3028), .Z(n3620) );
  NANDN U4725 ( .A(n3623), .B(n3620), .Z(n3029) );
  XOR U4726 ( .A(n3270), .B(n3029), .Z(out[322]) );
  XOR U4727 ( .A(in[75]), .B(n4455), .Z(n3151) );
  IV U4728 ( .A(n3151), .Z(n3273) );
  XOR U4729 ( .A(in[1320]), .B(n4288), .Z(n3627) );
  XNOR U4730 ( .A(in[1247]), .B(n3030), .Z(n3624) );
  NANDN U4731 ( .A(n3627), .B(n3624), .Z(n3031) );
  XOR U4732 ( .A(n3273), .B(n3031), .Z(out[323]) );
  XNOR U4733 ( .A(n4458), .B(in[76]), .Z(n3276) );
  XOR U4734 ( .A(in[1321]), .B(n4290), .Z(n3635) );
  XNOR U4735 ( .A(in[1248]), .B(n3032), .Z(n3632) );
  NANDN U4736 ( .A(n3635), .B(n3632), .Z(n3033) );
  XNOR U4737 ( .A(n3276), .B(n3033), .Z(out[324]) );
  XNOR U4738 ( .A(n4461), .B(in[77]), .Z(n3279) );
  XOR U4739 ( .A(in[1322]), .B(n4292), .Z(n3639) );
  XNOR U4740 ( .A(in[1249]), .B(n3034), .Z(n3636) );
  NANDN U4741 ( .A(n3639), .B(n3636), .Z(n3035) );
  XNOR U4742 ( .A(n3279), .B(n3035), .Z(out[325]) );
  XNOR U4743 ( .A(n4464), .B(in[78]), .Z(n3282) );
  XOR U4744 ( .A(in[1323]), .B(n4294), .Z(n3643) );
  XOR U4745 ( .A(in[1250]), .B(n4124), .Z(n3640) );
  NANDN U4746 ( .A(n3643), .B(n3640), .Z(n3036) );
  XNOR U4747 ( .A(n3282), .B(n3036), .Z(out[326]) );
  XNOR U4748 ( .A(n4467), .B(in[79]), .Z(n3285) );
  XOR U4749 ( .A(in[1324]), .B(n4296), .Z(n3647) );
  XNOR U4750 ( .A(in[1251]), .B(n3037), .Z(n3644) );
  NANDN U4751 ( .A(n3647), .B(n3644), .Z(n3038) );
  XNOR U4752 ( .A(n3285), .B(n3038), .Z(out[327]) );
  XNOR U4753 ( .A(n4470), .B(in[80]), .Z(n3288) );
  XOR U4754 ( .A(in[1325]), .B(n4298), .Z(n3651) );
  XNOR U4755 ( .A(in[1252]), .B(n3039), .Z(n3648) );
  NANDN U4756 ( .A(n3651), .B(n3648), .Z(n3040) );
  XNOR U4757 ( .A(n3288), .B(n3040), .Z(out[328]) );
  XNOR U4758 ( .A(n4477), .B(in[81]), .Z(n3291) );
  XNOR U4759 ( .A(in[1253]), .B(n4136), .Z(n3653) );
  XNOR U4760 ( .A(in[1326]), .B(n4300), .Z(n3655) );
  NANDN U4761 ( .A(n3653), .B(n3655), .Z(n3041) );
  XNOR U4762 ( .A(n3291), .B(n3041), .Z(out[329]) );
  OR U4763 ( .A(n5031), .B(n3042), .Z(n3043) );
  XOR U4764 ( .A(n5032), .B(n3043), .Z(out[32]) );
  XNOR U4765 ( .A(n4480), .B(in[82]), .Z(n3294) );
  XNOR U4766 ( .A(in[1254]), .B(n4140), .Z(n3657) );
  XNOR U4767 ( .A(in[1327]), .B(n4302), .Z(n3659) );
  NANDN U4768 ( .A(n3657), .B(n3659), .Z(n3044) );
  XNOR U4769 ( .A(n3294), .B(n3044), .Z(out[330]) );
  XNOR U4770 ( .A(n4483), .B(in[83]), .Z(n3297) );
  XNOR U4771 ( .A(in[1255]), .B(n4144), .Z(n3661) );
  XNOR U4772 ( .A(in[1328]), .B(n4309), .Z(n3663) );
  NANDN U4773 ( .A(n3661), .B(n3663), .Z(n3045) );
  XNOR U4774 ( .A(n3297), .B(n3045), .Z(out[331]) );
  XNOR U4775 ( .A(in[84]), .B(n4486), .Z(n3304) );
  XNOR U4776 ( .A(in[1256]), .B(n4148), .Z(n3665) );
  XNOR U4777 ( .A(in[1329]), .B(n4312), .Z(n3667) );
  NANDN U4778 ( .A(n3665), .B(n3667), .Z(n3046) );
  XNOR U4779 ( .A(n3304), .B(n3046), .Z(out[332]) );
  XNOR U4780 ( .A(in[85]), .B(n4489), .Z(n3307) );
  XNOR U4781 ( .A(in[1257]), .B(n4152), .Z(n3669) );
  XNOR U4782 ( .A(in[1330]), .B(n4315), .Z(n3671) );
  NANDN U4783 ( .A(n3669), .B(n3671), .Z(n3047) );
  XNOR U4784 ( .A(n3307), .B(n3047), .Z(out[333]) );
  XNOR U4785 ( .A(in[86]), .B(n4492), .Z(n3310) );
  XNOR U4786 ( .A(in[1258]), .B(n4162), .Z(n3677) );
  XNOR U4787 ( .A(in[1331]), .B(n4318), .Z(n3679) );
  NANDN U4788 ( .A(n3677), .B(n3679), .Z(n3048) );
  XNOR U4789 ( .A(n3310), .B(n3048), .Z(out[334]) );
  XNOR U4790 ( .A(in[87]), .B(n4495), .Z(n3313) );
  XNOR U4791 ( .A(in[1259]), .B(n4166), .Z(n3681) );
  XNOR U4792 ( .A(in[1332]), .B(n4321), .Z(n3683) );
  NANDN U4793 ( .A(n3681), .B(n3683), .Z(n3049) );
  XNOR U4794 ( .A(n3313), .B(n3049), .Z(out[335]) );
  XNOR U4795 ( .A(in[88]), .B(n4498), .Z(n3316) );
  XNOR U4796 ( .A(in[1260]), .B(n4170), .Z(n3685) );
  XNOR U4797 ( .A(in[1333]), .B(n4324), .Z(n3687) );
  NANDN U4798 ( .A(n3685), .B(n3687), .Z(n3050) );
  XNOR U4799 ( .A(n3316), .B(n3050), .Z(out[336]) );
  XNOR U4800 ( .A(in[89]), .B(n4501), .Z(n3319) );
  XNOR U4801 ( .A(in[1261]), .B(n4174), .Z(n3689) );
  XNOR U4802 ( .A(in[1334]), .B(n4327), .Z(n3691) );
  NANDN U4803 ( .A(n3689), .B(n3691), .Z(n3051) );
  XNOR U4804 ( .A(n3319), .B(n3051), .Z(out[337]) );
  XNOR U4805 ( .A(in[90]), .B(n4504), .Z(n3321) );
  XNOR U4806 ( .A(in[1262]), .B(n3898), .Z(n3693) );
  XNOR U4807 ( .A(in[1335]), .B(n4330), .Z(n3695) );
  NANDN U4808 ( .A(n3693), .B(n3695), .Z(n3052) );
  XNOR U4809 ( .A(n3321), .B(n3052), .Z(out[338]) );
  XOR U4810 ( .A(in[91]), .B(n4511), .Z(n3323) );
  XNOR U4811 ( .A(in[1263]), .B(n3902), .Z(n3697) );
  XNOR U4812 ( .A(in[1336]), .B(n4178), .Z(n3699) );
  NANDN U4813 ( .A(n3697), .B(n3699), .Z(n3053) );
  XNOR U4814 ( .A(n3323), .B(n3053), .Z(out[339]) );
  OR U4815 ( .A(n5072), .B(n3054), .Z(n3055) );
  XOR U4816 ( .A(n5073), .B(n3055), .Z(out[33]) );
  XOR U4817 ( .A(in[92]), .B(n4514), .Z(n3325) );
  XNOR U4818 ( .A(in[1264]), .B(n3906), .Z(n3701) );
  XNOR U4819 ( .A(in[1337]), .B(n4181), .Z(n3703) );
  NANDN U4820 ( .A(n3701), .B(n3703), .Z(n3056) );
  XNOR U4821 ( .A(n3325), .B(n3056), .Z(out[340]) );
  XOR U4822 ( .A(in[93]), .B(n4517), .Z(n3327) );
  XNOR U4823 ( .A(in[1265]), .B(n3910), .Z(n3705) );
  XNOR U4824 ( .A(in[1338]), .B(n4184), .Z(n3707) );
  NANDN U4825 ( .A(n3705), .B(n3707), .Z(n3057) );
  XNOR U4826 ( .A(n3327), .B(n3057), .Z(out[341]) );
  XNOR U4827 ( .A(in[94]), .B(n4520), .Z(n3333) );
  XNOR U4828 ( .A(in[1266]), .B(n3914), .Z(n3709) );
  XNOR U4829 ( .A(in[1339]), .B(n4187), .Z(n3711) );
  NANDN U4830 ( .A(n3709), .B(n3711), .Z(n3058) );
  XNOR U4831 ( .A(n3333), .B(n3058), .Z(out[342]) );
  XNOR U4832 ( .A(in[95]), .B(n4524), .Z(n3335) );
  XOR U4833 ( .A(in[1267]), .B(n3918), .Z(n3713) );
  XNOR U4834 ( .A(in[1340]), .B(n3059), .Z(n3715) );
  NANDN U4835 ( .A(n3713), .B(n3715), .Z(n3060) );
  XNOR U4836 ( .A(n3335), .B(n3060), .Z(out[343]) );
  XNOR U4837 ( .A(in[96]), .B(n4528), .Z(n3337) );
  XOR U4838 ( .A(in[1268]), .B(n3922), .Z(n3723) );
  XNOR U4839 ( .A(in[1341]), .B(n3061), .Z(n3725) );
  NANDN U4840 ( .A(n3723), .B(n3725), .Z(n3062) );
  XNOR U4841 ( .A(n3337), .B(n3062), .Z(out[344]) );
  XNOR U4842 ( .A(in[97]), .B(n4532), .Z(n3339) );
  XOR U4843 ( .A(in[1269]), .B(n3926), .Z(n3727) );
  XNOR U4844 ( .A(in[1342]), .B(n3063), .Z(n3729) );
  NANDN U4845 ( .A(n3727), .B(n3729), .Z(n3064) );
  XNOR U4846 ( .A(n3339), .B(n3064), .Z(out[345]) );
  XNOR U4847 ( .A(in[98]), .B(n4536), .Z(n3341) );
  IV U4848 ( .A(n3065), .Z(n3930) );
  XOR U4849 ( .A(in[1270]), .B(n3930), .Z(n3731) );
  XNOR U4850 ( .A(in[1343]), .B(n4199), .Z(n3733) );
  NANDN U4851 ( .A(n3731), .B(n3733), .Z(n3066) );
  XNOR U4852 ( .A(n3341), .B(n3066), .Z(out[346]) );
  XNOR U4853 ( .A(in[99]), .B(n4540), .Z(n3343) );
  IV U4854 ( .A(n3067), .Z(n3934) );
  XOR U4855 ( .A(in[1271]), .B(n3934), .Z(n3735) );
  XNOR U4856 ( .A(in[1280]), .B(n3068), .Z(n3737) );
  NANDN U4857 ( .A(n3735), .B(n3737), .Z(n3069) );
  XNOR U4858 ( .A(n3343), .B(n3069), .Z(out[347]) );
  XOR U4859 ( .A(in[100]), .B(n4544), .Z(n3197) );
  IV U4860 ( .A(n3197), .Z(n3346) );
  IV U4861 ( .A(n3070), .Z(n3941) );
  XOR U4862 ( .A(in[1272]), .B(n3941), .Z(n3739) );
  XNOR U4863 ( .A(in[1281]), .B(n3071), .Z(n3741) );
  NANDN U4864 ( .A(n3739), .B(n3741), .Z(n3072) );
  XOR U4865 ( .A(n3346), .B(n3072), .Z(out[348]) );
  XOR U4866 ( .A(in[101]), .B(n4550), .Z(n3200) );
  IV U4867 ( .A(n3200), .Z(n3349) );
  XOR U4868 ( .A(in[1273]), .B(n3945), .Z(n3743) );
  XNOR U4869 ( .A(in[1282]), .B(n3073), .Z(n3745) );
  NANDN U4870 ( .A(n3743), .B(n3745), .Z(n3074) );
  XOR U4871 ( .A(n3349), .B(n3074), .Z(out[349]) );
  OR U4872 ( .A(n5108), .B(n3075), .Z(n3076) );
  XNOR U4873 ( .A(n5107), .B(n3076), .Z(out[34]) );
  XOR U4874 ( .A(in[102]), .B(n4552), .Z(n3203) );
  IV U4875 ( .A(n3203), .Z(n3352) );
  XOR U4876 ( .A(in[1274]), .B(n3949), .Z(n3747) );
  XNOR U4877 ( .A(in[1283]), .B(n3077), .Z(n3749) );
  NANDN U4878 ( .A(n3747), .B(n3749), .Z(n3078) );
  XOR U4879 ( .A(n3352), .B(n3078), .Z(out[350]) );
  XOR U4880 ( .A(in[103]), .B(n4333), .Z(n3206) );
  IV U4881 ( .A(n3206), .Z(n3355) );
  XNOR U4882 ( .A(in[1275]), .B(n3953), .Z(n3751) );
  XNOR U4883 ( .A(in[1284]), .B(n3079), .Z(n3753) );
  NANDN U4884 ( .A(n3751), .B(n3753), .Z(n3080) );
  XOR U4885 ( .A(n3355), .B(n3080), .Z(out[351]) );
  XOR U4886 ( .A(in[104]), .B(n4335), .Z(n3209) );
  IV U4887 ( .A(n3209), .Z(n3362) );
  XNOR U4888 ( .A(in[1276]), .B(n3957), .Z(n3755) );
  XNOR U4889 ( .A(in[1285]), .B(n3081), .Z(n3757) );
  NANDN U4890 ( .A(n3755), .B(n3757), .Z(n3082) );
  XOR U4891 ( .A(n3362), .B(n3082), .Z(out[352]) );
  XOR U4892 ( .A(in[105]), .B(n4341), .Z(n3211) );
  IV U4893 ( .A(n3211), .Z(n3365) );
  XNOR U4894 ( .A(in[1277]), .B(n3961), .Z(n3759) );
  XNOR U4895 ( .A(in[1286]), .B(n3083), .Z(n3761) );
  NANDN U4896 ( .A(n3759), .B(n3761), .Z(n3084) );
  XOR U4897 ( .A(n3365), .B(n3084), .Z(out[353]) );
  XOR U4898 ( .A(in[106]), .B(n4343), .Z(n3214) );
  IV U4899 ( .A(n3214), .Z(n3368) );
  XNOR U4900 ( .A(in[1278]), .B(n3965), .Z(n3767) );
  XNOR U4901 ( .A(in[1287]), .B(n3085), .Z(n3769) );
  NANDN U4902 ( .A(n3767), .B(n3769), .Z(n3086) );
  XOR U4903 ( .A(n3368), .B(n3086), .Z(out[354]) );
  XOR U4904 ( .A(in[107]), .B(n4345), .Z(n3217) );
  IV U4905 ( .A(n3217), .Z(n3371) );
  XNOR U4906 ( .A(in[1279]), .B(n3969), .Z(n3771) );
  XNOR U4907 ( .A(in[1288]), .B(n4216), .Z(n3773) );
  NANDN U4908 ( .A(n3771), .B(n3773), .Z(n3087) );
  XOR U4909 ( .A(n3371), .B(n3087), .Z(out[355]) );
  XOR U4910 ( .A(in[108]), .B(n4348), .Z(n3223) );
  IV U4911 ( .A(n3223), .Z(n3373) );
  XNOR U4912 ( .A(in[1216]), .B(n3973), .Z(n3775) );
  XNOR U4913 ( .A(in[1289]), .B(n3088), .Z(n3777) );
  NANDN U4914 ( .A(n3775), .B(n3777), .Z(n3089) );
  XOR U4915 ( .A(n3373), .B(n3089), .Z(out[356]) );
  XOR U4916 ( .A(in[109]), .B(n4351), .Z(n3225) );
  IV U4917 ( .A(n3225), .Z(n3375) );
  XNOR U4918 ( .A(in[1217]), .B(n3977), .Z(n3779) );
  XNOR U4919 ( .A(in[1290]), .B(n3090), .Z(n3781) );
  NANDN U4920 ( .A(n3779), .B(n3781), .Z(n3091) );
  XOR U4921 ( .A(n3375), .B(n3091), .Z(out[357]) );
  XOR U4922 ( .A(in[110]), .B(n4354), .Z(n3227) );
  IV U4923 ( .A(n3227), .Z(n3377) );
  XNOR U4924 ( .A(in[1218]), .B(n3984), .Z(n3783) );
  XNOR U4925 ( .A(in[1291]), .B(n3092), .Z(n3785) );
  NANDN U4926 ( .A(n3783), .B(n3785), .Z(n3093) );
  XOR U4927 ( .A(n3377), .B(n3093), .Z(out[358]) );
  XOR U4928 ( .A(in[111]), .B(n4356), .Z(n3229) );
  IV U4929 ( .A(n3229), .Z(n3379) );
  XNOR U4930 ( .A(in[1219]), .B(n3988), .Z(n3787) );
  XNOR U4931 ( .A(in[1292]), .B(n3094), .Z(n3789) );
  NANDN U4932 ( .A(n3787), .B(n3789), .Z(n3095) );
  XOR U4933 ( .A(n3379), .B(n3095), .Z(out[359]) );
  OR U4934 ( .A(n5150), .B(n3096), .Z(n3097) );
  XNOR U4935 ( .A(n5149), .B(n3097), .Z(out[35]) );
  XOR U4936 ( .A(in[112]), .B(n4359), .Z(n3231) );
  IV U4937 ( .A(n3231), .Z(n3381) );
  XOR U4938 ( .A(in[1293]), .B(n3098), .Z(n3793) );
  XOR U4939 ( .A(in[1220]), .B(n3992), .Z(n3790) );
  NANDN U4940 ( .A(n3793), .B(n3790), .Z(n3099) );
  XOR U4941 ( .A(n3381), .B(n3099), .Z(out[360]) );
  XOR U4942 ( .A(in[113]), .B(n4362), .Z(n3233) );
  IV U4943 ( .A(n3233), .Z(n3383) );
  XOR U4944 ( .A(in[1294]), .B(n3100), .Z(n3797) );
  XOR U4945 ( .A(in[1221]), .B(n3996), .Z(n3794) );
  NANDN U4946 ( .A(n3797), .B(n3794), .Z(n3101) );
  XOR U4947 ( .A(n3383), .B(n3101), .Z(out[361]) );
  XOR U4948 ( .A(in[114]), .B(n4365), .Z(n3235) );
  IV U4949 ( .A(n3235), .Z(n3389) );
  XOR U4950 ( .A(in[1295]), .B(n4237), .Z(n3801) );
  XOR U4951 ( .A(in[1222]), .B(n4000), .Z(n3798) );
  NANDN U4952 ( .A(n3801), .B(n3798), .Z(n3102) );
  XOR U4953 ( .A(n3389), .B(n3102), .Z(out[362]) );
  XOR U4954 ( .A(in[115]), .B(n4372), .Z(n3237) );
  IV U4955 ( .A(n3237), .Z(n3391) );
  XOR U4956 ( .A(in[1296]), .B(n3103), .Z(n3805) );
  XOR U4957 ( .A(in[1223]), .B(n4004), .Z(n3802) );
  NANDN U4958 ( .A(n3805), .B(n3802), .Z(n3104) );
  XOR U4959 ( .A(n3391), .B(n3104), .Z(out[363]) );
  XOR U4960 ( .A(in[116]), .B(n4375), .Z(n3239) );
  IV U4961 ( .A(n3239), .Z(n3394) );
  XOR U4962 ( .A(in[1297]), .B(n3105), .Z(n3813) );
  XOR U4963 ( .A(in[1224]), .B(n4008), .Z(n3810) );
  NANDN U4964 ( .A(n3813), .B(n3810), .Z(n3106) );
  XOR U4965 ( .A(n3394), .B(n3106), .Z(out[364]) );
  XOR U4966 ( .A(in[117]), .B(n4378), .Z(n3241) );
  IV U4967 ( .A(n3241), .Z(n3398) );
  XOR U4968 ( .A(in[1298]), .B(n3107), .Z(n3817) );
  XOR U4969 ( .A(in[1225]), .B(n4012), .Z(n3814) );
  NANDN U4970 ( .A(n3817), .B(n3814), .Z(n3108) );
  XOR U4971 ( .A(n3398), .B(n3108), .Z(out[365]) );
  XOR U4972 ( .A(in[118]), .B(n4381), .Z(n3247) );
  IV U4973 ( .A(n3247), .Z(n3402) );
  XOR U4974 ( .A(in[1299]), .B(n3109), .Z(n3821) );
  XOR U4975 ( .A(in[1226]), .B(n4016), .Z(n3818) );
  NANDN U4976 ( .A(n3821), .B(n3818), .Z(n3110) );
  XOR U4977 ( .A(n3402), .B(n3110), .Z(out[366]) );
  XOR U4978 ( .A(in[119]), .B(n4384), .Z(n3249) );
  IV U4979 ( .A(n3249), .Z(n3406) );
  XOR U4980 ( .A(in[1300]), .B(n4248), .Z(n3825) );
  XNOR U4981 ( .A(in[1227]), .B(n4020), .Z(n3822) );
  NANDN U4982 ( .A(n3825), .B(n3822), .Z(n3111) );
  XOR U4983 ( .A(n3406), .B(n3111), .Z(out[367]) );
  XOR U4984 ( .A(in[120]), .B(n4386), .Z(n3251) );
  IV U4985 ( .A(n3251), .Z(n3409) );
  XOR U4986 ( .A(in[1301]), .B(n4249), .Z(n3829) );
  XOR U4987 ( .A(in[1228]), .B(n4028), .Z(n3826) );
  NANDN U4988 ( .A(n3829), .B(n3826), .Z(n3112) );
  XOR U4989 ( .A(n3409), .B(n3112), .Z(out[368]) );
  XOR U4990 ( .A(in[121]), .B(n4389), .Z(n3253) );
  IV U4991 ( .A(n3253), .Z(n3412) );
  XOR U4992 ( .A(in[1302]), .B(n4250), .Z(n3833) );
  XNOR U4993 ( .A(in[1229]), .B(n4032), .Z(n3830) );
  NANDN U4994 ( .A(n3833), .B(n3830), .Z(n3113) );
  XOR U4995 ( .A(n3412), .B(n3113), .Z(out[369]) );
  ANDN U4996 ( .B(n3115), .A(n3114), .Z(n3116) );
  XOR U4997 ( .A(n3117), .B(n3116), .Z(out[36]) );
  XOR U4998 ( .A(in[122]), .B(n4392), .Z(n3415) );
  XOR U4999 ( .A(in[1303]), .B(n4251), .Z(n3837) );
  XNOR U5000 ( .A(in[1230]), .B(n3118), .Z(n3834) );
  NANDN U5001 ( .A(n3837), .B(n3834), .Z(n3119) );
  XOR U5002 ( .A(n3415), .B(n3119), .Z(out[370]) );
  XOR U5003 ( .A(in[123]), .B(n4395), .Z(n3418) );
  XOR U5004 ( .A(in[1304]), .B(n4252), .Z(n3841) );
  XNOR U5005 ( .A(in[1231]), .B(n4040), .Z(n3838) );
  NANDN U5006 ( .A(n3841), .B(n3838), .Z(n3120) );
  XOR U5007 ( .A(n3418), .B(n3120), .Z(out[371]) );
  XOR U5008 ( .A(in[124]), .B(n4398), .Z(n3426) );
  XOR U5009 ( .A(in[1305]), .B(n4253), .Z(n3845) );
  XNOR U5010 ( .A(in[1232]), .B(n4044), .Z(n3842) );
  NANDN U5011 ( .A(n3845), .B(n3842), .Z(n3121) );
  XNOR U5012 ( .A(n3426), .B(n3121), .Z(out[372]) );
  XOR U5013 ( .A(in[125]), .B(n4405), .Z(n3429) );
  XOR U5014 ( .A(in[1306]), .B(n4254), .Z(n3849) );
  XOR U5015 ( .A(in[1233]), .B(n4048), .Z(n3846) );
  NANDN U5016 ( .A(n3849), .B(n3846), .Z(n3122) );
  XNOR U5017 ( .A(n3429), .B(n3122), .Z(out[373]) );
  XOR U5018 ( .A(in[126]), .B(n4408), .Z(n3432) );
  XOR U5019 ( .A(in[1307]), .B(n4255), .Z(n3857) );
  XOR U5020 ( .A(in[1234]), .B(n4052), .Z(n3854) );
  NANDN U5021 ( .A(n3857), .B(n3854), .Z(n3123) );
  XNOR U5022 ( .A(n3432), .B(n3123), .Z(out[374]) );
  XOR U5023 ( .A(in[127]), .B(n4411), .Z(n3435) );
  XOR U5024 ( .A(in[1308]), .B(n4258), .Z(n3861) );
  XNOR U5025 ( .A(in[1235]), .B(n3124), .Z(n3858) );
  NANDN U5026 ( .A(n3861), .B(n3858), .Z(n3125) );
  XNOR U5027 ( .A(n3435), .B(n3125), .Z(out[375]) );
  XOR U5028 ( .A(in[64]), .B(n4414), .Z(n3438) );
  XOR U5029 ( .A(in[1309]), .B(n4259), .Z(n3865) );
  XNOR U5030 ( .A(in[1236]), .B(n3126), .Z(n3862) );
  NANDN U5031 ( .A(n3865), .B(n3862), .Z(n3127) );
  XNOR U5032 ( .A(n3438), .B(n3127), .Z(out[376]) );
  XOR U5033 ( .A(in[65]), .B(n4417), .Z(n3441) );
  XOR U5034 ( .A(in[1310]), .B(n4260), .Z(n3869) );
  XNOR U5035 ( .A(in[1237]), .B(n3128), .Z(n3866) );
  NANDN U5036 ( .A(n3869), .B(n3866), .Z(n3129) );
  XNOR U5037 ( .A(n3441), .B(n3129), .Z(out[377]) );
  XOR U5038 ( .A(in[66]), .B(n4420), .Z(n3444) );
  XOR U5039 ( .A(in[1311]), .B(n4261), .Z(n3873) );
  XNOR U5040 ( .A(in[1238]), .B(n3130), .Z(n3870) );
  NANDN U5041 ( .A(n3873), .B(n3870), .Z(n3131) );
  XNOR U5042 ( .A(n3444), .B(n3131), .Z(out[378]) );
  XOR U5043 ( .A(in[67]), .B(n4423), .Z(n3447) );
  XOR U5044 ( .A(in[1312]), .B(n4264), .Z(n3877) );
  XNOR U5045 ( .A(in[1239]), .B(n3132), .Z(n3874) );
  NANDN U5046 ( .A(n3877), .B(n3874), .Z(n3133) );
  XNOR U5047 ( .A(n3447), .B(n3133), .Z(out[379]) );
  ANDN U5048 ( .B(n3135), .A(n3134), .Z(n3136) );
  XOR U5049 ( .A(n3137), .B(n3136), .Z(out[37]) );
  XOR U5050 ( .A(in[68]), .B(n4426), .Z(n3450) );
  XOR U5051 ( .A(in[1313]), .B(n4267), .Z(n3881) );
  XNOR U5052 ( .A(in[1240]), .B(n3138), .Z(n3878) );
  NANDN U5053 ( .A(n3881), .B(n3878), .Z(n3139) );
  XNOR U5054 ( .A(n3450), .B(n3139), .Z(out[380]) );
  XOR U5055 ( .A(in[69]), .B(n4429), .Z(n3453) );
  XOR U5056 ( .A(in[1314]), .B(n4270), .Z(n3885) );
  XNOR U5057 ( .A(in[1241]), .B(n3140), .Z(n3882) );
  NANDN U5058 ( .A(n3885), .B(n3882), .Z(n3141) );
  XNOR U5059 ( .A(n3453), .B(n3141), .Z(out[381]) );
  XOR U5060 ( .A(in[70]), .B(n4432), .Z(n3460) );
  XOR U5061 ( .A(in[1315]), .B(n3142), .Z(n3889) );
  XNOR U5062 ( .A(in[1242]), .B(n3143), .Z(n3886) );
  NANDN U5063 ( .A(n3889), .B(n3886), .Z(n3144) );
  XOR U5064 ( .A(n3460), .B(n3144), .Z(out[382]) );
  XOR U5065 ( .A(in[71]), .B(n4443), .Z(n3463) );
  XOR U5066 ( .A(in[1316]), .B(n4276), .Z(n3893) );
  XNOR U5067 ( .A(in[1243]), .B(n3145), .Z(n3890) );
  NANDN U5068 ( .A(n3893), .B(n3890), .Z(n3146) );
  XNOR U5069 ( .A(n3463), .B(n3146), .Z(out[383]) );
  XOR U5070 ( .A(in[497]), .B(n4137), .Z(n3465) );
  XOR U5071 ( .A(in[498]), .B(n4141), .Z(n3467) );
  ANDN U5072 ( .B(n3619), .A(n3147), .Z(n3148) );
  XNOR U5073 ( .A(n3467), .B(n3148), .Z(out[385]) );
  XOR U5074 ( .A(in[499]), .B(n4145), .Z(n3469) );
  ANDN U5075 ( .B(n3623), .A(n3149), .Z(n3150) );
  XNOR U5076 ( .A(n3469), .B(n3150), .Z(out[386]) );
  XOR U5077 ( .A(in[500]), .B(n4149), .Z(n3471) );
  ANDN U5078 ( .B(n3627), .A(n3151), .Z(n3152) );
  XNOR U5079 ( .A(n3471), .B(n3152), .Z(out[387]) );
  XOR U5080 ( .A(in[501]), .B(n4153), .Z(n3473) );
  XOR U5081 ( .A(in[502]), .B(n4163), .Z(n3474) );
  NOR U5082 ( .A(n3154), .B(n3153), .Z(n3155) );
  XOR U5083 ( .A(n3156), .B(n3155), .Z(out[38]) );
  XOR U5084 ( .A(in[503]), .B(n4167), .Z(n3475) );
  XOR U5085 ( .A(in[504]), .B(n4171), .Z(n3476) );
  XOR U5086 ( .A(in[505]), .B(n4175), .Z(n3481) );
  XOR U5087 ( .A(in[506]), .B(n3899), .Z(n3482) );
  NOR U5088 ( .A(n3655), .B(n3291), .Z(n3157) );
  XNOR U5089 ( .A(n3482), .B(n3157), .Z(out[393]) );
  XOR U5090 ( .A(in[507]), .B(n3903), .Z(n3484) );
  NOR U5091 ( .A(n3659), .B(n3294), .Z(n3158) );
  XNOR U5092 ( .A(n3484), .B(n3158), .Z(out[394]) );
  XOR U5093 ( .A(in[508]), .B(n3907), .Z(n3486) );
  NOR U5094 ( .A(n3663), .B(n3297), .Z(n3159) );
  XNOR U5095 ( .A(n3486), .B(n3159), .Z(out[395]) );
  XOR U5096 ( .A(in[509]), .B(n3911), .Z(n3488) );
  NOR U5097 ( .A(n3667), .B(n3304), .Z(n3160) );
  XNOR U5098 ( .A(n3488), .B(n3160), .Z(out[396]) );
  XOR U5099 ( .A(in[510]), .B(n3915), .Z(n3490) );
  NOR U5100 ( .A(n3671), .B(n3307), .Z(n3161) );
  XNOR U5101 ( .A(n3490), .B(n3161), .Z(out[397]) );
  XOR U5102 ( .A(in[511]), .B(n3919), .Z(n3492) );
  NOR U5103 ( .A(n3679), .B(n3310), .Z(n3162) );
  XNOR U5104 ( .A(n3492), .B(n3162), .Z(out[398]) );
  XOR U5105 ( .A(in[448]), .B(n3923), .Z(n3494) );
  NOR U5106 ( .A(n3683), .B(n3313), .Z(n3163) );
  XNOR U5107 ( .A(n3494), .B(n3163), .Z(out[399]) );
  ANDN U5108 ( .B(n3165), .A(n3164), .Z(n3166) );
  XOR U5109 ( .A(n3167), .B(n3166), .Z(out[39]) );
  OR U5110 ( .A(n4069), .B(n3168), .Z(n3169) );
  XNOR U5111 ( .A(n4068), .B(n3169), .Z(out[3]) );
  XOR U5112 ( .A(in[449]), .B(n3927), .Z(n3496) );
  NOR U5113 ( .A(n3687), .B(n3316), .Z(n3170) );
  XNOR U5114 ( .A(n3496), .B(n3170), .Z(out[400]) );
  XOR U5115 ( .A(n3171), .B(in[450]), .Z(n3498) );
  NOR U5116 ( .A(n3691), .B(n3319), .Z(n3172) );
  XOR U5117 ( .A(n3498), .B(n3172), .Z(out[401]) );
  XOR U5118 ( .A(n3173), .B(in[451]), .Z(n3503) );
  NOR U5119 ( .A(n3695), .B(n3321), .Z(n3174) );
  XOR U5120 ( .A(n3503), .B(n3174), .Z(out[402]) );
  XOR U5121 ( .A(n3175), .B(in[452]), .Z(n3504) );
  NOR U5122 ( .A(n3699), .B(n3323), .Z(n3176) );
  XOR U5123 ( .A(n3504), .B(n3176), .Z(out[403]) );
  XOR U5124 ( .A(n3177), .B(in[453]), .Z(n3505) );
  NOR U5125 ( .A(n3703), .B(n3325), .Z(n3178) );
  XOR U5126 ( .A(n3505), .B(n3178), .Z(out[404]) );
  XOR U5127 ( .A(n3179), .B(in[454]), .Z(n3506) );
  NOR U5128 ( .A(n3707), .B(n3327), .Z(n3180) );
  XOR U5129 ( .A(n3506), .B(n3180), .Z(out[405]) );
  XOR U5130 ( .A(n3181), .B(in[455]), .Z(n3507) );
  NOR U5131 ( .A(n3711), .B(n3333), .Z(n3182) );
  XOR U5132 ( .A(n3507), .B(n3182), .Z(out[406]) );
  XOR U5133 ( .A(n3183), .B(in[456]), .Z(n3508) );
  NOR U5134 ( .A(n3715), .B(n3335), .Z(n3184) );
  XOR U5135 ( .A(n3508), .B(n3184), .Z(out[407]) );
  XOR U5136 ( .A(in[457]), .B(n3185), .Z(n3509) );
  NOR U5137 ( .A(n3725), .B(n3337), .Z(n3186) );
  XOR U5138 ( .A(n3509), .B(n3186), .Z(out[408]) );
  XOR U5139 ( .A(n3187), .B(in[458]), .Z(n3510) );
  NOR U5140 ( .A(n3729), .B(n3339), .Z(n3188) );
  XOR U5141 ( .A(n3510), .B(n3188), .Z(out[409]) );
  ANDN U5142 ( .B(n3190), .A(n3189), .Z(n3191) );
  XNOR U5143 ( .A(n3192), .B(n3191), .Z(out[40]) );
  XOR U5144 ( .A(n3971), .B(in[459]), .Z(n3511) );
  NOR U5145 ( .A(n3733), .B(n3341), .Z(n3193) );
  XNOR U5146 ( .A(n3511), .B(n3193), .Z(out[410]) );
  XOR U5147 ( .A(in[460]), .B(n3194), .Z(n3513) );
  NOR U5148 ( .A(n3737), .B(n3343), .Z(n3195) );
  XOR U5149 ( .A(n3513), .B(n3195), .Z(out[411]) );
  XOR U5150 ( .A(in[461]), .B(n3196), .Z(n3345) );
  NOR U5151 ( .A(n3197), .B(n3741), .Z(n3198) );
  XOR U5152 ( .A(n3345), .B(n3198), .Z(out[412]) );
  XOR U5153 ( .A(in[462]), .B(n3199), .Z(n3348) );
  NOR U5154 ( .A(n3200), .B(n3745), .Z(n3201) );
  XOR U5155 ( .A(n3348), .B(n3201), .Z(out[413]) );
  XOR U5156 ( .A(in[463]), .B(n3202), .Z(n3351) );
  NOR U5157 ( .A(n3203), .B(n3749), .Z(n3204) );
  XOR U5158 ( .A(n3351), .B(n3204), .Z(out[414]) );
  XOR U5159 ( .A(in[464]), .B(n3205), .Z(n3354) );
  NOR U5160 ( .A(n3206), .B(n3753), .Z(n3207) );
  XOR U5161 ( .A(n3354), .B(n3207), .Z(out[415]) );
  XOR U5162 ( .A(in[465]), .B(n3208), .Z(n3361) );
  NOR U5163 ( .A(n3209), .B(n3757), .Z(n3210) );
  XOR U5164 ( .A(n3361), .B(n3210), .Z(out[416]) );
  XOR U5165 ( .A(in[466]), .B(n4002), .Z(n3364) );
  NOR U5166 ( .A(n3211), .B(n3761), .Z(n3212) );
  XOR U5167 ( .A(n3364), .B(n3212), .Z(out[417]) );
  XOR U5168 ( .A(in[467]), .B(n3213), .Z(n3367) );
  NOR U5169 ( .A(n3214), .B(n3769), .Z(n3215) );
  XOR U5170 ( .A(n3367), .B(n3215), .Z(out[418]) );
  XOR U5171 ( .A(in[468]), .B(n3216), .Z(n3370) );
  NOR U5172 ( .A(n3217), .B(n3773), .Z(n3218) );
  XOR U5173 ( .A(n3370), .B(n3218), .Z(out[419]) );
  AND U5174 ( .A(n3220), .B(n3219), .Z(n3221) );
  XNOR U5175 ( .A(n3222), .B(n3221), .Z(out[41]) );
  XOR U5176 ( .A(in[469]), .B(n4014), .Z(n3539) );
  NOR U5177 ( .A(n3223), .B(n3777), .Z(n3224) );
  XNOR U5178 ( .A(n3539), .B(n3224), .Z(out[420]) );
  XOR U5179 ( .A(in[470]), .B(n4018), .Z(n3542) );
  NOR U5180 ( .A(n3225), .B(n3781), .Z(n3226) );
  XNOR U5181 ( .A(n3542), .B(n3226), .Z(out[421]) );
  XOR U5182 ( .A(in[471]), .B(n4022), .Z(n3549) );
  NOR U5183 ( .A(n3227), .B(n3785), .Z(n3228) );
  XNOR U5184 ( .A(n3549), .B(n3228), .Z(out[422]) );
  XOR U5185 ( .A(in[472]), .B(n4030), .Z(n3552) );
  NOR U5186 ( .A(n3229), .B(n3789), .Z(n3230) );
  XNOR U5187 ( .A(n3552), .B(n3230), .Z(out[423]) );
  XOR U5188 ( .A(in[473]), .B(n4034), .Z(n3555) );
  ANDN U5189 ( .B(n3793), .A(n3231), .Z(n3232) );
  XNOR U5190 ( .A(n3555), .B(n3232), .Z(out[424]) );
  XOR U5191 ( .A(in[474]), .B(n4038), .Z(n3558) );
  ANDN U5192 ( .B(n3797), .A(n3233), .Z(n3234) );
  XNOR U5193 ( .A(n3558), .B(n3234), .Z(out[425]) );
  XOR U5194 ( .A(in[475]), .B(n4042), .Z(n3561) );
  ANDN U5195 ( .B(n3801), .A(n3235), .Z(n3236) );
  XNOR U5196 ( .A(n3561), .B(n3236), .Z(out[426]) );
  XOR U5197 ( .A(in[476]), .B(n4046), .Z(n3564) );
  ANDN U5198 ( .B(n3805), .A(n3237), .Z(n3238) );
  XNOR U5199 ( .A(n3564), .B(n3238), .Z(out[427]) );
  XOR U5200 ( .A(in[477]), .B(n4050), .Z(n3566) );
  ANDN U5201 ( .B(n3813), .A(n3239), .Z(n3240) );
  XNOR U5202 ( .A(n3566), .B(n3240), .Z(out[428]) );
  XOR U5203 ( .A(in[478]), .B(n4054), .Z(n3397) );
  ANDN U5204 ( .B(n3817), .A(n3241), .Z(n3242) );
  XOR U5205 ( .A(n3397), .B(n3242), .Z(out[429]) );
  AND U5206 ( .A(n3244), .B(n3243), .Z(n3245) );
  XNOR U5207 ( .A(n3246), .B(n3245), .Z(out[42]) );
  XOR U5208 ( .A(in[479]), .B(n4058), .Z(n3401) );
  ANDN U5209 ( .B(n3821), .A(n3247), .Z(n3248) );
  XOR U5210 ( .A(n3401), .B(n3248), .Z(out[430]) );
  XOR U5211 ( .A(in[480]), .B(n4062), .Z(n3405) );
  ANDN U5212 ( .B(n3825), .A(n3249), .Z(n3250) );
  XOR U5213 ( .A(n3405), .B(n3250), .Z(out[431]) );
  XOR U5214 ( .A(in[481]), .B(n4066), .Z(n3408) );
  ANDN U5215 ( .B(n3829), .A(n3251), .Z(n3252) );
  XOR U5216 ( .A(n3408), .B(n3252), .Z(out[432]) );
  XOR U5217 ( .A(in[482]), .B(n4074), .Z(n3411) );
  ANDN U5218 ( .B(n3833), .A(n3253), .Z(n3254) );
  XOR U5219 ( .A(n3411), .B(n3254), .Z(out[433]) );
  XOR U5220 ( .A(in[483]), .B(n4078), .Z(n3414) );
  XOR U5221 ( .A(in[484]), .B(n4082), .Z(n3417) );
  XOR U5222 ( .A(in[485]), .B(n4086), .Z(n3586) );
  XOR U5223 ( .A(in[486]), .B(n4089), .Z(n3588) );
  XOR U5224 ( .A(in[487]), .B(n4093), .Z(n3590) );
  XOR U5225 ( .A(in[488]), .B(n4097), .Z(n3592) );
  AND U5226 ( .A(n3256), .B(n3255), .Z(n3257) );
  XNOR U5227 ( .A(n3258), .B(n3257), .Z(out[43]) );
  XOR U5228 ( .A(in[489]), .B(n4101), .Z(n3594) );
  XOR U5229 ( .A(in[490]), .B(n4105), .Z(n3596) );
  XOR U5230 ( .A(in[491]), .B(n4109), .Z(n3602) );
  XOR U5231 ( .A(in[492]), .B(n4117), .Z(n3603) );
  XOR U5232 ( .A(in[493]), .B(n4121), .Z(n3604) );
  XOR U5233 ( .A(in[494]), .B(n4125), .Z(n3606) );
  XOR U5234 ( .A(in[495]), .B(n4129), .Z(n3608) );
  XOR U5235 ( .A(in[496]), .B(n4133), .Z(n3610) );
  XOR U5236 ( .A(in[886]), .B(n3259), .Z(n3613) );
  NAND U5237 ( .A(n3260), .B(n3465), .Z(n3261) );
  XOR U5238 ( .A(n3613), .B(n3261), .Z(out[448]) );
  XOR U5239 ( .A(in[887]), .B(n3262), .Z(n3617) );
  NANDN U5240 ( .A(n3263), .B(n3467), .Z(n3264) );
  XOR U5241 ( .A(n3617), .B(n3264), .Z(out[449]) );
  AND U5242 ( .A(n3266), .B(n3265), .Z(n3267) );
  XNOR U5243 ( .A(n3268), .B(n3267), .Z(out[44]) );
  XOR U5244 ( .A(in[888]), .B(n3269), .Z(n3621) );
  NANDN U5245 ( .A(n3270), .B(n3469), .Z(n3271) );
  XOR U5246 ( .A(n3621), .B(n3271), .Z(out[450]) );
  XOR U5247 ( .A(in[889]), .B(n3272), .Z(n3625) );
  NANDN U5248 ( .A(n3273), .B(n3471), .Z(n3274) );
  XOR U5249 ( .A(n3625), .B(n3274), .Z(out[451]) );
  XOR U5250 ( .A(in[890]), .B(n3275), .Z(n3633) );
  NANDN U5251 ( .A(n3473), .B(n3276), .Z(n3277) );
  XOR U5252 ( .A(n3633), .B(n3277), .Z(out[452]) );
  XOR U5253 ( .A(in[891]), .B(n3278), .Z(n3637) );
  NANDN U5254 ( .A(n3474), .B(n3279), .Z(n3280) );
  XNOR U5255 ( .A(n3637), .B(n3280), .Z(out[453]) );
  XOR U5256 ( .A(in[892]), .B(n3281), .Z(n3641) );
  NANDN U5257 ( .A(n3475), .B(n3282), .Z(n3283) );
  XNOR U5258 ( .A(n3641), .B(n3283), .Z(out[454]) );
  XOR U5259 ( .A(in[893]), .B(n3284), .Z(n3645) );
  NANDN U5260 ( .A(n3476), .B(n3285), .Z(n3286) );
  XNOR U5261 ( .A(n3645), .B(n3286), .Z(out[455]) );
  XOR U5262 ( .A(in[894]), .B(n3287), .Z(n3649) );
  NANDN U5263 ( .A(n3481), .B(n3288), .Z(n3289) );
  XOR U5264 ( .A(n3649), .B(n3289), .Z(out[456]) );
  IV U5265 ( .A(n3290), .Z(n3900) );
  XOR U5266 ( .A(in[895]), .B(n3900), .Z(n3652) );
  NAND U5267 ( .A(n3291), .B(n3482), .Z(n3292) );
  XNOR U5268 ( .A(n3652), .B(n3292), .Z(out[457]) );
  IV U5269 ( .A(n3293), .Z(n3904) );
  XOR U5270 ( .A(in[832]), .B(n3904), .Z(n3656) );
  NAND U5271 ( .A(n3294), .B(n3484), .Z(n3295) );
  XNOR U5272 ( .A(n3656), .B(n3295), .Z(out[458]) );
  IV U5273 ( .A(n3296), .Z(n3908) );
  XOR U5274 ( .A(in[833]), .B(n3908), .Z(n3660) );
  NAND U5275 ( .A(n3297), .B(n3486), .Z(n3298) );
  XNOR U5276 ( .A(n3660), .B(n3298), .Z(out[459]) );
  AND U5277 ( .A(n3300), .B(n3299), .Z(n3301) );
  XNOR U5278 ( .A(n3302), .B(n3301), .Z(out[45]) );
  IV U5279 ( .A(n3303), .Z(n3912) );
  XOR U5280 ( .A(in[834]), .B(n3912), .Z(n3664) );
  NAND U5281 ( .A(n3304), .B(n3488), .Z(n3305) );
  XNOR U5282 ( .A(n3664), .B(n3305), .Z(out[460]) );
  IV U5283 ( .A(n3306), .Z(n3916) );
  XOR U5284 ( .A(in[835]), .B(n3916), .Z(n3668) );
  NAND U5285 ( .A(n3307), .B(n3490), .Z(n3308) );
  XNOR U5286 ( .A(n3668), .B(n3308), .Z(out[461]) );
  IV U5287 ( .A(n3309), .Z(n3920) );
  XOR U5288 ( .A(in[836]), .B(n3920), .Z(n3676) );
  NAND U5289 ( .A(n3310), .B(n3492), .Z(n3311) );
  XNOR U5290 ( .A(n3676), .B(n3311), .Z(out[462]) );
  IV U5291 ( .A(n3312), .Z(n3924) );
  XOR U5292 ( .A(in[837]), .B(n3924), .Z(n3680) );
  NAND U5293 ( .A(n3313), .B(n3494), .Z(n3314) );
  XNOR U5294 ( .A(n3680), .B(n3314), .Z(out[463]) );
  IV U5295 ( .A(n3315), .Z(n3928) );
  XOR U5296 ( .A(in[838]), .B(n3928), .Z(n3684) );
  NAND U5297 ( .A(n3316), .B(n3496), .Z(n3317) );
  XNOR U5298 ( .A(n3684), .B(n3317), .Z(out[464]) );
  XNOR U5299 ( .A(in[839]), .B(n3318), .Z(n3688) );
  NANDN U5300 ( .A(n3498), .B(n3319), .Z(n3320) );
  XNOR U5301 ( .A(n3688), .B(n3320), .Z(out[465]) );
  XNOR U5302 ( .A(in[840]), .B(n3935), .Z(n3692) );
  NANDN U5303 ( .A(n3503), .B(n3321), .Z(n3322) );
  XNOR U5304 ( .A(n3692), .B(n3322), .Z(out[466]) );
  XNOR U5305 ( .A(in[841]), .B(n3942), .Z(n3696) );
  NANDN U5306 ( .A(n3504), .B(n3323), .Z(n3324) );
  XNOR U5307 ( .A(n3696), .B(n3324), .Z(out[467]) );
  XNOR U5308 ( .A(in[842]), .B(n3946), .Z(n3700) );
  NANDN U5309 ( .A(n3505), .B(n3325), .Z(n3326) );
  XNOR U5310 ( .A(n3700), .B(n3326), .Z(out[468]) );
  XNOR U5311 ( .A(in[843]), .B(n3950), .Z(n3704) );
  NANDN U5312 ( .A(n3506), .B(n3327), .Z(n3328) );
  XNOR U5313 ( .A(n3704), .B(n3328), .Z(out[469]) );
  AND U5314 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U5315 ( .A(n3332), .B(n3331), .Z(out[46]) );
  XNOR U5316 ( .A(in[844]), .B(n3954), .Z(n3708) );
  NANDN U5317 ( .A(n3507), .B(n3333), .Z(n3334) );
  XNOR U5318 ( .A(n3708), .B(n3334), .Z(out[470]) );
  XNOR U5319 ( .A(in[845]), .B(n3958), .Z(n3712) );
  NANDN U5320 ( .A(n3508), .B(n3335), .Z(n3336) );
  XNOR U5321 ( .A(n3712), .B(n3336), .Z(out[471]) );
  XNOR U5322 ( .A(in[846]), .B(n3962), .Z(n3722) );
  NANDN U5323 ( .A(n3509), .B(n3337), .Z(n3338) );
  XNOR U5324 ( .A(n3722), .B(n3338), .Z(out[472]) );
  XNOR U5325 ( .A(in[847]), .B(n3966), .Z(n3726) );
  NANDN U5326 ( .A(n3510), .B(n3339), .Z(n3340) );
  XNOR U5327 ( .A(n3726), .B(n3340), .Z(out[473]) );
  XNOR U5328 ( .A(in[848]), .B(n3970), .Z(n3730) );
  NAND U5329 ( .A(n3341), .B(n3511), .Z(n3342) );
  XNOR U5330 ( .A(n3730), .B(n3342), .Z(out[474]) );
  XNOR U5331 ( .A(in[849]), .B(n3974), .Z(n3734) );
  NANDN U5332 ( .A(n3513), .B(n3343), .Z(n3344) );
  XNOR U5333 ( .A(n3734), .B(n3344), .Z(out[475]) );
  XNOR U5334 ( .A(in[850]), .B(n3978), .Z(n3738) );
  IV U5335 ( .A(n3345), .Z(n3518) );
  NANDN U5336 ( .A(n3346), .B(n3518), .Z(n3347) );
  XNOR U5337 ( .A(n3738), .B(n3347), .Z(out[476]) );
  XOR U5338 ( .A(in[851]), .B(n3985), .Z(n3520) );
  IV U5339 ( .A(n3348), .Z(n3521) );
  NANDN U5340 ( .A(n3349), .B(n3521), .Z(n3350) );
  XNOR U5341 ( .A(n3520), .B(n3350), .Z(out[477]) );
  XOR U5342 ( .A(in[852]), .B(n3989), .Z(n3523) );
  IV U5343 ( .A(n3351), .Z(n3524) );
  NANDN U5344 ( .A(n3352), .B(n3524), .Z(n3353) );
  XNOR U5345 ( .A(n3523), .B(n3353), .Z(out[478]) );
  XOR U5346 ( .A(in[853]), .B(n3993), .Z(n3750) );
  IV U5347 ( .A(n3354), .Z(n3526) );
  NANDN U5348 ( .A(n3355), .B(n3526), .Z(n3356) );
  XOR U5349 ( .A(n3750), .B(n3356), .Z(out[479]) );
  ANDN U5350 ( .B(n3358), .A(n3357), .Z(n3359) );
  XNOR U5351 ( .A(n3360), .B(n3359), .Z(out[47]) );
  XOR U5352 ( .A(in[854]), .B(n3997), .Z(n3528) );
  IV U5353 ( .A(n3361), .Z(n3529) );
  NANDN U5354 ( .A(n3362), .B(n3529), .Z(n3363) );
  XNOR U5355 ( .A(n3528), .B(n3363), .Z(out[480]) );
  XOR U5356 ( .A(in[855]), .B(n4001), .Z(n3531) );
  IV U5357 ( .A(n3364), .Z(n3532) );
  NANDN U5358 ( .A(n3365), .B(n3532), .Z(n3366) );
  XNOR U5359 ( .A(n3531), .B(n3366), .Z(out[481]) );
  XOR U5360 ( .A(in[856]), .B(n4005), .Z(n3766) );
  IV U5361 ( .A(n3367), .Z(n3534) );
  NANDN U5362 ( .A(n3368), .B(n3534), .Z(n3369) );
  XOR U5363 ( .A(n3766), .B(n3369), .Z(out[482]) );
  XOR U5364 ( .A(in[857]), .B(n4009), .Z(n3770) );
  IV U5365 ( .A(n3370), .Z(n3536) );
  NANDN U5366 ( .A(n3371), .B(n3536), .Z(n3372) );
  XOR U5367 ( .A(n3770), .B(n3372), .Z(out[483]) );
  XOR U5368 ( .A(in[858]), .B(n4013), .Z(n3538) );
  NANDN U5369 ( .A(n3373), .B(n3539), .Z(n3374) );
  XNOR U5370 ( .A(n3538), .B(n3374), .Z(out[484]) );
  XOR U5371 ( .A(in[859]), .B(n4017), .Z(n3541) );
  NANDN U5372 ( .A(n3375), .B(n3542), .Z(n3376) );
  XNOR U5373 ( .A(n3541), .B(n3376), .Z(out[485]) );
  XOR U5374 ( .A(in[860]), .B(n4021), .Z(n3548) );
  NANDN U5375 ( .A(n3377), .B(n3549), .Z(n3378) );
  XNOR U5376 ( .A(n3548), .B(n3378), .Z(out[486]) );
  XOR U5377 ( .A(in[861]), .B(n4029), .Z(n3551) );
  NANDN U5378 ( .A(n3379), .B(n3552), .Z(n3380) );
  XNOR U5379 ( .A(n3551), .B(n3380), .Z(out[487]) );
  XOR U5380 ( .A(in[862]), .B(n4033), .Z(n3554) );
  NANDN U5381 ( .A(n3381), .B(n3555), .Z(n3382) );
  XNOR U5382 ( .A(n3554), .B(n3382), .Z(out[488]) );
  XOR U5383 ( .A(in[863]), .B(n4037), .Z(n3557) );
  NANDN U5384 ( .A(n3383), .B(n3558), .Z(n3384) );
  XNOR U5385 ( .A(n3557), .B(n3384), .Z(out[489]) );
  AND U5386 ( .A(n3386), .B(n3385), .Z(n3387) );
  XNOR U5387 ( .A(n3388), .B(n3387), .Z(out[48]) );
  XOR U5388 ( .A(in[864]), .B(n4041), .Z(n3560) );
  NANDN U5389 ( .A(n3389), .B(n3561), .Z(n3390) );
  XNOR U5390 ( .A(n3560), .B(n3390), .Z(out[490]) );
  XOR U5391 ( .A(in[865]), .B(n4045), .Z(n3563) );
  NANDN U5392 ( .A(n3391), .B(n3564), .Z(n3392) );
  XNOR U5393 ( .A(n3563), .B(n3392), .Z(out[491]) );
  XNOR U5394 ( .A(n3393), .B(in[866]), .Z(n3811) );
  NANDN U5395 ( .A(n3394), .B(n3566), .Z(n3395) );
  XNOR U5396 ( .A(n3811), .B(n3395), .Z(out[492]) );
  XNOR U5397 ( .A(n3396), .B(in[867]), .Z(n3815) );
  IV U5398 ( .A(n3397), .Z(n3568) );
  NANDN U5399 ( .A(n3398), .B(n3568), .Z(n3399) );
  XNOR U5400 ( .A(n3815), .B(n3399), .Z(out[493]) );
  XNOR U5401 ( .A(n3400), .B(in[868]), .Z(n3819) );
  IV U5402 ( .A(n3401), .Z(n3570) );
  NANDN U5403 ( .A(n3402), .B(n3570), .Z(n3403) );
  XNOR U5404 ( .A(n3819), .B(n3403), .Z(out[494]) );
  XNOR U5405 ( .A(n3404), .B(in[869]), .Z(n3823) );
  IV U5406 ( .A(n3405), .Z(n3572) );
  NANDN U5407 ( .A(n3406), .B(n3572), .Z(n3407) );
  XNOR U5408 ( .A(n3823), .B(n3407), .Z(out[495]) );
  XOR U5409 ( .A(in[870]), .B(n4065), .Z(n3827) );
  IV U5410 ( .A(n3408), .Z(n3578) );
  NANDN U5411 ( .A(n3409), .B(n3578), .Z(n3410) );
  XOR U5412 ( .A(n3827), .B(n3410), .Z(out[496]) );
  XOR U5413 ( .A(in[871]), .B(n4073), .Z(n3831) );
  IV U5414 ( .A(n3411), .Z(n3580) );
  NANDN U5415 ( .A(n3412), .B(n3580), .Z(n3413) );
  XOR U5416 ( .A(n3831), .B(n3413), .Z(out[497]) );
  XOR U5417 ( .A(in[872]), .B(n4077), .Z(n3835) );
  IV U5418 ( .A(n3414), .Z(n3582) );
  NANDN U5419 ( .A(n3415), .B(n3582), .Z(n3416) );
  XOR U5420 ( .A(n3835), .B(n3416), .Z(out[498]) );
  XOR U5421 ( .A(in[873]), .B(n4081), .Z(n3839) );
  IV U5422 ( .A(n3417), .Z(n3584) );
  NANDN U5423 ( .A(n3418), .B(n3584), .Z(n3419) );
  XOR U5424 ( .A(n3839), .B(n3419), .Z(out[499]) );
  ANDN U5425 ( .B(n3421), .A(n3420), .Z(n3422) );
  XNOR U5426 ( .A(n3423), .B(n3422), .Z(out[49]) );
  OR U5427 ( .A(n4113), .B(n3424), .Z(n3425) );
  XNOR U5428 ( .A(n4112), .B(n3425), .Z(out[4]) );
  XOR U5429 ( .A(in[874]), .B(n4085), .Z(n3843) );
  NAND U5430 ( .A(n3426), .B(n3586), .Z(n3427) );
  XOR U5431 ( .A(n3843), .B(n3427), .Z(out[500]) );
  XOR U5432 ( .A(in[875]), .B(n3428), .Z(n3847) );
  NAND U5433 ( .A(n3429), .B(n3588), .Z(n3430) );
  XOR U5434 ( .A(n3847), .B(n3430), .Z(out[501]) );
  XOR U5435 ( .A(in[876]), .B(n3431), .Z(n3855) );
  NAND U5436 ( .A(n3432), .B(n3590), .Z(n3433) );
  XOR U5437 ( .A(n3855), .B(n3433), .Z(out[502]) );
  XOR U5438 ( .A(in[877]), .B(n3434), .Z(n3859) );
  NAND U5439 ( .A(n3435), .B(n3592), .Z(n3436) );
  XOR U5440 ( .A(n3859), .B(n3436), .Z(out[503]) );
  XOR U5441 ( .A(in[878]), .B(n3437), .Z(n3863) );
  NAND U5442 ( .A(n3438), .B(n3594), .Z(n3439) );
  XOR U5443 ( .A(n3863), .B(n3439), .Z(out[504]) );
  XOR U5444 ( .A(in[879]), .B(n3440), .Z(n3867) );
  NAND U5445 ( .A(n3441), .B(n3596), .Z(n3442) );
  XOR U5446 ( .A(n3867), .B(n3442), .Z(out[505]) );
  XOR U5447 ( .A(in[880]), .B(n3443), .Z(n3871) );
  NANDN U5448 ( .A(n3602), .B(n3444), .Z(n3445) );
  XOR U5449 ( .A(n3871), .B(n3445), .Z(out[506]) );
  XOR U5450 ( .A(in[881]), .B(n3446), .Z(n3875) );
  NANDN U5451 ( .A(n3603), .B(n3447), .Z(n3448) );
  XOR U5452 ( .A(n3875), .B(n3448), .Z(out[507]) );
  XOR U5453 ( .A(in[882]), .B(n3449), .Z(n3879) );
  NAND U5454 ( .A(n3450), .B(n3604), .Z(n3451) );
  XOR U5455 ( .A(n3879), .B(n3451), .Z(out[508]) );
  XOR U5456 ( .A(in[883]), .B(n3452), .Z(n3883) );
  NAND U5457 ( .A(n3453), .B(n3606), .Z(n3454) );
  XOR U5458 ( .A(n3883), .B(n3454), .Z(out[509]) );
  ANDN U5459 ( .B(n3456), .A(n3455), .Z(n3457) );
  XNOR U5460 ( .A(n3458), .B(n3457), .Z(out[50]) );
  XOR U5461 ( .A(in[884]), .B(n3459), .Z(n3887) );
  NANDN U5462 ( .A(n3460), .B(n3608), .Z(n3461) );
  XOR U5463 ( .A(n3887), .B(n3461), .Z(out[510]) );
  XOR U5464 ( .A(in[885]), .B(n3462), .Z(n3891) );
  NAND U5465 ( .A(n3463), .B(n3610), .Z(n3464) );
  XOR U5466 ( .A(n3891), .B(n3464), .Z(out[511]) );
  NANDN U5467 ( .A(n3465), .B(n3613), .Z(n3466) );
  XNOR U5468 ( .A(n3612), .B(n3466), .Z(out[512]) );
  NANDN U5469 ( .A(n3467), .B(n3617), .Z(n3468) );
  XNOR U5470 ( .A(n3616), .B(n3468), .Z(out[513]) );
  NANDN U5471 ( .A(n3469), .B(n3621), .Z(n3470) );
  XNOR U5472 ( .A(n3620), .B(n3470), .Z(out[514]) );
  NANDN U5473 ( .A(n3471), .B(n3625), .Z(n3472) );
  XNOR U5474 ( .A(n3624), .B(n3472), .Z(out[515]) );
  ANDN U5475 ( .B(n3478), .A(n3477), .Z(n3479) );
  XNOR U5476 ( .A(n3480), .B(n3479), .Z(out[51]) );
  OR U5477 ( .A(n3652), .B(n3482), .Z(n3483) );
  XOR U5478 ( .A(n3653), .B(n3483), .Z(out[521]) );
  OR U5479 ( .A(n3656), .B(n3484), .Z(n3485) );
  XOR U5480 ( .A(n3657), .B(n3485), .Z(out[522]) );
  OR U5481 ( .A(n3660), .B(n3486), .Z(n3487) );
  XOR U5482 ( .A(n3661), .B(n3487), .Z(out[523]) );
  OR U5483 ( .A(n3664), .B(n3488), .Z(n3489) );
  XOR U5484 ( .A(n3665), .B(n3489), .Z(out[524]) );
  OR U5485 ( .A(n3668), .B(n3490), .Z(n3491) );
  XOR U5486 ( .A(n3669), .B(n3491), .Z(out[525]) );
  OR U5487 ( .A(n3676), .B(n3492), .Z(n3493) );
  XOR U5488 ( .A(n3677), .B(n3493), .Z(out[526]) );
  OR U5489 ( .A(n3680), .B(n3494), .Z(n3495) );
  XOR U5490 ( .A(n3681), .B(n3495), .Z(out[527]) );
  OR U5491 ( .A(n3684), .B(n3496), .Z(n3497) );
  XOR U5492 ( .A(n3685), .B(n3497), .Z(out[528]) );
  ANDN U5493 ( .B(n3500), .A(n3499), .Z(n3501) );
  XNOR U5494 ( .A(n3502), .B(n3501), .Z(out[52]) );
  OR U5495 ( .A(n3730), .B(n3511), .Z(n3512) );
  XOR U5496 ( .A(n3731), .B(n3512), .Z(out[538]) );
  ANDN U5497 ( .B(n3515), .A(n3514), .Z(n3516) );
  XNOR U5498 ( .A(n3517), .B(n3516), .Z(out[53]) );
  OR U5499 ( .A(n3738), .B(n3518), .Z(n3519) );
  XOR U5500 ( .A(n3739), .B(n3519), .Z(out[540]) );
  IV U5501 ( .A(n3520), .Z(n3742) );
  NANDN U5502 ( .A(n3521), .B(n3742), .Z(n3522) );
  XOR U5503 ( .A(n3743), .B(n3522), .Z(out[541]) );
  IV U5504 ( .A(n3523), .Z(n3746) );
  NANDN U5505 ( .A(n3524), .B(n3746), .Z(n3525) );
  XOR U5506 ( .A(n3747), .B(n3525), .Z(out[542]) );
  NANDN U5507 ( .A(n3526), .B(n3750), .Z(n3527) );
  XOR U5508 ( .A(n3751), .B(n3527), .Z(out[543]) );
  IV U5509 ( .A(n3528), .Z(n3754) );
  NANDN U5510 ( .A(n3529), .B(n3754), .Z(n3530) );
  XOR U5511 ( .A(n3755), .B(n3530), .Z(out[544]) );
  IV U5512 ( .A(n3531), .Z(n3758) );
  NANDN U5513 ( .A(n3532), .B(n3758), .Z(n3533) );
  XOR U5514 ( .A(n3759), .B(n3533), .Z(out[545]) );
  NANDN U5515 ( .A(n3534), .B(n3766), .Z(n3535) );
  XOR U5516 ( .A(n3767), .B(n3535), .Z(out[546]) );
  NANDN U5517 ( .A(n3536), .B(n3770), .Z(n3537) );
  XOR U5518 ( .A(n3771), .B(n3537), .Z(out[547]) );
  IV U5519 ( .A(n3538), .Z(n3774) );
  NANDN U5520 ( .A(n3539), .B(n3774), .Z(n3540) );
  XOR U5521 ( .A(n3775), .B(n3540), .Z(out[548]) );
  IV U5522 ( .A(n3541), .Z(n3778) );
  NANDN U5523 ( .A(n3542), .B(n3778), .Z(n3543) );
  XOR U5524 ( .A(n3779), .B(n3543), .Z(out[549]) );
  ANDN U5525 ( .B(n3545), .A(n3544), .Z(n3546) );
  XNOR U5526 ( .A(n3547), .B(n3546), .Z(out[54]) );
  IV U5527 ( .A(n3548), .Z(n3782) );
  NANDN U5528 ( .A(n3549), .B(n3782), .Z(n3550) );
  XOR U5529 ( .A(n3783), .B(n3550), .Z(out[550]) );
  IV U5530 ( .A(n3551), .Z(n3786) );
  NANDN U5531 ( .A(n3552), .B(n3786), .Z(n3553) );
  XOR U5532 ( .A(n3787), .B(n3553), .Z(out[551]) );
  IV U5533 ( .A(n3554), .Z(n3791) );
  NANDN U5534 ( .A(n3555), .B(n3791), .Z(n3556) );
  XNOR U5535 ( .A(n3790), .B(n3556), .Z(out[552]) );
  IV U5536 ( .A(n3557), .Z(n3795) );
  NANDN U5537 ( .A(n3558), .B(n3795), .Z(n3559) );
  XNOR U5538 ( .A(n3794), .B(n3559), .Z(out[553]) );
  IV U5539 ( .A(n3560), .Z(n3799) );
  NANDN U5540 ( .A(n3561), .B(n3799), .Z(n3562) );
  XNOR U5541 ( .A(n3798), .B(n3562), .Z(out[554]) );
  IV U5542 ( .A(n3563), .Z(n3803) );
  NANDN U5543 ( .A(n3564), .B(n3803), .Z(n3565) );
  XNOR U5544 ( .A(n3802), .B(n3565), .Z(out[555]) );
  OR U5545 ( .A(n3811), .B(n3566), .Z(n3567) );
  XNOR U5546 ( .A(n3810), .B(n3567), .Z(out[556]) );
  OR U5547 ( .A(n3815), .B(n3568), .Z(n3569) );
  XNOR U5548 ( .A(n3814), .B(n3569), .Z(out[557]) );
  OR U5549 ( .A(n3819), .B(n3570), .Z(n3571) );
  XNOR U5550 ( .A(n3818), .B(n3571), .Z(out[558]) );
  OR U5551 ( .A(n3823), .B(n3572), .Z(n3573) );
  XNOR U5552 ( .A(n3822), .B(n3573), .Z(out[559]) );
  ANDN U5553 ( .B(n3575), .A(n3574), .Z(n3576) );
  XNOR U5554 ( .A(n3577), .B(n3576), .Z(out[55]) );
  NANDN U5555 ( .A(n3578), .B(n3827), .Z(n3579) );
  XNOR U5556 ( .A(n3826), .B(n3579), .Z(out[560]) );
  NANDN U5557 ( .A(n3580), .B(n3831), .Z(n3581) );
  XNOR U5558 ( .A(n3830), .B(n3581), .Z(out[561]) );
  NANDN U5559 ( .A(n3582), .B(n3835), .Z(n3583) );
  XNOR U5560 ( .A(n3834), .B(n3583), .Z(out[562]) );
  NANDN U5561 ( .A(n3584), .B(n3839), .Z(n3585) );
  XNOR U5562 ( .A(n3838), .B(n3585), .Z(out[563]) );
  NANDN U5563 ( .A(n3586), .B(n3843), .Z(n3587) );
  XNOR U5564 ( .A(n3842), .B(n3587), .Z(out[564]) );
  NANDN U5565 ( .A(n3588), .B(n3847), .Z(n3589) );
  XNOR U5566 ( .A(n3846), .B(n3589), .Z(out[565]) );
  NANDN U5567 ( .A(n3590), .B(n3855), .Z(n3591) );
  XNOR U5568 ( .A(n3854), .B(n3591), .Z(out[566]) );
  NANDN U5569 ( .A(n3592), .B(n3859), .Z(n3593) );
  XNOR U5570 ( .A(n3858), .B(n3593), .Z(out[567]) );
  NANDN U5571 ( .A(n3594), .B(n3863), .Z(n3595) );
  XNOR U5572 ( .A(n3862), .B(n3595), .Z(out[568]) );
  NANDN U5573 ( .A(n3596), .B(n3867), .Z(n3597) );
  XNOR U5574 ( .A(n3866), .B(n3597), .Z(out[569]) );
  ANDN U5575 ( .B(n3599), .A(n3598), .Z(n3600) );
  XNOR U5576 ( .A(n3601), .B(n3600), .Z(out[56]) );
  NANDN U5577 ( .A(n3604), .B(n3879), .Z(n3605) );
  XNOR U5578 ( .A(n3878), .B(n3605), .Z(out[572]) );
  NANDN U5579 ( .A(n3606), .B(n3883), .Z(n3607) );
  XNOR U5580 ( .A(n3882), .B(n3607), .Z(out[573]) );
  NANDN U5581 ( .A(n3608), .B(n3887), .Z(n3609) );
  XNOR U5582 ( .A(n3886), .B(n3609), .Z(out[574]) );
  NANDN U5583 ( .A(n3610), .B(n3891), .Z(n3611) );
  XNOR U5584 ( .A(n3890), .B(n3611), .Z(out[575]) );
  NOR U5585 ( .A(n3613), .B(n3612), .Z(n3614) );
  XOR U5586 ( .A(n3615), .B(n3614), .Z(out[576]) );
  NOR U5587 ( .A(n3617), .B(n3616), .Z(n3618) );
  XOR U5588 ( .A(n3619), .B(n3618), .Z(out[577]) );
  NOR U5589 ( .A(n3621), .B(n3620), .Z(n3622) );
  XOR U5590 ( .A(n3623), .B(n3622), .Z(out[578]) );
  NOR U5591 ( .A(n3625), .B(n3624), .Z(n3626) );
  XOR U5592 ( .A(n3627), .B(n3626), .Z(out[579]) );
  ANDN U5593 ( .B(n3629), .A(n3628), .Z(n3630) );
  XNOR U5594 ( .A(n3631), .B(n3630), .Z(out[57]) );
  NOR U5595 ( .A(n3633), .B(n3632), .Z(n3634) );
  XOR U5596 ( .A(n3635), .B(n3634), .Z(out[580]) );
  ANDN U5597 ( .B(n3637), .A(n3636), .Z(n3638) );
  XOR U5598 ( .A(n3639), .B(n3638), .Z(out[581]) );
  ANDN U5599 ( .B(n3641), .A(n3640), .Z(n3642) );
  XOR U5600 ( .A(n3643), .B(n3642), .Z(out[582]) );
  ANDN U5601 ( .B(n3645), .A(n3644), .Z(n3646) );
  XOR U5602 ( .A(n3647), .B(n3646), .Z(out[583]) );
  NOR U5603 ( .A(n3649), .B(n3648), .Z(n3650) );
  XOR U5604 ( .A(n3651), .B(n3650), .Z(out[584]) );
  AND U5605 ( .A(n3653), .B(n3652), .Z(n3654) );
  XNOR U5606 ( .A(n3655), .B(n3654), .Z(out[585]) );
  AND U5607 ( .A(n3657), .B(n3656), .Z(n3658) );
  XNOR U5608 ( .A(n3659), .B(n3658), .Z(out[586]) );
  AND U5609 ( .A(n3661), .B(n3660), .Z(n3662) );
  XNOR U5610 ( .A(n3663), .B(n3662), .Z(out[587]) );
  AND U5611 ( .A(n3665), .B(n3664), .Z(n3666) );
  XNOR U5612 ( .A(n3667), .B(n3666), .Z(out[588]) );
  AND U5613 ( .A(n3669), .B(n3668), .Z(n3670) );
  XNOR U5614 ( .A(n3671), .B(n3670), .Z(out[589]) );
  ANDN U5615 ( .B(n3673), .A(n3672), .Z(n3674) );
  XNOR U5616 ( .A(n3675), .B(n3674), .Z(out[58]) );
  AND U5617 ( .A(n3677), .B(n3676), .Z(n3678) );
  XNOR U5618 ( .A(n3679), .B(n3678), .Z(out[590]) );
  AND U5619 ( .A(n3681), .B(n3680), .Z(n3682) );
  XNOR U5620 ( .A(n3683), .B(n3682), .Z(out[591]) );
  AND U5621 ( .A(n3685), .B(n3684), .Z(n3686) );
  XNOR U5622 ( .A(n3687), .B(n3686), .Z(out[592]) );
  AND U5623 ( .A(n3689), .B(n3688), .Z(n3690) );
  XNOR U5624 ( .A(n3691), .B(n3690), .Z(out[593]) );
  AND U5625 ( .A(n3693), .B(n3692), .Z(n3694) );
  XNOR U5626 ( .A(n3695), .B(n3694), .Z(out[594]) );
  AND U5627 ( .A(n3697), .B(n3696), .Z(n3698) );
  XNOR U5628 ( .A(n3699), .B(n3698), .Z(out[595]) );
  AND U5629 ( .A(n3701), .B(n3700), .Z(n3702) );
  XNOR U5630 ( .A(n3703), .B(n3702), .Z(out[596]) );
  AND U5631 ( .A(n3705), .B(n3704), .Z(n3706) );
  XNOR U5632 ( .A(n3707), .B(n3706), .Z(out[597]) );
  AND U5633 ( .A(n3709), .B(n3708), .Z(n3710) );
  XNOR U5634 ( .A(n3711), .B(n3710), .Z(out[598]) );
  AND U5635 ( .A(n3713), .B(n3712), .Z(n3714) );
  XNOR U5636 ( .A(n3715), .B(n3714), .Z(out[599]) );
  ANDN U5637 ( .B(n3717), .A(n3716), .Z(n3718) );
  XNOR U5638 ( .A(n3719), .B(n3718), .Z(out[59]) );
  OR U5639 ( .A(n4157), .B(n3720), .Z(n3721) );
  XNOR U5640 ( .A(n4156), .B(n3721), .Z(out[5]) );
  AND U5641 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U5642 ( .A(n3725), .B(n3724), .Z(out[600]) );
  AND U5643 ( .A(n3727), .B(n3726), .Z(n3728) );
  XNOR U5644 ( .A(n3729), .B(n3728), .Z(out[601]) );
  AND U5645 ( .A(n3731), .B(n3730), .Z(n3732) );
  XNOR U5646 ( .A(n3733), .B(n3732), .Z(out[602]) );
  AND U5647 ( .A(n3735), .B(n3734), .Z(n3736) );
  XNOR U5648 ( .A(n3737), .B(n3736), .Z(out[603]) );
  AND U5649 ( .A(n3739), .B(n3738), .Z(n3740) );
  XNOR U5650 ( .A(n3741), .B(n3740), .Z(out[604]) );
  ANDN U5651 ( .B(n3743), .A(n3742), .Z(n3744) );
  XNOR U5652 ( .A(n3745), .B(n3744), .Z(out[605]) );
  ANDN U5653 ( .B(n3747), .A(n3746), .Z(n3748) );
  XNOR U5654 ( .A(n3749), .B(n3748), .Z(out[606]) );
  ANDN U5655 ( .B(n3751), .A(n3750), .Z(n3752) );
  XNOR U5656 ( .A(n3753), .B(n3752), .Z(out[607]) );
  ANDN U5657 ( .B(n3755), .A(n3754), .Z(n3756) );
  XNOR U5658 ( .A(n3757), .B(n3756), .Z(out[608]) );
  ANDN U5659 ( .B(n3759), .A(n3758), .Z(n3760) );
  XNOR U5660 ( .A(n3761), .B(n3760), .Z(out[609]) );
  ANDN U5661 ( .B(n3763), .A(n3762), .Z(n3764) );
  XNOR U5662 ( .A(n3765), .B(n3764), .Z(out[60]) );
  ANDN U5663 ( .B(n3767), .A(n3766), .Z(n3768) );
  XNOR U5664 ( .A(n3769), .B(n3768), .Z(out[610]) );
  ANDN U5665 ( .B(n3771), .A(n3770), .Z(n3772) );
  XNOR U5666 ( .A(n3773), .B(n3772), .Z(out[611]) );
  ANDN U5667 ( .B(n3775), .A(n3774), .Z(n3776) );
  XNOR U5668 ( .A(n3777), .B(n3776), .Z(out[612]) );
  ANDN U5669 ( .B(n3779), .A(n3778), .Z(n3780) );
  XNOR U5670 ( .A(n3781), .B(n3780), .Z(out[613]) );
  ANDN U5671 ( .B(n3783), .A(n3782), .Z(n3784) );
  XNOR U5672 ( .A(n3785), .B(n3784), .Z(out[614]) );
  ANDN U5673 ( .B(n3787), .A(n3786), .Z(n3788) );
  XNOR U5674 ( .A(n3789), .B(n3788), .Z(out[615]) );
  NOR U5675 ( .A(n3791), .B(n3790), .Z(n3792) );
  XOR U5676 ( .A(n3793), .B(n3792), .Z(out[616]) );
  NOR U5677 ( .A(n3795), .B(n3794), .Z(n3796) );
  XOR U5678 ( .A(n3797), .B(n3796), .Z(out[617]) );
  NOR U5679 ( .A(n3799), .B(n3798), .Z(n3800) );
  XOR U5680 ( .A(n3801), .B(n3800), .Z(out[618]) );
  NOR U5681 ( .A(n3803), .B(n3802), .Z(n3804) );
  XOR U5682 ( .A(n3805), .B(n3804), .Z(out[619]) );
  ANDN U5683 ( .B(n3807), .A(n3806), .Z(n3808) );
  XOR U5684 ( .A(n3809), .B(n3808), .Z(out[61]) );
  ANDN U5685 ( .B(n3811), .A(n3810), .Z(n3812) );
  XOR U5686 ( .A(n3813), .B(n3812), .Z(out[620]) );
  ANDN U5687 ( .B(n3815), .A(n3814), .Z(n3816) );
  XOR U5688 ( .A(n3817), .B(n3816), .Z(out[621]) );
  ANDN U5689 ( .B(n3819), .A(n3818), .Z(n3820) );
  XOR U5690 ( .A(n3821), .B(n3820), .Z(out[622]) );
  ANDN U5691 ( .B(n3823), .A(n3822), .Z(n3824) );
  XOR U5692 ( .A(n3825), .B(n3824), .Z(out[623]) );
  NOR U5693 ( .A(n3827), .B(n3826), .Z(n3828) );
  XOR U5694 ( .A(n3829), .B(n3828), .Z(out[624]) );
  NOR U5695 ( .A(n3831), .B(n3830), .Z(n3832) );
  XOR U5696 ( .A(n3833), .B(n3832), .Z(out[625]) );
  NOR U5697 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U5698 ( .A(n3837), .B(n3836), .Z(out[626]) );
  NOR U5699 ( .A(n3839), .B(n3838), .Z(n3840) );
  XOR U5700 ( .A(n3841), .B(n3840), .Z(out[627]) );
  NOR U5701 ( .A(n3843), .B(n3842), .Z(n3844) );
  XOR U5702 ( .A(n3845), .B(n3844), .Z(out[628]) );
  NOR U5703 ( .A(n3847), .B(n3846), .Z(n3848) );
  XOR U5704 ( .A(n3849), .B(n3848), .Z(out[629]) );
  ANDN U5705 ( .B(n3851), .A(n3850), .Z(n3852) );
  XOR U5706 ( .A(n3853), .B(n3852), .Z(out[62]) );
  NOR U5707 ( .A(n3855), .B(n3854), .Z(n3856) );
  XOR U5708 ( .A(n3857), .B(n3856), .Z(out[630]) );
  NOR U5709 ( .A(n3859), .B(n3858), .Z(n3860) );
  XOR U5710 ( .A(n3861), .B(n3860), .Z(out[631]) );
  NOR U5711 ( .A(n3863), .B(n3862), .Z(n3864) );
  XOR U5712 ( .A(n3865), .B(n3864), .Z(out[632]) );
  NOR U5713 ( .A(n3867), .B(n3866), .Z(n3868) );
  XOR U5714 ( .A(n3869), .B(n3868), .Z(out[633]) );
  NOR U5715 ( .A(n3871), .B(n3870), .Z(n3872) );
  XOR U5716 ( .A(n3873), .B(n3872), .Z(out[634]) );
  NOR U5717 ( .A(n3875), .B(n3874), .Z(n3876) );
  XOR U5718 ( .A(n3877), .B(n3876), .Z(out[635]) );
  NOR U5719 ( .A(n3879), .B(n3878), .Z(n3880) );
  XOR U5720 ( .A(n3881), .B(n3880), .Z(out[636]) );
  NOR U5721 ( .A(n3883), .B(n3882), .Z(n3884) );
  XOR U5722 ( .A(n3885), .B(n3884), .Z(out[637]) );
  NOR U5723 ( .A(n3887), .B(n3886), .Z(n3888) );
  XOR U5724 ( .A(n3889), .B(n3888), .Z(out[638]) );
  NOR U5725 ( .A(n3891), .B(n3890), .Z(n3892) );
  XOR U5726 ( .A(n3893), .B(n3892), .Z(out[639]) );
  ANDN U5727 ( .B(n3895), .A(n3894), .Z(n3896) );
  XOR U5728 ( .A(n3897), .B(n3896), .Z(out[63]) );
  XOR U5729 ( .A(in[302]), .B(n3898), .Z(n4179) );
  IV U5730 ( .A(n4179), .Z(n4334) );
  XOR U5731 ( .A(in[1146]), .B(n3899), .Z(n4706) );
  XOR U5732 ( .A(in[1535]), .B(n3900), .Z(n4708) );
  OR U5733 ( .A(n4706), .B(n4708), .Z(n3901) );
  XOR U5734 ( .A(n4334), .B(n3901), .Z(out[640]) );
  XOR U5735 ( .A(in[303]), .B(n3902), .Z(n4182) );
  IV U5736 ( .A(n4182), .Z(n4336) );
  XOR U5737 ( .A(in[1147]), .B(n3903), .Z(n4710) );
  XOR U5738 ( .A(in[1472]), .B(n3904), .Z(n4712) );
  OR U5739 ( .A(n4710), .B(n4712), .Z(n3905) );
  XOR U5740 ( .A(n4336), .B(n3905), .Z(out[641]) );
  XOR U5741 ( .A(in[304]), .B(n3906), .Z(n4185) );
  IV U5742 ( .A(n4185), .Z(n4342) );
  XOR U5743 ( .A(in[1148]), .B(n3907), .Z(n4714) );
  XOR U5744 ( .A(in[1473]), .B(n3908), .Z(n4716) );
  OR U5745 ( .A(n4714), .B(n4716), .Z(n3909) );
  XOR U5746 ( .A(n4342), .B(n3909), .Z(out[642]) );
  XOR U5747 ( .A(in[305]), .B(n3910), .Z(n4188) );
  IV U5748 ( .A(n4188), .Z(n4344) );
  XOR U5749 ( .A(in[1149]), .B(n3911), .Z(n4718) );
  XOR U5750 ( .A(in[1474]), .B(n3912), .Z(n4720) );
  OR U5751 ( .A(n4718), .B(n4720), .Z(n3913) );
  XOR U5752 ( .A(n4344), .B(n3913), .Z(out[643]) );
  XOR U5753 ( .A(in[306]), .B(n3914), .Z(n4191) );
  IV U5754 ( .A(n4191), .Z(n4346) );
  XOR U5755 ( .A(in[1150]), .B(n3915), .Z(n4730) );
  XOR U5756 ( .A(in[1475]), .B(n3916), .Z(n4732) );
  OR U5757 ( .A(n4730), .B(n4732), .Z(n3917) );
  XOR U5758 ( .A(n4346), .B(n3917), .Z(out[644]) );
  XOR U5759 ( .A(in[307]), .B(n3918), .Z(n4349) );
  XOR U5760 ( .A(in[1151]), .B(n3919), .Z(n4734) );
  XOR U5761 ( .A(in[1476]), .B(n3920), .Z(n4736) );
  OR U5762 ( .A(n4734), .B(n4736), .Z(n3921) );
  XOR U5763 ( .A(n4349), .B(n3921), .Z(out[645]) );
  XOR U5764 ( .A(in[308]), .B(n3922), .Z(n4352) );
  XOR U5765 ( .A(in[1088]), .B(n3923), .Z(n4738) );
  XOR U5766 ( .A(in[1477]), .B(n3924), .Z(n4740) );
  OR U5767 ( .A(n4738), .B(n4740), .Z(n3925) );
  XOR U5768 ( .A(n4352), .B(n3925), .Z(out[646]) );
  XOR U5769 ( .A(in[309]), .B(n3926), .Z(n4355) );
  XOR U5770 ( .A(in[1089]), .B(n3927), .Z(n4742) );
  XOR U5771 ( .A(in[1478]), .B(n3928), .Z(n4744) );
  OR U5772 ( .A(n4742), .B(n4744), .Z(n3929) );
  XOR U5773 ( .A(n4355), .B(n3929), .Z(out[647]) );
  XOR U5774 ( .A(in[310]), .B(n3930), .Z(n4357) );
  XOR U5775 ( .A(in[1479]), .B(n3931), .Z(n4748) );
  XNOR U5776 ( .A(n3932), .B(in[1090]), .Z(n4745) );
  NANDN U5777 ( .A(n4748), .B(n4745), .Z(n3933) );
  XOR U5778 ( .A(n4357), .B(n3933), .Z(out[648]) );
  XOR U5779 ( .A(in[311]), .B(n3934), .Z(n4360) );
  XNOR U5780 ( .A(n3936), .B(in[1091]), .Z(n4749) );
  NANDN U5781 ( .A(n4752), .B(n4749), .Z(n3937) );
  XOR U5782 ( .A(n4360), .B(n3937), .Z(out[649]) );
  XOR U5783 ( .A(in[312]), .B(n3941), .Z(n4363) );
  XNOR U5784 ( .A(n3943), .B(in[1092]), .Z(n4753) );
  NANDN U5785 ( .A(n4756), .B(n4753), .Z(n3944) );
  XOR U5786 ( .A(n4363), .B(n3944), .Z(out[650]) );
  XOR U5787 ( .A(in[313]), .B(n3945), .Z(n4366) );
  XNOR U5788 ( .A(n3947), .B(in[1093]), .Z(n4757) );
  NANDN U5789 ( .A(n4760), .B(n4757), .Z(n3948) );
  XOR U5790 ( .A(n4366), .B(n3948), .Z(out[651]) );
  XOR U5791 ( .A(in[314]), .B(n3949), .Z(n4373) );
  XNOR U5792 ( .A(n3951), .B(in[1094]), .Z(n4761) );
  NANDN U5793 ( .A(n4764), .B(n4761), .Z(n3952) );
  XOR U5794 ( .A(n4373), .B(n3952), .Z(out[652]) );
  XOR U5795 ( .A(in[315]), .B(n3953), .Z(n4206) );
  IV U5796 ( .A(n4206), .Z(n4376) );
  XNOR U5797 ( .A(n3955), .B(in[1095]), .Z(n4765) );
  NANDN U5798 ( .A(n4768), .B(n4765), .Z(n3956) );
  XOR U5799 ( .A(n4376), .B(n3956), .Z(out[653]) );
  XOR U5800 ( .A(in[316]), .B(n3957), .Z(n4209) );
  IV U5801 ( .A(n4209), .Z(n4379) );
  XNOR U5802 ( .A(n3959), .B(in[1096]), .Z(n4772) );
  NANDN U5803 ( .A(n4775), .B(n4772), .Z(n3960) );
  XOR U5804 ( .A(n4379), .B(n3960), .Z(out[654]) );
  XOR U5805 ( .A(in[317]), .B(n3961), .Z(n4212) );
  IV U5806 ( .A(n4212), .Z(n4382) );
  XNOR U5807 ( .A(in[1097]), .B(n3963), .Z(n4776) );
  NANDN U5808 ( .A(n4779), .B(n4776), .Z(n3964) );
  XOR U5809 ( .A(n4382), .B(n3964), .Z(out[655]) );
  XOR U5810 ( .A(in[318]), .B(n3965), .Z(n4217) );
  IV U5811 ( .A(n4217), .Z(n4385) );
  XNOR U5812 ( .A(n3967), .B(in[1098]), .Z(n4780) );
  NANDN U5813 ( .A(n4783), .B(n4780), .Z(n3968) );
  XOR U5814 ( .A(n4385), .B(n3968), .Z(out[656]) );
  XOR U5815 ( .A(in[319]), .B(n3969), .Z(n4220) );
  IV U5816 ( .A(n4220), .Z(n4387) );
  XNOR U5817 ( .A(n3971), .B(in[1099]), .Z(n4784) );
  NANDN U5818 ( .A(n4787), .B(n4784), .Z(n3972) );
  XOR U5819 ( .A(n4387), .B(n3972), .Z(out[657]) );
  XOR U5820 ( .A(in[256]), .B(n3973), .Z(n4223) );
  IV U5821 ( .A(n4223), .Z(n4390) );
  XNOR U5822 ( .A(in[1100]), .B(n3975), .Z(n4788) );
  NANDN U5823 ( .A(n4791), .B(n4788), .Z(n3976) );
  XOR U5824 ( .A(n4390), .B(n3976), .Z(out[658]) );
  XOR U5825 ( .A(in[257]), .B(n3977), .Z(n4226) );
  IV U5826 ( .A(n4226), .Z(n4393) );
  XNOR U5827 ( .A(in[1101]), .B(n3979), .Z(n4792) );
  NANDN U5828 ( .A(n4795), .B(n4792), .Z(n3980) );
  XOR U5829 ( .A(n4393), .B(n3980), .Z(out[659]) );
  XOR U5830 ( .A(in[258]), .B(n3984), .Z(n4229) );
  IV U5831 ( .A(n4229), .Z(n4396) );
  XOR U5832 ( .A(in[1491]), .B(n3985), .Z(n4799) );
  XNOR U5833 ( .A(in[1102]), .B(n3986), .Z(n4796) );
  NANDN U5834 ( .A(n4799), .B(n4796), .Z(n3987) );
  XOR U5835 ( .A(n4396), .B(n3987), .Z(out[660]) );
  XOR U5836 ( .A(in[259]), .B(n3988), .Z(n4232) );
  IV U5837 ( .A(n4232), .Z(n4399) );
  XOR U5838 ( .A(in[1492]), .B(n3989), .Z(n4803) );
  XNOR U5839 ( .A(in[1103]), .B(n3990), .Z(n4800) );
  NANDN U5840 ( .A(n4803), .B(n4800), .Z(n3991) );
  XOR U5841 ( .A(n4399), .B(n3991), .Z(out[661]) );
  XOR U5842 ( .A(in[260]), .B(n3992), .Z(n4406) );
  XOR U5843 ( .A(in[1493]), .B(n3993), .Z(n4235) );
  IV U5844 ( .A(n4235), .Z(n4807) );
  XNOR U5845 ( .A(in[1104]), .B(n3994), .Z(n4804) );
  NANDN U5846 ( .A(n4807), .B(n4804), .Z(n3995) );
  XNOR U5847 ( .A(n4406), .B(n3995), .Z(out[662]) );
  XOR U5848 ( .A(in[261]), .B(n3996), .Z(n4409) );
  XOR U5849 ( .A(in[1494]), .B(n3997), .Z(n4811) );
  XNOR U5850 ( .A(in[1105]), .B(n3998), .Z(n4808) );
  NANDN U5851 ( .A(n4811), .B(n4808), .Z(n3999) );
  XNOR U5852 ( .A(n4409), .B(n3999), .Z(out[663]) );
  XOR U5853 ( .A(in[262]), .B(n4000), .Z(n4412) );
  XOR U5854 ( .A(in[1495]), .B(n4001), .Z(n4818) );
  XOR U5855 ( .A(in[1106]), .B(n4002), .Z(n4815) );
  NANDN U5856 ( .A(n4818), .B(n4815), .Z(n4003) );
  XNOR U5857 ( .A(n4412), .B(n4003), .Z(out[664]) );
  XOR U5858 ( .A(in[263]), .B(n4004), .Z(n4415) );
  XOR U5859 ( .A(in[1496]), .B(n4005), .Z(n4240) );
  IV U5860 ( .A(n4240), .Z(n4822) );
  XNOR U5861 ( .A(in[1107]), .B(n4006), .Z(n4819) );
  NANDN U5862 ( .A(n4822), .B(n4819), .Z(n4007) );
  XNOR U5863 ( .A(n4415), .B(n4007), .Z(out[665]) );
  XOR U5864 ( .A(in[264]), .B(n4008), .Z(n4418) );
  XOR U5865 ( .A(in[1497]), .B(n4009), .Z(n4245) );
  IV U5866 ( .A(n4245), .Z(n4826) );
  XNOR U5867 ( .A(in[1108]), .B(n4010), .Z(n4823) );
  NANDN U5868 ( .A(n4826), .B(n4823), .Z(n4011) );
  XNOR U5869 ( .A(n4418), .B(n4011), .Z(out[666]) );
  XOR U5870 ( .A(in[265]), .B(n4012), .Z(n4421) );
  XOR U5871 ( .A(in[1498]), .B(n4013), .Z(n4830) );
  XNOR U5872 ( .A(in[1109]), .B(n4014), .Z(n4827) );
  NANDN U5873 ( .A(n4830), .B(n4827), .Z(n4015) );
  XNOR U5874 ( .A(n4421), .B(n4015), .Z(out[667]) );
  XOR U5875 ( .A(in[266]), .B(n4016), .Z(n4424) );
  XOR U5876 ( .A(in[1499]), .B(n4017), .Z(n4834) );
  XNOR U5877 ( .A(in[1110]), .B(n4018), .Z(n4831) );
  NANDN U5878 ( .A(n4834), .B(n4831), .Z(n4019) );
  XNOR U5879 ( .A(n4424), .B(n4019), .Z(out[668]) );
  XNOR U5880 ( .A(in[267]), .B(n4020), .Z(n4427) );
  XOR U5881 ( .A(in[1500]), .B(n4021), .Z(n4838) );
  XNOR U5882 ( .A(in[1111]), .B(n4022), .Z(n4835) );
  NANDN U5883 ( .A(n4838), .B(n4835), .Z(n4023) );
  XNOR U5884 ( .A(n4427), .B(n4023), .Z(out[669]) );
  ANDN U5885 ( .B(n4025), .A(n4024), .Z(n4026) );
  XOR U5886 ( .A(n4027), .B(n4026), .Z(out[66]) );
  XOR U5887 ( .A(in[268]), .B(n4028), .Z(n4430) );
  XOR U5888 ( .A(in[1501]), .B(n4029), .Z(n4842) );
  XNOR U5889 ( .A(in[1112]), .B(n4030), .Z(n4839) );
  NANDN U5890 ( .A(n4842), .B(n4839), .Z(n4031) );
  XNOR U5891 ( .A(n4430), .B(n4031), .Z(out[670]) );
  XNOR U5892 ( .A(in[269]), .B(n4032), .Z(n4433) );
  XOR U5893 ( .A(in[1502]), .B(n4033), .Z(n4846) );
  XNOR U5894 ( .A(in[1113]), .B(n4034), .Z(n4843) );
  NANDN U5895 ( .A(n4846), .B(n4843), .Z(n4035) );
  XNOR U5896 ( .A(n4433), .B(n4035), .Z(out[671]) );
  XOR U5897 ( .A(in[270]), .B(n4036), .Z(n4444) );
  XOR U5898 ( .A(in[1503]), .B(n4037), .Z(n4850) );
  XNOR U5899 ( .A(in[1114]), .B(n4038), .Z(n4847) );
  NANDN U5900 ( .A(n4850), .B(n4847), .Z(n4039) );
  XNOR U5901 ( .A(n4444), .B(n4039), .Z(out[672]) );
  XNOR U5902 ( .A(in[271]), .B(n4040), .Z(n4447) );
  XOR U5903 ( .A(in[1504]), .B(n4041), .Z(n4854) );
  XNOR U5904 ( .A(in[1115]), .B(n4042), .Z(n4851) );
  NANDN U5905 ( .A(n4854), .B(n4851), .Z(n4043) );
  XNOR U5906 ( .A(n4447), .B(n4043), .Z(out[673]) );
  XNOR U5907 ( .A(in[272]), .B(n4044), .Z(n4450) );
  XOR U5908 ( .A(in[1505]), .B(n4045), .Z(n4862) );
  XNOR U5909 ( .A(in[1116]), .B(n4046), .Z(n4859) );
  NANDN U5910 ( .A(n4862), .B(n4859), .Z(n4047) );
  XNOR U5911 ( .A(n4450), .B(n4047), .Z(out[674]) );
  XOR U5912 ( .A(in[273]), .B(n4048), .Z(n4453) );
  XOR U5913 ( .A(n4049), .B(in[1506]), .Z(n4866) );
  XNOR U5914 ( .A(in[1117]), .B(n4050), .Z(n4863) );
  NANDN U5915 ( .A(n4866), .B(n4863), .Z(n4051) );
  XNOR U5916 ( .A(n4453), .B(n4051), .Z(out[675]) );
  XOR U5917 ( .A(in[274]), .B(n4052), .Z(n4456) );
  XOR U5918 ( .A(n4053), .B(in[1507]), .Z(n4870) );
  XOR U5919 ( .A(in[1118]), .B(n4054), .Z(n4867) );
  NANDN U5920 ( .A(n4870), .B(n4867), .Z(n4055) );
  XNOR U5921 ( .A(n4456), .B(n4055), .Z(out[676]) );
  XOR U5922 ( .A(in[275]), .B(n4056), .Z(n4459) );
  XOR U5923 ( .A(n4057), .B(in[1508]), .Z(n4874) );
  XOR U5924 ( .A(in[1119]), .B(n4058), .Z(n4871) );
  NANDN U5925 ( .A(n4874), .B(n4871), .Z(n4059) );
  XNOR U5926 ( .A(n4459), .B(n4059), .Z(out[677]) );
  XOR U5927 ( .A(in[276]), .B(n4060), .Z(n4462) );
  XOR U5928 ( .A(n4061), .B(in[1509]), .Z(n4878) );
  XOR U5929 ( .A(in[1120]), .B(n4062), .Z(n4875) );
  NANDN U5930 ( .A(n4878), .B(n4875), .Z(n4063) );
  XNOR U5931 ( .A(n4462), .B(n4063), .Z(out[678]) );
  XOR U5932 ( .A(in[277]), .B(n4064), .Z(n4465) );
  XOR U5933 ( .A(in[1510]), .B(n4065), .Z(n4262) );
  IV U5934 ( .A(n4262), .Z(n4882) );
  XOR U5935 ( .A(in[1121]), .B(n4066), .Z(n4879) );
  NANDN U5936 ( .A(n4882), .B(n4879), .Z(n4067) );
  XNOR U5937 ( .A(n4465), .B(n4067), .Z(out[679]) );
  ANDN U5938 ( .B(n4069), .A(n4068), .Z(n4070) );
  XOR U5939 ( .A(n4071), .B(n4070), .Z(out[67]) );
  XOR U5940 ( .A(in[278]), .B(n4072), .Z(n4468) );
  XOR U5941 ( .A(in[1511]), .B(n4073), .Z(n4265) );
  IV U5942 ( .A(n4265), .Z(n4886) );
  XOR U5943 ( .A(in[1122]), .B(n4074), .Z(n4883) );
  NANDN U5944 ( .A(n4886), .B(n4883), .Z(n4075) );
  XNOR U5945 ( .A(n4468), .B(n4075), .Z(out[680]) );
  XOR U5946 ( .A(in[279]), .B(n4076), .Z(n4471) );
  XOR U5947 ( .A(in[1512]), .B(n4077), .Z(n4268) );
  IV U5948 ( .A(n4268), .Z(n4890) );
  XOR U5949 ( .A(in[1123]), .B(n4078), .Z(n4887) );
  NANDN U5950 ( .A(n4890), .B(n4887), .Z(n4079) );
  XNOR U5951 ( .A(n4471), .B(n4079), .Z(out[681]) );
  XOR U5952 ( .A(in[280]), .B(n4080), .Z(n4478) );
  XOR U5953 ( .A(in[1513]), .B(n4081), .Z(n4271) );
  IV U5954 ( .A(n4271), .Z(n4894) );
  XOR U5955 ( .A(in[1124]), .B(n4082), .Z(n4891) );
  NANDN U5956 ( .A(n4894), .B(n4891), .Z(n4083) );
  XNOR U5957 ( .A(n4478), .B(n4083), .Z(out[682]) );
  XOR U5958 ( .A(in[281]), .B(n4084), .Z(n4481) );
  XOR U5959 ( .A(in[1514]), .B(n4085), .Z(n4274) );
  IV U5960 ( .A(n4274), .Z(n4898) );
  XNOR U5961 ( .A(in[1125]), .B(n4086), .Z(n4895) );
  NANDN U5962 ( .A(n4898), .B(n4895), .Z(n4087) );
  XNOR U5963 ( .A(n4481), .B(n4087), .Z(out[683]) );
  XOR U5964 ( .A(in[282]), .B(n4088), .Z(n4484) );
  XOR U5965 ( .A(in[1126]), .B(n4089), .Z(n4904) );
  XNOR U5966 ( .A(in[1515]), .B(n4090), .Z(n4906) );
  NANDN U5967 ( .A(n4904), .B(n4906), .Z(n4091) );
  XNOR U5968 ( .A(n4484), .B(n4091), .Z(out[684]) );
  XOR U5969 ( .A(in[283]), .B(n4092), .Z(n4487) );
  XOR U5970 ( .A(in[1127]), .B(n4093), .Z(n4908) );
  XNOR U5971 ( .A(in[1516]), .B(n4094), .Z(n4910) );
  NANDN U5972 ( .A(n4908), .B(n4910), .Z(n4095) );
  XNOR U5973 ( .A(n4487), .B(n4095), .Z(out[685]) );
  XOR U5974 ( .A(in[284]), .B(n4096), .Z(n4490) );
  XOR U5975 ( .A(in[1128]), .B(n4097), .Z(n4912) );
  XNOR U5976 ( .A(in[1517]), .B(n4098), .Z(n4914) );
  NANDN U5977 ( .A(n4912), .B(n4914), .Z(n4099) );
  XNOR U5978 ( .A(n4490), .B(n4099), .Z(out[686]) );
  XOR U5979 ( .A(in[285]), .B(n4100), .Z(n4493) );
  XOR U5980 ( .A(in[1129]), .B(n4101), .Z(n4916) );
  XNOR U5981 ( .A(in[1518]), .B(n4102), .Z(n4918) );
  NANDN U5982 ( .A(n4916), .B(n4918), .Z(n4103) );
  XNOR U5983 ( .A(n4493), .B(n4103), .Z(out[687]) );
  XOR U5984 ( .A(in[286]), .B(n4104), .Z(n4496) );
  XOR U5985 ( .A(in[1130]), .B(n4105), .Z(n4920) );
  XNOR U5986 ( .A(in[1519]), .B(n4106), .Z(n4922) );
  NANDN U5987 ( .A(n4920), .B(n4922), .Z(n4107) );
  XNOR U5988 ( .A(n4496), .B(n4107), .Z(out[688]) );
  XOR U5989 ( .A(in[287]), .B(n4108), .Z(n4499) );
  XNOR U5990 ( .A(in[1131]), .B(n4109), .Z(n4924) );
  XNOR U5991 ( .A(in[1520]), .B(n4110), .Z(n4926) );
  NANDN U5992 ( .A(n4924), .B(n4926), .Z(n4111) );
  XNOR U5993 ( .A(n4499), .B(n4111), .Z(out[689]) );
  ANDN U5994 ( .B(n4113), .A(n4112), .Z(n4114) );
  XOR U5995 ( .A(n4115), .B(n4114), .Z(out[68]) );
  XOR U5996 ( .A(in[288]), .B(n4116), .Z(n4502) );
  XNOR U5997 ( .A(in[1132]), .B(n4117), .Z(n4928) );
  XNOR U5998 ( .A(in[1521]), .B(n4118), .Z(n4930) );
  NANDN U5999 ( .A(n4928), .B(n4930), .Z(n4119) );
  XNOR U6000 ( .A(n4502), .B(n4119), .Z(out[690]) );
  XOR U6001 ( .A(in[289]), .B(n4120), .Z(n4505) );
  XOR U6002 ( .A(in[1133]), .B(n4121), .Z(n4932) );
  XNOR U6003 ( .A(in[1522]), .B(n4122), .Z(n4934) );
  NANDN U6004 ( .A(n4932), .B(n4934), .Z(n4123) );
  XNOR U6005 ( .A(n4505), .B(n4123), .Z(out[691]) );
  XOR U6006 ( .A(in[290]), .B(n4124), .Z(n4512) );
  XOR U6007 ( .A(in[1134]), .B(n4125), .Z(n4936) );
  XNOR U6008 ( .A(in[1523]), .B(n4126), .Z(n4938) );
  NANDN U6009 ( .A(n4936), .B(n4938), .Z(n4127) );
  XNOR U6010 ( .A(n4512), .B(n4127), .Z(out[692]) );
  XOR U6011 ( .A(in[291]), .B(n4128), .Z(n4515) );
  XOR U6012 ( .A(in[1135]), .B(n4129), .Z(n4940) );
  XNOR U6013 ( .A(in[1524]), .B(n4130), .Z(n4942) );
  NANDN U6014 ( .A(n4940), .B(n4942), .Z(n4131) );
  XNOR U6015 ( .A(n4515), .B(n4131), .Z(out[693]) );
  XOR U6016 ( .A(in[292]), .B(n4132), .Z(n4518) );
  XOR U6017 ( .A(in[1136]), .B(n4133), .Z(n4948) );
  XNOR U6018 ( .A(in[1525]), .B(n4134), .Z(n4950) );
  NANDN U6019 ( .A(n4948), .B(n4950), .Z(n4135) );
  XNOR U6020 ( .A(n4518), .B(n4135), .Z(out[694]) );
  XOR U6021 ( .A(in[293]), .B(n4136), .Z(n4303) );
  IV U6022 ( .A(n4303), .Z(n4522) );
  XOR U6023 ( .A(in[1137]), .B(n4137), .Z(n4952) );
  XNOR U6024 ( .A(in[1526]), .B(n4138), .Z(n4954) );
  NANDN U6025 ( .A(n4952), .B(n4954), .Z(n4139) );
  XOR U6026 ( .A(n4522), .B(n4139), .Z(out[695]) );
  XOR U6027 ( .A(in[294]), .B(n4140), .Z(n4310) );
  IV U6028 ( .A(n4310), .Z(n4526) );
  XOR U6029 ( .A(in[1138]), .B(n4141), .Z(n4956) );
  XNOR U6030 ( .A(in[1527]), .B(n4142), .Z(n4958) );
  NANDN U6031 ( .A(n4956), .B(n4958), .Z(n4143) );
  XOR U6032 ( .A(n4526), .B(n4143), .Z(out[696]) );
  XOR U6033 ( .A(in[295]), .B(n4144), .Z(n4313) );
  IV U6034 ( .A(n4313), .Z(n4530) );
  XOR U6035 ( .A(in[1139]), .B(n4145), .Z(n4960) );
  XNOR U6036 ( .A(in[1528]), .B(n4146), .Z(n4962) );
  NANDN U6037 ( .A(n4960), .B(n4962), .Z(n4147) );
  XOR U6038 ( .A(n4530), .B(n4147), .Z(out[697]) );
  XOR U6039 ( .A(in[296]), .B(n4148), .Z(n4316) );
  IV U6040 ( .A(n4316), .Z(n4534) );
  XOR U6041 ( .A(in[1140]), .B(n4149), .Z(n4964) );
  XNOR U6042 ( .A(in[1529]), .B(n4150), .Z(n4966) );
  NANDN U6043 ( .A(n4964), .B(n4966), .Z(n4151) );
  XOR U6044 ( .A(n4534), .B(n4151), .Z(out[698]) );
  XOR U6045 ( .A(in[297]), .B(n4152), .Z(n4319) );
  IV U6046 ( .A(n4319), .Z(n4538) );
  XNOR U6047 ( .A(in[1141]), .B(n4153), .Z(n4968) );
  XNOR U6048 ( .A(in[1530]), .B(n4154), .Z(n4970) );
  NANDN U6049 ( .A(n4968), .B(n4970), .Z(n4155) );
  XOR U6050 ( .A(n4538), .B(n4155), .Z(out[699]) );
  ANDN U6051 ( .B(n4157), .A(n4156), .Z(n4158) );
  XOR U6052 ( .A(n4159), .B(n4158), .Z(out[69]) );
  OR U6053 ( .A(n4195), .B(n4160), .Z(n4161) );
  XNOR U6054 ( .A(n4194), .B(n4161), .Z(out[6]) );
  XOR U6055 ( .A(in[298]), .B(n4162), .Z(n4322) );
  IV U6056 ( .A(n4322), .Z(n4542) );
  XNOR U6057 ( .A(in[1142]), .B(n4163), .Z(n4972) );
  XNOR U6058 ( .A(in[1531]), .B(n4164), .Z(n4974) );
  OR U6059 ( .A(n4972), .B(n4974), .Z(n4165) );
  XOR U6060 ( .A(n4542), .B(n4165), .Z(out[700]) );
  XOR U6061 ( .A(in[299]), .B(n4166), .Z(n4325) );
  IV U6062 ( .A(n4325), .Z(n4545) );
  XNOR U6063 ( .A(in[1143]), .B(n4167), .Z(n4976) );
  XNOR U6064 ( .A(in[1532]), .B(n4168), .Z(n4978) );
  OR U6065 ( .A(n4976), .B(n4978), .Z(n4169) );
  XOR U6066 ( .A(n4545), .B(n4169), .Z(out[701]) );
  XOR U6067 ( .A(in[300]), .B(n4170), .Z(n4328) );
  IV U6068 ( .A(n4328), .Z(n4551) );
  XNOR U6069 ( .A(in[1144]), .B(n4171), .Z(n4980) );
  XNOR U6070 ( .A(in[1533]), .B(n4172), .Z(n4982) );
  OR U6071 ( .A(n4980), .B(n4982), .Z(n4173) );
  XOR U6072 ( .A(n4551), .B(n4173), .Z(out[702]) );
  XOR U6073 ( .A(in[301]), .B(n4174), .Z(n4331) );
  IV U6074 ( .A(n4331), .Z(n4553) );
  XNOR U6075 ( .A(in[1145]), .B(n4175), .Z(n4984) );
  XNOR U6076 ( .A(in[1534]), .B(n4176), .Z(n4986) );
  NANDN U6077 ( .A(n4984), .B(n4986), .Z(n4177) );
  XOR U6078 ( .A(n4553), .B(n4177), .Z(out[703]) );
  XOR U6079 ( .A(in[376]), .B(n4178), .Z(n4554) );
  ANDN U6080 ( .B(n4708), .A(n4179), .Z(n4180) );
  XOR U6081 ( .A(n4554), .B(n4180), .Z(out[704]) );
  XOR U6082 ( .A(in[377]), .B(n4181), .Z(n4557) );
  ANDN U6083 ( .B(n4712), .A(n4182), .Z(n4183) );
  XOR U6084 ( .A(n4557), .B(n4183), .Z(out[705]) );
  XOR U6085 ( .A(in[378]), .B(n4184), .Z(n4560) );
  ANDN U6086 ( .B(n4716), .A(n4185), .Z(n4186) );
  XOR U6087 ( .A(n4560), .B(n4186), .Z(out[706]) );
  XOR U6088 ( .A(in[379]), .B(n4187), .Z(n4563) );
  ANDN U6089 ( .B(n4720), .A(n4188), .Z(n4189) );
  XOR U6090 ( .A(n4563), .B(n4189), .Z(out[707]) );
  XOR U6091 ( .A(in[380]), .B(n4190), .Z(n4566) );
  ANDN U6092 ( .B(n4732), .A(n4191), .Z(n4192) );
  XNOR U6093 ( .A(n4566), .B(n4192), .Z(out[708]) );
  XOR U6094 ( .A(in[381]), .B(n4193), .Z(n4568) );
  ANDN U6095 ( .B(n4195), .A(n4194), .Z(n4196) );
  XOR U6096 ( .A(n4197), .B(n4196), .Z(out[70]) );
  XOR U6097 ( .A(in[382]), .B(n4198), .Z(n4570) );
  XOR U6098 ( .A(in[383]), .B(n4199), .Z(n4572) );
  XOR U6099 ( .A(in[320]), .B(n4200), .Z(n4579) );
  XOR U6100 ( .A(in[321]), .B(n4201), .Z(n4581) );
  XOR U6101 ( .A(in[322]), .B(n4202), .Z(n4583) );
  XOR U6102 ( .A(in[323]), .B(n4203), .Z(n4585) );
  XOR U6103 ( .A(in[324]), .B(n4204), .Z(n4587) );
  XOR U6104 ( .A(in[325]), .B(n4205), .Z(n4589) );
  ANDN U6105 ( .B(n4768), .A(n4206), .Z(n4207) );
  XNOR U6106 ( .A(n4589), .B(n4207), .Z(out[717]) );
  XOR U6107 ( .A(in[326]), .B(n4208), .Z(n4591) );
  ANDN U6108 ( .B(n4775), .A(n4209), .Z(n4210) );
  XNOR U6109 ( .A(n4591), .B(n4210), .Z(out[718]) );
  XOR U6110 ( .A(in[327]), .B(n4211), .Z(n4593) );
  ANDN U6111 ( .B(n4779), .A(n4212), .Z(n4213) );
  XNOR U6112 ( .A(n4593), .B(n4213), .Z(out[719]) );
  ANDN U6113 ( .B(n4440), .A(n4442), .Z(n4214) );
  XOR U6114 ( .A(n4215), .B(n4214), .Z(out[71]) );
  XOR U6115 ( .A(in[328]), .B(n4216), .Z(n4595) );
  ANDN U6116 ( .B(n4783), .A(n4217), .Z(n4218) );
  XOR U6117 ( .A(n4595), .B(n4218), .Z(out[720]) );
  XOR U6118 ( .A(in[329]), .B(n4219), .Z(n4598) );
  ANDN U6119 ( .B(n4787), .A(n4220), .Z(n4221) );
  XNOR U6120 ( .A(n4598), .B(n4221), .Z(out[721]) );
  XOR U6121 ( .A(in[330]), .B(n4222), .Z(n4604) );
  ANDN U6122 ( .B(n4791), .A(n4223), .Z(n4224) );
  XNOR U6123 ( .A(n4604), .B(n4224), .Z(out[722]) );
  XOR U6124 ( .A(in[331]), .B(n4225), .Z(n4606) );
  ANDN U6125 ( .B(n4795), .A(n4226), .Z(n4227) );
  XNOR U6126 ( .A(n4606), .B(n4227), .Z(out[723]) );
  XOR U6127 ( .A(in[332]), .B(n4228), .Z(n4608) );
  ANDN U6128 ( .B(n4799), .A(n4229), .Z(n4230) );
  XNOR U6129 ( .A(n4608), .B(n4230), .Z(out[724]) );
  XOR U6130 ( .A(in[333]), .B(n4231), .Z(n4610) );
  ANDN U6131 ( .B(n4803), .A(n4232), .Z(n4233) );
  XNOR U6132 ( .A(n4610), .B(n4233), .Z(out[725]) );
  XOR U6133 ( .A(in[334]), .B(n4234), .Z(n4612) );
  NOR U6134 ( .A(n4235), .B(n4406), .Z(n4236) );
  XNOR U6135 ( .A(n4612), .B(n4236), .Z(out[726]) );
  XOR U6136 ( .A(in[335]), .B(n4237), .Z(n4614) );
  XOR U6137 ( .A(in[336]), .B(n4238), .Z(n4617) );
  XOR U6138 ( .A(in[337]), .B(n4239), .Z(n4619) );
  NOR U6139 ( .A(n4240), .B(n4415), .Z(n4241) );
  XNOR U6140 ( .A(n4619), .B(n4241), .Z(out[729]) );
  ANDN U6141 ( .B(n4726), .A(n4728), .Z(n4242) );
  XOR U6142 ( .A(n4243), .B(n4242), .Z(out[72]) );
  XOR U6143 ( .A(in[338]), .B(n4244), .Z(n4621) );
  NOR U6144 ( .A(n4245), .B(n4418), .Z(n4246) );
  XNOR U6145 ( .A(n4621), .B(n4246), .Z(out[730]) );
  XOR U6146 ( .A(in[339]), .B(n4247), .Z(n4623) );
  XOR U6147 ( .A(in[340]), .B(n4248), .Z(n4629) );
  XOR U6148 ( .A(in[341]), .B(n4249), .Z(n4632) );
  XOR U6149 ( .A(in[342]), .B(n4250), .Z(n4635) );
  XOR U6150 ( .A(in[343]), .B(n4251), .Z(n4638) );
  XOR U6151 ( .A(in[344]), .B(n4252), .Z(n4639) );
  XOR U6152 ( .A(in[345]), .B(n4253), .Z(n4642) );
  XOR U6153 ( .A(in[346]), .B(n4254), .Z(n4645) );
  XOR U6154 ( .A(in[347]), .B(n4255), .Z(n4648) );
  ANDN U6155 ( .B(n5154), .A(n5156), .Z(n4256) );
  XOR U6156 ( .A(n4257), .B(n4256), .Z(out[73]) );
  XOR U6157 ( .A(in[348]), .B(n4258), .Z(n4651) );
  XOR U6158 ( .A(in[349]), .B(n4259), .Z(n4654) );
  XOR U6159 ( .A(in[350]), .B(n4260), .Z(n4659) );
  XOR U6160 ( .A(in[351]), .B(n4261), .Z(n4660) );
  NOR U6161 ( .A(n4262), .B(n4465), .Z(n4263) );
  XOR U6162 ( .A(n4660), .B(n4263), .Z(out[743]) );
  XOR U6163 ( .A(in[352]), .B(n4264), .Z(n4661) );
  NOR U6164 ( .A(n4265), .B(n4468), .Z(n4266) );
  XOR U6165 ( .A(n4661), .B(n4266), .Z(out[744]) );
  XOR U6166 ( .A(in[353]), .B(n4267), .Z(n4662) );
  NOR U6167 ( .A(n4268), .B(n4471), .Z(n4269) );
  XOR U6168 ( .A(n4662), .B(n4269), .Z(out[745]) );
  XOR U6169 ( .A(in[354]), .B(n4270), .Z(n4663) );
  NOR U6170 ( .A(n4271), .B(n4478), .Z(n4272) );
  XOR U6171 ( .A(n4663), .B(n4272), .Z(out[746]) );
  XOR U6172 ( .A(in[355]), .B(n4273), .Z(n4664) );
  NOR U6173 ( .A(n4274), .B(n4481), .Z(n4275) );
  XNOR U6174 ( .A(n4664), .B(n4275), .Z(out[747]) );
  XOR U6175 ( .A(in[356]), .B(n4276), .Z(n4666) );
  NOR U6176 ( .A(n4906), .B(n4484), .Z(n4277) );
  XOR U6177 ( .A(n4666), .B(n4277), .Z(out[748]) );
  XOR U6178 ( .A(in[357]), .B(n4278), .Z(n4667) );
  NOR U6179 ( .A(n4910), .B(n4487), .Z(n4279) );
  XOR U6180 ( .A(n4667), .B(n4279), .Z(out[749]) );
  ANDN U6181 ( .B(n4281), .A(n4280), .Z(n4282) );
  XOR U6182 ( .A(n4283), .B(n4282), .Z(out[74]) );
  XOR U6183 ( .A(in[358]), .B(n4284), .Z(n4668) );
  NOR U6184 ( .A(n4914), .B(n4490), .Z(n4285) );
  XOR U6185 ( .A(n4668), .B(n4285), .Z(out[750]) );
  XOR U6186 ( .A(in[359]), .B(n4286), .Z(n4669) );
  NOR U6187 ( .A(n4918), .B(n4493), .Z(n4287) );
  XOR U6188 ( .A(n4669), .B(n4287), .Z(out[751]) );
  XOR U6189 ( .A(in[360]), .B(n4288), .Z(n4673) );
  NOR U6190 ( .A(n4922), .B(n4496), .Z(n4289) );
  XOR U6191 ( .A(n4673), .B(n4289), .Z(out[752]) );
  XOR U6192 ( .A(in[361]), .B(n4290), .Z(n4674) );
  NOR U6193 ( .A(n4926), .B(n4499), .Z(n4291) );
  XOR U6194 ( .A(n4674), .B(n4291), .Z(out[753]) );
  XOR U6195 ( .A(in[362]), .B(n4292), .Z(n4675) );
  NOR U6196 ( .A(n4930), .B(n4502), .Z(n4293) );
  XOR U6197 ( .A(n4675), .B(n4293), .Z(out[754]) );
  XOR U6198 ( .A(in[363]), .B(n4294), .Z(n4676) );
  NOR U6199 ( .A(n4934), .B(n4505), .Z(n4295) );
  XOR U6200 ( .A(n4676), .B(n4295), .Z(out[755]) );
  XOR U6201 ( .A(in[364]), .B(n4296), .Z(n4677) );
  NOR U6202 ( .A(n4938), .B(n4512), .Z(n4297) );
  XOR U6203 ( .A(n4677), .B(n4297), .Z(out[756]) );
  XOR U6204 ( .A(in[365]), .B(n4298), .Z(n4678) );
  NOR U6205 ( .A(n4942), .B(n4515), .Z(n4299) );
  XOR U6206 ( .A(n4678), .B(n4299), .Z(out[757]) );
  XOR U6207 ( .A(in[366]), .B(n4300), .Z(n4679) );
  NOR U6208 ( .A(n4950), .B(n4518), .Z(n4301) );
  XOR U6209 ( .A(n4679), .B(n4301), .Z(out[758]) );
  XOR U6210 ( .A(in[367]), .B(n4302), .Z(n4521) );
  NOR U6211 ( .A(n4303), .B(n4954), .Z(n4304) );
  XOR U6212 ( .A(n4521), .B(n4304), .Z(out[759]) );
  ANDN U6213 ( .B(n4306), .A(n4305), .Z(n4307) );
  XOR U6214 ( .A(n4308), .B(n4307), .Z(out[75]) );
  XOR U6215 ( .A(in[368]), .B(n4309), .Z(n4525) );
  NOR U6216 ( .A(n4310), .B(n4958), .Z(n4311) );
  XOR U6217 ( .A(n4525), .B(n4311), .Z(out[760]) );
  XOR U6218 ( .A(in[369]), .B(n4312), .Z(n4529) );
  NOR U6219 ( .A(n4313), .B(n4962), .Z(n4314) );
  XOR U6220 ( .A(n4529), .B(n4314), .Z(out[761]) );
  XOR U6221 ( .A(in[370]), .B(n4315), .Z(n4533) );
  NOR U6222 ( .A(n4316), .B(n4966), .Z(n4317) );
  XOR U6223 ( .A(n4533), .B(n4317), .Z(out[762]) );
  XOR U6224 ( .A(in[371]), .B(n4318), .Z(n4537) );
  NOR U6225 ( .A(n4319), .B(n4970), .Z(n4320) );
  XOR U6226 ( .A(n4537), .B(n4320), .Z(out[763]) );
  XOR U6227 ( .A(in[372]), .B(n4321), .Z(n4541) );
  ANDN U6228 ( .B(n4974), .A(n4322), .Z(n4323) );
  XOR U6229 ( .A(n4541), .B(n4323), .Z(out[764]) );
  XOR U6230 ( .A(in[373]), .B(n4324), .Z(n4696) );
  ANDN U6231 ( .B(n4978), .A(n4325), .Z(n4326) );
  XOR U6232 ( .A(n4696), .B(n4326), .Z(out[765]) );
  XOR U6233 ( .A(in[374]), .B(n4327), .Z(n4699) );
  ANDN U6234 ( .B(n4982), .A(n4328), .Z(n4329) );
  XOR U6235 ( .A(n4699), .B(n4329), .Z(out[766]) );
  XOR U6236 ( .A(in[375]), .B(n4330), .Z(n4702) );
  NOR U6237 ( .A(n4331), .B(n4986), .Z(n4332) );
  XOR U6238 ( .A(n4702), .B(n4332), .Z(out[767]) );
  XOR U6239 ( .A(in[743]), .B(n4333), .Z(n4555) );
  IV U6240 ( .A(n4555), .Z(n4705) );
  XOR U6241 ( .A(in[744]), .B(n4335), .Z(n4558) );
  IV U6242 ( .A(n4558), .Z(n4709) );
  ANDN U6243 ( .B(n4338), .A(n4337), .Z(n4339) );
  XOR U6244 ( .A(n4340), .B(n4339), .Z(out[76]) );
  XOR U6245 ( .A(in[745]), .B(n4341), .Z(n4561) );
  IV U6246 ( .A(n4561), .Z(n4713) );
  XOR U6247 ( .A(in[746]), .B(n4343), .Z(n4564) );
  IV U6248 ( .A(n4564), .Z(n4717) );
  XNOR U6249 ( .A(in[747]), .B(n4345), .Z(n4729) );
  NANDN U6250 ( .A(n4346), .B(n4566), .Z(n4347) );
  XOR U6251 ( .A(n4729), .B(n4347), .Z(out[772]) );
  XNOR U6252 ( .A(in[748]), .B(n4348), .Z(n4733) );
  NANDN U6253 ( .A(n4349), .B(n4568), .Z(n4350) );
  XOR U6254 ( .A(n4733), .B(n4350), .Z(out[773]) );
  XNOR U6255 ( .A(in[749]), .B(n4351), .Z(n4737) );
  NANDN U6256 ( .A(n4352), .B(n4570), .Z(n4353) );
  XOR U6257 ( .A(n4737), .B(n4353), .Z(out[774]) );
  XOR U6258 ( .A(in[750]), .B(n4354), .Z(n4573) );
  IV U6259 ( .A(n4573), .Z(n4741) );
  XNOR U6260 ( .A(in[751]), .B(n4356), .Z(n4746) );
  NANDN U6261 ( .A(n4357), .B(n4579), .Z(n4358) );
  XOR U6262 ( .A(n4746), .B(n4358), .Z(out[776]) );
  XNOR U6263 ( .A(in[752]), .B(n4359), .Z(n4750) );
  NANDN U6264 ( .A(n4360), .B(n4581), .Z(n4361) );
  XOR U6265 ( .A(n4750), .B(n4361), .Z(out[777]) );
  XNOR U6266 ( .A(in[753]), .B(n4362), .Z(n4754) );
  NANDN U6267 ( .A(n4363), .B(n4583), .Z(n4364) );
  XOR U6268 ( .A(n4754), .B(n4364), .Z(out[778]) );
  XNOR U6269 ( .A(in[754]), .B(n4365), .Z(n4758) );
  NANDN U6270 ( .A(n4366), .B(n4585), .Z(n4367) );
  XOR U6271 ( .A(n4758), .B(n4367), .Z(out[779]) );
  ANDN U6272 ( .B(n4369), .A(n4368), .Z(n4370) );
  XOR U6273 ( .A(n4371), .B(n4370), .Z(out[77]) );
  XNOR U6274 ( .A(in[755]), .B(n4372), .Z(n4762) );
  NANDN U6275 ( .A(n4373), .B(n4587), .Z(n4374) );
  XOR U6276 ( .A(n4762), .B(n4374), .Z(out[780]) );
  XNOR U6277 ( .A(in[756]), .B(n4375), .Z(n4766) );
  NANDN U6278 ( .A(n4376), .B(n4589), .Z(n4377) );
  XOR U6279 ( .A(n4766), .B(n4377), .Z(out[781]) );
  XNOR U6280 ( .A(in[757]), .B(n4378), .Z(n4773) );
  NANDN U6281 ( .A(n4379), .B(n4591), .Z(n4380) );
  XOR U6282 ( .A(n4773), .B(n4380), .Z(out[782]) );
  XNOR U6283 ( .A(in[758]), .B(n4381), .Z(n4777) );
  NANDN U6284 ( .A(n4382), .B(n4593), .Z(n4383) );
  XOR U6285 ( .A(n4777), .B(n4383), .Z(out[783]) );
  XOR U6286 ( .A(in[759]), .B(n4384), .Z(n4596) );
  IV U6287 ( .A(n4596), .Z(n4781) );
  XNOR U6288 ( .A(in[760]), .B(n4386), .Z(n4785) );
  NANDN U6289 ( .A(n4387), .B(n4598), .Z(n4388) );
  XOR U6290 ( .A(n4785), .B(n4388), .Z(out[785]) );
  XNOR U6291 ( .A(in[761]), .B(n4389), .Z(n4789) );
  NANDN U6292 ( .A(n4390), .B(n4604), .Z(n4391) );
  XOR U6293 ( .A(n4789), .B(n4391), .Z(out[786]) );
  XOR U6294 ( .A(in[762]), .B(n4392), .Z(n4793) );
  NANDN U6295 ( .A(n4393), .B(n4606), .Z(n4394) );
  XOR U6296 ( .A(n4793), .B(n4394), .Z(out[787]) );
  XOR U6297 ( .A(in[763]), .B(n4395), .Z(n4797) );
  NANDN U6298 ( .A(n4396), .B(n4608), .Z(n4397) );
  XOR U6299 ( .A(n4797), .B(n4397), .Z(out[788]) );
  XNOR U6300 ( .A(in[764]), .B(n4398), .Z(n4801) );
  NANDN U6301 ( .A(n4399), .B(n4610), .Z(n4400) );
  XOR U6302 ( .A(n4801), .B(n4400), .Z(out[789]) );
  ANDN U6303 ( .B(n4402), .A(n4401), .Z(n4403) );
  XOR U6304 ( .A(n4404), .B(n4403), .Z(out[78]) );
  XNOR U6305 ( .A(in[765]), .B(n4405), .Z(n4805) );
  NAND U6306 ( .A(n4406), .B(n4612), .Z(n4407) );
  XOR U6307 ( .A(n4805), .B(n4407), .Z(out[790]) );
  XOR U6308 ( .A(in[766]), .B(n4408), .Z(n4615) );
  IV U6309 ( .A(n4615), .Z(n4809) );
  NANDN U6310 ( .A(n4614), .B(n4409), .Z(n4410) );
  XOR U6311 ( .A(n4809), .B(n4410), .Z(out[791]) );
  XNOR U6312 ( .A(in[767]), .B(n4411), .Z(n4816) );
  NAND U6313 ( .A(n4412), .B(n4617), .Z(n4413) );
  XOR U6314 ( .A(n4816), .B(n4413), .Z(out[792]) );
  XNOR U6315 ( .A(in[704]), .B(n4414), .Z(n4820) );
  NAND U6316 ( .A(n4415), .B(n4619), .Z(n4416) );
  XOR U6317 ( .A(n4820), .B(n4416), .Z(out[793]) );
  XNOR U6318 ( .A(in[705]), .B(n4417), .Z(n4824) );
  NAND U6319 ( .A(n4418), .B(n4621), .Z(n4419) );
  XOR U6320 ( .A(n4824), .B(n4419), .Z(out[794]) );
  XNOR U6321 ( .A(in[706]), .B(n4420), .Z(n4828) );
  NAND U6322 ( .A(n4421), .B(n4623), .Z(n4422) );
  XOR U6323 ( .A(n4828), .B(n4422), .Z(out[795]) );
  XOR U6324 ( .A(in[707]), .B(n4423), .Z(n4630) );
  IV U6325 ( .A(n4630), .Z(n4832) );
  NANDN U6326 ( .A(n4629), .B(n4424), .Z(n4425) );
  XOR U6327 ( .A(n4832), .B(n4425), .Z(out[796]) );
  XOR U6328 ( .A(in[708]), .B(n4426), .Z(n4633) );
  IV U6329 ( .A(n4633), .Z(n4836) );
  NANDN U6330 ( .A(n4632), .B(n4427), .Z(n4428) );
  XOR U6331 ( .A(n4836), .B(n4428), .Z(out[797]) );
  XOR U6332 ( .A(in[709]), .B(n4429), .Z(n4636) );
  IV U6333 ( .A(n4636), .Z(n4840) );
  NANDN U6334 ( .A(n4635), .B(n4430), .Z(n4431) );
  XOR U6335 ( .A(n4840), .B(n4431), .Z(out[798]) );
  XOR U6336 ( .A(in[710]), .B(n4432), .Z(n4844) );
  NANDN U6337 ( .A(n4638), .B(n4433), .Z(n4434) );
  XOR U6338 ( .A(n4844), .B(n4434), .Z(out[799]) );
  ANDN U6339 ( .B(n4436), .A(n4435), .Z(n4437) );
  XOR U6340 ( .A(n4438), .B(n4437), .Z(out[79]) );
  OR U6341 ( .A(n4440), .B(n4439), .Z(n4441) );
  XNOR U6342 ( .A(n4442), .B(n4441), .Z(out[7]) );
  XOR U6343 ( .A(in[711]), .B(n4443), .Z(n4640) );
  IV U6344 ( .A(n4640), .Z(n4848) );
  NANDN U6345 ( .A(n4639), .B(n4444), .Z(n4445) );
  XOR U6346 ( .A(n4848), .B(n4445), .Z(out[800]) );
  XOR U6347 ( .A(in[712]), .B(n4446), .Z(n4643) );
  IV U6348 ( .A(n4643), .Z(n4852) );
  NANDN U6349 ( .A(n4642), .B(n4447), .Z(n4448) );
  XOR U6350 ( .A(n4852), .B(n4448), .Z(out[801]) );
  XOR U6351 ( .A(in[713]), .B(n4449), .Z(n4646) );
  IV U6352 ( .A(n4646), .Z(n4860) );
  NANDN U6353 ( .A(n4645), .B(n4450), .Z(n4451) );
  XOR U6354 ( .A(n4860), .B(n4451), .Z(out[802]) );
  XOR U6355 ( .A(in[714]), .B(n4452), .Z(n4649) );
  IV U6356 ( .A(n4649), .Z(n4864) );
  NANDN U6357 ( .A(n4648), .B(n4453), .Z(n4454) );
  XOR U6358 ( .A(n4864), .B(n4454), .Z(out[803]) );
  XOR U6359 ( .A(in[715]), .B(n4455), .Z(n4652) );
  IV U6360 ( .A(n4652), .Z(n4868) );
  NANDN U6361 ( .A(n4651), .B(n4456), .Z(n4457) );
  XOR U6362 ( .A(n4868), .B(n4457), .Z(out[804]) );
  XNOR U6363 ( .A(n4458), .B(in[716]), .Z(n4872) );
  NANDN U6364 ( .A(n4654), .B(n4459), .Z(n4460) );
  XNOR U6365 ( .A(n4872), .B(n4460), .Z(out[805]) );
  XNOR U6366 ( .A(n4461), .B(in[717]), .Z(n4876) );
  NANDN U6367 ( .A(n4659), .B(n4462), .Z(n4463) );
  XNOR U6368 ( .A(n4876), .B(n4463), .Z(out[806]) );
  XNOR U6369 ( .A(n4464), .B(in[718]), .Z(n4880) );
  NANDN U6370 ( .A(n4660), .B(n4465), .Z(n4466) );
  XNOR U6371 ( .A(n4880), .B(n4466), .Z(out[807]) );
  XNOR U6372 ( .A(n4467), .B(in[719]), .Z(n4884) );
  NANDN U6373 ( .A(n4661), .B(n4468), .Z(n4469) );
  XNOR U6374 ( .A(n4884), .B(n4469), .Z(out[808]) );
  XNOR U6375 ( .A(n4470), .B(in[720]), .Z(n4888) );
  NANDN U6376 ( .A(n4662), .B(n4471), .Z(n4472) );
  XNOR U6377 ( .A(n4888), .B(n4472), .Z(out[809]) );
  ANDN U6378 ( .B(n4474), .A(n4473), .Z(n4475) );
  XOR U6379 ( .A(n4476), .B(n4475), .Z(out[80]) );
  XNOR U6380 ( .A(n4477), .B(in[721]), .Z(n4892) );
  NANDN U6381 ( .A(n4663), .B(n4478), .Z(n4479) );
  XNOR U6382 ( .A(n4892), .B(n4479), .Z(out[810]) );
  XNOR U6383 ( .A(n4480), .B(in[722]), .Z(n4896) );
  NAND U6384 ( .A(n4481), .B(n4664), .Z(n4482) );
  XNOR U6385 ( .A(n4896), .B(n4482), .Z(out[811]) );
  XNOR U6386 ( .A(n4483), .B(in[723]), .Z(n4903) );
  NANDN U6387 ( .A(n4666), .B(n4484), .Z(n4485) );
  XNOR U6388 ( .A(n4903), .B(n4485), .Z(out[812]) );
  XNOR U6389 ( .A(in[724]), .B(n4486), .Z(n4907) );
  NANDN U6390 ( .A(n4667), .B(n4487), .Z(n4488) );
  XNOR U6391 ( .A(n4907), .B(n4488), .Z(out[813]) );
  XNOR U6392 ( .A(in[725]), .B(n4489), .Z(n4911) );
  NANDN U6393 ( .A(n4668), .B(n4490), .Z(n4491) );
  XNOR U6394 ( .A(n4911), .B(n4491), .Z(out[814]) );
  XNOR U6395 ( .A(in[726]), .B(n4492), .Z(n4915) );
  NANDN U6396 ( .A(n4669), .B(n4493), .Z(n4494) );
  XNOR U6397 ( .A(n4915), .B(n4494), .Z(out[815]) );
  XNOR U6398 ( .A(in[727]), .B(n4495), .Z(n4919) );
  NANDN U6399 ( .A(n4673), .B(n4496), .Z(n4497) );
  XNOR U6400 ( .A(n4919), .B(n4497), .Z(out[816]) );
  XNOR U6401 ( .A(in[728]), .B(n4498), .Z(n4923) );
  NANDN U6402 ( .A(n4674), .B(n4499), .Z(n4500) );
  XNOR U6403 ( .A(n4923), .B(n4500), .Z(out[817]) );
  XNOR U6404 ( .A(in[729]), .B(n4501), .Z(n4927) );
  NANDN U6405 ( .A(n4675), .B(n4502), .Z(n4503) );
  XNOR U6406 ( .A(n4927), .B(n4503), .Z(out[818]) );
  XNOR U6407 ( .A(in[730]), .B(n4504), .Z(n4931) );
  NANDN U6408 ( .A(n4676), .B(n4505), .Z(n4506) );
  XNOR U6409 ( .A(n4931), .B(n4506), .Z(out[819]) );
  ANDN U6410 ( .B(n4508), .A(n4507), .Z(n4509) );
  XOR U6411 ( .A(n4510), .B(n4509), .Z(out[81]) );
  XOR U6412 ( .A(in[731]), .B(n4511), .Z(n4935) );
  NANDN U6413 ( .A(n4677), .B(n4512), .Z(n4513) );
  XNOR U6414 ( .A(n4935), .B(n4513), .Z(out[820]) );
  XOR U6415 ( .A(in[732]), .B(n4514), .Z(n4939) );
  NANDN U6416 ( .A(n4678), .B(n4515), .Z(n4516) );
  XNOR U6417 ( .A(n4939), .B(n4516), .Z(out[821]) );
  XOR U6418 ( .A(in[733]), .B(n4517), .Z(n4947) );
  NANDN U6419 ( .A(n4679), .B(n4518), .Z(n4519) );
  XNOR U6420 ( .A(n4947), .B(n4519), .Z(out[822]) );
  XNOR U6421 ( .A(in[734]), .B(n4520), .Z(n4951) );
  IV U6422 ( .A(n4521), .Z(n4680) );
  NANDN U6423 ( .A(n4522), .B(n4680), .Z(n4523) );
  XNOR U6424 ( .A(n4951), .B(n4523), .Z(out[823]) );
  XNOR U6425 ( .A(in[735]), .B(n4524), .Z(n4955) );
  IV U6426 ( .A(n4525), .Z(n4682) );
  NANDN U6427 ( .A(n4526), .B(n4682), .Z(n4527) );
  XNOR U6428 ( .A(n4955), .B(n4527), .Z(out[824]) );
  XNOR U6429 ( .A(in[736]), .B(n4528), .Z(n4959) );
  IV U6430 ( .A(n4529), .Z(n4684) );
  NANDN U6431 ( .A(n4530), .B(n4684), .Z(n4531) );
  XNOR U6432 ( .A(n4959), .B(n4531), .Z(out[825]) );
  XNOR U6433 ( .A(in[737]), .B(n4532), .Z(n4963) );
  IV U6434 ( .A(n4533), .Z(n4690) );
  NANDN U6435 ( .A(n4534), .B(n4690), .Z(n4535) );
  XNOR U6436 ( .A(n4963), .B(n4535), .Z(out[826]) );
  XNOR U6437 ( .A(in[738]), .B(n4536), .Z(n4967) );
  IV U6438 ( .A(n4537), .Z(n4692) );
  NANDN U6439 ( .A(n4538), .B(n4692), .Z(n4539) );
  XNOR U6440 ( .A(n4967), .B(n4539), .Z(out[827]) );
  XNOR U6441 ( .A(in[739]), .B(n4540), .Z(n4971) );
  IV U6442 ( .A(n4541), .Z(n4694) );
  NANDN U6443 ( .A(n4542), .B(n4694), .Z(n4543) );
  XNOR U6444 ( .A(n4971), .B(n4543), .Z(out[828]) );
  XOR U6445 ( .A(in[740]), .B(n4544), .Z(n4697) );
  IV U6446 ( .A(n4697), .Z(n4975) );
  ANDN U6447 ( .B(n4547), .A(n4546), .Z(n4548) );
  XOR U6448 ( .A(n4549), .B(n4548), .Z(out[82]) );
  XOR U6449 ( .A(in[741]), .B(n4550), .Z(n4700) );
  IV U6450 ( .A(n4700), .Z(n4979) );
  XOR U6451 ( .A(in[742]), .B(n4552), .Z(n4703) );
  IV U6452 ( .A(n4703), .Z(n4983) );
  NANDN U6453 ( .A(n4555), .B(n4554), .Z(n4556) );
  XOR U6454 ( .A(n4706), .B(n4556), .Z(out[832]) );
  NANDN U6455 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U6456 ( .A(n4710), .B(n4559), .Z(out[833]) );
  NANDN U6457 ( .A(n4561), .B(n4560), .Z(n4562) );
  XOR U6458 ( .A(n4714), .B(n4562), .Z(out[834]) );
  NANDN U6459 ( .A(n4564), .B(n4563), .Z(n4565) );
  XOR U6460 ( .A(n4718), .B(n4565), .Z(out[835]) );
  NANDN U6461 ( .A(n4566), .B(n4729), .Z(n4567) );
  XOR U6462 ( .A(n4730), .B(n4567), .Z(out[836]) );
  NANDN U6463 ( .A(n4568), .B(n4733), .Z(n4569) );
  XOR U6464 ( .A(n4734), .B(n4569), .Z(out[837]) );
  NANDN U6465 ( .A(n4570), .B(n4737), .Z(n4571) );
  XOR U6466 ( .A(n4738), .B(n4571), .Z(out[838]) );
  NANDN U6467 ( .A(n4573), .B(n4572), .Z(n4574) );
  XOR U6468 ( .A(n4742), .B(n4574), .Z(out[839]) );
  ANDN U6469 ( .B(n4576), .A(n4575), .Z(n4577) );
  XOR U6470 ( .A(n4578), .B(n4577), .Z(out[83]) );
  NANDN U6471 ( .A(n4579), .B(n4746), .Z(n4580) );
  XNOR U6472 ( .A(n4745), .B(n4580), .Z(out[840]) );
  NANDN U6473 ( .A(n4581), .B(n4750), .Z(n4582) );
  XNOR U6474 ( .A(n4749), .B(n4582), .Z(out[841]) );
  NANDN U6475 ( .A(n4583), .B(n4754), .Z(n4584) );
  XNOR U6476 ( .A(n4753), .B(n4584), .Z(out[842]) );
  NANDN U6477 ( .A(n4585), .B(n4758), .Z(n4586) );
  XNOR U6478 ( .A(n4757), .B(n4586), .Z(out[843]) );
  NANDN U6479 ( .A(n4587), .B(n4762), .Z(n4588) );
  XNOR U6480 ( .A(n4761), .B(n4588), .Z(out[844]) );
  NANDN U6481 ( .A(n4589), .B(n4766), .Z(n4590) );
  XNOR U6482 ( .A(n4765), .B(n4590), .Z(out[845]) );
  NANDN U6483 ( .A(n4591), .B(n4773), .Z(n4592) );
  XNOR U6484 ( .A(n4772), .B(n4592), .Z(out[846]) );
  NANDN U6485 ( .A(n4593), .B(n4777), .Z(n4594) );
  XNOR U6486 ( .A(n4776), .B(n4594), .Z(out[847]) );
  NANDN U6487 ( .A(n4596), .B(n4595), .Z(n4597) );
  XNOR U6488 ( .A(n4780), .B(n4597), .Z(out[848]) );
  NANDN U6489 ( .A(n4598), .B(n4785), .Z(n4599) );
  XNOR U6490 ( .A(n4784), .B(n4599), .Z(out[849]) );
  ANDN U6491 ( .B(n4601), .A(n4600), .Z(n4602) );
  XOR U6492 ( .A(n4603), .B(n4602), .Z(out[84]) );
  NANDN U6493 ( .A(n4604), .B(n4789), .Z(n4605) );
  XNOR U6494 ( .A(n4788), .B(n4605), .Z(out[850]) );
  NANDN U6495 ( .A(n4606), .B(n4793), .Z(n4607) );
  XNOR U6496 ( .A(n4792), .B(n4607), .Z(out[851]) );
  NANDN U6497 ( .A(n4608), .B(n4797), .Z(n4609) );
  XNOR U6498 ( .A(n4796), .B(n4609), .Z(out[852]) );
  NANDN U6499 ( .A(n4610), .B(n4801), .Z(n4611) );
  XNOR U6500 ( .A(n4800), .B(n4611), .Z(out[853]) );
  NANDN U6501 ( .A(n4612), .B(n4805), .Z(n4613) );
  XNOR U6502 ( .A(n4804), .B(n4613), .Z(out[854]) );
  NANDN U6503 ( .A(n4615), .B(n4614), .Z(n4616) );
  XNOR U6504 ( .A(n4808), .B(n4616), .Z(out[855]) );
  NANDN U6505 ( .A(n4617), .B(n4816), .Z(n4618) );
  XNOR U6506 ( .A(n4815), .B(n4618), .Z(out[856]) );
  NANDN U6507 ( .A(n4619), .B(n4820), .Z(n4620) );
  XNOR U6508 ( .A(n4819), .B(n4620), .Z(out[857]) );
  NANDN U6509 ( .A(n4621), .B(n4824), .Z(n4622) );
  XNOR U6510 ( .A(n4823), .B(n4622), .Z(out[858]) );
  NANDN U6511 ( .A(n4623), .B(n4828), .Z(n4624) );
  XNOR U6512 ( .A(n4827), .B(n4624), .Z(out[859]) );
  ANDN U6513 ( .B(n4626), .A(n4625), .Z(n4627) );
  XOR U6514 ( .A(n4628), .B(n4627), .Z(out[85]) );
  NANDN U6515 ( .A(n4630), .B(n4629), .Z(n4631) );
  XNOR U6516 ( .A(n4831), .B(n4631), .Z(out[860]) );
  NANDN U6517 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U6518 ( .A(n4835), .B(n4634), .Z(out[861]) );
  NANDN U6519 ( .A(n4636), .B(n4635), .Z(n4637) );
  XNOR U6520 ( .A(n4839), .B(n4637), .Z(out[862]) );
  NANDN U6521 ( .A(n4640), .B(n4639), .Z(n4641) );
  XNOR U6522 ( .A(n4847), .B(n4641), .Z(out[864]) );
  NANDN U6523 ( .A(n4643), .B(n4642), .Z(n4644) );
  XNOR U6524 ( .A(n4851), .B(n4644), .Z(out[865]) );
  NANDN U6525 ( .A(n4646), .B(n4645), .Z(n4647) );
  XNOR U6526 ( .A(n4859), .B(n4647), .Z(out[866]) );
  NANDN U6527 ( .A(n4649), .B(n4648), .Z(n4650) );
  XNOR U6528 ( .A(n4863), .B(n4650), .Z(out[867]) );
  NANDN U6529 ( .A(n4652), .B(n4651), .Z(n4653) );
  XNOR U6530 ( .A(n4867), .B(n4653), .Z(out[868]) );
  ANDN U6531 ( .B(n4656), .A(n4655), .Z(n4657) );
  XOR U6532 ( .A(n4658), .B(n4657), .Z(out[86]) );
  OR U6533 ( .A(n4896), .B(n4664), .Z(n4665) );
  XNOR U6534 ( .A(n4895), .B(n4665), .Z(out[875]) );
  OR U6535 ( .A(n4951), .B(n4680), .Z(n4681) );
  XOR U6536 ( .A(n4952), .B(n4681), .Z(out[887]) );
  OR U6537 ( .A(n4955), .B(n4682), .Z(n4683) );
  XOR U6538 ( .A(n4956), .B(n4683), .Z(out[888]) );
  OR U6539 ( .A(n4959), .B(n4684), .Z(n4685) );
  XOR U6540 ( .A(n4960), .B(n4685), .Z(out[889]) );
  ANDN U6541 ( .B(n4687), .A(n4686), .Z(n4688) );
  XOR U6542 ( .A(n4689), .B(n4688), .Z(out[88]) );
  OR U6543 ( .A(n4963), .B(n4690), .Z(n4691) );
  XOR U6544 ( .A(n4964), .B(n4691), .Z(out[890]) );
  OR U6545 ( .A(n4967), .B(n4692), .Z(n4693) );
  XOR U6546 ( .A(n4968), .B(n4693), .Z(out[891]) );
  OR U6547 ( .A(n4971), .B(n4694), .Z(n4695) );
  XOR U6548 ( .A(n4972), .B(n4695), .Z(out[892]) );
  NANDN U6549 ( .A(n4697), .B(n4696), .Z(n4698) );
  XOR U6550 ( .A(n4976), .B(n4698), .Z(out[893]) );
  NANDN U6551 ( .A(n4700), .B(n4699), .Z(n4701) );
  XOR U6552 ( .A(n4980), .B(n4701), .Z(out[894]) );
  NANDN U6553 ( .A(n4703), .B(n4702), .Z(n4704) );
  XOR U6554 ( .A(n4984), .B(n4704), .Z(out[895]) );
  ANDN U6555 ( .B(n4706), .A(n4705), .Z(n4707) );
  XOR U6556 ( .A(n4708), .B(n4707), .Z(out[896]) );
  ANDN U6557 ( .B(n4710), .A(n4709), .Z(n4711) );
  XOR U6558 ( .A(n4712), .B(n4711), .Z(out[897]) );
  ANDN U6559 ( .B(n4714), .A(n4713), .Z(n4715) );
  XOR U6560 ( .A(n4716), .B(n4715), .Z(out[898]) );
  ANDN U6561 ( .B(n4718), .A(n4717), .Z(n4719) );
  XOR U6562 ( .A(n4720), .B(n4719), .Z(out[899]) );
  ANDN U6563 ( .B(n4722), .A(n4721), .Z(n4723) );
  XOR U6564 ( .A(n4724), .B(n4723), .Z(out[89]) );
  OR U6565 ( .A(n4726), .B(n4725), .Z(n4727) );
  XNOR U6566 ( .A(n4728), .B(n4727), .Z(out[8]) );
  ANDN U6567 ( .B(n4730), .A(n4729), .Z(n4731) );
  XOR U6568 ( .A(n4732), .B(n4731), .Z(out[900]) );
  ANDN U6569 ( .B(n4734), .A(n4733), .Z(n4735) );
  XOR U6570 ( .A(n4736), .B(n4735), .Z(out[901]) );
  ANDN U6571 ( .B(n4738), .A(n4737), .Z(n4739) );
  XOR U6572 ( .A(n4740), .B(n4739), .Z(out[902]) );
  ANDN U6573 ( .B(n4742), .A(n4741), .Z(n4743) );
  XOR U6574 ( .A(n4744), .B(n4743), .Z(out[903]) );
  NOR U6575 ( .A(n4746), .B(n4745), .Z(n4747) );
  XOR U6576 ( .A(n4748), .B(n4747), .Z(out[904]) );
  NOR U6577 ( .A(n4750), .B(n4749), .Z(n4751) );
  XOR U6578 ( .A(n4752), .B(n4751), .Z(out[905]) );
  NOR U6579 ( .A(n4754), .B(n4753), .Z(n4755) );
  XOR U6580 ( .A(n4756), .B(n4755), .Z(out[906]) );
  NOR U6581 ( .A(n4758), .B(n4757), .Z(n4759) );
  XOR U6582 ( .A(n4760), .B(n4759), .Z(out[907]) );
  NOR U6583 ( .A(n4762), .B(n4761), .Z(n4763) );
  XOR U6584 ( .A(n4764), .B(n4763), .Z(out[908]) );
  NOR U6585 ( .A(n4766), .B(n4765), .Z(n4767) );
  XOR U6586 ( .A(n4768), .B(n4767), .Z(out[909]) );
  NOR U6587 ( .A(n4773), .B(n4772), .Z(n4774) );
  XOR U6588 ( .A(n4775), .B(n4774), .Z(out[910]) );
  NOR U6589 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U6590 ( .A(n4779), .B(n4778), .Z(out[911]) );
  NOR U6591 ( .A(n4781), .B(n4780), .Z(n4782) );
  XOR U6592 ( .A(n4783), .B(n4782), .Z(out[912]) );
  NOR U6593 ( .A(n4785), .B(n4784), .Z(n4786) );
  XOR U6594 ( .A(n4787), .B(n4786), .Z(out[913]) );
  NOR U6595 ( .A(n4789), .B(n4788), .Z(n4790) );
  XOR U6596 ( .A(n4791), .B(n4790), .Z(out[914]) );
  NOR U6597 ( .A(n4793), .B(n4792), .Z(n4794) );
  XOR U6598 ( .A(n4795), .B(n4794), .Z(out[915]) );
  NOR U6599 ( .A(n4797), .B(n4796), .Z(n4798) );
  XOR U6600 ( .A(n4799), .B(n4798), .Z(out[916]) );
  NOR U6601 ( .A(n4801), .B(n4800), .Z(n4802) );
  XOR U6602 ( .A(n4803), .B(n4802), .Z(out[917]) );
  NOR U6603 ( .A(n4805), .B(n4804), .Z(n4806) );
  XOR U6604 ( .A(n4807), .B(n4806), .Z(out[918]) );
  NOR U6605 ( .A(n4809), .B(n4808), .Z(n4810) );
  XOR U6606 ( .A(n4811), .B(n4810), .Z(out[919]) );
  NOR U6607 ( .A(n4816), .B(n4815), .Z(n4817) );
  XOR U6608 ( .A(n4818), .B(n4817), .Z(out[920]) );
  NOR U6609 ( .A(n4820), .B(n4819), .Z(n4821) );
  XOR U6610 ( .A(n4822), .B(n4821), .Z(out[921]) );
  NOR U6611 ( .A(n4824), .B(n4823), .Z(n4825) );
  XOR U6612 ( .A(n4826), .B(n4825), .Z(out[922]) );
  NOR U6613 ( .A(n4828), .B(n4827), .Z(n4829) );
  XOR U6614 ( .A(n4830), .B(n4829), .Z(out[923]) );
  NOR U6615 ( .A(n4832), .B(n4831), .Z(n4833) );
  XOR U6616 ( .A(n4834), .B(n4833), .Z(out[924]) );
  NOR U6617 ( .A(n4836), .B(n4835), .Z(n4837) );
  XOR U6618 ( .A(n4838), .B(n4837), .Z(out[925]) );
  NOR U6619 ( .A(n4840), .B(n4839), .Z(n4841) );
  XOR U6620 ( .A(n4842), .B(n4841), .Z(out[926]) );
  NOR U6621 ( .A(n4844), .B(n4843), .Z(n4845) );
  XOR U6622 ( .A(n4846), .B(n4845), .Z(out[927]) );
  NOR U6623 ( .A(n4848), .B(n4847), .Z(n4849) );
  XOR U6624 ( .A(n4850), .B(n4849), .Z(out[928]) );
  NOR U6625 ( .A(n4852), .B(n4851), .Z(n4853) );
  XOR U6626 ( .A(n4854), .B(n4853), .Z(out[929]) );
  AND U6627 ( .A(n4856), .B(n4855), .Z(n4857) );
  XNOR U6628 ( .A(n4858), .B(n4857), .Z(out[92]) );
  NOR U6629 ( .A(n4860), .B(n4859), .Z(n4861) );
  XOR U6630 ( .A(n4862), .B(n4861), .Z(out[930]) );
  NOR U6631 ( .A(n4864), .B(n4863), .Z(n4865) );
  XOR U6632 ( .A(n4866), .B(n4865), .Z(out[931]) );
  NOR U6633 ( .A(n4868), .B(n4867), .Z(n4869) );
  XOR U6634 ( .A(n4870), .B(n4869), .Z(out[932]) );
  ANDN U6635 ( .B(n4872), .A(n4871), .Z(n4873) );
  XOR U6636 ( .A(n4874), .B(n4873), .Z(out[933]) );
  ANDN U6637 ( .B(n4876), .A(n4875), .Z(n4877) );
  XOR U6638 ( .A(n4878), .B(n4877), .Z(out[934]) );
  ANDN U6639 ( .B(n4880), .A(n4879), .Z(n4881) );
  XOR U6640 ( .A(n4882), .B(n4881), .Z(out[935]) );
  ANDN U6641 ( .B(n4884), .A(n4883), .Z(n4885) );
  XOR U6642 ( .A(n4886), .B(n4885), .Z(out[936]) );
  ANDN U6643 ( .B(n4888), .A(n4887), .Z(n4889) );
  XOR U6644 ( .A(n4890), .B(n4889), .Z(out[937]) );
  ANDN U6645 ( .B(n4892), .A(n4891), .Z(n4893) );
  XOR U6646 ( .A(n4894), .B(n4893), .Z(out[938]) );
  ANDN U6647 ( .B(n4896), .A(n4895), .Z(n4897) );
  XOR U6648 ( .A(n4898), .B(n4897), .Z(out[939]) );
  AND U6649 ( .A(n4900), .B(n4899), .Z(n4901) );
  XNOR U6650 ( .A(n4902), .B(n4901), .Z(out[93]) );
  AND U6651 ( .A(n4904), .B(n4903), .Z(n4905) );
  XNOR U6652 ( .A(n4906), .B(n4905), .Z(out[940]) );
  AND U6653 ( .A(n4908), .B(n4907), .Z(n4909) );
  XNOR U6654 ( .A(n4910), .B(n4909), .Z(out[941]) );
  AND U6655 ( .A(n4912), .B(n4911), .Z(n4913) );
  XNOR U6656 ( .A(n4914), .B(n4913), .Z(out[942]) );
  AND U6657 ( .A(n4916), .B(n4915), .Z(n4917) );
  XNOR U6658 ( .A(n4918), .B(n4917), .Z(out[943]) );
  AND U6659 ( .A(n4920), .B(n4919), .Z(n4921) );
  XNOR U6660 ( .A(n4922), .B(n4921), .Z(out[944]) );
  AND U6661 ( .A(n4924), .B(n4923), .Z(n4925) );
  XNOR U6662 ( .A(n4926), .B(n4925), .Z(out[945]) );
  AND U6663 ( .A(n4928), .B(n4927), .Z(n4929) );
  XNOR U6664 ( .A(n4930), .B(n4929), .Z(out[946]) );
  AND U6665 ( .A(n4932), .B(n4931), .Z(n4933) );
  XNOR U6666 ( .A(n4934), .B(n4933), .Z(out[947]) );
  AND U6667 ( .A(n4936), .B(n4935), .Z(n4937) );
  XNOR U6668 ( .A(n4938), .B(n4937), .Z(out[948]) );
  AND U6669 ( .A(n4940), .B(n4939), .Z(n4941) );
  XNOR U6670 ( .A(n4942), .B(n4941), .Z(out[949]) );
  AND U6671 ( .A(n4944), .B(n4943), .Z(n4945) );
  XNOR U6672 ( .A(n4946), .B(n4945), .Z(out[94]) );
  AND U6673 ( .A(n4948), .B(n4947), .Z(n4949) );
  XNOR U6674 ( .A(n4950), .B(n4949), .Z(out[950]) );
  AND U6675 ( .A(n4952), .B(n4951), .Z(n4953) );
  XNOR U6676 ( .A(n4954), .B(n4953), .Z(out[951]) );
  AND U6677 ( .A(n4956), .B(n4955), .Z(n4957) );
  XNOR U6678 ( .A(n4958), .B(n4957), .Z(out[952]) );
  AND U6679 ( .A(n4960), .B(n4959), .Z(n4961) );
  XNOR U6680 ( .A(n4962), .B(n4961), .Z(out[953]) );
  AND U6681 ( .A(n4964), .B(n4963), .Z(n4965) );
  XNOR U6682 ( .A(n4966), .B(n4965), .Z(out[954]) );
  AND U6683 ( .A(n4968), .B(n4967), .Z(n4969) );
  XNOR U6684 ( .A(n4970), .B(n4969), .Z(out[955]) );
  AND U6685 ( .A(n4972), .B(n4971), .Z(n4973) );
  XOR U6686 ( .A(n4974), .B(n4973), .Z(out[956]) );
  ANDN U6687 ( .B(n4976), .A(n4975), .Z(n4977) );
  XOR U6688 ( .A(n4978), .B(n4977), .Z(out[957]) );
  ANDN U6689 ( .B(n4980), .A(n4979), .Z(n4981) );
  XOR U6690 ( .A(n4982), .B(n4981), .Z(out[958]) );
  ANDN U6691 ( .B(n4984), .A(n4983), .Z(n4985) );
  XNOR U6692 ( .A(n4986), .B(n4985), .Z(out[959]) );
  AND U6693 ( .A(n4988), .B(n4987), .Z(n4989) );
  XNOR U6694 ( .A(n4990), .B(n4989), .Z(out[95]) );
  ANDN U6695 ( .B(n4992), .A(n4991), .Z(n4993) );
  XOR U6696 ( .A(n4994), .B(n4993), .Z(out[960]) );
  ANDN U6697 ( .B(n4996), .A(n4995), .Z(n4997) );
  XOR U6698 ( .A(n4998), .B(n4997), .Z(out[961]) );
  ANDN U6699 ( .B(n5000), .A(n4999), .Z(n5001) );
  XOR U6700 ( .A(n5002), .B(n5001), .Z(out[962]) );
  ANDN U6701 ( .B(n5004), .A(n5003), .Z(n5005) );
  XOR U6702 ( .A(n5006), .B(n5005), .Z(out[963]) );
  ANDN U6703 ( .B(n5008), .A(n5007), .Z(n5009) );
  XOR U6704 ( .A(n5010), .B(n5009), .Z(out[964]) );
  ANDN U6705 ( .B(n5012), .A(n5011), .Z(n5013) );
  XOR U6706 ( .A(n5014), .B(n5013), .Z(out[965]) );
  ANDN U6707 ( .B(n5016), .A(n5015), .Z(n5017) );
  XOR U6708 ( .A(n5018), .B(n5017), .Z(out[966]) );
  ANDN U6709 ( .B(n5020), .A(n5019), .Z(n5021) );
  XOR U6710 ( .A(n5022), .B(n5021), .Z(out[967]) );
  ANDN U6711 ( .B(n5024), .A(n5023), .Z(n5025) );
  XOR U6712 ( .A(n5026), .B(n5025), .Z(out[968]) );
  ANDN U6713 ( .B(n5028), .A(n5027), .Z(n5029) );
  XOR U6714 ( .A(n5030), .B(n5029), .Z(out[969]) );
  AND U6715 ( .A(n5032), .B(n5031), .Z(n5033) );
  XNOR U6716 ( .A(n5034), .B(n5033), .Z(out[96]) );
  ANDN U6717 ( .B(n5036), .A(n5035), .Z(n5037) );
  XOR U6718 ( .A(n5038), .B(n5037), .Z(out[970]) );
  ANDN U6719 ( .B(n5040), .A(n5039), .Z(n5041) );
  XOR U6720 ( .A(n5042), .B(n5041), .Z(out[971]) );
  ANDN U6721 ( .B(n5044), .A(n5043), .Z(n5045) );
  XOR U6722 ( .A(n5046), .B(n5045), .Z(out[972]) );
  ANDN U6723 ( .B(n5048), .A(n5047), .Z(n5049) );
  XOR U6724 ( .A(n5050), .B(n5049), .Z(out[973]) );
  ANDN U6725 ( .B(n5052), .A(n5051), .Z(n5053) );
  XOR U6726 ( .A(n5054), .B(n5053), .Z(out[974]) );
  ANDN U6727 ( .B(n5056), .A(n5055), .Z(n5057) );
  XOR U6728 ( .A(n5058), .B(n5057), .Z(out[975]) );
  ANDN U6729 ( .B(n5069), .A(n5068), .Z(n5070) );
  XOR U6730 ( .A(n5071), .B(n5070), .Z(out[979]) );
  AND U6731 ( .A(n5073), .B(n5072), .Z(n5074) );
  XNOR U6732 ( .A(n5075), .B(n5074), .Z(out[97]) );
  ANDN U6733 ( .B(n5101), .A(n5100), .Z(n5102) );
  XOR U6734 ( .A(n5103), .B(n5102), .Z(out[988]) );
  ANDN U6735 ( .B(n5108), .A(n5107), .Z(n5109) );
  XNOR U6736 ( .A(n5110), .B(n5109), .Z(out[98]) );
  ANDN U6737 ( .B(n5115), .A(n5114), .Z(n5116) );
  XOR U6738 ( .A(n5117), .B(n5116), .Z(out[991]) );
  ANDN U6739 ( .B(n5119), .A(n5118), .Z(n5120) );
  XOR U6740 ( .A(n5121), .B(n5120), .Z(out[992]) );
  ANDN U6741 ( .B(n5123), .A(n5122), .Z(n5124) );
  XOR U6742 ( .A(n5125), .B(n5124), .Z(out[993]) );
  ANDN U6743 ( .B(n5127), .A(n5126), .Z(n5128) );
  XOR U6744 ( .A(n5129), .B(n5128), .Z(out[994]) );
  ANDN U6745 ( .B(n5131), .A(n5130), .Z(n5132) );
  XNOR U6746 ( .A(n5133), .B(n5132), .Z(out[995]) );
  ANDN U6747 ( .B(n5135), .A(n5134), .Z(n5136) );
  XNOR U6748 ( .A(n5137), .B(n5136), .Z(out[996]) );
  AND U6749 ( .A(n5142), .B(n5141), .Z(n5143) );
  XNOR U6750 ( .A(n5144), .B(n5143), .Z(out[998]) );
  ANDN U6751 ( .B(n5146), .A(n5145), .Z(n5147) );
  XNOR U6752 ( .A(n5148), .B(n5147), .Z(out[999]) );
  ANDN U6753 ( .B(n5150), .A(n5149), .Z(n5151) );
  XNOR U6754 ( .A(n5152), .B(n5151), .Z(out[99]) );
  OR U6755 ( .A(n5154), .B(n5153), .Z(n5155) );
  XNOR U6756 ( .A(n5156), .B(n5155), .Z(out[9]) );
endmodule


module round_5 ( in, round_const, out );
  input [1599:0] in;
  input [63:0] round_const;
  output [1599:0] out;
  wire   round_const_63, round_const_31, round_const_15, round_const_7,
         round_const_3, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164;
  assign round_const_63 = round_const[63];
  assign round_const_31 = round_const[31];
  assign round_const_15 = round_const[15];
  assign round_const_7 = round_const[7];
  assign round_const_3 = round_const[3];

  XNOR U1 ( .A(n1481), .B(n1147), .Z(n4056) );
  XOR U2 ( .A(n1396), .B(n1433), .Z(n4467) );
  NANDN U3 ( .A(n3281), .B(n3641), .Z(n1) );
  XNOR U4 ( .A(n3475), .B(n1), .Z(out[390]) );
  NANDN U5 ( .A(n3287), .B(n3649), .Z(n2) );
  XNOR U6 ( .A(n3481), .B(n2), .Z(out[392]) );
  ANDN U7 ( .B(n2508), .A(n2218), .Z(n3) );
  XNOR U8 ( .A(n2359), .B(n3), .Z(out[1363]) );
  ANDN U9 ( .B(n2529), .A(n2229), .Z(n4) );
  XNOR U10 ( .A(n2369), .B(n4), .Z(out[1368]) );
  NANDN U11 ( .A(n2250), .B(n2572), .Z(n5) );
  XNOR U12 ( .A(n2389), .B(n5), .Z(out[1378]) );
  NAND U13 ( .A(n2563), .B(n2388), .Z(n6) );
  XNOR U14 ( .A(n2564), .B(n6), .Z(out[1505]) );
  NANDN U15 ( .A(n2883), .B(n2882), .Z(n7) );
  XNOR U16 ( .A(n4338), .B(n7), .Z(out[268]) );
  XNOR U17 ( .A(n1449), .B(n1008), .Z(n2754) );
  XNOR U18 ( .A(n1461), .B(n1073), .Z(n2838) );
  XNOR U19 ( .A(n1475), .B(n1121), .Z(n2919) );
  XNOR U20 ( .A(n1728), .B(n1729), .Z(n3096) );
  XNOR U21 ( .A(n1405), .B(n1680), .Z(n3169) );
  XNOR U22 ( .A(n1411), .B(n1688), .Z(n3173) );
  XOR U23 ( .A(n794), .B(n1450), .Z(n4495) );
  XOR U24 ( .A(n820), .B(n1452), .Z(n4498) );
  XOR U25 ( .A(n1487), .B(n813), .Z(n4540) );
  XOR U26 ( .A(n1444), .B(n749), .Z(n4486) );
  XNOR U27 ( .A(n3940), .B(in[1481]), .Z(n4761) );
  XNOR U28 ( .A(n3964), .B(in[1487]), .Z(n4789) );
  NAND U29 ( .A(n4640), .B(n4851), .Z(n8) );
  XNOR U30 ( .A(n4850), .B(n8), .Z(out[863]) );
  NANDN U31 ( .A(n3284), .B(n3645), .Z(n9) );
  XNOR U32 ( .A(n3476), .B(n9), .Z(out[391]) );
  ANDN U33 ( .B(n2500), .A(n2214), .Z(n10) );
  XNOR U34 ( .A(n2354), .B(n10), .Z(out[1361]) );
  NANDN U35 ( .A(n4895), .B(n4668), .Z(n11) );
  XNOR U36 ( .A(n4894), .B(n11), .Z(out[873]) );
  ANDN U37 ( .B(n4675), .A(n4922), .Z(n12) );
  XNOR U38 ( .A(n4923), .B(n12), .Z(out[879]) );
  ANDN U39 ( .B(n4681), .A(n4934), .Z(n13) );
  XNOR U40 ( .A(n4935), .B(n13), .Z(out[882]) );
  ANDN U41 ( .B(n4682), .A(n4938), .Z(n14) );
  XNOR U42 ( .A(n4939), .B(n14), .Z(out[883]) );
  ANDN U43 ( .B(n2553), .A(n2241), .Z(n15) );
  XNOR U44 ( .A(n2382), .B(n15), .Z(out[1374]) );
  ANDN U45 ( .B(n5053), .A(n1644), .Z(n16) );
  XNOR U46 ( .A(n1839), .B(n16), .Z(out[1100]) );
  ANDN U47 ( .B(n2646), .A(n2288), .Z(n17) );
  XNOR U48 ( .A(n2410), .B(n17), .Z(out[1396]) );
  NAND U49 ( .A(n2569), .B(n2389), .Z(n18) );
  XNOR U50 ( .A(n2570), .B(n18), .Z(out[1506]) );
  NANDN U51 ( .A(n3275), .B(n3633), .Z(n19) );
  XNOR U52 ( .A(n3473), .B(n19), .Z(out[388]) );
  XNOR U53 ( .A(n1447), .B(n1754), .Z(n3215) );
  XNOR U54 ( .A(n1432), .B(n1725), .Z(n3194) );
  XNOR U55 ( .A(n1457), .B(n1047), .Z(n2792) );
  XNOR U56 ( .A(n1459), .B(n1060), .Z(n2815) );
  XNOR U57 ( .A(n1465), .B(n1088), .Z(n2862) );
  XNOR U58 ( .A(n1471), .B(n1101), .Z(n2886) );
  XNOR U59 ( .A(n1484), .B(n1160), .Z(n4060) );
  XNOR U60 ( .A(n1489), .B(n1190), .Z(n4072) );
  XNOR U61 ( .A(n1220), .B(n1495), .Z(n4080) );
  XNOR U62 ( .A(n1462), .B(n880), .Z(n4514) );
  XNOR U63 ( .A(n1466), .B(n895), .Z(n4517) );
  XNOR U64 ( .A(n1749), .B(n1750), .Z(n3102) );
  XNOR U65 ( .A(n1413), .B(n1692), .Z(n3175) );
  XOR U66 ( .A(n1392), .B(n1431), .Z(n4464) );
  XOR U67 ( .A(n1437), .B(n1404), .Z(n4477) );
  XNOR U68 ( .A(n3968), .B(in[1488]), .Z(n4793) );
  XNOR U69 ( .A(n3933), .B(in[1480]), .Z(n4757) );
  XNOR U70 ( .A(n3944), .B(in[1482]), .Z(n4765) );
  XNOR U71 ( .A(n3948), .B(in[1483]), .Z(n4769) );
  XNOR U72 ( .A(n3952), .B(in[1484]), .Z(n4773) );
  XNOR U73 ( .A(n3956), .B(in[1485]), .Z(n4781) );
  AND U74 ( .A(n2000), .B(n1591), .Z(n20) );
  XNOR U75 ( .A(n1806), .B(n20), .Z(out[1087]) );
  AND U76 ( .A(n4761), .B(n4363), .Z(n21) );
  XNOR U77 ( .A(n4583), .B(n21), .Z(out[714]) );
  AND U78 ( .A(n3420), .B(n2982), .Z(n22) );
  XNOR U79 ( .A(n3421), .B(n22), .Z(out[305]) );
  NAND U80 ( .A(n2601), .B(n2398), .Z(n23) );
  XNOR U81 ( .A(n2602), .B(n23), .Z(out[1514]) );
  ANDN U82 ( .B(n4672), .A(n4910), .Z(n24) );
  XNOR U83 ( .A(n4911), .B(n24), .Z(out[876]) );
  ANDN U84 ( .B(n4673), .A(n4914), .Z(n25) );
  XNOR U85 ( .A(n4915), .B(n25), .Z(out[877]) );
  ANDN U86 ( .B(n4679), .A(n4926), .Z(n26) );
  XNOR U87 ( .A(n4927), .B(n26), .Z(out[880]) );
  ANDN U88 ( .B(n4680), .A(n4930), .Z(n27) );
  XNOR U89 ( .A(n4931), .B(n27), .Z(out[881]) );
  NANDN U90 ( .A(n2847), .B(n3807), .Z(n28) );
  XNOR U91 ( .A(n3013), .B(n28), .Z(out[189]) );
  NANDN U92 ( .A(n2849), .B(n3851), .Z(n29) );
  XNOR U93 ( .A(n3014), .B(n29), .Z(out[190]) );
  AND U94 ( .A(n2493), .B(n2353), .Z(n30) );
  XNOR U95 ( .A(n2494), .B(n30), .Z(out[1488]) );
  AND U96 ( .A(n5065), .B(n1656), .Z(n31) );
  XNOR U97 ( .A(n1847), .B(n31), .Z(out[1103]) );
  ANDN U98 ( .B(n5085), .A(n1677), .Z(n32) );
  XNOR U99 ( .A(n1857), .B(n32), .Z(out[1108]) );
  NAND U100 ( .A(n2538), .B(n2375), .Z(n33) );
  XNOR U101 ( .A(n2539), .B(n33), .Z(out[1499]) );
  ANDN U102 ( .B(n2650), .A(n2290), .Z(n34) );
  XNOR U103 ( .A(n2412), .B(n34), .Z(out[1397]) );
  NAND U104 ( .A(n2581), .B(n2392), .Z(n35) );
  XNOR U105 ( .A(n2582), .B(n35), .Z(out[1509]) );
  ANDN U106 ( .B(n2672), .A(n2301), .Z(n36) );
  XNOR U107 ( .A(n2420), .B(n36), .Z(out[1402]) );
  AND U108 ( .A(n2619), .B(n2402), .Z(n37) );
  XNOR U109 ( .A(n2620), .B(n37), .Z(out[1518]) );
  AND U110 ( .A(n2623), .B(n2403), .Z(n38) );
  XNOR U111 ( .A(n2624), .B(n38), .Z(out[1519]) );
  NANDN U112 ( .A(n3278), .B(n3637), .Z(n39) );
  XNOR U113 ( .A(n3474), .B(n39), .Z(out[389]) );
  NOR U114 ( .A(n4572), .B(n4355), .Z(n40) );
  XNOR U115 ( .A(n4746), .B(n40), .Z(out[775]) );
  NANDN U116 ( .A(n2885), .B(n2884), .Z(n41) );
  XNOR U117 ( .A(n4369), .B(n41), .Z(out[269]) );
  NANDN U118 ( .A(n3980), .B(n3979), .Z(n42) );
  XNOR U119 ( .A(n3981), .B(n42), .Z(out[65]) );
  AND U120 ( .A(n4693), .B(n4692), .Z(n43) );
  XNOR U121 ( .A(n4694), .B(n43), .Z(out[88]) );
  ANDN U122 ( .B(n2433), .A(n2432), .Z(n44) );
  XNOR U123 ( .A(n2434), .B(round_const[0]), .Z(n45) );
  XOR U124 ( .A(n44), .B(n45), .Z(out[1536]) );
  ANDN U125 ( .B(n2467), .A(n2466), .Z(n46) );
  XNOR U126 ( .A(n2465), .B(n46), .Z(out[1544]) );
  ANDN U127 ( .B(n2473), .A(n2472), .Z(n47) );
  XNOR U128 ( .A(n2471), .B(n47), .Z(out[1546]) );
  XNOR U129 ( .A(n1445), .B(n1750), .Z(n3212) );
  XNOR U130 ( .A(n1658), .B(n1659), .Z(n3057) );
  XNOR U131 ( .A(n1675), .B(n1676), .Z(n3066) );
  XNOR U132 ( .A(n1428), .B(n1717), .Z(n2292) );
  XNOR U133 ( .A(n1439), .B(n1741), .Z(n3206) );
  XNOR U134 ( .A(n1443), .B(n1745), .Z(n3209) );
  XNOR U135 ( .A(n1691), .B(n1692), .Z(n3077) );
  XNOR U136 ( .A(n1703), .B(n1704), .Z(n3083) );
  XNOR U137 ( .A(n1479), .B(n1134), .Z(n4052) );
  XNOR U138 ( .A(n1460), .B(n865), .Z(n4511) );
  XNOR U139 ( .A(n1409), .B(n1684), .Z(n3171) );
  XNOR U140 ( .A(n1415), .B(n1696), .Z(n3177) );
  XNOR U141 ( .A(n1417), .B(n1700), .Z(n3179) );
  XNOR U142 ( .A(n1426), .B(n1713), .Z(n3185) );
  XNOR U143 ( .A(n1430), .B(n1721), .Z(n3192) );
  XNOR U144 ( .A(n1708), .B(n1350), .Z(n3929) );
  XOR U145 ( .A(n1384), .B(n1427), .Z(n4458) );
  XOR U146 ( .A(n1435), .B(n1400), .Z(n4470) );
  XOR U147 ( .A(n1482), .B(n685), .Z(n4532) );
  XNOR U148 ( .A(n3960), .B(in[1486]), .Z(n4785) );
  AND U149 ( .A(n4741), .B(n4349), .Z(n48) );
  XNOR U150 ( .A(n4568), .B(n48), .Z(out[709]) );
  NAND U151 ( .A(n4749), .B(n4355), .Z(n49) );
  XNOR U152 ( .A(n4572), .B(n49), .Z(out[711]) );
  NANDN U153 ( .A(n4459), .B(n4881), .Z(n50) );
  XNOR U154 ( .A(n4656), .B(n50), .Z(out[741]) );
  AND U155 ( .A(n4757), .B(n4360), .Z(n51) );
  XNOR U156 ( .A(n4581), .B(n51), .Z(out[713]) );
  NAND U157 ( .A(n2585), .B(n2394), .Z(n52) );
  XNOR U158 ( .A(n2586), .B(n52), .Z(out[1510]) );
  AND U159 ( .A(n2589), .B(n2395), .Z(n53) );
  XNOR U160 ( .A(n2590), .B(n53), .Z(out[1511]) );
  AND U161 ( .A(n2593), .B(n2396), .Z(n54) );
  XNOR U162 ( .A(n2594), .B(n54), .Z(out[1512]) );
  AND U163 ( .A(n2597), .B(n2397), .Z(n55) );
  XNOR U164 ( .A(n2598), .B(n55), .Z(out[1513]) );
  AND U165 ( .A(n3013), .B(n3804), .Z(n56) );
  XNOR U166 ( .A(n3805), .B(n56), .Z(out[317]) );
  ANDN U167 ( .B(n2512), .A(n2220), .Z(n57) );
  XNOR U168 ( .A(n2361), .B(n57), .Z(out[1364]) );
  ANDN U169 ( .B(n4674), .A(n4918), .Z(n58) );
  XNOR U170 ( .A(n4919), .B(n58), .Z(out[878]) );
  ANDN U171 ( .B(n4684), .A(n4946), .Z(n59) );
  XNOR U172 ( .A(n4947), .B(n59), .Z(out[885]) );
  ANDN U173 ( .B(n4685), .A(n4954), .Z(n60) );
  XNOR U174 ( .A(n4955), .B(n60), .Z(out[886]) );
  ANDN U175 ( .B(n2533), .A(n2231), .Z(n61) );
  XNOR U176 ( .A(n2371), .B(n61), .Z(out[1369]) );
  ANDN U177 ( .B(n5005), .A(n1599), .Z(n62) );
  XNOR U178 ( .A(n1812), .B(n62), .Z(out[1089]) );
  ANDN U179 ( .B(n5009), .A(n1603), .Z(n63) );
  XNOR U180 ( .A(n1815), .B(n63), .Z(out[1090]) );
  ANDN U181 ( .B(n5021), .A(n1615), .Z(n64) );
  XNOR U182 ( .A(n1826), .B(n64), .Z(out[1093]) );
  ANDN U183 ( .B(n5025), .A(n1619), .Z(n65) );
  XNOR U184 ( .A(n1828), .B(n65), .Z(out[1094]) );
  ANDN U185 ( .B(n2562), .A(n2246), .Z(n66) );
  XNOR U186 ( .A(n2386), .B(n66), .Z(out[1376]) );
  NANDN U187 ( .A(n2851), .B(n3895), .Z(n67) );
  XNOR U188 ( .A(n3017), .B(n67), .Z(out[191]) );
  ANDN U189 ( .B(n5045), .A(n1636), .Z(n68) );
  XNOR U190 ( .A(n1835), .B(n68), .Z(out[1098]) );
  NAND U191 ( .A(n2489), .B(n2351), .Z(n69) );
  XNOR U192 ( .A(n2488), .B(n69), .Z(out[1487]) );
  AND U193 ( .A(n5071), .B(n1664), .Z(n70) );
  XNOR U194 ( .A(n1851), .B(n70), .Z(out[1105]) );
  ANDN U195 ( .B(n5088), .A(n1681), .Z(n71) );
  XNOR U196 ( .A(n1859), .B(n71), .Z(out[1109]) );
  ANDN U197 ( .B(n5091), .A(n1685), .Z(n72) );
  XNOR U198 ( .A(n1861), .B(n72), .Z(out[1110]) );
  ANDN U199 ( .B(n5097), .A(n1693), .Z(n73) );
  XNOR U200 ( .A(n1867), .B(n73), .Z(out[1112]) );
  ANDN U201 ( .B(n5100), .A(n1697), .Z(n74) );
  XNOR U202 ( .A(n1869), .B(n74), .Z(out[1113]) );
  NAND U203 ( .A(n3835), .B(n3415), .Z(n75) );
  XNOR U204 ( .A(n3414), .B(n75), .Z(out[434]) );
  ANDN U205 ( .B(n2642), .A(n2285), .Z(n76) );
  XNOR U206 ( .A(n2408), .B(n76), .Z(out[1395]) );
  ANDN U207 ( .B(n3843), .A(n3426), .Z(n77) );
  XNOR U208 ( .A(n3584), .B(n77), .Z(out[436]) );
  ANDN U209 ( .B(n3847), .A(n3429), .Z(n78) );
  XNOR U210 ( .A(n3586), .B(n78), .Z(out[437]) );
  ANDN U211 ( .B(n3855), .A(n3432), .Z(n79) );
  XNOR U212 ( .A(n3588), .B(n79), .Z(out[438]) );
  NAND U213 ( .A(n2573), .B(n2390), .Z(n80) );
  XNOR U214 ( .A(n2574), .B(n80), .Z(out[1507]) );
  NAND U215 ( .A(n2577), .B(n2391), .Z(n81) );
  XNOR U216 ( .A(n2578), .B(n81), .Z(out[1508]) );
  ANDN U217 ( .B(n3867), .A(n3441), .Z(n82) );
  XNOR U218 ( .A(n3594), .B(n82), .Z(out[441]) );
  NANDN U219 ( .A(n3444), .B(n3871), .Z(n83) );
  XNOR U220 ( .A(n3600), .B(n83), .Z(out[442]) );
  ANDN U221 ( .B(n5136), .A(n1734), .Z(n84) );
  XNOR U222 ( .A(n1889), .B(n84), .Z(out[1122]) );
  NANDN U223 ( .A(n3447), .B(n3875), .Z(n85) );
  XNOR U224 ( .A(n3601), .B(n85), .Z(out[443]) );
  ANDN U225 ( .B(n3883), .A(n3453), .Z(n86) );
  XNOR U226 ( .A(n3604), .B(n86), .Z(out[445]) );
  AND U227 ( .A(n2605), .B(n2399), .Z(n87) );
  XNOR U228 ( .A(n2606), .B(n87), .Z(out[1515]) );
  AND U229 ( .A(n2611), .B(n2400), .Z(n88) );
  XNOR U230 ( .A(n2612), .B(n88), .Z(out[1516]) );
  ANDN U231 ( .B(n2401), .A(n2615), .Z(n89) );
  XNOR U232 ( .A(n2616), .B(n89), .Z(out[1517]) );
  ANDN U233 ( .B(n1996), .A(n1589), .Z(n90) );
  XNOR U234 ( .A(n1804), .B(n90), .Z(out[1086]) );
  AND U235 ( .A(n4745), .B(n4352), .Z(n91) );
  XNOR U236 ( .A(n4570), .B(n91), .Z(out[710]) );
  NAND U237 ( .A(n2896), .B(n4476), .Z(n92) );
  XNOR U238 ( .A(n2895), .B(n92), .Z(out[208]) );
  NAND U239 ( .A(n2899), .B(n4510), .Z(n93) );
  XNOR U240 ( .A(n2898), .B(n93), .Z(out[209]) );
  NANDN U241 ( .A(n2926), .B(n4729), .Z(n94) );
  XNOR U242 ( .A(n2925), .B(n94), .Z(out[217]) );
  NAND U243 ( .A(n3937), .B(n3936), .Z(n95) );
  XNOR U244 ( .A(n3938), .B(n95), .Z(out[64]) );
  AND U245 ( .A(n4629), .B(n4628), .Z(n96) );
  XNOR U246 ( .A(n4630), .B(n96), .Z(out[85]) );
  ANDN U247 ( .B(n2476), .A(n2475), .Z(n97) );
  XNOR U248 ( .A(n2474), .B(n97), .Z(out[1547]) );
  ANDN U249 ( .B(n2479), .A(n2478), .Z(n98) );
  XNOR U250 ( .A(n2477), .B(n98), .Z(out[1548]) );
  ANDN U251 ( .B(n2482), .A(n2481), .Z(n99) );
  XNOR U252 ( .A(n2480), .B(n99), .Z(out[1549]) );
  OR U253 ( .A(n5092), .B(n5093), .Z(n100) );
  XNOR U254 ( .A(n5094), .B(n100), .Z(out[983]) );
  XNOR U255 ( .A(n1662), .B(n1663), .Z(n3059) );
  XNOR U256 ( .A(n1436), .B(n1733), .Z(n3200) );
  XNOR U257 ( .A(n1683), .B(n1684), .Z(n3071) );
  XNOR U258 ( .A(n1451), .B(n1021), .Z(n2771) );
  XNOR U259 ( .A(n1695), .B(n1696), .Z(n3079) );
  XNOR U260 ( .A(n1699), .B(n1700), .Z(n3081) );
  XNOR U261 ( .A(n1716), .B(n1717), .Z(n3088) );
  XNOR U262 ( .A(n1492), .B(n1205), .Z(n4076) );
  XNOR U263 ( .A(n1753), .B(n1754), .Z(n3104) );
  XNOR U264 ( .A(n568), .B(n685), .Z(n4047) );
  XOR U265 ( .A(n1438), .B(n719), .Z(n4480) );
  XNOR U266 ( .A(n1422), .B(n1704), .Z(n3181) );
  XOR U267 ( .A(n1446), .B(n764), .Z(n4489) );
  XNOR U268 ( .A(n1424), .B(n1709), .Z(n3183) );
  XOR U269 ( .A(n1480), .B(n940), .Z(n4528) );
  XOR U270 ( .A(n702), .B(n1485), .Z(n4536) );
  XOR U271 ( .A(n734), .B(n1440), .Z(n4483) );
  XNOR U272 ( .A(n3972), .B(in[1489]), .Z(n4797) );
  ANDN U273 ( .B(n2545), .A(n2237), .Z(n101) );
  XNOR U274 ( .A(n2378), .B(n101), .Z(out[1372]) );
  ANDN U275 ( .B(n2549), .A(n2239), .Z(n102) );
  XNOR U276 ( .A(n2380), .B(n102), .Z(out[1373]) );
  AND U277 ( .A(n4765), .B(n4366), .Z(n103) );
  XNOR U278 ( .A(n4585), .B(n103), .Z(out[715]) );
  NAND U279 ( .A(n2854), .B(n2853), .Z(n104) );
  XNOR U280 ( .A(n3937), .B(n104), .Z(out[256]) );
  OR U281 ( .A(n5023), .B(n1828), .Z(n105) );
  XNOR U282 ( .A(n5022), .B(n105), .Z(out[1222]) );
  NANDN U283 ( .A(n4887), .B(n4666), .Z(n106) );
  XNOR U284 ( .A(n4886), .B(n106), .Z(out[871]) );
  NANDN U285 ( .A(n4891), .B(n4667), .Z(n107) );
  XNOR U286 ( .A(n4890), .B(n107), .Z(out[872]) );
  NANDN U287 ( .A(n4899), .B(n4669), .Z(n108) );
  XNOR U288 ( .A(n4898), .B(n108), .Z(out[874]) );
  ANDN U289 ( .B(n5001), .A(n1595), .Z(n109) );
  XNOR U290 ( .A(n1809), .B(n109), .Z(out[1088]) );
  ANDN U291 ( .B(n2537), .A(n2233), .Z(n110) );
  XNOR U292 ( .A(n2373), .B(n110), .Z(out[1370]) );
  ANDN U293 ( .B(n5017), .A(n1611), .Z(n111) );
  XNOR U294 ( .A(n1823), .B(n111), .Z(out[1092]) );
  ANDN U295 ( .B(n2556), .A(n2243), .Z(n112) );
  XNOR U296 ( .A(n2384), .B(n112), .Z(out[1375]) );
  ANDN U297 ( .B(n5037), .A(n1632), .Z(n113) );
  XNOR U298 ( .A(n1833), .B(n113), .Z(out[1097]) );
  ANDN U299 ( .B(n5049), .A(n1640), .Z(n114) );
  XNOR U300 ( .A(n1837), .B(n114), .Z(out[1099]) );
  ANDN U301 ( .B(n5057), .A(n1648), .Z(n115) );
  XNOR U302 ( .A(n1841), .B(n115), .Z(out[1101]) );
  AND U303 ( .A(n5068), .B(n1660), .Z(n116) );
  XNOR U304 ( .A(n1849), .B(n116), .Z(out[1104]) );
  ANDN U305 ( .B(n2452), .A(n2451), .Z(n117) );
  XNOR U306 ( .A(n2450), .B(n117), .Z(out[1540]) );
  ANDN U307 ( .B(n2455), .A(n2454), .Z(n118) );
  XNOR U308 ( .A(n2453), .B(n118), .Z(out[1541]) );
  ANDN U309 ( .B(n5103), .A(n1701), .Z(n119) );
  XNOR U310 ( .A(n1871), .B(n119), .Z(out[1114]) );
  ANDN U311 ( .B(n3859), .A(n3435), .Z(n120) );
  XNOR U312 ( .A(n3590), .B(n120), .Z(out[439]) );
  ANDN U313 ( .B(n3879), .A(n3450), .Z(n121) );
  XNOR U314 ( .A(n3602), .B(n121), .Z(out[444]) );
  AND U315 ( .A(n2627), .B(n2405), .Z(n122) );
  XNOR U316 ( .A(n2628), .B(n122), .Z(out[1520]) );
  AND U317 ( .A(n2653), .B(n2414), .Z(n123) );
  XNOR U318 ( .A(n2654), .B(n123), .Z(out[1526]) );
  AND U319 ( .A(n2661), .B(n2416), .Z(n124) );
  XNOR U320 ( .A(n2662), .B(n124), .Z(out[1528]) );
  NANDN U321 ( .A(n2209), .B(n2490), .Z(n125) );
  XNOR U322 ( .A(n2351), .B(n125), .Z(out[1359]) );
  NOR U323 ( .A(n4701), .B(n4545), .Z(n126) );
  XNOR U324 ( .A(n4982), .B(n126), .Z(out[829]) );
  NOR U325 ( .A(n4557), .B(n4336), .Z(n127) );
  XNOR U326 ( .A(n4714), .B(n127), .Z(out[769]) );
  NOR U327 ( .A(n4560), .B(n4342), .Z(n128) );
  XNOR U328 ( .A(n4718), .B(n128), .Z(out[770]) );
  NOR U329 ( .A(n4563), .B(n4344), .Z(n129) );
  XNOR U330 ( .A(n4722), .B(n129), .Z(out[771]) );
  ANDN U331 ( .B(n1984), .A(n1577), .Z(n130) );
  XNOR U332 ( .A(n1798), .B(n130), .Z(out[1083]) );
  NAND U333 ( .A(n2902), .B(n4549), .Z(n131) );
  XNOR U334 ( .A(n2901), .B(n131), .Z(out[210]) );
  NAND U335 ( .A(n2905), .B(n4578), .Z(n132) );
  XNOR U336 ( .A(n2904), .B(n132), .Z(out[211]) );
  NAND U337 ( .A(n2908), .B(n4603), .Z(n133) );
  XNOR U338 ( .A(n2907), .B(n133), .Z(out[212]) );
  NANDN U339 ( .A(n2914), .B(n4662), .Z(n134) );
  XNOR U340 ( .A(n2913), .B(n134), .Z(out[214]) );
  NANDN U341 ( .A(n2932), .B(n4821), .Z(n135) );
  XNOR U342 ( .A(n2931), .B(n135), .Z(out[219]) );
  ANDN U343 ( .B(n1904), .A(n1497), .Z(n136) );
  XNOR U344 ( .A(n1757), .B(n136), .Z(out[1064]) );
  ANDN U345 ( .B(n1908), .A(n1501), .Z(n137) );
  XNOR U346 ( .A(n1759), .B(n137), .Z(out[1065]) );
  ANDN U347 ( .B(n2950), .A(n5160), .Z(n138) );
  XNOR U348 ( .A(n3094), .B(n138), .Z(out[227]) );
  ANDN U349 ( .B(n1946), .A(n1539), .Z(n139) );
  XNOR U350 ( .A(n1778), .B(n139), .Z(out[1074]) );
  ANDN U351 ( .B(n1950), .A(n1543), .Z(n140) );
  XNOR U352 ( .A(n1780), .B(n140), .Z(out[1075]) );
  ANDN U353 ( .B(n1954), .A(n1549), .Z(n141) );
  XNOR U354 ( .A(n1782), .B(n141), .Z(out[1076]) );
  ANDN U355 ( .B(n1958), .A(n1553), .Z(n142) );
  XNOR U356 ( .A(n1784), .B(n142), .Z(out[1077]) );
  ANDN U357 ( .B(n1964), .A(n1557), .Z(n143) );
  XNOR U358 ( .A(n1786), .B(n143), .Z(out[1078]) );
  ANDN U359 ( .B(n1980), .A(n1573), .Z(n144) );
  XNOR U360 ( .A(n1796), .B(n144), .Z(out[1082]) );
  AND U361 ( .A(n4677), .B(n4676), .Z(n145) );
  XNOR U362 ( .A(n4678), .B(n145), .Z(out[87]) );
  NANDN U363 ( .A(n2881), .B(n2880), .Z(n146) );
  XNOR U364 ( .A(n4306), .B(n146), .Z(out[267]) );
  AND U365 ( .A(n4769), .B(n4373), .Z(n147) );
  XNOR U366 ( .A(n4587), .B(n147), .Z(out[716]) );
  OR U367 ( .A(n5072), .B(n5073), .Z(n148) );
  XNOR U368 ( .A(n5074), .B(n148), .Z(out[978]) );
  OR U369 ( .A(n5083), .B(n5084), .Z(n149) );
  XNOR U370 ( .A(n5085), .B(n149), .Z(out[980]) );
  OR U371 ( .A(n5086), .B(n5087), .Z(n150) );
  XNOR U372 ( .A(n5088), .B(n150), .Z(out[981]) );
  NANDN U373 ( .A(n1914), .B(n1763), .Z(n151) );
  XNOR U374 ( .A(n1913), .B(n151), .Z(out[1195]) );
  OR U375 ( .A(n5111), .B(n5112), .Z(n152) );
  XNOR U376 ( .A(n5113), .B(n152), .Z(out[989]) );
  NANDN U377 ( .A(n4430), .B(n4849), .Z(n153) );
  XNOR U378 ( .A(n4637), .B(n153), .Z(out[734]) );
  NANDN U379 ( .A(n4444), .B(n4857), .Z(n154) );
  XNOR U380 ( .A(n4641), .B(n154), .Z(out[736]) );
  NANDN U381 ( .A(n4450), .B(n4869), .Z(n155) );
  XNOR U382 ( .A(n4647), .B(n155), .Z(out[738]) );
  ANDN U383 ( .B(n3506), .A(n3702), .Z(n156) );
  XNOR U384 ( .A(n3703), .B(n156), .Z(out[533]) );
  ANDN U385 ( .B(n3510), .A(n3724), .Z(n157) );
  XNOR U386 ( .A(n3725), .B(n157), .Z(out[537]) );
  XNOR U387 ( .A(n1667), .B(n1668), .Z(n3061) );
  XNOR U388 ( .A(n1679), .B(n1680), .Z(n3069) );
  XNOR U389 ( .A(n1434), .B(n1729), .Z(n3197) );
  XNOR U390 ( .A(n1687), .B(n1688), .Z(n3075) );
  XNOR U391 ( .A(n1453), .B(n1034), .Z(n2778) );
  XNOR U392 ( .A(n1712), .B(n1713), .Z(n3086) );
  XNOR U393 ( .A(n1720), .B(n1721), .Z(n3090) );
  XNOR U394 ( .A(n1724), .B(n1725), .Z(n3092) );
  XNOR U395 ( .A(n1499), .B(n1235), .Z(n2211) );
  XOR U396 ( .A(n779), .B(n1448), .Z(n4492) );
  XOR U397 ( .A(n1454), .B(n835), .Z(n4501) );
  XOR U398 ( .A(n1458), .B(n850), .Z(n4504) );
  XOR U399 ( .A(n1388), .B(n1429), .Z(n4461) );
  XOR U400 ( .A(n1472), .B(n910), .Z(n4520) );
  XOR U401 ( .A(n1476), .B(n925), .Z(n4524) );
  XNOR U402 ( .A(n3976), .B(in[1490]), .Z(n4801) );
  NANDN U403 ( .A(n2235), .B(n2541), .Z(n158) );
  XNOR U404 ( .A(n2375), .B(n158), .Z(out[1371]) );
  AND U405 ( .A(n4753), .B(n4357), .Z(n159) );
  XNOR U406 ( .A(n4579), .B(n159), .Z(out[712]) );
  NANDN U407 ( .A(n4456), .B(n4877), .Z(n160) );
  XNOR U408 ( .A(n4653), .B(n160), .Z(out[740]) );
  NANDN U409 ( .A(n4462), .B(n4885), .Z(n161) );
  XNOR U410 ( .A(n4663), .B(n161), .Z(out[742]) );
  NANDN U411 ( .A(n2212), .B(n2496), .Z(n162) );
  XNOR U412 ( .A(n2353), .B(n162), .Z(out[1360]) );
  ANDN U413 ( .B(n4683), .A(n4942), .Z(n163) );
  XNOR U414 ( .A(n4943), .B(n163), .Z(out[884]) );
  ANDN U415 ( .B(n5013), .A(n1607), .Z(n164) );
  XNOR U416 ( .A(n1818), .B(n164), .Z(out[1091]) );
  ANDN U417 ( .B(n5029), .A(n1623), .Z(n165) );
  XNOR U418 ( .A(n1829), .B(n165), .Z(out[1095]) );
  ANDN U419 ( .B(n5033), .A(n1628), .Z(n166) );
  XNOR U420 ( .A(n1831), .B(n166), .Z(out[1096]) );
  ANDN U421 ( .B(n5061), .A(n1652), .Z(n167) );
  XNOR U422 ( .A(n1845), .B(n167), .Z(out[1102]) );
  AND U423 ( .A(n5074), .B(n1669), .Z(n168) );
  XNOR U424 ( .A(n1853), .B(n168), .Z(out[1106]) );
  ANDN U425 ( .B(n5078), .A(n1673), .Z(n169) );
  XNOR U426 ( .A(n1855), .B(n169), .Z(out[1107]) );
  ANDN U427 ( .B(n5094), .A(n1689), .Z(n170) );
  XNOR U428 ( .A(n1863), .B(n170), .Z(out[1111]) );
  NAND U429 ( .A(n3839), .B(n3418), .Z(n171) );
  XNOR U430 ( .A(n3417), .B(n171), .Z(out[435]) );
  ANDN U431 ( .B(n5110), .A(n1710), .Z(n172) );
  XNOR U432 ( .A(n1875), .B(n172), .Z(out[1116]) );
  ANDN U433 ( .B(n5113), .A(n1714), .Z(n173) );
  XNOR U434 ( .A(n1877), .B(n173), .Z(out[1117]) );
  ANDN U435 ( .B(n3863), .A(n3438), .Z(n174) );
  XNOR U436 ( .A(n3592), .B(n174), .Z(out[440]) );
  ANDN U437 ( .B(n2668), .A(n2299), .Z(n175) );
  XNOR U438 ( .A(n2417), .B(n175), .Z(out[1401]) );
  AND U439 ( .A(n3887), .B(n3460), .Z(n176) );
  XNOR U440 ( .A(n3606), .B(n176), .Z(out[446]) );
  ANDN U441 ( .B(n3891), .A(n3463), .Z(n177) );
  XNOR U442 ( .A(n3608), .B(n177), .Z(out[447]) );
  ANDN U443 ( .B(n3613), .A(n3259), .Z(n178) );
  XNOR U444 ( .A(n3465), .B(n178), .Z(out[384]) );
  AND U445 ( .A(n2631), .B(n2406), .Z(n179) );
  XNOR U446 ( .A(n2632), .B(n179), .Z(out[1521]) );
  AND U447 ( .A(n2635), .B(n2407), .Z(n180) );
  XNOR U448 ( .A(n2636), .B(n180), .Z(out[1522]) );
  AND U449 ( .A(n2657), .B(n2415), .Z(n181) );
  XNOR U450 ( .A(n2658), .B(n181), .Z(out[1527]) );
  NOR U451 ( .A(n4704), .B(n4551), .Z(n182) );
  XNOR U452 ( .A(n4986), .B(n182), .Z(out[830]) );
  NOR U453 ( .A(n4707), .B(n4553), .Z(n183) );
  XNOR U454 ( .A(n4990), .B(n183), .Z(out[831]) );
  NOR U455 ( .A(n4554), .B(n4334), .Z(n184) );
  XNOR U456 ( .A(n4710), .B(n184), .Z(out[768]) );
  NOR U457 ( .A(n4595), .B(n4385), .Z(n185) );
  XNOR U458 ( .A(n4787), .B(n185), .Z(out[784]) );
  ANDN U459 ( .B(n1988), .A(n1581), .Z(n186) );
  XNOR U460 ( .A(n1800), .B(n186), .Z(out[1084]) );
  ANDN U461 ( .B(n1992), .A(n1585), .Z(n187) );
  XNOR U462 ( .A(n1802), .B(n187), .Z(out[1085]) );
  NAND U463 ( .A(n2890), .B(n4404), .Z(n188) );
  XNOR U464 ( .A(n2889), .B(n188), .Z(out[206]) );
  NAND U465 ( .A(n2893), .B(n4438), .Z(n189) );
  XNOR U466 ( .A(n2892), .B(n189), .Z(out[207]) );
  NANDN U467 ( .A(n2929), .B(n4777), .Z(n190) );
  XNOR U468 ( .A(n2928), .B(n190), .Z(out[218]) );
  ANDN U469 ( .B(n1912), .A(n1507), .Z(n191) );
  XNOR U470 ( .A(n1761), .B(n191), .Z(out[1066]) );
  NANDN U471 ( .A(n1511), .B(n1916), .Z(n192) );
  XNOR U472 ( .A(n1763), .B(n192), .Z(out[1067]) );
  ANDN U473 ( .B(n1922), .A(n1515), .Z(n193) );
  XNOR U474 ( .A(n1764), .B(n193), .Z(out[1068]) );
  ANDN U475 ( .B(n1926), .A(n1519), .Z(n194) );
  XNOR U476 ( .A(n1766), .B(n194), .Z(out[1069]) );
  ANDN U477 ( .B(n1930), .A(n1523), .Z(n195) );
  XNOR U478 ( .A(n1768), .B(n195), .Z(out[1070]) );
  ANDN U479 ( .B(n1934), .A(n1527), .Z(n196) );
  XNOR U480 ( .A(n1770), .B(n196), .Z(out[1071]) );
  ANDN U481 ( .B(n1938), .A(n1531), .Z(n197) );
  XNOR U482 ( .A(n1774), .B(n197), .Z(out[1072]) );
  ANDN U483 ( .B(n1942), .A(n1535), .Z(n198) );
  XNOR U484 ( .A(n1776), .B(n198), .Z(out[1073]) );
  ANDN U485 ( .B(n2470), .A(n2469), .Z(n199) );
  XNOR U486 ( .A(n2468), .B(n199), .Z(out[1545]) );
  OR U487 ( .A(n5066), .B(n5067), .Z(n200) );
  XNOR U488 ( .A(n5068), .B(n200), .Z(out[976]) );
  OR U489 ( .A(n5069), .B(n5070), .Z(n201) );
  XNOR U490 ( .A(n5071), .B(n201), .Z(out[977]) );
  NAND U491 ( .A(n3600), .B(n3869), .Z(n202) );
  XNOR U492 ( .A(n3868), .B(n202), .Z(out[570]) );
  NAND U493 ( .A(n3601), .B(n3873), .Z(n203) );
  XNOR U494 ( .A(n3872), .B(n203), .Z(out[571]) );
  OR U495 ( .A(n5089), .B(n5090), .Z(n204) );
  XNOR U496 ( .A(n5091), .B(n204), .Z(out[982]) );
  OR U497 ( .A(n5095), .B(n5096), .Z(n205) );
  XNOR U498 ( .A(n5097), .B(n205), .Z(out[984]) );
  OR U499 ( .A(n5098), .B(n5099), .Z(n206) );
  XNOR U500 ( .A(n5100), .B(n206), .Z(out[985]) );
  OR U501 ( .A(n5101), .B(n5102), .Z(n207) );
  XNOR U502 ( .A(n5103), .B(n207), .Z(out[986]) );
  OR U503 ( .A(n5104), .B(n5105), .Z(n208) );
  XNOR U504 ( .A(n5106), .B(n208), .Z(out[987]) );
  NANDN U505 ( .A(n4412), .B(n4825), .Z(n209) );
  XNOR U506 ( .A(n4618), .B(n209), .Z(out[728]) );
  NAND U507 ( .A(n3473), .B(n3631), .Z(n210) );
  XNOR U508 ( .A(n3630), .B(n210), .Z(out[516]) );
  NANDN U509 ( .A(n4415), .B(n4829), .Z(n211) );
  XNOR U510 ( .A(n4621), .B(n211), .Z(out[729]) );
  NANDN U511 ( .A(n3635), .B(n3474), .Z(n212) );
  XNOR U512 ( .A(n3634), .B(n212), .Z(out[517]) );
  OR U513 ( .A(n5118), .B(n5119), .Z(n213) );
  XNOR U514 ( .A(n5120), .B(n213), .Z(out[990]) );
  ANDN U515 ( .B(n4833), .A(n4418), .Z(n214) );
  XNOR U516 ( .A(n4624), .B(n214), .Z(out[730]) );
  NANDN U517 ( .A(n3639), .B(n3475), .Z(n215) );
  XNOR U518 ( .A(n3638), .B(n215), .Z(out[518]) );
  NANDN U519 ( .A(n3643), .B(n3476), .Z(n216) );
  XNOR U520 ( .A(n3642), .B(n216), .Z(out[519]) );
  NAND U521 ( .A(n3481), .B(n3647), .Z(n217) );
  XNOR U522 ( .A(n3646), .B(n217), .Z(out[520]) );
  NANDN U523 ( .A(n4427), .B(n4845), .Z(n218) );
  XNOR U524 ( .A(n4634), .B(n218), .Z(out[733]) );
  NANDN U525 ( .A(n4433), .B(n4853), .Z(n219) );
  XNOR U526 ( .A(n4640), .B(n219), .Z(out[735]) );
  NANDN U527 ( .A(n4447), .B(n4861), .Z(n220) );
  XNOR U528 ( .A(n4644), .B(n220), .Z(out[737]) );
  NANDN U529 ( .A(n4453), .B(n4873), .Z(n221) );
  XNOR U530 ( .A(n4650), .B(n221), .Z(out[739]) );
  ANDN U531 ( .B(n3498), .A(n3686), .Z(n222) );
  XNOR U532 ( .A(n3687), .B(n222), .Z(out[529]) );
  ANDN U533 ( .B(n3503), .A(n3690), .Z(n223) );
  XNOR U534 ( .A(n3691), .B(n223), .Z(out[530]) );
  ANDN U535 ( .B(n3504), .A(n3694), .Z(n224) );
  XNOR U536 ( .A(n3695), .B(n224), .Z(out[531]) );
  ANDN U537 ( .B(n3505), .A(n3698), .Z(n225) );
  XNOR U538 ( .A(n3699), .B(n225), .Z(out[532]) );
  ANDN U539 ( .B(n3507), .A(n3706), .Z(n226) );
  XNOR U540 ( .A(n3707), .B(n226), .Z(out[534]) );
  ANDN U541 ( .B(n3508), .A(n3710), .Z(n227) );
  XNOR U542 ( .A(n3711), .B(n227), .Z(out[535]) );
  ANDN U543 ( .B(n3509), .A(n3720), .Z(n228) );
  XNOR U544 ( .A(n3721), .B(n228), .Z(out[536]) );
  ANDN U545 ( .B(n3513), .A(n3732), .Z(n229) );
  XNOR U546 ( .A(n3733), .B(n229), .Z(out[539]) );
  XNOR U547 ( .A(in[1168]), .B(n932), .Z(n230) );
  XNOR U548 ( .A(in[545]), .B(n1174), .Z(n231) );
  XOR U549 ( .A(in[1469]), .B(in[509]), .Z(n233) );
  XNOR U550 ( .A(in[829]), .B(in[189]), .Z(n232) );
  XNOR U551 ( .A(n233), .B(n232), .Z(n234) );
  XNOR U552 ( .A(in[1149]), .B(n234), .Z(n1103) );
  XOR U553 ( .A(in[1598]), .B(in[638]), .Z(n236) );
  XNOR U554 ( .A(in[958]), .B(in[318]), .Z(n235) );
  XNOR U555 ( .A(n236), .B(n235), .Z(n237) );
  XNOR U556 ( .A(in[1278]), .B(n237), .Z(n1672) );
  XNOR U557 ( .A(n1103), .B(n1672), .Z(n3286) );
  XOR U558 ( .A(in[254]), .B(n3286), .Z(n3936) );
  XOR U559 ( .A(in[1345]), .B(in[65]), .Z(n239) );
  XNOR U560 ( .A(in[1025]), .B(in[385]), .Z(n238) );
  XNOR U561 ( .A(n239), .B(n238), .Z(n240) );
  XNOR U562 ( .A(in[705]), .B(n240), .Z(n1680) );
  XOR U563 ( .A(in[1474]), .B(in[514]), .Z(n242) );
  XNOR U564 ( .A(in[834]), .B(in[194]), .Z(n241) );
  XNOR U565 ( .A(n242), .B(n241), .Z(n243) );
  XOR U566 ( .A(in[1154]), .B(n243), .Z(n1405) );
  XOR U567 ( .A(in[1410]), .B(n3169), .Z(n3937) );
  XOR U568 ( .A(in[137]), .B(in[457]), .Z(n245) );
  XNOR U569 ( .A(in[777]), .B(in[1417]), .Z(n244) );
  XNOR U570 ( .A(n245), .B(n244), .Z(n246) );
  XNOR U571 ( .A(in[1097]), .B(n246), .Z(n1362) );
  XOR U572 ( .A(in[328]), .B(in[8]), .Z(n248) );
  XNOR U573 ( .A(in[968]), .B(in[648]), .Z(n247) );
  XNOR U574 ( .A(n248), .B(n247), .Z(n249) );
  XNOR U575 ( .A(in[1288]), .B(n249), .Z(n1418) );
  XOR U576 ( .A(n1362), .B(n1418), .Z(n4449) );
  XNOR U577 ( .A(in[1033]), .B(n4449), .Z(n2854) );
  OR U578 ( .A(n3937), .B(n2854), .Z(n250) );
  XOR U579 ( .A(n3936), .B(n250), .Z(out[0]) );
  XOR U580 ( .A(in[1386]), .B(in[106]), .Z(n252) );
  XNOR U581 ( .A(in[1066]), .B(in[746]), .Z(n251) );
  XNOR U582 ( .A(n252), .B(n251), .Z(n253) );
  XNOR U583 ( .A(in[426]), .B(n253), .Z(n706) );
  XOR U584 ( .A(in[1515]), .B(in[555]), .Z(n255) );
  XNOR U585 ( .A(in[875]), .B(in[235]), .Z(n254) );
  XNOR U586 ( .A(n255), .B(n254), .Z(n256) );
  XNOR U587 ( .A(in[1195]), .B(n256), .Z(n1526) );
  XOR U588 ( .A(n706), .B(n1526), .Z(n4107) );
  XOR U589 ( .A(in[171]), .B(n4107), .Z(n1497) );
  XOR U590 ( .A(in[971]), .B(in[1291]), .Z(n258) );
  XNOR U591 ( .A(in[11]), .B(in[331]), .Z(n257) );
  XNOR U592 ( .A(n258), .B(n257), .Z(n259) );
  XNOR U593 ( .A(in[651]), .B(n259), .Z(n1427) );
  XOR U594 ( .A(in[140]), .B(in[460]), .Z(n261) );
  XNOR U595 ( .A(in[1100]), .B(in[1420]), .Z(n260) );
  XNOR U596 ( .A(n261), .B(n260), .Z(n262) );
  XOR U597 ( .A(in[780]), .B(n262), .Z(n1384) );
  XNOR U598 ( .A(in[1356]), .B(n4458), .Z(n1904) );
  XOR U599 ( .A(in[1364]), .B(in[724]), .Z(n264) );
  XNOR U600 ( .A(in[84]), .B(in[404]), .Z(n263) );
  XNOR U601 ( .A(n264), .B(n263), .Z(n265) );
  XNOR U602 ( .A(in[1044]), .B(n265), .Z(n1008) );
  XOR U603 ( .A(in[1555]), .B(in[595]), .Z(n267) );
  XNOR U604 ( .A(in[915]), .B(in[275]), .Z(n266) );
  XNOR U605 ( .A(n267), .B(n266), .Z(n268) );
  XNOR U606 ( .A(in[1235]), .B(n268), .Z(n720) );
  XOR U607 ( .A(n1008), .B(n720), .Z(n4246) );
  XOR U608 ( .A(in[980]), .B(n4246), .Z(n1901) );
  NANDN U609 ( .A(n1904), .B(n1901), .Z(n269) );
  XNOR U610 ( .A(n1497), .B(n269), .Z(out[1000]) );
  XOR U611 ( .A(in[1387]), .B(in[107]), .Z(n271) );
  XNOR U612 ( .A(in[1067]), .B(in[747]), .Z(n270) );
  XNOR U613 ( .A(n271), .B(n270), .Z(n272) );
  XNOR U614 ( .A(in[427]), .B(n272), .Z(n717) );
  XOR U615 ( .A(in[1516]), .B(in[556]), .Z(n274) );
  XNOR U616 ( .A(in[876]), .B(in[236]), .Z(n273) );
  XNOR U617 ( .A(n274), .B(n273), .Z(n275) );
  XNOR U618 ( .A(in[1196]), .B(n275), .Z(n1530) );
  XOR U619 ( .A(n717), .B(n1530), .Z(n4115) );
  XOR U620 ( .A(in[172]), .B(n4115), .Z(n1501) );
  XOR U621 ( .A(in[972]), .B(in[12]), .Z(n277) );
  XNOR U622 ( .A(in[1292]), .B(in[332]), .Z(n276) );
  XNOR U623 ( .A(n277), .B(n276), .Z(n278) );
  XNOR U624 ( .A(in[652]), .B(n278), .Z(n1429) );
  XOR U625 ( .A(in[141]), .B(in[461]), .Z(n280) );
  XNOR U626 ( .A(in[1101]), .B(in[1421]), .Z(n279) );
  XNOR U627 ( .A(n280), .B(n279), .Z(n281) );
  XOR U628 ( .A(in[781]), .B(n281), .Z(n1388) );
  XNOR U629 ( .A(in[1357]), .B(n4461), .Z(n1908) );
  XOR U630 ( .A(in[1365]), .B(in[725]), .Z(n283) );
  XNOR U631 ( .A(in[85]), .B(in[405]), .Z(n282) );
  XNOR U632 ( .A(n283), .B(n282), .Z(n284) );
  XNOR U633 ( .A(in[1045]), .B(n284), .Z(n1021) );
  XOR U634 ( .A(in[1556]), .B(in[596]), .Z(n286) );
  XNOR U635 ( .A(in[916]), .B(in[276]), .Z(n285) );
  XNOR U636 ( .A(n286), .B(n285), .Z(n287) );
  XNOR U637 ( .A(in[1236]), .B(n287), .Z(n735) );
  XOR U638 ( .A(n1021), .B(n735), .Z(n4249) );
  XOR U639 ( .A(in[981]), .B(n4249), .Z(n1905) );
  NANDN U640 ( .A(n1908), .B(n1905), .Z(n288) );
  XNOR U641 ( .A(n1501), .B(n288), .Z(out[1001]) );
  XOR U642 ( .A(in[1388]), .B(in[108]), .Z(n290) );
  XNOR U643 ( .A(in[1068]), .B(in[748]), .Z(n289) );
  XNOR U644 ( .A(n290), .B(n289), .Z(n291) );
  XNOR U645 ( .A(in[428]), .B(n291), .Z(n1594) );
  XOR U646 ( .A(in[1517]), .B(in[557]), .Z(n293) );
  XNOR U647 ( .A(in[877]), .B(in[237]), .Z(n292) );
  XNOR U648 ( .A(n293), .B(n292), .Z(n294) );
  XNOR U649 ( .A(in[1197]), .B(n294), .Z(n1534) );
  XOR U650 ( .A(n1594), .B(n1534), .Z(n1367) );
  XOR U651 ( .A(in[173]), .B(n1367), .Z(n1507) );
  XOR U652 ( .A(in[973]), .B(in[13]), .Z(n296) );
  XNOR U653 ( .A(in[1293]), .B(in[333]), .Z(n295) );
  XNOR U654 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U655 ( .A(in[653]), .B(n297), .Z(n1431) );
  XOR U656 ( .A(in[142]), .B(in[1422]), .Z(n299) );
  XNOR U657 ( .A(in[1102]), .B(in[782]), .Z(n298) );
  XNOR U658 ( .A(n299), .B(n298), .Z(n300) );
  XOR U659 ( .A(in[462]), .B(n300), .Z(n1392) );
  XNOR U660 ( .A(in[1358]), .B(n4464), .Z(n1912) );
  XOR U661 ( .A(in[1366]), .B(in[726]), .Z(n302) );
  XNOR U662 ( .A(in[86]), .B(in[406]), .Z(n301) );
  XNOR U663 ( .A(n302), .B(n301), .Z(n303) );
  XNOR U664 ( .A(in[1046]), .B(n303), .Z(n1034) );
  XOR U665 ( .A(in[1557]), .B(in[597]), .Z(n305) );
  XNOR U666 ( .A(in[917]), .B(in[277]), .Z(n304) );
  XNOR U667 ( .A(n305), .B(n304), .Z(n306) );
  XNOR U668 ( .A(in[1237]), .B(n306), .Z(n750) );
  XOR U669 ( .A(n1034), .B(n750), .Z(n4250) );
  XOR U670 ( .A(in[982]), .B(n4250), .Z(n1909) );
  NANDN U671 ( .A(n1912), .B(n1909), .Z(n307) );
  XNOR U672 ( .A(n1507), .B(n307), .Z(out[1002]) );
  XOR U673 ( .A(in[1389]), .B(in[109]), .Z(n309) );
  XNOR U674 ( .A(in[1069]), .B(in[749]), .Z(n308) );
  XNOR U675 ( .A(n309), .B(n308), .Z(n310) );
  XNOR U676 ( .A(in[429]), .B(n310), .Z(n1598) );
  XOR U677 ( .A(in[1518]), .B(in[558]), .Z(n312) );
  XNOR U678 ( .A(in[878]), .B(in[238]), .Z(n311) );
  XNOR U679 ( .A(n312), .B(n311), .Z(n313) );
  XNOR U680 ( .A(in[1198]), .B(n313), .Z(n1538) );
  XOR U681 ( .A(n1598), .B(n1538), .Z(n1407) );
  XOR U682 ( .A(in[174]), .B(n1407), .Z(n1511) );
  XOR U683 ( .A(in[974]), .B(in[14]), .Z(n315) );
  XNOR U684 ( .A(in[1294]), .B(in[334]), .Z(n314) );
  XNOR U685 ( .A(n315), .B(n314), .Z(n316) );
  XNOR U686 ( .A(in[654]), .B(n316), .Z(n1433) );
  XOR U687 ( .A(in[143]), .B(in[1423]), .Z(n318) );
  XNOR U688 ( .A(in[1103]), .B(in[783]), .Z(n317) );
  XNOR U689 ( .A(n318), .B(n317), .Z(n319) );
  XOR U690 ( .A(in[463]), .B(n319), .Z(n1396) );
  XNOR U691 ( .A(in[1359]), .B(n4467), .Z(n1916) );
  XOR U692 ( .A(in[1367]), .B(in[727]), .Z(n321) );
  XNOR U693 ( .A(in[87]), .B(in[407]), .Z(n320) );
  XNOR U694 ( .A(n321), .B(n320), .Z(n322) );
  XNOR U695 ( .A(in[1047]), .B(n322), .Z(n1047) );
  XOR U696 ( .A(in[1558]), .B(in[598]), .Z(n324) );
  XNOR U697 ( .A(in[918]), .B(in[278]), .Z(n323) );
  XNOR U698 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U699 ( .A(in[1238]), .B(n325), .Z(n765) );
  XOR U700 ( .A(n1047), .B(n765), .Z(n4251) );
  XOR U701 ( .A(in[983]), .B(n4251), .Z(n1913) );
  NANDN U702 ( .A(n1916), .B(n1913), .Z(n326) );
  XNOR U703 ( .A(n1511), .B(n326), .Z(out[1003]) );
  XOR U704 ( .A(in[1390]), .B(in[110]), .Z(n328) );
  XNOR U705 ( .A(in[1070]), .B(in[750]), .Z(n327) );
  XNOR U706 ( .A(n328), .B(n327), .Z(n329) );
  XNOR U707 ( .A(in[430]), .B(n329), .Z(n1602) );
  XOR U708 ( .A(in[1519]), .B(in[559]), .Z(n331) );
  XNOR U709 ( .A(in[879]), .B(in[239]), .Z(n330) );
  XNOR U710 ( .A(n331), .B(n330), .Z(n332) );
  XNOR U711 ( .A(in[1199]), .B(n332), .Z(n1542) );
  XOR U712 ( .A(n1602), .B(n1542), .Z(n1419) );
  XOR U713 ( .A(in[175]), .B(n1419), .Z(n1515) );
  XOR U714 ( .A(in[144]), .B(in[1424]), .Z(n334) );
  XNOR U715 ( .A(in[1104]), .B(in[784]), .Z(n333) );
  XNOR U716 ( .A(n334), .B(n333), .Z(n335) );
  XNOR U717 ( .A(in[464]), .B(n335), .Z(n1400) );
  XOR U718 ( .A(in[975]), .B(in[15]), .Z(n337) );
  XNOR U719 ( .A(in[1295]), .B(in[335]), .Z(n336) );
  XNOR U720 ( .A(n337), .B(n336), .Z(n338) );
  XOR U721 ( .A(in[655]), .B(n338), .Z(n1435) );
  XNOR U722 ( .A(in[1360]), .B(n4470), .Z(n1922) );
  XOR U723 ( .A(in[1368]), .B(in[728]), .Z(n340) );
  XNOR U724 ( .A(in[88]), .B(in[408]), .Z(n339) );
  XNOR U725 ( .A(n340), .B(n339), .Z(n341) );
  XNOR U726 ( .A(in[1048]), .B(n341), .Z(n1060) );
  XOR U727 ( .A(in[1559]), .B(in[599]), .Z(n343) );
  XNOR U728 ( .A(in[919]), .B(in[279]), .Z(n342) );
  XNOR U729 ( .A(n343), .B(n342), .Z(n344) );
  XNOR U730 ( .A(in[1239]), .B(n344), .Z(n780) );
  XOR U731 ( .A(n1060), .B(n780), .Z(n4252) );
  XOR U732 ( .A(in[984]), .B(n4252), .Z(n1919) );
  NANDN U733 ( .A(n1922), .B(n1919), .Z(n345) );
  XNOR U734 ( .A(n1515), .B(n345), .Z(out[1004]) );
  XOR U735 ( .A(in[1391]), .B(in[111]), .Z(n347) );
  XNOR U736 ( .A(in[1071]), .B(in[751]), .Z(n346) );
  XNOR U737 ( .A(n347), .B(n346), .Z(n348) );
  XNOR U738 ( .A(in[431]), .B(n348), .Z(n1606) );
  XOR U739 ( .A(in[1520]), .B(in[560]), .Z(n350) );
  XNOR U740 ( .A(in[880]), .B(in[240]), .Z(n349) );
  XNOR U741 ( .A(n350), .B(n349), .Z(n351) );
  XNOR U742 ( .A(in[1200]), .B(n351), .Z(n1548) );
  XOR U743 ( .A(n1606), .B(n1548), .Z(n1441) );
  XOR U744 ( .A(in[176]), .B(n1441), .Z(n1519) );
  XOR U745 ( .A(in[145]), .B(in[1425]), .Z(n353) );
  XNOR U746 ( .A(in[1105]), .B(in[785]), .Z(n352) );
  XNOR U747 ( .A(n353), .B(n352), .Z(n354) );
  XNOR U748 ( .A(in[465]), .B(n354), .Z(n1404) );
  XOR U749 ( .A(in[976]), .B(in[16]), .Z(n356) );
  XNOR U750 ( .A(in[1296]), .B(in[336]), .Z(n355) );
  XNOR U751 ( .A(n356), .B(n355), .Z(n357) );
  XOR U752 ( .A(in[656]), .B(n357), .Z(n1437) );
  XNOR U753 ( .A(in[1361]), .B(n4477), .Z(n1926) );
  XOR U754 ( .A(in[1369]), .B(in[729]), .Z(n359) );
  XNOR U755 ( .A(in[89]), .B(in[409]), .Z(n358) );
  XNOR U756 ( .A(n359), .B(n358), .Z(n360) );
  XNOR U757 ( .A(in[1049]), .B(n360), .Z(n1073) );
  XOR U758 ( .A(in[1560]), .B(in[600]), .Z(n362) );
  XNOR U759 ( .A(in[920]), .B(in[280]), .Z(n361) );
  XNOR U760 ( .A(n362), .B(n361), .Z(n363) );
  XNOR U761 ( .A(in[1240]), .B(n363), .Z(n795) );
  XOR U762 ( .A(n1073), .B(n795), .Z(n4253) );
  XOR U763 ( .A(in[985]), .B(n4253), .Z(n1923) );
  NANDN U764 ( .A(n1926), .B(n1923), .Z(n364) );
  XNOR U765 ( .A(n1519), .B(n364), .Z(out[1005]) );
  XOR U766 ( .A(in[1392]), .B(in[112]), .Z(n366) );
  XNOR U767 ( .A(in[1072]), .B(in[752]), .Z(n365) );
  XNOR U768 ( .A(n366), .B(n365), .Z(n367) );
  XNOR U769 ( .A(in[432]), .B(n367), .Z(n1610) );
  XOR U770 ( .A(in[1521]), .B(in[561]), .Z(n369) );
  XNOR U771 ( .A(in[881]), .B(in[241]), .Z(n368) );
  XNOR U772 ( .A(n369), .B(n368), .Z(n370) );
  XNOR U773 ( .A(in[1201]), .B(n370), .Z(n1552) );
  XOR U774 ( .A(n1610), .B(n1552), .Z(n1469) );
  XOR U775 ( .A(in[177]), .B(n1469), .Z(n1523) );
  XOR U776 ( .A(in[1426]), .B(in[466]), .Z(n372) );
  XNOR U777 ( .A(in[786]), .B(in[146]), .Z(n371) );
  XNOR U778 ( .A(n372), .B(n371), .Z(n373) );
  XNOR U779 ( .A(in[1106]), .B(n373), .Z(n719) );
  XOR U780 ( .A(in[17]), .B(in[657]), .Z(n375) );
  XNOR U781 ( .A(in[977]), .B(in[337]), .Z(n374) );
  XNOR U782 ( .A(n375), .B(n374), .Z(n376) );
  XOR U783 ( .A(in[1297]), .B(n376), .Z(n1438) );
  XNOR U784 ( .A(n4480), .B(in[1362]), .Z(n1930) );
  XOR U785 ( .A(in[1370]), .B(in[730]), .Z(n378) );
  XNOR U786 ( .A(in[90]), .B(in[410]), .Z(n377) );
  XNOR U787 ( .A(n378), .B(n377), .Z(n379) );
  XNOR U788 ( .A(in[1050]), .B(n379), .Z(n1088) );
  XOR U789 ( .A(in[1561]), .B(in[601]), .Z(n381) );
  XNOR U790 ( .A(in[921]), .B(in[281]), .Z(n380) );
  XNOR U791 ( .A(n381), .B(n380), .Z(n382) );
  XNOR U792 ( .A(in[1241]), .B(n382), .Z(n821) );
  XOR U793 ( .A(n1088), .B(n821), .Z(n4254) );
  XOR U794 ( .A(in[986]), .B(n4254), .Z(n1927) );
  NANDN U795 ( .A(n1930), .B(n1927), .Z(n383) );
  XNOR U796 ( .A(n1523), .B(n383), .Z(out[1006]) );
  XOR U797 ( .A(in[1393]), .B(in[113]), .Z(n385) );
  XNOR U798 ( .A(in[1073]), .B(in[753]), .Z(n384) );
  XNOR U799 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U800 ( .A(in[433]), .B(n386), .Z(n1614) );
  XOR U801 ( .A(in[1522]), .B(in[562]), .Z(n388) );
  XNOR U802 ( .A(in[882]), .B(in[242]), .Z(n387) );
  XNOR U803 ( .A(n388), .B(n387), .Z(n389) );
  XNOR U804 ( .A(in[1202]), .B(n389), .Z(n1556) );
  XOR U805 ( .A(n1614), .B(n1556), .Z(n1503) );
  XOR U806 ( .A(in[178]), .B(n1503), .Z(n1527) );
  XOR U807 ( .A(in[978]), .B(in[18]), .Z(n391) );
  XNOR U808 ( .A(in[1298]), .B(in[338]), .Z(n390) );
  XNOR U809 ( .A(n391), .B(n390), .Z(n392) );
  XNOR U810 ( .A(in[658]), .B(n392), .Z(n1440) );
  XOR U811 ( .A(in[147]), .B(in[1427]), .Z(n394) );
  XNOR U812 ( .A(in[1107]), .B(in[787]), .Z(n393) );
  XNOR U813 ( .A(n394), .B(n393), .Z(n395) );
  XOR U814 ( .A(in[467]), .B(n395), .Z(n734) );
  XNOR U815 ( .A(in[1363]), .B(n4483), .Z(n1934) );
  XOR U816 ( .A(in[1371]), .B(in[731]), .Z(n397) );
  XNOR U817 ( .A(in[91]), .B(in[411]), .Z(n396) );
  XNOR U818 ( .A(n397), .B(n396), .Z(n398) );
  XNOR U819 ( .A(in[1051]), .B(n398), .Z(n1101) );
  XOR U820 ( .A(in[1562]), .B(in[602]), .Z(n400) );
  XNOR U821 ( .A(in[922]), .B(in[282]), .Z(n399) );
  XNOR U822 ( .A(n400), .B(n399), .Z(n401) );
  XNOR U823 ( .A(in[1242]), .B(n401), .Z(n836) );
  XOR U824 ( .A(n1101), .B(n836), .Z(n4255) );
  XOR U825 ( .A(in[987]), .B(n4255), .Z(n1931) );
  NANDN U826 ( .A(n1934), .B(n1931), .Z(n402) );
  XNOR U827 ( .A(n1527), .B(n402), .Z(out[1007]) );
  XOR U828 ( .A(in[1394]), .B(in[114]), .Z(n404) );
  XNOR U829 ( .A(in[1074]), .B(in[754]), .Z(n403) );
  XNOR U830 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U831 ( .A(in[434]), .B(n405), .Z(n1618) );
  XOR U832 ( .A(in[1523]), .B(in[563]), .Z(n407) );
  XNOR U833 ( .A(in[883]), .B(in[243]), .Z(n406) );
  XNOR U834 ( .A(n407), .B(n406), .Z(n408) );
  XNOR U835 ( .A(in[1203]), .B(n408), .Z(n1560) );
  XOR U836 ( .A(n1618), .B(n1560), .Z(n1545) );
  XOR U837 ( .A(in[179]), .B(n1545), .Z(n1531) );
  XOR U838 ( .A(in[148]), .B(in[1428]), .Z(n410) );
  XNOR U839 ( .A(in[1108]), .B(in[788]), .Z(n409) );
  XNOR U840 ( .A(n410), .B(n409), .Z(n411) );
  XNOR U841 ( .A(in[468]), .B(n411), .Z(n749) );
  XOR U842 ( .A(in[979]), .B(in[19]), .Z(n413) );
  XNOR U843 ( .A(in[1299]), .B(in[339]), .Z(n412) );
  XNOR U844 ( .A(n413), .B(n412), .Z(n414) );
  XOR U845 ( .A(in[659]), .B(n414), .Z(n1444) );
  XNOR U846 ( .A(in[1364]), .B(n4486), .Z(n1938) );
  XOR U847 ( .A(in[1372]), .B(in[732]), .Z(n416) );
  XNOR U848 ( .A(in[92]), .B(in[412]), .Z(n415) );
  XNOR U849 ( .A(n416), .B(n415), .Z(n417) );
  XNOR U850 ( .A(in[1052]), .B(n417), .Z(n1121) );
  XOR U851 ( .A(in[1563]), .B(in[603]), .Z(n419) );
  XNOR U852 ( .A(in[923]), .B(in[283]), .Z(n418) );
  XNOR U853 ( .A(n419), .B(n418), .Z(n420) );
  XNOR U854 ( .A(in[1243]), .B(n420), .Z(n851) );
  XOR U855 ( .A(n1121), .B(n851), .Z(n4258) );
  XOR U856 ( .A(in[988]), .B(n4258), .Z(n1935) );
  NANDN U857 ( .A(n1938), .B(n1935), .Z(n421) );
  XNOR U858 ( .A(n1531), .B(n421), .Z(out[1008]) );
  XOR U859 ( .A(in[1395]), .B(in[115]), .Z(n423) );
  XNOR U860 ( .A(in[1075]), .B(in[755]), .Z(n422) );
  XNOR U861 ( .A(n423), .B(n422), .Z(n424) );
  XNOR U862 ( .A(in[435]), .B(n424), .Z(n1622) );
  XOR U863 ( .A(in[1524]), .B(in[564]), .Z(n426) );
  XNOR U864 ( .A(in[884]), .B(in[244]), .Z(n425) );
  XNOR U865 ( .A(n426), .B(n425), .Z(n427) );
  XNOR U866 ( .A(in[1204]), .B(n427), .Z(n1564) );
  XOR U867 ( .A(n1622), .B(n1564), .Z(n1587) );
  XOR U868 ( .A(in[180]), .B(n1587), .Z(n1535) );
  XOR U869 ( .A(in[149]), .B(in[1429]), .Z(n429) );
  XNOR U870 ( .A(in[1109]), .B(in[789]), .Z(n428) );
  XNOR U871 ( .A(n429), .B(n428), .Z(n430) );
  XNOR U872 ( .A(in[469]), .B(n430), .Z(n764) );
  XOR U873 ( .A(in[340]), .B(in[660]), .Z(n432) );
  XNOR U874 ( .A(in[20]), .B(in[1300]), .Z(n431) );
  XNOR U875 ( .A(n432), .B(n431), .Z(n433) );
  XOR U876 ( .A(in[980]), .B(n433), .Z(n1446) );
  XNOR U877 ( .A(in[1365]), .B(n4489), .Z(n1942) );
  XOR U878 ( .A(in[1373]), .B(in[733]), .Z(n435) );
  XNOR U879 ( .A(in[93]), .B(in[413]), .Z(n434) );
  XNOR U880 ( .A(n435), .B(n434), .Z(n436) );
  XNOR U881 ( .A(in[1053]), .B(n436), .Z(n1134) );
  XOR U882 ( .A(in[1564]), .B(in[604]), .Z(n438) );
  XNOR U883 ( .A(in[924]), .B(in[284]), .Z(n437) );
  XNOR U884 ( .A(n438), .B(n437), .Z(n439) );
  XNOR U885 ( .A(in[1244]), .B(n439), .Z(n866) );
  XOR U886 ( .A(n1134), .B(n866), .Z(n4259) );
  XOR U887 ( .A(in[989]), .B(n4259), .Z(n1939) );
  NANDN U888 ( .A(n1942), .B(n1939), .Z(n440) );
  XNOR U889 ( .A(n1535), .B(n440), .Z(out[1009]) );
  XOR U890 ( .A(in[1339]), .B(in[59]), .Z(n442) );
  XNOR U891 ( .A(in[699]), .B(in[379]), .Z(n441) );
  XNOR U892 ( .A(n442), .B(n441), .Z(n443) );
  XNOR U893 ( .A(in[1019]), .B(n443), .Z(n1092) );
  XOR U894 ( .A(in[1530]), .B(in[570]), .Z(n445) );
  XNOR U895 ( .A(in[1210]), .B(in[250]), .Z(n444) );
  XNOR U896 ( .A(n445), .B(n444), .Z(n446) );
  XNOR U897 ( .A(in[890]), .B(n446), .Z(n558) );
  XOR U898 ( .A(n1092), .B(n558), .Z(n3951) );
  XOR U899 ( .A(in[635]), .B(n3951), .Z(n2702) );
  IV U900 ( .A(n2702), .Z(n2788) );
  XOR U901 ( .A(in[161]), .B(in[1441]), .Z(n448) );
  XNOR U902 ( .A(in[801]), .B(in[1121]), .Z(n447) );
  XNOR U903 ( .A(n448), .B(n447), .Z(n449) );
  XNOR U904 ( .A(in[481]), .B(n449), .Z(n685) );
  XOR U905 ( .A(in[1570]), .B(in[610]), .Z(n451) );
  XNOR U906 ( .A(in[930]), .B(in[290]), .Z(n450) );
  XNOR U907 ( .A(n451), .B(n450), .Z(n452) );
  XOR U908 ( .A(in[1250]), .B(n452), .Z(n568) );
  XOR U909 ( .A(in[226]), .B(n4047), .Z(n3113) );
  XOR U910 ( .A(in[1510]), .B(in[550]), .Z(n454) );
  XNOR U911 ( .A(in[870]), .B(in[230]), .Z(n453) );
  XNOR U912 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U913 ( .A(in[1190]), .B(n455), .Z(n1506) );
  XOR U914 ( .A(in[1061]), .B(in[421]), .Z(n457) );
  XNOR U915 ( .A(in[741]), .B(in[1381]), .Z(n456) );
  XNOR U916 ( .A(n457), .B(n456), .Z(n458) );
  XNOR U917 ( .A(in[101]), .B(n458), .Z(n604) );
  XNOR U918 ( .A(n1506), .B(n604), .Z(n4087) );
  IV U919 ( .A(n4087), .Z(n1247) );
  XOR U920 ( .A(in[1446]), .B(n1247), .Z(n3110) );
  NANDN U921 ( .A(n3113), .B(n3110), .Z(n459) );
  XOR U922 ( .A(n2788), .B(n459), .Z(out[100]) );
  XOR U923 ( .A(in[1396]), .B(in[116]), .Z(n461) );
  XNOR U924 ( .A(in[1076]), .B(in[756]), .Z(n460) );
  XNOR U925 ( .A(n461), .B(n460), .Z(n462) );
  XNOR U926 ( .A(in[436]), .B(n462), .Z(n1627) );
  XOR U927 ( .A(in[1525]), .B(in[565]), .Z(n464) );
  XNOR U928 ( .A(in[885]), .B(in[245]), .Z(n463) );
  XNOR U929 ( .A(n464), .B(n463), .Z(n465) );
  XNOR U930 ( .A(in[1205]), .B(n465), .Z(n1568) );
  XOR U931 ( .A(n1627), .B(n1568), .Z(n4151) );
  XOR U932 ( .A(in[181]), .B(n4151), .Z(n1539) );
  XOR U933 ( .A(in[341]), .B(in[661]), .Z(n467) );
  XNOR U934 ( .A(in[21]), .B(in[1301]), .Z(n466) );
  XNOR U935 ( .A(n467), .B(n466), .Z(n468) );
  XNOR U936 ( .A(in[981]), .B(n468), .Z(n1448) );
  XOR U937 ( .A(in[150]), .B(in[1430]), .Z(n470) );
  XNOR U938 ( .A(in[1110]), .B(in[790]), .Z(n469) );
  XNOR U939 ( .A(n470), .B(n469), .Z(n471) );
  XOR U940 ( .A(in[470]), .B(n471), .Z(n779) );
  XNOR U941 ( .A(in[1366]), .B(n4492), .Z(n1946) );
  XOR U942 ( .A(in[1374]), .B(in[734]), .Z(n473) );
  XNOR U943 ( .A(in[94]), .B(in[414]), .Z(n472) );
  XNOR U944 ( .A(n473), .B(n472), .Z(n474) );
  XNOR U945 ( .A(in[1054]), .B(n474), .Z(n1147) );
  XOR U946 ( .A(in[1565]), .B(in[605]), .Z(n476) );
  XNOR U947 ( .A(in[925]), .B(in[285]), .Z(n475) );
  XNOR U948 ( .A(n476), .B(n475), .Z(n477) );
  XNOR U949 ( .A(in[1245]), .B(n477), .Z(n881) );
  XOR U950 ( .A(n1147), .B(n881), .Z(n4260) );
  XOR U951 ( .A(in[990]), .B(n4260), .Z(n1943) );
  NANDN U952 ( .A(n1946), .B(n1943), .Z(n478) );
  XNOR U953 ( .A(n1539), .B(n478), .Z(out[1010]) );
  XOR U954 ( .A(in[1526]), .B(in[566]), .Z(n480) );
  XNOR U955 ( .A(in[886]), .B(in[246]), .Z(n479) );
  XNOR U956 ( .A(n480), .B(n479), .Z(n481) );
  XNOR U957 ( .A(in[1206]), .B(n481), .Z(n1572) );
  XOR U958 ( .A(in[1397]), .B(in[117]), .Z(n483) );
  XNOR U959 ( .A(in[1077]), .B(in[757]), .Z(n482) );
  XNOR U960 ( .A(n483), .B(n482), .Z(n484) );
  XNOR U961 ( .A(in[437]), .B(n484), .Z(n1631) );
  XOR U962 ( .A(n1572), .B(n1631), .Z(n4161) );
  XOR U963 ( .A(in[182]), .B(n4161), .Z(n1543) );
  XOR U964 ( .A(in[342]), .B(in[662]), .Z(n486) );
  XNOR U965 ( .A(in[22]), .B(in[1302]), .Z(n485) );
  XNOR U966 ( .A(n486), .B(n485), .Z(n487) );
  XNOR U967 ( .A(in[982]), .B(n487), .Z(n1450) );
  XOR U968 ( .A(in[151]), .B(in[1431]), .Z(n489) );
  XNOR U969 ( .A(in[1111]), .B(in[791]), .Z(n488) );
  XNOR U970 ( .A(n489), .B(n488), .Z(n490) );
  XOR U971 ( .A(in[471]), .B(n490), .Z(n794) );
  XNOR U972 ( .A(in[1367]), .B(n4495), .Z(n1950) );
  XOR U973 ( .A(in[1375]), .B(in[735]), .Z(n492) );
  XNOR U974 ( .A(in[95]), .B(in[415]), .Z(n491) );
  XNOR U975 ( .A(n492), .B(n491), .Z(n493) );
  XNOR U976 ( .A(in[1055]), .B(n493), .Z(n1160) );
  XOR U977 ( .A(in[1566]), .B(in[606]), .Z(n495) );
  XNOR U978 ( .A(in[926]), .B(in[286]), .Z(n494) );
  XNOR U979 ( .A(n495), .B(n494), .Z(n496) );
  XNOR U980 ( .A(in[1246]), .B(n496), .Z(n896) );
  XOR U981 ( .A(n1160), .B(n896), .Z(n4261) );
  XOR U982 ( .A(in[991]), .B(n4261), .Z(n1947) );
  NANDN U983 ( .A(n1950), .B(n1947), .Z(n497) );
  XNOR U984 ( .A(n1543), .B(n497), .Z(out[1011]) );
  XOR U985 ( .A(in[1527]), .B(in[567]), .Z(n499) );
  XNOR U986 ( .A(in[887]), .B(in[247]), .Z(n498) );
  XNOR U987 ( .A(n499), .B(n498), .Z(n500) );
  XNOR U988 ( .A(in[1207]), .B(n500), .Z(n1576) );
  XOR U989 ( .A(in[1398]), .B(in[118]), .Z(n502) );
  XNOR U990 ( .A(in[1078]), .B(in[758]), .Z(n501) );
  XNOR U991 ( .A(n502), .B(n501), .Z(n503) );
  XNOR U992 ( .A(in[438]), .B(n503), .Z(n1635) );
  XOR U993 ( .A(n1576), .B(n1635), .Z(n4165) );
  XOR U994 ( .A(in[183]), .B(n4165), .Z(n1549) );
  XOR U995 ( .A(in[343]), .B(in[663]), .Z(n505) );
  XNOR U996 ( .A(in[23]), .B(in[1303]), .Z(n504) );
  XNOR U997 ( .A(n505), .B(n504), .Z(n506) );
  XNOR U998 ( .A(in[983]), .B(n506), .Z(n1452) );
  XOR U999 ( .A(in[152]), .B(in[1432]), .Z(n508) );
  XNOR U1000 ( .A(in[1112]), .B(in[792]), .Z(n507) );
  XNOR U1001 ( .A(n508), .B(n507), .Z(n509) );
  XOR U1002 ( .A(in[472]), .B(n509), .Z(n820) );
  XNOR U1003 ( .A(in[1368]), .B(n4498), .Z(n1954) );
  XOR U1004 ( .A(in[1376]), .B(in[736]), .Z(n511) );
  XNOR U1005 ( .A(in[96]), .B(in[416]), .Z(n510) );
  XNOR U1006 ( .A(n511), .B(n510), .Z(n512) );
  XNOR U1007 ( .A(in[1056]), .B(n512), .Z(n1175) );
  XOR U1008 ( .A(in[1567]), .B(in[607]), .Z(n514) );
  XNOR U1009 ( .A(in[927]), .B(in[287]), .Z(n513) );
  XNOR U1010 ( .A(n514), .B(n513), .Z(n515) );
  XNOR U1011 ( .A(in[1247]), .B(n515), .Z(n911) );
  XOR U1012 ( .A(n1175), .B(n911), .Z(n4264) );
  XOR U1013 ( .A(in[992]), .B(n4264), .Z(n1951) );
  NANDN U1014 ( .A(n1954), .B(n1951), .Z(n516) );
  XNOR U1015 ( .A(n1549), .B(n516), .Z(out[1012]) );
  XOR U1016 ( .A(in[1528]), .B(in[568]), .Z(n518) );
  XNOR U1017 ( .A(in[888]), .B(in[248]), .Z(n517) );
  XNOR U1018 ( .A(n518), .B(n517), .Z(n519) );
  XNOR U1019 ( .A(in[1208]), .B(n519), .Z(n1580) );
  XOR U1020 ( .A(in[1399]), .B(in[119]), .Z(n521) );
  XNOR U1021 ( .A(in[1079]), .B(in[759]), .Z(n520) );
  XNOR U1022 ( .A(n521), .B(n520), .Z(n522) );
  XNOR U1023 ( .A(in[439]), .B(n522), .Z(n1639) );
  XOR U1024 ( .A(n1580), .B(n1639), .Z(n4169) );
  XOR U1025 ( .A(in[184]), .B(n4169), .Z(n1553) );
  XOR U1026 ( .A(in[153]), .B(in[1433]), .Z(n524) );
  XNOR U1027 ( .A(in[1113]), .B(in[793]), .Z(n523) );
  XNOR U1028 ( .A(n524), .B(n523), .Z(n525) );
  XNOR U1029 ( .A(in[473]), .B(n525), .Z(n835) );
  XOR U1030 ( .A(in[344]), .B(in[664]), .Z(n527) );
  XNOR U1031 ( .A(in[24]), .B(in[1304]), .Z(n526) );
  XNOR U1032 ( .A(n527), .B(n526), .Z(n528) );
  XOR U1033 ( .A(in[984]), .B(n528), .Z(n1454) );
  XNOR U1034 ( .A(in[1369]), .B(n4501), .Z(n1958) );
  XOR U1035 ( .A(in[1377]), .B(in[737]), .Z(n530) );
  XNOR U1036 ( .A(in[97]), .B(in[417]), .Z(n529) );
  XNOR U1037 ( .A(n530), .B(n529), .Z(n531) );
  XNOR U1038 ( .A(in[1057]), .B(n531), .Z(n1190) );
  XOR U1039 ( .A(in[1568]), .B(in[608]), .Z(n533) );
  XNOR U1040 ( .A(in[928]), .B(in[288]), .Z(n532) );
  XNOR U1041 ( .A(n533), .B(n532), .Z(n534) );
  XNOR U1042 ( .A(in[1248]), .B(n534), .Z(n926) );
  XOR U1043 ( .A(n1190), .B(n926), .Z(n4267) );
  XOR U1044 ( .A(in[993]), .B(n4267), .Z(n1955) );
  NANDN U1045 ( .A(n1958), .B(n1955), .Z(n535) );
  XNOR U1046 ( .A(n1553), .B(n535), .Z(out[1013]) );
  XOR U1047 ( .A(in[1529]), .B(in[569]), .Z(n537) );
  XNOR U1048 ( .A(in[889]), .B(in[249]), .Z(n536) );
  XNOR U1049 ( .A(n537), .B(n536), .Z(n538) );
  XNOR U1050 ( .A(in[1209]), .B(n538), .Z(n1584) );
  XOR U1051 ( .A(in[1400]), .B(in[120]), .Z(n540) );
  XNOR U1052 ( .A(in[1080]), .B(in[760]), .Z(n539) );
  XNOR U1053 ( .A(n540), .B(n539), .Z(n541) );
  XNOR U1054 ( .A(in[440]), .B(n541), .Z(n1643) );
  XOR U1055 ( .A(n1584), .B(n1643), .Z(n4173) );
  XOR U1056 ( .A(in[185]), .B(n4173), .Z(n1557) );
  XOR U1057 ( .A(in[154]), .B(in[1434]), .Z(n543) );
  XNOR U1058 ( .A(in[1114]), .B(in[794]), .Z(n542) );
  XNOR U1059 ( .A(n543), .B(n542), .Z(n544) );
  XNOR U1060 ( .A(in[474]), .B(n544), .Z(n850) );
  XOR U1061 ( .A(in[345]), .B(in[665]), .Z(n546) );
  XNOR U1062 ( .A(in[25]), .B(in[1305]), .Z(n545) );
  XNOR U1063 ( .A(n546), .B(n545), .Z(n547) );
  XOR U1064 ( .A(in[985]), .B(n547), .Z(n1458) );
  XNOR U1065 ( .A(in[1370]), .B(n4504), .Z(n1964) );
  XOR U1066 ( .A(in[1569]), .B(in[609]), .Z(n549) );
  XNOR U1067 ( .A(in[929]), .B(in[289]), .Z(n548) );
  XNOR U1068 ( .A(n549), .B(n548), .Z(n550) );
  XNOR U1069 ( .A(in[1249]), .B(n550), .Z(n941) );
  XOR U1070 ( .A(in[1378]), .B(in[738]), .Z(n552) );
  XNOR U1071 ( .A(in[98]), .B(in[418]), .Z(n551) );
  XNOR U1072 ( .A(n552), .B(n551), .Z(n553) );
  XNOR U1073 ( .A(in[1058]), .B(n553), .Z(n1205) );
  XOR U1074 ( .A(n941), .B(n1205), .Z(n4270) );
  XOR U1075 ( .A(in[994]), .B(n4270), .Z(n1961) );
  NANDN U1076 ( .A(n1964), .B(n1961), .Z(n554) );
  XNOR U1077 ( .A(n1557), .B(n554), .Z(out[1014]) );
  XOR U1078 ( .A(in[1401]), .B(in[121]), .Z(n556) );
  XNOR U1079 ( .A(in[1081]), .B(in[761]), .Z(n555) );
  XNOR U1080 ( .A(n556), .B(n555), .Z(n557) );
  XNOR U1081 ( .A(in[441]), .B(n557), .Z(n1647) );
  XOR U1082 ( .A(n558), .B(n1647), .Z(n1794) );
  XOR U1083 ( .A(in[186]), .B(n1794), .Z(n1561) );
  XOR U1084 ( .A(in[155]), .B(in[1435]), .Z(n560) );
  XNOR U1085 ( .A(in[1115]), .B(in[795]), .Z(n559) );
  XNOR U1086 ( .A(n560), .B(n559), .Z(n561) );
  XNOR U1087 ( .A(in[475]), .B(n561), .Z(n865) );
  XOR U1088 ( .A(in[346]), .B(in[666]), .Z(n563) );
  XNOR U1089 ( .A(in[26]), .B(in[1306]), .Z(n562) );
  XNOR U1090 ( .A(n563), .B(n562), .Z(n564) );
  XOR U1091 ( .A(in[986]), .B(n564), .Z(n1460) );
  IV U1092 ( .A(n4511), .Z(n2738) );
  XOR U1093 ( .A(in[1371]), .B(n2738), .Z(n1363) );
  IV U1094 ( .A(n1363), .Z(n1968) );
  XOR U1095 ( .A(in[1379]), .B(in[739]), .Z(n566) );
  XNOR U1096 ( .A(in[99]), .B(in[419]), .Z(n565) );
  XNOR U1097 ( .A(n566), .B(n565), .Z(n567) );
  XOR U1098 ( .A(in[1059]), .B(n567), .Z(n1220) );
  XNOR U1099 ( .A(n568), .B(n1220), .Z(n4273) );
  XNOR U1100 ( .A(in[995]), .B(n4273), .Z(n1965) );
  NANDN U1101 ( .A(n1968), .B(n1965), .Z(n569) );
  XNOR U1102 ( .A(n1561), .B(n569), .Z(out[1015]) );
  XOR U1103 ( .A(in[1402]), .B(in[122]), .Z(n571) );
  XNOR U1104 ( .A(in[1082]), .B(in[762]), .Z(n570) );
  XNOR U1105 ( .A(n571), .B(n570), .Z(n572) );
  XNOR U1106 ( .A(in[442]), .B(n572), .Z(n1651) );
  XOR U1107 ( .A(in[1531]), .B(in[571]), .Z(n574) );
  XNOR U1108 ( .A(in[1211]), .B(in[251]), .Z(n573) );
  XNOR U1109 ( .A(n574), .B(n573), .Z(n575) );
  XNOR U1110 ( .A(in[891]), .B(n575), .Z(n647) );
  XOR U1111 ( .A(n1651), .B(n647), .Z(n1820) );
  XOR U1112 ( .A(in[187]), .B(n1820), .Z(n1565) );
  XOR U1113 ( .A(in[156]), .B(in[1436]), .Z(n577) );
  XNOR U1114 ( .A(in[1116]), .B(in[796]), .Z(n576) );
  XNOR U1115 ( .A(n577), .B(n576), .Z(n578) );
  XNOR U1116 ( .A(in[476]), .B(n578), .Z(n880) );
  XOR U1117 ( .A(in[347]), .B(in[667]), .Z(n580) );
  XNOR U1118 ( .A(in[27]), .B(in[1307]), .Z(n579) );
  XNOR U1119 ( .A(n580), .B(n579), .Z(n581) );
  XOR U1120 ( .A(in[987]), .B(n581), .Z(n1462) );
  IV U1121 ( .A(n4514), .Z(n2755) );
  XOR U1122 ( .A(in[1372]), .B(n2755), .Z(n1373) );
  IV U1123 ( .A(n1373), .Z(n1972) );
  XOR U1124 ( .A(in[1060]), .B(in[420]), .Z(n583) );
  XNOR U1125 ( .A(in[740]), .B(in[1380]), .Z(n582) );
  XNOR U1126 ( .A(n583), .B(n582), .Z(n584) );
  XNOR U1127 ( .A(in[100]), .B(n584), .Z(n1235) );
  XOR U1128 ( .A(in[1571]), .B(in[611]), .Z(n586) );
  XNOR U1129 ( .A(in[931]), .B(in[291]), .Z(n585) );
  XNOR U1130 ( .A(n586), .B(n585), .Z(n587) );
  XNOR U1131 ( .A(in[1251]), .B(n587), .Z(n651) );
  XOR U1132 ( .A(n1235), .B(n651), .Z(n4276) );
  XOR U1133 ( .A(in[996]), .B(n4276), .Z(n1969) );
  NANDN U1134 ( .A(n1972), .B(n1969), .Z(n588) );
  XNOR U1135 ( .A(n1565), .B(n588), .Z(out[1016]) );
  XOR U1136 ( .A(in[1403]), .B(in[123]), .Z(n590) );
  XNOR U1137 ( .A(in[1083]), .B(in[763]), .Z(n589) );
  XNOR U1138 ( .A(n590), .B(n589), .Z(n591) );
  XNOR U1139 ( .A(in[443]), .B(n591), .Z(n1655) );
  XOR U1140 ( .A(in[1532]), .B(in[572]), .Z(n593) );
  XNOR U1141 ( .A(in[1212]), .B(in[252]), .Z(n592) );
  XNOR U1142 ( .A(n593), .B(n592), .Z(n594) );
  XNOR U1143 ( .A(in[892]), .B(n594), .Z(n812) );
  XOR U1144 ( .A(n1655), .B(n812), .Z(n1843) );
  XOR U1145 ( .A(in[188]), .B(n1843), .Z(n1569) );
  XOR U1146 ( .A(in[157]), .B(in[1437]), .Z(n596) );
  XNOR U1147 ( .A(in[1117]), .B(in[797]), .Z(n595) );
  XNOR U1148 ( .A(n596), .B(n595), .Z(n597) );
  XNOR U1149 ( .A(in[477]), .B(n597), .Z(n895) );
  XOR U1150 ( .A(in[348]), .B(in[668]), .Z(n599) );
  XNOR U1151 ( .A(in[28]), .B(in[1308]), .Z(n598) );
  XNOR U1152 ( .A(n599), .B(n598), .Z(n600) );
  XOR U1153 ( .A(in[988]), .B(n600), .Z(n1466) );
  IV U1154 ( .A(n4517), .Z(n2772) );
  XOR U1155 ( .A(in[1373]), .B(n2772), .Z(n1379) );
  IV U1156 ( .A(n1379), .Z(n1976) );
  XOR U1157 ( .A(in[1572]), .B(in[612]), .Z(n602) );
  XNOR U1158 ( .A(in[932]), .B(in[292]), .Z(n601) );
  XNOR U1159 ( .A(n602), .B(n601), .Z(n603) );
  XNOR U1160 ( .A(in[1252]), .B(n603), .Z(n814) );
  XOR U1161 ( .A(n604), .B(n814), .Z(n4278) );
  XOR U1162 ( .A(in[997]), .B(n4278), .Z(n1973) );
  NANDN U1163 ( .A(n1976), .B(n1973), .Z(n605) );
  XNOR U1164 ( .A(n1569), .B(n605), .Z(out[1017]) );
  XOR U1165 ( .A(in[1404]), .B(in[124]), .Z(n607) );
  XNOR U1166 ( .A(in[1084]), .B(in[764]), .Z(n606) );
  XNOR U1167 ( .A(n607), .B(n606), .Z(n608) );
  XNOR U1168 ( .A(in[444]), .B(n608), .Z(n1659) );
  XOR U1169 ( .A(in[1533]), .B(in[573]), .Z(n610) );
  XNOR U1170 ( .A(in[1213]), .B(in[253]), .Z(n609) );
  XNOR U1171 ( .A(n610), .B(n609), .Z(n611) );
  XNOR U1172 ( .A(in[893]), .B(n611), .Z(n971) );
  XOR U1173 ( .A(n1659), .B(n971), .Z(n1865) );
  XOR U1174 ( .A(in[189]), .B(n1865), .Z(n1573) );
  XOR U1175 ( .A(in[158]), .B(in[1438]), .Z(n613) );
  XNOR U1176 ( .A(in[1118]), .B(in[798]), .Z(n612) );
  XNOR U1177 ( .A(n613), .B(n612), .Z(n614) );
  XNOR U1178 ( .A(in[478]), .B(n614), .Z(n910) );
  XOR U1179 ( .A(in[349]), .B(in[669]), .Z(n616) );
  XNOR U1180 ( .A(in[29]), .B(in[1309]), .Z(n615) );
  XNOR U1181 ( .A(n616), .B(n615), .Z(n617) );
  XOR U1182 ( .A(in[989]), .B(n617), .Z(n1472) );
  XNOR U1183 ( .A(in[1374]), .B(n4520), .Z(n1980) );
  XOR U1184 ( .A(in[1062]), .B(in[422]), .Z(n619) );
  XNOR U1185 ( .A(in[742]), .B(in[1382]), .Z(n618) );
  XNOR U1186 ( .A(n619), .B(n618), .Z(n620) );
  XNOR U1187 ( .A(in[102]), .B(n620), .Z(n655) );
  XOR U1188 ( .A(in[1573]), .B(in[613]), .Z(n622) );
  XNOR U1189 ( .A(in[933]), .B(in[293]), .Z(n621) );
  XNOR U1190 ( .A(n622), .B(n621), .Z(n623) );
  XNOR U1191 ( .A(in[1253]), .B(n623), .Z(n973) );
  XOR U1192 ( .A(n655), .B(n973), .Z(n4284) );
  XOR U1193 ( .A(in[998]), .B(n4284), .Z(n1977) );
  NANDN U1194 ( .A(n1980), .B(n1977), .Z(n624) );
  XNOR U1195 ( .A(n1573), .B(n624), .Z(out[1018]) );
  XOR U1196 ( .A(in[1405]), .B(in[125]), .Z(n626) );
  XNOR U1197 ( .A(in[1085]), .B(in[765]), .Z(n625) );
  XNOR U1198 ( .A(n626), .B(n625), .Z(n627) );
  XNOR U1199 ( .A(in[445]), .B(n627), .Z(n1663) );
  XOR U1200 ( .A(in[1534]), .B(in[894]), .Z(n629) );
  XNOR U1201 ( .A(in[574]), .B(in[1214]), .Z(n628) );
  XNOR U1202 ( .A(n629), .B(n628), .Z(n630) );
  XNOR U1203 ( .A(in[254]), .B(n630), .Z(n1108) );
  XOR U1204 ( .A(n1663), .B(n1108), .Z(n1887) );
  XOR U1205 ( .A(in[190]), .B(n1887), .Z(n1577) );
  XOR U1206 ( .A(in[1439]), .B(in[479]), .Z(n632) );
  XNOR U1207 ( .A(in[799]), .B(in[159]), .Z(n631) );
  XNOR U1208 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U1209 ( .A(in[1119]), .B(n633), .Z(n925) );
  XOR U1210 ( .A(in[350]), .B(in[670]), .Z(n635) );
  XNOR U1211 ( .A(in[30]), .B(in[1310]), .Z(n634) );
  XNOR U1212 ( .A(n635), .B(n634), .Z(n636) );
  XOR U1213 ( .A(in[990]), .B(n636), .Z(n1476) );
  XNOR U1214 ( .A(in[1375]), .B(n4524), .Z(n1984) );
  XOR U1215 ( .A(in[1063]), .B(in[423]), .Z(n638) );
  XNOR U1216 ( .A(in[743]), .B(in[1383]), .Z(n637) );
  XNOR U1217 ( .A(n638), .B(n637), .Z(n639) );
  XNOR U1218 ( .A(in[103]), .B(n639), .Z(n818) );
  XOR U1219 ( .A(in[1574]), .B(in[614]), .Z(n641) );
  XNOR U1220 ( .A(in[934]), .B(in[294]), .Z(n640) );
  XNOR U1221 ( .A(n641), .B(n640), .Z(n642) );
  XNOR U1222 ( .A(in[1254]), .B(n642), .Z(n1017) );
  XOR U1223 ( .A(n818), .B(n1017), .Z(n4286) );
  XOR U1224 ( .A(in[999]), .B(n4286), .Z(n1981) );
  NANDN U1225 ( .A(n1984), .B(n1981), .Z(n643) );
  XNOR U1226 ( .A(n1577), .B(n643), .Z(out[1019]) );
  XOR U1227 ( .A(in[1340]), .B(in[60]), .Z(n645) );
  XNOR U1228 ( .A(in[700]), .B(in[380]), .Z(n644) );
  XNOR U1229 ( .A(n645), .B(n644), .Z(n646) );
  XNOR U1230 ( .A(in[1020]), .B(n646), .Z(n1102) );
  XOR U1231 ( .A(n647), .B(n1102), .Z(n3955) );
  XOR U1232 ( .A(in[636]), .B(n3955), .Z(n2704) );
  IV U1233 ( .A(n2704), .Z(n2790) );
  XOR U1234 ( .A(in[162]), .B(in[1442]), .Z(n649) );
  XNOR U1235 ( .A(in[802]), .B(in[1122]), .Z(n648) );
  XNOR U1236 ( .A(n649), .B(n648), .Z(n650) );
  XOR U1237 ( .A(in[482]), .B(n650), .Z(n702) );
  XOR U1238 ( .A(n651), .B(n702), .Z(n3396) );
  IV U1239 ( .A(n3396), .Z(n4051) );
  XOR U1240 ( .A(in[227]), .B(n4051), .Z(n3135) );
  XOR U1241 ( .A(in[1511]), .B(in[551]), .Z(n653) );
  XNOR U1242 ( .A(in[871]), .B(in[231]), .Z(n652) );
  XNOR U1243 ( .A(n653), .B(n652), .Z(n654) );
  XNOR U1244 ( .A(in[1191]), .B(n654), .Z(n1510) );
  XNOR U1245 ( .A(n655), .B(n1510), .Z(n4091) );
  IV U1246 ( .A(n4091), .Z(n1262) );
  XOR U1247 ( .A(in[1447]), .B(n1262), .Z(n3132) );
  NANDN U1248 ( .A(n3135), .B(n3132), .Z(n656) );
  XOR U1249 ( .A(n2790), .B(n656), .Z(out[101]) );
  XOR U1250 ( .A(in[1406]), .B(in[126]), .Z(n658) );
  XNOR U1251 ( .A(in[1086]), .B(in[766]), .Z(n657) );
  XNOR U1252 ( .A(n658), .B(n657), .Z(n659) );
  XNOR U1253 ( .A(in[446]), .B(n659), .Z(n1668) );
  XOR U1254 ( .A(in[1535]), .B(in[575]), .Z(n661) );
  XNOR U1255 ( .A(in[895]), .B(in[255]), .Z(n660) );
  XNOR U1256 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U1257 ( .A(in[1215]), .B(n662), .Z(n1256) );
  XOR U1258 ( .A(n1668), .B(n1256), .Z(n1917) );
  XOR U1259 ( .A(in[191]), .B(n1917), .Z(n1581) );
  XOR U1260 ( .A(in[1440]), .B(in[480]), .Z(n664) );
  XNOR U1261 ( .A(in[800]), .B(in[160]), .Z(n663) );
  XNOR U1262 ( .A(n664), .B(n663), .Z(n665) );
  XNOR U1263 ( .A(in[1120]), .B(n665), .Z(n940) );
  XOR U1264 ( .A(in[351]), .B(in[671]), .Z(n667) );
  XNOR U1265 ( .A(in[31]), .B(in[1311]), .Z(n666) );
  XNOR U1266 ( .A(n667), .B(n666), .Z(n668) );
  XOR U1267 ( .A(in[991]), .B(n668), .Z(n1480) );
  XNOR U1268 ( .A(in[1376]), .B(n4528), .Z(n1988) );
  XOR U1269 ( .A(in[1064]), .B(in[424]), .Z(n670) );
  XNOR U1270 ( .A(in[744]), .B(in[1384]), .Z(n669) );
  XNOR U1271 ( .A(n670), .B(n669), .Z(n671) );
  XNOR U1272 ( .A(in[104]), .B(n671), .Z(n977) );
  XOR U1273 ( .A(in[1575]), .B(in[615]), .Z(n673) );
  XNOR U1274 ( .A(in[935]), .B(in[295]), .Z(n672) );
  XNOR U1275 ( .A(n673), .B(n672), .Z(n674) );
  XNOR U1276 ( .A(in[1255]), .B(n674), .Z(n1030) );
  XOR U1277 ( .A(n977), .B(n1030), .Z(n4288) );
  XOR U1278 ( .A(in[1000]), .B(n4288), .Z(n1985) );
  NANDN U1279 ( .A(n1988), .B(n1985), .Z(n675) );
  XNOR U1280 ( .A(n1581), .B(n675), .Z(out[1020]) );
  XOR U1281 ( .A(in[1407]), .B(in[127]), .Z(n677) );
  XNOR U1282 ( .A(in[1087]), .B(in[767]), .Z(n676) );
  XNOR U1283 ( .A(n677), .B(n676), .Z(n678) );
  XNOR U1284 ( .A(in[447]), .B(n678), .Z(n1671) );
  XOR U1285 ( .A(in[1472]), .B(in[512]), .Z(n680) );
  XNOR U1286 ( .A(in[832]), .B(in[192]), .Z(n679) );
  XNOR U1287 ( .A(n680), .B(n679), .Z(n681) );
  XNOR U1288 ( .A(in[1152]), .B(n681), .Z(n1321) );
  XOR U1289 ( .A(n1671), .B(n1321), .Z(n1959) );
  XOR U1290 ( .A(in[128]), .B(n1959), .Z(n1585) );
  XOR U1291 ( .A(in[352]), .B(in[672]), .Z(n683) );
  XNOR U1292 ( .A(in[32]), .B(in[1312]), .Z(n682) );
  XNOR U1293 ( .A(n683), .B(n682), .Z(n684) );
  XOR U1294 ( .A(in[992]), .B(n684), .Z(n1482) );
  XNOR U1295 ( .A(in[1377]), .B(n4532), .Z(n1992) );
  XOR U1296 ( .A(in[1065]), .B(in[425]), .Z(n687) );
  XNOR U1297 ( .A(in[745]), .B(in[1385]), .Z(n686) );
  XNOR U1298 ( .A(n687), .B(n686), .Z(n688) );
  XNOR U1299 ( .A(in[105]), .B(n688), .Z(n1112) );
  XOR U1300 ( .A(in[1576]), .B(in[616]), .Z(n690) );
  XNOR U1301 ( .A(in[936]), .B(in[296]), .Z(n689) );
  XNOR U1302 ( .A(n690), .B(n689), .Z(n691) );
  XNOR U1303 ( .A(in[1256]), .B(n691), .Z(n1043) );
  XOR U1304 ( .A(n1112), .B(n1043), .Z(n4290) );
  XOR U1305 ( .A(in[1001]), .B(n4290), .Z(n1989) );
  NANDN U1306 ( .A(n1992), .B(n1989), .Z(n692) );
  XNOR U1307 ( .A(n1585), .B(n692), .Z(out[1021]) );
  XOR U1308 ( .A(in[1344]), .B(in[64]), .Z(n694) );
  XNOR U1309 ( .A(in[1024]), .B(in[384]), .Z(n693) );
  XNOR U1310 ( .A(n694), .B(n693), .Z(n695) );
  XNOR U1311 ( .A(in[704]), .B(n695), .Z(n1676) );
  XOR U1312 ( .A(in[1473]), .B(in[513]), .Z(n697) );
  XNOR U1313 ( .A(in[833]), .B(in[193]), .Z(n696) );
  XNOR U1314 ( .A(n697), .B(n696), .Z(n698) );
  XNOR U1315 ( .A(in[1153]), .B(n698), .Z(n1366) );
  XOR U1316 ( .A(n1676), .B(n1366), .Z(n2001) );
  XOR U1317 ( .A(in[129]), .B(n2001), .Z(n1589) );
  XOR U1318 ( .A(in[353]), .B(in[673]), .Z(n700) );
  XNOR U1319 ( .A(in[33]), .B(in[1313]), .Z(n699) );
  XNOR U1320 ( .A(n700), .B(n699), .Z(n701) );
  XNOR U1321 ( .A(in[993]), .B(n701), .Z(n1485) );
  XNOR U1322 ( .A(in[1378]), .B(n4536), .Z(n1996) );
  XOR U1323 ( .A(in[1577]), .B(in[617]), .Z(n704) );
  XNOR U1324 ( .A(in[937]), .B(in[297]), .Z(n703) );
  XNOR U1325 ( .A(n704), .B(n703), .Z(n705) );
  XNOR U1326 ( .A(in[1257]), .B(n705), .Z(n1056) );
  XOR U1327 ( .A(n706), .B(n1056), .Z(n4292) );
  XOR U1328 ( .A(in[1002]), .B(n4292), .Z(n1993) );
  NANDN U1329 ( .A(n1996), .B(n1993), .Z(n707) );
  XNOR U1330 ( .A(n1589), .B(n707), .Z(out[1022]) );
  IV U1331 ( .A(n3169), .Z(n3930) );
  XOR U1332 ( .A(n3930), .B(in[130]), .Z(n1591) );
  XOR U1333 ( .A(in[163]), .B(in[1443]), .Z(n709) );
  XNOR U1334 ( .A(in[803]), .B(in[1123]), .Z(n708) );
  XNOR U1335 ( .A(n709), .B(n708), .Z(n710) );
  XNOR U1336 ( .A(in[483]), .B(n710), .Z(n813) );
  XOR U1337 ( .A(in[354]), .B(in[674]), .Z(n712) );
  XNOR U1338 ( .A(in[34]), .B(in[1314]), .Z(n711) );
  XNOR U1339 ( .A(n712), .B(n711), .Z(n713) );
  XOR U1340 ( .A(in[994]), .B(n713), .Z(n1487) );
  XNOR U1341 ( .A(in[1379]), .B(n4540), .Z(n2000) );
  XOR U1342 ( .A(in[1578]), .B(in[618]), .Z(n715) );
  XNOR U1343 ( .A(in[938]), .B(in[298]), .Z(n714) );
  XNOR U1344 ( .A(n715), .B(n714), .Z(n716) );
  XNOR U1345 ( .A(in[1258]), .B(n716), .Z(n1069) );
  XOR U1346 ( .A(n717), .B(n1069), .Z(n4294) );
  XOR U1347 ( .A(in[1003]), .B(n4294), .Z(n1997) );
  NANDN U1348 ( .A(n2000), .B(n1997), .Z(n718) );
  XOR U1349 ( .A(n1591), .B(n718), .Z(out[1023]) );
  XOR U1350 ( .A(n720), .B(n719), .Z(n3983) );
  XOR U1351 ( .A(in[531]), .B(n3983), .Z(n1595) );
  XOR U1352 ( .A(in[35]), .B(in[675]), .Z(n722) );
  XNOR U1353 ( .A(in[355]), .B(in[1315]), .Z(n721) );
  XNOR U1354 ( .A(n722), .B(n721), .Z(n723) );
  XNOR U1355 ( .A(in[995]), .B(n723), .Z(n1490) );
  XOR U1356 ( .A(in[164]), .B(in[1444]), .Z(n725) );
  XNOR U1357 ( .A(in[804]), .B(in[1124]), .Z(n724) );
  XNOR U1358 ( .A(n725), .B(n724), .Z(n726) );
  XNOR U1359 ( .A(in[484]), .B(n726), .Z(n972) );
  XOR U1360 ( .A(n1490), .B(n972), .Z(n4544) );
  XNOR U1361 ( .A(in[1380]), .B(n4544), .Z(n4999) );
  XOR U1362 ( .A(in[1346]), .B(in[66]), .Z(n728) );
  XNOR U1363 ( .A(in[1026]), .B(in[386]), .Z(n727) );
  XNOR U1364 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U1365 ( .A(in[706]), .B(n729), .Z(n1684) );
  XOR U1366 ( .A(in[1475]), .B(in[515]), .Z(n731) );
  XNOR U1367 ( .A(in[835]), .B(in[195]), .Z(n730) );
  XNOR U1368 ( .A(n731), .B(n730), .Z(n732) );
  XOR U1369 ( .A(in[1155]), .B(n732), .Z(n1409) );
  XOR U1370 ( .A(in[131]), .B(n3171), .Z(n5001) );
  OR U1371 ( .A(n4999), .B(n5001), .Z(n733) );
  XNOR U1372 ( .A(n1595), .B(n733), .Z(out[1024]) );
  XNOR U1373 ( .A(n735), .B(n734), .Z(n3987) );
  XOR U1374 ( .A(in[532]), .B(n3987), .Z(n1599) );
  XOR U1375 ( .A(in[36]), .B(in[676]), .Z(n737) );
  XNOR U1376 ( .A(in[356]), .B(in[1316]), .Z(n736) );
  XNOR U1377 ( .A(n737), .B(n736), .Z(n738) );
  XNOR U1378 ( .A(in[996]), .B(n738), .Z(n1493) );
  XOR U1379 ( .A(in[1445]), .B(in[165]), .Z(n740) );
  XNOR U1380 ( .A(in[805]), .B(in[1125]), .Z(n739) );
  XNOR U1381 ( .A(n740), .B(n739), .Z(n741) );
  XNOR U1382 ( .A(in[485]), .B(n741), .Z(n1016) );
  XOR U1383 ( .A(n1493), .B(n1016), .Z(n4550) );
  XNOR U1384 ( .A(in[1381]), .B(n4550), .Z(n5003) );
  XOR U1385 ( .A(in[1347]), .B(in[67]), .Z(n743) );
  XNOR U1386 ( .A(in[1027]), .B(in[387]), .Z(n742) );
  XNOR U1387 ( .A(n743), .B(n742), .Z(n744) );
  XNOR U1388 ( .A(in[707]), .B(n744), .Z(n1688) );
  XOR U1389 ( .A(in[1476]), .B(in[516]), .Z(n746) );
  XNOR U1390 ( .A(in[836]), .B(in[196]), .Z(n745) );
  XNOR U1391 ( .A(n746), .B(n745), .Z(n747) );
  XOR U1392 ( .A(in[1156]), .B(n747), .Z(n1411) );
  XOR U1393 ( .A(in[132]), .B(n3173), .Z(n5005) );
  OR U1394 ( .A(n5003), .B(n5005), .Z(n748) );
  XNOR U1395 ( .A(n1599), .B(n748), .Z(out[1025]) );
  XOR U1396 ( .A(n750), .B(n749), .Z(n2004) );
  XOR U1397 ( .A(in[533]), .B(n2004), .Z(n1603) );
  XOR U1398 ( .A(in[166]), .B(in[806]), .Z(n752) );
  XNOR U1399 ( .A(in[1126]), .B(in[486]), .Z(n751) );
  XNOR U1400 ( .A(n752), .B(n751), .Z(n753) );
  XNOR U1401 ( .A(in[1446]), .B(n753), .Z(n1029) );
  XOR U1402 ( .A(in[37]), .B(in[677]), .Z(n755) );
  XNOR U1403 ( .A(in[357]), .B(in[1317]), .Z(n754) );
  XNOR U1404 ( .A(n755), .B(n754), .Z(n756) );
  XNOR U1405 ( .A(in[997]), .B(n756), .Z(n1496) );
  XOR U1406 ( .A(n1029), .B(n1496), .Z(n4552) );
  XNOR U1407 ( .A(in[1382]), .B(n4552), .Z(n5007) );
  XOR U1408 ( .A(in[1348]), .B(in[68]), .Z(n758) );
  XNOR U1409 ( .A(in[1028]), .B(in[388]), .Z(n757) );
  XNOR U1410 ( .A(n758), .B(n757), .Z(n759) );
  XNOR U1411 ( .A(in[708]), .B(n759), .Z(n1692) );
  XOR U1412 ( .A(in[1477]), .B(in[517]), .Z(n761) );
  XNOR U1413 ( .A(in[837]), .B(in[197]), .Z(n760) );
  XNOR U1414 ( .A(n761), .B(n760), .Z(n762) );
  XOR U1415 ( .A(in[1157]), .B(n762), .Z(n1413) );
  XOR U1416 ( .A(in[133]), .B(n3175), .Z(n5009) );
  OR U1417 ( .A(n5007), .B(n5009), .Z(n763) );
  XNOR U1418 ( .A(n1603), .B(n763), .Z(out[1026]) );
  XOR U1419 ( .A(n765), .B(n764), .Z(n2006) );
  XOR U1420 ( .A(in[534]), .B(n2006), .Z(n1607) );
  XOR U1421 ( .A(in[38]), .B(in[678]), .Z(n767) );
  XNOR U1422 ( .A(in[358]), .B(in[1318]), .Z(n766) );
  XNOR U1423 ( .A(n767), .B(n766), .Z(n768) );
  XNOR U1424 ( .A(in[998]), .B(n768), .Z(n1500) );
  XOR U1425 ( .A(in[167]), .B(in[807]), .Z(n770) );
  XNOR U1426 ( .A(in[1127]), .B(in[487]), .Z(n769) );
  XNOR U1427 ( .A(n770), .B(n769), .Z(n771) );
  XNOR U1428 ( .A(in[1447]), .B(n771), .Z(n1042) );
  XOR U1429 ( .A(n1500), .B(n1042), .Z(n4333) );
  XNOR U1430 ( .A(in[1383]), .B(n4333), .Z(n5011) );
  XOR U1431 ( .A(in[1349]), .B(in[69]), .Z(n773) );
  XNOR U1432 ( .A(in[1029]), .B(in[389]), .Z(n772) );
  XNOR U1433 ( .A(n773), .B(n772), .Z(n774) );
  XNOR U1434 ( .A(in[709]), .B(n774), .Z(n1696) );
  XOR U1435 ( .A(in[1478]), .B(in[518]), .Z(n776) );
  XNOR U1436 ( .A(in[838]), .B(in[198]), .Z(n775) );
  XNOR U1437 ( .A(n776), .B(n775), .Z(n777) );
  XOR U1438 ( .A(in[1158]), .B(n777), .Z(n1415) );
  XOR U1439 ( .A(in[134]), .B(n3177), .Z(n5013) );
  OR U1440 ( .A(n5011), .B(n5013), .Z(n778) );
  XNOR U1441 ( .A(n1607), .B(n778), .Z(out[1027]) );
  XNOR U1442 ( .A(n780), .B(n779), .Z(n3999) );
  XOR U1443 ( .A(in[535]), .B(n3999), .Z(n1611) );
  XOR U1444 ( .A(in[168]), .B(in[1448]), .Z(n782) );
  XNOR U1445 ( .A(in[1128]), .B(in[808]), .Z(n781) );
  XNOR U1446 ( .A(n782), .B(n781), .Z(n783) );
  XNOR U1447 ( .A(in[488]), .B(n783), .Z(n1055) );
  XOR U1448 ( .A(in[39]), .B(in[679]), .Z(n785) );
  XNOR U1449 ( .A(in[359]), .B(in[1319]), .Z(n784) );
  XNOR U1450 ( .A(n785), .B(n784), .Z(n786) );
  XNOR U1451 ( .A(in[999]), .B(n786), .Z(n1505) );
  XOR U1452 ( .A(n1055), .B(n1505), .Z(n4335) );
  XNOR U1453 ( .A(in[1384]), .B(n4335), .Z(n5015) );
  XOR U1454 ( .A(in[1350]), .B(in[70]), .Z(n788) );
  XNOR U1455 ( .A(in[1030]), .B(in[390]), .Z(n787) );
  XNOR U1456 ( .A(n788), .B(n787), .Z(n789) );
  XNOR U1457 ( .A(in[710]), .B(n789), .Z(n1700) );
  XOR U1458 ( .A(in[199]), .B(in[1479]), .Z(n791) );
  XNOR U1459 ( .A(in[1159]), .B(in[839]), .Z(n790) );
  XNOR U1460 ( .A(n791), .B(n790), .Z(n792) );
  XOR U1461 ( .A(in[519]), .B(n792), .Z(n1417) );
  XOR U1462 ( .A(in[135]), .B(n3179), .Z(n5017) );
  OR U1463 ( .A(n5015), .B(n5017), .Z(n793) );
  XNOR U1464 ( .A(n1611), .B(n793), .Z(out[1028]) );
  XNOR U1465 ( .A(n795), .B(n794), .Z(n4003) );
  XOR U1466 ( .A(in[536]), .B(n4003), .Z(n1615) );
  XOR U1467 ( .A(in[169]), .B(in[1449]), .Z(n797) );
  XNOR U1468 ( .A(in[1129]), .B(in[809]), .Z(n796) );
  XNOR U1469 ( .A(n797), .B(n796), .Z(n798) );
  XNOR U1470 ( .A(in[489]), .B(n798), .Z(n1068) );
  XOR U1471 ( .A(in[680]), .B(in[1320]), .Z(n800) );
  XNOR U1472 ( .A(in[40]), .B(in[360]), .Z(n799) );
  XNOR U1473 ( .A(n800), .B(n799), .Z(n801) );
  XNOR U1474 ( .A(in[1000]), .B(n801), .Z(n1509) );
  XOR U1475 ( .A(n1068), .B(n1509), .Z(n4341) );
  XNOR U1476 ( .A(in[1385]), .B(n4341), .Z(n5019) );
  XOR U1477 ( .A(in[1351]), .B(in[711]), .Z(n803) );
  XNOR U1478 ( .A(in[1031]), .B(in[391]), .Z(n802) );
  XNOR U1479 ( .A(n803), .B(n802), .Z(n804) );
  XNOR U1480 ( .A(in[71]), .B(n804), .Z(n1704) );
  XOR U1481 ( .A(in[1480]), .B(in[520]), .Z(n806) );
  XNOR U1482 ( .A(in[840]), .B(in[200]), .Z(n805) );
  XNOR U1483 ( .A(n806), .B(n805), .Z(n807) );
  XOR U1484 ( .A(in[1160]), .B(n807), .Z(n1422) );
  XOR U1485 ( .A(in[136]), .B(n3181), .Z(n5021) );
  OR U1486 ( .A(n5019), .B(n5021), .Z(n808) );
  XNOR U1487 ( .A(n1615), .B(n808), .Z(out[1029]) );
  XOR U1488 ( .A(in[1341]), .B(in[61]), .Z(n810) );
  XNOR U1489 ( .A(in[701]), .B(in[381]), .Z(n809) );
  XNOR U1490 ( .A(n810), .B(n809), .Z(n811) );
  XNOR U1491 ( .A(in[1021]), .B(n811), .Z(n1125) );
  XOR U1492 ( .A(n812), .B(n1125), .Z(n3959) );
  XOR U1493 ( .A(in[637]), .B(n3959), .Z(n2706) );
  IV U1494 ( .A(n2706), .Z(n2795) );
  XOR U1495 ( .A(n814), .B(n813), .Z(n4055) );
  XOR U1496 ( .A(in[228]), .B(n4055), .Z(n3154) );
  XOR U1497 ( .A(in[1512]), .B(in[552]), .Z(n816) );
  XNOR U1498 ( .A(in[872]), .B(in[232]), .Z(n815) );
  XNOR U1499 ( .A(n816), .B(n815), .Z(n817) );
  XNOR U1500 ( .A(in[1192]), .B(n817), .Z(n1514) );
  XNOR U1501 ( .A(n818), .B(n1514), .Z(n4095) );
  IV U1502 ( .A(n4095), .Z(n1274) );
  XOR U1503 ( .A(in[1448]), .B(n1274), .Z(n3152) );
  NANDN U1504 ( .A(n3154), .B(n3152), .Z(n819) );
  XOR U1505 ( .A(n2795), .B(n819), .Z(out[102]) );
  XNOR U1506 ( .A(n821), .B(n820), .Z(n4007) );
  XOR U1507 ( .A(in[537]), .B(n4007), .Z(n1619) );
  XOR U1508 ( .A(in[1352]), .B(in[712]), .Z(n823) );
  XNOR U1509 ( .A(in[1032]), .B(in[392]), .Z(n822) );
  XNOR U1510 ( .A(n823), .B(n822), .Z(n824) );
  XNOR U1511 ( .A(in[72]), .B(n824), .Z(n1709) );
  XOR U1512 ( .A(in[1481]), .B(in[521]), .Z(n826) );
  XNOR U1513 ( .A(in[841]), .B(in[201]), .Z(n825) );
  XNOR U1514 ( .A(n826), .B(n825), .Z(n827) );
  XOR U1515 ( .A(in[1161]), .B(n827), .Z(n1424) );
  XOR U1516 ( .A(in[137]), .B(n3183), .Z(n5025) );
  XOR U1517 ( .A(in[681]), .B(in[1321]), .Z(n829) );
  XNOR U1518 ( .A(in[41]), .B(in[361]), .Z(n828) );
  XNOR U1519 ( .A(n829), .B(n828), .Z(n830) );
  XNOR U1520 ( .A(in[1001]), .B(n830), .Z(n1513) );
  XOR U1521 ( .A(in[170]), .B(in[1450]), .Z(n832) );
  XNOR U1522 ( .A(in[1130]), .B(in[810]), .Z(n831) );
  XNOR U1523 ( .A(n832), .B(n831), .Z(n833) );
  XNOR U1524 ( .A(in[490]), .B(n833), .Z(n1084) );
  XOR U1525 ( .A(n1513), .B(n1084), .Z(n4343) );
  XOR U1526 ( .A(in[1386]), .B(n4343), .Z(n5022) );
  NANDN U1527 ( .A(n5025), .B(n5022), .Z(n834) );
  XNOR U1528 ( .A(n1619), .B(n834), .Z(out[1030]) );
  XOR U1529 ( .A(n836), .B(n835), .Z(n2013) );
  XOR U1530 ( .A(in[538]), .B(n2013), .Z(n1623) );
  XOR U1531 ( .A(in[1353]), .B(in[393]), .Z(n838) );
  XNOR U1532 ( .A(in[713]), .B(in[73]), .Z(n837) );
  XNOR U1533 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U1534 ( .A(in[1033]), .B(n839), .Z(n1713) );
  XOR U1535 ( .A(in[1482]), .B(in[522]), .Z(n841) );
  XNOR U1536 ( .A(in[842]), .B(in[202]), .Z(n840) );
  XNOR U1537 ( .A(n841), .B(n840), .Z(n842) );
  XOR U1538 ( .A(in[1162]), .B(n842), .Z(n1426) );
  XOR U1539 ( .A(in[138]), .B(n3185), .Z(n5029) );
  XOR U1540 ( .A(in[811]), .B(in[491]), .Z(n844) );
  XNOR U1541 ( .A(in[1451]), .B(in[1131]), .Z(n843) );
  XNOR U1542 ( .A(n844), .B(n843), .Z(n845) );
  XNOR U1543 ( .A(in[171]), .B(n845), .Z(n1097) );
  XOR U1544 ( .A(in[682]), .B(in[1322]), .Z(n847) );
  XNOR U1545 ( .A(in[42]), .B(in[362]), .Z(n846) );
  XNOR U1546 ( .A(n847), .B(n846), .Z(n848) );
  XNOR U1547 ( .A(in[1002]), .B(n848), .Z(n1518) );
  XOR U1548 ( .A(n1097), .B(n1518), .Z(n4345) );
  XOR U1549 ( .A(in[1387]), .B(n4345), .Z(n5026) );
  NANDN U1550 ( .A(n5029), .B(n5026), .Z(n849) );
  XNOR U1551 ( .A(n1623), .B(n849), .Z(out[1031]) );
  XOR U1552 ( .A(n851), .B(n850), .Z(n2016) );
  XOR U1553 ( .A(in[539]), .B(n2016), .Z(n1628) );
  XOR U1554 ( .A(in[1354]), .B(in[714]), .Z(n853) );
  XNOR U1555 ( .A(in[74]), .B(in[394]), .Z(n852) );
  XNOR U1556 ( .A(n853), .B(n852), .Z(n854) );
  XNOR U1557 ( .A(in[1034]), .B(n854), .Z(n1717) );
  XOR U1558 ( .A(in[1483]), .B(in[523]), .Z(n856) );
  XNOR U1559 ( .A(in[843]), .B(in[203]), .Z(n855) );
  XNOR U1560 ( .A(n856), .B(n855), .Z(n857) );
  XOR U1561 ( .A(in[1163]), .B(n857), .Z(n1428) );
  XOR U1562 ( .A(n2292), .B(in[139]), .Z(n5033) );
  XOR U1563 ( .A(in[812]), .B(in[492]), .Z(n859) );
  XNOR U1564 ( .A(in[1452]), .B(in[1132]), .Z(n858) );
  XNOR U1565 ( .A(n859), .B(n858), .Z(n860) );
  XNOR U1566 ( .A(in[172]), .B(n860), .Z(n1117) );
  XOR U1567 ( .A(in[683]), .B(in[1323]), .Z(n862) );
  XNOR U1568 ( .A(in[43]), .B(in[363]), .Z(n861) );
  XNOR U1569 ( .A(n862), .B(n861), .Z(n863) );
  XNOR U1570 ( .A(in[1003]), .B(n863), .Z(n1522) );
  XOR U1571 ( .A(n1117), .B(n1522), .Z(n4348) );
  XOR U1572 ( .A(in[1388]), .B(n4348), .Z(n5030) );
  NANDN U1573 ( .A(n5033), .B(n5030), .Z(n864) );
  XNOR U1574 ( .A(n1628), .B(n864), .Z(out[1032]) );
  XOR U1575 ( .A(n866), .B(n865), .Z(n4019) );
  XOR U1576 ( .A(in[540]), .B(n4019), .Z(n1632) );
  XOR U1577 ( .A(in[1355]), .B(in[715]), .Z(n868) );
  XNOR U1578 ( .A(in[1035]), .B(in[395]), .Z(n867) );
  XNOR U1579 ( .A(n868), .B(n867), .Z(n869) );
  XNOR U1580 ( .A(in[75]), .B(n869), .Z(n1721) );
  XOR U1581 ( .A(in[1484]), .B(in[524]), .Z(n871) );
  XNOR U1582 ( .A(in[844]), .B(in[204]), .Z(n870) );
  XNOR U1583 ( .A(n871), .B(n870), .Z(n872) );
  XOR U1584 ( .A(in[1164]), .B(n872), .Z(n1430) );
  XOR U1585 ( .A(in[140]), .B(n3192), .Z(n5037) );
  XOR U1586 ( .A(in[1324]), .B(in[44]), .Z(n874) );
  XNOR U1587 ( .A(in[684]), .B(in[364]), .Z(n873) );
  XNOR U1588 ( .A(n874), .B(n873), .Z(n875) );
  XNOR U1589 ( .A(in[1004]), .B(n875), .Z(n1525) );
  XOR U1590 ( .A(in[813]), .B(in[493]), .Z(n877) );
  XNOR U1591 ( .A(in[1453]), .B(in[1133]), .Z(n876) );
  XNOR U1592 ( .A(n877), .B(n876), .Z(n878) );
  XNOR U1593 ( .A(in[173]), .B(n878), .Z(n1130) );
  XOR U1594 ( .A(n1525), .B(n1130), .Z(n4351) );
  XOR U1595 ( .A(in[1389]), .B(n4351), .Z(n5034) );
  NANDN U1596 ( .A(n5037), .B(n5034), .Z(n879) );
  XNOR U1597 ( .A(n1632), .B(n879), .Z(out[1033]) );
  XOR U1598 ( .A(n881), .B(n880), .Z(n4027) );
  XOR U1599 ( .A(in[541]), .B(n4027), .Z(n1636) );
  XOR U1600 ( .A(in[76]), .B(in[1036]), .Z(n883) );
  XNOR U1601 ( .A(in[716]), .B(in[396]), .Z(n882) );
  XNOR U1602 ( .A(n883), .B(n882), .Z(n884) );
  XNOR U1603 ( .A(in[1356]), .B(n884), .Z(n1725) );
  XOR U1604 ( .A(in[1485]), .B(in[525]), .Z(n886) );
  XNOR U1605 ( .A(in[845]), .B(in[205]), .Z(n885) );
  XNOR U1606 ( .A(n886), .B(n885), .Z(n887) );
  XOR U1607 ( .A(in[1165]), .B(n887), .Z(n1432) );
  XOR U1608 ( .A(in[141]), .B(n3194), .Z(n5045) );
  XOR U1609 ( .A(in[1325]), .B(in[45]), .Z(n889) );
  XNOR U1610 ( .A(in[685]), .B(in[365]), .Z(n888) );
  XNOR U1611 ( .A(n889), .B(n888), .Z(n890) );
  XNOR U1612 ( .A(in[1005]), .B(n890), .Z(n1529) );
  XOR U1613 ( .A(in[814]), .B(in[494]), .Z(n892) );
  XNOR U1614 ( .A(in[1454]), .B(in[1134]), .Z(n891) );
  XNOR U1615 ( .A(n892), .B(n891), .Z(n893) );
  XNOR U1616 ( .A(in[174]), .B(n893), .Z(n1143) );
  XOR U1617 ( .A(n1529), .B(n1143), .Z(n4354) );
  XOR U1618 ( .A(in[1390]), .B(n4354), .Z(n5042) );
  NANDN U1619 ( .A(n5045), .B(n5042), .Z(n894) );
  XNOR U1620 ( .A(n1636), .B(n894), .Z(out[1034]) );
  XOR U1621 ( .A(n896), .B(n895), .Z(n4031) );
  XOR U1622 ( .A(in[542]), .B(n4031), .Z(n1640) );
  XOR U1623 ( .A(in[77]), .B(in[1037]), .Z(n898) );
  XNOR U1624 ( .A(in[717]), .B(in[397]), .Z(n897) );
  XNOR U1625 ( .A(n898), .B(n897), .Z(n899) );
  XNOR U1626 ( .A(in[1357]), .B(n899), .Z(n1729) );
  XOR U1627 ( .A(in[1486]), .B(in[526]), .Z(n901) );
  XNOR U1628 ( .A(in[846]), .B(in[206]), .Z(n900) );
  XNOR U1629 ( .A(n901), .B(n900), .Z(n902) );
  XOR U1630 ( .A(in[1166]), .B(n902), .Z(n1434) );
  XOR U1631 ( .A(in[142]), .B(n3197), .Z(n5049) );
  XOR U1632 ( .A(in[1326]), .B(in[46]), .Z(n904) );
  XNOR U1633 ( .A(in[686]), .B(in[366]), .Z(n903) );
  XNOR U1634 ( .A(n904), .B(n903), .Z(n905) );
  XNOR U1635 ( .A(in[1006]), .B(n905), .Z(n1533) );
  XOR U1636 ( .A(in[815]), .B(in[495]), .Z(n907) );
  XNOR U1637 ( .A(in[1455]), .B(in[1135]), .Z(n906) );
  XNOR U1638 ( .A(n907), .B(n906), .Z(n908) );
  XNOR U1639 ( .A(in[175]), .B(n908), .Z(n1156) );
  XOR U1640 ( .A(n1533), .B(n1156), .Z(n4356) );
  XOR U1641 ( .A(in[1391]), .B(n4356), .Z(n5046) );
  NANDN U1642 ( .A(n5049), .B(n5046), .Z(n909) );
  XNOR U1643 ( .A(n1640), .B(n909), .Z(out[1035]) );
  XOR U1644 ( .A(n911), .B(n910), .Z(n4035) );
  XOR U1645 ( .A(in[543]), .B(n4035), .Z(n1644) );
  XOR U1646 ( .A(in[78]), .B(in[1038]), .Z(n913) );
  XNOR U1647 ( .A(in[718]), .B(in[398]), .Z(n912) );
  XNOR U1648 ( .A(n913), .B(n912), .Z(n914) );
  XNOR U1649 ( .A(in[1358]), .B(n914), .Z(n1733) );
  XOR U1650 ( .A(in[1487]), .B(in[527]), .Z(n916) );
  XNOR U1651 ( .A(in[847]), .B(in[207]), .Z(n915) );
  XNOR U1652 ( .A(n916), .B(n915), .Z(n917) );
  XOR U1653 ( .A(in[1167]), .B(n917), .Z(n1436) );
  XOR U1654 ( .A(in[143]), .B(n3200), .Z(n5053) );
  XOR U1655 ( .A(in[816]), .B(in[496]), .Z(n919) );
  XNOR U1656 ( .A(in[1456]), .B(in[1136]), .Z(n918) );
  XNOR U1657 ( .A(n919), .B(n918), .Z(n920) );
  XNOR U1658 ( .A(in[176]), .B(n920), .Z(n1171) );
  XOR U1659 ( .A(in[1327]), .B(in[47]), .Z(n922) );
  XNOR U1660 ( .A(in[687]), .B(in[367]), .Z(n921) );
  XNOR U1661 ( .A(n922), .B(n921), .Z(n923) );
  XNOR U1662 ( .A(in[1007]), .B(n923), .Z(n1537) );
  XOR U1663 ( .A(n1171), .B(n1537), .Z(n4359) );
  XOR U1664 ( .A(in[1392]), .B(n4359), .Z(n5050) );
  NANDN U1665 ( .A(n5053), .B(n5050), .Z(n924) );
  XNOR U1666 ( .A(n1644), .B(n924), .Z(out[1036]) );
  XOR U1667 ( .A(n926), .B(n925), .Z(n4039) );
  XOR U1668 ( .A(in[544]), .B(n4039), .Z(n1648) );
  XOR U1669 ( .A(in[79]), .B(in[1039]), .Z(n928) );
  XNOR U1670 ( .A(in[719]), .B(in[399]), .Z(n927) );
  XNOR U1671 ( .A(n928), .B(n927), .Z(n929) );
  XNOR U1672 ( .A(in[1359]), .B(n929), .Z(n1737) );
  XOR U1673 ( .A(in[1488]), .B(in[528]), .Z(n931) );
  XNOR U1674 ( .A(in[848]), .B(in[208]), .Z(n930) );
  XNOR U1675 ( .A(n931), .B(n930), .Z(n932) );
  XOR U1676 ( .A(n1737), .B(n230), .Z(n3203) );
  XOR U1677 ( .A(in[144]), .B(n3203), .Z(n5057) );
  XOR U1678 ( .A(in[817]), .B(in[497]), .Z(n934) );
  XNOR U1679 ( .A(in[1457]), .B(in[1137]), .Z(n933) );
  XNOR U1680 ( .A(n934), .B(n933), .Z(n935) );
  XNOR U1681 ( .A(in[177]), .B(n935), .Z(n1186) );
  XOR U1682 ( .A(in[1328]), .B(in[48]), .Z(n937) );
  XNOR U1683 ( .A(in[688]), .B(in[368]), .Z(n936) );
  XNOR U1684 ( .A(n937), .B(n936), .Z(n938) );
  XNOR U1685 ( .A(in[1008]), .B(n938), .Z(n1541) );
  XOR U1686 ( .A(n1186), .B(n1541), .Z(n4362) );
  XOR U1687 ( .A(in[1393]), .B(n4362), .Z(n5054) );
  NANDN U1688 ( .A(n5057), .B(n5054), .Z(n939) );
  XNOR U1689 ( .A(n1648), .B(n939), .Z(out[1037]) );
  XOR U1690 ( .A(n941), .B(n940), .Z(n4043) );
  XOR U1691 ( .A(in[545]), .B(n4043), .Z(n1652) );
  XOR U1692 ( .A(in[80]), .B(in[1040]), .Z(n943) );
  XNOR U1693 ( .A(in[720]), .B(in[400]), .Z(n942) );
  XNOR U1694 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U1695 ( .A(in[1360]), .B(n944), .Z(n1741) );
  XOR U1696 ( .A(in[1489]), .B(in[529]), .Z(n946) );
  XNOR U1697 ( .A(in[849]), .B(in[209]), .Z(n945) );
  XNOR U1698 ( .A(n946), .B(n945), .Z(n947) );
  XOR U1699 ( .A(in[1169]), .B(n947), .Z(n1439) );
  XOR U1700 ( .A(in[145]), .B(n3206), .Z(n5061) );
  XOR U1701 ( .A(in[818]), .B(in[498]), .Z(n949) );
  XNOR U1702 ( .A(in[1458]), .B(in[1138]), .Z(n948) );
  XNOR U1703 ( .A(n949), .B(n948), .Z(n950) );
  XNOR U1704 ( .A(in[178]), .B(n950), .Z(n1201) );
  XOR U1705 ( .A(in[1329]), .B(in[49]), .Z(n952) );
  XNOR U1706 ( .A(in[689]), .B(in[369]), .Z(n951) );
  XNOR U1707 ( .A(n952), .B(n951), .Z(n953) );
  XNOR U1708 ( .A(in[1009]), .B(n953), .Z(n1547) );
  XOR U1709 ( .A(n1201), .B(n1547), .Z(n4365) );
  XOR U1710 ( .A(in[1394]), .B(n4365), .Z(n5058) );
  NANDN U1711 ( .A(n5061), .B(n5058), .Z(n954) );
  XNOR U1712 ( .A(n1652), .B(n954), .Z(out[1038]) );
  IV U1713 ( .A(n4047), .Z(n3393) );
  XOR U1714 ( .A(n3393), .B(in[546]), .Z(n1656) );
  XOR U1715 ( .A(in[81]), .B(in[1041]), .Z(n956) );
  XNOR U1716 ( .A(in[721]), .B(in[401]), .Z(n955) );
  XNOR U1717 ( .A(n956), .B(n955), .Z(n957) );
  XNOR U1718 ( .A(in[1361]), .B(n957), .Z(n1745) );
  XOR U1719 ( .A(in[1490]), .B(in[530]), .Z(n959) );
  XNOR U1720 ( .A(in[850]), .B(in[210]), .Z(n958) );
  XNOR U1721 ( .A(n959), .B(n958), .Z(n960) );
  XOR U1722 ( .A(in[1170]), .B(n960), .Z(n1443) );
  XOR U1723 ( .A(in[146]), .B(n3209), .Z(n5065) );
  XOR U1724 ( .A(in[1330]), .B(in[50]), .Z(n962) );
  XNOR U1725 ( .A(in[690]), .B(in[370]), .Z(n961) );
  XNOR U1726 ( .A(n962), .B(n961), .Z(n963) );
  XNOR U1727 ( .A(in[1010]), .B(n963), .Z(n1551) );
  XOR U1728 ( .A(in[819]), .B(in[499]), .Z(n965) );
  XNOR U1729 ( .A(in[1459]), .B(in[1139]), .Z(n964) );
  XNOR U1730 ( .A(n965), .B(n964), .Z(n966) );
  XNOR U1731 ( .A(in[179]), .B(n966), .Z(n1216) );
  XOR U1732 ( .A(n1551), .B(n1216), .Z(n4372) );
  XOR U1733 ( .A(in[1395]), .B(n4372), .Z(n5062) );
  NANDN U1734 ( .A(n5065), .B(n5062), .Z(n967) );
  XOR U1735 ( .A(n1656), .B(n967), .Z(out[1039]) );
  XOR U1736 ( .A(in[1342]), .B(in[62]), .Z(n969) );
  XNOR U1737 ( .A(in[702]), .B(in[382]), .Z(n968) );
  XNOR U1738 ( .A(n969), .B(n968), .Z(n970) );
  XNOR U1739 ( .A(in[1022]), .B(n970), .Z(n1138) );
  XOR U1740 ( .A(n971), .B(n1138), .Z(n3963) );
  XOR U1741 ( .A(in[638]), .B(n3963), .Z(n2708) );
  IV U1742 ( .A(n2708), .Z(n2797) );
  XOR U1743 ( .A(n973), .B(n972), .Z(n4059) );
  XOR U1744 ( .A(in[229]), .B(n4059), .Z(n3165) );
  XOR U1745 ( .A(in[1513]), .B(in[553]), .Z(n975) );
  XNOR U1746 ( .A(in[873]), .B(in[233]), .Z(n974) );
  XNOR U1747 ( .A(n975), .B(n974), .Z(n976) );
  XNOR U1748 ( .A(in[1193]), .B(n976), .Z(n1517) );
  XNOR U1749 ( .A(n977), .B(n1517), .Z(n4099) );
  IV U1750 ( .A(n4099), .Z(n1286) );
  XOR U1751 ( .A(in[1449]), .B(n1286), .Z(n3162) );
  NANDN U1752 ( .A(n3165), .B(n3162), .Z(n978) );
  XOR U1753 ( .A(n2797), .B(n978), .Z(out[103]) );
  XOR U1754 ( .A(n3396), .B(in[547]), .Z(n1660) );
  XOR U1755 ( .A(in[1042]), .B(in[402]), .Z(n980) );
  XNOR U1756 ( .A(in[722]), .B(in[82]), .Z(n979) );
  XNOR U1757 ( .A(n980), .B(n979), .Z(n981) );
  XNOR U1758 ( .A(in[1362]), .B(n981), .Z(n1750) );
  XOR U1759 ( .A(in[851]), .B(in[1171]), .Z(n983) );
  XNOR U1760 ( .A(in[1491]), .B(in[211]), .Z(n982) );
  XNOR U1761 ( .A(n983), .B(n982), .Z(n984) );
  XOR U1762 ( .A(in[531]), .B(n984), .Z(n1445) );
  IV U1763 ( .A(n3212), .Z(n4004) );
  XNOR U1764 ( .A(in[147]), .B(n4004), .Z(n5068) );
  XOR U1765 ( .A(in[820]), .B(in[500]), .Z(n986) );
  XNOR U1766 ( .A(in[1460]), .B(in[1140]), .Z(n985) );
  XNOR U1767 ( .A(n986), .B(n985), .Z(n987) );
  XNOR U1768 ( .A(in[180]), .B(n987), .Z(n1231) );
  XOR U1769 ( .A(in[1331]), .B(in[51]), .Z(n989) );
  XNOR U1770 ( .A(in[691]), .B(in[371]), .Z(n988) );
  XNOR U1771 ( .A(n989), .B(n988), .Z(n990) );
  XNOR U1772 ( .A(in[1011]), .B(n990), .Z(n1555) );
  XOR U1773 ( .A(n1231), .B(n1555), .Z(n4375) );
  XOR U1774 ( .A(in[1396]), .B(n4375), .Z(n5067) );
  NANDN U1775 ( .A(n5068), .B(n5067), .Z(n991) );
  XOR U1776 ( .A(n1660), .B(n991), .Z(out[1040]) );
  IV U1777 ( .A(n4055), .Z(n3400) );
  XOR U1778 ( .A(n3400), .B(in[548]), .Z(n1664) );
  XOR U1779 ( .A(in[83]), .B(in[1043]), .Z(n993) );
  XNOR U1780 ( .A(in[723]), .B(in[403]), .Z(n992) );
  XNOR U1781 ( .A(n993), .B(n992), .Z(n994) );
  XNOR U1782 ( .A(in[1363]), .B(n994), .Z(n1754) );
  XOR U1783 ( .A(in[852]), .B(in[1172]), .Z(n996) );
  XNOR U1784 ( .A(in[1492]), .B(in[212]), .Z(n995) );
  XNOR U1785 ( .A(n996), .B(n995), .Z(n997) );
  XOR U1786 ( .A(in[532]), .B(n997), .Z(n1447) );
  IV U1787 ( .A(n3215), .Z(n4008) );
  XNOR U1788 ( .A(in[148]), .B(n4008), .Z(n5071) );
  XOR U1789 ( .A(in[821]), .B(in[501]), .Z(n999) );
  XNOR U1790 ( .A(in[1461]), .B(in[1141]), .Z(n998) );
  XNOR U1791 ( .A(n999), .B(n998), .Z(n1000) );
  XNOR U1792 ( .A(in[181]), .B(n1000), .Z(n1246) );
  XOR U1793 ( .A(in[1332]), .B(in[52]), .Z(n1002) );
  XNOR U1794 ( .A(in[692]), .B(in[372]), .Z(n1001) );
  XNOR U1795 ( .A(n1002), .B(n1001), .Z(n1003) );
  XNOR U1796 ( .A(in[1012]), .B(n1003), .Z(n1559) );
  XOR U1797 ( .A(n1246), .B(n1559), .Z(n4378) );
  XOR U1798 ( .A(in[1397]), .B(n4378), .Z(n5070) );
  NANDN U1799 ( .A(n5071), .B(n5070), .Z(n1004) );
  XOR U1800 ( .A(n1664), .B(n1004), .Z(out[1041]) );
  IV U1801 ( .A(n4059), .Z(n3404) );
  XOR U1802 ( .A(n3404), .B(in[549]), .Z(n1669) );
  XOR U1803 ( .A(in[853]), .B(in[1173]), .Z(n1006) );
  XNOR U1804 ( .A(in[1493]), .B(in[213]), .Z(n1005) );
  XNOR U1805 ( .A(n1006), .B(n1005), .Z(n1007) );
  XOR U1806 ( .A(in[533]), .B(n1007), .Z(n1449) );
  IV U1807 ( .A(n2754), .Z(n4012) );
  XNOR U1808 ( .A(in[149]), .B(n4012), .Z(n5074) );
  XOR U1809 ( .A(in[822]), .B(in[502]), .Z(n1010) );
  XNOR U1810 ( .A(in[1462]), .B(in[1142]), .Z(n1009) );
  XNOR U1811 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR U1812 ( .A(in[182]), .B(n1011), .Z(n1261) );
  XOR U1813 ( .A(in[1333]), .B(in[53]), .Z(n1013) );
  XNOR U1814 ( .A(in[693]), .B(in[373]), .Z(n1012) );
  XNOR U1815 ( .A(n1013), .B(n1012), .Z(n1014) );
  XNOR U1816 ( .A(in[1013]), .B(n1014), .Z(n1563) );
  XOR U1817 ( .A(n1261), .B(n1563), .Z(n4381) );
  XOR U1818 ( .A(in[1398]), .B(n4381), .Z(n5073) );
  NANDN U1819 ( .A(n5074), .B(n5073), .Z(n1015) );
  XOR U1820 ( .A(n1669), .B(n1015), .Z(out[1042]) );
  XOR U1821 ( .A(n1017), .B(n1016), .Z(n2035) );
  XOR U1822 ( .A(in[550]), .B(n2035), .Z(n1673) );
  XOR U1823 ( .A(in[854]), .B(in[1174]), .Z(n1019) );
  XNOR U1824 ( .A(in[1494]), .B(in[214]), .Z(n1018) );
  XNOR U1825 ( .A(n1019), .B(n1018), .Z(n1020) );
  XOR U1826 ( .A(in[534]), .B(n1020), .Z(n1451) );
  XOR U1827 ( .A(in[150]), .B(n2771), .Z(n5078) );
  XOR U1828 ( .A(in[823]), .B(in[503]), .Z(n1023) );
  XNOR U1829 ( .A(in[1463]), .B(in[1143]), .Z(n1022) );
  XNOR U1830 ( .A(n1023), .B(n1022), .Z(n1024) );
  XNOR U1831 ( .A(in[183]), .B(n1024), .Z(n1273) );
  XOR U1832 ( .A(in[1334]), .B(in[54]), .Z(n1026) );
  XNOR U1833 ( .A(in[694]), .B(in[374]), .Z(n1025) );
  XNOR U1834 ( .A(n1026), .B(n1025), .Z(n1027) );
  XNOR U1835 ( .A(in[1014]), .B(n1027), .Z(n1567) );
  XOR U1836 ( .A(n1273), .B(n1567), .Z(n4384) );
  XOR U1837 ( .A(in[1399]), .B(n4384), .Z(n5075) );
  NANDN U1838 ( .A(n5078), .B(n5075), .Z(n1028) );
  XNOR U1839 ( .A(n1673), .B(n1028), .Z(out[1043]) );
  XOR U1840 ( .A(n1030), .B(n1029), .Z(n2038) );
  XOR U1841 ( .A(in[551]), .B(n2038), .Z(n1677) );
  XOR U1842 ( .A(in[855]), .B(in[1175]), .Z(n1032) );
  XNOR U1843 ( .A(in[1495]), .B(in[215]), .Z(n1031) );
  XNOR U1844 ( .A(n1032), .B(n1031), .Z(n1033) );
  XOR U1845 ( .A(in[535]), .B(n1033), .Z(n1453) );
  XOR U1846 ( .A(in[151]), .B(n2778), .Z(n5085) );
  XOR U1847 ( .A(in[824]), .B(in[504]), .Z(n1036) );
  XNOR U1848 ( .A(in[1464]), .B(in[1144]), .Z(n1035) );
  XNOR U1849 ( .A(n1036), .B(n1035), .Z(n1037) );
  XNOR U1850 ( .A(in[184]), .B(n1037), .Z(n1279) );
  XOR U1851 ( .A(in[1335]), .B(in[55]), .Z(n1039) );
  XNOR U1852 ( .A(in[695]), .B(in[375]), .Z(n1038) );
  XNOR U1853 ( .A(n1039), .B(n1038), .Z(n1040) );
  XNOR U1854 ( .A(in[1015]), .B(n1040), .Z(n1571) );
  XOR U1855 ( .A(n1279), .B(n1571), .Z(n4386) );
  XOR U1856 ( .A(in[1400]), .B(n4386), .Z(n5084) );
  NANDN U1857 ( .A(n5085), .B(n5084), .Z(n1041) );
  XNOR U1858 ( .A(n1677), .B(n1041), .Z(out[1044]) );
  XOR U1859 ( .A(n1043), .B(n1042), .Z(n2042) );
  XOR U1860 ( .A(in[552]), .B(n2042), .Z(n1681) );
  XOR U1861 ( .A(in[856]), .B(in[1176]), .Z(n1045) );
  XNOR U1862 ( .A(in[1496]), .B(in[216]), .Z(n1044) );
  XNOR U1863 ( .A(n1045), .B(n1044), .Z(n1046) );
  XOR U1864 ( .A(in[536]), .B(n1046), .Z(n1457) );
  XOR U1865 ( .A(in[152]), .B(n2792), .Z(n5088) );
  XOR U1866 ( .A(in[825]), .B(in[505]), .Z(n1049) );
  XNOR U1867 ( .A(in[1465]), .B(in[1145]), .Z(n1048) );
  XNOR U1868 ( .A(n1049), .B(n1048), .Z(n1050) );
  XNOR U1869 ( .A(in[185]), .B(n1050), .Z(n1291) );
  XOR U1870 ( .A(in[1336]), .B(in[56]), .Z(n1052) );
  XNOR U1871 ( .A(in[696]), .B(in[376]), .Z(n1051) );
  XNOR U1872 ( .A(n1052), .B(n1051), .Z(n1053) );
  XNOR U1873 ( .A(in[1016]), .B(n1053), .Z(n1575) );
  XOR U1874 ( .A(n1291), .B(n1575), .Z(n4389) );
  XOR U1875 ( .A(in[1401]), .B(n4389), .Z(n5087) );
  NANDN U1876 ( .A(n5088), .B(n5087), .Z(n1054) );
  XNOR U1877 ( .A(n1681), .B(n1054), .Z(out[1045]) );
  XOR U1878 ( .A(n1056), .B(n1055), .Z(n2044) );
  XOR U1879 ( .A(in[553]), .B(n2044), .Z(n1685) );
  XOR U1880 ( .A(in[857]), .B(in[1177]), .Z(n1058) );
  XNOR U1881 ( .A(in[1497]), .B(in[217]), .Z(n1057) );
  XNOR U1882 ( .A(n1058), .B(n1057), .Z(n1059) );
  XOR U1883 ( .A(in[537]), .B(n1059), .Z(n1459) );
  XOR U1884 ( .A(in[153]), .B(n2815), .Z(n5091) );
  XOR U1885 ( .A(in[1337]), .B(in[57]), .Z(n1062) );
  XNOR U1886 ( .A(in[697]), .B(in[377]), .Z(n1061) );
  XNOR U1887 ( .A(n1062), .B(n1061), .Z(n1063) );
  XNOR U1888 ( .A(in[1017]), .B(n1063), .Z(n1579) );
  XOR U1889 ( .A(in[826]), .B(in[506]), .Z(n1065) );
  XNOR U1890 ( .A(in[1466]), .B(in[1146]), .Z(n1064) );
  XNOR U1891 ( .A(n1065), .B(n1064), .Z(n1066) );
  XNOR U1892 ( .A(in[186]), .B(n1066), .Z(n1303) );
  XOR U1893 ( .A(n1579), .B(n1303), .Z(n2114) );
  IV U1894 ( .A(n2114), .Z(n4392) );
  XNOR U1895 ( .A(in[1402]), .B(n4392), .Z(n5090) );
  NANDN U1896 ( .A(n5091), .B(n5090), .Z(n1067) );
  XNOR U1897 ( .A(n1685), .B(n1067), .Z(out[1046]) );
  XOR U1898 ( .A(n1069), .B(n1068), .Z(n2046) );
  XOR U1899 ( .A(in[554]), .B(n2046), .Z(n1689) );
  XOR U1900 ( .A(in[858]), .B(in[1178]), .Z(n1071) );
  XNOR U1901 ( .A(in[1498]), .B(in[218]), .Z(n1070) );
  XNOR U1902 ( .A(n1071), .B(n1070), .Z(n1072) );
  XOR U1903 ( .A(in[538]), .B(n1072), .Z(n1461) );
  XOR U1904 ( .A(in[154]), .B(n2838), .Z(n5094) );
  XOR U1905 ( .A(in[1338]), .B(in[58]), .Z(n1075) );
  XNOR U1906 ( .A(in[698]), .B(in[378]), .Z(n1074) );
  XNOR U1907 ( .A(n1075), .B(n1074), .Z(n1076) );
  XNOR U1908 ( .A(in[1018]), .B(n1076), .Z(n1583) );
  XOR U1909 ( .A(in[827]), .B(in[507]), .Z(n1078) );
  XNOR U1910 ( .A(in[1467]), .B(in[1147]), .Z(n1077) );
  XNOR U1911 ( .A(n1078), .B(n1077), .Z(n1079) );
  XNOR U1912 ( .A(in[187]), .B(n1079), .Z(n1307) );
  XOR U1913 ( .A(n1583), .B(n1307), .Z(n2116) );
  IV U1914 ( .A(n2116), .Z(n4395) );
  XNOR U1915 ( .A(in[1403]), .B(n4395), .Z(n5093) );
  NANDN U1916 ( .A(n5094), .B(n5093), .Z(n1080) );
  XNOR U1917 ( .A(n1689), .B(n1080), .Z(out[1047]) );
  XOR U1918 ( .A(in[1579]), .B(in[619]), .Z(n1082) );
  XNOR U1919 ( .A(in[939]), .B(in[299]), .Z(n1081) );
  XNOR U1920 ( .A(n1082), .B(n1081), .Z(n1083) );
  XNOR U1921 ( .A(in[1259]), .B(n1083), .Z(n1593) );
  XNOR U1922 ( .A(n1084), .B(n1593), .Z(n3428) );
  IV U1923 ( .A(n3428), .Z(n4088) );
  XOR U1924 ( .A(in[555]), .B(n4088), .Z(n1693) );
  XOR U1925 ( .A(in[859]), .B(in[1179]), .Z(n1086) );
  XNOR U1926 ( .A(in[1499]), .B(in[219]), .Z(n1085) );
  XNOR U1927 ( .A(n1086), .B(n1085), .Z(n1087) );
  XOR U1928 ( .A(in[539]), .B(n1087), .Z(n1465) );
  XOR U1929 ( .A(in[155]), .B(n2862), .Z(n5097) );
  XOR U1930 ( .A(in[828]), .B(in[508]), .Z(n1090) );
  XNOR U1931 ( .A(in[1468]), .B(in[1148]), .Z(n1089) );
  XNOR U1932 ( .A(n1090), .B(n1089), .Z(n1091) );
  XNOR U1933 ( .A(in[188]), .B(n1091), .Z(n1311) );
  XOR U1934 ( .A(n1092), .B(n1311), .Z(n4398) );
  XOR U1935 ( .A(in[1404]), .B(n4398), .Z(n5096) );
  NANDN U1936 ( .A(n5097), .B(n5096), .Z(n1093) );
  XNOR U1937 ( .A(n1693), .B(n1093), .Z(out[1048]) );
  XOR U1938 ( .A(in[1580]), .B(in[620]), .Z(n1095) );
  XNOR U1939 ( .A(in[940]), .B(in[300]), .Z(n1094) );
  XNOR U1940 ( .A(n1095), .B(n1094), .Z(n1096) );
  XNOR U1941 ( .A(in[1260]), .B(n1096), .Z(n1597) );
  XNOR U1942 ( .A(n1097), .B(n1597), .Z(n3431) );
  IV U1943 ( .A(n3431), .Z(n4092) );
  XOR U1944 ( .A(in[556]), .B(n4092), .Z(n1697) );
  XOR U1945 ( .A(in[860]), .B(in[1180]), .Z(n1099) );
  XNOR U1946 ( .A(in[1500]), .B(in[220]), .Z(n1098) );
  XNOR U1947 ( .A(n1099), .B(n1098), .Z(n1100) );
  XOR U1948 ( .A(in[540]), .B(n1100), .Z(n1471) );
  XOR U1949 ( .A(in[156]), .B(n2886), .Z(n5100) );
  XOR U1950 ( .A(n1103), .B(n1102), .Z(n4405) );
  XOR U1951 ( .A(in[1405]), .B(n4405), .Z(n5099) );
  NANDN U1952 ( .A(n5100), .B(n5099), .Z(n1104) );
  XNOR U1953 ( .A(n1697), .B(n1104), .Z(out[1049]) );
  XOR U1954 ( .A(in[1343]), .B(in[63]), .Z(n1106) );
  XNOR U1955 ( .A(in[703]), .B(in[383]), .Z(n1105) );
  XNOR U1956 ( .A(n1106), .B(n1105), .Z(n1107) );
  XNOR U1957 ( .A(in[1023]), .B(n1107), .Z(n1151) );
  XOR U1958 ( .A(n1108), .B(n1151), .Z(n3967) );
  XOR U1959 ( .A(in[639]), .B(n3967), .Z(n2710) );
  IV U1960 ( .A(n2710), .Z(n2799) );
  XNOR U1961 ( .A(in[230]), .B(n2035), .Z(n3190) );
  XOR U1962 ( .A(in[874]), .B(in[1194]), .Z(n1110) );
  XNOR U1963 ( .A(in[1514]), .B(in[234]), .Z(n1109) );
  XNOR U1964 ( .A(n1110), .B(n1109), .Z(n1111) );
  XNOR U1965 ( .A(in[554]), .B(n1111), .Z(n1521) );
  XNOR U1966 ( .A(n1112), .B(n1521), .Z(n4103) );
  IV U1967 ( .A(n4103), .Z(n1292) );
  XOR U1968 ( .A(in[1450]), .B(n1292), .Z(n3187) );
  NAND U1969 ( .A(n3190), .B(n3187), .Z(n1113) );
  XOR U1970 ( .A(n2799), .B(n1113), .Z(out[104]) );
  XOR U1971 ( .A(in[1581]), .B(in[621]), .Z(n1115) );
  XNOR U1972 ( .A(in[941]), .B(in[301]), .Z(n1114) );
  XNOR U1973 ( .A(n1115), .B(n1114), .Z(n1116) );
  XNOR U1974 ( .A(in[1261]), .B(n1116), .Z(n1601) );
  XNOR U1975 ( .A(n1117), .B(n1601), .Z(n3434) );
  IV U1976 ( .A(n3434), .Z(n4096) );
  XOR U1977 ( .A(in[557]), .B(n4096), .Z(n1701) );
  XOR U1978 ( .A(in[861]), .B(in[1181]), .Z(n1119) );
  XNOR U1979 ( .A(in[1501]), .B(in[221]), .Z(n1118) );
  XNOR U1980 ( .A(n1119), .B(n1118), .Z(n1120) );
  XOR U1981 ( .A(in[541]), .B(n1120), .Z(n1475) );
  XOR U1982 ( .A(in[157]), .B(n2919), .Z(n5103) );
  XOR U1983 ( .A(in[830]), .B(in[510]), .Z(n1123) );
  XNOR U1984 ( .A(in[1470]), .B(in[1150]), .Z(n1122) );
  XNOR U1985 ( .A(n1123), .B(n1122), .Z(n1124) );
  XNOR U1986 ( .A(in[190]), .B(n1124), .Z(n1315) );
  XOR U1987 ( .A(n1125), .B(n1315), .Z(n4408) );
  XOR U1988 ( .A(in[1406]), .B(n4408), .Z(n5102) );
  NANDN U1989 ( .A(n5103), .B(n5102), .Z(n1126) );
  XNOR U1990 ( .A(n1701), .B(n1126), .Z(out[1050]) );
  XOR U1991 ( .A(in[1582]), .B(in[622]), .Z(n1128) );
  XNOR U1992 ( .A(in[942]), .B(in[302]), .Z(n1127) );
  XNOR U1993 ( .A(n1128), .B(n1127), .Z(n1129) );
  XNOR U1994 ( .A(in[1262]), .B(n1129), .Z(n1605) );
  XNOR U1995 ( .A(n1130), .B(n1605), .Z(n3437) );
  IV U1996 ( .A(n3437), .Z(n4100) );
  XOR U1997 ( .A(in[558]), .B(n4100), .Z(n1705) );
  XOR U1998 ( .A(in[862]), .B(in[1182]), .Z(n1132) );
  XNOR U1999 ( .A(in[1502]), .B(in[222]), .Z(n1131) );
  XNOR U2000 ( .A(n1132), .B(n1131), .Z(n1133) );
  XOR U2001 ( .A(in[542]), .B(n1133), .Z(n1479) );
  XNOR U2002 ( .A(in[158]), .B(n4052), .Z(n1455) );
  IV U2003 ( .A(n1455), .Z(n5106) );
  XOR U2004 ( .A(in[831]), .B(in[511]), .Z(n1136) );
  XNOR U2005 ( .A(in[1471]), .B(in[1151]), .Z(n1135) );
  XNOR U2006 ( .A(n1136), .B(n1135), .Z(n1137) );
  XNOR U2007 ( .A(in[191]), .B(n1137), .Z(n1319) );
  XOR U2008 ( .A(n1138), .B(n1319), .Z(n4411) );
  XOR U2009 ( .A(in[1407]), .B(n4411), .Z(n5105) );
  NANDN U2010 ( .A(n5106), .B(n5105), .Z(n1139) );
  XNOR U2011 ( .A(n1705), .B(n1139), .Z(out[1051]) );
  XOR U2012 ( .A(in[1583]), .B(in[623]), .Z(n1141) );
  XNOR U2013 ( .A(in[943]), .B(in[303]), .Z(n1140) );
  XNOR U2014 ( .A(n1141), .B(n1140), .Z(n1142) );
  XNOR U2015 ( .A(in[1263]), .B(n1142), .Z(n1609) );
  XNOR U2016 ( .A(n1143), .B(n1609), .Z(n3440) );
  IV U2017 ( .A(n3440), .Z(n4104) );
  XOR U2018 ( .A(in[559]), .B(n4104), .Z(n1710) );
  XOR U2019 ( .A(in[863]), .B(in[1183]), .Z(n1145) );
  XNOR U2020 ( .A(in[1503]), .B(in[223]), .Z(n1144) );
  XNOR U2021 ( .A(n1145), .B(n1144), .Z(n1146) );
  XOR U2022 ( .A(in[543]), .B(n1146), .Z(n1481) );
  XOR U2023 ( .A(in[159]), .B(n4056), .Z(n5110) );
  XOR U2024 ( .A(in[768]), .B(in[1088]), .Z(n1149) );
  XNOR U2025 ( .A(in[448]), .B(in[1408]), .Z(n1148) );
  XNOR U2026 ( .A(n1149), .B(n1148), .Z(n1150) );
  XNOR U2027 ( .A(in[128]), .B(n1150), .Z(n1326) );
  XOR U2028 ( .A(n1151), .B(n1326), .Z(n4414) );
  XOR U2029 ( .A(in[1344]), .B(n4414), .Z(n5107) );
  NANDN U2030 ( .A(n5110), .B(n5107), .Z(n1152) );
  XNOR U2031 ( .A(n1710), .B(n1152), .Z(out[1052]) );
  XOR U2032 ( .A(in[1584]), .B(in[624]), .Z(n1154) );
  XNOR U2033 ( .A(in[944]), .B(in[304]), .Z(n1153) );
  XNOR U2034 ( .A(n1154), .B(n1153), .Z(n1155) );
  XNOR U2035 ( .A(in[1264]), .B(n1155), .Z(n1613) );
  XNOR U2036 ( .A(n1156), .B(n1613), .Z(n3443) );
  IV U2037 ( .A(n3443), .Z(n4108) );
  XOR U2038 ( .A(in[560]), .B(n4108), .Z(n1714) );
  XOR U2039 ( .A(in[224]), .B(in[864]), .Z(n1158) );
  XNOR U2040 ( .A(in[1184]), .B(in[1504]), .Z(n1157) );
  XNOR U2041 ( .A(n1158), .B(n1157), .Z(n1159) );
  XOR U2042 ( .A(in[544]), .B(n1159), .Z(n1484) );
  XOR U2043 ( .A(in[160]), .B(n4060), .Z(n5113) );
  XOR U2044 ( .A(in[769]), .B(in[1089]), .Z(n1162) );
  XNOR U2045 ( .A(in[449]), .B(in[1409]), .Z(n1161) );
  XNOR U2046 ( .A(n1162), .B(n1161), .Z(n1163) );
  XNOR U2047 ( .A(in[129]), .B(n1163), .Z(n1330) );
  XOR U2048 ( .A(in[1280]), .B(in[640]), .Z(n1165) );
  XNOR U2049 ( .A(in[960]), .B(in[320]), .Z(n1164) );
  XNOR U2050 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U2051 ( .A(in[0]), .B(n1166), .Z(n1255) );
  XOR U2052 ( .A(n1330), .B(n1255), .Z(n4417) );
  XOR U2053 ( .A(in[1345]), .B(n4417), .Z(n5112) );
  NANDN U2054 ( .A(n5113), .B(n5112), .Z(n1167) );
  XNOR U2055 ( .A(n1714), .B(n1167), .Z(out[1053]) );
  XOR U2056 ( .A(in[1585]), .B(in[625]), .Z(n1169) );
  XNOR U2057 ( .A(in[945]), .B(in[305]), .Z(n1168) );
  XNOR U2058 ( .A(n1169), .B(n1168), .Z(n1170) );
  XNOR U2059 ( .A(in[1265]), .B(n1170), .Z(n1617) );
  XNOR U2060 ( .A(n1171), .B(n1617), .Z(n3446) );
  IV U2061 ( .A(n3446), .Z(n4116) );
  XOR U2062 ( .A(in[561]), .B(n4116), .Z(n1718) );
  XOR U2063 ( .A(in[225]), .B(in[865]), .Z(n1173) );
  XNOR U2064 ( .A(in[1185]), .B(in[1505]), .Z(n1172) );
  XNOR U2065 ( .A(n1173), .B(n1172), .Z(n1174) );
  XOR U2066 ( .A(n1175), .B(n231), .Z(n4064) );
  XNOR U2067 ( .A(in[161]), .B(n4064), .Z(n1463) );
  IV U2068 ( .A(n1463), .Z(n5120) );
  XOR U2069 ( .A(in[1]), .B(in[641]), .Z(n1177) );
  XNOR U2070 ( .A(in[961]), .B(in[321]), .Z(n1176) );
  XNOR U2071 ( .A(n1177), .B(n1176), .Z(n1178) );
  XNOR U2072 ( .A(in[1281]), .B(n1178), .Z(n1320) );
  XOR U2073 ( .A(in[1090]), .B(in[450]), .Z(n1180) );
  XNOR U2074 ( .A(in[130]), .B(in[770]), .Z(n1179) );
  XNOR U2075 ( .A(n1180), .B(n1179), .Z(n1181) );
  XNOR U2076 ( .A(in[1410]), .B(n1181), .Z(n1334) );
  XOR U2077 ( .A(n1320), .B(n1334), .Z(n4420) );
  XOR U2078 ( .A(in[1346]), .B(n4420), .Z(n5119) );
  NANDN U2079 ( .A(n5120), .B(n5119), .Z(n1182) );
  XNOR U2080 ( .A(n1718), .B(n1182), .Z(out[1054]) );
  XOR U2081 ( .A(in[1586]), .B(in[626]), .Z(n1184) );
  XNOR U2082 ( .A(in[946]), .B(in[306]), .Z(n1183) );
  XNOR U2083 ( .A(n1184), .B(n1183), .Z(n1185) );
  XNOR U2084 ( .A(in[1266]), .B(n1185), .Z(n1621) );
  XNOR U2085 ( .A(n1186), .B(n1621), .Z(n3449) );
  IV U2086 ( .A(n3449), .Z(n4120) );
  XOR U2087 ( .A(in[562]), .B(n4120), .Z(n1722) );
  XOR U2088 ( .A(in[1186]), .B(in[1506]), .Z(n1188) );
  XNOR U2089 ( .A(in[546]), .B(in[866]), .Z(n1187) );
  XNOR U2090 ( .A(n1188), .B(n1187), .Z(n1189) );
  XOR U2091 ( .A(in[226]), .B(n1189), .Z(n1489) );
  XNOR U2092 ( .A(in[162]), .B(n4072), .Z(n1467) );
  IV U2093 ( .A(n1467), .Z(n5124) );
  XOR U2094 ( .A(in[2]), .B(in[642]), .Z(n1192) );
  XNOR U2095 ( .A(in[962]), .B(in[322]), .Z(n1191) );
  XNOR U2096 ( .A(n1192), .B(n1191), .Z(n1193) );
  XNOR U2097 ( .A(in[1282]), .B(n1193), .Z(n1365) );
  XOR U2098 ( .A(in[771]), .B(in[1091]), .Z(n1195) );
  XNOR U2099 ( .A(in[451]), .B(in[1411]), .Z(n1194) );
  XNOR U2100 ( .A(n1195), .B(n1194), .Z(n1196) );
  XNOR U2101 ( .A(in[131]), .B(n1196), .Z(n1338) );
  XOR U2102 ( .A(n1365), .B(n1338), .Z(n4423) );
  XOR U2103 ( .A(in[1347]), .B(n4423), .Z(n5121) );
  NANDN U2104 ( .A(n5124), .B(n5121), .Z(n1197) );
  XNOR U2105 ( .A(n1722), .B(n1197), .Z(out[1055]) );
  XOR U2106 ( .A(in[1587]), .B(in[627]), .Z(n1199) );
  XNOR U2107 ( .A(in[947]), .B(in[307]), .Z(n1198) );
  XNOR U2108 ( .A(n1199), .B(n1198), .Z(n1200) );
  XNOR U2109 ( .A(in[1267]), .B(n1200), .Z(n1626) );
  XNOR U2110 ( .A(n1201), .B(n1626), .Z(n3452) );
  IV U2111 ( .A(n3452), .Z(n4124) );
  XOR U2112 ( .A(in[563]), .B(n4124), .Z(n1726) );
  XOR U2113 ( .A(in[1187]), .B(in[1507]), .Z(n1203) );
  XNOR U2114 ( .A(in[547]), .B(in[867]), .Z(n1202) );
  XNOR U2115 ( .A(n1203), .B(n1202), .Z(n1204) );
  XOR U2116 ( .A(in[227]), .B(n1204), .Z(n1492) );
  XNOR U2117 ( .A(in[163]), .B(n4076), .Z(n1473) );
  IV U2118 ( .A(n1473), .Z(n5128) );
  XOR U2119 ( .A(in[772]), .B(in[1092]), .Z(n1207) );
  XNOR U2120 ( .A(in[452]), .B(in[1412]), .Z(n1206) );
  XNOR U2121 ( .A(n1207), .B(n1206), .Z(n1208) );
  XNOR U2122 ( .A(in[132]), .B(n1208), .Z(n1342) );
  XOR U2123 ( .A(in[323]), .B(in[643]), .Z(n1210) );
  XNOR U2124 ( .A(in[963]), .B(in[3]), .Z(n1209) );
  XNOR U2125 ( .A(n1210), .B(n1209), .Z(n1211) );
  XNOR U2126 ( .A(in[1283]), .B(n1211), .Z(n1406) );
  XOR U2127 ( .A(n1342), .B(n1406), .Z(n4426) );
  XOR U2128 ( .A(in[1348]), .B(n4426), .Z(n5125) );
  NANDN U2129 ( .A(n5128), .B(n5125), .Z(n1212) );
  XNOR U2130 ( .A(n1726), .B(n1212), .Z(out[1056]) );
  XOR U2131 ( .A(in[1588]), .B(in[628]), .Z(n1214) );
  XNOR U2132 ( .A(in[948]), .B(in[308]), .Z(n1213) );
  XNOR U2133 ( .A(n1214), .B(n1213), .Z(n1215) );
  XNOR U2134 ( .A(in[1268]), .B(n1215), .Z(n1630) );
  XNOR U2135 ( .A(n1216), .B(n1630), .Z(n3459) );
  IV U2136 ( .A(n3459), .Z(n4128) );
  XOR U2137 ( .A(in[564]), .B(n4128), .Z(n1730) );
  XOR U2138 ( .A(in[1188]), .B(in[1508]), .Z(n1218) );
  XNOR U2139 ( .A(in[548]), .B(in[868]), .Z(n1217) );
  XNOR U2140 ( .A(n1218), .B(n1217), .Z(n1219) );
  XNOR U2141 ( .A(in[228]), .B(n1219), .Z(n1495) );
  XNOR U2142 ( .A(in[164]), .B(n4080), .Z(n1477) );
  IV U2143 ( .A(n1477), .Z(n5132) );
  XOR U2144 ( .A(in[324]), .B(in[644]), .Z(n1222) );
  XNOR U2145 ( .A(in[964]), .B(in[4]), .Z(n1221) );
  XNOR U2146 ( .A(n1222), .B(n1221), .Z(n1223) );
  XNOR U2147 ( .A(in[1284]), .B(n1223), .Z(n1410) );
  XOR U2148 ( .A(in[773]), .B(in[1093]), .Z(n1225) );
  XNOR U2149 ( .A(in[453]), .B(in[1413]), .Z(n1224) );
  XNOR U2150 ( .A(n1225), .B(n1224), .Z(n1226) );
  XNOR U2151 ( .A(in[133]), .B(n1226), .Z(n1346) );
  XOR U2152 ( .A(n1410), .B(n1346), .Z(n4429) );
  XOR U2153 ( .A(in[1349]), .B(n4429), .Z(n5129) );
  NANDN U2154 ( .A(n5132), .B(n5129), .Z(n1227) );
  XNOR U2155 ( .A(n1730), .B(n1227), .Z(out[1057]) );
  XOR U2156 ( .A(in[1589]), .B(in[629]), .Z(n1229) );
  XNOR U2157 ( .A(in[949]), .B(in[309]), .Z(n1228) );
  XNOR U2158 ( .A(n1229), .B(n1228), .Z(n1230) );
  XNOR U2159 ( .A(in[1269]), .B(n1230), .Z(n1634) );
  XNOR U2160 ( .A(n1231), .B(n1634), .Z(n3462) );
  IV U2161 ( .A(n3462), .Z(n4132) );
  XOR U2162 ( .A(in[565]), .B(n4132), .Z(n1734) );
  XOR U2163 ( .A(in[1189]), .B(in[1509]), .Z(n1233) );
  XNOR U2164 ( .A(in[549]), .B(in[869]), .Z(n1232) );
  XNOR U2165 ( .A(n1233), .B(n1232), .Z(n1234) );
  XOR U2166 ( .A(in[229]), .B(n1234), .Z(n1499) );
  XOR U2167 ( .A(in[165]), .B(n2211), .Z(n5136) );
  XOR U2168 ( .A(in[774]), .B(in[1094]), .Z(n1237) );
  XNOR U2169 ( .A(in[454]), .B(in[1414]), .Z(n1236) );
  XNOR U2170 ( .A(n1237), .B(n1236), .Z(n1238) );
  XNOR U2171 ( .A(in[134]), .B(n1238), .Z(n1350) );
  XOR U2172 ( .A(in[325]), .B(in[645]), .Z(n1240) );
  XNOR U2173 ( .A(in[965]), .B(in[5]), .Z(n1239) );
  XNOR U2174 ( .A(n1240), .B(n1239), .Z(n1241) );
  XNOR U2175 ( .A(in[1285]), .B(n1241), .Z(n1412) );
  XOR U2176 ( .A(n1350), .B(n1412), .Z(n2126) );
  IV U2177 ( .A(n2126), .Z(n4432) );
  XNOR U2178 ( .A(in[1350]), .B(n4432), .Z(n5133) );
  NANDN U2179 ( .A(n5136), .B(n5133), .Z(n1242) );
  XNOR U2180 ( .A(n1734), .B(n1242), .Z(out[1058]) );
  XOR U2181 ( .A(in[1590]), .B(in[630]), .Z(n1244) );
  XNOR U2182 ( .A(in[950]), .B(in[310]), .Z(n1243) );
  XNOR U2183 ( .A(n1244), .B(n1243), .Z(n1245) );
  XNOR U2184 ( .A(in[1270]), .B(n1245), .Z(n1638) );
  XNOR U2185 ( .A(n1246), .B(n1638), .Z(n3258) );
  IV U2186 ( .A(n3258), .Z(n4136) );
  XOR U2187 ( .A(in[566]), .B(n4136), .Z(n1738) );
  XNOR U2188 ( .A(in[166]), .B(n1247), .Z(n5140) );
  XOR U2189 ( .A(in[775]), .B(in[1095]), .Z(n1249) );
  XNOR U2190 ( .A(in[455]), .B(in[1415]), .Z(n1248) );
  XNOR U2191 ( .A(n1249), .B(n1248), .Z(n1250) );
  XNOR U2192 ( .A(in[135]), .B(n1250), .Z(n1354) );
  XOR U2193 ( .A(in[326]), .B(in[6]), .Z(n1252) );
  XNOR U2194 ( .A(in[966]), .B(in[646]), .Z(n1251) );
  XNOR U2195 ( .A(n1252), .B(n1251), .Z(n1253) );
  XNOR U2196 ( .A(in[1286]), .B(n1253), .Z(n1414) );
  XOR U2197 ( .A(n1354), .B(n1414), .Z(n4443) );
  XOR U2198 ( .A(in[1351]), .B(n4443), .Z(n5137) );
  NAND U2199 ( .A(n5140), .B(n5137), .Z(n1254) );
  XNOR U2200 ( .A(n1738), .B(n1254), .Z(out[1059]) );
  XOR U2201 ( .A(n1256), .B(n1255), .Z(n3971) );
  XOR U2202 ( .A(in[576]), .B(n3971), .Z(n2712) );
  IV U2203 ( .A(n2712), .Z(n2801) );
  XNOR U2204 ( .A(in[1451]), .B(n4107), .Z(n3219) );
  XNOR U2205 ( .A(in[231]), .B(n2038), .Z(n3221) );
  NANDN U2206 ( .A(n3219), .B(n3221), .Z(n1257) );
  XOR U2207 ( .A(n2801), .B(n1257), .Z(out[105]) );
  XOR U2208 ( .A(in[1591]), .B(in[631]), .Z(n1259) );
  XNOR U2209 ( .A(in[951]), .B(in[311]), .Z(n1258) );
  XNOR U2210 ( .A(n1259), .B(n1258), .Z(n1260) );
  XNOR U2211 ( .A(in[1271]), .B(n1260), .Z(n1642) );
  XNOR U2212 ( .A(n1261), .B(n1642), .Z(n3261) );
  IV U2213 ( .A(n3261), .Z(n4140) );
  XOR U2214 ( .A(in[567]), .B(n4140), .Z(n1742) );
  XNOR U2215 ( .A(in[167]), .B(n1262), .Z(n5144) );
  XOR U2216 ( .A(in[776]), .B(in[1096]), .Z(n1264) );
  XNOR U2217 ( .A(in[456]), .B(in[1416]), .Z(n1263) );
  XNOR U2218 ( .A(n1264), .B(n1263), .Z(n1265) );
  XNOR U2219 ( .A(in[136]), .B(n1265), .Z(n1358) );
  XOR U2220 ( .A(in[327]), .B(in[7]), .Z(n1267) );
  XNOR U2221 ( .A(in[967]), .B(in[647]), .Z(n1266) );
  XNOR U2222 ( .A(n1267), .B(n1266), .Z(n1268) );
  XNOR U2223 ( .A(in[1287]), .B(n1268), .Z(n1416) );
  XOR U2224 ( .A(n1358), .B(n1416), .Z(n4446) );
  XOR U2225 ( .A(in[1352]), .B(n4446), .Z(n5141) );
  NAND U2226 ( .A(n5144), .B(n5141), .Z(n1269) );
  XNOR U2227 ( .A(n1742), .B(n1269), .Z(out[1060]) );
  XOR U2228 ( .A(in[632]), .B(in[1592]), .Z(n1271) );
  XNOR U2229 ( .A(in[1272]), .B(in[312]), .Z(n1270) );
  XNOR U2230 ( .A(n1271), .B(n1270), .Z(n1272) );
  XNOR U2231 ( .A(in[952]), .B(n1272), .Z(n1646) );
  XNOR U2232 ( .A(n1273), .B(n1646), .Z(n3268) );
  IV U2233 ( .A(n3268), .Z(n4144) );
  XOR U2234 ( .A(in[568]), .B(n4144), .Z(n1746) );
  XNOR U2235 ( .A(in[168]), .B(n1274), .Z(n5148) );
  XOR U2236 ( .A(in[1353]), .B(n4449), .Z(n5145) );
  NAND U2237 ( .A(n5148), .B(n5145), .Z(n1275) );
  XNOR U2238 ( .A(n1746), .B(n1275), .Z(out[1061]) );
  XOR U2239 ( .A(in[633]), .B(in[1593]), .Z(n1277) );
  XNOR U2240 ( .A(in[1273]), .B(in[313]), .Z(n1276) );
  XNOR U2241 ( .A(n1277), .B(n1276), .Z(n1278) );
  XNOR U2242 ( .A(in[953]), .B(n1278), .Z(n1650) );
  XNOR U2243 ( .A(n1279), .B(n1650), .Z(n3271) );
  IV U2244 ( .A(n3271), .Z(n4148) );
  XOR U2245 ( .A(in[569]), .B(n4148), .Z(n1751) );
  XOR U2246 ( .A(in[329]), .B(in[969]), .Z(n1281) );
  XNOR U2247 ( .A(in[9]), .B(in[649]), .Z(n1280) );
  XNOR U2248 ( .A(n1281), .B(n1280), .Z(n1282) );
  XNOR U2249 ( .A(in[1289]), .B(n1282), .Z(n1423) );
  XOR U2250 ( .A(in[778]), .B(in[1098]), .Z(n1284) );
  XNOR U2251 ( .A(in[458]), .B(in[1418]), .Z(n1283) );
  XNOR U2252 ( .A(n1284), .B(n1283), .Z(n1285) );
  XNOR U2253 ( .A(in[138]), .B(n1285), .Z(n1372) );
  XOR U2254 ( .A(n1423), .B(n1372), .Z(n4452) );
  XNOR U2255 ( .A(in[1354]), .B(n4452), .Z(n5150) );
  XNOR U2256 ( .A(in[169]), .B(n1286), .Z(n5152) );
  NANDN U2257 ( .A(n5150), .B(n5152), .Z(n1287) );
  XNOR U2258 ( .A(n1751), .B(n1287), .Z(out[1062]) );
  XOR U2259 ( .A(in[634]), .B(in[1594]), .Z(n1289) );
  XNOR U2260 ( .A(in[1274]), .B(in[314]), .Z(n1288) );
  XNOR U2261 ( .A(n1289), .B(n1288), .Z(n1290) );
  XNOR U2262 ( .A(in[954]), .B(n1290), .Z(n1654) );
  XNOR U2263 ( .A(n1291), .B(n1654), .Z(n3274) );
  IV U2264 ( .A(n3274), .Z(n4152) );
  XOR U2265 ( .A(in[570]), .B(n4152), .Z(n1755) );
  XNOR U2266 ( .A(in[170]), .B(n1292), .Z(n5156) );
  XOR U2267 ( .A(in[1419]), .B(in[779]), .Z(n1294) );
  XNOR U2268 ( .A(in[1099]), .B(in[459]), .Z(n1293) );
  XNOR U2269 ( .A(n1294), .B(n1293), .Z(n1295) );
  XNOR U2270 ( .A(in[139]), .B(n1295), .Z(n1378) );
  XOR U2271 ( .A(in[1290]), .B(in[650]), .Z(n1297) );
  XNOR U2272 ( .A(in[970]), .B(in[330]), .Z(n1296) );
  XNOR U2273 ( .A(n1297), .B(n1296), .Z(n1298) );
  XNOR U2274 ( .A(in[10]), .B(n1298), .Z(n1425) );
  XOR U2275 ( .A(n1378), .B(n1425), .Z(n4455) );
  XOR U2276 ( .A(in[1355]), .B(n4455), .Z(n5153) );
  NAND U2277 ( .A(n5156), .B(n5153), .Z(n1299) );
  XNOR U2278 ( .A(n1755), .B(n1299), .Z(out[1063]) );
  XOR U2279 ( .A(in[955]), .B(in[1275]), .Z(n1301) );
  XNOR U2280 ( .A(in[1595]), .B(in[315]), .Z(n1300) );
  XNOR U2281 ( .A(n1301), .B(n1300), .Z(n1302) );
  XOR U2282 ( .A(in[635]), .B(n1302), .Z(n1658) );
  XOR U2283 ( .A(n1303), .B(n1658), .Z(n4162) );
  XOR U2284 ( .A(in[571]), .B(n4162), .Z(n1757) );
  XOR U2285 ( .A(in[956]), .B(in[1276]), .Z(n1305) );
  XNOR U2286 ( .A(in[1596]), .B(in[316]), .Z(n1304) );
  XNOR U2287 ( .A(n1305), .B(n1304), .Z(n1306) );
  XOR U2288 ( .A(in[636]), .B(n1306), .Z(n1662) );
  XOR U2289 ( .A(n1307), .B(n1662), .Z(n4166) );
  XOR U2290 ( .A(in[572]), .B(n4166), .Z(n1759) );
  XOR U2291 ( .A(in[957]), .B(in[1277]), .Z(n1309) );
  XNOR U2292 ( .A(in[1597]), .B(in[317]), .Z(n1308) );
  XNOR U2293 ( .A(n1309), .B(n1308), .Z(n1310) );
  XOR U2294 ( .A(in[637]), .B(n1310), .Z(n1667) );
  XOR U2295 ( .A(n1311), .B(n1667), .Z(n4170) );
  XOR U2296 ( .A(in[573]), .B(n4170), .Z(n1761) );
  IV U2297 ( .A(n3286), .Z(n4174) );
  XOR U2298 ( .A(in[574]), .B(n4174), .Z(n1763) );
  XOR U2299 ( .A(in[959]), .B(in[1279]), .Z(n1313) );
  XNOR U2300 ( .A(in[1599]), .B(in[319]), .Z(n1312) );
  XNOR U2301 ( .A(n1313), .B(n1312), .Z(n1314) );
  XOR U2302 ( .A(in[639]), .B(n1314), .Z(n1675) );
  XOR U2303 ( .A(n1315), .B(n1675), .Z(n3289) );
  XOR U2304 ( .A(in[575]), .B(n3289), .Z(n1764) );
  XOR U2305 ( .A(in[896]), .B(in[1216]), .Z(n1317) );
  XNOR U2306 ( .A(in[1536]), .B(in[256]), .Z(n1316) );
  XNOR U2307 ( .A(n1317), .B(n1316), .Z(n1318) );
  XOR U2308 ( .A(in[576]), .B(n1318), .Z(n1679) );
  XOR U2309 ( .A(n1319), .B(n1679), .Z(n3292) );
  XOR U2310 ( .A(in[512]), .B(n3292), .Z(n1766) );
  XOR U2311 ( .A(n1321), .B(n1320), .Z(n3975) );
  XOR U2312 ( .A(in[577]), .B(n3975), .Z(n2715) );
  IV U2313 ( .A(n2715), .Z(n2803) );
  XNOR U2314 ( .A(in[1452]), .B(n4115), .Z(n3243) );
  XNOR U2315 ( .A(in[232]), .B(n2042), .Z(n3245) );
  NANDN U2316 ( .A(n3243), .B(n3245), .Z(n1322) );
  XOR U2317 ( .A(n2803), .B(n1322), .Z(out[106]) );
  XOR U2318 ( .A(in[897]), .B(in[1217]), .Z(n1324) );
  XNOR U2319 ( .A(in[1537]), .B(in[257]), .Z(n1323) );
  XNOR U2320 ( .A(n1324), .B(n1323), .Z(n1325) );
  XOR U2321 ( .A(in[577]), .B(n1325), .Z(n1683) );
  XOR U2322 ( .A(n1326), .B(n1683), .Z(n3295) );
  XOR U2323 ( .A(in[513]), .B(n3295), .Z(n1768) );
  XOR U2324 ( .A(in[1538]), .B(in[578]), .Z(n1328) );
  XNOR U2325 ( .A(in[898]), .B(in[258]), .Z(n1327) );
  XNOR U2326 ( .A(n1328), .B(n1327), .Z(n1329) );
  XOR U2327 ( .A(in[1218]), .B(n1329), .Z(n1687) );
  XOR U2328 ( .A(n1330), .B(n1687), .Z(n3302) );
  XOR U2329 ( .A(in[514]), .B(n3302), .Z(n1770) );
  XOR U2330 ( .A(in[1539]), .B(in[579]), .Z(n1332) );
  XNOR U2331 ( .A(in[899]), .B(in[259]), .Z(n1331) );
  XNOR U2332 ( .A(n1332), .B(n1331), .Z(n1333) );
  XOR U2333 ( .A(in[1219]), .B(n1333), .Z(n1691) );
  XOR U2334 ( .A(n1334), .B(n1691), .Z(n3305) );
  XOR U2335 ( .A(in[515]), .B(n3305), .Z(n1774) );
  XOR U2336 ( .A(in[1540]), .B(in[580]), .Z(n1336) );
  XNOR U2337 ( .A(in[900]), .B(in[260]), .Z(n1335) );
  XNOR U2338 ( .A(n1336), .B(n1335), .Z(n1337) );
  XOR U2339 ( .A(in[1220]), .B(n1337), .Z(n1695) );
  XOR U2340 ( .A(n1338), .B(n1695), .Z(n3308) );
  XOR U2341 ( .A(in[516]), .B(n3308), .Z(n1776) );
  XOR U2342 ( .A(in[1541]), .B(in[581]), .Z(n1340) );
  XNOR U2343 ( .A(in[901]), .B(in[261]), .Z(n1339) );
  XNOR U2344 ( .A(n1340), .B(n1339), .Z(n1341) );
  XOR U2345 ( .A(in[1221]), .B(n1341), .Z(n1699) );
  XOR U2346 ( .A(n1342), .B(n1699), .Z(n3311) );
  XOR U2347 ( .A(in[517]), .B(n3311), .Z(n1778) );
  XOR U2348 ( .A(in[1542]), .B(in[582]), .Z(n1344) );
  XNOR U2349 ( .A(in[902]), .B(in[262]), .Z(n1343) );
  XNOR U2350 ( .A(n1344), .B(n1343), .Z(n1345) );
  XOR U2351 ( .A(in[1222]), .B(n1345), .Z(n1703) );
  XOR U2352 ( .A(n1346), .B(n1703), .Z(n3314) );
  XOR U2353 ( .A(in[518]), .B(n3314), .Z(n1780) );
  XOR U2354 ( .A(in[1543]), .B(in[583]), .Z(n1348) );
  XNOR U2355 ( .A(in[903]), .B(in[263]), .Z(n1347) );
  XNOR U2356 ( .A(n1348), .B(n1347), .Z(n1349) );
  XOR U2357 ( .A(in[1223]), .B(n1349), .Z(n1708) );
  IV U2358 ( .A(n3929), .Z(n3317) );
  XOR U2359 ( .A(in[519]), .B(n3317), .Z(n1782) );
  XOR U2360 ( .A(in[1544]), .B(in[584]), .Z(n1352) );
  XNOR U2361 ( .A(in[904]), .B(in[264]), .Z(n1351) );
  XNOR U2362 ( .A(n1352), .B(n1351), .Z(n1353) );
  XOR U2363 ( .A(in[1224]), .B(n1353), .Z(n1712) );
  XOR U2364 ( .A(n1354), .B(n1712), .Z(n3933) );
  XOR U2365 ( .A(in[520]), .B(n3933), .Z(n1784) );
  XOR U2366 ( .A(in[1545]), .B(in[585]), .Z(n1356) );
  XNOR U2367 ( .A(in[905]), .B(in[265]), .Z(n1355) );
  XNOR U2368 ( .A(n1356), .B(n1355), .Z(n1357) );
  XOR U2369 ( .A(in[1225]), .B(n1357), .Z(n1716) );
  XOR U2370 ( .A(n1358), .B(n1716), .Z(n3940) );
  XOR U2371 ( .A(in[521]), .B(n3940), .Z(n1786) );
  XOR U2372 ( .A(in[1546]), .B(in[586]), .Z(n1360) );
  XNOR U2373 ( .A(in[906]), .B(in[266]), .Z(n1359) );
  XNOR U2374 ( .A(n1360), .B(n1359), .Z(n1361) );
  XOR U2375 ( .A(in[1226]), .B(n1361), .Z(n1720) );
  XOR U2376 ( .A(n1362), .B(n1720), .Z(n3944) );
  XOR U2377 ( .A(in[522]), .B(n3944), .Z(n1788) );
  NOR U2378 ( .A(n1363), .B(n1561), .Z(n1364) );
  XNOR U2379 ( .A(n1788), .B(n1364), .Z(out[1079]) );
  XOR U2380 ( .A(n1366), .B(n1365), .Z(n3982) );
  XOR U2381 ( .A(in[578]), .B(n3982), .Z(n2717) );
  IV U2382 ( .A(n2717), .Z(n2805) );
  IV U2383 ( .A(n1367), .Z(n4119) );
  XOR U2384 ( .A(in[1453]), .B(n4119), .Z(n3255) );
  XNOR U2385 ( .A(in[233]), .B(n2044), .Z(n3257) );
  NANDN U2386 ( .A(n3255), .B(n3257), .Z(n1368) );
  XOR U2387 ( .A(n2805), .B(n1368), .Z(out[107]) );
  XOR U2388 ( .A(in[1547]), .B(in[587]), .Z(n1370) );
  XNOR U2389 ( .A(in[907]), .B(in[267]), .Z(n1369) );
  XNOR U2390 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U2391 ( .A(in[1227]), .B(n1371), .Z(n1724) );
  XOR U2392 ( .A(n1372), .B(n1724), .Z(n3948) );
  XOR U2393 ( .A(in[523]), .B(n3948), .Z(n1790) );
  NOR U2394 ( .A(n1373), .B(n1565), .Z(n1374) );
  XNOR U2395 ( .A(n1790), .B(n1374), .Z(out[1080]) );
  XOR U2396 ( .A(in[1548]), .B(in[588]), .Z(n1376) );
  XNOR U2397 ( .A(in[908]), .B(in[268]), .Z(n1375) );
  XNOR U2398 ( .A(n1376), .B(n1375), .Z(n1377) );
  XOR U2399 ( .A(in[1228]), .B(n1377), .Z(n1728) );
  XOR U2400 ( .A(n1378), .B(n1728), .Z(n3952) );
  XOR U2401 ( .A(in[524]), .B(n3952), .Z(n1792) );
  NOR U2402 ( .A(n1379), .B(n1569), .Z(n1380) );
  XNOR U2403 ( .A(n1792), .B(n1380), .Z(out[1081]) );
  XOR U2404 ( .A(in[1549]), .B(in[589]), .Z(n1382) );
  XNOR U2405 ( .A(in[909]), .B(in[269]), .Z(n1381) );
  XNOR U2406 ( .A(n1382), .B(n1381), .Z(n1383) );
  XNOR U2407 ( .A(in[1229]), .B(n1383), .Z(n1732) );
  XOR U2408 ( .A(n1732), .B(n1384), .Z(n3956) );
  XOR U2409 ( .A(in[525]), .B(n3956), .Z(n1796) );
  XOR U2410 ( .A(in[1550]), .B(in[590]), .Z(n1386) );
  XNOR U2411 ( .A(in[910]), .B(in[270]), .Z(n1385) );
  XNOR U2412 ( .A(n1386), .B(n1385), .Z(n1387) );
  XNOR U2413 ( .A(in[1230]), .B(n1387), .Z(n1736) );
  XOR U2414 ( .A(n1736), .B(n1388), .Z(n3960) );
  XOR U2415 ( .A(in[526]), .B(n3960), .Z(n1798) );
  XOR U2416 ( .A(in[1551]), .B(in[591]), .Z(n1390) );
  XNOR U2417 ( .A(in[911]), .B(in[271]), .Z(n1389) );
  XNOR U2418 ( .A(n1390), .B(n1389), .Z(n1391) );
  XNOR U2419 ( .A(in[1231]), .B(n1391), .Z(n1740) );
  XOR U2420 ( .A(n1740), .B(n1392), .Z(n3964) );
  XOR U2421 ( .A(in[527]), .B(n3964), .Z(n1800) );
  XOR U2422 ( .A(in[1552]), .B(in[592]), .Z(n1394) );
  XNOR U2423 ( .A(in[912]), .B(in[272]), .Z(n1393) );
  XNOR U2424 ( .A(n1394), .B(n1393), .Z(n1395) );
  XNOR U2425 ( .A(in[1232]), .B(n1395), .Z(n1744) );
  XOR U2426 ( .A(n1744), .B(n1396), .Z(n3968) );
  XOR U2427 ( .A(in[528]), .B(n3968), .Z(n1802) );
  XOR U2428 ( .A(in[1553]), .B(in[593]), .Z(n1398) );
  XNOR U2429 ( .A(in[913]), .B(in[273]), .Z(n1397) );
  XNOR U2430 ( .A(n1398), .B(n1397), .Z(n1399) );
  XOR U2431 ( .A(in[1233]), .B(n1399), .Z(n1749) );
  XOR U2432 ( .A(n1400), .B(n1749), .Z(n3972) );
  XOR U2433 ( .A(in[529]), .B(n3972), .Z(n1804) );
  XOR U2434 ( .A(in[1554]), .B(in[594]), .Z(n1402) );
  XNOR U2435 ( .A(in[914]), .B(in[274]), .Z(n1401) );
  XNOR U2436 ( .A(n1402), .B(n1401), .Z(n1403) );
  XOR U2437 ( .A(in[1234]), .B(n1403), .Z(n1753) );
  XOR U2438 ( .A(n1404), .B(n1753), .Z(n3976) );
  XOR U2439 ( .A(in[530]), .B(n3976), .Z(n1806) );
  XNOR U2440 ( .A(in[957]), .B(n3959), .Z(n1809) );
  XNOR U2441 ( .A(in[958]), .B(n3963), .Z(n1812) );
  XNOR U2442 ( .A(n1406), .B(n1405), .Z(n3986) );
  XOR U2443 ( .A(in[579]), .B(n3986), .Z(n2719) );
  IV U2444 ( .A(n2719), .Z(n2807) );
  IV U2445 ( .A(n1407), .Z(n4123) );
  XOR U2446 ( .A(in[1454]), .B(n4123), .Z(n3265) );
  XNOR U2447 ( .A(in[234]), .B(n2046), .Z(n3267) );
  NANDN U2448 ( .A(n3265), .B(n3267), .Z(n1408) );
  XOR U2449 ( .A(n2807), .B(n1408), .Z(out[108]) );
  XNOR U2450 ( .A(in[959]), .B(n3967), .Z(n1815) );
  XNOR U2451 ( .A(in[896]), .B(n3971), .Z(n1818) );
  XNOR U2452 ( .A(in[897]), .B(n3975), .Z(n1823) );
  XNOR U2453 ( .A(in[898]), .B(n3982), .Z(n1826) );
  XNOR U2454 ( .A(in[899]), .B(n3986), .Z(n1828) );
  XOR U2455 ( .A(n1410), .B(n1409), .Z(n2009) );
  XOR U2456 ( .A(in[900]), .B(n2009), .Z(n1829) );
  XOR U2457 ( .A(n1412), .B(n1411), .Z(n2011) );
  XOR U2458 ( .A(in[901]), .B(n2011), .Z(n1831) );
  XOR U2459 ( .A(n1414), .B(n1413), .Z(n2014) );
  XOR U2460 ( .A(in[902]), .B(n2014), .Z(n1833) );
  XOR U2461 ( .A(n1416), .B(n1415), .Z(n2017) );
  XOR U2462 ( .A(in[903]), .B(n2017), .Z(n1835) );
  XOR U2463 ( .A(n1418), .B(n1417), .Z(n2019) );
  XOR U2464 ( .A(in[904]), .B(n2019), .Z(n1837) );
  IV U2465 ( .A(n2009), .Z(n3990) );
  XOR U2466 ( .A(in[580]), .B(n3990), .Z(n2809) );
  IV U2467 ( .A(n1419), .Z(n4127) );
  XOR U2468 ( .A(in[1455]), .B(n4127), .Z(n3299) );
  XNOR U2469 ( .A(in[235]), .B(n4088), .Z(n3301) );
  NANDN U2470 ( .A(n3299), .B(n3301), .Z(n1420) );
  XNOR U2471 ( .A(n2809), .B(n1420), .Z(out[109]) );
  XNOR U2472 ( .A(in[200]), .B(n3933), .Z(n4280) );
  XOR U2473 ( .A(in[1420]), .B(n3192), .Z(n4281) );
  XNOR U2474 ( .A(n4483), .B(in[1043]), .Z(n2877) );
  NANDN U2475 ( .A(n4281), .B(n2877), .Z(n1421) );
  XNOR U2476 ( .A(n4280), .B(n1421), .Z(out[10]) );
  XOR U2477 ( .A(n1423), .B(n1422), .Z(n2021) );
  XOR U2478 ( .A(in[905]), .B(n2021), .Z(n1839) );
  XOR U2479 ( .A(n1425), .B(n1424), .Z(n2024) );
  XOR U2480 ( .A(in[906]), .B(n2024), .Z(n1841) );
  XOR U2481 ( .A(n1427), .B(n1426), .Z(n2026) );
  XOR U2482 ( .A(in[907]), .B(n2026), .Z(n1845) );
  XOR U2483 ( .A(n1429), .B(n1428), .Z(n2028) );
  XOR U2484 ( .A(in[908]), .B(n2028), .Z(n1847) );
  XOR U2485 ( .A(n1431), .B(n1430), .Z(n3108) );
  XOR U2486 ( .A(in[909]), .B(n3108), .Z(n1849) );
  XOR U2487 ( .A(n1433), .B(n1432), .Z(n3114) );
  XOR U2488 ( .A(in[910]), .B(n3114), .Z(n1851) );
  XNOR U2489 ( .A(n1435), .B(n1434), .Z(n3116) );
  XOR U2490 ( .A(in[911]), .B(n3116), .Z(n1853) );
  XNOR U2491 ( .A(n1437), .B(n1436), .Z(n3118) );
  XOR U2492 ( .A(in[912]), .B(n3118), .Z(n1855) );
  XOR U2493 ( .A(n1438), .B(n230), .Z(n4046) );
  XOR U2494 ( .A(in[913]), .B(n4046), .Z(n1857) );
  XOR U2495 ( .A(n1440), .B(n1439), .Z(n2036) );
  XOR U2496 ( .A(in[914]), .B(n2036), .Z(n1859) );
  IV U2497 ( .A(n2011), .Z(n3994) );
  XOR U2498 ( .A(in[581]), .B(n3994), .Z(n2811) );
  IV U2499 ( .A(n1441), .Z(n4131) );
  XOR U2500 ( .A(in[1456]), .B(n4131), .Z(n3329) );
  XNOR U2501 ( .A(in[236]), .B(n4092), .Z(n3331) );
  NANDN U2502 ( .A(n3329), .B(n3331), .Z(n1442) );
  XNOR U2503 ( .A(n2811), .B(n1442), .Z(out[110]) );
  XNOR U2504 ( .A(n1444), .B(n1443), .Z(n3122) );
  XOR U2505 ( .A(in[915]), .B(n3122), .Z(n1861) );
  XNOR U2506 ( .A(n1446), .B(n1445), .Z(n3124) );
  XOR U2507 ( .A(in[916]), .B(n3124), .Z(n1863) );
  XOR U2508 ( .A(n1448), .B(n1447), .Z(n3126) );
  XOR U2509 ( .A(in[917]), .B(n3126), .Z(n1867) );
  XOR U2510 ( .A(n1450), .B(n1449), .Z(n3128) );
  XOR U2511 ( .A(in[918]), .B(n3128), .Z(n1869) );
  XOR U2512 ( .A(n1452), .B(n1451), .Z(n3130) );
  XOR U2513 ( .A(in[919]), .B(n3130), .Z(n1871) );
  XNOR U2514 ( .A(n1454), .B(n1453), .Z(n3136) );
  XOR U2515 ( .A(in[920]), .B(n3136), .Z(n1873) );
  NOR U2516 ( .A(n1455), .B(n1705), .Z(n1456) );
  XNOR U2517 ( .A(n1873), .B(n1456), .Z(out[1115]) );
  XNOR U2518 ( .A(n1458), .B(n1457), .Z(n3138) );
  XOR U2519 ( .A(in[921]), .B(n3138), .Z(n1875) );
  XNOR U2520 ( .A(n1460), .B(n1459), .Z(n3141) );
  XOR U2521 ( .A(in[922]), .B(n3141), .Z(n1877) );
  XNOR U2522 ( .A(n1462), .B(n1461), .Z(n3143) );
  XOR U2523 ( .A(in[923]), .B(n3143), .Z(n1879) );
  NOR U2524 ( .A(n1463), .B(n1718), .Z(n1464) );
  XNOR U2525 ( .A(n1879), .B(n1464), .Z(out[1118]) );
  XNOR U2526 ( .A(n1466), .B(n1465), .Z(n3022) );
  XOR U2527 ( .A(in[924]), .B(n3022), .Z(n1881) );
  NOR U2528 ( .A(n1467), .B(n1722), .Z(n1468) );
  XNOR U2529 ( .A(n1881), .B(n1468), .Z(out[1119]) );
  IV U2530 ( .A(n2014), .Z(n3998) );
  XOR U2531 ( .A(in[582]), .B(n3998), .Z(n2813) );
  IV U2532 ( .A(n1469), .Z(n4135) );
  XOR U2533 ( .A(in[1457]), .B(n4135), .Z(n3358) );
  XNOR U2534 ( .A(in[237]), .B(n4096), .Z(n3360) );
  NANDN U2535 ( .A(n3358), .B(n3360), .Z(n1470) );
  XNOR U2536 ( .A(n2813), .B(n1470), .Z(out[111]) );
  XNOR U2537 ( .A(n1472), .B(n1471), .Z(n3024) );
  XOR U2538 ( .A(in[925]), .B(n3024), .Z(n1883) );
  NOR U2539 ( .A(n1473), .B(n1726), .Z(n1474) );
  XNOR U2540 ( .A(n1883), .B(n1474), .Z(out[1120]) );
  XNOR U2541 ( .A(n1476), .B(n1475), .Z(n3026) );
  XOR U2542 ( .A(in[926]), .B(n3026), .Z(n1885) );
  NOR U2543 ( .A(n1477), .B(n1730), .Z(n1478) );
  XNOR U2544 ( .A(n1885), .B(n1478), .Z(out[1121]) );
  XNOR U2545 ( .A(n1480), .B(n1479), .Z(n3028) );
  XOR U2546 ( .A(in[927]), .B(n3028), .Z(n1889) );
  XNOR U2547 ( .A(n1482), .B(n1481), .Z(n3030) );
  XOR U2548 ( .A(in[928]), .B(n3030), .Z(n1891) );
  NOR U2549 ( .A(n5140), .B(n1738), .Z(n1483) );
  XNOR U2550 ( .A(n1891), .B(n1483), .Z(out[1123]) );
  XOR U2551 ( .A(n1485), .B(n1484), .Z(n3032) );
  XOR U2552 ( .A(in[929]), .B(n3032), .Z(n1893) );
  NOR U2553 ( .A(n5144), .B(n1742), .Z(n1486) );
  XNOR U2554 ( .A(n1893), .B(n1486), .Z(out[1124]) );
  XOR U2555 ( .A(n1487), .B(n231), .Z(n4122) );
  XOR U2556 ( .A(in[930]), .B(n4122), .Z(n1895) );
  NOR U2557 ( .A(n5148), .B(n1746), .Z(n1488) );
  XNOR U2558 ( .A(n1895), .B(n1488), .Z(out[1125]) );
  XOR U2559 ( .A(n1490), .B(n1489), .Z(n3035) );
  XOR U2560 ( .A(in[931]), .B(n3035), .Z(n1897) );
  NOR U2561 ( .A(n5152), .B(n1751), .Z(n1491) );
  XNOR U2562 ( .A(n1897), .B(n1491), .Z(out[1126]) );
  XOR U2563 ( .A(n1493), .B(n1492), .Z(n3037) );
  XOR U2564 ( .A(in[932]), .B(n3037), .Z(n1899) );
  NOR U2565 ( .A(n5156), .B(n1755), .Z(n1494) );
  XNOR U2566 ( .A(n1899), .B(n1494), .Z(out[1127]) );
  XOR U2567 ( .A(n1496), .B(n1495), .Z(n4134) );
  XOR U2568 ( .A(in[933]), .B(n4134), .Z(n1902) );
  NAND U2569 ( .A(n1497), .B(n1757), .Z(n1498) );
  XNOR U2570 ( .A(n1902), .B(n1498), .Z(out[1128]) );
  XNOR U2571 ( .A(n1500), .B(n1499), .Z(n4138) );
  XOR U2572 ( .A(in[934]), .B(n4138), .Z(n1906) );
  NAND U2573 ( .A(n1501), .B(n1759), .Z(n1502) );
  XNOR U2574 ( .A(n1906), .B(n1502), .Z(out[1129]) );
  IV U2575 ( .A(n2017), .Z(n4002) );
  XOR U2576 ( .A(in[583]), .B(n4002), .Z(n2818) );
  IV U2577 ( .A(n1503), .Z(n4139) );
  XOR U2578 ( .A(in[1458]), .B(n4139), .Z(n3386) );
  XNOR U2579 ( .A(in[238]), .B(n4100), .Z(n3388) );
  NANDN U2580 ( .A(n3386), .B(n3388), .Z(n1504) );
  XNOR U2581 ( .A(n2818), .B(n1504), .Z(out[112]) );
  XOR U2582 ( .A(n1506), .B(n1505), .Z(n4142) );
  XOR U2583 ( .A(in[935]), .B(n4142), .Z(n1910) );
  NAND U2584 ( .A(n1507), .B(n1761), .Z(n1508) );
  XNOR U2585 ( .A(n1910), .B(n1508), .Z(out[1130]) );
  XOR U2586 ( .A(n1510), .B(n1509), .Z(n4146) );
  XOR U2587 ( .A(in[936]), .B(n4146), .Z(n1914) );
  NANDN U2588 ( .A(n1763), .B(n1511), .Z(n1512) );
  XNOR U2589 ( .A(n1914), .B(n1512), .Z(out[1131]) );
  XOR U2590 ( .A(n1514), .B(n1513), .Z(n4150) );
  XOR U2591 ( .A(in[937]), .B(n4150), .Z(n1920) );
  NAND U2592 ( .A(n1515), .B(n1764), .Z(n1516) );
  XNOR U2593 ( .A(n1920), .B(n1516), .Z(out[1132]) );
  XOR U2594 ( .A(n1518), .B(n1517), .Z(n4160) );
  XOR U2595 ( .A(in[938]), .B(n4160), .Z(n1924) );
  NAND U2596 ( .A(n1519), .B(n1766), .Z(n1520) );
  XNOR U2597 ( .A(n1924), .B(n1520), .Z(out[1133]) );
  XOR U2598 ( .A(n1522), .B(n1521), .Z(n4164) );
  XOR U2599 ( .A(in[939]), .B(n4164), .Z(n1928) );
  NAND U2600 ( .A(n1523), .B(n1768), .Z(n1524) );
  XNOR U2601 ( .A(n1928), .B(n1524), .Z(out[1134]) );
  XOR U2602 ( .A(n1526), .B(n1525), .Z(n4168) );
  XOR U2603 ( .A(in[940]), .B(n4168), .Z(n1932) );
  NAND U2604 ( .A(n1527), .B(n1770), .Z(n1528) );
  XNOR U2605 ( .A(n1932), .B(n1528), .Z(out[1135]) );
  XOR U2606 ( .A(n1530), .B(n1529), .Z(n4172) );
  XOR U2607 ( .A(in[941]), .B(n4172), .Z(n1936) );
  NAND U2608 ( .A(n1531), .B(n1774), .Z(n1532) );
  XNOR U2609 ( .A(n1936), .B(n1532), .Z(out[1136]) );
  XOR U2610 ( .A(n1534), .B(n1533), .Z(n3896) );
  XOR U2611 ( .A(in[942]), .B(n3896), .Z(n1940) );
  NAND U2612 ( .A(n1535), .B(n1776), .Z(n1536) );
  XNOR U2613 ( .A(n1940), .B(n1536), .Z(out[1137]) );
  XOR U2614 ( .A(n1538), .B(n1537), .Z(n3900) );
  XOR U2615 ( .A(in[943]), .B(n3900), .Z(n1944) );
  NAND U2616 ( .A(n1539), .B(n1778), .Z(n1540) );
  XNOR U2617 ( .A(n1944), .B(n1540), .Z(out[1138]) );
  XOR U2618 ( .A(n1542), .B(n1541), .Z(n3904) );
  XOR U2619 ( .A(in[944]), .B(n3904), .Z(n1948) );
  NAND U2620 ( .A(n1543), .B(n1780), .Z(n1544) );
  XNOR U2621 ( .A(n1948), .B(n1544), .Z(out[1139]) );
  IV U2622 ( .A(n2019), .Z(n4006) );
  XOR U2623 ( .A(in[584]), .B(n4006), .Z(n2820) );
  IV U2624 ( .A(n1545), .Z(n4143) );
  XOR U2625 ( .A(in[1459]), .B(n4143), .Z(n3421) );
  XNOR U2626 ( .A(in[239]), .B(n4104), .Z(n3423) );
  NANDN U2627 ( .A(n3421), .B(n3423), .Z(n1546) );
  XNOR U2628 ( .A(n2820), .B(n1546), .Z(out[113]) );
  XOR U2629 ( .A(n1548), .B(n1547), .Z(n3908) );
  XOR U2630 ( .A(in[945]), .B(n3908), .Z(n1952) );
  NAND U2631 ( .A(n1549), .B(n1782), .Z(n1550) );
  XNOR U2632 ( .A(n1952), .B(n1550), .Z(out[1140]) );
  XOR U2633 ( .A(n1552), .B(n1551), .Z(n3912) );
  XOR U2634 ( .A(in[946]), .B(n3912), .Z(n1956) );
  NAND U2635 ( .A(n1553), .B(n1784), .Z(n1554) );
  XNOR U2636 ( .A(n1956), .B(n1554), .Z(out[1141]) );
  XNOR U2637 ( .A(n1556), .B(n1555), .Z(n3916) );
  IV U2638 ( .A(n3916), .Z(n2567) );
  XOR U2639 ( .A(in[947]), .B(n2567), .Z(n1962) );
  NAND U2640 ( .A(n1557), .B(n1786), .Z(n1558) );
  XNOR U2641 ( .A(n1962), .B(n1558), .Z(out[1142]) );
  XNOR U2642 ( .A(n1560), .B(n1559), .Z(n3920) );
  IV U2643 ( .A(n3920), .Z(n2609) );
  XOR U2644 ( .A(in[948]), .B(n2609), .Z(n1966) );
  NAND U2645 ( .A(n1561), .B(n1788), .Z(n1562) );
  XNOR U2646 ( .A(n1966), .B(n1562), .Z(out[1143]) );
  XNOR U2647 ( .A(n1564), .B(n1563), .Z(n3924) );
  IV U2648 ( .A(n3924), .Z(n2651) );
  XOR U2649 ( .A(in[949]), .B(n2651), .Z(n1970) );
  NAND U2650 ( .A(n1565), .B(n1790), .Z(n1566) );
  XNOR U2651 ( .A(n1970), .B(n1566), .Z(out[1144]) );
  XOR U2652 ( .A(n1568), .B(n1567), .Z(n3063) );
  XOR U2653 ( .A(in[950]), .B(n3063), .Z(n1974) );
  NAND U2654 ( .A(n1569), .B(n1792), .Z(n1570) );
  XNOR U2655 ( .A(n1974), .B(n1570), .Z(out[1145]) );
  XOR U2656 ( .A(n1572), .B(n1571), .Z(n3065) );
  XOR U2657 ( .A(in[951]), .B(n3065), .Z(n1978) );
  NAND U2658 ( .A(n1573), .B(n1796), .Z(n1574) );
  XNOR U2659 ( .A(n1978), .B(n1574), .Z(out[1146]) );
  XOR U2660 ( .A(n1576), .B(n1575), .Z(n3068) );
  XOR U2661 ( .A(in[952]), .B(n3068), .Z(n1982) );
  NAND U2662 ( .A(n1577), .B(n1798), .Z(n1578) );
  XNOR U2663 ( .A(n1982), .B(n1578), .Z(out[1147]) );
  XNOR U2664 ( .A(n1580), .B(n1579), .Z(n3943) );
  IV U2665 ( .A(n3943), .Z(n2698) );
  XOR U2666 ( .A(in[953]), .B(n2698), .Z(n1986) );
  NAND U2667 ( .A(n1581), .B(n1800), .Z(n1582) );
  XNOR U2668 ( .A(n1986), .B(n1582), .Z(out[1148]) );
  XNOR U2669 ( .A(n1584), .B(n1583), .Z(n3947) );
  IV U2670 ( .A(n3947), .Z(n2700) );
  XOR U2671 ( .A(in[954]), .B(n2700), .Z(n1990) );
  NAND U2672 ( .A(n1585), .B(n1802), .Z(n1586) );
  XNOR U2673 ( .A(n1990), .B(n1586), .Z(out[1149]) );
  IV U2674 ( .A(n2021), .Z(n4010) );
  XOR U2675 ( .A(in[585]), .B(n4010), .Z(n2822) );
  IV U2676 ( .A(n1587), .Z(n4147) );
  XOR U2677 ( .A(in[1460]), .B(n4147), .Z(n3456) );
  XNOR U2678 ( .A(in[240]), .B(n4108), .Z(n3458) );
  NANDN U2679 ( .A(n3456), .B(n3458), .Z(n1588) );
  XNOR U2680 ( .A(n2822), .B(n1588), .Z(out[114]) );
  XOR U2681 ( .A(in[955]), .B(n3951), .Z(n1994) );
  NAND U2682 ( .A(n1589), .B(n1804), .Z(n1590) );
  XNOR U2683 ( .A(n1994), .B(n1590), .Z(out[1150]) );
  XOR U2684 ( .A(in[956]), .B(n3955), .Z(n1998) );
  NANDN U2685 ( .A(n1591), .B(n1806), .Z(n1592) );
  XNOR U2686 ( .A(n1998), .B(n1592), .Z(out[1151]) );
  XOR U2687 ( .A(n1594), .B(n1593), .Z(n4296) );
  XOR U2688 ( .A(in[1004]), .B(n4296), .Z(n1808) );
  NAND U2689 ( .A(n1595), .B(n1809), .Z(n1596) );
  XNOR U2690 ( .A(n1808), .B(n1596), .Z(out[1152]) );
  XOR U2691 ( .A(n1598), .B(n1597), .Z(n4298) );
  XOR U2692 ( .A(in[1005]), .B(n4298), .Z(n1811) );
  NAND U2693 ( .A(n1599), .B(n1812), .Z(n1600) );
  XNOR U2694 ( .A(n1811), .B(n1600), .Z(out[1153]) );
  XOR U2695 ( .A(n1602), .B(n1601), .Z(n4300) );
  XOR U2696 ( .A(in[1006]), .B(n4300), .Z(n1814) );
  NAND U2697 ( .A(n1603), .B(n1815), .Z(n1604) );
  XNOR U2698 ( .A(n1814), .B(n1604), .Z(out[1154]) );
  XOR U2699 ( .A(n1606), .B(n1605), .Z(n4302) );
  XOR U2700 ( .A(in[1007]), .B(n4302), .Z(n1817) );
  NAND U2701 ( .A(n1607), .B(n1818), .Z(n1608) );
  XNOR U2702 ( .A(n1817), .B(n1608), .Z(out[1155]) );
  XOR U2703 ( .A(n1610), .B(n1609), .Z(n4309) );
  XOR U2704 ( .A(in[1008]), .B(n4309), .Z(n1822) );
  NAND U2705 ( .A(n1611), .B(n1823), .Z(n1612) );
  XNOR U2706 ( .A(n1822), .B(n1612), .Z(out[1156]) );
  XOR U2707 ( .A(n1614), .B(n1613), .Z(n4312) );
  XOR U2708 ( .A(in[1009]), .B(n4312), .Z(n1825) );
  NAND U2709 ( .A(n1615), .B(n1826), .Z(n1616) );
  XNOR U2710 ( .A(n1825), .B(n1616), .Z(out[1157]) );
  XOR U2711 ( .A(n1618), .B(n1617), .Z(n4315) );
  XOR U2712 ( .A(in[1010]), .B(n4315), .Z(n5023) );
  NAND U2713 ( .A(n1619), .B(n1828), .Z(n1620) );
  XNOR U2714 ( .A(n5023), .B(n1620), .Z(out[1158]) );
  XOR U2715 ( .A(n1622), .B(n1621), .Z(n4318) );
  XOR U2716 ( .A(in[1011]), .B(n4318), .Z(n5027) );
  NAND U2717 ( .A(n1623), .B(n1829), .Z(n1624) );
  XNOR U2718 ( .A(n5027), .B(n1624), .Z(out[1159]) );
  IV U2719 ( .A(n2024), .Z(n4014) );
  XOR U2720 ( .A(in[586]), .B(n4014), .Z(n2824) );
  XNOR U2721 ( .A(in[1461]), .B(n4151), .Z(n3478) );
  XNOR U2722 ( .A(in[241]), .B(n4116), .Z(n3480) );
  NANDN U2723 ( .A(n3478), .B(n3480), .Z(n1625) );
  XNOR U2724 ( .A(n2824), .B(n1625), .Z(out[115]) );
  XOR U2725 ( .A(n1627), .B(n1626), .Z(n4321) );
  XOR U2726 ( .A(in[1012]), .B(n4321), .Z(n5031) );
  NAND U2727 ( .A(n1628), .B(n1831), .Z(n1629) );
  XNOR U2728 ( .A(n5031), .B(n1629), .Z(out[1160]) );
  XOR U2729 ( .A(n1631), .B(n1630), .Z(n4324) );
  XOR U2730 ( .A(in[1013]), .B(n4324), .Z(n5035) );
  NAND U2731 ( .A(n1632), .B(n1833), .Z(n1633) );
  XNOR U2732 ( .A(n5035), .B(n1633), .Z(out[1161]) );
  XOR U2733 ( .A(n1635), .B(n1634), .Z(n4327) );
  XOR U2734 ( .A(in[1014]), .B(n4327), .Z(n5043) );
  NAND U2735 ( .A(n1636), .B(n1835), .Z(n1637) );
  XNOR U2736 ( .A(n5043), .B(n1637), .Z(out[1162]) );
  XOR U2737 ( .A(n1639), .B(n1638), .Z(n4330) );
  XOR U2738 ( .A(in[1015]), .B(n4330), .Z(n5047) );
  NAND U2739 ( .A(n1640), .B(n1837), .Z(n1641) );
  XNOR U2740 ( .A(n5047), .B(n1641), .Z(out[1163]) );
  XOR U2741 ( .A(n1643), .B(n1642), .Z(n4176) );
  XOR U2742 ( .A(in[1016]), .B(n4176), .Z(n5051) );
  NAND U2743 ( .A(n1644), .B(n1839), .Z(n1645) );
  XNOR U2744 ( .A(n5051), .B(n1645), .Z(out[1164]) );
  XOR U2745 ( .A(n1647), .B(n1646), .Z(n4179) );
  XOR U2746 ( .A(in[1017]), .B(n4179), .Z(n5055) );
  NAND U2747 ( .A(n1648), .B(n1841), .Z(n1649) );
  XNOR U2748 ( .A(n5055), .B(n1649), .Z(out[1165]) );
  XOR U2749 ( .A(n1651), .B(n1650), .Z(n4182) );
  XOR U2750 ( .A(in[1018]), .B(n4182), .Z(n5059) );
  NAND U2751 ( .A(n1652), .B(n1845), .Z(n1653) );
  XNOR U2752 ( .A(n5059), .B(n1653), .Z(out[1166]) );
  XOR U2753 ( .A(n1655), .B(n1654), .Z(n4185) );
  XOR U2754 ( .A(in[1019]), .B(n4185), .Z(n5063) );
  NANDN U2755 ( .A(n1656), .B(n1847), .Z(n1657) );
  XNOR U2756 ( .A(n5063), .B(n1657), .Z(out[1167]) );
  IV U2757 ( .A(n3057), .Z(n4188) );
  XOR U2758 ( .A(in[1020]), .B(n4188), .Z(n5066) );
  NANDN U2759 ( .A(n1660), .B(n1849), .Z(n1661) );
  XOR U2760 ( .A(n5066), .B(n1661), .Z(out[1168]) );
  IV U2761 ( .A(n3059), .Z(n4191) );
  XOR U2762 ( .A(in[1021]), .B(n4191), .Z(n5069) );
  NANDN U2763 ( .A(n1664), .B(n1851), .Z(n1665) );
  XOR U2764 ( .A(n5069), .B(n1665), .Z(out[1169]) );
  IV U2765 ( .A(n2026), .Z(n4018) );
  XOR U2766 ( .A(in[587]), .B(n4018), .Z(n2826) );
  XNOR U2767 ( .A(in[1462]), .B(n4161), .Z(n3500) );
  XNOR U2768 ( .A(in[242]), .B(n4120), .Z(n3502) );
  NANDN U2769 ( .A(n3500), .B(n3502), .Z(n1666) );
  XNOR U2770 ( .A(n2826), .B(n1666), .Z(out[116]) );
  IV U2771 ( .A(n3061), .Z(n4196) );
  XOR U2772 ( .A(in[1022]), .B(n4196), .Z(n5072) );
  NANDN U2773 ( .A(n1669), .B(n1853), .Z(n1670) );
  XOR U2774 ( .A(n5072), .B(n1670), .Z(out[1170]) );
  XOR U2775 ( .A(n1672), .B(n1671), .Z(n4197) );
  XOR U2776 ( .A(in[1023]), .B(n4197), .Z(n5076) );
  NAND U2777 ( .A(n1673), .B(n1855), .Z(n1674) );
  XNOR U2778 ( .A(n5076), .B(n1674), .Z(out[1171]) );
  IV U2779 ( .A(n3066), .Z(n4198) );
  XOR U2780 ( .A(in[960]), .B(n4198), .Z(n5083) );
  NAND U2781 ( .A(n1677), .B(n1857), .Z(n1678) );
  XOR U2782 ( .A(n5083), .B(n1678), .Z(out[1172]) );
  IV U2783 ( .A(n3069), .Z(n4199) );
  XOR U2784 ( .A(in[961]), .B(n4199), .Z(n5086) );
  NAND U2785 ( .A(n1681), .B(n1859), .Z(n1682) );
  XOR U2786 ( .A(n5086), .B(n1682), .Z(out[1173]) );
  IV U2787 ( .A(n3071), .Z(n4200) );
  XOR U2788 ( .A(in[962]), .B(n4200), .Z(n5089) );
  NAND U2789 ( .A(n1685), .B(n1861), .Z(n1686) );
  XOR U2790 ( .A(n5089), .B(n1686), .Z(out[1174]) );
  IV U2791 ( .A(n3075), .Z(n4201) );
  XOR U2792 ( .A(in[963]), .B(n4201), .Z(n5092) );
  NAND U2793 ( .A(n1689), .B(n1863), .Z(n1690) );
  XOR U2794 ( .A(n5092), .B(n1690), .Z(out[1175]) );
  IV U2795 ( .A(n3077), .Z(n4202) );
  XOR U2796 ( .A(in[964]), .B(n4202), .Z(n5095) );
  NAND U2797 ( .A(n1693), .B(n1867), .Z(n1694) );
  XOR U2798 ( .A(n5095), .B(n1694), .Z(out[1176]) );
  IV U2799 ( .A(n3079), .Z(n4203) );
  XOR U2800 ( .A(in[965]), .B(n4203), .Z(n5098) );
  NAND U2801 ( .A(n1697), .B(n1869), .Z(n1698) );
  XOR U2802 ( .A(n5098), .B(n1698), .Z(out[1177]) );
  IV U2803 ( .A(n3081), .Z(n4206) );
  XOR U2804 ( .A(in[966]), .B(n4206), .Z(n5101) );
  NAND U2805 ( .A(n1701), .B(n1871), .Z(n1702) );
  XOR U2806 ( .A(n5101), .B(n1702), .Z(out[1178]) );
  IV U2807 ( .A(n3083), .Z(n4209) );
  XOR U2808 ( .A(in[967]), .B(n4209), .Z(n5104) );
  NAND U2809 ( .A(n1705), .B(n1873), .Z(n1706) );
  XOR U2810 ( .A(n5104), .B(n1706), .Z(out[1179]) );
  IV U2811 ( .A(n2028), .Z(n4026) );
  XOR U2812 ( .A(in[588]), .B(n4026), .Z(n2828) );
  XNOR U2813 ( .A(in[1463]), .B(n4165), .Z(n3515) );
  XNOR U2814 ( .A(in[243]), .B(n4124), .Z(n3517) );
  NANDN U2815 ( .A(n3515), .B(n3517), .Z(n1707) );
  XNOR U2816 ( .A(n2828), .B(n1707), .Z(out[117]) );
  XNOR U2817 ( .A(n1709), .B(n1708), .Z(n4214) );
  XOR U2818 ( .A(in[968]), .B(n4214), .Z(n5108) );
  NAND U2819 ( .A(n1710), .B(n1875), .Z(n1711) );
  XNOR U2820 ( .A(n5108), .B(n1711), .Z(out[1180]) );
  IV U2821 ( .A(n3086), .Z(n4217) );
  XOR U2822 ( .A(in[969]), .B(n4217), .Z(n5111) );
  NAND U2823 ( .A(n1714), .B(n1877), .Z(n1715) );
  XOR U2824 ( .A(n5111), .B(n1715), .Z(out[1181]) );
  IV U2825 ( .A(n3088), .Z(n4220) );
  XOR U2826 ( .A(in[970]), .B(n4220), .Z(n5118) );
  NAND U2827 ( .A(n1718), .B(n1879), .Z(n1719) );
  XOR U2828 ( .A(n5118), .B(n1719), .Z(out[1182]) );
  XOR U2829 ( .A(in[971]), .B(n3090), .Z(n5122) );
  NAND U2830 ( .A(n1722), .B(n1881), .Z(n1723) );
  XNOR U2831 ( .A(n5122), .B(n1723), .Z(out[1183]) );
  XOR U2832 ( .A(in[972]), .B(n3092), .Z(n5126) );
  NAND U2833 ( .A(n1726), .B(n1883), .Z(n1727) );
  XNOR U2834 ( .A(n5126), .B(n1727), .Z(out[1184]) );
  XOR U2835 ( .A(in[973]), .B(n3096), .Z(n5130) );
  NAND U2836 ( .A(n1730), .B(n1885), .Z(n1731) );
  XNOR U2837 ( .A(n5130), .B(n1731), .Z(out[1185]) );
  XOR U2838 ( .A(n1733), .B(n1732), .Z(n4232) );
  XOR U2839 ( .A(in[974]), .B(n4232), .Z(n5134) );
  NAND U2840 ( .A(n1734), .B(n1889), .Z(n1735) );
  XNOR U2841 ( .A(n5134), .B(n1735), .Z(out[1186]) );
  XOR U2842 ( .A(n1737), .B(n1736), .Z(n4235) );
  XOR U2843 ( .A(in[975]), .B(n4235), .Z(n5138) );
  NAND U2844 ( .A(n1738), .B(n1891), .Z(n1739) );
  XNOR U2845 ( .A(n5138), .B(n1739), .Z(out[1187]) );
  XOR U2846 ( .A(n1741), .B(n1740), .Z(n4238) );
  XOR U2847 ( .A(in[976]), .B(n4238), .Z(n5142) );
  NAND U2848 ( .A(n1742), .B(n1893), .Z(n1743) );
  XNOR U2849 ( .A(n5142), .B(n1743), .Z(out[1188]) );
  XOR U2850 ( .A(n1745), .B(n1744), .Z(n4239) );
  XOR U2851 ( .A(in[977]), .B(n4239), .Z(n5146) );
  NAND U2852 ( .A(n1746), .B(n1895), .Z(n1747) );
  XNOR U2853 ( .A(n5146), .B(n1747), .Z(out[1189]) );
  IV U2854 ( .A(n3108), .Z(n4030) );
  XOR U2855 ( .A(in[589]), .B(n4030), .Z(n2830) );
  XNOR U2856 ( .A(in[1464]), .B(n4169), .Z(n3543) );
  XNOR U2857 ( .A(in[244]), .B(n4128), .Z(n3545) );
  NANDN U2858 ( .A(n3543), .B(n3545), .Z(n1748) );
  XNOR U2859 ( .A(n2830), .B(n1748), .Z(out[118]) );
  XOR U2860 ( .A(in[978]), .B(n3102), .Z(n5149) );
  NAND U2861 ( .A(n1751), .B(n1897), .Z(n1752) );
  XNOR U2862 ( .A(n5149), .B(n1752), .Z(out[1190]) );
  XOR U2863 ( .A(in[979]), .B(n3104), .Z(n5154) );
  NAND U2864 ( .A(n1755), .B(n1899), .Z(n1756) );
  XNOR U2865 ( .A(n5154), .B(n1756), .Z(out[1191]) );
  OR U2866 ( .A(n1902), .B(n1757), .Z(n1758) );
  XNOR U2867 ( .A(n1901), .B(n1758), .Z(out[1192]) );
  OR U2868 ( .A(n1906), .B(n1759), .Z(n1760) );
  XNOR U2869 ( .A(n1905), .B(n1760), .Z(out[1193]) );
  OR U2870 ( .A(n1910), .B(n1761), .Z(n1762) );
  XNOR U2871 ( .A(n1909), .B(n1762), .Z(out[1194]) );
  OR U2872 ( .A(n1920), .B(n1764), .Z(n1765) );
  XNOR U2873 ( .A(n1919), .B(n1765), .Z(out[1196]) );
  OR U2874 ( .A(n1924), .B(n1766), .Z(n1767) );
  XNOR U2875 ( .A(n1923), .B(n1767), .Z(out[1197]) );
  OR U2876 ( .A(n1928), .B(n1768), .Z(n1769) );
  XNOR U2877 ( .A(n1927), .B(n1769), .Z(out[1198]) );
  OR U2878 ( .A(n1932), .B(n1770), .Z(n1771) );
  XNOR U2879 ( .A(n1931), .B(n1771), .Z(out[1199]) );
  IV U2880 ( .A(n3114), .Z(n4034) );
  XOR U2881 ( .A(in[590]), .B(n4034), .Z(n2832) );
  XNOR U2882 ( .A(in[1465]), .B(n4173), .Z(n3573) );
  XNOR U2883 ( .A(in[245]), .B(n4132), .Z(n3575) );
  NANDN U2884 ( .A(n3573), .B(n3575), .Z(n1772) );
  XNOR U2885 ( .A(n2832), .B(n1772), .Z(out[119]) );
  XNOR U2886 ( .A(in[201]), .B(n3940), .Z(n4305) );
  XOR U2887 ( .A(in[1421]), .B(n3194), .Z(n4306) );
  XNOR U2888 ( .A(in[1044]), .B(n4486), .Z(n2881) );
  NANDN U2889 ( .A(n4306), .B(n2881), .Z(n1773) );
  XNOR U2890 ( .A(n4305), .B(n1773), .Z(out[11]) );
  OR U2891 ( .A(n1936), .B(n1774), .Z(n1775) );
  XNOR U2892 ( .A(n1935), .B(n1775), .Z(out[1200]) );
  OR U2893 ( .A(n1940), .B(n1776), .Z(n1777) );
  XNOR U2894 ( .A(n1939), .B(n1777), .Z(out[1201]) );
  OR U2895 ( .A(n1944), .B(n1778), .Z(n1779) );
  XNOR U2896 ( .A(n1943), .B(n1779), .Z(out[1202]) );
  OR U2897 ( .A(n1948), .B(n1780), .Z(n1781) );
  XNOR U2898 ( .A(n1947), .B(n1781), .Z(out[1203]) );
  OR U2899 ( .A(n1952), .B(n1782), .Z(n1783) );
  XNOR U2900 ( .A(n1951), .B(n1783), .Z(out[1204]) );
  OR U2901 ( .A(n1956), .B(n1784), .Z(n1785) );
  XNOR U2902 ( .A(n1955), .B(n1785), .Z(out[1205]) );
  OR U2903 ( .A(n1962), .B(n1786), .Z(n1787) );
  XNOR U2904 ( .A(n1961), .B(n1787), .Z(out[1206]) );
  OR U2905 ( .A(n1966), .B(n1788), .Z(n1789) );
  XNOR U2906 ( .A(n1965), .B(n1789), .Z(out[1207]) );
  OR U2907 ( .A(n1970), .B(n1790), .Z(n1791) );
  XNOR U2908 ( .A(n1969), .B(n1791), .Z(out[1208]) );
  OR U2909 ( .A(n1974), .B(n1792), .Z(n1793) );
  XNOR U2910 ( .A(n1973), .B(n1793), .Z(out[1209]) );
  IV U2911 ( .A(n3116), .Z(n4038) );
  XOR U2912 ( .A(in[591]), .B(n4038), .Z(n2834) );
  IV U2913 ( .A(n1794), .Z(n3897) );
  XOR U2914 ( .A(in[1466]), .B(n3897), .Z(n3597) );
  XNOR U2915 ( .A(in[246]), .B(n4136), .Z(n3599) );
  NANDN U2916 ( .A(n3597), .B(n3599), .Z(n1795) );
  XNOR U2917 ( .A(n2834), .B(n1795), .Z(out[120]) );
  OR U2918 ( .A(n1978), .B(n1796), .Z(n1797) );
  XNOR U2919 ( .A(n1977), .B(n1797), .Z(out[1210]) );
  OR U2920 ( .A(n1982), .B(n1798), .Z(n1799) );
  XNOR U2921 ( .A(n1981), .B(n1799), .Z(out[1211]) );
  OR U2922 ( .A(n1986), .B(n1800), .Z(n1801) );
  XNOR U2923 ( .A(n1985), .B(n1801), .Z(out[1212]) );
  OR U2924 ( .A(n1990), .B(n1802), .Z(n1803) );
  XNOR U2925 ( .A(n1989), .B(n1803), .Z(out[1213]) );
  OR U2926 ( .A(n1994), .B(n1804), .Z(n1805) );
  XNOR U2927 ( .A(n1993), .B(n1805), .Z(out[1214]) );
  OR U2928 ( .A(n1998), .B(n1806), .Z(n1807) );
  XNOR U2929 ( .A(n1997), .B(n1807), .Z(out[1215]) );
  IV U2930 ( .A(n1808), .Z(n4998) );
  NANDN U2931 ( .A(n1809), .B(n4998), .Z(n1810) );
  XOR U2932 ( .A(n4999), .B(n1810), .Z(out[1216]) );
  IV U2933 ( .A(n1811), .Z(n5002) );
  NANDN U2934 ( .A(n1812), .B(n5002), .Z(n1813) );
  XOR U2935 ( .A(n5003), .B(n1813), .Z(out[1217]) );
  IV U2936 ( .A(n1814), .Z(n5006) );
  NANDN U2937 ( .A(n1815), .B(n5006), .Z(n1816) );
  XOR U2938 ( .A(n5007), .B(n1816), .Z(out[1218]) );
  IV U2939 ( .A(n1817), .Z(n5010) );
  NANDN U2940 ( .A(n1818), .B(n5010), .Z(n1819) );
  XOR U2941 ( .A(n5011), .B(n1819), .Z(out[1219]) );
  IV U2942 ( .A(n3118), .Z(n4042) );
  XOR U2943 ( .A(in[592]), .B(n4042), .Z(n2836) );
  IV U2944 ( .A(n1820), .Z(n3901) );
  XOR U2945 ( .A(in[1467]), .B(n3901), .Z(n3627) );
  XNOR U2946 ( .A(in[247]), .B(n4140), .Z(n3629) );
  NANDN U2947 ( .A(n3627), .B(n3629), .Z(n1821) );
  XNOR U2948 ( .A(n2836), .B(n1821), .Z(out[121]) );
  IV U2949 ( .A(n1822), .Z(n5014) );
  NANDN U2950 ( .A(n1823), .B(n5014), .Z(n1824) );
  XOR U2951 ( .A(n5015), .B(n1824), .Z(out[1220]) );
  IV U2952 ( .A(n1825), .Z(n5018) );
  NANDN U2953 ( .A(n1826), .B(n5018), .Z(n1827) );
  XOR U2954 ( .A(n5019), .B(n1827), .Z(out[1221]) );
  OR U2955 ( .A(n5027), .B(n1829), .Z(n1830) );
  XNOR U2956 ( .A(n5026), .B(n1830), .Z(out[1223]) );
  OR U2957 ( .A(n5031), .B(n1831), .Z(n1832) );
  XNOR U2958 ( .A(n5030), .B(n1832), .Z(out[1224]) );
  OR U2959 ( .A(n5035), .B(n1833), .Z(n1834) );
  XNOR U2960 ( .A(n5034), .B(n1834), .Z(out[1225]) );
  OR U2961 ( .A(n5043), .B(n1835), .Z(n1836) );
  XNOR U2962 ( .A(n5042), .B(n1836), .Z(out[1226]) );
  OR U2963 ( .A(n5047), .B(n1837), .Z(n1838) );
  XNOR U2964 ( .A(n5046), .B(n1838), .Z(out[1227]) );
  OR U2965 ( .A(n5051), .B(n1839), .Z(n1840) );
  XNOR U2966 ( .A(n5050), .B(n1840), .Z(out[1228]) );
  OR U2967 ( .A(n5055), .B(n1841), .Z(n1842) );
  XNOR U2968 ( .A(n5054), .B(n1842), .Z(out[1229]) );
  XNOR U2969 ( .A(in[593]), .B(n4046), .Z(n2841) );
  IV U2970 ( .A(n1843), .Z(n3905) );
  XOR U2971 ( .A(in[1468]), .B(n3905), .Z(n3671) );
  XNOR U2972 ( .A(in[248]), .B(n4144), .Z(n3673) );
  NANDN U2973 ( .A(n3671), .B(n3673), .Z(n1844) );
  XNOR U2974 ( .A(n2841), .B(n1844), .Z(out[122]) );
  OR U2975 ( .A(n5059), .B(n1845), .Z(n1846) );
  XNOR U2976 ( .A(n5058), .B(n1846), .Z(out[1230]) );
  OR U2977 ( .A(n5063), .B(n1847), .Z(n1848) );
  XNOR U2978 ( .A(n5062), .B(n1848), .Z(out[1231]) );
  NANDN U2979 ( .A(n1849), .B(n5066), .Z(n1850) );
  XNOR U2980 ( .A(n5067), .B(n1850), .Z(out[1232]) );
  NANDN U2981 ( .A(n1851), .B(n5069), .Z(n1852) );
  XNOR U2982 ( .A(n5070), .B(n1852), .Z(out[1233]) );
  NANDN U2983 ( .A(n1853), .B(n5072), .Z(n1854) );
  XNOR U2984 ( .A(n5073), .B(n1854), .Z(out[1234]) );
  OR U2985 ( .A(n5076), .B(n1855), .Z(n1856) );
  XNOR U2986 ( .A(n5075), .B(n1856), .Z(out[1235]) );
  NANDN U2987 ( .A(n1857), .B(n5083), .Z(n1858) );
  XNOR U2988 ( .A(n5084), .B(n1858), .Z(out[1236]) );
  NANDN U2989 ( .A(n1859), .B(n5086), .Z(n1860) );
  XNOR U2990 ( .A(n5087), .B(n1860), .Z(out[1237]) );
  NANDN U2991 ( .A(n1861), .B(n5089), .Z(n1862) );
  XNOR U2992 ( .A(n5090), .B(n1862), .Z(out[1238]) );
  NANDN U2993 ( .A(n1863), .B(n5092), .Z(n1864) );
  XNOR U2994 ( .A(n5093), .B(n1864), .Z(out[1239]) );
  IV U2995 ( .A(n2036), .Z(n4050) );
  XOR U2996 ( .A(in[594]), .B(n4050), .Z(n2843) );
  IV U2997 ( .A(n1865), .Z(n3909) );
  XOR U2998 ( .A(in[1469]), .B(n3909), .Z(n3715) );
  XNOR U2999 ( .A(in[249]), .B(n4148), .Z(n3717) );
  NANDN U3000 ( .A(n3715), .B(n3717), .Z(n1866) );
  XNOR U3001 ( .A(n2843), .B(n1866), .Z(out[123]) );
  NANDN U3002 ( .A(n1867), .B(n5095), .Z(n1868) );
  XNOR U3003 ( .A(n5096), .B(n1868), .Z(out[1240]) );
  NANDN U3004 ( .A(n1869), .B(n5098), .Z(n1870) );
  XNOR U3005 ( .A(n5099), .B(n1870), .Z(out[1241]) );
  NANDN U3006 ( .A(n1871), .B(n5101), .Z(n1872) );
  XNOR U3007 ( .A(n5102), .B(n1872), .Z(out[1242]) );
  NANDN U3008 ( .A(n1873), .B(n5104), .Z(n1874) );
  XNOR U3009 ( .A(n5105), .B(n1874), .Z(out[1243]) );
  OR U3010 ( .A(n5108), .B(n1875), .Z(n1876) );
  XNOR U3011 ( .A(n5107), .B(n1876), .Z(out[1244]) );
  NANDN U3012 ( .A(n1877), .B(n5111), .Z(n1878) );
  XNOR U3013 ( .A(n5112), .B(n1878), .Z(out[1245]) );
  NANDN U3014 ( .A(n1879), .B(n5118), .Z(n1880) );
  XNOR U3015 ( .A(n5119), .B(n1880), .Z(out[1246]) );
  OR U3016 ( .A(n5122), .B(n1881), .Z(n1882) );
  XNOR U3017 ( .A(n5121), .B(n1882), .Z(out[1247]) );
  OR U3018 ( .A(n5126), .B(n1883), .Z(n1884) );
  XNOR U3019 ( .A(n5125), .B(n1884), .Z(out[1248]) );
  OR U3020 ( .A(n5130), .B(n1885), .Z(n1886) );
  XNOR U3021 ( .A(n5129), .B(n1886), .Z(out[1249]) );
  IV U3022 ( .A(n3122), .Z(n4054) );
  XOR U3023 ( .A(in[595]), .B(n4054), .Z(n2845) );
  IV U3024 ( .A(n1887), .Z(n3913) );
  XOR U3025 ( .A(in[1470]), .B(n3913), .Z(n3761) );
  XNOR U3026 ( .A(in[250]), .B(n4152), .Z(n3763) );
  NANDN U3027 ( .A(n3761), .B(n3763), .Z(n1888) );
  XNOR U3028 ( .A(n2845), .B(n1888), .Z(out[124]) );
  OR U3029 ( .A(n5134), .B(n1889), .Z(n1890) );
  XNOR U3030 ( .A(n5133), .B(n1890), .Z(out[1250]) );
  OR U3031 ( .A(n5138), .B(n1891), .Z(n1892) );
  XNOR U3032 ( .A(n5137), .B(n1892), .Z(out[1251]) );
  OR U3033 ( .A(n5142), .B(n1893), .Z(n1894) );
  XNOR U3034 ( .A(n5141), .B(n1894), .Z(out[1252]) );
  OR U3035 ( .A(n5146), .B(n1895), .Z(n1896) );
  XNOR U3036 ( .A(n5145), .B(n1896), .Z(out[1253]) );
  OR U3037 ( .A(n5149), .B(n1897), .Z(n1898) );
  XOR U3038 ( .A(n5150), .B(n1898), .Z(out[1254]) );
  OR U3039 ( .A(n5154), .B(n1899), .Z(n1900) );
  XNOR U3040 ( .A(n5153), .B(n1900), .Z(out[1255]) );
  ANDN U3041 ( .B(n1902), .A(n1901), .Z(n1903) );
  XOR U3042 ( .A(n1904), .B(n1903), .Z(out[1256]) );
  ANDN U3043 ( .B(n1906), .A(n1905), .Z(n1907) );
  XOR U3044 ( .A(n1908), .B(n1907), .Z(out[1257]) );
  ANDN U3045 ( .B(n1910), .A(n1909), .Z(n1911) );
  XOR U3046 ( .A(n1912), .B(n1911), .Z(out[1258]) );
  ANDN U3047 ( .B(n1914), .A(n1913), .Z(n1915) );
  XOR U3048 ( .A(n1916), .B(n1915), .Z(out[1259]) );
  IV U3049 ( .A(n3124), .Z(n4058) );
  XOR U3050 ( .A(in[596]), .B(n4058), .Z(n2847) );
  IV U3051 ( .A(n1917), .Z(n3917) );
  XOR U3052 ( .A(in[1471]), .B(n3917), .Z(n3805) );
  IV U3053 ( .A(n4162), .Z(n3277) );
  XOR U3054 ( .A(in[251]), .B(n3277), .Z(n3807) );
  OR U3055 ( .A(n3805), .B(n3807), .Z(n1918) );
  XNOR U3056 ( .A(n2847), .B(n1918), .Z(out[125]) );
  ANDN U3057 ( .B(n1920), .A(n1919), .Z(n1921) );
  XOR U3058 ( .A(n1922), .B(n1921), .Z(out[1260]) );
  ANDN U3059 ( .B(n1924), .A(n1923), .Z(n1925) );
  XOR U3060 ( .A(n1926), .B(n1925), .Z(out[1261]) );
  ANDN U3061 ( .B(n1928), .A(n1927), .Z(n1929) );
  XOR U3062 ( .A(n1930), .B(n1929), .Z(out[1262]) );
  ANDN U3063 ( .B(n1932), .A(n1931), .Z(n1933) );
  XOR U3064 ( .A(n1934), .B(n1933), .Z(out[1263]) );
  ANDN U3065 ( .B(n1936), .A(n1935), .Z(n1937) );
  XOR U3066 ( .A(n1938), .B(n1937), .Z(out[1264]) );
  ANDN U3067 ( .B(n1940), .A(n1939), .Z(n1941) );
  XOR U3068 ( .A(n1942), .B(n1941), .Z(out[1265]) );
  ANDN U3069 ( .B(n1944), .A(n1943), .Z(n1945) );
  XOR U3070 ( .A(n1946), .B(n1945), .Z(out[1266]) );
  ANDN U3071 ( .B(n1948), .A(n1947), .Z(n1949) );
  XOR U3072 ( .A(n1950), .B(n1949), .Z(out[1267]) );
  ANDN U3073 ( .B(n1952), .A(n1951), .Z(n1953) );
  XOR U3074 ( .A(n1954), .B(n1953), .Z(out[1268]) );
  ANDN U3075 ( .B(n1956), .A(n1955), .Z(n1957) );
  XOR U3076 ( .A(n1958), .B(n1957), .Z(out[1269]) );
  IV U3077 ( .A(n3126), .Z(n4062) );
  XOR U3078 ( .A(in[597]), .B(n4062), .Z(n2849) );
  IV U3079 ( .A(n1959), .Z(n3921) );
  XOR U3080 ( .A(in[1408]), .B(n3921), .Z(n3849) );
  IV U3081 ( .A(n4166), .Z(n3280) );
  XOR U3082 ( .A(in[252]), .B(n3280), .Z(n3851) );
  OR U3083 ( .A(n3849), .B(n3851), .Z(n1960) );
  XNOR U3084 ( .A(n2849), .B(n1960), .Z(out[126]) );
  ANDN U3085 ( .B(n1962), .A(n1961), .Z(n1963) );
  XOR U3086 ( .A(n1964), .B(n1963), .Z(out[1270]) );
  ANDN U3087 ( .B(n1966), .A(n1965), .Z(n1967) );
  XOR U3088 ( .A(n1968), .B(n1967), .Z(out[1271]) );
  ANDN U3089 ( .B(n1970), .A(n1969), .Z(n1971) );
  XOR U3090 ( .A(n1972), .B(n1971), .Z(out[1272]) );
  ANDN U3091 ( .B(n1974), .A(n1973), .Z(n1975) );
  XOR U3092 ( .A(n1976), .B(n1975), .Z(out[1273]) );
  ANDN U3093 ( .B(n1978), .A(n1977), .Z(n1979) );
  XOR U3094 ( .A(n1980), .B(n1979), .Z(out[1274]) );
  ANDN U3095 ( .B(n1982), .A(n1981), .Z(n1983) );
  XOR U3096 ( .A(n1984), .B(n1983), .Z(out[1275]) );
  ANDN U3097 ( .B(n1986), .A(n1985), .Z(n1987) );
  XOR U3098 ( .A(n1988), .B(n1987), .Z(out[1276]) );
  ANDN U3099 ( .B(n1990), .A(n1989), .Z(n1991) );
  XOR U3100 ( .A(n1992), .B(n1991), .Z(out[1277]) );
  ANDN U3101 ( .B(n1994), .A(n1993), .Z(n1995) );
  XOR U3102 ( .A(n1996), .B(n1995), .Z(out[1278]) );
  ANDN U3103 ( .B(n1998), .A(n1997), .Z(n1999) );
  XOR U3104 ( .A(n2000), .B(n1999), .Z(out[1279]) );
  IV U3105 ( .A(n3128), .Z(n4070) );
  XOR U3106 ( .A(in[598]), .B(n4070), .Z(n2851) );
  IV U3107 ( .A(n2001), .Z(n3925) );
  XOR U3108 ( .A(in[1409]), .B(n3925), .Z(n3893) );
  IV U3109 ( .A(n4170), .Z(n3283) );
  XOR U3110 ( .A(in[253]), .B(n3283), .Z(n3895) );
  OR U3111 ( .A(n3893), .B(n3895), .Z(n2002) );
  XNOR U3112 ( .A(n2851), .B(n2002), .Z(out[127]) );
  XOR U3113 ( .A(in[50]), .B(n4315), .Z(n2177) );
  XNOR U3114 ( .A(in[1172]), .B(n3987), .Z(n2433) );
  XNOR U3115 ( .A(in[1536]), .B(n3971), .Z(n2434) );
  NANDN U3116 ( .A(n2433), .B(n2434), .Z(n2003) );
  XNOR U3117 ( .A(n2177), .B(n2003), .Z(out[1280]) );
  XOR U3118 ( .A(in[51]), .B(n4318), .Z(n2179) );
  IV U3119 ( .A(n2004), .Z(n3991) );
  XOR U3120 ( .A(in[1173]), .B(n3991), .Z(n2436) );
  XNOR U3121 ( .A(in[1537]), .B(n3975), .Z(n2094) );
  IV U3122 ( .A(n2094), .Z(n2437) );
  OR U3123 ( .A(n2436), .B(n2437), .Z(n2005) );
  XNOR U3124 ( .A(n2179), .B(n2005), .Z(out[1281]) );
  XOR U3125 ( .A(in[52]), .B(n4321), .Z(n2182) );
  IV U3126 ( .A(n2006), .Z(n3995) );
  XOR U3127 ( .A(in[1174]), .B(n3995), .Z(n2441) );
  XNOR U3128 ( .A(in[1538]), .B(n3982), .Z(n2096) );
  IV U3129 ( .A(n2096), .Z(n2443) );
  OR U3130 ( .A(n2441), .B(n2443), .Z(n2007) );
  XNOR U3131 ( .A(n2182), .B(n2007), .Z(out[1282]) );
  XOR U3132 ( .A(in[53]), .B(n4324), .Z(n2184) );
  XNOR U3133 ( .A(in[1175]), .B(n3999), .Z(n2445) );
  XNOR U3134 ( .A(in[1539]), .B(n3986), .Z(n2446) );
  NANDN U3135 ( .A(n2445), .B(n2446), .Z(n2008) );
  XNOR U3136 ( .A(n2184), .B(n2008), .Z(out[1283]) );
  XOR U3137 ( .A(in[54]), .B(n4327), .Z(n2186) );
  XNOR U3138 ( .A(in[1176]), .B(n4003), .Z(n2452) );
  XOR U3139 ( .A(in[1540]), .B(n2009), .Z(n2450) );
  NANDN U3140 ( .A(n2452), .B(n2450), .Z(n2010) );
  XNOR U3141 ( .A(n2186), .B(n2010), .Z(out[1284]) );
  XOR U3142 ( .A(in[55]), .B(n4330), .Z(n2188) );
  XNOR U3143 ( .A(in[1177]), .B(n4007), .Z(n2455) );
  XOR U3144 ( .A(in[1541]), .B(n2011), .Z(n2453) );
  NANDN U3145 ( .A(n2455), .B(n2453), .Z(n2012) );
  XNOR U3146 ( .A(n2188), .B(n2012), .Z(out[1285]) );
  XOR U3147 ( .A(in[56]), .B(n4176), .Z(n2190) );
  IV U3148 ( .A(n2013), .Z(n4011) );
  XOR U3149 ( .A(in[1178]), .B(n4011), .Z(n2457) );
  XOR U3150 ( .A(in[1542]), .B(n2014), .Z(n2102) );
  IV U3151 ( .A(n2102), .Z(n2459) );
  OR U3152 ( .A(n2457), .B(n2459), .Z(n2015) );
  XNOR U3153 ( .A(n2190), .B(n2015), .Z(out[1286]) );
  XOR U3154 ( .A(in[57]), .B(n4179), .Z(n2192) );
  IV U3155 ( .A(n2016), .Z(n4015) );
  XOR U3156 ( .A(in[1179]), .B(n4015), .Z(n2461) );
  XOR U3157 ( .A(in[1543]), .B(n2017), .Z(n2104) );
  IV U3158 ( .A(n2104), .Z(n2462) );
  OR U3159 ( .A(n2461), .B(n2462), .Z(n2018) );
  XNOR U3160 ( .A(n2192), .B(n2018), .Z(out[1287]) );
  XOR U3161 ( .A(in[58]), .B(n4182), .Z(n2194) );
  XNOR U3162 ( .A(in[1180]), .B(n4019), .Z(n2467) );
  XOR U3163 ( .A(in[1544]), .B(n2019), .Z(n2465) );
  NANDN U3164 ( .A(n2467), .B(n2465), .Z(n2020) );
  XNOR U3165 ( .A(n2194), .B(n2020), .Z(out[1288]) );
  XOR U3166 ( .A(in[59]), .B(n4185), .Z(n2196) );
  XNOR U3167 ( .A(in[1181]), .B(n4027), .Z(n2470) );
  XOR U3168 ( .A(in[1545]), .B(n2021), .Z(n2468) );
  NANDN U3169 ( .A(n2470), .B(n2468), .Z(n2022) );
  XNOR U3170 ( .A(n2196), .B(n2022), .Z(out[1289]) );
  XOR U3171 ( .A(in[665]), .B(n4253), .Z(n2853) );
  IV U3172 ( .A(n3130), .Z(n4074) );
  XOR U3173 ( .A(in[599]), .B(n4074), .Z(n3938) );
  OR U3174 ( .A(n3938), .B(n3936), .Z(n2023) );
  XNOR U3175 ( .A(n2853), .B(n2023), .Z(out[128]) );
  XOR U3176 ( .A(in[60]), .B(n3057), .Z(n2198) );
  XNOR U3177 ( .A(in[1182]), .B(n4031), .Z(n2473) );
  XOR U3178 ( .A(in[1546]), .B(n2024), .Z(n2471) );
  NANDN U3179 ( .A(n2473), .B(n2471), .Z(n2025) );
  XNOR U3180 ( .A(n2198), .B(n2025), .Z(out[1290]) );
  XOR U3181 ( .A(in[61]), .B(n3059), .Z(n2200) );
  XNOR U3182 ( .A(in[1183]), .B(n4035), .Z(n2476) );
  XOR U3183 ( .A(in[1547]), .B(n2026), .Z(n2474) );
  NANDN U3184 ( .A(n2476), .B(n2474), .Z(n2027) );
  XNOR U3185 ( .A(n2200), .B(n2027), .Z(out[1291]) );
  XOR U3186 ( .A(in[62]), .B(n3061), .Z(n2203) );
  XNOR U3187 ( .A(in[1184]), .B(n4039), .Z(n2479) );
  XOR U3188 ( .A(in[1548]), .B(n2028), .Z(n2477) );
  NANDN U3189 ( .A(n2479), .B(n2477), .Z(n2029) );
  XNOR U3190 ( .A(n2203), .B(n2029), .Z(out[1292]) );
  XOR U3191 ( .A(in[63]), .B(n4197), .Z(n2205) );
  XNOR U3192 ( .A(in[1185]), .B(n4043), .Z(n2482) );
  XOR U3193 ( .A(in[1549]), .B(n3108), .Z(n2480) );
  NANDN U3194 ( .A(n2482), .B(n2480), .Z(n2030) );
  XNOR U3195 ( .A(n2205), .B(n2030), .Z(out[1293]) );
  XOR U3196 ( .A(in[0]), .B(n3066), .Z(n2207) );
  XOR U3197 ( .A(in[1550]), .B(n3114), .Z(n2112) );
  IV U3198 ( .A(n2112), .Z(n2487) );
  XNOR U3199 ( .A(n3393), .B(in[1186]), .Z(n2484) );
  NANDN U3200 ( .A(n2487), .B(n2484), .Z(n2031) );
  XNOR U3201 ( .A(n2207), .B(n2031), .Z(out[1294]) );
  XOR U3202 ( .A(in[1]), .B(n3069), .Z(n2209) );
  XOR U3203 ( .A(in[1551]), .B(n4038), .Z(n2490) );
  XNOR U3204 ( .A(n3396), .B(in[1187]), .Z(n2488) );
  NANDN U3205 ( .A(n2490), .B(n2488), .Z(n2032) );
  XNOR U3206 ( .A(n2209), .B(n2032), .Z(out[1295]) );
  XOR U3207 ( .A(in[2]), .B(n3071), .Z(n2212) );
  XOR U3208 ( .A(n3400), .B(in[1188]), .Z(n2494) );
  XOR U3209 ( .A(in[1552]), .B(n4042), .Z(n2496) );
  OR U3210 ( .A(n2494), .B(n2496), .Z(n2033) );
  XNOR U3211 ( .A(n2212), .B(n2033), .Z(out[1296]) );
  XOR U3212 ( .A(in[3]), .B(n3075), .Z(n2214) );
  XOR U3213 ( .A(n3404), .B(in[1189]), .Z(n2498) );
  XNOR U3214 ( .A(in[1553]), .B(n4046), .Z(n2500) );
  OR U3215 ( .A(n2498), .B(n2500), .Z(n2034) );
  XNOR U3216 ( .A(n2214), .B(n2034), .Z(out[1297]) );
  XOR U3217 ( .A(in[4]), .B(n3077), .Z(n2216) );
  IV U3218 ( .A(n2035), .Z(n4063) );
  XOR U3219 ( .A(in[1190]), .B(n4063), .Z(n2502) );
  XOR U3220 ( .A(in[1554]), .B(n2036), .Z(n2117) );
  IV U3221 ( .A(n2117), .Z(n2504) );
  OR U3222 ( .A(n2502), .B(n2504), .Z(n2037) );
  XNOR U3223 ( .A(n2216), .B(n2037), .Z(out[1298]) );
  XOR U3224 ( .A(in[5]), .B(n3079), .Z(n2218) );
  IV U3225 ( .A(n2038), .Z(n4071) );
  XOR U3226 ( .A(in[1191]), .B(n4071), .Z(n2506) );
  XOR U3227 ( .A(in[1555]), .B(n4054), .Z(n2508) );
  OR U3228 ( .A(n2506), .B(n2508), .Z(n2039) );
  XNOR U3229 ( .A(n2218), .B(n2039), .Z(out[1299]) );
  XOR U3230 ( .A(in[666]), .B(n4254), .Z(n2856) );
  IV U3231 ( .A(n3136), .Z(n4078) );
  XOR U3232 ( .A(in[600]), .B(n4078), .Z(n3981) );
  XNOR U3233 ( .A(in[255]), .B(n3289), .Z(n3980) );
  NANDN U3234 ( .A(n3981), .B(n3980), .Z(n2040) );
  XNOR U3235 ( .A(n2856), .B(n2040), .Z(out[129]) );
  XNOR U3236 ( .A(in[202]), .B(n3944), .Z(n4337) );
  XOR U3237 ( .A(in[1422]), .B(n3197), .Z(n4338) );
  XNOR U3238 ( .A(in[1045]), .B(n4489), .Z(n2883) );
  NANDN U3239 ( .A(n4338), .B(n2883), .Z(n2041) );
  XNOR U3240 ( .A(n4337), .B(n2041), .Z(out[12]) );
  XOR U3241 ( .A(in[6]), .B(n3081), .Z(n2220) );
  IV U3242 ( .A(n2042), .Z(n4075) );
  XOR U3243 ( .A(in[1192]), .B(n4075), .Z(n2510) );
  XOR U3244 ( .A(in[1556]), .B(n4058), .Z(n2512) );
  OR U3245 ( .A(n2510), .B(n2512), .Z(n2043) );
  XNOR U3246 ( .A(n2220), .B(n2043), .Z(out[1300]) );
  XOR U3247 ( .A(in[7]), .B(n3083), .Z(n2222) );
  IV U3248 ( .A(n2044), .Z(n4079) );
  XOR U3249 ( .A(in[1193]), .B(n4079), .Z(n2514) );
  XOR U3250 ( .A(in[1557]), .B(n3126), .Z(n2119) );
  IV U3251 ( .A(n2119), .Z(n2516) );
  OR U3252 ( .A(n2514), .B(n2516), .Z(n2045) );
  XNOR U3253 ( .A(n2222), .B(n2045), .Z(out[1301]) );
  XOR U3254 ( .A(in[8]), .B(n4214), .Z(n2225) );
  IV U3255 ( .A(n2046), .Z(n4083) );
  XOR U3256 ( .A(in[1194]), .B(n4083), .Z(n2518) );
  XOR U3257 ( .A(in[1558]), .B(n3128), .Z(n2121) );
  IV U3258 ( .A(n2121), .Z(n2520) );
  OR U3259 ( .A(n2518), .B(n2520), .Z(n2047) );
  XNOR U3260 ( .A(n2225), .B(n2047), .Z(out[1302]) );
  XOR U3261 ( .A(in[9]), .B(n3086), .Z(n2227) );
  XOR U3262 ( .A(in[1559]), .B(n3130), .Z(n2123) );
  IV U3263 ( .A(n2123), .Z(n2524) );
  XOR U3264 ( .A(in[1195]), .B(n4088), .Z(n2522) );
  NANDN U3265 ( .A(n2524), .B(n2522), .Z(n2048) );
  XNOR U3266 ( .A(n2227), .B(n2048), .Z(out[1303]) );
  XOR U3267 ( .A(in[10]), .B(n3088), .Z(n2229) );
  XOR U3268 ( .A(in[1560]), .B(n4078), .Z(n2529) );
  XOR U3269 ( .A(in[1196]), .B(n4092), .Z(n2527) );
  NANDN U3270 ( .A(n2529), .B(n2527), .Z(n2049) );
  XNOR U3271 ( .A(n2229), .B(n2049), .Z(out[1304]) );
  XOR U3272 ( .A(in[11]), .B(n3090), .Z(n2231) );
  IV U3273 ( .A(n3138), .Z(n4082) );
  XOR U3274 ( .A(in[1561]), .B(n4082), .Z(n2533) );
  XOR U3275 ( .A(in[1197]), .B(n4096), .Z(n2531) );
  NANDN U3276 ( .A(n2533), .B(n2531), .Z(n2050) );
  XNOR U3277 ( .A(n2231), .B(n2050), .Z(out[1305]) );
  XOR U3278 ( .A(in[12]), .B(n3092), .Z(n2233) );
  IV U3279 ( .A(n3141), .Z(n4086) );
  XOR U3280 ( .A(in[1562]), .B(n4086), .Z(n2537) );
  XOR U3281 ( .A(in[1198]), .B(n4100), .Z(n2535) );
  NANDN U3282 ( .A(n2537), .B(n2535), .Z(n2051) );
  XNOR U3283 ( .A(n2233), .B(n2051), .Z(out[1306]) );
  XOR U3284 ( .A(in[13]), .B(n3096), .Z(n2235) );
  IV U3285 ( .A(n3143), .Z(n4090) );
  XOR U3286 ( .A(in[1563]), .B(n4090), .Z(n2541) );
  XOR U3287 ( .A(in[1199]), .B(n4104), .Z(n2539) );
  NANDN U3288 ( .A(n2541), .B(n2539), .Z(n2052) );
  XNOR U3289 ( .A(n2235), .B(n2052), .Z(out[1307]) );
  XOR U3290 ( .A(in[14]), .B(n4232), .Z(n2237) );
  IV U3291 ( .A(n3022), .Z(n4094) );
  XOR U3292 ( .A(in[1564]), .B(n4094), .Z(n2545) );
  XOR U3293 ( .A(in[1200]), .B(n4108), .Z(n2543) );
  NANDN U3294 ( .A(n2545), .B(n2543), .Z(n2053) );
  XNOR U3295 ( .A(n2237), .B(n2053), .Z(out[1308]) );
  XOR U3296 ( .A(in[15]), .B(n4235), .Z(n2239) );
  IV U3297 ( .A(n3024), .Z(n4098) );
  XOR U3298 ( .A(in[1565]), .B(n4098), .Z(n2549) );
  XOR U3299 ( .A(in[1201]), .B(n4116), .Z(n2547) );
  NANDN U3300 ( .A(n2549), .B(n2547), .Z(n2054) );
  XNOR U3301 ( .A(n2239), .B(n2054), .Z(out[1309]) );
  XOR U3302 ( .A(in[667]), .B(n4255), .Z(n2742) );
  IV U3303 ( .A(n2742), .Z(n2858) );
  XOR U3304 ( .A(in[601]), .B(n4082), .Z(n4025) );
  XNOR U3305 ( .A(in[192]), .B(n3292), .Z(n4022) );
  NANDN U3306 ( .A(n4025), .B(n4022), .Z(n2055) );
  XOR U3307 ( .A(n2858), .B(n2055), .Z(out[130]) );
  XOR U3308 ( .A(in[16]), .B(n4238), .Z(n2241) );
  IV U3309 ( .A(n3026), .Z(n4102) );
  XOR U3310 ( .A(in[1566]), .B(n4102), .Z(n2553) );
  XOR U3311 ( .A(in[1202]), .B(n4120), .Z(n2551) );
  NANDN U3312 ( .A(n2553), .B(n2551), .Z(n2056) );
  XNOR U3313 ( .A(n2241), .B(n2056), .Z(out[1310]) );
  XOR U3314 ( .A(in[17]), .B(n4239), .Z(n2243) );
  IV U3315 ( .A(n3028), .Z(n4106) );
  XOR U3316 ( .A(in[1567]), .B(n4106), .Z(n2556) );
  XOR U3317 ( .A(in[1203]), .B(n4124), .Z(n2555) );
  NANDN U3318 ( .A(n2556), .B(n2555), .Z(n2057) );
  XNOR U3319 ( .A(n2243), .B(n2057), .Z(out[1311]) );
  XOR U3320 ( .A(in[18]), .B(n3102), .Z(n2246) );
  IV U3321 ( .A(n3030), .Z(n4114) );
  XOR U3322 ( .A(in[1568]), .B(n4114), .Z(n2562) );
  XOR U3323 ( .A(in[1204]), .B(n4128), .Z(n2560) );
  NANDN U3324 ( .A(n2562), .B(n2560), .Z(n2058) );
  XNOR U3325 ( .A(n2246), .B(n2058), .Z(out[1312]) );
  XOR U3326 ( .A(in[19]), .B(n3104), .Z(n2248) );
  XOR U3327 ( .A(in[1569]), .B(n3032), .Z(n2127) );
  IV U3328 ( .A(n2127), .Z(n2566) );
  XOR U3329 ( .A(in[1205]), .B(n4132), .Z(n2564) );
  NANDN U3330 ( .A(n2566), .B(n2564), .Z(n2059) );
  XNOR U3331 ( .A(n2248), .B(n2059), .Z(out[1313]) );
  XOR U3332 ( .A(in[20]), .B(n4246), .Z(n2250) );
  XNOR U3333 ( .A(in[1570]), .B(n4122), .Z(n2572) );
  XOR U3334 ( .A(in[1206]), .B(n4136), .Z(n2570) );
  NANDN U3335 ( .A(n2572), .B(n2570), .Z(n2060) );
  XNOR U3336 ( .A(n2250), .B(n2060), .Z(out[1314]) );
  XOR U3337 ( .A(in[21]), .B(n4249), .Z(n2252) );
  XOR U3338 ( .A(in[1571]), .B(n3035), .Z(n2129) );
  IV U3339 ( .A(n2129), .Z(n2576) );
  XOR U3340 ( .A(in[1207]), .B(n4140), .Z(n2574) );
  NANDN U3341 ( .A(n2576), .B(n2574), .Z(n2061) );
  XNOR U3342 ( .A(n2252), .B(n2061), .Z(out[1315]) );
  XOR U3343 ( .A(in[22]), .B(n4250), .Z(n2254) );
  XOR U3344 ( .A(in[1572]), .B(n3037), .Z(n2132) );
  IV U3345 ( .A(n2132), .Z(n2580) );
  XOR U3346 ( .A(in[1208]), .B(n4144), .Z(n2578) );
  NANDN U3347 ( .A(n2580), .B(n2578), .Z(n2062) );
  XNOR U3348 ( .A(n2254), .B(n2062), .Z(out[1316]) );
  XOR U3349 ( .A(in[23]), .B(n4251), .Z(n2256) );
  XNOR U3350 ( .A(in[1573]), .B(n4134), .Z(n2134) );
  IV U3351 ( .A(n2134), .Z(n2584) );
  XOR U3352 ( .A(in[1209]), .B(n4148), .Z(n2582) );
  NANDN U3353 ( .A(n2584), .B(n2582), .Z(n2063) );
  XNOR U3354 ( .A(n2256), .B(n2063), .Z(out[1317]) );
  XOR U3355 ( .A(in[24]), .B(n4252), .Z(n2258) );
  XNOR U3356 ( .A(in[1574]), .B(n4138), .Z(n2588) );
  XOR U3357 ( .A(in[1210]), .B(n4152), .Z(n2586) );
  NAND U3358 ( .A(n2588), .B(n2586), .Z(n2064) );
  XNOR U3359 ( .A(n2258), .B(n2064), .Z(out[1318]) );
  XOR U3360 ( .A(in[25]), .B(n4253), .Z(n2260) );
  XOR U3361 ( .A(in[1211]), .B(n4162), .Z(n2590) );
  XNOR U3362 ( .A(in[1575]), .B(n4142), .Z(n2137) );
  IV U3363 ( .A(n2137), .Z(n2592) );
  OR U3364 ( .A(n2590), .B(n2592), .Z(n2065) );
  XNOR U3365 ( .A(n2260), .B(n2065), .Z(out[1319]) );
  XOR U3366 ( .A(in[668]), .B(n4258), .Z(n2744) );
  IV U3367 ( .A(n2744), .Z(n2860) );
  XOR U3368 ( .A(in[602]), .B(n4086), .Z(n4069) );
  XNOR U3369 ( .A(in[193]), .B(n3295), .Z(n4066) );
  NANDN U3370 ( .A(n4069), .B(n4066), .Z(n2066) );
  XOR U3371 ( .A(n2860), .B(n2066), .Z(out[131]) );
  XOR U3372 ( .A(in[26]), .B(n4254), .Z(n2262) );
  XOR U3373 ( .A(in[1212]), .B(n4166), .Z(n2594) );
  XNOR U3374 ( .A(in[1576]), .B(n4146), .Z(n2139) );
  IV U3375 ( .A(n2139), .Z(n2596) );
  OR U3376 ( .A(n2594), .B(n2596), .Z(n2067) );
  XNOR U3377 ( .A(n2262), .B(n2067), .Z(out[1320]) );
  XOR U3378 ( .A(in[27]), .B(n4255), .Z(n2264) );
  XOR U3379 ( .A(in[1213]), .B(n4170), .Z(n2598) );
  XNOR U3380 ( .A(in[1577]), .B(n4150), .Z(n2141) );
  IV U3381 ( .A(n2141), .Z(n2600) );
  OR U3382 ( .A(n2598), .B(n2600), .Z(n2068) );
  XNOR U3383 ( .A(n2264), .B(n2068), .Z(out[1321]) );
  XOR U3384 ( .A(in[28]), .B(n4258), .Z(n2267) );
  XNOR U3385 ( .A(in[1578]), .B(n4160), .Z(n2143) );
  IV U3386 ( .A(n2143), .Z(n2604) );
  XOR U3387 ( .A(in[1214]), .B(n4174), .Z(n2602) );
  NANDN U3388 ( .A(n2604), .B(n2602), .Z(n2069) );
  XNOR U3389 ( .A(n2267), .B(n2069), .Z(out[1322]) );
  XOR U3390 ( .A(in[29]), .B(n4259), .Z(n2269) );
  XOR U3391 ( .A(in[1215]), .B(n3289), .Z(n2606) );
  XNOR U3392 ( .A(in[1579]), .B(n4164), .Z(n2145) );
  IV U3393 ( .A(n2145), .Z(n2608) );
  OR U3394 ( .A(n2606), .B(n2608), .Z(n2070) );
  XNOR U3395 ( .A(n2269), .B(n2070), .Z(out[1323]) );
  XOR U3396 ( .A(in[30]), .B(n4260), .Z(n2271) );
  XOR U3397 ( .A(in[1152]), .B(n3292), .Z(n2612) );
  XNOR U3398 ( .A(in[1580]), .B(n4168), .Z(n2147) );
  IV U3399 ( .A(n2147), .Z(n2614) );
  OR U3400 ( .A(n2612), .B(n2614), .Z(n2071) );
  XNOR U3401 ( .A(n2271), .B(n2071), .Z(out[1324]) );
  XOR U3402 ( .A(in[31]), .B(n4261), .Z(n2273) );
  XOR U3403 ( .A(in[1153]), .B(n3295), .Z(n2616) );
  XNOR U3404 ( .A(in[1581]), .B(n4172), .Z(n2149) );
  IV U3405 ( .A(n2149), .Z(n2618) );
  OR U3406 ( .A(n2616), .B(n2618), .Z(n2072) );
  XNOR U3407 ( .A(n2273), .B(n2072), .Z(out[1325]) );
  XOR U3408 ( .A(in[32]), .B(n4264), .Z(n2275) );
  XOR U3409 ( .A(in[1154]), .B(n3302), .Z(n2620) );
  XNOR U3410 ( .A(in[1582]), .B(n3896), .Z(n2152) );
  IV U3411 ( .A(n2152), .Z(n2622) );
  OR U3412 ( .A(n2620), .B(n2622), .Z(n2073) );
  XNOR U3413 ( .A(n2275), .B(n2073), .Z(out[1326]) );
  XOR U3414 ( .A(in[33]), .B(n4267), .Z(n2277) );
  XOR U3415 ( .A(in[1155]), .B(n3305), .Z(n2624) );
  XNOR U3416 ( .A(in[1583]), .B(n3900), .Z(n2154) );
  IV U3417 ( .A(n2154), .Z(n2626) );
  OR U3418 ( .A(n2624), .B(n2626), .Z(n2074) );
  XNOR U3419 ( .A(n2277), .B(n2074), .Z(out[1327]) );
  XOR U3420 ( .A(in[34]), .B(n4270), .Z(n2279) );
  XOR U3421 ( .A(in[1156]), .B(n3308), .Z(n2628) );
  XNOR U3422 ( .A(in[1584]), .B(n3904), .Z(n2156) );
  IV U3423 ( .A(n2156), .Z(n2630) );
  OR U3424 ( .A(n2628), .B(n2630), .Z(n2075) );
  XNOR U3425 ( .A(n2279), .B(n2075), .Z(out[1328]) );
  IV U3426 ( .A(n4273), .Z(n3140) );
  XOR U3427 ( .A(in[35]), .B(n3140), .Z(n2281) );
  XOR U3428 ( .A(in[1157]), .B(n3311), .Z(n2632) );
  XNOR U3429 ( .A(in[1585]), .B(n3908), .Z(n2158) );
  IV U3430 ( .A(n2158), .Z(n2634) );
  OR U3431 ( .A(n2632), .B(n2634), .Z(n2076) );
  XNOR U3432 ( .A(n2281), .B(n2076), .Z(out[1329]) );
  XOR U3433 ( .A(in[669]), .B(n4259), .Z(n2746) );
  IV U3434 ( .A(n2746), .Z(n2865) );
  XOR U3435 ( .A(in[603]), .B(n4090), .Z(n4113) );
  XNOR U3436 ( .A(in[194]), .B(n3302), .Z(n4110) );
  NANDN U3437 ( .A(n4113), .B(n4110), .Z(n2077) );
  XOR U3438 ( .A(n2865), .B(n2077), .Z(out[132]) );
  XOR U3439 ( .A(in[36]), .B(n4276), .Z(n2283) );
  XOR U3440 ( .A(in[1158]), .B(n3314), .Z(n2636) );
  XNOR U3441 ( .A(in[1586]), .B(n3912), .Z(n2160) );
  IV U3442 ( .A(n2160), .Z(n2638) );
  OR U3443 ( .A(n2636), .B(n2638), .Z(n2078) );
  XNOR U3444 ( .A(n2283), .B(n2078), .Z(out[1330]) );
  XOR U3445 ( .A(in[37]), .B(n4278), .Z(n2285) );
  XOR U3446 ( .A(in[1159]), .B(n3317), .Z(n2640) );
  XOR U3447 ( .A(in[1587]), .B(n2567), .Z(n2642) );
  OR U3448 ( .A(n2640), .B(n2642), .Z(n2079) );
  XNOR U3449 ( .A(n2285), .B(n2079), .Z(out[1331]) );
  XOR U3450 ( .A(in[38]), .B(n4284), .Z(n2288) );
  XOR U3451 ( .A(in[1160]), .B(n3933), .Z(n2644) );
  XOR U3452 ( .A(in[1588]), .B(n2609), .Z(n2646) );
  OR U3453 ( .A(n2644), .B(n2646), .Z(n2080) );
  XNOR U3454 ( .A(n2288), .B(n2080), .Z(out[1332]) );
  XOR U3455 ( .A(in[39]), .B(n4286), .Z(n2290) );
  XOR U3456 ( .A(in[1161]), .B(n3940), .Z(n2648) );
  XOR U3457 ( .A(in[1589]), .B(n2651), .Z(n2650) );
  OR U3458 ( .A(n2648), .B(n2650), .Z(n2081) );
  XNOR U3459 ( .A(n2290), .B(n2081), .Z(out[1333]) );
  XOR U3460 ( .A(in[40]), .B(n4288), .Z(n2293) );
  XOR U3461 ( .A(in[1162]), .B(n3944), .Z(n2654) );
  XNOR U3462 ( .A(in[1590]), .B(n3063), .Z(n2656) );
  NANDN U3463 ( .A(n2654), .B(n2656), .Z(n2082) );
  XNOR U3464 ( .A(n2293), .B(n2082), .Z(out[1334]) );
  XOR U3465 ( .A(in[41]), .B(n4290), .Z(n2295) );
  XOR U3466 ( .A(in[1163]), .B(n3948), .Z(n2658) );
  XNOR U3467 ( .A(in[1591]), .B(n3065), .Z(n2660) );
  NANDN U3468 ( .A(n2658), .B(n2660), .Z(n2083) );
  XNOR U3469 ( .A(n2295), .B(n2083), .Z(out[1335]) );
  XOR U3470 ( .A(in[42]), .B(n4292), .Z(n2297) );
  XOR U3471 ( .A(in[1164]), .B(n3952), .Z(n2662) );
  XNOR U3472 ( .A(in[1592]), .B(n3068), .Z(n2664) );
  NANDN U3473 ( .A(n2662), .B(n2664), .Z(n2084) );
  XNOR U3474 ( .A(n2297), .B(n2084), .Z(out[1336]) );
  XOR U3475 ( .A(in[43]), .B(n4294), .Z(n2299) );
  XOR U3476 ( .A(in[1165]), .B(n3956), .Z(n2666) );
  XOR U3477 ( .A(in[1593]), .B(n2698), .Z(n2668) );
  OR U3478 ( .A(n2666), .B(n2668), .Z(n2085) );
  XNOR U3479 ( .A(n2299), .B(n2085), .Z(out[1337]) );
  XOR U3480 ( .A(in[44]), .B(n4296), .Z(n2301) );
  XOR U3481 ( .A(in[1166]), .B(n3960), .Z(n2670) );
  XOR U3482 ( .A(in[1594]), .B(n2700), .Z(n2672) );
  OR U3483 ( .A(n2670), .B(n2672), .Z(n2086) );
  XNOR U3484 ( .A(n2301), .B(n2086), .Z(out[1338]) );
  XOR U3485 ( .A(in[45]), .B(n4298), .Z(n2303) );
  XOR U3486 ( .A(in[1167]), .B(n3964), .Z(n2674) );
  XNOR U3487 ( .A(in[1595]), .B(n3951), .Z(n2167) );
  IV U3488 ( .A(n2167), .Z(n2676) );
  OR U3489 ( .A(n2674), .B(n2676), .Z(n2087) );
  XNOR U3490 ( .A(n2303), .B(n2087), .Z(out[1339]) );
  XOR U3491 ( .A(in[670]), .B(n4260), .Z(n2748) );
  IV U3492 ( .A(n2748), .Z(n2867) );
  XOR U3493 ( .A(in[604]), .B(n4094), .Z(n4157) );
  XNOR U3494 ( .A(in[195]), .B(n3305), .Z(n4154) );
  NANDN U3495 ( .A(n4157), .B(n4154), .Z(n2088) );
  XOR U3496 ( .A(n2867), .B(n2088), .Z(out[133]) );
  XOR U3497 ( .A(in[46]), .B(n4300), .Z(n2305) );
  XOR U3498 ( .A(in[1168]), .B(n3968), .Z(n2678) );
  XNOR U3499 ( .A(in[1596]), .B(n3955), .Z(n2169) );
  IV U3500 ( .A(n2169), .Z(n2680) );
  OR U3501 ( .A(n2678), .B(n2680), .Z(n2089) );
  XNOR U3502 ( .A(n2305), .B(n2089), .Z(out[1340]) );
  XOR U3503 ( .A(in[47]), .B(n4302), .Z(n2307) );
  XOR U3504 ( .A(in[1169]), .B(n3972), .Z(n2682) );
  XNOR U3505 ( .A(in[1597]), .B(n3959), .Z(n2171) );
  IV U3506 ( .A(n2171), .Z(n2684) );
  OR U3507 ( .A(n2682), .B(n2684), .Z(n2090) );
  XNOR U3508 ( .A(n2307), .B(n2090), .Z(out[1341]) );
  XOR U3509 ( .A(in[48]), .B(n4309), .Z(n2310) );
  XOR U3510 ( .A(in[1170]), .B(n3976), .Z(n2686) );
  XNOR U3511 ( .A(in[1598]), .B(n3963), .Z(n2173) );
  IV U3512 ( .A(n2173), .Z(n2688) );
  OR U3513 ( .A(n2686), .B(n2688), .Z(n2091) );
  XNOR U3514 ( .A(n2310), .B(n2091), .Z(out[1342]) );
  XOR U3515 ( .A(in[49]), .B(n4312), .Z(n2312) );
  IV U3516 ( .A(n3983), .Z(n3347) );
  XOR U3517 ( .A(in[1171]), .B(n3347), .Z(n2690) );
  XNOR U3518 ( .A(in[1599]), .B(n3967), .Z(n2175) );
  IV U3519 ( .A(n2175), .Z(n2691) );
  OR U3520 ( .A(n2690), .B(n2691), .Z(n2092) );
  XNOR U3521 ( .A(n2312), .B(n2092), .Z(out[1343]) );
  XNOR U3522 ( .A(in[427]), .B(n4345), .Z(n2314) );
  NOR U3523 ( .A(n2434), .B(n2177), .Z(n2093) );
  XNOR U3524 ( .A(n2314), .B(n2093), .Z(out[1344]) );
  XNOR U3525 ( .A(in[428]), .B(n4348), .Z(n2316) );
  NOR U3526 ( .A(n2094), .B(n2179), .Z(n2095) );
  XNOR U3527 ( .A(n2316), .B(n2095), .Z(out[1345]) );
  XNOR U3528 ( .A(in[429]), .B(n4351), .Z(n2318) );
  NOR U3529 ( .A(n2096), .B(n2182), .Z(n2097) );
  XNOR U3530 ( .A(n2318), .B(n2097), .Z(out[1346]) );
  XNOR U3531 ( .A(in[430]), .B(n4354), .Z(n2320) );
  NOR U3532 ( .A(n2446), .B(n2184), .Z(n2098) );
  XNOR U3533 ( .A(n2320), .B(n2098), .Z(out[1347]) );
  XNOR U3534 ( .A(in[431]), .B(n4356), .Z(n2322) );
  NOR U3535 ( .A(n2450), .B(n2186), .Z(n2099) );
  XNOR U3536 ( .A(n2322), .B(n2099), .Z(out[1348]) );
  XNOR U3537 ( .A(in[432]), .B(n4359), .Z(n2324) );
  NOR U3538 ( .A(n2453), .B(n2188), .Z(n2100) );
  XNOR U3539 ( .A(n2324), .B(n2100), .Z(out[1349]) );
  XOR U3540 ( .A(in[671]), .B(n4261), .Z(n2750) );
  IV U3541 ( .A(n2750), .Z(n2869) );
  XOR U3542 ( .A(in[605]), .B(n4098), .Z(n4195) );
  XNOR U3543 ( .A(in[196]), .B(n3308), .Z(n4192) );
  NANDN U3544 ( .A(n4195), .B(n4192), .Z(n2101) );
  XOR U3545 ( .A(n2869), .B(n2101), .Z(out[134]) );
  XNOR U3546 ( .A(in[433]), .B(n4362), .Z(n2326) );
  NOR U3547 ( .A(n2102), .B(n2190), .Z(n2103) );
  XNOR U3548 ( .A(n2326), .B(n2103), .Z(out[1350]) );
  XNOR U3549 ( .A(in[434]), .B(n4365), .Z(n2328) );
  NOR U3550 ( .A(n2104), .B(n2192), .Z(n2105) );
  XNOR U3551 ( .A(n2328), .B(n2105), .Z(out[1351]) );
  XNOR U3552 ( .A(in[435]), .B(n4372), .Z(n2331) );
  NOR U3553 ( .A(n2465), .B(n2194), .Z(n2106) );
  XNOR U3554 ( .A(n2331), .B(n2106), .Z(out[1352]) );
  XNOR U3555 ( .A(in[436]), .B(n4375), .Z(n2334) );
  NOR U3556 ( .A(n2468), .B(n2196), .Z(n2107) );
  XNOR U3557 ( .A(n2334), .B(n2107), .Z(out[1353]) );
  XNOR U3558 ( .A(in[437]), .B(n4378), .Z(n2337) );
  NOR U3559 ( .A(n2471), .B(n2198), .Z(n2108) );
  XNOR U3560 ( .A(n2337), .B(n2108), .Z(out[1354]) );
  XNOR U3561 ( .A(in[438]), .B(n4381), .Z(n2340) );
  NOR U3562 ( .A(n2474), .B(n2200), .Z(n2109) );
  XNOR U3563 ( .A(n2340), .B(n2109), .Z(out[1355]) );
  XNOR U3564 ( .A(in[439]), .B(n4384), .Z(n2343) );
  NOR U3565 ( .A(n2477), .B(n2203), .Z(n2110) );
  XNOR U3566 ( .A(n2343), .B(n2110), .Z(out[1356]) );
  XNOR U3567 ( .A(in[440]), .B(n4386), .Z(n2346) );
  NOR U3568 ( .A(n2480), .B(n2205), .Z(n2111) );
  XNOR U3569 ( .A(n2346), .B(n2111), .Z(out[1357]) );
  XNOR U3570 ( .A(in[441]), .B(n4389), .Z(n2349) );
  NOR U3571 ( .A(n2112), .B(n2207), .Z(n2113) );
  XNOR U3572 ( .A(n2349), .B(n2113), .Z(out[1358]) );
  XOR U3573 ( .A(in[442]), .B(n2114), .Z(n2351) );
  XOR U3574 ( .A(in[672]), .B(n4264), .Z(n2752) );
  IV U3575 ( .A(n2752), .Z(n2871) );
  XOR U3576 ( .A(in[606]), .B(n4102), .Z(n4213) );
  XNOR U3577 ( .A(in[197]), .B(n3311), .Z(n4442) );
  NANDN U3578 ( .A(n4213), .B(n4442), .Z(n2115) );
  XOR U3579 ( .A(n2871), .B(n2115), .Z(out[135]) );
  XOR U3580 ( .A(in[443]), .B(n2116), .Z(n2353) );
  XNOR U3581 ( .A(in[444]), .B(n4398), .Z(n2354) );
  XNOR U3582 ( .A(in[445]), .B(n4405), .Z(n2357) );
  NOR U3583 ( .A(n2117), .B(n2216), .Z(n2118) );
  XNOR U3584 ( .A(n2357), .B(n2118), .Z(out[1362]) );
  XNOR U3585 ( .A(in[446]), .B(n4408), .Z(n2359) );
  XNOR U3586 ( .A(in[447]), .B(n4411), .Z(n2361) );
  XNOR U3587 ( .A(in[384]), .B(n4414), .Z(n2363) );
  NOR U3588 ( .A(n2119), .B(n2222), .Z(n2120) );
  XNOR U3589 ( .A(n2363), .B(n2120), .Z(out[1365]) );
  XNOR U3590 ( .A(in[385]), .B(n4417), .Z(n2365) );
  NOR U3591 ( .A(n2121), .B(n2225), .Z(n2122) );
  XNOR U3592 ( .A(n2365), .B(n2122), .Z(out[1366]) );
  XNOR U3593 ( .A(in[386]), .B(n4420), .Z(n2367) );
  NOR U3594 ( .A(n2123), .B(n2227), .Z(n2124) );
  XNOR U3595 ( .A(n2367), .B(n2124), .Z(out[1367]) );
  XNOR U3596 ( .A(in[387]), .B(n4423), .Z(n2369) );
  XNOR U3597 ( .A(in[388]), .B(n4426), .Z(n2371) );
  XOR U3598 ( .A(in[673]), .B(n4267), .Z(n2759) );
  IV U3599 ( .A(n2759), .Z(n2873) );
  XOR U3600 ( .A(in[607]), .B(n4106), .Z(n4241) );
  XNOR U3601 ( .A(in[198]), .B(n3314), .Z(n4733) );
  NANDN U3602 ( .A(n4241), .B(n4733), .Z(n2125) );
  XOR U3603 ( .A(n2873), .B(n2125), .Z(out[136]) );
  XNOR U3604 ( .A(in[389]), .B(n4429), .Z(n2373) );
  XOR U3605 ( .A(in[390]), .B(n2126), .Z(n2375) );
  XNOR U3606 ( .A(in[391]), .B(n4443), .Z(n2378) );
  XNOR U3607 ( .A(in[392]), .B(n4446), .Z(n2380) );
  XNOR U3608 ( .A(in[393]), .B(n4449), .Z(n2382) );
  XNOR U3609 ( .A(in[394]), .B(n4452), .Z(n2384) );
  XNOR U3610 ( .A(in[395]), .B(n4455), .Z(n2386) );
  XNOR U3611 ( .A(n4458), .B(in[396]), .Z(n2388) );
  NOR U3612 ( .A(n2127), .B(n2248), .Z(n2128) );
  XOR U3613 ( .A(n2388), .B(n2128), .Z(out[1377]) );
  XNOR U3614 ( .A(n4461), .B(in[397]), .Z(n2389) );
  XNOR U3615 ( .A(n4464), .B(in[398]), .Z(n2390) );
  NOR U3616 ( .A(n2129), .B(n2252), .Z(n2130) );
  XOR U3617 ( .A(n2390), .B(n2130), .Z(out[1379]) );
  XOR U3618 ( .A(in[674]), .B(n4270), .Z(n2761) );
  IV U3619 ( .A(n2761), .Z(n2875) );
  XOR U3620 ( .A(in[608]), .B(n4114), .Z(n4257) );
  XNOR U3621 ( .A(in[199]), .B(n3317), .Z(n5164) );
  NANDN U3622 ( .A(n4257), .B(n5164), .Z(n2131) );
  XOR U3623 ( .A(n2875), .B(n2131), .Z(out[137]) );
  XNOR U3624 ( .A(n4467), .B(in[399]), .Z(n2391) );
  NOR U3625 ( .A(n2132), .B(n2254), .Z(n2133) );
  XOR U3626 ( .A(n2391), .B(n2133), .Z(out[1380]) );
  XNOR U3627 ( .A(n4470), .B(in[400]), .Z(n2392) );
  NOR U3628 ( .A(n2134), .B(n2256), .Z(n2135) );
  XOR U3629 ( .A(n2392), .B(n2135), .Z(out[1381]) );
  XNOR U3630 ( .A(n4477), .B(in[401]), .Z(n2394) );
  NOR U3631 ( .A(n2588), .B(n2258), .Z(n2136) );
  XOR U3632 ( .A(n2394), .B(n2136), .Z(out[1382]) );
  XNOR U3633 ( .A(n4480), .B(in[402]), .Z(n2395) );
  NOR U3634 ( .A(n2137), .B(n2260), .Z(n2138) );
  XOR U3635 ( .A(n2395), .B(n2138), .Z(out[1383]) );
  XNOR U3636 ( .A(n4483), .B(in[403]), .Z(n2396) );
  NOR U3637 ( .A(n2139), .B(n2262), .Z(n2140) );
  XOR U3638 ( .A(n2396), .B(n2140), .Z(out[1384]) );
  XNOR U3639 ( .A(in[404]), .B(n4486), .Z(n2397) );
  NOR U3640 ( .A(n2141), .B(n2264), .Z(n2142) );
  XOR U3641 ( .A(n2397), .B(n2142), .Z(out[1385]) );
  XNOR U3642 ( .A(in[405]), .B(n4489), .Z(n2398) );
  NOR U3643 ( .A(n2143), .B(n2267), .Z(n2144) );
  XOR U3644 ( .A(n2398), .B(n2144), .Z(out[1386]) );
  XNOR U3645 ( .A(in[406]), .B(n4492), .Z(n2399) );
  NOR U3646 ( .A(n2145), .B(n2269), .Z(n2146) );
  XOR U3647 ( .A(n2399), .B(n2146), .Z(out[1387]) );
  XNOR U3648 ( .A(in[407]), .B(n4495), .Z(n2400) );
  NOR U3649 ( .A(n2147), .B(n2271), .Z(n2148) );
  XOR U3650 ( .A(n2400), .B(n2148), .Z(out[1388]) );
  XNOR U3651 ( .A(in[408]), .B(n4498), .Z(n2401) );
  NOR U3652 ( .A(n2149), .B(n2273), .Z(n2150) );
  XOR U3653 ( .A(n2401), .B(n2150), .Z(out[1389]) );
  XOR U3654 ( .A(in[675]), .B(n4273), .Z(n2878) );
  IV U3655 ( .A(n3032), .Z(n4118) );
  XOR U3656 ( .A(in[609]), .B(n4118), .Z(n4283) );
  NANDN U3657 ( .A(n4283), .B(n4280), .Z(n2151) );
  XOR U3658 ( .A(n2878), .B(n2151), .Z(out[138]) );
  XNOR U3659 ( .A(in[409]), .B(n4501), .Z(n2402) );
  NOR U3660 ( .A(n2152), .B(n2275), .Z(n2153) );
  XOR U3661 ( .A(n2402), .B(n2153), .Z(out[1390]) );
  XNOR U3662 ( .A(in[410]), .B(n4504), .Z(n2403) );
  NOR U3663 ( .A(n2154), .B(n2277), .Z(n2155) );
  XOR U3664 ( .A(n2403), .B(n2155), .Z(out[1391]) );
  XOR U3665 ( .A(in[411]), .B(n4511), .Z(n2405) );
  NOR U3666 ( .A(n2156), .B(n2279), .Z(n2157) );
  XOR U3667 ( .A(n2405), .B(n2157), .Z(out[1392]) );
  XOR U3668 ( .A(in[412]), .B(n4514), .Z(n2406) );
  NOR U3669 ( .A(n2158), .B(n2281), .Z(n2159) );
  XOR U3670 ( .A(n2406), .B(n2159), .Z(out[1393]) );
  XOR U3671 ( .A(in[413]), .B(n4517), .Z(n2407) );
  NOR U3672 ( .A(n2160), .B(n2283), .Z(n2161) );
  XOR U3673 ( .A(n2407), .B(n2161), .Z(out[1394]) );
  XOR U3674 ( .A(in[414]), .B(n4520), .Z(n2408) );
  XOR U3675 ( .A(in[415]), .B(n4524), .Z(n2410) );
  XOR U3676 ( .A(in[416]), .B(n4528), .Z(n2412) );
  XNOR U3677 ( .A(in[417]), .B(n4532), .Z(n2414) );
  NOR U3678 ( .A(n2656), .B(n2293), .Z(n2162) );
  XOR U3679 ( .A(n2414), .B(n2162), .Z(out[1398]) );
  XNOR U3680 ( .A(in[418]), .B(n4536), .Z(n2415) );
  NOR U3681 ( .A(n2660), .B(n2295), .Z(n2163) );
  XOR U3682 ( .A(n2415), .B(n2163), .Z(out[1399]) );
  XOR U3683 ( .A(in[676]), .B(n4276), .Z(n2880) );
  XNOR U3684 ( .A(in[610]), .B(n4122), .Z(n4308) );
  NANDN U3685 ( .A(n4308), .B(n4305), .Z(n2164) );
  XNOR U3686 ( .A(n2880), .B(n2164), .Z(out[139]) );
  XNOR U3687 ( .A(in[203]), .B(n3948), .Z(n4368) );
  XOR U3688 ( .A(in[1423]), .B(n3200), .Z(n4369) );
  XNOR U3689 ( .A(in[1046]), .B(n4492), .Z(n2885) );
  NANDN U3690 ( .A(n4369), .B(n2885), .Z(n2165) );
  XNOR U3691 ( .A(n4368), .B(n2165), .Z(out[13]) );
  XNOR U3692 ( .A(in[419]), .B(n4540), .Z(n2416) );
  NOR U3693 ( .A(n2664), .B(n2297), .Z(n2166) );
  XOR U3694 ( .A(n2416), .B(n2166), .Z(out[1400]) );
  XNOR U3695 ( .A(in[420]), .B(n4544), .Z(n2417) );
  XNOR U3696 ( .A(in[421]), .B(n4550), .Z(n2420) );
  XNOR U3697 ( .A(in[422]), .B(n4552), .Z(n2422) );
  NOR U3698 ( .A(n2167), .B(n2303), .Z(n2168) );
  XNOR U3699 ( .A(n2422), .B(n2168), .Z(out[1403]) );
  XNOR U3700 ( .A(in[423]), .B(n4333), .Z(n2424) );
  NOR U3701 ( .A(n2169), .B(n2305), .Z(n2170) );
  XNOR U3702 ( .A(n2424), .B(n2170), .Z(out[1404]) );
  XNOR U3703 ( .A(in[424]), .B(n4335), .Z(n2426) );
  NOR U3704 ( .A(n2171), .B(n2307), .Z(n2172) );
  XNOR U3705 ( .A(n2426), .B(n2172), .Z(out[1405]) );
  XNOR U3706 ( .A(in[425]), .B(n4341), .Z(n2428) );
  NOR U3707 ( .A(n2173), .B(n2310), .Z(n2174) );
  XNOR U3708 ( .A(n2428), .B(n2174), .Z(out[1406]) );
  XNOR U3709 ( .A(in[426]), .B(n4343), .Z(n2430) );
  NOR U3710 ( .A(n2175), .B(n2312), .Z(n2176) );
  XNOR U3711 ( .A(n2430), .B(n2176), .Z(out[1407]) );
  XOR U3712 ( .A(in[789]), .B(n4012), .Z(n2432) );
  NAND U3713 ( .A(n2177), .B(n2314), .Z(n2178) );
  XOR U3714 ( .A(n2432), .B(n2178), .Z(out[1408]) );
  IV U3715 ( .A(n2771), .Z(n4016) );
  XOR U3716 ( .A(in[790]), .B(n4016), .Z(n2435) );
  NAND U3717 ( .A(n2179), .B(n2316), .Z(n2180) );
  XOR U3718 ( .A(n2435), .B(n2180), .Z(out[1409]) );
  XOR U3719 ( .A(in[677]), .B(n4278), .Z(n2882) );
  IV U3720 ( .A(n3035), .Z(n4126) );
  XOR U3721 ( .A(in[611]), .B(n4126), .Z(n4340) );
  NANDN U3722 ( .A(n4340), .B(n4337), .Z(n2181) );
  XNOR U3723 ( .A(n2882), .B(n2181), .Z(out[140]) );
  IV U3724 ( .A(n2778), .Z(n4020) );
  XOR U3725 ( .A(in[791]), .B(n4020), .Z(n2440) );
  NAND U3726 ( .A(n2182), .B(n2318), .Z(n2183) );
  XOR U3727 ( .A(n2440), .B(n2183), .Z(out[1410]) );
  IV U3728 ( .A(n2792), .Z(n4028) );
  XOR U3729 ( .A(in[792]), .B(n4028), .Z(n2444) );
  NAND U3730 ( .A(n2184), .B(n2320), .Z(n2185) );
  XOR U3731 ( .A(n2444), .B(n2185), .Z(out[1411]) );
  IV U3732 ( .A(n2815), .Z(n4032) );
  XOR U3733 ( .A(in[793]), .B(n4032), .Z(n2451) );
  NAND U3734 ( .A(n2186), .B(n2322), .Z(n2187) );
  XOR U3735 ( .A(n2451), .B(n2187), .Z(out[1412]) );
  IV U3736 ( .A(n2838), .Z(n4036) );
  XOR U3737 ( .A(in[794]), .B(n4036), .Z(n2454) );
  NAND U3738 ( .A(n2188), .B(n2324), .Z(n2189) );
  XOR U3739 ( .A(n2454), .B(n2189), .Z(out[1413]) );
  IV U3740 ( .A(n2862), .Z(n4040) );
  XOR U3741 ( .A(in[795]), .B(n4040), .Z(n2456) );
  NAND U3742 ( .A(n2190), .B(n2326), .Z(n2191) );
  XOR U3743 ( .A(n2456), .B(n2191), .Z(out[1414]) );
  IV U3744 ( .A(n2886), .Z(n4044) );
  XOR U3745 ( .A(in[796]), .B(n4044), .Z(n2460) );
  NAND U3746 ( .A(n2192), .B(n2328), .Z(n2193) );
  XOR U3747 ( .A(n2460), .B(n2193), .Z(out[1415]) );
  IV U3748 ( .A(n2919), .Z(n4048) );
  XOR U3749 ( .A(in[797]), .B(n4048), .Z(n2466) );
  NAND U3750 ( .A(n2194), .B(n2331), .Z(n2195) );
  XOR U3751 ( .A(n2466), .B(n2195), .Z(out[1416]) );
  XOR U3752 ( .A(in[798]), .B(n4052), .Z(n2333) );
  NAND U3753 ( .A(n2196), .B(n2334), .Z(n2197) );
  XNOR U3754 ( .A(n2333), .B(n2197), .Z(out[1417]) );
  XOR U3755 ( .A(in[799]), .B(n4056), .Z(n2336) );
  NAND U3756 ( .A(n2198), .B(n2337), .Z(n2199) );
  XNOR U3757 ( .A(n2336), .B(n2199), .Z(out[1418]) );
  XOR U3758 ( .A(in[800]), .B(n4060), .Z(n2339) );
  NAND U3759 ( .A(n2200), .B(n2340), .Z(n2201) );
  XNOR U3760 ( .A(n2339), .B(n2201), .Z(out[1419]) );
  XOR U3761 ( .A(in[678]), .B(n4284), .Z(n2884) );
  IV U3762 ( .A(n3037), .Z(n4130) );
  XOR U3763 ( .A(in[612]), .B(n4130), .Z(n4371) );
  NANDN U3764 ( .A(n4371), .B(n4368), .Z(n2202) );
  XNOR U3765 ( .A(n2884), .B(n2202), .Z(out[141]) );
  XOR U3766 ( .A(in[801]), .B(n4064), .Z(n2342) );
  NAND U3767 ( .A(n2203), .B(n2343), .Z(n2204) );
  XNOR U3768 ( .A(n2342), .B(n2204), .Z(out[1420]) );
  XOR U3769 ( .A(in[802]), .B(n4072), .Z(n2345) );
  NAND U3770 ( .A(n2205), .B(n2346), .Z(n2206) );
  XNOR U3771 ( .A(n2345), .B(n2206), .Z(out[1421]) );
  XOR U3772 ( .A(in[803]), .B(n4076), .Z(n2348) );
  NAND U3773 ( .A(n2207), .B(n2349), .Z(n2208) );
  XNOR U3774 ( .A(n2348), .B(n2208), .Z(out[1422]) );
  XOR U3775 ( .A(in[804]), .B(n4080), .Z(n2352) );
  NANDN U3776 ( .A(n2351), .B(n2209), .Z(n2210) );
  XNOR U3777 ( .A(n2352), .B(n2210), .Z(out[1423]) );
  IV U3778 ( .A(n2211), .Z(n4084) );
  XOR U3779 ( .A(in[805]), .B(n4084), .Z(n2493) );
  NANDN U3780 ( .A(n2353), .B(n2212), .Z(n2213) );
  XOR U3781 ( .A(n2493), .B(n2213), .Z(out[1424]) );
  XNOR U3782 ( .A(in[806]), .B(n4087), .Z(n2497) );
  NAND U3783 ( .A(n2214), .B(n2354), .Z(n2215) );
  XNOR U3784 ( .A(n2497), .B(n2215), .Z(out[1425]) );
  XNOR U3785 ( .A(in[807]), .B(n4091), .Z(n2501) );
  NAND U3786 ( .A(n2216), .B(n2357), .Z(n2217) );
  XNOR U3787 ( .A(n2501), .B(n2217), .Z(out[1426]) );
  XNOR U3788 ( .A(in[808]), .B(n4095), .Z(n2505) );
  NAND U3789 ( .A(n2218), .B(n2359), .Z(n2219) );
  XNOR U3790 ( .A(n2505), .B(n2219), .Z(out[1427]) );
  XNOR U3791 ( .A(in[809]), .B(n4099), .Z(n2509) );
  NAND U3792 ( .A(n2220), .B(n2361), .Z(n2221) );
  XNOR U3793 ( .A(n2509), .B(n2221), .Z(out[1428]) );
  XNOR U3794 ( .A(in[810]), .B(n4103), .Z(n2513) );
  NAND U3795 ( .A(n2222), .B(n2363), .Z(n2223) );
  XNOR U3796 ( .A(n2513), .B(n2223), .Z(out[1429]) );
  XOR U3797 ( .A(in[679]), .B(n4286), .Z(n2767) );
  XOR U3798 ( .A(in[613]), .B(n4134), .Z(n4404) );
  XNOR U3799 ( .A(in[204]), .B(n3952), .Z(n4401) );
  NANDN U3800 ( .A(n4404), .B(n4401), .Z(n2224) );
  XNOR U3801 ( .A(n2767), .B(n2224), .Z(out[142]) );
  XNOR U3802 ( .A(in[811]), .B(n4107), .Z(n2517) );
  NAND U3803 ( .A(n2225), .B(n2365), .Z(n2226) );
  XOR U3804 ( .A(n2517), .B(n2226), .Z(out[1430]) );
  XNOR U3805 ( .A(in[812]), .B(n4115), .Z(n2521) );
  NAND U3806 ( .A(n2227), .B(n2367), .Z(n2228) );
  XOR U3807 ( .A(n2521), .B(n2228), .Z(out[1431]) );
  XOR U3808 ( .A(in[813]), .B(n4119), .Z(n2526) );
  NAND U3809 ( .A(n2229), .B(n2369), .Z(n2230) );
  XOR U3810 ( .A(n2526), .B(n2230), .Z(out[1432]) );
  XOR U3811 ( .A(in[814]), .B(n4123), .Z(n2530) );
  NAND U3812 ( .A(n2231), .B(n2371), .Z(n2232) );
  XOR U3813 ( .A(n2530), .B(n2232), .Z(out[1433]) );
  XOR U3814 ( .A(in[815]), .B(n4127), .Z(n2534) );
  NAND U3815 ( .A(n2233), .B(n2373), .Z(n2234) );
  XOR U3816 ( .A(n2534), .B(n2234), .Z(out[1434]) );
  XOR U3817 ( .A(in[816]), .B(n4131), .Z(n2538) );
  NANDN U3818 ( .A(n2375), .B(n2235), .Z(n2236) );
  XOR U3819 ( .A(n2538), .B(n2236), .Z(out[1435]) );
  XOR U3820 ( .A(in[817]), .B(n4135), .Z(n2542) );
  NAND U3821 ( .A(n2237), .B(n2378), .Z(n2238) );
  XOR U3822 ( .A(n2542), .B(n2238), .Z(out[1436]) );
  XOR U3823 ( .A(in[818]), .B(n4139), .Z(n2546) );
  NAND U3824 ( .A(n2239), .B(n2380), .Z(n2240) );
  XOR U3825 ( .A(n2546), .B(n2240), .Z(out[1437]) );
  XOR U3826 ( .A(in[819]), .B(n4143), .Z(n2550) );
  NAND U3827 ( .A(n2241), .B(n2382), .Z(n2242) );
  XOR U3828 ( .A(n2550), .B(n2242), .Z(out[1438]) );
  XOR U3829 ( .A(in[820]), .B(n4147), .Z(n2554) );
  NAND U3830 ( .A(n2243), .B(n2384), .Z(n2244) );
  XOR U3831 ( .A(n2554), .B(n2244), .Z(out[1439]) );
  XOR U3832 ( .A(in[680]), .B(n4288), .Z(n2768) );
  XOR U3833 ( .A(in[614]), .B(n4138), .Z(n4438) );
  XNOR U3834 ( .A(in[205]), .B(n3956), .Z(n4435) );
  NANDN U3835 ( .A(n4438), .B(n4435), .Z(n2245) );
  XNOR U3836 ( .A(n2768), .B(n2245), .Z(out[143]) );
  XNOR U3837 ( .A(in[821]), .B(n4151), .Z(n2559) );
  NAND U3838 ( .A(n2246), .B(n2386), .Z(n2247) );
  XOR U3839 ( .A(n2559), .B(n2247), .Z(out[1440]) );
  XNOR U3840 ( .A(in[822]), .B(n4161), .Z(n2563) );
  NANDN U3841 ( .A(n2388), .B(n2248), .Z(n2249) );
  XOR U3842 ( .A(n2563), .B(n2249), .Z(out[1441]) );
  XNOR U3843 ( .A(in[823]), .B(n4165), .Z(n2569) );
  NANDN U3844 ( .A(n2389), .B(n2250), .Z(n2251) );
  XOR U3845 ( .A(n2569), .B(n2251), .Z(out[1442]) );
  XNOR U3846 ( .A(in[824]), .B(n4169), .Z(n2573) );
  NANDN U3847 ( .A(n2390), .B(n2252), .Z(n2253) );
  XOR U3848 ( .A(n2573), .B(n2253), .Z(out[1443]) );
  XNOR U3849 ( .A(in[825]), .B(n4173), .Z(n2577) );
  NANDN U3850 ( .A(n2391), .B(n2254), .Z(n2255) );
  XOR U3851 ( .A(n2577), .B(n2255), .Z(out[1444]) );
  XOR U3852 ( .A(in[826]), .B(n3897), .Z(n2581) );
  NANDN U3853 ( .A(n2392), .B(n2256), .Z(n2257) );
  XOR U3854 ( .A(n2581), .B(n2257), .Z(out[1445]) );
  XOR U3855 ( .A(in[827]), .B(n3901), .Z(n2585) );
  NANDN U3856 ( .A(n2394), .B(n2258), .Z(n2259) );
  XOR U3857 ( .A(n2585), .B(n2259), .Z(out[1446]) );
  XOR U3858 ( .A(in[828]), .B(n3905), .Z(n2589) );
  NANDN U3859 ( .A(n2395), .B(n2260), .Z(n2261) );
  XOR U3860 ( .A(n2589), .B(n2261), .Z(out[1447]) );
  XOR U3861 ( .A(in[829]), .B(n3909), .Z(n2593) );
  NANDN U3862 ( .A(n2396), .B(n2262), .Z(n2263) );
  XOR U3863 ( .A(n2593), .B(n2263), .Z(out[1448]) );
  XOR U3864 ( .A(in[830]), .B(n3913), .Z(n2597) );
  NANDN U3865 ( .A(n2397), .B(n2264), .Z(n2265) );
  XOR U3866 ( .A(n2597), .B(n2265), .Z(out[1449]) );
  XOR U3867 ( .A(in[681]), .B(n4290), .Z(n2769) );
  XOR U3868 ( .A(in[615]), .B(n4142), .Z(n4476) );
  XNOR U3869 ( .A(in[206]), .B(n3960), .Z(n4473) );
  NANDN U3870 ( .A(n4476), .B(n4473), .Z(n2266) );
  XNOR U3871 ( .A(n2769), .B(n2266), .Z(out[144]) );
  XOR U3872 ( .A(in[831]), .B(n3917), .Z(n2601) );
  NANDN U3873 ( .A(n2398), .B(n2267), .Z(n2268) );
  XOR U3874 ( .A(n2601), .B(n2268), .Z(out[1450]) );
  XOR U3875 ( .A(in[768]), .B(n3921), .Z(n2605) );
  NANDN U3876 ( .A(n2399), .B(n2269), .Z(n2270) );
  XOR U3877 ( .A(n2605), .B(n2270), .Z(out[1451]) );
  XOR U3878 ( .A(in[769]), .B(n3925), .Z(n2611) );
  NANDN U3879 ( .A(n2400), .B(n2271), .Z(n2272) );
  XOR U3880 ( .A(n2611), .B(n2272), .Z(out[1452]) );
  XNOR U3881 ( .A(n3930), .B(in[770]), .Z(n2615) );
  NANDN U3882 ( .A(n2401), .B(n2273), .Z(n2274) );
  XNOR U3883 ( .A(n2615), .B(n2274), .Z(out[1453]) );
  IV U3884 ( .A(n3171), .Z(n3934) );
  XOR U3885 ( .A(n3934), .B(in[771]), .Z(n2619) );
  NANDN U3886 ( .A(n2402), .B(n2275), .Z(n2276) );
  XOR U3887 ( .A(n2619), .B(n2276), .Z(out[1454]) );
  IV U3888 ( .A(n3173), .Z(n3941) );
  XOR U3889 ( .A(n3941), .B(in[772]), .Z(n2623) );
  NANDN U3890 ( .A(n2403), .B(n2277), .Z(n2278) );
  XOR U3891 ( .A(n2623), .B(n2278), .Z(out[1455]) );
  IV U3892 ( .A(n3175), .Z(n3945) );
  XOR U3893 ( .A(n3945), .B(in[773]), .Z(n2627) );
  NANDN U3894 ( .A(n2405), .B(n2279), .Z(n2280) );
  XOR U3895 ( .A(n2627), .B(n2280), .Z(out[1456]) );
  IV U3896 ( .A(n3177), .Z(n3949) );
  XOR U3897 ( .A(n3949), .B(in[774]), .Z(n2631) );
  NANDN U3898 ( .A(n2406), .B(n2281), .Z(n2282) );
  XOR U3899 ( .A(n2631), .B(n2282), .Z(out[1457]) );
  IV U3900 ( .A(n3179), .Z(n3953) );
  XOR U3901 ( .A(n3953), .B(in[775]), .Z(n2635) );
  NANDN U3902 ( .A(n2407), .B(n2283), .Z(n2284) );
  XOR U3903 ( .A(n2635), .B(n2284), .Z(out[1458]) );
  IV U3904 ( .A(n3181), .Z(n3957) );
  XOR U3905 ( .A(n3957), .B(in[776]), .Z(n2639) );
  NAND U3906 ( .A(n2285), .B(n2408), .Z(n2286) );
  XOR U3907 ( .A(n2639), .B(n2286), .Z(out[1459]) );
  XOR U3908 ( .A(in[682]), .B(n4292), .Z(n2770) );
  XOR U3909 ( .A(in[616]), .B(n4146), .Z(n4510) );
  XNOR U3910 ( .A(in[207]), .B(n3964), .Z(n4507) );
  NANDN U3911 ( .A(n4510), .B(n4507), .Z(n2287) );
  XNOR U3912 ( .A(n2770), .B(n2287), .Z(out[145]) );
  IV U3913 ( .A(n3183), .Z(n3961) );
  XOR U3914 ( .A(in[777]), .B(n3961), .Z(n2643) );
  NAND U3915 ( .A(n2288), .B(n2410), .Z(n2289) );
  XOR U3916 ( .A(n2643), .B(n2289), .Z(out[1460]) );
  IV U3917 ( .A(n3185), .Z(n3965) );
  XOR U3918 ( .A(n3965), .B(in[778]), .Z(n2647) );
  NAND U3919 ( .A(n2290), .B(n2412), .Z(n2291) );
  XOR U3920 ( .A(n2647), .B(n2291), .Z(out[1461]) );
  IV U3921 ( .A(n2292), .Z(n3969) );
  XOR U3922 ( .A(n3969), .B(in[779]), .Z(n2653) );
  NANDN U3923 ( .A(n2414), .B(n2293), .Z(n2294) );
  XOR U3924 ( .A(n2653), .B(n2294), .Z(out[1462]) );
  IV U3925 ( .A(n3192), .Z(n3973) );
  XOR U3926 ( .A(in[780]), .B(n3973), .Z(n2657) );
  NANDN U3927 ( .A(n2415), .B(n2295), .Z(n2296) );
  XOR U3928 ( .A(n2657), .B(n2296), .Z(out[1463]) );
  IV U3929 ( .A(n3194), .Z(n3977) );
  XOR U3930 ( .A(in[781]), .B(n3977), .Z(n2661) );
  NANDN U3931 ( .A(n2416), .B(n2297), .Z(n2298) );
  XOR U3932 ( .A(n2661), .B(n2298), .Z(out[1464]) );
  IV U3933 ( .A(n3197), .Z(n3984) );
  XOR U3934 ( .A(in[782]), .B(n3984), .Z(n2665) );
  NAND U3935 ( .A(n2299), .B(n2417), .Z(n2300) );
  XOR U3936 ( .A(n2665), .B(n2300), .Z(out[1465]) );
  IV U3937 ( .A(n3200), .Z(n3988) );
  XOR U3938 ( .A(in[783]), .B(n3988), .Z(n2669) );
  NAND U3939 ( .A(n2301), .B(n2420), .Z(n2302) );
  XOR U3940 ( .A(n2669), .B(n2302), .Z(out[1466]) );
  IV U3941 ( .A(n3203), .Z(n3992) );
  XOR U3942 ( .A(in[784]), .B(n3992), .Z(n2673) );
  NAND U3943 ( .A(n2303), .B(n2422), .Z(n2304) );
  XOR U3944 ( .A(n2673), .B(n2304), .Z(out[1467]) );
  IV U3945 ( .A(n3206), .Z(n3996) );
  XOR U3946 ( .A(in[785]), .B(n3996), .Z(n2677) );
  NAND U3947 ( .A(n2305), .B(n2424), .Z(n2306) );
  XOR U3948 ( .A(n2677), .B(n2306), .Z(out[1468]) );
  IV U3949 ( .A(n3209), .Z(n4000) );
  XOR U3950 ( .A(in[786]), .B(n4000), .Z(n2681) );
  NAND U3951 ( .A(n2307), .B(n2426), .Z(n2308) );
  XOR U3952 ( .A(n2681), .B(n2308), .Z(out[1469]) );
  XOR U3953 ( .A(in[683]), .B(n4294), .Z(n2774) );
  XOR U3954 ( .A(in[617]), .B(n4150), .Z(n4549) );
  XNOR U3955 ( .A(in[208]), .B(n3968), .Z(n4546) );
  NANDN U3956 ( .A(n4549), .B(n4546), .Z(n2309) );
  XNOR U3957 ( .A(n2774), .B(n2309), .Z(out[146]) );
  XOR U3958 ( .A(in[787]), .B(n4004), .Z(n2685) );
  NAND U3959 ( .A(n2310), .B(n2428), .Z(n2311) );
  XOR U3960 ( .A(n2685), .B(n2311), .Z(out[1470]) );
  XOR U3961 ( .A(in[788]), .B(n4008), .Z(n2689) );
  NAND U3962 ( .A(n2312), .B(n2430), .Z(n2313) );
  XOR U3963 ( .A(n2689), .B(n2313), .Z(out[1471]) );
  NANDN U3964 ( .A(n2314), .B(n2432), .Z(n2315) );
  XOR U3965 ( .A(n2433), .B(n2315), .Z(out[1472]) );
  NANDN U3966 ( .A(n2316), .B(n2435), .Z(n2317) );
  XOR U3967 ( .A(n2436), .B(n2317), .Z(out[1473]) );
  NANDN U3968 ( .A(n2318), .B(n2440), .Z(n2319) );
  XOR U3969 ( .A(n2441), .B(n2319), .Z(out[1474]) );
  NANDN U3970 ( .A(n2320), .B(n2444), .Z(n2321) );
  XOR U3971 ( .A(n2445), .B(n2321), .Z(out[1475]) );
  NANDN U3972 ( .A(n2322), .B(n2451), .Z(n2323) );
  XOR U3973 ( .A(n2452), .B(n2323), .Z(out[1476]) );
  NANDN U3974 ( .A(n2324), .B(n2454), .Z(n2325) );
  XOR U3975 ( .A(n2455), .B(n2325), .Z(out[1477]) );
  NANDN U3976 ( .A(n2326), .B(n2456), .Z(n2327) );
  XOR U3977 ( .A(n2457), .B(n2327), .Z(out[1478]) );
  NANDN U3978 ( .A(n2328), .B(n2460), .Z(n2329) );
  XOR U3979 ( .A(n2461), .B(n2329), .Z(out[1479]) );
  XNOR U3980 ( .A(in[684]), .B(n4296), .Z(n2905) );
  XOR U3981 ( .A(in[618]), .B(n4160), .Z(n4578) );
  XNOR U3982 ( .A(in[209]), .B(n3972), .Z(n4575) );
  NANDN U3983 ( .A(n4578), .B(n4575), .Z(n2330) );
  XOR U3984 ( .A(n2905), .B(n2330), .Z(out[147]) );
  NANDN U3985 ( .A(n2331), .B(n2466), .Z(n2332) );
  XOR U3986 ( .A(n2467), .B(n2332), .Z(out[1480]) );
  IV U3987 ( .A(n2333), .Z(n2469) );
  NANDN U3988 ( .A(n2334), .B(n2469), .Z(n2335) );
  XOR U3989 ( .A(n2470), .B(n2335), .Z(out[1481]) );
  IV U3990 ( .A(n2336), .Z(n2472) );
  NANDN U3991 ( .A(n2337), .B(n2472), .Z(n2338) );
  XOR U3992 ( .A(n2473), .B(n2338), .Z(out[1482]) );
  IV U3993 ( .A(n2339), .Z(n2475) );
  NANDN U3994 ( .A(n2340), .B(n2475), .Z(n2341) );
  XOR U3995 ( .A(n2476), .B(n2341), .Z(out[1483]) );
  IV U3996 ( .A(n2342), .Z(n2478) );
  NANDN U3997 ( .A(n2343), .B(n2478), .Z(n2344) );
  XOR U3998 ( .A(n2479), .B(n2344), .Z(out[1484]) );
  IV U3999 ( .A(n2345), .Z(n2481) );
  NANDN U4000 ( .A(n2346), .B(n2481), .Z(n2347) );
  XOR U4001 ( .A(n2482), .B(n2347), .Z(out[1485]) );
  IV U4002 ( .A(n2348), .Z(n2485) );
  NANDN U4003 ( .A(n2349), .B(n2485), .Z(n2350) );
  XNOR U4004 ( .A(n2484), .B(n2350), .Z(out[1486]) );
  IV U4005 ( .A(n2352), .Z(n2489) );
  OR U4006 ( .A(n2497), .B(n2354), .Z(n2355) );
  XOR U4007 ( .A(n2498), .B(n2355), .Z(out[1489]) );
  XNOR U4008 ( .A(in[685]), .B(n4298), .Z(n2908) );
  XOR U4009 ( .A(in[619]), .B(n4164), .Z(n4603) );
  XNOR U4010 ( .A(in[210]), .B(n3976), .Z(n4600) );
  NANDN U4011 ( .A(n4603), .B(n4600), .Z(n2356) );
  XOR U4012 ( .A(n2908), .B(n2356), .Z(out[148]) );
  OR U4013 ( .A(n2501), .B(n2357), .Z(n2358) );
  XOR U4014 ( .A(n2502), .B(n2358), .Z(out[1490]) );
  OR U4015 ( .A(n2505), .B(n2359), .Z(n2360) );
  XOR U4016 ( .A(n2506), .B(n2360), .Z(out[1491]) );
  OR U4017 ( .A(n2509), .B(n2361), .Z(n2362) );
  XOR U4018 ( .A(n2510), .B(n2362), .Z(out[1492]) );
  OR U4019 ( .A(n2513), .B(n2363), .Z(n2364) );
  XOR U4020 ( .A(n2514), .B(n2364), .Z(out[1493]) );
  NANDN U4021 ( .A(n2365), .B(n2517), .Z(n2366) );
  XOR U4022 ( .A(n2518), .B(n2366), .Z(out[1494]) );
  NANDN U4023 ( .A(n2367), .B(n2521), .Z(n2368) );
  XNOR U4024 ( .A(n2522), .B(n2368), .Z(out[1495]) );
  NANDN U4025 ( .A(n2369), .B(n2526), .Z(n2370) );
  XNOR U4026 ( .A(n2527), .B(n2370), .Z(out[1496]) );
  NANDN U4027 ( .A(n2371), .B(n2530), .Z(n2372) );
  XNOR U4028 ( .A(n2531), .B(n2372), .Z(out[1497]) );
  NANDN U4029 ( .A(n2373), .B(n2534), .Z(n2374) );
  XNOR U4030 ( .A(n2535), .B(n2374), .Z(out[1498]) );
  XOR U4031 ( .A(in[686]), .B(n4300), .Z(n2911) );
  XOR U4032 ( .A(in[211]), .B(n3347), .Z(n4628) );
  XNOR U4033 ( .A(in[620]), .B(n4168), .Z(n4630) );
  NANDN U4034 ( .A(n4628), .B(n4630), .Z(n2376) );
  XNOR U4035 ( .A(n2911), .B(n2376), .Z(out[149]) );
  XOR U4036 ( .A(in[1424]), .B(n3203), .Z(n4402) );
  XNOR U4037 ( .A(in[1047]), .B(n4495), .Z(n2889) );
  NANDN U4038 ( .A(n4402), .B(n2889), .Z(n2377) );
  XNOR U4039 ( .A(n4401), .B(n2377), .Z(out[14]) );
  NANDN U4040 ( .A(n2378), .B(n2542), .Z(n2379) );
  XNOR U4041 ( .A(n2543), .B(n2379), .Z(out[1500]) );
  NANDN U4042 ( .A(n2380), .B(n2546), .Z(n2381) );
  XNOR U4043 ( .A(n2547), .B(n2381), .Z(out[1501]) );
  NANDN U4044 ( .A(n2382), .B(n2550), .Z(n2383) );
  XNOR U4045 ( .A(n2551), .B(n2383), .Z(out[1502]) );
  NANDN U4046 ( .A(n2384), .B(n2554), .Z(n2385) );
  XNOR U4047 ( .A(n2555), .B(n2385), .Z(out[1503]) );
  NANDN U4048 ( .A(n2386), .B(n2559), .Z(n2387) );
  XNOR U4049 ( .A(n2560), .B(n2387), .Z(out[1504]) );
  XOR U4050 ( .A(in[687]), .B(n4302), .Z(n2914) );
  XOR U4051 ( .A(in[621]), .B(n4172), .Z(n4662) );
  XOR U4052 ( .A(in[212]), .B(n3987), .Z(n4659) );
  NANDN U4053 ( .A(n4662), .B(n4659), .Z(n2393) );
  XNOR U4054 ( .A(n2914), .B(n2393), .Z(out[150]) );
  XOR U4055 ( .A(in[688]), .B(n4309), .Z(n2917) );
  XOR U4056 ( .A(in[213]), .B(n3991), .Z(n4676) );
  XNOR U4057 ( .A(in[622]), .B(n3896), .Z(n4678) );
  NANDN U4058 ( .A(n4676), .B(n4678), .Z(n2404) );
  XNOR U4059 ( .A(n2917), .B(n2404), .Z(out[151]) );
  NANDN U4060 ( .A(n2408), .B(n2639), .Z(n2409) );
  XOR U4061 ( .A(n2640), .B(n2409), .Z(out[1523]) );
  NANDN U4062 ( .A(n2410), .B(n2643), .Z(n2411) );
  XOR U4063 ( .A(n2644), .B(n2411), .Z(out[1524]) );
  NANDN U4064 ( .A(n2412), .B(n2647), .Z(n2413) );
  XOR U4065 ( .A(n2648), .B(n2413), .Z(out[1525]) );
  NANDN U4066 ( .A(n2417), .B(n2665), .Z(n2418) );
  XOR U4067 ( .A(n2666), .B(n2418), .Z(out[1529]) );
  XOR U4068 ( .A(in[689]), .B(n4312), .Z(n2923) );
  XOR U4069 ( .A(in[214]), .B(n3995), .Z(n4692) );
  XNOR U4070 ( .A(in[623]), .B(n3900), .Z(n4694) );
  NANDN U4071 ( .A(n4692), .B(n4694), .Z(n2419) );
  XNOR U4072 ( .A(n2923), .B(n2419), .Z(out[152]) );
  NANDN U4073 ( .A(n2420), .B(n2669), .Z(n2421) );
  XOR U4074 ( .A(n2670), .B(n2421), .Z(out[1530]) );
  NANDN U4075 ( .A(n2422), .B(n2673), .Z(n2423) );
  XOR U4076 ( .A(n2674), .B(n2423), .Z(out[1531]) );
  NANDN U4077 ( .A(n2424), .B(n2677), .Z(n2425) );
  XOR U4078 ( .A(n2678), .B(n2425), .Z(out[1532]) );
  NANDN U4079 ( .A(n2426), .B(n2681), .Z(n2427) );
  XOR U4080 ( .A(n2682), .B(n2427), .Z(out[1533]) );
  NANDN U4081 ( .A(n2428), .B(n2685), .Z(n2429) );
  XOR U4082 ( .A(n2686), .B(n2429), .Z(out[1534]) );
  NANDN U4083 ( .A(n2430), .B(n2689), .Z(n2431) );
  XOR U4084 ( .A(n2690), .B(n2431), .Z(out[1535]) );
  ANDN U4085 ( .B(n2436), .A(n2435), .Z(n2439) );
  XNOR U4086 ( .A(n2437), .B(round_const[1]), .Z(n2438) );
  XNOR U4087 ( .A(n2439), .B(n2438), .Z(out[1537]) );
  ANDN U4088 ( .B(n2441), .A(n2440), .Z(n2442) );
  XOR U4089 ( .A(n2443), .B(n2442), .Z(out[1538]) );
  ANDN U4090 ( .B(n2445), .A(n2444), .Z(n2448) );
  XOR U4091 ( .A(n2446), .B(round_const_3), .Z(n2447) );
  XNOR U4092 ( .A(n2448), .B(n2447), .Z(out[1539]) );
  XOR U4093 ( .A(in[690]), .B(n4315), .Z(n2926) );
  XOR U4094 ( .A(in[624]), .B(n3904), .Z(n4729) );
  XOR U4095 ( .A(in[215]), .B(n3999), .Z(n4726) );
  NANDN U4096 ( .A(n4729), .B(n4726), .Z(n2449) );
  XNOR U4097 ( .A(n2926), .B(n2449), .Z(out[153]) );
  ANDN U4098 ( .B(n2457), .A(n2456), .Z(n2458) );
  XOR U4099 ( .A(n2459), .B(n2458), .Z(out[1542]) );
  ANDN U4100 ( .B(n2461), .A(n2460), .Z(n2464) );
  XNOR U4101 ( .A(n2462), .B(round_const_7), .Z(n2463) );
  XNOR U4102 ( .A(n2464), .B(n2463), .Z(out[1543]) );
  XOR U4103 ( .A(in[691]), .B(n4318), .Z(n2929) );
  XOR U4104 ( .A(in[625]), .B(n3908), .Z(n4777) );
  XOR U4105 ( .A(in[216]), .B(n4003), .Z(n4774) );
  NANDN U4106 ( .A(n4777), .B(n4774), .Z(n2483) );
  XNOR U4107 ( .A(n2929), .B(n2483), .Z(out[154]) );
  NOR U4108 ( .A(n2485), .B(n2484), .Z(n2486) );
  XOR U4109 ( .A(n2487), .B(n2486), .Z(out[1550]) );
  NOR U4110 ( .A(n2489), .B(n2488), .Z(n2492) );
  XNOR U4111 ( .A(n2490), .B(round_const_15), .Z(n2491) );
  XNOR U4112 ( .A(n2492), .B(n2491), .Z(out[1551]) );
  ANDN U4113 ( .B(n2494), .A(n2493), .Z(n2495) );
  XOR U4114 ( .A(n2496), .B(n2495), .Z(out[1552]) );
  AND U4115 ( .A(n2498), .B(n2497), .Z(n2499) );
  XOR U4116 ( .A(n2500), .B(n2499), .Z(out[1553]) );
  AND U4117 ( .A(n2502), .B(n2501), .Z(n2503) );
  XOR U4118 ( .A(n2504), .B(n2503), .Z(out[1554]) );
  AND U4119 ( .A(n2506), .B(n2505), .Z(n2507) );
  XOR U4120 ( .A(n2508), .B(n2507), .Z(out[1555]) );
  AND U4121 ( .A(n2510), .B(n2509), .Z(n2511) );
  XOR U4122 ( .A(n2512), .B(n2511), .Z(out[1556]) );
  AND U4123 ( .A(n2514), .B(n2513), .Z(n2515) );
  XOR U4124 ( .A(n2516), .B(n2515), .Z(out[1557]) );
  ANDN U4125 ( .B(n2518), .A(n2517), .Z(n2519) );
  XOR U4126 ( .A(n2520), .B(n2519), .Z(out[1558]) );
  NOR U4127 ( .A(n2522), .B(n2521), .Z(n2523) );
  XOR U4128 ( .A(n2524), .B(n2523), .Z(out[1559]) );
  XOR U4129 ( .A(in[692]), .B(n4321), .Z(n2932) );
  XOR U4130 ( .A(in[626]), .B(n3912), .Z(n4821) );
  XOR U4131 ( .A(in[217]), .B(n4007), .Z(n4818) );
  NANDN U4132 ( .A(n4821), .B(n4818), .Z(n2525) );
  XNOR U4133 ( .A(n2932), .B(n2525), .Z(out[155]) );
  NOR U4134 ( .A(n2527), .B(n2526), .Z(n2528) );
  XOR U4135 ( .A(n2529), .B(n2528), .Z(out[1560]) );
  NOR U4136 ( .A(n2531), .B(n2530), .Z(n2532) );
  XOR U4137 ( .A(n2533), .B(n2532), .Z(out[1561]) );
  NOR U4138 ( .A(n2535), .B(n2534), .Z(n2536) );
  XOR U4139 ( .A(n2537), .B(n2536), .Z(out[1562]) );
  NOR U4140 ( .A(n2539), .B(n2538), .Z(n2540) );
  XOR U4141 ( .A(n2541), .B(n2540), .Z(out[1563]) );
  NOR U4142 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U4143 ( .A(n2545), .B(n2544), .Z(out[1564]) );
  NOR U4144 ( .A(n2547), .B(n2546), .Z(n2548) );
  XOR U4145 ( .A(n2549), .B(n2548), .Z(out[1565]) );
  NOR U4146 ( .A(n2551), .B(n2550), .Z(n2552) );
  XOR U4147 ( .A(n2553), .B(n2552), .Z(out[1566]) );
  NOR U4148 ( .A(n2555), .B(n2554), .Z(n2558) );
  XNOR U4149 ( .A(n2556), .B(round_const_31), .Z(n2557) );
  XNOR U4150 ( .A(n2558), .B(n2557), .Z(out[1567]) );
  NOR U4151 ( .A(n2560), .B(n2559), .Z(n2561) );
  XOR U4152 ( .A(n2562), .B(n2561), .Z(out[1568]) );
  NOR U4153 ( .A(n2564), .B(n2563), .Z(n2565) );
  XOR U4154 ( .A(n2566), .B(n2565), .Z(out[1569]) );
  XOR U4155 ( .A(in[693]), .B(n4324), .Z(n2934) );
  XOR U4156 ( .A(in[218]), .B(n4011), .Z(n4863) );
  XNOR U4157 ( .A(in[627]), .B(n2567), .Z(n4865) );
  NANDN U4158 ( .A(n4863), .B(n4865), .Z(n2568) );
  XNOR U4159 ( .A(n2934), .B(n2568), .Z(out[156]) );
  NOR U4160 ( .A(n2570), .B(n2569), .Z(n2571) );
  XOR U4161 ( .A(n2572), .B(n2571), .Z(out[1570]) );
  NOR U4162 ( .A(n2574), .B(n2573), .Z(n2575) );
  XOR U4163 ( .A(n2576), .B(n2575), .Z(out[1571]) );
  NOR U4164 ( .A(n2578), .B(n2577), .Z(n2579) );
  XOR U4165 ( .A(n2580), .B(n2579), .Z(out[1572]) );
  NOR U4166 ( .A(n2582), .B(n2581), .Z(n2583) );
  XOR U4167 ( .A(n2584), .B(n2583), .Z(out[1573]) );
  NOR U4168 ( .A(n2586), .B(n2585), .Z(n2587) );
  XNOR U4169 ( .A(n2588), .B(n2587), .Z(out[1574]) );
  ANDN U4170 ( .B(n2590), .A(n2589), .Z(n2591) );
  XOR U4171 ( .A(n2592), .B(n2591), .Z(out[1575]) );
  ANDN U4172 ( .B(n2594), .A(n2593), .Z(n2595) );
  XOR U4173 ( .A(n2596), .B(n2595), .Z(out[1576]) );
  ANDN U4174 ( .B(n2598), .A(n2597), .Z(n2599) );
  XOR U4175 ( .A(n2600), .B(n2599), .Z(out[1577]) );
  NOR U4176 ( .A(n2602), .B(n2601), .Z(n2603) );
  XOR U4177 ( .A(n2604), .B(n2603), .Z(out[1578]) );
  ANDN U4178 ( .B(n2606), .A(n2605), .Z(n2607) );
  XOR U4179 ( .A(n2608), .B(n2607), .Z(out[1579]) );
  XOR U4180 ( .A(in[694]), .B(n4327), .Z(n2936) );
  XOR U4181 ( .A(in[219]), .B(n4015), .Z(n4907) );
  XNOR U4182 ( .A(in[628]), .B(n2609), .Z(n4909) );
  NANDN U4183 ( .A(n4907), .B(n4909), .Z(n2610) );
  XNOR U4184 ( .A(n2936), .B(n2610), .Z(out[157]) );
  ANDN U4185 ( .B(n2612), .A(n2611), .Z(n2613) );
  XOR U4186 ( .A(n2614), .B(n2613), .Z(out[1580]) );
  AND U4187 ( .A(n2616), .B(n2615), .Z(n2617) );
  XOR U4188 ( .A(n2618), .B(n2617), .Z(out[1581]) );
  ANDN U4189 ( .B(n2620), .A(n2619), .Z(n2621) );
  XOR U4190 ( .A(n2622), .B(n2621), .Z(out[1582]) );
  ANDN U4191 ( .B(n2624), .A(n2623), .Z(n2625) );
  XOR U4192 ( .A(n2626), .B(n2625), .Z(out[1583]) );
  ANDN U4193 ( .B(n2628), .A(n2627), .Z(n2629) );
  XOR U4194 ( .A(n2630), .B(n2629), .Z(out[1584]) );
  ANDN U4195 ( .B(n2632), .A(n2631), .Z(n2633) );
  XOR U4196 ( .A(n2634), .B(n2633), .Z(out[1585]) );
  ANDN U4197 ( .B(n2636), .A(n2635), .Z(n2637) );
  XOR U4198 ( .A(n2638), .B(n2637), .Z(out[1586]) );
  ANDN U4199 ( .B(n2640), .A(n2639), .Z(n2641) );
  XOR U4200 ( .A(n2642), .B(n2641), .Z(out[1587]) );
  ANDN U4201 ( .B(n2644), .A(n2643), .Z(n2645) );
  XOR U4202 ( .A(n2646), .B(n2645), .Z(out[1588]) );
  ANDN U4203 ( .B(n2648), .A(n2647), .Z(n2649) );
  XOR U4204 ( .A(n2650), .B(n2649), .Z(out[1589]) );
  XOR U4205 ( .A(in[695]), .B(n4330), .Z(n2938) );
  XNOR U4206 ( .A(in[220]), .B(n4019), .Z(n4951) );
  XNOR U4207 ( .A(in[629]), .B(n2651), .Z(n4953) );
  NANDN U4208 ( .A(n4951), .B(n4953), .Z(n2652) );
  XNOR U4209 ( .A(n2938), .B(n2652), .Z(out[158]) );
  ANDN U4210 ( .B(n2654), .A(n2653), .Z(n2655) );
  XNOR U4211 ( .A(n2656), .B(n2655), .Z(out[1590]) );
  ANDN U4212 ( .B(n2658), .A(n2657), .Z(n2659) );
  XNOR U4213 ( .A(n2660), .B(n2659), .Z(out[1591]) );
  ANDN U4214 ( .B(n2662), .A(n2661), .Z(n2663) );
  XNOR U4215 ( .A(n2664), .B(n2663), .Z(out[1592]) );
  ANDN U4216 ( .B(n2666), .A(n2665), .Z(n2667) );
  XOR U4217 ( .A(n2668), .B(n2667), .Z(out[1593]) );
  ANDN U4218 ( .B(n2670), .A(n2669), .Z(n2671) );
  XOR U4219 ( .A(n2672), .B(n2671), .Z(out[1594]) );
  ANDN U4220 ( .B(n2674), .A(n2673), .Z(n2675) );
  XOR U4221 ( .A(n2676), .B(n2675), .Z(out[1595]) );
  ANDN U4222 ( .B(n2678), .A(n2677), .Z(n2679) );
  XOR U4223 ( .A(n2680), .B(n2679), .Z(out[1596]) );
  ANDN U4224 ( .B(n2682), .A(n2681), .Z(n2683) );
  XOR U4225 ( .A(n2684), .B(n2683), .Z(out[1597]) );
  ANDN U4226 ( .B(n2686), .A(n2685), .Z(n2687) );
  XOR U4227 ( .A(n2688), .B(n2687), .Z(out[1598]) );
  ANDN U4228 ( .B(n2690), .A(n2689), .Z(n2693) );
  XNOR U4229 ( .A(n2691), .B(round_const_63), .Z(n2692) );
  XNOR U4230 ( .A(n2693), .B(n2692), .Z(out[1599]) );
  XOR U4231 ( .A(in[696]), .B(n4176), .Z(n2940) );
  XNOR U4232 ( .A(in[221]), .B(n4027), .Z(n4995) );
  XNOR U4233 ( .A(in[630]), .B(n3063), .Z(n4997) );
  NANDN U4234 ( .A(n4995), .B(n4997), .Z(n2694) );
  XNOR U4235 ( .A(n2940), .B(n2694), .Z(out[159]) );
  XOR U4236 ( .A(in[1425]), .B(n3206), .Z(n4436) );
  XNOR U4237 ( .A(in[1048]), .B(n4498), .Z(n2892) );
  NANDN U4238 ( .A(n4436), .B(n2892), .Z(n2695) );
  XNOR U4239 ( .A(n4435), .B(n2695), .Z(out[15]) );
  XOR U4240 ( .A(in[697]), .B(n4179), .Z(n2942) );
  XNOR U4241 ( .A(in[222]), .B(n4031), .Z(n5039) );
  XNOR U4242 ( .A(in[631]), .B(n3065), .Z(n5041) );
  NANDN U4243 ( .A(n5039), .B(n5041), .Z(n2696) );
  XNOR U4244 ( .A(n2942), .B(n2696), .Z(out[160]) );
  XOR U4245 ( .A(in[698]), .B(n4182), .Z(n2944) );
  XNOR U4246 ( .A(in[223]), .B(n4035), .Z(n5080) );
  XNOR U4247 ( .A(in[632]), .B(n3068), .Z(n5082) );
  NANDN U4248 ( .A(n5080), .B(n5082), .Z(n2697) );
  XNOR U4249 ( .A(n2944), .B(n2697), .Z(out[161]) );
  XOR U4250 ( .A(in[699]), .B(n4185), .Z(n2948) );
  XNOR U4251 ( .A(in[633]), .B(n2698), .Z(n5117) );
  XOR U4252 ( .A(in[224]), .B(n4039), .Z(n5114) );
  NAND U4253 ( .A(n5117), .B(n5114), .Z(n2699) );
  XNOR U4254 ( .A(n2948), .B(n2699), .Z(out[162]) );
  XOR U4255 ( .A(in[700]), .B(n4188), .Z(n2950) );
  XNOR U4256 ( .A(in[634]), .B(n2700), .Z(n5160) );
  XOR U4257 ( .A(in[225]), .B(n4043), .Z(n5157) );
  NAND U4258 ( .A(n5160), .B(n5157), .Z(n2701) );
  XOR U4259 ( .A(n2950), .B(n2701), .Z(out[163]) );
  XOR U4260 ( .A(in[701]), .B(n4191), .Z(n2952) );
  ANDN U4261 ( .B(n3113), .A(n2702), .Z(n2703) );
  XNOR U4262 ( .A(n2952), .B(n2703), .Z(out[164]) );
  XOR U4263 ( .A(in[702]), .B(n4196), .Z(n2954) );
  ANDN U4264 ( .B(n3135), .A(n2704), .Z(n2705) );
  XNOR U4265 ( .A(n2954), .B(n2705), .Z(out[165]) );
  XNOR U4266 ( .A(in[703]), .B(n4197), .Z(n2956) );
  ANDN U4267 ( .B(n3154), .A(n2706), .Z(n2707) );
  XNOR U4268 ( .A(n2956), .B(n2707), .Z(out[166]) );
  XOR U4269 ( .A(in[640]), .B(n4198), .Z(n2958) );
  ANDN U4270 ( .B(n3165), .A(n2708), .Z(n2709) );
  XNOR U4271 ( .A(n2958), .B(n2709), .Z(out[167]) );
  XOR U4272 ( .A(in[641]), .B(n4199), .Z(n2960) );
  NOR U4273 ( .A(n2710), .B(n3190), .Z(n2711) );
  XNOR U4274 ( .A(n2960), .B(n2711), .Z(out[168]) );
  XOR U4275 ( .A(in[642]), .B(n4200), .Z(n2962) );
  NOR U4276 ( .A(n2712), .B(n3221), .Z(n2713) );
  XNOR U4277 ( .A(n2962), .B(n2713), .Z(out[169]) );
  XOR U4278 ( .A(in[1426]), .B(n3209), .Z(n4474) );
  XNOR U4279 ( .A(in[1049]), .B(n4501), .Z(n2895) );
  NANDN U4280 ( .A(n4474), .B(n2895), .Z(n2714) );
  XNOR U4281 ( .A(n4473), .B(n2714), .Z(out[16]) );
  XOR U4282 ( .A(in[643]), .B(n4201), .Z(n2964) );
  NOR U4283 ( .A(n2715), .B(n3245), .Z(n2716) );
  XNOR U4284 ( .A(n2964), .B(n2716), .Z(out[170]) );
  XOR U4285 ( .A(in[644]), .B(n4202), .Z(n2966) );
  NOR U4286 ( .A(n2717), .B(n3257), .Z(n2718) );
  XNOR U4287 ( .A(n2966), .B(n2718), .Z(out[171]) );
  XOR U4288 ( .A(in[645]), .B(n4203), .Z(n2972) );
  NOR U4289 ( .A(n2719), .B(n3267), .Z(n2720) );
  XNOR U4290 ( .A(n2972), .B(n2720), .Z(out[172]) );
  XOR U4291 ( .A(in[646]), .B(n4206), .Z(n2974) );
  NOR U4292 ( .A(n3301), .B(n2809), .Z(n2721) );
  XNOR U4293 ( .A(n2974), .B(n2721), .Z(out[173]) );
  XOR U4294 ( .A(in[647]), .B(n4209), .Z(n2976) );
  NOR U4295 ( .A(n3331), .B(n2811), .Z(n2722) );
  XNOR U4296 ( .A(n2976), .B(n2722), .Z(out[174]) );
  XNOR U4297 ( .A(in[648]), .B(n4214), .Z(n2978) );
  NOR U4298 ( .A(n3360), .B(n2813), .Z(n2723) );
  XNOR U4299 ( .A(n2978), .B(n2723), .Z(out[175]) );
  XOR U4300 ( .A(in[649]), .B(n4217), .Z(n2980) );
  NOR U4301 ( .A(n3388), .B(n2818), .Z(n2724) );
  XNOR U4302 ( .A(n2980), .B(n2724), .Z(out[176]) );
  XOR U4303 ( .A(in[650]), .B(n3088), .Z(n2982) );
  NOR U4304 ( .A(n3423), .B(n2820), .Z(n2725) );
  XOR U4305 ( .A(n2982), .B(n2725), .Z(out[177]) );
  IV U4306 ( .A(n3090), .Z(n4223) );
  XOR U4307 ( .A(in[651]), .B(n4223), .Z(n2983) );
  NOR U4308 ( .A(n3458), .B(n2822), .Z(n2726) );
  XNOR U4309 ( .A(n2983), .B(n2726), .Z(out[178]) );
  IV U4310 ( .A(n3092), .Z(n4226) );
  XOR U4311 ( .A(in[652]), .B(n4226), .Z(n2985) );
  NOR U4312 ( .A(n3480), .B(n2824), .Z(n2727) );
  XNOR U4313 ( .A(n2985), .B(n2727), .Z(out[179]) );
  XOR U4314 ( .A(in[1427]), .B(n3212), .Z(n4508) );
  XNOR U4315 ( .A(in[1050]), .B(n4504), .Z(n2898) );
  NANDN U4316 ( .A(n4508), .B(n2898), .Z(n2728) );
  XNOR U4317 ( .A(n4507), .B(n2728), .Z(out[17]) );
  IV U4318 ( .A(n3096), .Z(n4229) );
  XOR U4319 ( .A(in[653]), .B(n4229), .Z(n2987) );
  NOR U4320 ( .A(n3502), .B(n2826), .Z(n2729) );
  XNOR U4321 ( .A(n2987), .B(n2729), .Z(out[180]) );
  XNOR U4322 ( .A(in[654]), .B(n4232), .Z(n2990) );
  NOR U4323 ( .A(n3517), .B(n2828), .Z(n2730) );
  XNOR U4324 ( .A(n2990), .B(n2730), .Z(out[181]) );
  XNOR U4325 ( .A(in[655]), .B(n4235), .Z(n2995) );
  NOR U4326 ( .A(n3545), .B(n2830), .Z(n2731) );
  XNOR U4327 ( .A(n2995), .B(n2731), .Z(out[182]) );
  XNOR U4328 ( .A(in[656]), .B(n4238), .Z(n2998) );
  NOR U4329 ( .A(n3575), .B(n2832), .Z(n2732) );
  XNOR U4330 ( .A(n2998), .B(n2732), .Z(out[183]) );
  XNOR U4331 ( .A(in[657]), .B(n4239), .Z(n3001) );
  NOR U4332 ( .A(n3599), .B(n2834), .Z(n2733) );
  XNOR U4333 ( .A(n3001), .B(n2733), .Z(out[184]) );
  IV U4334 ( .A(n3102), .Z(n4242) );
  XOR U4335 ( .A(in[658]), .B(n4242), .Z(n3003) );
  NOR U4336 ( .A(n3629), .B(n2836), .Z(n2734) );
  XNOR U4337 ( .A(n3003), .B(n2734), .Z(out[185]) );
  IV U4338 ( .A(n3104), .Z(n4243) );
  XOR U4339 ( .A(in[659]), .B(n4243), .Z(n3005) );
  NOR U4340 ( .A(n3673), .B(n2841), .Z(n2735) );
  XNOR U4341 ( .A(n3005), .B(n2735), .Z(out[186]) );
  XOR U4342 ( .A(in[660]), .B(n4246), .Z(n3007) );
  NOR U4343 ( .A(n3717), .B(n2843), .Z(n2736) );
  XOR U4344 ( .A(n3007), .B(n2736), .Z(out[187]) );
  XOR U4345 ( .A(in[661]), .B(n4249), .Z(n3010) );
  NOR U4346 ( .A(n3763), .B(n2845), .Z(n2737) );
  XOR U4347 ( .A(n3010), .B(n2737), .Z(out[188]) );
  XOR U4348 ( .A(in[662]), .B(n4250), .Z(n3013) );
  XOR U4349 ( .A(in[1428]), .B(n3215), .Z(n4547) );
  XNOR U4350 ( .A(in[1051]), .B(n2738), .Z(n2901) );
  NANDN U4351 ( .A(n4547), .B(n2901), .Z(n2739) );
  XNOR U4352 ( .A(n4546), .B(n2739), .Z(out[18]) );
  XOR U4353 ( .A(in[663]), .B(n4251), .Z(n3014) );
  XOR U4354 ( .A(in[664]), .B(n4252), .Z(n3017) );
  NANDN U4355 ( .A(n2853), .B(n3938), .Z(n2740) );
  XOR U4356 ( .A(n2854), .B(n2740), .Z(out[192]) );
  XNOR U4357 ( .A(in[1034]), .B(n4452), .Z(n2757) );
  ANDN U4358 ( .B(n3981), .A(n2856), .Z(n2741) );
  XNOR U4359 ( .A(n2757), .B(n2741), .Z(out[193]) );
  XNOR U4360 ( .A(in[1035]), .B(n4455), .Z(n2970) );
  ANDN U4361 ( .B(n4025), .A(n2742), .Z(n2743) );
  XNOR U4362 ( .A(n2970), .B(n2743), .Z(out[194]) );
  XOR U4363 ( .A(n4458), .B(in[1036]), .Z(n3166) );
  ANDN U4364 ( .B(n4069), .A(n2744), .Z(n2745) );
  XNOR U4365 ( .A(n3166), .B(n2745), .Z(out[195]) );
  XOR U4366 ( .A(n4461), .B(in[1037]), .Z(n3424) );
  ANDN U4367 ( .B(n4113), .A(n2746), .Z(n2747) );
  XNOR U4368 ( .A(n3424), .B(n2747), .Z(out[196]) );
  XOR U4369 ( .A(n4464), .B(in[1038]), .Z(n3718) );
  ANDN U4370 ( .B(n4157), .A(n2748), .Z(n2749) );
  XNOR U4371 ( .A(n3718), .B(n2749), .Z(out[197]) );
  XOR U4372 ( .A(n4467), .B(in[1039]), .Z(n4158) );
  ANDN U4373 ( .B(n4195), .A(n2750), .Z(n2751) );
  XNOR U4374 ( .A(n4158), .B(n2751), .Z(out[198]) );
  XOR U4375 ( .A(n4470), .B(in[1040]), .Z(n4439) );
  ANDN U4376 ( .B(n4213), .A(n2752), .Z(n2753) );
  XNOR U4377 ( .A(n4439), .B(n2753), .Z(out[199]) );
  XOR U4378 ( .A(in[1429]), .B(n2754), .Z(n4576) );
  XNOR U4379 ( .A(in[1052]), .B(n2755), .Z(n2904) );
  NANDN U4380 ( .A(n4576), .B(n2904), .Z(n2756) );
  XNOR U4381 ( .A(n4575), .B(n2756), .Z(out[19]) );
  XOR U4382 ( .A(n3171), .B(in[1411]), .Z(n3979) );
  IV U4383 ( .A(n2757), .Z(n2855) );
  NANDN U4384 ( .A(n3979), .B(n2855), .Z(n2758) );
  XNOR U4385 ( .A(n3980), .B(n2758), .Z(out[1]) );
  XOR U4386 ( .A(n4477), .B(in[1041]), .Z(n4730) );
  ANDN U4387 ( .B(n4241), .A(n2759), .Z(n2760) );
  XNOR U4388 ( .A(n4730), .B(n2760), .Z(out[200]) );
  XOR U4389 ( .A(n4480), .B(in[1042]), .Z(n5161) );
  ANDN U4390 ( .B(n4257), .A(n2761), .Z(n2762) );
  XNOR U4391 ( .A(n5161), .B(n2762), .Z(out[201]) );
  NAND U4392 ( .A(n4283), .B(n2878), .Z(n2763) );
  XNOR U4393 ( .A(n2877), .B(n2763), .Z(out[202]) );
  NANDN U4394 ( .A(n2880), .B(n4308), .Z(n2764) );
  XNOR U4395 ( .A(n2881), .B(n2764), .Z(out[203]) );
  NANDN U4396 ( .A(n2882), .B(n4340), .Z(n2765) );
  XNOR U4397 ( .A(n2883), .B(n2765), .Z(out[204]) );
  NANDN U4398 ( .A(n2884), .B(n4371), .Z(n2766) );
  XNOR U4399 ( .A(n2885), .B(n2766), .Z(out[205]) );
  IV U4400 ( .A(n2767), .Z(n2890) );
  IV U4401 ( .A(n2768), .Z(n2893) );
  IV U4402 ( .A(n2769), .Z(n2896) );
  IV U4403 ( .A(n2770), .Z(n2899) );
  XOR U4404 ( .A(in[1430]), .B(n2771), .Z(n4601) );
  XNOR U4405 ( .A(in[1053]), .B(n2772), .Z(n2907) );
  NANDN U4406 ( .A(n4601), .B(n2907), .Z(n2773) );
  XNOR U4407 ( .A(n4600), .B(n2773), .Z(out[20]) );
  IV U4408 ( .A(n2774), .Z(n2902) );
  XOR U4409 ( .A(in[1054]), .B(n4520), .Z(n2779) );
  IV U4410 ( .A(n2779), .Z(n2910) );
  NOR U4411 ( .A(n4630), .B(n2911), .Z(n2775) );
  XOR U4412 ( .A(n2910), .B(n2775), .Z(out[213]) );
  XOR U4413 ( .A(in[1055]), .B(n4524), .Z(n2793) );
  IV U4414 ( .A(n2793), .Z(n2913) );
  XOR U4415 ( .A(in[1056]), .B(n4528), .Z(n2816) );
  IV U4416 ( .A(n2816), .Z(n2916) );
  NOR U4417 ( .A(n4678), .B(n2917), .Z(n2776) );
  XOR U4418 ( .A(n2916), .B(n2776), .Z(out[215]) );
  XOR U4419 ( .A(in[1057]), .B(n4532), .Z(n2839) );
  IV U4420 ( .A(n2839), .Z(n2922) );
  NOR U4421 ( .A(n4694), .B(n2923), .Z(n2777) );
  XOR U4422 ( .A(n2922), .B(n2777), .Z(out[216]) );
  XOR U4423 ( .A(in[1058]), .B(n4536), .Z(n2863) );
  IV U4424 ( .A(n2863), .Z(n2925) );
  XOR U4425 ( .A(in[1059]), .B(n4540), .Z(n2887) );
  IV U4426 ( .A(n2887), .Z(n2928) );
  XNOR U4427 ( .A(in[1060]), .B(n4544), .Z(n2920) );
  IV U4428 ( .A(n2920), .Z(n2931) );
  XOR U4429 ( .A(in[1431]), .B(n2778), .Z(n4629) );
  OR U4430 ( .A(n4629), .B(n2779), .Z(n2780) );
  XOR U4431 ( .A(n4628), .B(n2780), .Z(out[21]) );
  XNOR U4432 ( .A(in[1061]), .B(n4550), .Z(n2946) );
  NOR U4433 ( .A(n4865), .B(n2934), .Z(n2781) );
  XNOR U4434 ( .A(n2946), .B(n2781), .Z(out[220]) );
  XNOR U4435 ( .A(in[1062]), .B(n4552), .Z(n2968) );
  NOR U4436 ( .A(n4909), .B(n2936), .Z(n2782) );
  XNOR U4437 ( .A(n2968), .B(n2782), .Z(out[221]) );
  XNOR U4438 ( .A(in[1063]), .B(n4333), .Z(n2992) );
  NOR U4439 ( .A(n4953), .B(n2938), .Z(n2783) );
  XNOR U4440 ( .A(n2992), .B(n2783), .Z(out[222]) );
  XNOR U4441 ( .A(in[1064]), .B(n4335), .Z(n3020) );
  NOR U4442 ( .A(n4997), .B(n2940), .Z(n2784) );
  XNOR U4443 ( .A(n3020), .B(n2784), .Z(out[223]) );
  XNOR U4444 ( .A(in[1065]), .B(n4341), .Z(n3040) );
  NOR U4445 ( .A(n5041), .B(n2942), .Z(n2785) );
  XNOR U4446 ( .A(n3040), .B(n2785), .Z(out[224]) );
  XNOR U4447 ( .A(in[1066]), .B(n4343), .Z(n3052) );
  NOR U4448 ( .A(n5082), .B(n2944), .Z(n2786) );
  XNOR U4449 ( .A(n3052), .B(n2786), .Z(out[225]) );
  XNOR U4450 ( .A(in[1067]), .B(n4345), .Z(n3073) );
  NOR U4451 ( .A(n5117), .B(n2948), .Z(n2787) );
  XNOR U4452 ( .A(n3073), .B(n2787), .Z(out[226]) );
  XNOR U4453 ( .A(in[1068]), .B(n4348), .Z(n3094) );
  XOR U4454 ( .A(in[1069]), .B(n4351), .Z(n3111) );
  NANDN U4455 ( .A(n2788), .B(n2952), .Z(n2789) );
  XNOR U4456 ( .A(n3111), .B(n2789), .Z(out[228]) );
  XOR U4457 ( .A(in[1070]), .B(n4354), .Z(n3133) );
  NANDN U4458 ( .A(n2790), .B(n2954), .Z(n2791) );
  XNOR U4459 ( .A(n3133), .B(n2791), .Z(out[229]) );
  XOR U4460 ( .A(in[1432]), .B(n2792), .Z(n4660) );
  OR U4461 ( .A(n4660), .B(n2793), .Z(n2794) );
  XNOR U4462 ( .A(n4659), .B(n2794), .Z(out[22]) );
  XNOR U4463 ( .A(in[1071]), .B(n4356), .Z(n3151) );
  NANDN U4464 ( .A(n2795), .B(n2956), .Z(n2796) );
  XOR U4465 ( .A(n3151), .B(n2796), .Z(out[230]) );
  XOR U4466 ( .A(in[1072]), .B(n4359), .Z(n3163) );
  NANDN U4467 ( .A(n2797), .B(n2958), .Z(n2798) );
  XNOR U4468 ( .A(n3163), .B(n2798), .Z(out[231]) );
  XOR U4469 ( .A(in[1073]), .B(n4362), .Z(n3188) );
  NANDN U4470 ( .A(n2799), .B(n2960), .Z(n2800) );
  XNOR U4471 ( .A(n3188), .B(n2800), .Z(out[232]) );
  XOR U4472 ( .A(in[1074]), .B(n4365), .Z(n3218) );
  NANDN U4473 ( .A(n2801), .B(n2962), .Z(n2802) );
  XNOR U4474 ( .A(n3218), .B(n2802), .Z(out[233]) );
  XOR U4475 ( .A(in[1075]), .B(n4372), .Z(n3242) );
  NANDN U4476 ( .A(n2803), .B(n2964), .Z(n2804) );
  XNOR U4477 ( .A(n3242), .B(n2804), .Z(out[234]) );
  XOR U4478 ( .A(in[1076]), .B(n4375), .Z(n3254) );
  NANDN U4479 ( .A(n2805), .B(n2966), .Z(n2806) );
  XNOR U4480 ( .A(n3254), .B(n2806), .Z(out[235]) );
  XOR U4481 ( .A(in[1077]), .B(n4378), .Z(n3264) );
  NANDN U4482 ( .A(n2807), .B(n2972), .Z(n2808) );
  XNOR U4483 ( .A(n3264), .B(n2808), .Z(out[236]) );
  XOR U4484 ( .A(in[1078]), .B(n4381), .Z(n3298) );
  NAND U4485 ( .A(n2809), .B(n2974), .Z(n2810) );
  XNOR U4486 ( .A(n3298), .B(n2810), .Z(out[237]) );
  XOR U4487 ( .A(in[1079]), .B(n4384), .Z(n3328) );
  NAND U4488 ( .A(n2811), .B(n2976), .Z(n2812) );
  XNOR U4489 ( .A(n3328), .B(n2812), .Z(out[238]) );
  XNOR U4490 ( .A(in[1080]), .B(n4386), .Z(n3357) );
  NAND U4491 ( .A(n2813), .B(n2978), .Z(n2814) );
  XOR U4492 ( .A(n3357), .B(n2814), .Z(out[239]) );
  XOR U4493 ( .A(in[1433]), .B(n2815), .Z(n4677) );
  OR U4494 ( .A(n4677), .B(n2816), .Z(n2817) );
  XOR U4495 ( .A(n4676), .B(n2817), .Z(out[23]) );
  XOR U4496 ( .A(in[1081]), .B(n4389), .Z(n3385) );
  NAND U4497 ( .A(n2818), .B(n2980), .Z(n2819) );
  XNOR U4498 ( .A(n3385), .B(n2819), .Z(out[240]) );
  XOR U4499 ( .A(in[1082]), .B(n4392), .Z(n3420) );
  NANDN U4500 ( .A(n2982), .B(n2820), .Z(n2821) );
  XOR U4501 ( .A(n3420), .B(n2821), .Z(out[241]) );
  XOR U4502 ( .A(in[1083]), .B(n4395), .Z(n3455) );
  NAND U4503 ( .A(n2822), .B(n2983), .Z(n2823) );
  XOR U4504 ( .A(n3455), .B(n2823), .Z(out[242]) );
  XNOR U4505 ( .A(in[1084]), .B(n4398), .Z(n3477) );
  NAND U4506 ( .A(n2824), .B(n2985), .Z(n2825) );
  XOR U4507 ( .A(n3477), .B(n2825), .Z(out[243]) );
  XNOR U4508 ( .A(in[1085]), .B(n4405), .Z(n3499) );
  NAND U4509 ( .A(n2826), .B(n2987), .Z(n2827) );
  XOR U4510 ( .A(n3499), .B(n2827), .Z(out[244]) );
  XOR U4511 ( .A(in[1086]), .B(n4408), .Z(n2989) );
  NAND U4512 ( .A(n2828), .B(n2990), .Z(n2829) );
  XNOR U4513 ( .A(n2989), .B(n2829), .Z(out[245]) );
  XOR U4514 ( .A(in[1087]), .B(n4411), .Z(n2994) );
  NAND U4515 ( .A(n2830), .B(n2995), .Z(n2831) );
  XNOR U4516 ( .A(n2994), .B(n2831), .Z(out[246]) );
  XOR U4517 ( .A(in[1024]), .B(n4414), .Z(n2997) );
  NAND U4518 ( .A(n2832), .B(n2998), .Z(n2833) );
  XNOR U4519 ( .A(n2997), .B(n2833), .Z(out[247]) );
  XOR U4520 ( .A(in[1025]), .B(n4417), .Z(n3000) );
  NAND U4521 ( .A(n2834), .B(n3001), .Z(n2835) );
  XNOR U4522 ( .A(n3000), .B(n2835), .Z(out[248]) );
  XNOR U4523 ( .A(in[1026]), .B(n4420), .Z(n3626) );
  NAND U4524 ( .A(n2836), .B(n3003), .Z(n2837) );
  XOR U4525 ( .A(n3626), .B(n2837), .Z(out[249]) );
  XOR U4526 ( .A(in[1434]), .B(n2838), .Z(n4693) );
  OR U4527 ( .A(n4693), .B(n2839), .Z(n2840) );
  XOR U4528 ( .A(n4692), .B(n2840), .Z(out[24]) );
  XNOR U4529 ( .A(in[1027]), .B(n4423), .Z(n3670) );
  NAND U4530 ( .A(n2841), .B(n3005), .Z(n2842) );
  XOR U4531 ( .A(n3670), .B(n2842), .Z(out[250]) );
  XOR U4532 ( .A(in[1028]), .B(n4426), .Z(n3008) );
  IV U4533 ( .A(n3008), .Z(n3714) );
  NANDN U4534 ( .A(n3007), .B(n2843), .Z(n2844) );
  XOR U4535 ( .A(n3714), .B(n2844), .Z(out[251]) );
  XOR U4536 ( .A(in[1029]), .B(n4429), .Z(n3011) );
  IV U4537 ( .A(n3011), .Z(n3760) );
  NANDN U4538 ( .A(n3010), .B(n2845), .Z(n2846) );
  XOR U4539 ( .A(n3760), .B(n2846), .Z(out[252]) );
  XOR U4540 ( .A(in[1030]), .B(n4432), .Z(n3804) );
  NANDN U4541 ( .A(n3013), .B(n2847), .Z(n2848) );
  XOR U4542 ( .A(n3804), .B(n2848), .Z(out[253]) );
  XOR U4543 ( .A(in[1031]), .B(n4443), .Z(n3015) );
  IV U4544 ( .A(n3015), .Z(n3848) );
  NANDN U4545 ( .A(n3014), .B(n2849), .Z(n2850) );
  XOR U4546 ( .A(n3848), .B(n2850), .Z(out[254]) );
  XOR U4547 ( .A(in[1032]), .B(n4446), .Z(n3018) );
  IV U4548 ( .A(n3018), .Z(n3892) );
  NANDN U4549 ( .A(n3017), .B(n2851), .Z(n2852) );
  XOR U4550 ( .A(n3892), .B(n2852), .Z(out[255]) );
  ANDN U4551 ( .B(n2856), .A(n2855), .Z(n2857) );
  XOR U4552 ( .A(n3979), .B(n2857), .Z(out[257]) );
  XNOR U4553 ( .A(n3941), .B(in[1412]), .Z(n4023) );
  NANDN U4554 ( .A(n2858), .B(n2970), .Z(n2859) );
  XNOR U4555 ( .A(n4023), .B(n2859), .Z(out[258]) );
  XNOR U4556 ( .A(n3945), .B(in[1413]), .Z(n4067) );
  NANDN U4557 ( .A(n2860), .B(n3166), .Z(n2861) );
  XNOR U4558 ( .A(n4067), .B(n2861), .Z(out[259]) );
  XOR U4559 ( .A(in[1435]), .B(n2862), .Z(n4727) );
  OR U4560 ( .A(n4727), .B(n2863), .Z(n2864) );
  XNOR U4561 ( .A(n4726), .B(n2864), .Z(out[25]) );
  XNOR U4562 ( .A(n3949), .B(in[1414]), .Z(n4111) );
  NANDN U4563 ( .A(n2865), .B(n3424), .Z(n2866) );
  XNOR U4564 ( .A(n4111), .B(n2866), .Z(out[260]) );
  XNOR U4565 ( .A(n3953), .B(in[1415]), .Z(n4155) );
  NANDN U4566 ( .A(n2867), .B(n3718), .Z(n2868) );
  XNOR U4567 ( .A(n4155), .B(n2868), .Z(out[261]) );
  XNOR U4568 ( .A(n3957), .B(in[1416]), .Z(n4193) );
  NANDN U4569 ( .A(n2869), .B(n4158), .Z(n2870) );
  XNOR U4570 ( .A(n4193), .B(n2870), .Z(out[262]) );
  XNOR U4571 ( .A(in[1417]), .B(n3961), .Z(n4440) );
  NANDN U4572 ( .A(n2871), .B(n4439), .Z(n2872) );
  XNOR U4573 ( .A(n4440), .B(n2872), .Z(out[263]) );
  XNOR U4574 ( .A(n3965), .B(in[1418]), .Z(n4731) );
  NANDN U4575 ( .A(n2873), .B(n4730), .Z(n2874) );
  XNOR U4576 ( .A(n4731), .B(n2874), .Z(out[264]) );
  XNOR U4577 ( .A(n3969), .B(in[1419]), .Z(n5162) );
  NANDN U4578 ( .A(n2875), .B(n5161), .Z(n2876) );
  XNOR U4579 ( .A(n5162), .B(n2876), .Z(out[265]) );
  NOR U4580 ( .A(n2878), .B(n2877), .Z(n2879) );
  XOR U4581 ( .A(n4281), .B(n2879), .Z(out[266]) );
  XOR U4582 ( .A(in[1436]), .B(n2886), .Z(n4775) );
  OR U4583 ( .A(n4775), .B(n2887), .Z(n2888) );
  XNOR U4584 ( .A(n4774), .B(n2888), .Z(out[26]) );
  NOR U4585 ( .A(n2890), .B(n2889), .Z(n2891) );
  XOR U4586 ( .A(n4402), .B(n2891), .Z(out[270]) );
  NOR U4587 ( .A(n2893), .B(n2892), .Z(n2894) );
  XOR U4588 ( .A(n4436), .B(n2894), .Z(out[271]) );
  NOR U4589 ( .A(n2896), .B(n2895), .Z(n2897) );
  XOR U4590 ( .A(n4474), .B(n2897), .Z(out[272]) );
  NOR U4591 ( .A(n2899), .B(n2898), .Z(n2900) );
  XOR U4592 ( .A(n4508), .B(n2900), .Z(out[273]) );
  NOR U4593 ( .A(n2902), .B(n2901), .Z(n2903) );
  XOR U4594 ( .A(n4547), .B(n2903), .Z(out[274]) );
  NOR U4595 ( .A(n2905), .B(n2904), .Z(n2906) );
  XOR U4596 ( .A(n4576), .B(n2906), .Z(out[275]) );
  NOR U4597 ( .A(n2908), .B(n2907), .Z(n2909) );
  XOR U4598 ( .A(n4601), .B(n2909), .Z(out[276]) );
  ANDN U4599 ( .B(n2911), .A(n2910), .Z(n2912) );
  XOR U4600 ( .A(n4629), .B(n2912), .Z(out[277]) );
  ANDN U4601 ( .B(n2914), .A(n2913), .Z(n2915) );
  XOR U4602 ( .A(n4660), .B(n2915), .Z(out[278]) );
  ANDN U4603 ( .B(n2917), .A(n2916), .Z(n2918) );
  XOR U4604 ( .A(n4677), .B(n2918), .Z(out[279]) );
  XOR U4605 ( .A(in[1437]), .B(n2919), .Z(n4819) );
  OR U4606 ( .A(n4819), .B(n2920), .Z(n2921) );
  XNOR U4607 ( .A(n4818), .B(n2921), .Z(out[27]) );
  ANDN U4608 ( .B(n2923), .A(n2922), .Z(n2924) );
  XOR U4609 ( .A(n4693), .B(n2924), .Z(out[280]) );
  ANDN U4610 ( .B(n2926), .A(n2925), .Z(n2927) );
  XOR U4611 ( .A(n4727), .B(n2927), .Z(out[281]) );
  ANDN U4612 ( .B(n2929), .A(n2928), .Z(n2930) );
  XOR U4613 ( .A(n4775), .B(n2930), .Z(out[282]) );
  ANDN U4614 ( .B(n2932), .A(n2931), .Z(n2933) );
  XOR U4615 ( .A(n4819), .B(n2933), .Z(out[283]) );
  XOR U4616 ( .A(in[1438]), .B(n4052), .Z(n4862) );
  NAND U4617 ( .A(n2934), .B(n2946), .Z(n2935) );
  XNOR U4618 ( .A(n4862), .B(n2935), .Z(out[284]) );
  XOR U4619 ( .A(in[1439]), .B(n4056), .Z(n4906) );
  NAND U4620 ( .A(n2936), .B(n2968), .Z(n2937) );
  XNOR U4621 ( .A(n4906), .B(n2937), .Z(out[285]) );
  XOR U4622 ( .A(in[1440]), .B(n4060), .Z(n4950) );
  NAND U4623 ( .A(n2938), .B(n2992), .Z(n2939) );
  XNOR U4624 ( .A(n4950), .B(n2939), .Z(out[286]) );
  XOR U4625 ( .A(in[1441]), .B(n4064), .Z(n4994) );
  NAND U4626 ( .A(n2940), .B(n3020), .Z(n2941) );
  XNOR U4627 ( .A(n4994), .B(n2941), .Z(out[287]) );
  XOR U4628 ( .A(in[1442]), .B(n4072), .Z(n5038) );
  NAND U4629 ( .A(n2942), .B(n3040), .Z(n2943) );
  XNOR U4630 ( .A(n5038), .B(n2943), .Z(out[288]) );
  XOR U4631 ( .A(in[1443]), .B(n4076), .Z(n5079) );
  NAND U4632 ( .A(n2944), .B(n3052), .Z(n2945) );
  XNOR U4633 ( .A(n5079), .B(n2945), .Z(out[289]) );
  OR U4634 ( .A(n4862), .B(n2946), .Z(n2947) );
  XOR U4635 ( .A(n4863), .B(n2947), .Z(out[28]) );
  XOR U4636 ( .A(in[1444]), .B(n4080), .Z(n5115) );
  NAND U4637 ( .A(n2948), .B(n3073), .Z(n2949) );
  XNOR U4638 ( .A(n5115), .B(n2949), .Z(out[290]) );
  XNOR U4639 ( .A(in[1445]), .B(n4084), .Z(n5158) );
  NANDN U4640 ( .A(n2950), .B(n3094), .Z(n2951) );
  XNOR U4641 ( .A(n5158), .B(n2951), .Z(out[291]) );
  OR U4642 ( .A(n3111), .B(n2952), .Z(n2953) );
  XNOR U4643 ( .A(n3110), .B(n2953), .Z(out[292]) );
  OR U4644 ( .A(n3133), .B(n2954), .Z(n2955) );
  XNOR U4645 ( .A(n3132), .B(n2955), .Z(out[293]) );
  NANDN U4646 ( .A(n2956), .B(n3151), .Z(n2957) );
  XNOR U4647 ( .A(n3152), .B(n2957), .Z(out[294]) );
  OR U4648 ( .A(n3163), .B(n2958), .Z(n2959) );
  XNOR U4649 ( .A(n3162), .B(n2959), .Z(out[295]) );
  OR U4650 ( .A(n3188), .B(n2960), .Z(n2961) );
  XNOR U4651 ( .A(n3187), .B(n2961), .Z(out[296]) );
  OR U4652 ( .A(n3218), .B(n2962), .Z(n2963) );
  XOR U4653 ( .A(n3219), .B(n2963), .Z(out[297]) );
  OR U4654 ( .A(n3242), .B(n2964), .Z(n2965) );
  XOR U4655 ( .A(n3243), .B(n2965), .Z(out[298]) );
  OR U4656 ( .A(n3254), .B(n2966), .Z(n2967) );
  XOR U4657 ( .A(n3255), .B(n2967), .Z(out[299]) );
  OR U4658 ( .A(n4906), .B(n2968), .Z(n2969) );
  XOR U4659 ( .A(n4907), .B(n2969), .Z(out[29]) );
  OR U4660 ( .A(n4023), .B(n2970), .Z(n2971) );
  XNOR U4661 ( .A(n4022), .B(n2971), .Z(out[2]) );
  OR U4662 ( .A(n3264), .B(n2972), .Z(n2973) );
  XOR U4663 ( .A(n3265), .B(n2973), .Z(out[300]) );
  OR U4664 ( .A(n3298), .B(n2974), .Z(n2975) );
  XOR U4665 ( .A(n3299), .B(n2975), .Z(out[301]) );
  OR U4666 ( .A(n3328), .B(n2976), .Z(n2977) );
  XOR U4667 ( .A(n3329), .B(n2977), .Z(out[302]) );
  NANDN U4668 ( .A(n2978), .B(n3357), .Z(n2979) );
  XOR U4669 ( .A(n3358), .B(n2979), .Z(out[303]) );
  OR U4670 ( .A(n3385), .B(n2980), .Z(n2981) );
  XOR U4671 ( .A(n3386), .B(n2981), .Z(out[304]) );
  NANDN U4672 ( .A(n2983), .B(n3455), .Z(n2984) );
  XOR U4673 ( .A(n3456), .B(n2984), .Z(out[306]) );
  NANDN U4674 ( .A(n2985), .B(n3477), .Z(n2986) );
  XOR U4675 ( .A(n3478), .B(n2986), .Z(out[307]) );
  NANDN U4676 ( .A(n2987), .B(n3499), .Z(n2988) );
  XOR U4677 ( .A(n3500), .B(n2988), .Z(out[308]) );
  IV U4678 ( .A(n2989), .Z(n3514) );
  NANDN U4679 ( .A(n2990), .B(n3514), .Z(n2991) );
  XOR U4680 ( .A(n3515), .B(n2991), .Z(out[309]) );
  OR U4681 ( .A(n4950), .B(n2992), .Z(n2993) );
  XOR U4682 ( .A(n4951), .B(n2993), .Z(out[30]) );
  IV U4683 ( .A(n2994), .Z(n3542) );
  NANDN U4684 ( .A(n2995), .B(n3542), .Z(n2996) );
  XOR U4685 ( .A(n3543), .B(n2996), .Z(out[310]) );
  IV U4686 ( .A(n2997), .Z(n3572) );
  NANDN U4687 ( .A(n2998), .B(n3572), .Z(n2999) );
  XOR U4688 ( .A(n3573), .B(n2999), .Z(out[311]) );
  IV U4689 ( .A(n3000), .Z(n3596) );
  NANDN U4690 ( .A(n3001), .B(n3596), .Z(n3002) );
  XOR U4691 ( .A(n3597), .B(n3002), .Z(out[312]) );
  NANDN U4692 ( .A(n3003), .B(n3626), .Z(n3004) );
  XOR U4693 ( .A(n3627), .B(n3004), .Z(out[313]) );
  NANDN U4694 ( .A(n3005), .B(n3670), .Z(n3006) );
  XOR U4695 ( .A(n3671), .B(n3006), .Z(out[314]) );
  NANDN U4696 ( .A(n3008), .B(n3007), .Z(n3009) );
  XOR U4697 ( .A(n3715), .B(n3009), .Z(out[315]) );
  NANDN U4698 ( .A(n3011), .B(n3010), .Z(n3012) );
  XOR U4699 ( .A(n3761), .B(n3012), .Z(out[316]) );
  NANDN U4700 ( .A(n3015), .B(n3014), .Z(n3016) );
  XOR U4701 ( .A(n3849), .B(n3016), .Z(out[318]) );
  NANDN U4702 ( .A(n3018), .B(n3017), .Z(n3019) );
  XOR U4703 ( .A(n3893), .B(n3019), .Z(out[319]) );
  OR U4704 ( .A(n4994), .B(n3020), .Z(n3021) );
  XOR U4705 ( .A(n4995), .B(n3021), .Z(out[31]) );
  XOR U4706 ( .A(in[72]), .B(n4446), .Z(n3259) );
  XOR U4707 ( .A(in[1317]), .B(n4278), .Z(n3613) );
  XNOR U4708 ( .A(in[1244]), .B(n3022), .Z(n3610) );
  NANDN U4709 ( .A(n3613), .B(n3610), .Z(n3023) );
  XNOR U4710 ( .A(n3259), .B(n3023), .Z(out[320]) );
  XOR U4711 ( .A(in[73]), .B(n4449), .Z(n3145) );
  IV U4712 ( .A(n3145), .Z(n3262) );
  XOR U4713 ( .A(in[1318]), .B(n4284), .Z(n3617) );
  XNOR U4714 ( .A(in[1245]), .B(n3024), .Z(n3614) );
  NANDN U4715 ( .A(n3617), .B(n3614), .Z(n3025) );
  XOR U4716 ( .A(n3262), .B(n3025), .Z(out[321]) );
  XOR U4717 ( .A(in[74]), .B(n4452), .Z(n3147) );
  IV U4718 ( .A(n3147), .Z(n3269) );
  XOR U4719 ( .A(in[1319]), .B(n4286), .Z(n3621) );
  XNOR U4720 ( .A(in[1246]), .B(n3026), .Z(n3618) );
  NANDN U4721 ( .A(n3621), .B(n3618), .Z(n3027) );
  XOR U4722 ( .A(n3269), .B(n3027), .Z(out[322]) );
  XOR U4723 ( .A(in[75]), .B(n4455), .Z(n3149) );
  IV U4724 ( .A(n3149), .Z(n3272) );
  XOR U4725 ( .A(in[1320]), .B(n4288), .Z(n3625) );
  XNOR U4726 ( .A(in[1247]), .B(n3028), .Z(n3622) );
  NANDN U4727 ( .A(n3625), .B(n3622), .Z(n3029) );
  XOR U4728 ( .A(n3272), .B(n3029), .Z(out[323]) );
  XNOR U4729 ( .A(n4458), .B(in[76]), .Z(n3275) );
  XOR U4730 ( .A(in[1321]), .B(n4290), .Z(n3633) );
  XNOR U4731 ( .A(in[1248]), .B(n3030), .Z(n3630) );
  NANDN U4732 ( .A(n3633), .B(n3630), .Z(n3031) );
  XNOR U4733 ( .A(n3275), .B(n3031), .Z(out[324]) );
  XNOR U4734 ( .A(n4461), .B(in[77]), .Z(n3278) );
  XOR U4735 ( .A(in[1322]), .B(n4292), .Z(n3637) );
  XNOR U4736 ( .A(in[1249]), .B(n3032), .Z(n3634) );
  NANDN U4737 ( .A(n3637), .B(n3634), .Z(n3033) );
  XNOR U4738 ( .A(n3278), .B(n3033), .Z(out[325]) );
  XNOR U4739 ( .A(n4464), .B(in[78]), .Z(n3281) );
  XOR U4740 ( .A(in[1323]), .B(n4294), .Z(n3641) );
  XNOR U4741 ( .A(in[1250]), .B(n4122), .Z(n3638) );
  NANDN U4742 ( .A(n3641), .B(n3638), .Z(n3034) );
  XNOR U4743 ( .A(n3281), .B(n3034), .Z(out[326]) );
  XNOR U4744 ( .A(n4467), .B(in[79]), .Z(n3284) );
  XOR U4745 ( .A(in[1324]), .B(n4296), .Z(n3645) );
  XNOR U4746 ( .A(in[1251]), .B(n3035), .Z(n3642) );
  NANDN U4747 ( .A(n3645), .B(n3642), .Z(n3036) );
  XNOR U4748 ( .A(n3284), .B(n3036), .Z(out[327]) );
  XNOR U4749 ( .A(n4470), .B(in[80]), .Z(n3287) );
  XOR U4750 ( .A(in[1325]), .B(n4298), .Z(n3649) );
  XNOR U4751 ( .A(in[1252]), .B(n3037), .Z(n3646) );
  NANDN U4752 ( .A(n3649), .B(n3646), .Z(n3038) );
  XNOR U4753 ( .A(n3287), .B(n3038), .Z(out[328]) );
  XNOR U4754 ( .A(n4477), .B(in[81]), .Z(n3290) );
  XNOR U4755 ( .A(in[1253]), .B(n4134), .Z(n3651) );
  XNOR U4756 ( .A(in[1326]), .B(n4300), .Z(n3653) );
  NANDN U4757 ( .A(n3651), .B(n3653), .Z(n3039) );
  XNOR U4758 ( .A(n3290), .B(n3039), .Z(out[329]) );
  OR U4759 ( .A(n5038), .B(n3040), .Z(n3041) );
  XOR U4760 ( .A(n5039), .B(n3041), .Z(out[32]) );
  XNOR U4761 ( .A(n4480), .B(in[82]), .Z(n3293) );
  XNOR U4762 ( .A(in[1254]), .B(n4138), .Z(n3655) );
  XNOR U4763 ( .A(in[1327]), .B(n4302), .Z(n3657) );
  NANDN U4764 ( .A(n3655), .B(n3657), .Z(n3042) );
  XNOR U4765 ( .A(n3293), .B(n3042), .Z(out[330]) );
  XNOR U4766 ( .A(n4483), .B(in[83]), .Z(n3296) );
  XNOR U4767 ( .A(in[1255]), .B(n4142), .Z(n3659) );
  XNOR U4768 ( .A(in[1328]), .B(n4309), .Z(n3661) );
  NANDN U4769 ( .A(n3659), .B(n3661), .Z(n3043) );
  XNOR U4770 ( .A(n3296), .B(n3043), .Z(out[331]) );
  XNOR U4771 ( .A(in[84]), .B(n4486), .Z(n3303) );
  XNOR U4772 ( .A(in[1256]), .B(n4146), .Z(n3663) );
  XNOR U4773 ( .A(in[1329]), .B(n4312), .Z(n3665) );
  NANDN U4774 ( .A(n3663), .B(n3665), .Z(n3044) );
  XNOR U4775 ( .A(n3303), .B(n3044), .Z(out[332]) );
  XNOR U4776 ( .A(in[85]), .B(n4489), .Z(n3306) );
  XNOR U4777 ( .A(in[1257]), .B(n4150), .Z(n3667) );
  XNOR U4778 ( .A(in[1330]), .B(n4315), .Z(n3669) );
  NANDN U4779 ( .A(n3667), .B(n3669), .Z(n3045) );
  XNOR U4780 ( .A(n3306), .B(n3045), .Z(out[333]) );
  XNOR U4781 ( .A(in[86]), .B(n4492), .Z(n3309) );
  XNOR U4782 ( .A(in[1258]), .B(n4160), .Z(n3675) );
  XNOR U4783 ( .A(in[1331]), .B(n4318), .Z(n3677) );
  NANDN U4784 ( .A(n3675), .B(n3677), .Z(n3046) );
  XNOR U4785 ( .A(n3309), .B(n3046), .Z(out[334]) );
  XNOR U4786 ( .A(in[87]), .B(n4495), .Z(n3312) );
  XNOR U4787 ( .A(in[1259]), .B(n4164), .Z(n3679) );
  XNOR U4788 ( .A(in[1332]), .B(n4321), .Z(n3681) );
  NANDN U4789 ( .A(n3679), .B(n3681), .Z(n3047) );
  XNOR U4790 ( .A(n3312), .B(n3047), .Z(out[335]) );
  XNOR U4791 ( .A(in[88]), .B(n4498), .Z(n3315) );
  XNOR U4792 ( .A(in[1260]), .B(n4168), .Z(n3683) );
  XNOR U4793 ( .A(in[1333]), .B(n4324), .Z(n3685) );
  NANDN U4794 ( .A(n3683), .B(n3685), .Z(n3048) );
  XNOR U4795 ( .A(n3315), .B(n3048), .Z(out[336]) );
  XNOR U4796 ( .A(in[89]), .B(n4501), .Z(n3318) );
  XNOR U4797 ( .A(in[1261]), .B(n4172), .Z(n3687) );
  XNOR U4798 ( .A(in[1334]), .B(n4327), .Z(n3689) );
  NANDN U4799 ( .A(n3687), .B(n3689), .Z(n3049) );
  XNOR U4800 ( .A(n3318), .B(n3049), .Z(out[337]) );
  XNOR U4801 ( .A(in[90]), .B(n4504), .Z(n3320) );
  XNOR U4802 ( .A(in[1262]), .B(n3896), .Z(n3691) );
  XNOR U4803 ( .A(in[1335]), .B(n4330), .Z(n3693) );
  NANDN U4804 ( .A(n3691), .B(n3693), .Z(n3050) );
  XNOR U4805 ( .A(n3320), .B(n3050), .Z(out[338]) );
  XOR U4806 ( .A(in[91]), .B(n4511), .Z(n3322) );
  XNOR U4807 ( .A(in[1263]), .B(n3900), .Z(n3695) );
  XNOR U4808 ( .A(in[1336]), .B(n4176), .Z(n3697) );
  NANDN U4809 ( .A(n3695), .B(n3697), .Z(n3051) );
  XNOR U4810 ( .A(n3322), .B(n3051), .Z(out[339]) );
  OR U4811 ( .A(n5079), .B(n3052), .Z(n3053) );
  XOR U4812 ( .A(n5080), .B(n3053), .Z(out[33]) );
  XOR U4813 ( .A(in[92]), .B(n4514), .Z(n3324) );
  XNOR U4814 ( .A(in[1264]), .B(n3904), .Z(n3699) );
  XNOR U4815 ( .A(in[1337]), .B(n4179), .Z(n3701) );
  NANDN U4816 ( .A(n3699), .B(n3701), .Z(n3054) );
  XNOR U4817 ( .A(n3324), .B(n3054), .Z(out[340]) );
  XOR U4818 ( .A(in[93]), .B(n4517), .Z(n3326) );
  XNOR U4819 ( .A(in[1265]), .B(n3908), .Z(n3703) );
  XNOR U4820 ( .A(in[1338]), .B(n4182), .Z(n3705) );
  NANDN U4821 ( .A(n3703), .B(n3705), .Z(n3055) );
  XNOR U4822 ( .A(n3326), .B(n3055), .Z(out[341]) );
  XNOR U4823 ( .A(in[94]), .B(n4520), .Z(n3332) );
  XNOR U4824 ( .A(in[1266]), .B(n3912), .Z(n3707) );
  XNOR U4825 ( .A(in[1339]), .B(n4185), .Z(n3709) );
  NANDN U4826 ( .A(n3707), .B(n3709), .Z(n3056) );
  XNOR U4827 ( .A(n3332), .B(n3056), .Z(out[342]) );
  XNOR U4828 ( .A(in[95]), .B(n4524), .Z(n3334) );
  XOR U4829 ( .A(in[1267]), .B(n3916), .Z(n3711) );
  XNOR U4830 ( .A(in[1340]), .B(n3057), .Z(n3713) );
  NANDN U4831 ( .A(n3711), .B(n3713), .Z(n3058) );
  XNOR U4832 ( .A(n3334), .B(n3058), .Z(out[343]) );
  XNOR U4833 ( .A(in[96]), .B(n4528), .Z(n3336) );
  XOR U4834 ( .A(in[1268]), .B(n3920), .Z(n3721) );
  XNOR U4835 ( .A(in[1341]), .B(n3059), .Z(n3723) );
  NANDN U4836 ( .A(n3721), .B(n3723), .Z(n3060) );
  XNOR U4837 ( .A(n3336), .B(n3060), .Z(out[344]) );
  XNOR U4838 ( .A(in[97]), .B(n4532), .Z(n3338) );
  XOR U4839 ( .A(in[1269]), .B(n3924), .Z(n3725) );
  XNOR U4840 ( .A(in[1342]), .B(n3061), .Z(n3727) );
  NANDN U4841 ( .A(n3725), .B(n3727), .Z(n3062) );
  XNOR U4842 ( .A(n3338), .B(n3062), .Z(out[345]) );
  XNOR U4843 ( .A(in[98]), .B(n4536), .Z(n3340) );
  IV U4844 ( .A(n3063), .Z(n3928) );
  XOR U4845 ( .A(in[1270]), .B(n3928), .Z(n3729) );
  XNOR U4846 ( .A(in[1343]), .B(n4197), .Z(n3731) );
  NANDN U4847 ( .A(n3729), .B(n3731), .Z(n3064) );
  XNOR U4848 ( .A(n3340), .B(n3064), .Z(out[346]) );
  XNOR U4849 ( .A(in[99]), .B(n4540), .Z(n3342) );
  IV U4850 ( .A(n3065), .Z(n3932) );
  XOR U4851 ( .A(in[1271]), .B(n3932), .Z(n3733) );
  XNOR U4852 ( .A(in[1280]), .B(n3066), .Z(n3735) );
  NANDN U4853 ( .A(n3733), .B(n3735), .Z(n3067) );
  XNOR U4854 ( .A(n3342), .B(n3067), .Z(out[347]) );
  XOR U4855 ( .A(in[100]), .B(n4544), .Z(n3195) );
  IV U4856 ( .A(n3195), .Z(n3345) );
  IV U4857 ( .A(n3068), .Z(n3939) );
  XOR U4858 ( .A(in[1272]), .B(n3939), .Z(n3737) );
  XNOR U4859 ( .A(in[1281]), .B(n3069), .Z(n3739) );
  NANDN U4860 ( .A(n3737), .B(n3739), .Z(n3070) );
  XOR U4861 ( .A(n3345), .B(n3070), .Z(out[348]) );
  XOR U4862 ( .A(in[101]), .B(n4550), .Z(n3198) );
  IV U4863 ( .A(n3198), .Z(n3349) );
  XOR U4864 ( .A(in[1273]), .B(n3943), .Z(n3741) );
  XNOR U4865 ( .A(in[1282]), .B(n3071), .Z(n3743) );
  NANDN U4866 ( .A(n3741), .B(n3743), .Z(n3072) );
  XOR U4867 ( .A(n3349), .B(n3072), .Z(out[349]) );
  OR U4868 ( .A(n5115), .B(n3073), .Z(n3074) );
  XNOR U4869 ( .A(n5114), .B(n3074), .Z(out[34]) );
  XOR U4870 ( .A(in[102]), .B(n4552), .Z(n3201) );
  IV U4871 ( .A(n3201), .Z(n3352) );
  XOR U4872 ( .A(in[1274]), .B(n3947), .Z(n3745) );
  XNOR U4873 ( .A(in[1283]), .B(n3075), .Z(n3747) );
  NANDN U4874 ( .A(n3745), .B(n3747), .Z(n3076) );
  XOR U4875 ( .A(n3352), .B(n3076), .Z(out[350]) );
  XOR U4876 ( .A(in[103]), .B(n4333), .Z(n3204) );
  IV U4877 ( .A(n3204), .Z(n3355) );
  XNOR U4878 ( .A(in[1275]), .B(n3951), .Z(n3749) );
  XNOR U4879 ( .A(in[1284]), .B(n3077), .Z(n3751) );
  NANDN U4880 ( .A(n3749), .B(n3751), .Z(n3078) );
  XOR U4881 ( .A(n3355), .B(n3078), .Z(out[351]) );
  XOR U4882 ( .A(in[104]), .B(n4335), .Z(n3207) );
  IV U4883 ( .A(n3207), .Z(n3362) );
  XNOR U4884 ( .A(in[1276]), .B(n3955), .Z(n3753) );
  XNOR U4885 ( .A(in[1285]), .B(n3079), .Z(n3755) );
  NANDN U4886 ( .A(n3753), .B(n3755), .Z(n3080) );
  XOR U4887 ( .A(n3362), .B(n3080), .Z(out[352]) );
  XOR U4888 ( .A(in[105]), .B(n4341), .Z(n3210) );
  IV U4889 ( .A(n3210), .Z(n3365) );
  XNOR U4890 ( .A(in[1277]), .B(n3959), .Z(n3757) );
  XNOR U4891 ( .A(in[1286]), .B(n3081), .Z(n3759) );
  NANDN U4892 ( .A(n3757), .B(n3759), .Z(n3082) );
  XOR U4893 ( .A(n3365), .B(n3082), .Z(out[353]) );
  XOR U4894 ( .A(in[106]), .B(n4343), .Z(n3213) );
  IV U4895 ( .A(n3213), .Z(n3368) );
  XNOR U4896 ( .A(in[1278]), .B(n3963), .Z(n3765) );
  XNOR U4897 ( .A(in[1287]), .B(n3083), .Z(n3767) );
  NANDN U4898 ( .A(n3765), .B(n3767), .Z(n3084) );
  XOR U4899 ( .A(n3368), .B(n3084), .Z(out[354]) );
  XOR U4900 ( .A(in[107]), .B(n4345), .Z(n3216) );
  IV U4901 ( .A(n3216), .Z(n3371) );
  XNOR U4902 ( .A(in[1279]), .B(n3967), .Z(n3769) );
  XNOR U4903 ( .A(in[1288]), .B(n4214), .Z(n3771) );
  NANDN U4904 ( .A(n3769), .B(n3771), .Z(n3085) );
  XOR U4905 ( .A(n3371), .B(n3085), .Z(out[355]) );
  XOR U4906 ( .A(in[108]), .B(n4348), .Z(n3222) );
  IV U4907 ( .A(n3222), .Z(n3373) );
  XNOR U4908 ( .A(in[1216]), .B(n3971), .Z(n3773) );
  XNOR U4909 ( .A(in[1289]), .B(n3086), .Z(n3775) );
  NANDN U4910 ( .A(n3773), .B(n3775), .Z(n3087) );
  XOR U4911 ( .A(n3373), .B(n3087), .Z(out[356]) );
  XOR U4912 ( .A(in[109]), .B(n4351), .Z(n3224) );
  IV U4913 ( .A(n3224), .Z(n3375) );
  XNOR U4914 ( .A(in[1217]), .B(n3975), .Z(n3777) );
  XNOR U4915 ( .A(in[1290]), .B(n3088), .Z(n3779) );
  NANDN U4916 ( .A(n3777), .B(n3779), .Z(n3089) );
  XOR U4917 ( .A(n3375), .B(n3089), .Z(out[357]) );
  XOR U4918 ( .A(in[110]), .B(n4354), .Z(n3226) );
  IV U4919 ( .A(n3226), .Z(n3377) );
  XNOR U4920 ( .A(in[1218]), .B(n3982), .Z(n3781) );
  XNOR U4921 ( .A(in[1291]), .B(n3090), .Z(n3783) );
  NANDN U4922 ( .A(n3781), .B(n3783), .Z(n3091) );
  XOR U4923 ( .A(n3377), .B(n3091), .Z(out[358]) );
  XOR U4924 ( .A(in[111]), .B(n4356), .Z(n3228) );
  IV U4925 ( .A(n3228), .Z(n3379) );
  XNOR U4926 ( .A(in[1219]), .B(n3986), .Z(n3785) );
  XNOR U4927 ( .A(in[1292]), .B(n3092), .Z(n3787) );
  NANDN U4928 ( .A(n3785), .B(n3787), .Z(n3093) );
  XOR U4929 ( .A(n3379), .B(n3093), .Z(out[359]) );
  OR U4930 ( .A(n5158), .B(n3094), .Z(n3095) );
  XNOR U4931 ( .A(n5157), .B(n3095), .Z(out[35]) );
  XOR U4932 ( .A(in[112]), .B(n4359), .Z(n3230) );
  IV U4933 ( .A(n3230), .Z(n3381) );
  XOR U4934 ( .A(in[1293]), .B(n3096), .Z(n3791) );
  XOR U4935 ( .A(in[1220]), .B(n3990), .Z(n3788) );
  NANDN U4936 ( .A(n3791), .B(n3788), .Z(n3097) );
  XOR U4937 ( .A(n3381), .B(n3097), .Z(out[360]) );
  XOR U4938 ( .A(in[113]), .B(n4362), .Z(n3232) );
  IV U4939 ( .A(n3232), .Z(n3383) );
  XOR U4940 ( .A(in[1294]), .B(n4232), .Z(n3795) );
  XOR U4941 ( .A(in[1221]), .B(n3994), .Z(n3792) );
  NANDN U4942 ( .A(n3795), .B(n3792), .Z(n3098) );
  XOR U4943 ( .A(n3383), .B(n3098), .Z(out[361]) );
  XOR U4944 ( .A(in[114]), .B(n4365), .Z(n3234) );
  IV U4945 ( .A(n3234), .Z(n3389) );
  XOR U4946 ( .A(in[1295]), .B(n4235), .Z(n3799) );
  XOR U4947 ( .A(in[1222]), .B(n3998), .Z(n3796) );
  NANDN U4948 ( .A(n3799), .B(n3796), .Z(n3099) );
  XOR U4949 ( .A(n3389), .B(n3099), .Z(out[362]) );
  XOR U4950 ( .A(in[115]), .B(n4372), .Z(n3236) );
  IV U4951 ( .A(n3236), .Z(n3391) );
  XOR U4952 ( .A(in[1296]), .B(n4238), .Z(n3803) );
  XOR U4953 ( .A(in[1223]), .B(n4002), .Z(n3800) );
  NANDN U4954 ( .A(n3803), .B(n3800), .Z(n3100) );
  XOR U4955 ( .A(n3391), .B(n3100), .Z(out[363]) );
  XOR U4956 ( .A(in[116]), .B(n4375), .Z(n3238) );
  IV U4957 ( .A(n3238), .Z(n3394) );
  XOR U4958 ( .A(in[1297]), .B(n4239), .Z(n3811) );
  XOR U4959 ( .A(in[1224]), .B(n4006), .Z(n3808) );
  NANDN U4960 ( .A(n3811), .B(n3808), .Z(n3101) );
  XOR U4961 ( .A(n3394), .B(n3101), .Z(out[364]) );
  XOR U4962 ( .A(in[117]), .B(n4378), .Z(n3240) );
  IV U4963 ( .A(n3240), .Z(n3398) );
  XOR U4964 ( .A(in[1298]), .B(n3102), .Z(n3815) );
  XOR U4965 ( .A(in[1225]), .B(n4010), .Z(n3812) );
  NANDN U4966 ( .A(n3815), .B(n3812), .Z(n3103) );
  XOR U4967 ( .A(n3398), .B(n3103), .Z(out[365]) );
  XOR U4968 ( .A(in[118]), .B(n4381), .Z(n3246) );
  IV U4969 ( .A(n3246), .Z(n3402) );
  XOR U4970 ( .A(in[1299]), .B(n3104), .Z(n3819) );
  XOR U4971 ( .A(in[1226]), .B(n4014), .Z(n3816) );
  NANDN U4972 ( .A(n3819), .B(n3816), .Z(n3105) );
  XOR U4973 ( .A(n3402), .B(n3105), .Z(out[366]) );
  XOR U4974 ( .A(in[119]), .B(n4384), .Z(n3248) );
  IV U4975 ( .A(n3248), .Z(n3406) );
  XOR U4976 ( .A(in[1300]), .B(n4246), .Z(n3823) );
  XOR U4977 ( .A(in[1227]), .B(n4018), .Z(n3820) );
  NANDN U4978 ( .A(n3823), .B(n3820), .Z(n3106) );
  XOR U4979 ( .A(n3406), .B(n3106), .Z(out[367]) );
  XOR U4980 ( .A(in[120]), .B(n4386), .Z(n3250) );
  IV U4981 ( .A(n3250), .Z(n3409) );
  XOR U4982 ( .A(in[1301]), .B(n4249), .Z(n3827) );
  XOR U4983 ( .A(in[1228]), .B(n4026), .Z(n3824) );
  NANDN U4984 ( .A(n3827), .B(n3824), .Z(n3107) );
  XOR U4985 ( .A(n3409), .B(n3107), .Z(out[368]) );
  XOR U4986 ( .A(in[121]), .B(n4389), .Z(n3252) );
  IV U4987 ( .A(n3252), .Z(n3412) );
  XOR U4988 ( .A(in[1302]), .B(n4250), .Z(n3831) );
  XNOR U4989 ( .A(in[1229]), .B(n3108), .Z(n3828) );
  NANDN U4990 ( .A(n3831), .B(n3828), .Z(n3109) );
  XOR U4991 ( .A(n3412), .B(n3109), .Z(out[369]) );
  ANDN U4992 ( .B(n3111), .A(n3110), .Z(n3112) );
  XOR U4993 ( .A(n3113), .B(n3112), .Z(out[36]) );
  XOR U4994 ( .A(in[122]), .B(n4392), .Z(n3415) );
  XOR U4995 ( .A(in[1303]), .B(n4251), .Z(n3835) );
  XNOR U4996 ( .A(in[1230]), .B(n3114), .Z(n3832) );
  NANDN U4997 ( .A(n3835), .B(n3832), .Z(n3115) );
  XOR U4998 ( .A(n3415), .B(n3115), .Z(out[370]) );
  XOR U4999 ( .A(in[123]), .B(n4395), .Z(n3418) );
  XOR U5000 ( .A(in[1304]), .B(n4252), .Z(n3839) );
  XNOR U5001 ( .A(in[1231]), .B(n3116), .Z(n3836) );
  NANDN U5002 ( .A(n3839), .B(n3836), .Z(n3117) );
  XOR U5003 ( .A(n3418), .B(n3117), .Z(out[371]) );
  XOR U5004 ( .A(in[124]), .B(n4398), .Z(n3426) );
  XOR U5005 ( .A(in[1305]), .B(n4253), .Z(n3843) );
  XNOR U5006 ( .A(in[1232]), .B(n3118), .Z(n3840) );
  NANDN U5007 ( .A(n3843), .B(n3840), .Z(n3119) );
  XNOR U5008 ( .A(n3426), .B(n3119), .Z(out[372]) );
  XOR U5009 ( .A(in[125]), .B(n4405), .Z(n3429) );
  XOR U5010 ( .A(in[1306]), .B(n4254), .Z(n3847) );
  XNOR U5011 ( .A(in[1233]), .B(n4046), .Z(n3844) );
  NANDN U5012 ( .A(n3847), .B(n3844), .Z(n3120) );
  XNOR U5013 ( .A(n3429), .B(n3120), .Z(out[373]) );
  XOR U5014 ( .A(in[126]), .B(n4408), .Z(n3432) );
  XOR U5015 ( .A(in[1307]), .B(n4255), .Z(n3855) );
  XOR U5016 ( .A(in[1234]), .B(n4050), .Z(n3852) );
  NANDN U5017 ( .A(n3855), .B(n3852), .Z(n3121) );
  XNOR U5018 ( .A(n3432), .B(n3121), .Z(out[374]) );
  XOR U5019 ( .A(in[127]), .B(n4411), .Z(n3435) );
  XOR U5020 ( .A(in[1308]), .B(n4258), .Z(n3859) );
  XNOR U5021 ( .A(in[1235]), .B(n3122), .Z(n3856) );
  NANDN U5022 ( .A(n3859), .B(n3856), .Z(n3123) );
  XNOR U5023 ( .A(n3435), .B(n3123), .Z(out[375]) );
  XOR U5024 ( .A(in[64]), .B(n4414), .Z(n3438) );
  XOR U5025 ( .A(in[1309]), .B(n4259), .Z(n3863) );
  XNOR U5026 ( .A(in[1236]), .B(n3124), .Z(n3860) );
  NANDN U5027 ( .A(n3863), .B(n3860), .Z(n3125) );
  XNOR U5028 ( .A(n3438), .B(n3125), .Z(out[376]) );
  XOR U5029 ( .A(in[65]), .B(n4417), .Z(n3441) );
  XOR U5030 ( .A(in[1310]), .B(n4260), .Z(n3867) );
  XNOR U5031 ( .A(in[1237]), .B(n3126), .Z(n3864) );
  NANDN U5032 ( .A(n3867), .B(n3864), .Z(n3127) );
  XNOR U5033 ( .A(n3441), .B(n3127), .Z(out[377]) );
  XOR U5034 ( .A(in[66]), .B(n4420), .Z(n3444) );
  XOR U5035 ( .A(in[1311]), .B(n4261), .Z(n3871) );
  XNOR U5036 ( .A(in[1238]), .B(n3128), .Z(n3868) );
  NANDN U5037 ( .A(n3871), .B(n3868), .Z(n3129) );
  XNOR U5038 ( .A(n3444), .B(n3129), .Z(out[378]) );
  XOR U5039 ( .A(in[67]), .B(n4423), .Z(n3447) );
  XOR U5040 ( .A(in[1312]), .B(n4264), .Z(n3875) );
  XNOR U5041 ( .A(in[1239]), .B(n3130), .Z(n3872) );
  NANDN U5042 ( .A(n3875), .B(n3872), .Z(n3131) );
  XNOR U5043 ( .A(n3447), .B(n3131), .Z(out[379]) );
  ANDN U5044 ( .B(n3133), .A(n3132), .Z(n3134) );
  XOR U5045 ( .A(n3135), .B(n3134), .Z(out[37]) );
  XOR U5046 ( .A(in[68]), .B(n4426), .Z(n3450) );
  XOR U5047 ( .A(in[1313]), .B(n4267), .Z(n3879) );
  XNOR U5048 ( .A(in[1240]), .B(n3136), .Z(n3876) );
  NANDN U5049 ( .A(n3879), .B(n3876), .Z(n3137) );
  XNOR U5050 ( .A(n3450), .B(n3137), .Z(out[380]) );
  XOR U5051 ( .A(in[69]), .B(n4429), .Z(n3453) );
  XOR U5052 ( .A(in[1314]), .B(n4270), .Z(n3883) );
  XNOR U5053 ( .A(in[1241]), .B(n3138), .Z(n3880) );
  NANDN U5054 ( .A(n3883), .B(n3880), .Z(n3139) );
  XNOR U5055 ( .A(n3453), .B(n3139), .Z(out[381]) );
  XOR U5056 ( .A(in[70]), .B(n4432), .Z(n3460) );
  XOR U5057 ( .A(in[1315]), .B(n3140), .Z(n3887) );
  XNOR U5058 ( .A(in[1242]), .B(n3141), .Z(n3884) );
  NANDN U5059 ( .A(n3887), .B(n3884), .Z(n3142) );
  XOR U5060 ( .A(n3460), .B(n3142), .Z(out[382]) );
  XOR U5061 ( .A(in[71]), .B(n4443), .Z(n3463) );
  XOR U5062 ( .A(in[1316]), .B(n4276), .Z(n3891) );
  XNOR U5063 ( .A(in[1243]), .B(n3143), .Z(n3888) );
  NANDN U5064 ( .A(n3891), .B(n3888), .Z(n3144) );
  XNOR U5065 ( .A(n3463), .B(n3144), .Z(out[383]) );
  XOR U5066 ( .A(in[497]), .B(n4135), .Z(n3465) );
  XOR U5067 ( .A(in[498]), .B(n4139), .Z(n3467) );
  ANDN U5068 ( .B(n3617), .A(n3145), .Z(n3146) );
  XNOR U5069 ( .A(n3467), .B(n3146), .Z(out[385]) );
  XOR U5070 ( .A(in[499]), .B(n4143), .Z(n3469) );
  ANDN U5071 ( .B(n3621), .A(n3147), .Z(n3148) );
  XNOR U5072 ( .A(n3469), .B(n3148), .Z(out[386]) );
  XOR U5073 ( .A(in[500]), .B(n4147), .Z(n3471) );
  ANDN U5074 ( .B(n3625), .A(n3149), .Z(n3150) );
  XNOR U5075 ( .A(n3471), .B(n3150), .Z(out[387]) );
  XOR U5076 ( .A(in[501]), .B(n4151), .Z(n3473) );
  XOR U5077 ( .A(in[502]), .B(n4161), .Z(n3474) );
  NOR U5078 ( .A(n3152), .B(n3151), .Z(n3153) );
  XOR U5079 ( .A(n3154), .B(n3153), .Z(out[38]) );
  XOR U5080 ( .A(in[503]), .B(n4165), .Z(n3475) );
  XOR U5081 ( .A(in[504]), .B(n4169), .Z(n3476) );
  XOR U5082 ( .A(in[505]), .B(n4173), .Z(n3481) );
  XOR U5083 ( .A(in[506]), .B(n3897), .Z(n3482) );
  NOR U5084 ( .A(n3653), .B(n3290), .Z(n3155) );
  XNOR U5085 ( .A(n3482), .B(n3155), .Z(out[393]) );
  XOR U5086 ( .A(in[507]), .B(n3901), .Z(n3484) );
  NOR U5087 ( .A(n3657), .B(n3293), .Z(n3156) );
  XNOR U5088 ( .A(n3484), .B(n3156), .Z(out[394]) );
  XOR U5089 ( .A(in[508]), .B(n3905), .Z(n3486) );
  NOR U5090 ( .A(n3661), .B(n3296), .Z(n3157) );
  XNOR U5091 ( .A(n3486), .B(n3157), .Z(out[395]) );
  XOR U5092 ( .A(in[509]), .B(n3909), .Z(n3488) );
  NOR U5093 ( .A(n3665), .B(n3303), .Z(n3158) );
  XNOR U5094 ( .A(n3488), .B(n3158), .Z(out[396]) );
  XOR U5095 ( .A(in[510]), .B(n3913), .Z(n3490) );
  NOR U5096 ( .A(n3669), .B(n3306), .Z(n3159) );
  XNOR U5097 ( .A(n3490), .B(n3159), .Z(out[397]) );
  XOR U5098 ( .A(in[511]), .B(n3917), .Z(n3492) );
  NOR U5099 ( .A(n3677), .B(n3309), .Z(n3160) );
  XNOR U5100 ( .A(n3492), .B(n3160), .Z(out[398]) );
  XOR U5101 ( .A(in[448]), .B(n3921), .Z(n3494) );
  NOR U5102 ( .A(n3681), .B(n3312), .Z(n3161) );
  XNOR U5103 ( .A(n3494), .B(n3161), .Z(out[399]) );
  ANDN U5104 ( .B(n3163), .A(n3162), .Z(n3164) );
  XOR U5105 ( .A(n3165), .B(n3164), .Z(out[39]) );
  OR U5106 ( .A(n4067), .B(n3166), .Z(n3167) );
  XNOR U5107 ( .A(n4066), .B(n3167), .Z(out[3]) );
  XOR U5108 ( .A(in[449]), .B(n3925), .Z(n3496) );
  NOR U5109 ( .A(n3685), .B(n3315), .Z(n3168) );
  XNOR U5110 ( .A(n3496), .B(n3168), .Z(out[400]) );
  XOR U5111 ( .A(n3169), .B(in[450]), .Z(n3498) );
  NOR U5112 ( .A(n3689), .B(n3318), .Z(n3170) );
  XOR U5113 ( .A(n3498), .B(n3170), .Z(out[401]) );
  XOR U5114 ( .A(n3171), .B(in[451]), .Z(n3503) );
  NOR U5115 ( .A(n3693), .B(n3320), .Z(n3172) );
  XOR U5116 ( .A(n3503), .B(n3172), .Z(out[402]) );
  XOR U5117 ( .A(n3173), .B(in[452]), .Z(n3504) );
  NOR U5118 ( .A(n3697), .B(n3322), .Z(n3174) );
  XOR U5119 ( .A(n3504), .B(n3174), .Z(out[403]) );
  XOR U5120 ( .A(n3175), .B(in[453]), .Z(n3505) );
  NOR U5121 ( .A(n3701), .B(n3324), .Z(n3176) );
  XOR U5122 ( .A(n3505), .B(n3176), .Z(out[404]) );
  XOR U5123 ( .A(n3177), .B(in[454]), .Z(n3506) );
  NOR U5124 ( .A(n3705), .B(n3326), .Z(n3178) );
  XOR U5125 ( .A(n3506), .B(n3178), .Z(out[405]) );
  XOR U5126 ( .A(n3179), .B(in[455]), .Z(n3507) );
  NOR U5127 ( .A(n3709), .B(n3332), .Z(n3180) );
  XOR U5128 ( .A(n3507), .B(n3180), .Z(out[406]) );
  XOR U5129 ( .A(n3181), .B(in[456]), .Z(n3508) );
  NOR U5130 ( .A(n3713), .B(n3334), .Z(n3182) );
  XOR U5131 ( .A(n3508), .B(n3182), .Z(out[407]) );
  XOR U5132 ( .A(in[457]), .B(n3183), .Z(n3509) );
  NOR U5133 ( .A(n3723), .B(n3336), .Z(n3184) );
  XOR U5134 ( .A(n3509), .B(n3184), .Z(out[408]) );
  XOR U5135 ( .A(n3185), .B(in[458]), .Z(n3510) );
  NOR U5136 ( .A(n3727), .B(n3338), .Z(n3186) );
  XOR U5137 ( .A(n3510), .B(n3186), .Z(out[409]) );
  ANDN U5138 ( .B(n3188), .A(n3187), .Z(n3189) );
  XNOR U5139 ( .A(n3190), .B(n3189), .Z(out[40]) );
  XOR U5140 ( .A(n3969), .B(in[459]), .Z(n3511) );
  NOR U5141 ( .A(n3731), .B(n3340), .Z(n3191) );
  XNOR U5142 ( .A(n3511), .B(n3191), .Z(out[410]) );
  XOR U5143 ( .A(in[460]), .B(n3192), .Z(n3513) );
  NOR U5144 ( .A(n3735), .B(n3342), .Z(n3193) );
  XOR U5145 ( .A(n3513), .B(n3193), .Z(out[411]) );
  XOR U5146 ( .A(in[461]), .B(n3194), .Z(n3344) );
  NOR U5147 ( .A(n3195), .B(n3739), .Z(n3196) );
  XOR U5148 ( .A(n3344), .B(n3196), .Z(out[412]) );
  XOR U5149 ( .A(in[462]), .B(n3197), .Z(n3348) );
  NOR U5150 ( .A(n3198), .B(n3743), .Z(n3199) );
  XOR U5151 ( .A(n3348), .B(n3199), .Z(out[413]) );
  XOR U5152 ( .A(in[463]), .B(n3200), .Z(n3351) );
  NOR U5153 ( .A(n3201), .B(n3747), .Z(n3202) );
  XOR U5154 ( .A(n3351), .B(n3202), .Z(out[414]) );
  XOR U5155 ( .A(in[464]), .B(n3203), .Z(n3354) );
  NOR U5156 ( .A(n3204), .B(n3751), .Z(n3205) );
  XOR U5157 ( .A(n3354), .B(n3205), .Z(out[415]) );
  XOR U5158 ( .A(in[465]), .B(n3206), .Z(n3361) );
  NOR U5159 ( .A(n3207), .B(n3755), .Z(n3208) );
  XOR U5160 ( .A(n3361), .B(n3208), .Z(out[416]) );
  XOR U5161 ( .A(in[466]), .B(n3209), .Z(n3364) );
  NOR U5162 ( .A(n3210), .B(n3759), .Z(n3211) );
  XOR U5163 ( .A(n3364), .B(n3211), .Z(out[417]) );
  XOR U5164 ( .A(in[467]), .B(n3212), .Z(n3367) );
  NOR U5165 ( .A(n3213), .B(n3767), .Z(n3214) );
  XOR U5166 ( .A(n3367), .B(n3214), .Z(out[418]) );
  XOR U5167 ( .A(in[468]), .B(n3215), .Z(n3370) );
  NOR U5168 ( .A(n3216), .B(n3771), .Z(n3217) );
  XOR U5169 ( .A(n3370), .B(n3217), .Z(out[419]) );
  AND U5170 ( .A(n3219), .B(n3218), .Z(n3220) );
  XNOR U5171 ( .A(n3221), .B(n3220), .Z(out[41]) );
  XOR U5172 ( .A(in[469]), .B(n4012), .Z(n3538) );
  NOR U5173 ( .A(n3222), .B(n3775), .Z(n3223) );
  XNOR U5174 ( .A(n3538), .B(n3223), .Z(out[420]) );
  XOR U5175 ( .A(in[470]), .B(n4016), .Z(n3540) );
  NOR U5176 ( .A(n3224), .B(n3779), .Z(n3225) );
  XNOR U5177 ( .A(n3540), .B(n3225), .Z(out[421]) );
  XOR U5178 ( .A(in[471]), .B(n4020), .Z(n3547) );
  NOR U5179 ( .A(n3226), .B(n3783), .Z(n3227) );
  XNOR U5180 ( .A(n3547), .B(n3227), .Z(out[422]) );
  XOR U5181 ( .A(in[472]), .B(n4028), .Z(n3550) );
  NOR U5182 ( .A(n3228), .B(n3787), .Z(n3229) );
  XNOR U5183 ( .A(n3550), .B(n3229), .Z(out[423]) );
  XOR U5184 ( .A(in[473]), .B(n4032), .Z(n3553) );
  ANDN U5185 ( .B(n3791), .A(n3230), .Z(n3231) );
  XNOR U5186 ( .A(n3553), .B(n3231), .Z(out[424]) );
  XOR U5187 ( .A(in[474]), .B(n4036), .Z(n3556) );
  ANDN U5188 ( .B(n3795), .A(n3232), .Z(n3233) );
  XNOR U5189 ( .A(n3556), .B(n3233), .Z(out[425]) );
  XOR U5190 ( .A(in[475]), .B(n4040), .Z(n3559) );
  ANDN U5191 ( .B(n3799), .A(n3234), .Z(n3235) );
  XNOR U5192 ( .A(n3559), .B(n3235), .Z(out[426]) );
  XOR U5193 ( .A(in[476]), .B(n4044), .Z(n3562) );
  ANDN U5194 ( .B(n3803), .A(n3236), .Z(n3237) );
  XNOR U5195 ( .A(n3562), .B(n3237), .Z(out[427]) );
  XOR U5196 ( .A(in[477]), .B(n4048), .Z(n3564) );
  ANDN U5197 ( .B(n3811), .A(n3238), .Z(n3239) );
  XNOR U5198 ( .A(n3564), .B(n3239), .Z(out[428]) );
  XOR U5199 ( .A(in[478]), .B(n4052), .Z(n3397) );
  ANDN U5200 ( .B(n3815), .A(n3240), .Z(n3241) );
  XOR U5201 ( .A(n3397), .B(n3241), .Z(out[429]) );
  AND U5202 ( .A(n3243), .B(n3242), .Z(n3244) );
  XNOR U5203 ( .A(n3245), .B(n3244), .Z(out[42]) );
  XOR U5204 ( .A(in[479]), .B(n4056), .Z(n3401) );
  ANDN U5205 ( .B(n3819), .A(n3246), .Z(n3247) );
  XOR U5206 ( .A(n3401), .B(n3247), .Z(out[430]) );
  XOR U5207 ( .A(in[480]), .B(n4060), .Z(n3405) );
  ANDN U5208 ( .B(n3823), .A(n3248), .Z(n3249) );
  XOR U5209 ( .A(n3405), .B(n3249), .Z(out[431]) );
  XOR U5210 ( .A(in[481]), .B(n4064), .Z(n3408) );
  ANDN U5211 ( .B(n3827), .A(n3250), .Z(n3251) );
  XOR U5212 ( .A(n3408), .B(n3251), .Z(out[432]) );
  XOR U5213 ( .A(in[482]), .B(n4072), .Z(n3411) );
  ANDN U5214 ( .B(n3831), .A(n3252), .Z(n3253) );
  XOR U5215 ( .A(n3411), .B(n3253), .Z(out[433]) );
  XOR U5216 ( .A(in[483]), .B(n4076), .Z(n3414) );
  XOR U5217 ( .A(in[484]), .B(n4080), .Z(n3417) );
  XOR U5218 ( .A(in[485]), .B(n4084), .Z(n3584) );
  XOR U5219 ( .A(in[486]), .B(n4087), .Z(n3586) );
  XOR U5220 ( .A(in[487]), .B(n4091), .Z(n3588) );
  XOR U5221 ( .A(in[488]), .B(n4095), .Z(n3590) );
  AND U5222 ( .A(n3255), .B(n3254), .Z(n3256) );
  XNOR U5223 ( .A(n3257), .B(n3256), .Z(out[43]) );
  XOR U5224 ( .A(in[489]), .B(n4099), .Z(n3592) );
  XOR U5225 ( .A(in[490]), .B(n4103), .Z(n3594) );
  XOR U5226 ( .A(in[491]), .B(n4107), .Z(n3600) );
  XOR U5227 ( .A(in[492]), .B(n4115), .Z(n3601) );
  XOR U5228 ( .A(in[493]), .B(n4119), .Z(n3602) );
  XOR U5229 ( .A(in[494]), .B(n4123), .Z(n3604) );
  XOR U5230 ( .A(in[495]), .B(n4127), .Z(n3606) );
  XOR U5231 ( .A(in[496]), .B(n4131), .Z(n3608) );
  XOR U5232 ( .A(in[886]), .B(n3258), .Z(n3611) );
  NAND U5233 ( .A(n3259), .B(n3465), .Z(n3260) );
  XOR U5234 ( .A(n3611), .B(n3260), .Z(out[448]) );
  XOR U5235 ( .A(in[887]), .B(n3261), .Z(n3615) );
  NANDN U5236 ( .A(n3262), .B(n3467), .Z(n3263) );
  XOR U5237 ( .A(n3615), .B(n3263), .Z(out[449]) );
  AND U5238 ( .A(n3265), .B(n3264), .Z(n3266) );
  XNOR U5239 ( .A(n3267), .B(n3266), .Z(out[44]) );
  XOR U5240 ( .A(in[888]), .B(n3268), .Z(n3619) );
  NANDN U5241 ( .A(n3269), .B(n3469), .Z(n3270) );
  XOR U5242 ( .A(n3619), .B(n3270), .Z(out[450]) );
  XOR U5243 ( .A(in[889]), .B(n3271), .Z(n3623) );
  NANDN U5244 ( .A(n3272), .B(n3471), .Z(n3273) );
  XOR U5245 ( .A(n3623), .B(n3273), .Z(out[451]) );
  XOR U5246 ( .A(in[890]), .B(n3274), .Z(n3631) );
  NANDN U5247 ( .A(n3473), .B(n3275), .Z(n3276) );
  XOR U5248 ( .A(n3631), .B(n3276), .Z(out[452]) );
  XOR U5249 ( .A(in[891]), .B(n3277), .Z(n3635) );
  NANDN U5250 ( .A(n3474), .B(n3278), .Z(n3279) );
  XNOR U5251 ( .A(n3635), .B(n3279), .Z(out[453]) );
  XOR U5252 ( .A(in[892]), .B(n3280), .Z(n3639) );
  NANDN U5253 ( .A(n3475), .B(n3281), .Z(n3282) );
  XNOR U5254 ( .A(n3639), .B(n3282), .Z(out[454]) );
  XOR U5255 ( .A(in[893]), .B(n3283), .Z(n3643) );
  NANDN U5256 ( .A(n3476), .B(n3284), .Z(n3285) );
  XNOR U5257 ( .A(n3643), .B(n3285), .Z(out[455]) );
  XOR U5258 ( .A(in[894]), .B(n3286), .Z(n3647) );
  NANDN U5259 ( .A(n3481), .B(n3287), .Z(n3288) );
  XOR U5260 ( .A(n3647), .B(n3288), .Z(out[456]) );
  IV U5261 ( .A(n3289), .Z(n3898) );
  XOR U5262 ( .A(in[895]), .B(n3898), .Z(n3650) );
  NAND U5263 ( .A(n3290), .B(n3482), .Z(n3291) );
  XNOR U5264 ( .A(n3650), .B(n3291), .Z(out[457]) );
  IV U5265 ( .A(n3292), .Z(n3902) );
  XOR U5266 ( .A(in[832]), .B(n3902), .Z(n3654) );
  NAND U5267 ( .A(n3293), .B(n3484), .Z(n3294) );
  XNOR U5268 ( .A(n3654), .B(n3294), .Z(out[458]) );
  IV U5269 ( .A(n3295), .Z(n3906) );
  XOR U5270 ( .A(in[833]), .B(n3906), .Z(n3658) );
  NAND U5271 ( .A(n3296), .B(n3486), .Z(n3297) );
  XNOR U5272 ( .A(n3658), .B(n3297), .Z(out[459]) );
  AND U5273 ( .A(n3299), .B(n3298), .Z(n3300) );
  XNOR U5274 ( .A(n3301), .B(n3300), .Z(out[45]) );
  IV U5275 ( .A(n3302), .Z(n3910) );
  XOR U5276 ( .A(in[834]), .B(n3910), .Z(n3662) );
  NAND U5277 ( .A(n3303), .B(n3488), .Z(n3304) );
  XNOR U5278 ( .A(n3662), .B(n3304), .Z(out[460]) );
  IV U5279 ( .A(n3305), .Z(n3914) );
  XOR U5280 ( .A(in[835]), .B(n3914), .Z(n3666) );
  NAND U5281 ( .A(n3306), .B(n3490), .Z(n3307) );
  XNOR U5282 ( .A(n3666), .B(n3307), .Z(out[461]) );
  IV U5283 ( .A(n3308), .Z(n3918) );
  XOR U5284 ( .A(in[836]), .B(n3918), .Z(n3674) );
  NAND U5285 ( .A(n3309), .B(n3492), .Z(n3310) );
  XNOR U5286 ( .A(n3674), .B(n3310), .Z(out[462]) );
  IV U5287 ( .A(n3311), .Z(n3922) );
  XOR U5288 ( .A(in[837]), .B(n3922), .Z(n3678) );
  NAND U5289 ( .A(n3312), .B(n3494), .Z(n3313) );
  XNOR U5290 ( .A(n3678), .B(n3313), .Z(out[463]) );
  IV U5291 ( .A(n3314), .Z(n3926) );
  XOR U5292 ( .A(in[838]), .B(n3926), .Z(n3682) );
  NAND U5293 ( .A(n3315), .B(n3496), .Z(n3316) );
  XNOR U5294 ( .A(n3682), .B(n3316), .Z(out[464]) );
  XNOR U5295 ( .A(in[839]), .B(n3317), .Z(n3686) );
  NANDN U5296 ( .A(n3498), .B(n3318), .Z(n3319) );
  XNOR U5297 ( .A(n3686), .B(n3319), .Z(out[465]) );
  XNOR U5298 ( .A(in[840]), .B(n3933), .Z(n3690) );
  NANDN U5299 ( .A(n3503), .B(n3320), .Z(n3321) );
  XNOR U5300 ( .A(n3690), .B(n3321), .Z(out[466]) );
  XNOR U5301 ( .A(in[841]), .B(n3940), .Z(n3694) );
  NANDN U5302 ( .A(n3504), .B(n3322), .Z(n3323) );
  XNOR U5303 ( .A(n3694), .B(n3323), .Z(out[467]) );
  XNOR U5304 ( .A(in[842]), .B(n3944), .Z(n3698) );
  NANDN U5305 ( .A(n3505), .B(n3324), .Z(n3325) );
  XNOR U5306 ( .A(n3698), .B(n3325), .Z(out[468]) );
  XNOR U5307 ( .A(in[843]), .B(n3948), .Z(n3702) );
  NANDN U5308 ( .A(n3506), .B(n3326), .Z(n3327) );
  XNOR U5309 ( .A(n3702), .B(n3327), .Z(out[469]) );
  AND U5310 ( .A(n3329), .B(n3328), .Z(n3330) );
  XNOR U5311 ( .A(n3331), .B(n3330), .Z(out[46]) );
  XNOR U5312 ( .A(in[844]), .B(n3952), .Z(n3706) );
  NANDN U5313 ( .A(n3507), .B(n3332), .Z(n3333) );
  XNOR U5314 ( .A(n3706), .B(n3333), .Z(out[470]) );
  XNOR U5315 ( .A(in[845]), .B(n3956), .Z(n3710) );
  NANDN U5316 ( .A(n3508), .B(n3334), .Z(n3335) );
  XNOR U5317 ( .A(n3710), .B(n3335), .Z(out[471]) );
  XNOR U5318 ( .A(in[846]), .B(n3960), .Z(n3720) );
  NANDN U5319 ( .A(n3509), .B(n3336), .Z(n3337) );
  XNOR U5320 ( .A(n3720), .B(n3337), .Z(out[472]) );
  XNOR U5321 ( .A(in[847]), .B(n3964), .Z(n3724) );
  NANDN U5322 ( .A(n3510), .B(n3338), .Z(n3339) );
  XNOR U5323 ( .A(n3724), .B(n3339), .Z(out[473]) );
  XNOR U5324 ( .A(in[848]), .B(n3968), .Z(n3728) );
  NAND U5325 ( .A(n3340), .B(n3511), .Z(n3341) );
  XNOR U5326 ( .A(n3728), .B(n3341), .Z(out[474]) );
  XNOR U5327 ( .A(in[849]), .B(n3972), .Z(n3732) );
  NANDN U5328 ( .A(n3513), .B(n3342), .Z(n3343) );
  XNOR U5329 ( .A(n3732), .B(n3343), .Z(out[475]) );
  XNOR U5330 ( .A(in[850]), .B(n3976), .Z(n3736) );
  IV U5331 ( .A(n3344), .Z(n3518) );
  NANDN U5332 ( .A(n3345), .B(n3518), .Z(n3346) );
  XNOR U5333 ( .A(n3736), .B(n3346), .Z(out[476]) );
  XOR U5334 ( .A(in[851]), .B(n3347), .Z(n3740) );
  IV U5335 ( .A(n3348), .Z(n3520) );
  NANDN U5336 ( .A(n3349), .B(n3520), .Z(n3350) );
  XOR U5337 ( .A(n3740), .B(n3350), .Z(out[477]) );
  XOR U5338 ( .A(in[852]), .B(n3987), .Z(n3522) );
  IV U5339 ( .A(n3351), .Z(n3523) );
  NANDN U5340 ( .A(n3352), .B(n3523), .Z(n3353) );
  XNOR U5341 ( .A(n3522), .B(n3353), .Z(out[478]) );
  XOR U5342 ( .A(in[853]), .B(n3991), .Z(n3748) );
  IV U5343 ( .A(n3354), .Z(n3525) );
  NANDN U5344 ( .A(n3355), .B(n3525), .Z(n3356) );
  XOR U5345 ( .A(n3748), .B(n3356), .Z(out[479]) );
  ANDN U5346 ( .B(n3358), .A(n3357), .Z(n3359) );
  XNOR U5347 ( .A(n3360), .B(n3359), .Z(out[47]) );
  XOR U5348 ( .A(in[854]), .B(n3995), .Z(n3752) );
  IV U5349 ( .A(n3361), .Z(n3527) );
  NANDN U5350 ( .A(n3362), .B(n3527), .Z(n3363) );
  XOR U5351 ( .A(n3752), .B(n3363), .Z(out[480]) );
  XOR U5352 ( .A(in[855]), .B(n3999), .Z(n3529) );
  IV U5353 ( .A(n3364), .Z(n3530) );
  NANDN U5354 ( .A(n3365), .B(n3530), .Z(n3366) );
  XNOR U5355 ( .A(n3529), .B(n3366), .Z(out[481]) );
  XOR U5356 ( .A(in[856]), .B(n4003), .Z(n3532) );
  IV U5357 ( .A(n3367), .Z(n3533) );
  NANDN U5358 ( .A(n3368), .B(n3533), .Z(n3369) );
  XNOR U5359 ( .A(n3532), .B(n3369), .Z(out[482]) );
  XOR U5360 ( .A(in[857]), .B(n4007), .Z(n3535) );
  IV U5361 ( .A(n3370), .Z(n3536) );
  NANDN U5362 ( .A(n3371), .B(n3536), .Z(n3372) );
  XNOR U5363 ( .A(n3535), .B(n3372), .Z(out[483]) );
  XOR U5364 ( .A(in[858]), .B(n4011), .Z(n3772) );
  NANDN U5365 ( .A(n3373), .B(n3538), .Z(n3374) );
  XOR U5366 ( .A(n3772), .B(n3374), .Z(out[484]) );
  XOR U5367 ( .A(in[859]), .B(n4015), .Z(n3776) );
  NANDN U5368 ( .A(n3375), .B(n3540), .Z(n3376) );
  XOR U5369 ( .A(n3776), .B(n3376), .Z(out[485]) );
  XOR U5370 ( .A(in[860]), .B(n4019), .Z(n3546) );
  NANDN U5371 ( .A(n3377), .B(n3547), .Z(n3378) );
  XNOR U5372 ( .A(n3546), .B(n3378), .Z(out[486]) );
  XOR U5373 ( .A(in[861]), .B(n4027), .Z(n3549) );
  NANDN U5374 ( .A(n3379), .B(n3550), .Z(n3380) );
  XNOR U5375 ( .A(n3549), .B(n3380), .Z(out[487]) );
  XOR U5376 ( .A(in[862]), .B(n4031), .Z(n3552) );
  NANDN U5377 ( .A(n3381), .B(n3553), .Z(n3382) );
  XNOR U5378 ( .A(n3552), .B(n3382), .Z(out[488]) );
  XOR U5379 ( .A(in[863]), .B(n4035), .Z(n3555) );
  NANDN U5380 ( .A(n3383), .B(n3556), .Z(n3384) );
  XNOR U5381 ( .A(n3555), .B(n3384), .Z(out[489]) );
  AND U5382 ( .A(n3386), .B(n3385), .Z(n3387) );
  XNOR U5383 ( .A(n3388), .B(n3387), .Z(out[48]) );
  XOR U5384 ( .A(in[864]), .B(n4039), .Z(n3558) );
  NANDN U5385 ( .A(n3389), .B(n3559), .Z(n3390) );
  XNOR U5386 ( .A(n3558), .B(n3390), .Z(out[490]) );
  XOR U5387 ( .A(in[865]), .B(n4043), .Z(n3561) );
  NANDN U5388 ( .A(n3391), .B(n3562), .Z(n3392) );
  XNOR U5389 ( .A(n3561), .B(n3392), .Z(out[491]) );
  XNOR U5390 ( .A(n3393), .B(in[866]), .Z(n3809) );
  NANDN U5391 ( .A(n3394), .B(n3564), .Z(n3395) );
  XNOR U5392 ( .A(n3809), .B(n3395), .Z(out[492]) );
  XNOR U5393 ( .A(n3396), .B(in[867]), .Z(n3813) );
  IV U5394 ( .A(n3397), .Z(n3566) );
  NANDN U5395 ( .A(n3398), .B(n3566), .Z(n3399) );
  XNOR U5396 ( .A(n3813), .B(n3399), .Z(out[493]) );
  XNOR U5397 ( .A(n3400), .B(in[868]), .Z(n3817) );
  IV U5398 ( .A(n3401), .Z(n3568) );
  NANDN U5399 ( .A(n3402), .B(n3568), .Z(n3403) );
  XNOR U5400 ( .A(n3817), .B(n3403), .Z(out[494]) );
  XNOR U5401 ( .A(n3404), .B(in[869]), .Z(n3821) );
  IV U5402 ( .A(n3405), .Z(n3570) );
  NANDN U5403 ( .A(n3406), .B(n3570), .Z(n3407) );
  XNOR U5404 ( .A(n3821), .B(n3407), .Z(out[495]) );
  XOR U5405 ( .A(in[870]), .B(n4063), .Z(n3825) );
  IV U5406 ( .A(n3408), .Z(n3576) );
  NANDN U5407 ( .A(n3409), .B(n3576), .Z(n3410) );
  XOR U5408 ( .A(n3825), .B(n3410), .Z(out[496]) );
  XOR U5409 ( .A(in[871]), .B(n4071), .Z(n3829) );
  IV U5410 ( .A(n3411), .Z(n3578) );
  NANDN U5411 ( .A(n3412), .B(n3578), .Z(n3413) );
  XOR U5412 ( .A(n3829), .B(n3413), .Z(out[497]) );
  XOR U5413 ( .A(in[872]), .B(n4075), .Z(n3833) );
  IV U5414 ( .A(n3414), .Z(n3580) );
  NANDN U5415 ( .A(n3415), .B(n3580), .Z(n3416) );
  XOR U5416 ( .A(n3833), .B(n3416), .Z(out[498]) );
  XOR U5417 ( .A(in[873]), .B(n4079), .Z(n3837) );
  IV U5418 ( .A(n3417), .Z(n3582) );
  NANDN U5419 ( .A(n3418), .B(n3582), .Z(n3419) );
  XOR U5420 ( .A(n3837), .B(n3419), .Z(out[499]) );
  ANDN U5421 ( .B(n3421), .A(n3420), .Z(n3422) );
  XNOR U5422 ( .A(n3423), .B(n3422), .Z(out[49]) );
  OR U5423 ( .A(n4111), .B(n3424), .Z(n3425) );
  XNOR U5424 ( .A(n4110), .B(n3425), .Z(out[4]) );
  XOR U5425 ( .A(in[874]), .B(n4083), .Z(n3841) );
  NAND U5426 ( .A(n3426), .B(n3584), .Z(n3427) );
  XOR U5427 ( .A(n3841), .B(n3427), .Z(out[500]) );
  XOR U5428 ( .A(in[875]), .B(n3428), .Z(n3845) );
  NAND U5429 ( .A(n3429), .B(n3586), .Z(n3430) );
  XOR U5430 ( .A(n3845), .B(n3430), .Z(out[501]) );
  XOR U5431 ( .A(in[876]), .B(n3431), .Z(n3853) );
  NAND U5432 ( .A(n3432), .B(n3588), .Z(n3433) );
  XOR U5433 ( .A(n3853), .B(n3433), .Z(out[502]) );
  XOR U5434 ( .A(in[877]), .B(n3434), .Z(n3857) );
  NAND U5435 ( .A(n3435), .B(n3590), .Z(n3436) );
  XOR U5436 ( .A(n3857), .B(n3436), .Z(out[503]) );
  XOR U5437 ( .A(in[878]), .B(n3437), .Z(n3861) );
  NAND U5438 ( .A(n3438), .B(n3592), .Z(n3439) );
  XOR U5439 ( .A(n3861), .B(n3439), .Z(out[504]) );
  XOR U5440 ( .A(in[879]), .B(n3440), .Z(n3865) );
  NAND U5441 ( .A(n3441), .B(n3594), .Z(n3442) );
  XOR U5442 ( .A(n3865), .B(n3442), .Z(out[505]) );
  XOR U5443 ( .A(in[880]), .B(n3443), .Z(n3869) );
  NANDN U5444 ( .A(n3600), .B(n3444), .Z(n3445) );
  XOR U5445 ( .A(n3869), .B(n3445), .Z(out[506]) );
  XOR U5446 ( .A(in[881]), .B(n3446), .Z(n3873) );
  NANDN U5447 ( .A(n3601), .B(n3447), .Z(n3448) );
  XOR U5448 ( .A(n3873), .B(n3448), .Z(out[507]) );
  XOR U5449 ( .A(in[882]), .B(n3449), .Z(n3877) );
  NAND U5450 ( .A(n3450), .B(n3602), .Z(n3451) );
  XOR U5451 ( .A(n3877), .B(n3451), .Z(out[508]) );
  XOR U5452 ( .A(in[883]), .B(n3452), .Z(n3881) );
  NAND U5453 ( .A(n3453), .B(n3604), .Z(n3454) );
  XOR U5454 ( .A(n3881), .B(n3454), .Z(out[509]) );
  ANDN U5455 ( .B(n3456), .A(n3455), .Z(n3457) );
  XNOR U5456 ( .A(n3458), .B(n3457), .Z(out[50]) );
  XOR U5457 ( .A(in[884]), .B(n3459), .Z(n3885) );
  NANDN U5458 ( .A(n3460), .B(n3606), .Z(n3461) );
  XOR U5459 ( .A(n3885), .B(n3461), .Z(out[510]) );
  XOR U5460 ( .A(in[885]), .B(n3462), .Z(n3889) );
  NAND U5461 ( .A(n3463), .B(n3608), .Z(n3464) );
  XOR U5462 ( .A(n3889), .B(n3464), .Z(out[511]) );
  NANDN U5463 ( .A(n3465), .B(n3611), .Z(n3466) );
  XNOR U5464 ( .A(n3610), .B(n3466), .Z(out[512]) );
  NANDN U5465 ( .A(n3467), .B(n3615), .Z(n3468) );
  XNOR U5466 ( .A(n3614), .B(n3468), .Z(out[513]) );
  NANDN U5467 ( .A(n3469), .B(n3619), .Z(n3470) );
  XNOR U5468 ( .A(n3618), .B(n3470), .Z(out[514]) );
  NANDN U5469 ( .A(n3471), .B(n3623), .Z(n3472) );
  XNOR U5470 ( .A(n3622), .B(n3472), .Z(out[515]) );
  ANDN U5471 ( .B(n3478), .A(n3477), .Z(n3479) );
  XNOR U5472 ( .A(n3480), .B(n3479), .Z(out[51]) );
  OR U5473 ( .A(n3650), .B(n3482), .Z(n3483) );
  XOR U5474 ( .A(n3651), .B(n3483), .Z(out[521]) );
  OR U5475 ( .A(n3654), .B(n3484), .Z(n3485) );
  XOR U5476 ( .A(n3655), .B(n3485), .Z(out[522]) );
  OR U5477 ( .A(n3658), .B(n3486), .Z(n3487) );
  XOR U5478 ( .A(n3659), .B(n3487), .Z(out[523]) );
  OR U5479 ( .A(n3662), .B(n3488), .Z(n3489) );
  XOR U5480 ( .A(n3663), .B(n3489), .Z(out[524]) );
  OR U5481 ( .A(n3666), .B(n3490), .Z(n3491) );
  XOR U5482 ( .A(n3667), .B(n3491), .Z(out[525]) );
  OR U5483 ( .A(n3674), .B(n3492), .Z(n3493) );
  XOR U5484 ( .A(n3675), .B(n3493), .Z(out[526]) );
  OR U5485 ( .A(n3678), .B(n3494), .Z(n3495) );
  XOR U5486 ( .A(n3679), .B(n3495), .Z(out[527]) );
  OR U5487 ( .A(n3682), .B(n3496), .Z(n3497) );
  XOR U5488 ( .A(n3683), .B(n3497), .Z(out[528]) );
  ANDN U5489 ( .B(n3500), .A(n3499), .Z(n3501) );
  XNOR U5490 ( .A(n3502), .B(n3501), .Z(out[52]) );
  OR U5491 ( .A(n3728), .B(n3511), .Z(n3512) );
  XOR U5492 ( .A(n3729), .B(n3512), .Z(out[538]) );
  ANDN U5493 ( .B(n3515), .A(n3514), .Z(n3516) );
  XNOR U5494 ( .A(n3517), .B(n3516), .Z(out[53]) );
  OR U5495 ( .A(n3736), .B(n3518), .Z(n3519) );
  XOR U5496 ( .A(n3737), .B(n3519), .Z(out[540]) );
  NANDN U5497 ( .A(n3520), .B(n3740), .Z(n3521) );
  XOR U5498 ( .A(n3741), .B(n3521), .Z(out[541]) );
  IV U5499 ( .A(n3522), .Z(n3744) );
  NANDN U5500 ( .A(n3523), .B(n3744), .Z(n3524) );
  XOR U5501 ( .A(n3745), .B(n3524), .Z(out[542]) );
  NANDN U5502 ( .A(n3525), .B(n3748), .Z(n3526) );
  XOR U5503 ( .A(n3749), .B(n3526), .Z(out[543]) );
  NANDN U5504 ( .A(n3527), .B(n3752), .Z(n3528) );
  XOR U5505 ( .A(n3753), .B(n3528), .Z(out[544]) );
  IV U5506 ( .A(n3529), .Z(n3756) );
  NANDN U5507 ( .A(n3530), .B(n3756), .Z(n3531) );
  XOR U5508 ( .A(n3757), .B(n3531), .Z(out[545]) );
  IV U5509 ( .A(n3532), .Z(n3764) );
  NANDN U5510 ( .A(n3533), .B(n3764), .Z(n3534) );
  XOR U5511 ( .A(n3765), .B(n3534), .Z(out[546]) );
  IV U5512 ( .A(n3535), .Z(n3768) );
  NANDN U5513 ( .A(n3536), .B(n3768), .Z(n3537) );
  XOR U5514 ( .A(n3769), .B(n3537), .Z(out[547]) );
  NANDN U5515 ( .A(n3538), .B(n3772), .Z(n3539) );
  XOR U5516 ( .A(n3773), .B(n3539), .Z(out[548]) );
  NANDN U5517 ( .A(n3540), .B(n3776), .Z(n3541) );
  XOR U5518 ( .A(n3777), .B(n3541), .Z(out[549]) );
  ANDN U5519 ( .B(n3543), .A(n3542), .Z(n3544) );
  XNOR U5520 ( .A(n3545), .B(n3544), .Z(out[54]) );
  IV U5521 ( .A(n3546), .Z(n3780) );
  NANDN U5522 ( .A(n3547), .B(n3780), .Z(n3548) );
  XOR U5523 ( .A(n3781), .B(n3548), .Z(out[550]) );
  IV U5524 ( .A(n3549), .Z(n3784) );
  NANDN U5525 ( .A(n3550), .B(n3784), .Z(n3551) );
  XOR U5526 ( .A(n3785), .B(n3551), .Z(out[551]) );
  IV U5527 ( .A(n3552), .Z(n3789) );
  NANDN U5528 ( .A(n3553), .B(n3789), .Z(n3554) );
  XNOR U5529 ( .A(n3788), .B(n3554), .Z(out[552]) );
  IV U5530 ( .A(n3555), .Z(n3793) );
  NANDN U5531 ( .A(n3556), .B(n3793), .Z(n3557) );
  XNOR U5532 ( .A(n3792), .B(n3557), .Z(out[553]) );
  IV U5533 ( .A(n3558), .Z(n3797) );
  NANDN U5534 ( .A(n3559), .B(n3797), .Z(n3560) );
  XNOR U5535 ( .A(n3796), .B(n3560), .Z(out[554]) );
  IV U5536 ( .A(n3561), .Z(n3801) );
  NANDN U5537 ( .A(n3562), .B(n3801), .Z(n3563) );
  XNOR U5538 ( .A(n3800), .B(n3563), .Z(out[555]) );
  OR U5539 ( .A(n3809), .B(n3564), .Z(n3565) );
  XNOR U5540 ( .A(n3808), .B(n3565), .Z(out[556]) );
  OR U5541 ( .A(n3813), .B(n3566), .Z(n3567) );
  XNOR U5542 ( .A(n3812), .B(n3567), .Z(out[557]) );
  OR U5543 ( .A(n3817), .B(n3568), .Z(n3569) );
  XNOR U5544 ( .A(n3816), .B(n3569), .Z(out[558]) );
  OR U5545 ( .A(n3821), .B(n3570), .Z(n3571) );
  XNOR U5546 ( .A(n3820), .B(n3571), .Z(out[559]) );
  ANDN U5547 ( .B(n3573), .A(n3572), .Z(n3574) );
  XNOR U5548 ( .A(n3575), .B(n3574), .Z(out[55]) );
  NANDN U5549 ( .A(n3576), .B(n3825), .Z(n3577) );
  XNOR U5550 ( .A(n3824), .B(n3577), .Z(out[560]) );
  NANDN U5551 ( .A(n3578), .B(n3829), .Z(n3579) );
  XNOR U5552 ( .A(n3828), .B(n3579), .Z(out[561]) );
  NANDN U5553 ( .A(n3580), .B(n3833), .Z(n3581) );
  XNOR U5554 ( .A(n3832), .B(n3581), .Z(out[562]) );
  NANDN U5555 ( .A(n3582), .B(n3837), .Z(n3583) );
  XNOR U5556 ( .A(n3836), .B(n3583), .Z(out[563]) );
  NANDN U5557 ( .A(n3584), .B(n3841), .Z(n3585) );
  XNOR U5558 ( .A(n3840), .B(n3585), .Z(out[564]) );
  NANDN U5559 ( .A(n3586), .B(n3845), .Z(n3587) );
  XNOR U5560 ( .A(n3844), .B(n3587), .Z(out[565]) );
  NANDN U5561 ( .A(n3588), .B(n3853), .Z(n3589) );
  XNOR U5562 ( .A(n3852), .B(n3589), .Z(out[566]) );
  NANDN U5563 ( .A(n3590), .B(n3857), .Z(n3591) );
  XNOR U5564 ( .A(n3856), .B(n3591), .Z(out[567]) );
  NANDN U5565 ( .A(n3592), .B(n3861), .Z(n3593) );
  XNOR U5566 ( .A(n3860), .B(n3593), .Z(out[568]) );
  NANDN U5567 ( .A(n3594), .B(n3865), .Z(n3595) );
  XNOR U5568 ( .A(n3864), .B(n3595), .Z(out[569]) );
  ANDN U5569 ( .B(n3597), .A(n3596), .Z(n3598) );
  XNOR U5570 ( .A(n3599), .B(n3598), .Z(out[56]) );
  NANDN U5571 ( .A(n3602), .B(n3877), .Z(n3603) );
  XNOR U5572 ( .A(n3876), .B(n3603), .Z(out[572]) );
  NANDN U5573 ( .A(n3604), .B(n3881), .Z(n3605) );
  XNOR U5574 ( .A(n3880), .B(n3605), .Z(out[573]) );
  NANDN U5575 ( .A(n3606), .B(n3885), .Z(n3607) );
  XNOR U5576 ( .A(n3884), .B(n3607), .Z(out[574]) );
  NANDN U5577 ( .A(n3608), .B(n3889), .Z(n3609) );
  XNOR U5578 ( .A(n3888), .B(n3609), .Z(out[575]) );
  NOR U5579 ( .A(n3611), .B(n3610), .Z(n3612) );
  XOR U5580 ( .A(n3613), .B(n3612), .Z(out[576]) );
  NOR U5581 ( .A(n3615), .B(n3614), .Z(n3616) );
  XOR U5582 ( .A(n3617), .B(n3616), .Z(out[577]) );
  NOR U5583 ( .A(n3619), .B(n3618), .Z(n3620) );
  XOR U5584 ( .A(n3621), .B(n3620), .Z(out[578]) );
  NOR U5585 ( .A(n3623), .B(n3622), .Z(n3624) );
  XOR U5586 ( .A(n3625), .B(n3624), .Z(out[579]) );
  ANDN U5587 ( .B(n3627), .A(n3626), .Z(n3628) );
  XNOR U5588 ( .A(n3629), .B(n3628), .Z(out[57]) );
  NOR U5589 ( .A(n3631), .B(n3630), .Z(n3632) );
  XOR U5590 ( .A(n3633), .B(n3632), .Z(out[580]) );
  ANDN U5591 ( .B(n3635), .A(n3634), .Z(n3636) );
  XOR U5592 ( .A(n3637), .B(n3636), .Z(out[581]) );
  ANDN U5593 ( .B(n3639), .A(n3638), .Z(n3640) );
  XOR U5594 ( .A(n3641), .B(n3640), .Z(out[582]) );
  ANDN U5595 ( .B(n3643), .A(n3642), .Z(n3644) );
  XOR U5596 ( .A(n3645), .B(n3644), .Z(out[583]) );
  NOR U5597 ( .A(n3647), .B(n3646), .Z(n3648) );
  XOR U5598 ( .A(n3649), .B(n3648), .Z(out[584]) );
  AND U5599 ( .A(n3651), .B(n3650), .Z(n3652) );
  XNOR U5600 ( .A(n3653), .B(n3652), .Z(out[585]) );
  AND U5601 ( .A(n3655), .B(n3654), .Z(n3656) );
  XNOR U5602 ( .A(n3657), .B(n3656), .Z(out[586]) );
  AND U5603 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U5604 ( .A(n3661), .B(n3660), .Z(out[587]) );
  AND U5605 ( .A(n3663), .B(n3662), .Z(n3664) );
  XNOR U5606 ( .A(n3665), .B(n3664), .Z(out[588]) );
  AND U5607 ( .A(n3667), .B(n3666), .Z(n3668) );
  XNOR U5608 ( .A(n3669), .B(n3668), .Z(out[589]) );
  ANDN U5609 ( .B(n3671), .A(n3670), .Z(n3672) );
  XNOR U5610 ( .A(n3673), .B(n3672), .Z(out[58]) );
  AND U5611 ( .A(n3675), .B(n3674), .Z(n3676) );
  XNOR U5612 ( .A(n3677), .B(n3676), .Z(out[590]) );
  AND U5613 ( .A(n3679), .B(n3678), .Z(n3680) );
  XNOR U5614 ( .A(n3681), .B(n3680), .Z(out[591]) );
  AND U5615 ( .A(n3683), .B(n3682), .Z(n3684) );
  XNOR U5616 ( .A(n3685), .B(n3684), .Z(out[592]) );
  AND U5617 ( .A(n3687), .B(n3686), .Z(n3688) );
  XNOR U5618 ( .A(n3689), .B(n3688), .Z(out[593]) );
  AND U5619 ( .A(n3691), .B(n3690), .Z(n3692) );
  XNOR U5620 ( .A(n3693), .B(n3692), .Z(out[594]) );
  AND U5621 ( .A(n3695), .B(n3694), .Z(n3696) );
  XNOR U5622 ( .A(n3697), .B(n3696), .Z(out[595]) );
  AND U5623 ( .A(n3699), .B(n3698), .Z(n3700) );
  XNOR U5624 ( .A(n3701), .B(n3700), .Z(out[596]) );
  AND U5625 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR U5626 ( .A(n3705), .B(n3704), .Z(out[597]) );
  AND U5627 ( .A(n3707), .B(n3706), .Z(n3708) );
  XNOR U5628 ( .A(n3709), .B(n3708), .Z(out[598]) );
  AND U5629 ( .A(n3711), .B(n3710), .Z(n3712) );
  XNOR U5630 ( .A(n3713), .B(n3712), .Z(out[599]) );
  ANDN U5631 ( .B(n3715), .A(n3714), .Z(n3716) );
  XNOR U5632 ( .A(n3717), .B(n3716), .Z(out[59]) );
  OR U5633 ( .A(n4155), .B(n3718), .Z(n3719) );
  XNOR U5634 ( .A(n4154), .B(n3719), .Z(out[5]) );
  AND U5635 ( .A(n3721), .B(n3720), .Z(n3722) );
  XNOR U5636 ( .A(n3723), .B(n3722), .Z(out[600]) );
  AND U5637 ( .A(n3725), .B(n3724), .Z(n3726) );
  XNOR U5638 ( .A(n3727), .B(n3726), .Z(out[601]) );
  AND U5639 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U5640 ( .A(n3731), .B(n3730), .Z(out[602]) );
  AND U5641 ( .A(n3733), .B(n3732), .Z(n3734) );
  XNOR U5642 ( .A(n3735), .B(n3734), .Z(out[603]) );
  AND U5643 ( .A(n3737), .B(n3736), .Z(n3738) );
  XNOR U5644 ( .A(n3739), .B(n3738), .Z(out[604]) );
  ANDN U5645 ( .B(n3741), .A(n3740), .Z(n3742) );
  XNOR U5646 ( .A(n3743), .B(n3742), .Z(out[605]) );
  ANDN U5647 ( .B(n3745), .A(n3744), .Z(n3746) );
  XNOR U5648 ( .A(n3747), .B(n3746), .Z(out[606]) );
  ANDN U5649 ( .B(n3749), .A(n3748), .Z(n3750) );
  XNOR U5650 ( .A(n3751), .B(n3750), .Z(out[607]) );
  ANDN U5651 ( .B(n3753), .A(n3752), .Z(n3754) );
  XNOR U5652 ( .A(n3755), .B(n3754), .Z(out[608]) );
  ANDN U5653 ( .B(n3757), .A(n3756), .Z(n3758) );
  XNOR U5654 ( .A(n3759), .B(n3758), .Z(out[609]) );
  ANDN U5655 ( .B(n3761), .A(n3760), .Z(n3762) );
  XNOR U5656 ( .A(n3763), .B(n3762), .Z(out[60]) );
  ANDN U5657 ( .B(n3765), .A(n3764), .Z(n3766) );
  XNOR U5658 ( .A(n3767), .B(n3766), .Z(out[610]) );
  ANDN U5659 ( .B(n3769), .A(n3768), .Z(n3770) );
  XNOR U5660 ( .A(n3771), .B(n3770), .Z(out[611]) );
  ANDN U5661 ( .B(n3773), .A(n3772), .Z(n3774) );
  XNOR U5662 ( .A(n3775), .B(n3774), .Z(out[612]) );
  ANDN U5663 ( .B(n3777), .A(n3776), .Z(n3778) );
  XNOR U5664 ( .A(n3779), .B(n3778), .Z(out[613]) );
  ANDN U5665 ( .B(n3781), .A(n3780), .Z(n3782) );
  XNOR U5666 ( .A(n3783), .B(n3782), .Z(out[614]) );
  ANDN U5667 ( .B(n3785), .A(n3784), .Z(n3786) );
  XNOR U5668 ( .A(n3787), .B(n3786), .Z(out[615]) );
  NOR U5669 ( .A(n3789), .B(n3788), .Z(n3790) );
  XOR U5670 ( .A(n3791), .B(n3790), .Z(out[616]) );
  NOR U5671 ( .A(n3793), .B(n3792), .Z(n3794) );
  XOR U5672 ( .A(n3795), .B(n3794), .Z(out[617]) );
  NOR U5673 ( .A(n3797), .B(n3796), .Z(n3798) );
  XOR U5674 ( .A(n3799), .B(n3798), .Z(out[618]) );
  NOR U5675 ( .A(n3801), .B(n3800), .Z(n3802) );
  XOR U5676 ( .A(n3803), .B(n3802), .Z(out[619]) );
  ANDN U5677 ( .B(n3805), .A(n3804), .Z(n3806) );
  XOR U5678 ( .A(n3807), .B(n3806), .Z(out[61]) );
  ANDN U5679 ( .B(n3809), .A(n3808), .Z(n3810) );
  XOR U5680 ( .A(n3811), .B(n3810), .Z(out[620]) );
  ANDN U5681 ( .B(n3813), .A(n3812), .Z(n3814) );
  XOR U5682 ( .A(n3815), .B(n3814), .Z(out[621]) );
  ANDN U5683 ( .B(n3817), .A(n3816), .Z(n3818) );
  XOR U5684 ( .A(n3819), .B(n3818), .Z(out[622]) );
  ANDN U5685 ( .B(n3821), .A(n3820), .Z(n3822) );
  XOR U5686 ( .A(n3823), .B(n3822), .Z(out[623]) );
  NOR U5687 ( .A(n3825), .B(n3824), .Z(n3826) );
  XOR U5688 ( .A(n3827), .B(n3826), .Z(out[624]) );
  NOR U5689 ( .A(n3829), .B(n3828), .Z(n3830) );
  XOR U5690 ( .A(n3831), .B(n3830), .Z(out[625]) );
  NOR U5691 ( .A(n3833), .B(n3832), .Z(n3834) );
  XOR U5692 ( .A(n3835), .B(n3834), .Z(out[626]) );
  NOR U5693 ( .A(n3837), .B(n3836), .Z(n3838) );
  XOR U5694 ( .A(n3839), .B(n3838), .Z(out[627]) );
  NOR U5695 ( .A(n3841), .B(n3840), .Z(n3842) );
  XOR U5696 ( .A(n3843), .B(n3842), .Z(out[628]) );
  NOR U5697 ( .A(n3845), .B(n3844), .Z(n3846) );
  XOR U5698 ( .A(n3847), .B(n3846), .Z(out[629]) );
  ANDN U5699 ( .B(n3849), .A(n3848), .Z(n3850) );
  XOR U5700 ( .A(n3851), .B(n3850), .Z(out[62]) );
  NOR U5701 ( .A(n3853), .B(n3852), .Z(n3854) );
  XOR U5702 ( .A(n3855), .B(n3854), .Z(out[630]) );
  NOR U5703 ( .A(n3857), .B(n3856), .Z(n3858) );
  XOR U5704 ( .A(n3859), .B(n3858), .Z(out[631]) );
  NOR U5705 ( .A(n3861), .B(n3860), .Z(n3862) );
  XOR U5706 ( .A(n3863), .B(n3862), .Z(out[632]) );
  NOR U5707 ( .A(n3865), .B(n3864), .Z(n3866) );
  XOR U5708 ( .A(n3867), .B(n3866), .Z(out[633]) );
  NOR U5709 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U5710 ( .A(n3871), .B(n3870), .Z(out[634]) );
  NOR U5711 ( .A(n3873), .B(n3872), .Z(n3874) );
  XOR U5712 ( .A(n3875), .B(n3874), .Z(out[635]) );
  NOR U5713 ( .A(n3877), .B(n3876), .Z(n3878) );
  XOR U5714 ( .A(n3879), .B(n3878), .Z(out[636]) );
  NOR U5715 ( .A(n3881), .B(n3880), .Z(n3882) );
  XOR U5716 ( .A(n3883), .B(n3882), .Z(out[637]) );
  NOR U5717 ( .A(n3885), .B(n3884), .Z(n3886) );
  XOR U5718 ( .A(n3887), .B(n3886), .Z(out[638]) );
  NOR U5719 ( .A(n3889), .B(n3888), .Z(n3890) );
  XOR U5720 ( .A(n3891), .B(n3890), .Z(out[639]) );
  ANDN U5721 ( .B(n3893), .A(n3892), .Z(n3894) );
  XOR U5722 ( .A(n3895), .B(n3894), .Z(out[63]) );
  XOR U5723 ( .A(in[302]), .B(n3896), .Z(n4177) );
  IV U5724 ( .A(n4177), .Z(n4334) );
  XOR U5725 ( .A(in[1146]), .B(n3897), .Z(n4711) );
  XOR U5726 ( .A(in[1535]), .B(n3898), .Z(n4713) );
  OR U5727 ( .A(n4711), .B(n4713), .Z(n3899) );
  XOR U5728 ( .A(n4334), .B(n3899), .Z(out[640]) );
  XOR U5729 ( .A(in[303]), .B(n3900), .Z(n4180) );
  IV U5730 ( .A(n4180), .Z(n4336) );
  XOR U5731 ( .A(in[1147]), .B(n3901), .Z(n4715) );
  XOR U5732 ( .A(in[1472]), .B(n3902), .Z(n4717) );
  OR U5733 ( .A(n4715), .B(n4717), .Z(n3903) );
  XOR U5734 ( .A(n4336), .B(n3903), .Z(out[641]) );
  XOR U5735 ( .A(in[304]), .B(n3904), .Z(n4183) );
  IV U5736 ( .A(n4183), .Z(n4342) );
  XOR U5737 ( .A(in[1148]), .B(n3905), .Z(n4719) );
  XOR U5738 ( .A(in[1473]), .B(n3906), .Z(n4721) );
  OR U5739 ( .A(n4719), .B(n4721), .Z(n3907) );
  XOR U5740 ( .A(n4342), .B(n3907), .Z(out[642]) );
  XOR U5741 ( .A(in[305]), .B(n3908), .Z(n4186) );
  IV U5742 ( .A(n4186), .Z(n4344) );
  XOR U5743 ( .A(in[1149]), .B(n3909), .Z(n4723) );
  XOR U5744 ( .A(in[1474]), .B(n3910), .Z(n4725) );
  OR U5745 ( .A(n4723), .B(n4725), .Z(n3911) );
  XOR U5746 ( .A(n4344), .B(n3911), .Z(out[643]) );
  XOR U5747 ( .A(in[306]), .B(n3912), .Z(n4189) );
  IV U5748 ( .A(n4189), .Z(n4346) );
  XOR U5749 ( .A(in[1150]), .B(n3913), .Z(n4735) );
  XOR U5750 ( .A(in[1475]), .B(n3914), .Z(n4737) );
  OR U5751 ( .A(n4735), .B(n4737), .Z(n3915) );
  XOR U5752 ( .A(n4346), .B(n3915), .Z(out[644]) );
  XOR U5753 ( .A(in[307]), .B(n3916), .Z(n4349) );
  XOR U5754 ( .A(in[1151]), .B(n3917), .Z(n4739) );
  XOR U5755 ( .A(in[1476]), .B(n3918), .Z(n4741) );
  OR U5756 ( .A(n4739), .B(n4741), .Z(n3919) );
  XOR U5757 ( .A(n4349), .B(n3919), .Z(out[645]) );
  XOR U5758 ( .A(in[308]), .B(n3920), .Z(n4352) );
  XOR U5759 ( .A(in[1088]), .B(n3921), .Z(n4743) );
  XOR U5760 ( .A(in[1477]), .B(n3922), .Z(n4745) );
  OR U5761 ( .A(n4743), .B(n4745), .Z(n3923) );
  XOR U5762 ( .A(n4352), .B(n3923), .Z(out[646]) );
  XOR U5763 ( .A(in[309]), .B(n3924), .Z(n4355) );
  XOR U5764 ( .A(in[1089]), .B(n3925), .Z(n4747) );
  XOR U5765 ( .A(in[1478]), .B(n3926), .Z(n4749) );
  OR U5766 ( .A(n4747), .B(n4749), .Z(n3927) );
  XOR U5767 ( .A(n4355), .B(n3927), .Z(out[647]) );
  XOR U5768 ( .A(in[310]), .B(n3928), .Z(n4357) );
  XOR U5769 ( .A(in[1479]), .B(n3929), .Z(n4753) );
  XNOR U5770 ( .A(n3930), .B(in[1090]), .Z(n4750) );
  NANDN U5771 ( .A(n4753), .B(n4750), .Z(n3931) );
  XOR U5772 ( .A(n4357), .B(n3931), .Z(out[648]) );
  XOR U5773 ( .A(in[311]), .B(n3932), .Z(n4360) );
  XNOR U5774 ( .A(n3934), .B(in[1091]), .Z(n4754) );
  NANDN U5775 ( .A(n4757), .B(n4754), .Z(n3935) );
  XOR U5776 ( .A(n4360), .B(n3935), .Z(out[649]) );
  XOR U5777 ( .A(in[312]), .B(n3939), .Z(n4363) );
  XNOR U5778 ( .A(n3941), .B(in[1092]), .Z(n4758) );
  NANDN U5779 ( .A(n4761), .B(n4758), .Z(n3942) );
  XOR U5780 ( .A(n4363), .B(n3942), .Z(out[650]) );
  XOR U5781 ( .A(in[313]), .B(n3943), .Z(n4366) );
  XNOR U5782 ( .A(n3945), .B(in[1093]), .Z(n4762) );
  NANDN U5783 ( .A(n4765), .B(n4762), .Z(n3946) );
  XOR U5784 ( .A(n4366), .B(n3946), .Z(out[651]) );
  XOR U5785 ( .A(in[314]), .B(n3947), .Z(n4373) );
  XNOR U5786 ( .A(n3949), .B(in[1094]), .Z(n4766) );
  NANDN U5787 ( .A(n4769), .B(n4766), .Z(n3950) );
  XOR U5788 ( .A(n4373), .B(n3950), .Z(out[652]) );
  XOR U5789 ( .A(in[315]), .B(n3951), .Z(n4204) );
  IV U5790 ( .A(n4204), .Z(n4376) );
  XNOR U5791 ( .A(n3953), .B(in[1095]), .Z(n4770) );
  NANDN U5792 ( .A(n4773), .B(n4770), .Z(n3954) );
  XOR U5793 ( .A(n4376), .B(n3954), .Z(out[653]) );
  XOR U5794 ( .A(in[316]), .B(n3955), .Z(n4207) );
  IV U5795 ( .A(n4207), .Z(n4379) );
  XNOR U5796 ( .A(n3957), .B(in[1096]), .Z(n4778) );
  NANDN U5797 ( .A(n4781), .B(n4778), .Z(n3958) );
  XOR U5798 ( .A(n4379), .B(n3958), .Z(out[654]) );
  XOR U5799 ( .A(in[317]), .B(n3959), .Z(n4210) );
  IV U5800 ( .A(n4210), .Z(n4382) );
  XNOR U5801 ( .A(in[1097]), .B(n3961), .Z(n4782) );
  NANDN U5802 ( .A(n4785), .B(n4782), .Z(n3962) );
  XOR U5803 ( .A(n4382), .B(n3962), .Z(out[655]) );
  XOR U5804 ( .A(in[318]), .B(n3963), .Z(n4215) );
  IV U5805 ( .A(n4215), .Z(n4385) );
  XNOR U5806 ( .A(n3965), .B(in[1098]), .Z(n4786) );
  NANDN U5807 ( .A(n4789), .B(n4786), .Z(n3966) );
  XOR U5808 ( .A(n4385), .B(n3966), .Z(out[656]) );
  XOR U5809 ( .A(in[319]), .B(n3967), .Z(n4218) );
  IV U5810 ( .A(n4218), .Z(n4387) );
  XNOR U5811 ( .A(n3969), .B(in[1099]), .Z(n4790) );
  NANDN U5812 ( .A(n4793), .B(n4790), .Z(n3970) );
  XOR U5813 ( .A(n4387), .B(n3970), .Z(out[657]) );
  XOR U5814 ( .A(in[256]), .B(n3971), .Z(n4221) );
  IV U5815 ( .A(n4221), .Z(n4390) );
  XNOR U5816 ( .A(in[1100]), .B(n3973), .Z(n4794) );
  NANDN U5817 ( .A(n4797), .B(n4794), .Z(n3974) );
  XOR U5818 ( .A(n4390), .B(n3974), .Z(out[658]) );
  XOR U5819 ( .A(in[257]), .B(n3975), .Z(n4224) );
  IV U5820 ( .A(n4224), .Z(n4393) );
  XNOR U5821 ( .A(in[1101]), .B(n3977), .Z(n4798) );
  NANDN U5822 ( .A(n4801), .B(n4798), .Z(n3978) );
  XOR U5823 ( .A(n4393), .B(n3978), .Z(out[659]) );
  XOR U5824 ( .A(in[258]), .B(n3982), .Z(n4227) );
  IV U5825 ( .A(n4227), .Z(n4396) );
  XOR U5826 ( .A(in[1491]), .B(n3983), .Z(n4805) );
  XNOR U5827 ( .A(in[1102]), .B(n3984), .Z(n4802) );
  NANDN U5828 ( .A(n4805), .B(n4802), .Z(n3985) );
  XOR U5829 ( .A(n4396), .B(n3985), .Z(out[660]) );
  XOR U5830 ( .A(in[259]), .B(n3986), .Z(n4230) );
  IV U5831 ( .A(n4230), .Z(n4399) );
  XOR U5832 ( .A(in[1492]), .B(n3987), .Z(n4809) );
  XNOR U5833 ( .A(in[1103]), .B(n3988), .Z(n4806) );
  NANDN U5834 ( .A(n4809), .B(n4806), .Z(n3989) );
  XOR U5835 ( .A(n4399), .B(n3989), .Z(out[661]) );
  XOR U5836 ( .A(in[260]), .B(n3990), .Z(n4406) );
  XOR U5837 ( .A(in[1493]), .B(n3991), .Z(n4233) );
  IV U5838 ( .A(n4233), .Z(n4813) );
  XNOR U5839 ( .A(in[1104]), .B(n3992), .Z(n4810) );
  NANDN U5840 ( .A(n4813), .B(n4810), .Z(n3993) );
  XNOR U5841 ( .A(n4406), .B(n3993), .Z(out[662]) );
  XOR U5842 ( .A(in[261]), .B(n3994), .Z(n4409) );
  XOR U5843 ( .A(in[1494]), .B(n3995), .Z(n4236) );
  IV U5844 ( .A(n4236), .Z(n4817) );
  XNOR U5845 ( .A(in[1105]), .B(n3996), .Z(n4814) );
  NANDN U5846 ( .A(n4817), .B(n4814), .Z(n3997) );
  XNOR U5847 ( .A(n4409), .B(n3997), .Z(out[663]) );
  XOR U5848 ( .A(in[262]), .B(n3998), .Z(n4412) );
  XOR U5849 ( .A(in[1495]), .B(n3999), .Z(n4825) );
  XNOR U5850 ( .A(in[1106]), .B(n4000), .Z(n4822) );
  NANDN U5851 ( .A(n4825), .B(n4822), .Z(n4001) );
  XNOR U5852 ( .A(n4412), .B(n4001), .Z(out[664]) );
  XOR U5853 ( .A(in[263]), .B(n4002), .Z(n4415) );
  XOR U5854 ( .A(in[1496]), .B(n4003), .Z(n4829) );
  XNOR U5855 ( .A(in[1107]), .B(n4004), .Z(n4826) );
  NANDN U5856 ( .A(n4829), .B(n4826), .Z(n4005) );
  XNOR U5857 ( .A(n4415), .B(n4005), .Z(out[665]) );
  XOR U5858 ( .A(in[264]), .B(n4006), .Z(n4418) );
  XOR U5859 ( .A(in[1497]), .B(n4007), .Z(n4833) );
  XNOR U5860 ( .A(in[1108]), .B(n4008), .Z(n4830) );
  NANDN U5861 ( .A(n4833), .B(n4830), .Z(n4009) );
  XNOR U5862 ( .A(n4418), .B(n4009), .Z(out[666]) );
  XOR U5863 ( .A(in[265]), .B(n4010), .Z(n4421) );
  XOR U5864 ( .A(in[1498]), .B(n4011), .Z(n4244) );
  IV U5865 ( .A(n4244), .Z(n4837) );
  XNOR U5866 ( .A(in[1109]), .B(n4012), .Z(n4834) );
  NANDN U5867 ( .A(n4837), .B(n4834), .Z(n4013) );
  XNOR U5868 ( .A(n4421), .B(n4013), .Z(out[667]) );
  XOR U5869 ( .A(in[266]), .B(n4014), .Z(n4424) );
  XOR U5870 ( .A(in[1499]), .B(n4015), .Z(n4247) );
  IV U5871 ( .A(n4247), .Z(n4841) );
  XNOR U5872 ( .A(in[1110]), .B(n4016), .Z(n4838) );
  NANDN U5873 ( .A(n4841), .B(n4838), .Z(n4017) );
  XNOR U5874 ( .A(n4424), .B(n4017), .Z(out[668]) );
  XOR U5875 ( .A(in[267]), .B(n4018), .Z(n4427) );
  XOR U5876 ( .A(in[1500]), .B(n4019), .Z(n4845) );
  XNOR U5877 ( .A(in[1111]), .B(n4020), .Z(n4842) );
  NANDN U5878 ( .A(n4845), .B(n4842), .Z(n4021) );
  XNOR U5879 ( .A(n4427), .B(n4021), .Z(out[669]) );
  ANDN U5880 ( .B(n4023), .A(n4022), .Z(n4024) );
  XOR U5881 ( .A(n4025), .B(n4024), .Z(out[66]) );
  XOR U5882 ( .A(in[268]), .B(n4026), .Z(n4430) );
  XOR U5883 ( .A(in[1501]), .B(n4027), .Z(n4849) );
  XNOR U5884 ( .A(in[1112]), .B(n4028), .Z(n4846) );
  NANDN U5885 ( .A(n4849), .B(n4846), .Z(n4029) );
  XNOR U5886 ( .A(n4430), .B(n4029), .Z(out[670]) );
  XOR U5887 ( .A(in[269]), .B(n4030), .Z(n4433) );
  XOR U5888 ( .A(in[1502]), .B(n4031), .Z(n4853) );
  XNOR U5889 ( .A(in[1113]), .B(n4032), .Z(n4850) );
  NANDN U5890 ( .A(n4853), .B(n4850), .Z(n4033) );
  XNOR U5891 ( .A(n4433), .B(n4033), .Z(out[671]) );
  XOR U5892 ( .A(in[270]), .B(n4034), .Z(n4444) );
  XOR U5893 ( .A(in[1503]), .B(n4035), .Z(n4857) );
  XNOR U5894 ( .A(in[1114]), .B(n4036), .Z(n4854) );
  NANDN U5895 ( .A(n4857), .B(n4854), .Z(n4037) );
  XNOR U5896 ( .A(n4444), .B(n4037), .Z(out[672]) );
  XOR U5897 ( .A(in[271]), .B(n4038), .Z(n4447) );
  XOR U5898 ( .A(in[1504]), .B(n4039), .Z(n4861) );
  XNOR U5899 ( .A(in[1115]), .B(n4040), .Z(n4858) );
  NANDN U5900 ( .A(n4861), .B(n4858), .Z(n4041) );
  XNOR U5901 ( .A(n4447), .B(n4041), .Z(out[673]) );
  XOR U5902 ( .A(in[272]), .B(n4042), .Z(n4450) );
  XOR U5903 ( .A(in[1505]), .B(n4043), .Z(n4869) );
  XNOR U5904 ( .A(in[1116]), .B(n4044), .Z(n4866) );
  NANDN U5905 ( .A(n4869), .B(n4866), .Z(n4045) );
  XNOR U5906 ( .A(n4450), .B(n4045), .Z(out[674]) );
  XNOR U5907 ( .A(in[273]), .B(n4046), .Z(n4453) );
  XOR U5908 ( .A(n4047), .B(in[1506]), .Z(n4873) );
  XNOR U5909 ( .A(in[1117]), .B(n4048), .Z(n4870) );
  NANDN U5910 ( .A(n4873), .B(n4870), .Z(n4049) );
  XNOR U5911 ( .A(n4453), .B(n4049), .Z(out[675]) );
  XOR U5912 ( .A(in[274]), .B(n4050), .Z(n4456) );
  XOR U5913 ( .A(n4051), .B(in[1507]), .Z(n4877) );
  XOR U5914 ( .A(in[1118]), .B(n4052), .Z(n4874) );
  NANDN U5915 ( .A(n4877), .B(n4874), .Z(n4053) );
  XNOR U5916 ( .A(n4456), .B(n4053), .Z(out[676]) );
  XOR U5917 ( .A(in[275]), .B(n4054), .Z(n4459) );
  XOR U5918 ( .A(n4055), .B(in[1508]), .Z(n4881) );
  XOR U5919 ( .A(in[1119]), .B(n4056), .Z(n4878) );
  NANDN U5920 ( .A(n4881), .B(n4878), .Z(n4057) );
  XNOR U5921 ( .A(n4459), .B(n4057), .Z(out[677]) );
  XOR U5922 ( .A(in[276]), .B(n4058), .Z(n4462) );
  XOR U5923 ( .A(n4059), .B(in[1509]), .Z(n4885) );
  XOR U5924 ( .A(in[1120]), .B(n4060), .Z(n4882) );
  NANDN U5925 ( .A(n4885), .B(n4882), .Z(n4061) );
  XNOR U5926 ( .A(n4462), .B(n4061), .Z(out[678]) );
  XOR U5927 ( .A(in[277]), .B(n4062), .Z(n4465) );
  XOR U5928 ( .A(in[1510]), .B(n4063), .Z(n4262) );
  IV U5929 ( .A(n4262), .Z(n4889) );
  XOR U5930 ( .A(in[1121]), .B(n4064), .Z(n4886) );
  NANDN U5931 ( .A(n4889), .B(n4886), .Z(n4065) );
  XNOR U5932 ( .A(n4465), .B(n4065), .Z(out[679]) );
  ANDN U5933 ( .B(n4067), .A(n4066), .Z(n4068) );
  XOR U5934 ( .A(n4069), .B(n4068), .Z(out[67]) );
  XOR U5935 ( .A(in[278]), .B(n4070), .Z(n4468) );
  XOR U5936 ( .A(in[1511]), .B(n4071), .Z(n4265) );
  IV U5937 ( .A(n4265), .Z(n4893) );
  XOR U5938 ( .A(in[1122]), .B(n4072), .Z(n4890) );
  NANDN U5939 ( .A(n4893), .B(n4890), .Z(n4073) );
  XNOR U5940 ( .A(n4468), .B(n4073), .Z(out[680]) );
  XOR U5941 ( .A(in[279]), .B(n4074), .Z(n4471) );
  XOR U5942 ( .A(in[1512]), .B(n4075), .Z(n4268) );
  IV U5943 ( .A(n4268), .Z(n4897) );
  XOR U5944 ( .A(in[1123]), .B(n4076), .Z(n4894) );
  NANDN U5945 ( .A(n4897), .B(n4894), .Z(n4077) );
  XNOR U5946 ( .A(n4471), .B(n4077), .Z(out[681]) );
  XOR U5947 ( .A(in[280]), .B(n4078), .Z(n4478) );
  XOR U5948 ( .A(in[1513]), .B(n4079), .Z(n4271) );
  IV U5949 ( .A(n4271), .Z(n4901) );
  XOR U5950 ( .A(in[1124]), .B(n4080), .Z(n4898) );
  NANDN U5951 ( .A(n4901), .B(n4898), .Z(n4081) );
  XNOR U5952 ( .A(n4478), .B(n4081), .Z(out[682]) );
  XOR U5953 ( .A(in[281]), .B(n4082), .Z(n4481) );
  XOR U5954 ( .A(in[1514]), .B(n4083), .Z(n4274) );
  IV U5955 ( .A(n4274), .Z(n4905) );
  XNOR U5956 ( .A(in[1125]), .B(n4084), .Z(n4902) );
  NANDN U5957 ( .A(n4905), .B(n4902), .Z(n4085) );
  XNOR U5958 ( .A(n4481), .B(n4085), .Z(out[683]) );
  XOR U5959 ( .A(in[282]), .B(n4086), .Z(n4484) );
  XOR U5960 ( .A(in[1126]), .B(n4087), .Z(n4911) );
  XNOR U5961 ( .A(in[1515]), .B(n4088), .Z(n4913) );
  NANDN U5962 ( .A(n4911), .B(n4913), .Z(n4089) );
  XNOR U5963 ( .A(n4484), .B(n4089), .Z(out[684]) );
  XOR U5964 ( .A(in[283]), .B(n4090), .Z(n4487) );
  XOR U5965 ( .A(in[1127]), .B(n4091), .Z(n4915) );
  XNOR U5966 ( .A(in[1516]), .B(n4092), .Z(n4917) );
  NANDN U5967 ( .A(n4915), .B(n4917), .Z(n4093) );
  XNOR U5968 ( .A(n4487), .B(n4093), .Z(out[685]) );
  XOR U5969 ( .A(in[284]), .B(n4094), .Z(n4490) );
  XOR U5970 ( .A(in[1128]), .B(n4095), .Z(n4919) );
  XNOR U5971 ( .A(in[1517]), .B(n4096), .Z(n4921) );
  NANDN U5972 ( .A(n4919), .B(n4921), .Z(n4097) );
  XNOR U5973 ( .A(n4490), .B(n4097), .Z(out[686]) );
  XOR U5974 ( .A(in[285]), .B(n4098), .Z(n4493) );
  XOR U5975 ( .A(in[1129]), .B(n4099), .Z(n4923) );
  XNOR U5976 ( .A(in[1518]), .B(n4100), .Z(n4925) );
  NANDN U5977 ( .A(n4923), .B(n4925), .Z(n4101) );
  XNOR U5978 ( .A(n4493), .B(n4101), .Z(out[687]) );
  XOR U5979 ( .A(in[286]), .B(n4102), .Z(n4496) );
  XOR U5980 ( .A(in[1130]), .B(n4103), .Z(n4927) );
  XNOR U5981 ( .A(in[1519]), .B(n4104), .Z(n4929) );
  NANDN U5982 ( .A(n4927), .B(n4929), .Z(n4105) );
  XNOR U5983 ( .A(n4496), .B(n4105), .Z(out[688]) );
  XOR U5984 ( .A(in[287]), .B(n4106), .Z(n4499) );
  XNOR U5985 ( .A(in[1131]), .B(n4107), .Z(n4931) );
  XNOR U5986 ( .A(in[1520]), .B(n4108), .Z(n4933) );
  NANDN U5987 ( .A(n4931), .B(n4933), .Z(n4109) );
  XNOR U5988 ( .A(n4499), .B(n4109), .Z(out[689]) );
  ANDN U5989 ( .B(n4111), .A(n4110), .Z(n4112) );
  XOR U5990 ( .A(n4113), .B(n4112), .Z(out[68]) );
  XOR U5991 ( .A(in[288]), .B(n4114), .Z(n4502) );
  XNOR U5992 ( .A(in[1132]), .B(n4115), .Z(n4935) );
  XNOR U5993 ( .A(in[1521]), .B(n4116), .Z(n4937) );
  NANDN U5994 ( .A(n4935), .B(n4937), .Z(n4117) );
  XNOR U5995 ( .A(n4502), .B(n4117), .Z(out[690]) );
  XOR U5996 ( .A(in[289]), .B(n4118), .Z(n4505) );
  XOR U5997 ( .A(in[1133]), .B(n4119), .Z(n4939) );
  XNOR U5998 ( .A(in[1522]), .B(n4120), .Z(n4941) );
  NANDN U5999 ( .A(n4939), .B(n4941), .Z(n4121) );
  XNOR U6000 ( .A(n4505), .B(n4121), .Z(out[691]) );
  XNOR U6001 ( .A(in[290]), .B(n4122), .Z(n4512) );
  XOR U6002 ( .A(in[1134]), .B(n4123), .Z(n4943) );
  XNOR U6003 ( .A(in[1523]), .B(n4124), .Z(n4945) );
  NANDN U6004 ( .A(n4943), .B(n4945), .Z(n4125) );
  XNOR U6005 ( .A(n4512), .B(n4125), .Z(out[692]) );
  XOR U6006 ( .A(in[291]), .B(n4126), .Z(n4515) );
  XOR U6007 ( .A(in[1135]), .B(n4127), .Z(n4947) );
  XNOR U6008 ( .A(in[1524]), .B(n4128), .Z(n4949) );
  NANDN U6009 ( .A(n4947), .B(n4949), .Z(n4129) );
  XNOR U6010 ( .A(n4515), .B(n4129), .Z(out[693]) );
  XOR U6011 ( .A(in[292]), .B(n4130), .Z(n4518) );
  XOR U6012 ( .A(in[1136]), .B(n4131), .Z(n4955) );
  XNOR U6013 ( .A(in[1525]), .B(n4132), .Z(n4957) );
  NANDN U6014 ( .A(n4955), .B(n4957), .Z(n4133) );
  XNOR U6015 ( .A(n4518), .B(n4133), .Z(out[694]) );
  XOR U6016 ( .A(in[293]), .B(n4134), .Z(n4303) );
  IV U6017 ( .A(n4303), .Z(n4522) );
  XOR U6018 ( .A(in[1137]), .B(n4135), .Z(n4959) );
  XNOR U6019 ( .A(in[1526]), .B(n4136), .Z(n4961) );
  NANDN U6020 ( .A(n4959), .B(n4961), .Z(n4137) );
  XOR U6021 ( .A(n4522), .B(n4137), .Z(out[695]) );
  XOR U6022 ( .A(in[294]), .B(n4138), .Z(n4310) );
  IV U6023 ( .A(n4310), .Z(n4526) );
  XOR U6024 ( .A(in[1138]), .B(n4139), .Z(n4963) );
  XNOR U6025 ( .A(in[1527]), .B(n4140), .Z(n4965) );
  NANDN U6026 ( .A(n4963), .B(n4965), .Z(n4141) );
  XOR U6027 ( .A(n4526), .B(n4141), .Z(out[696]) );
  XOR U6028 ( .A(in[295]), .B(n4142), .Z(n4313) );
  IV U6029 ( .A(n4313), .Z(n4530) );
  XOR U6030 ( .A(in[1139]), .B(n4143), .Z(n4967) );
  XNOR U6031 ( .A(in[1528]), .B(n4144), .Z(n4969) );
  NANDN U6032 ( .A(n4967), .B(n4969), .Z(n4145) );
  XOR U6033 ( .A(n4530), .B(n4145), .Z(out[697]) );
  XOR U6034 ( .A(in[296]), .B(n4146), .Z(n4316) );
  IV U6035 ( .A(n4316), .Z(n4534) );
  XOR U6036 ( .A(in[1140]), .B(n4147), .Z(n4971) );
  XNOR U6037 ( .A(in[1529]), .B(n4148), .Z(n4973) );
  NANDN U6038 ( .A(n4971), .B(n4973), .Z(n4149) );
  XOR U6039 ( .A(n4534), .B(n4149), .Z(out[698]) );
  XOR U6040 ( .A(in[297]), .B(n4150), .Z(n4319) );
  IV U6041 ( .A(n4319), .Z(n4538) );
  XNOR U6042 ( .A(in[1141]), .B(n4151), .Z(n4975) );
  XNOR U6043 ( .A(in[1530]), .B(n4152), .Z(n4977) );
  NANDN U6044 ( .A(n4975), .B(n4977), .Z(n4153) );
  XOR U6045 ( .A(n4538), .B(n4153), .Z(out[699]) );
  ANDN U6046 ( .B(n4155), .A(n4154), .Z(n4156) );
  XOR U6047 ( .A(n4157), .B(n4156), .Z(out[69]) );
  OR U6048 ( .A(n4193), .B(n4158), .Z(n4159) );
  XNOR U6049 ( .A(n4192), .B(n4159), .Z(out[6]) );
  XOR U6050 ( .A(in[298]), .B(n4160), .Z(n4322) );
  IV U6051 ( .A(n4322), .Z(n4542) );
  XNOR U6052 ( .A(in[1142]), .B(n4161), .Z(n4979) );
  XNOR U6053 ( .A(in[1531]), .B(n4162), .Z(n4981) );
  OR U6054 ( .A(n4979), .B(n4981), .Z(n4163) );
  XOR U6055 ( .A(n4542), .B(n4163), .Z(out[700]) );
  XOR U6056 ( .A(in[299]), .B(n4164), .Z(n4325) );
  IV U6057 ( .A(n4325), .Z(n4545) );
  XNOR U6058 ( .A(in[1143]), .B(n4165), .Z(n4983) );
  XNOR U6059 ( .A(in[1532]), .B(n4166), .Z(n4985) );
  OR U6060 ( .A(n4983), .B(n4985), .Z(n4167) );
  XOR U6061 ( .A(n4545), .B(n4167), .Z(out[701]) );
  XOR U6062 ( .A(in[300]), .B(n4168), .Z(n4328) );
  IV U6063 ( .A(n4328), .Z(n4551) );
  XNOR U6064 ( .A(in[1144]), .B(n4169), .Z(n4987) );
  XNOR U6065 ( .A(in[1533]), .B(n4170), .Z(n4989) );
  OR U6066 ( .A(n4987), .B(n4989), .Z(n4171) );
  XOR U6067 ( .A(n4551), .B(n4171), .Z(out[702]) );
  XOR U6068 ( .A(in[301]), .B(n4172), .Z(n4331) );
  IV U6069 ( .A(n4331), .Z(n4553) );
  XNOR U6070 ( .A(in[1145]), .B(n4173), .Z(n4991) );
  XNOR U6071 ( .A(in[1534]), .B(n4174), .Z(n4993) );
  NANDN U6072 ( .A(n4991), .B(n4993), .Z(n4175) );
  XOR U6073 ( .A(n4553), .B(n4175), .Z(out[703]) );
  XOR U6074 ( .A(in[376]), .B(n4176), .Z(n4554) );
  ANDN U6075 ( .B(n4713), .A(n4177), .Z(n4178) );
  XOR U6076 ( .A(n4554), .B(n4178), .Z(out[704]) );
  XOR U6077 ( .A(in[377]), .B(n4179), .Z(n4557) );
  ANDN U6078 ( .B(n4717), .A(n4180), .Z(n4181) );
  XOR U6079 ( .A(n4557), .B(n4181), .Z(out[705]) );
  XOR U6080 ( .A(in[378]), .B(n4182), .Z(n4560) );
  ANDN U6081 ( .B(n4721), .A(n4183), .Z(n4184) );
  XOR U6082 ( .A(n4560), .B(n4184), .Z(out[706]) );
  XOR U6083 ( .A(in[379]), .B(n4185), .Z(n4563) );
  ANDN U6084 ( .B(n4725), .A(n4186), .Z(n4187) );
  XOR U6085 ( .A(n4563), .B(n4187), .Z(out[707]) );
  XOR U6086 ( .A(in[380]), .B(n4188), .Z(n4566) );
  ANDN U6087 ( .B(n4737), .A(n4189), .Z(n4190) );
  XNOR U6088 ( .A(n4566), .B(n4190), .Z(out[708]) );
  XOR U6089 ( .A(in[381]), .B(n4191), .Z(n4568) );
  ANDN U6090 ( .B(n4193), .A(n4192), .Z(n4194) );
  XOR U6091 ( .A(n4195), .B(n4194), .Z(out[70]) );
  XOR U6092 ( .A(in[382]), .B(n4196), .Z(n4570) );
  XOR U6093 ( .A(in[383]), .B(n4197), .Z(n4572) );
  XOR U6094 ( .A(in[320]), .B(n4198), .Z(n4579) );
  XOR U6095 ( .A(in[321]), .B(n4199), .Z(n4581) );
  XOR U6096 ( .A(in[322]), .B(n4200), .Z(n4583) );
  XOR U6097 ( .A(in[323]), .B(n4201), .Z(n4585) );
  XOR U6098 ( .A(in[324]), .B(n4202), .Z(n4587) );
  XOR U6099 ( .A(in[325]), .B(n4203), .Z(n4589) );
  ANDN U6100 ( .B(n4773), .A(n4204), .Z(n4205) );
  XNOR U6101 ( .A(n4589), .B(n4205), .Z(out[717]) );
  XOR U6102 ( .A(in[326]), .B(n4206), .Z(n4591) );
  ANDN U6103 ( .B(n4781), .A(n4207), .Z(n4208) );
  XNOR U6104 ( .A(n4591), .B(n4208), .Z(out[718]) );
  XOR U6105 ( .A(in[327]), .B(n4209), .Z(n4593) );
  ANDN U6106 ( .B(n4785), .A(n4210), .Z(n4211) );
  XNOR U6107 ( .A(n4593), .B(n4211), .Z(out[719]) );
  ANDN U6108 ( .B(n4440), .A(n4442), .Z(n4212) );
  XOR U6109 ( .A(n4213), .B(n4212), .Z(out[71]) );
  XOR U6110 ( .A(in[328]), .B(n4214), .Z(n4595) );
  ANDN U6111 ( .B(n4789), .A(n4215), .Z(n4216) );
  XOR U6112 ( .A(n4595), .B(n4216), .Z(out[720]) );
  XOR U6113 ( .A(in[329]), .B(n4217), .Z(n4598) );
  ANDN U6114 ( .B(n4793), .A(n4218), .Z(n4219) );
  XNOR U6115 ( .A(n4598), .B(n4219), .Z(out[721]) );
  XOR U6116 ( .A(in[330]), .B(n4220), .Z(n4604) );
  ANDN U6117 ( .B(n4797), .A(n4221), .Z(n4222) );
  XNOR U6118 ( .A(n4604), .B(n4222), .Z(out[722]) );
  XOR U6119 ( .A(in[331]), .B(n4223), .Z(n4606) );
  ANDN U6120 ( .B(n4801), .A(n4224), .Z(n4225) );
  XNOR U6121 ( .A(n4606), .B(n4225), .Z(out[723]) );
  XOR U6122 ( .A(in[332]), .B(n4226), .Z(n4608) );
  ANDN U6123 ( .B(n4805), .A(n4227), .Z(n4228) );
  XNOR U6124 ( .A(n4608), .B(n4228), .Z(out[724]) );
  XOR U6125 ( .A(in[333]), .B(n4229), .Z(n4610) );
  ANDN U6126 ( .B(n4809), .A(n4230), .Z(n4231) );
  XNOR U6127 ( .A(n4610), .B(n4231), .Z(out[725]) );
  XOR U6128 ( .A(in[334]), .B(n4232), .Z(n4612) );
  NOR U6129 ( .A(n4233), .B(n4406), .Z(n4234) );
  XOR U6130 ( .A(n4612), .B(n4234), .Z(out[726]) );
  XOR U6131 ( .A(in[335]), .B(n4235), .Z(n4615) );
  NOR U6132 ( .A(n4236), .B(n4409), .Z(n4237) );
  XOR U6133 ( .A(n4615), .B(n4237), .Z(out[727]) );
  XOR U6134 ( .A(in[336]), .B(n4238), .Z(n4618) );
  XOR U6135 ( .A(in[337]), .B(n4239), .Z(n4621) );
  ANDN U6136 ( .B(n4731), .A(n4733), .Z(n4240) );
  XOR U6137 ( .A(n4241), .B(n4240), .Z(out[72]) );
  XOR U6138 ( .A(in[338]), .B(n4242), .Z(n4624) );
  XOR U6139 ( .A(in[339]), .B(n4243), .Z(n4626) );
  NOR U6140 ( .A(n4244), .B(n4421), .Z(n4245) );
  XNOR U6141 ( .A(n4626), .B(n4245), .Z(out[731]) );
  XOR U6142 ( .A(in[340]), .B(n4246), .Z(n4631) );
  NOR U6143 ( .A(n4247), .B(n4424), .Z(n4248) );
  XOR U6144 ( .A(n4631), .B(n4248), .Z(out[732]) );
  XOR U6145 ( .A(in[341]), .B(n4249), .Z(n4634) );
  XOR U6146 ( .A(in[342]), .B(n4250), .Z(n4637) );
  XOR U6147 ( .A(in[343]), .B(n4251), .Z(n4640) );
  XOR U6148 ( .A(in[344]), .B(n4252), .Z(n4641) );
  XOR U6149 ( .A(in[345]), .B(n4253), .Z(n4644) );
  XOR U6150 ( .A(in[346]), .B(n4254), .Z(n4647) );
  XOR U6151 ( .A(in[347]), .B(n4255), .Z(n4650) );
  ANDN U6152 ( .B(n5162), .A(n5164), .Z(n4256) );
  XOR U6153 ( .A(n4257), .B(n4256), .Z(out[73]) );
  XOR U6154 ( .A(in[348]), .B(n4258), .Z(n4653) );
  XOR U6155 ( .A(in[349]), .B(n4259), .Z(n4656) );
  XOR U6156 ( .A(in[350]), .B(n4260), .Z(n4663) );
  XOR U6157 ( .A(in[351]), .B(n4261), .Z(n4666) );
  NOR U6158 ( .A(n4262), .B(n4465), .Z(n4263) );
  XOR U6159 ( .A(n4666), .B(n4263), .Z(out[743]) );
  XOR U6160 ( .A(in[352]), .B(n4264), .Z(n4667) );
  NOR U6161 ( .A(n4265), .B(n4468), .Z(n4266) );
  XOR U6162 ( .A(n4667), .B(n4266), .Z(out[744]) );
  XOR U6163 ( .A(in[353]), .B(n4267), .Z(n4668) );
  NOR U6164 ( .A(n4268), .B(n4471), .Z(n4269) );
  XOR U6165 ( .A(n4668), .B(n4269), .Z(out[745]) );
  XOR U6166 ( .A(in[354]), .B(n4270), .Z(n4669) );
  NOR U6167 ( .A(n4271), .B(n4478), .Z(n4272) );
  XOR U6168 ( .A(n4669), .B(n4272), .Z(out[746]) );
  XOR U6169 ( .A(in[355]), .B(n4273), .Z(n4670) );
  NOR U6170 ( .A(n4274), .B(n4481), .Z(n4275) );
  XNOR U6171 ( .A(n4670), .B(n4275), .Z(out[747]) );
  XOR U6172 ( .A(in[356]), .B(n4276), .Z(n4672) );
  NOR U6173 ( .A(n4913), .B(n4484), .Z(n4277) );
  XOR U6174 ( .A(n4672), .B(n4277), .Z(out[748]) );
  XOR U6175 ( .A(in[357]), .B(n4278), .Z(n4673) );
  NOR U6176 ( .A(n4917), .B(n4487), .Z(n4279) );
  XOR U6177 ( .A(n4673), .B(n4279), .Z(out[749]) );
  ANDN U6178 ( .B(n4281), .A(n4280), .Z(n4282) );
  XOR U6179 ( .A(n4283), .B(n4282), .Z(out[74]) );
  XOR U6180 ( .A(in[358]), .B(n4284), .Z(n4674) );
  NOR U6181 ( .A(n4921), .B(n4490), .Z(n4285) );
  XOR U6182 ( .A(n4674), .B(n4285), .Z(out[750]) );
  XOR U6183 ( .A(in[359]), .B(n4286), .Z(n4675) );
  NOR U6184 ( .A(n4925), .B(n4493), .Z(n4287) );
  XOR U6185 ( .A(n4675), .B(n4287), .Z(out[751]) );
  XOR U6186 ( .A(in[360]), .B(n4288), .Z(n4679) );
  NOR U6187 ( .A(n4929), .B(n4496), .Z(n4289) );
  XOR U6188 ( .A(n4679), .B(n4289), .Z(out[752]) );
  XOR U6189 ( .A(in[361]), .B(n4290), .Z(n4680) );
  NOR U6190 ( .A(n4933), .B(n4499), .Z(n4291) );
  XOR U6191 ( .A(n4680), .B(n4291), .Z(out[753]) );
  XOR U6192 ( .A(in[362]), .B(n4292), .Z(n4681) );
  NOR U6193 ( .A(n4937), .B(n4502), .Z(n4293) );
  XOR U6194 ( .A(n4681), .B(n4293), .Z(out[754]) );
  XOR U6195 ( .A(in[363]), .B(n4294), .Z(n4682) );
  NOR U6196 ( .A(n4941), .B(n4505), .Z(n4295) );
  XOR U6197 ( .A(n4682), .B(n4295), .Z(out[755]) );
  XOR U6198 ( .A(in[364]), .B(n4296), .Z(n4683) );
  NOR U6199 ( .A(n4945), .B(n4512), .Z(n4297) );
  XOR U6200 ( .A(n4683), .B(n4297), .Z(out[756]) );
  XOR U6201 ( .A(in[365]), .B(n4298), .Z(n4684) );
  NOR U6202 ( .A(n4949), .B(n4515), .Z(n4299) );
  XOR U6203 ( .A(n4684), .B(n4299), .Z(out[757]) );
  XOR U6204 ( .A(in[366]), .B(n4300), .Z(n4685) );
  NOR U6205 ( .A(n4957), .B(n4518), .Z(n4301) );
  XOR U6206 ( .A(n4685), .B(n4301), .Z(out[758]) );
  XOR U6207 ( .A(in[367]), .B(n4302), .Z(n4521) );
  NOR U6208 ( .A(n4303), .B(n4961), .Z(n4304) );
  XOR U6209 ( .A(n4521), .B(n4304), .Z(out[759]) );
  ANDN U6210 ( .B(n4306), .A(n4305), .Z(n4307) );
  XOR U6211 ( .A(n4308), .B(n4307), .Z(out[75]) );
  XOR U6212 ( .A(in[368]), .B(n4309), .Z(n4525) );
  NOR U6213 ( .A(n4310), .B(n4965), .Z(n4311) );
  XOR U6214 ( .A(n4525), .B(n4311), .Z(out[760]) );
  XOR U6215 ( .A(in[369]), .B(n4312), .Z(n4529) );
  NOR U6216 ( .A(n4313), .B(n4969), .Z(n4314) );
  XOR U6217 ( .A(n4529), .B(n4314), .Z(out[761]) );
  XOR U6218 ( .A(in[370]), .B(n4315), .Z(n4533) );
  NOR U6219 ( .A(n4316), .B(n4973), .Z(n4317) );
  XOR U6220 ( .A(n4533), .B(n4317), .Z(out[762]) );
  XOR U6221 ( .A(in[371]), .B(n4318), .Z(n4537) );
  NOR U6222 ( .A(n4319), .B(n4977), .Z(n4320) );
  XOR U6223 ( .A(n4537), .B(n4320), .Z(out[763]) );
  XOR U6224 ( .A(in[372]), .B(n4321), .Z(n4541) );
  ANDN U6225 ( .B(n4981), .A(n4322), .Z(n4323) );
  XOR U6226 ( .A(n4541), .B(n4323), .Z(out[764]) );
  XOR U6227 ( .A(in[373]), .B(n4324), .Z(n4701) );
  ANDN U6228 ( .B(n4985), .A(n4325), .Z(n4326) );
  XOR U6229 ( .A(n4701), .B(n4326), .Z(out[765]) );
  XOR U6230 ( .A(in[374]), .B(n4327), .Z(n4704) );
  ANDN U6231 ( .B(n4989), .A(n4328), .Z(n4329) );
  XOR U6232 ( .A(n4704), .B(n4329), .Z(out[766]) );
  XOR U6233 ( .A(in[375]), .B(n4330), .Z(n4707) );
  NOR U6234 ( .A(n4331), .B(n4993), .Z(n4332) );
  XOR U6235 ( .A(n4707), .B(n4332), .Z(out[767]) );
  XOR U6236 ( .A(in[743]), .B(n4333), .Z(n4555) );
  IV U6237 ( .A(n4555), .Z(n4710) );
  XOR U6238 ( .A(in[744]), .B(n4335), .Z(n4558) );
  IV U6239 ( .A(n4558), .Z(n4714) );
  ANDN U6240 ( .B(n4338), .A(n4337), .Z(n4339) );
  XOR U6241 ( .A(n4340), .B(n4339), .Z(out[76]) );
  XOR U6242 ( .A(in[745]), .B(n4341), .Z(n4561) );
  IV U6243 ( .A(n4561), .Z(n4718) );
  XOR U6244 ( .A(in[746]), .B(n4343), .Z(n4564) );
  IV U6245 ( .A(n4564), .Z(n4722) );
  XNOR U6246 ( .A(in[747]), .B(n4345), .Z(n4734) );
  NANDN U6247 ( .A(n4346), .B(n4566), .Z(n4347) );
  XOR U6248 ( .A(n4734), .B(n4347), .Z(out[772]) );
  XNOR U6249 ( .A(in[748]), .B(n4348), .Z(n4738) );
  NANDN U6250 ( .A(n4349), .B(n4568), .Z(n4350) );
  XOR U6251 ( .A(n4738), .B(n4350), .Z(out[773]) );
  XNOR U6252 ( .A(in[749]), .B(n4351), .Z(n4742) );
  NANDN U6253 ( .A(n4352), .B(n4570), .Z(n4353) );
  XOR U6254 ( .A(n4742), .B(n4353), .Z(out[774]) );
  XOR U6255 ( .A(in[750]), .B(n4354), .Z(n4573) );
  IV U6256 ( .A(n4573), .Z(n4746) );
  XNOR U6257 ( .A(in[751]), .B(n4356), .Z(n4751) );
  NANDN U6258 ( .A(n4357), .B(n4579), .Z(n4358) );
  XOR U6259 ( .A(n4751), .B(n4358), .Z(out[776]) );
  XNOR U6260 ( .A(in[752]), .B(n4359), .Z(n4755) );
  NANDN U6261 ( .A(n4360), .B(n4581), .Z(n4361) );
  XOR U6262 ( .A(n4755), .B(n4361), .Z(out[777]) );
  XNOR U6263 ( .A(in[753]), .B(n4362), .Z(n4759) );
  NANDN U6264 ( .A(n4363), .B(n4583), .Z(n4364) );
  XOR U6265 ( .A(n4759), .B(n4364), .Z(out[778]) );
  XNOR U6266 ( .A(in[754]), .B(n4365), .Z(n4763) );
  NANDN U6267 ( .A(n4366), .B(n4585), .Z(n4367) );
  XOR U6268 ( .A(n4763), .B(n4367), .Z(out[779]) );
  ANDN U6269 ( .B(n4369), .A(n4368), .Z(n4370) );
  XOR U6270 ( .A(n4371), .B(n4370), .Z(out[77]) );
  XNOR U6271 ( .A(in[755]), .B(n4372), .Z(n4767) );
  NANDN U6272 ( .A(n4373), .B(n4587), .Z(n4374) );
  XOR U6273 ( .A(n4767), .B(n4374), .Z(out[780]) );
  XNOR U6274 ( .A(in[756]), .B(n4375), .Z(n4771) );
  NANDN U6275 ( .A(n4376), .B(n4589), .Z(n4377) );
  XOR U6276 ( .A(n4771), .B(n4377), .Z(out[781]) );
  XNOR U6277 ( .A(in[757]), .B(n4378), .Z(n4779) );
  NANDN U6278 ( .A(n4379), .B(n4591), .Z(n4380) );
  XOR U6279 ( .A(n4779), .B(n4380), .Z(out[782]) );
  XNOR U6280 ( .A(in[758]), .B(n4381), .Z(n4783) );
  NANDN U6281 ( .A(n4382), .B(n4593), .Z(n4383) );
  XOR U6282 ( .A(n4783), .B(n4383), .Z(out[783]) );
  XOR U6283 ( .A(in[759]), .B(n4384), .Z(n4596) );
  IV U6284 ( .A(n4596), .Z(n4787) );
  XNOR U6285 ( .A(in[760]), .B(n4386), .Z(n4791) );
  NANDN U6286 ( .A(n4387), .B(n4598), .Z(n4388) );
  XOR U6287 ( .A(n4791), .B(n4388), .Z(out[785]) );
  XNOR U6288 ( .A(in[761]), .B(n4389), .Z(n4795) );
  NANDN U6289 ( .A(n4390), .B(n4604), .Z(n4391) );
  XOR U6290 ( .A(n4795), .B(n4391), .Z(out[786]) );
  XOR U6291 ( .A(in[762]), .B(n4392), .Z(n4799) );
  NANDN U6292 ( .A(n4393), .B(n4606), .Z(n4394) );
  XOR U6293 ( .A(n4799), .B(n4394), .Z(out[787]) );
  XOR U6294 ( .A(in[763]), .B(n4395), .Z(n4803) );
  NANDN U6295 ( .A(n4396), .B(n4608), .Z(n4397) );
  XOR U6296 ( .A(n4803), .B(n4397), .Z(out[788]) );
  XNOR U6297 ( .A(in[764]), .B(n4398), .Z(n4807) );
  NANDN U6298 ( .A(n4399), .B(n4610), .Z(n4400) );
  XOR U6299 ( .A(n4807), .B(n4400), .Z(out[789]) );
  ANDN U6300 ( .B(n4402), .A(n4401), .Z(n4403) );
  XOR U6301 ( .A(n4404), .B(n4403), .Z(out[78]) );
  XOR U6302 ( .A(in[765]), .B(n4405), .Z(n4613) );
  IV U6303 ( .A(n4613), .Z(n4811) );
  NANDN U6304 ( .A(n4612), .B(n4406), .Z(n4407) );
  XOR U6305 ( .A(n4811), .B(n4407), .Z(out[790]) );
  XOR U6306 ( .A(in[766]), .B(n4408), .Z(n4616) );
  IV U6307 ( .A(n4616), .Z(n4815) );
  NANDN U6308 ( .A(n4615), .B(n4409), .Z(n4410) );
  XOR U6309 ( .A(n4815), .B(n4410), .Z(out[791]) );
  XOR U6310 ( .A(in[767]), .B(n4411), .Z(n4619) );
  IV U6311 ( .A(n4619), .Z(n4823) );
  NANDN U6312 ( .A(n4618), .B(n4412), .Z(n4413) );
  XOR U6313 ( .A(n4823), .B(n4413), .Z(out[792]) );
  XOR U6314 ( .A(in[704]), .B(n4414), .Z(n4622) );
  IV U6315 ( .A(n4622), .Z(n4827) );
  NANDN U6316 ( .A(n4621), .B(n4415), .Z(n4416) );
  XOR U6317 ( .A(n4827), .B(n4416), .Z(out[793]) );
  XNOR U6318 ( .A(in[705]), .B(n4417), .Z(n4831) );
  NAND U6319 ( .A(n4418), .B(n4624), .Z(n4419) );
  XOR U6320 ( .A(n4831), .B(n4419), .Z(out[794]) );
  XNOR U6321 ( .A(in[706]), .B(n4420), .Z(n4835) );
  NAND U6322 ( .A(n4421), .B(n4626), .Z(n4422) );
  XOR U6323 ( .A(n4835), .B(n4422), .Z(out[795]) );
  XOR U6324 ( .A(in[707]), .B(n4423), .Z(n4632) );
  IV U6325 ( .A(n4632), .Z(n4839) );
  NANDN U6326 ( .A(n4631), .B(n4424), .Z(n4425) );
  XOR U6327 ( .A(n4839), .B(n4425), .Z(out[796]) );
  XOR U6328 ( .A(in[708]), .B(n4426), .Z(n4635) );
  IV U6329 ( .A(n4635), .Z(n4843) );
  NANDN U6330 ( .A(n4634), .B(n4427), .Z(n4428) );
  XOR U6331 ( .A(n4843), .B(n4428), .Z(out[797]) );
  XOR U6332 ( .A(in[709]), .B(n4429), .Z(n4638) );
  IV U6333 ( .A(n4638), .Z(n4847) );
  NANDN U6334 ( .A(n4637), .B(n4430), .Z(n4431) );
  XOR U6335 ( .A(n4847), .B(n4431), .Z(out[798]) );
  XOR U6336 ( .A(in[710]), .B(n4432), .Z(n4851) );
  NANDN U6337 ( .A(n4640), .B(n4433), .Z(n4434) );
  XOR U6338 ( .A(n4851), .B(n4434), .Z(out[799]) );
  ANDN U6339 ( .B(n4436), .A(n4435), .Z(n4437) );
  XOR U6340 ( .A(n4438), .B(n4437), .Z(out[79]) );
  OR U6341 ( .A(n4440), .B(n4439), .Z(n4441) );
  XNOR U6342 ( .A(n4442), .B(n4441), .Z(out[7]) );
  XOR U6343 ( .A(in[711]), .B(n4443), .Z(n4642) );
  IV U6344 ( .A(n4642), .Z(n4855) );
  NANDN U6345 ( .A(n4641), .B(n4444), .Z(n4445) );
  XOR U6346 ( .A(n4855), .B(n4445), .Z(out[800]) );
  XOR U6347 ( .A(in[712]), .B(n4446), .Z(n4645) );
  IV U6348 ( .A(n4645), .Z(n4859) );
  NANDN U6349 ( .A(n4644), .B(n4447), .Z(n4448) );
  XOR U6350 ( .A(n4859), .B(n4448), .Z(out[801]) );
  XOR U6351 ( .A(in[713]), .B(n4449), .Z(n4648) );
  IV U6352 ( .A(n4648), .Z(n4867) );
  NANDN U6353 ( .A(n4647), .B(n4450), .Z(n4451) );
  XOR U6354 ( .A(n4867), .B(n4451), .Z(out[802]) );
  XOR U6355 ( .A(in[714]), .B(n4452), .Z(n4651) );
  IV U6356 ( .A(n4651), .Z(n4871) );
  NANDN U6357 ( .A(n4650), .B(n4453), .Z(n4454) );
  XOR U6358 ( .A(n4871), .B(n4454), .Z(out[803]) );
  XOR U6359 ( .A(in[715]), .B(n4455), .Z(n4654) );
  IV U6360 ( .A(n4654), .Z(n4875) );
  NANDN U6361 ( .A(n4653), .B(n4456), .Z(n4457) );
  XOR U6362 ( .A(n4875), .B(n4457), .Z(out[804]) );
  XNOR U6363 ( .A(n4458), .B(in[716]), .Z(n4879) );
  NANDN U6364 ( .A(n4656), .B(n4459), .Z(n4460) );
  XNOR U6365 ( .A(n4879), .B(n4460), .Z(out[805]) );
  XNOR U6366 ( .A(n4461), .B(in[717]), .Z(n4883) );
  NANDN U6367 ( .A(n4663), .B(n4462), .Z(n4463) );
  XNOR U6368 ( .A(n4883), .B(n4463), .Z(out[806]) );
  XNOR U6369 ( .A(n4464), .B(in[718]), .Z(n4887) );
  NANDN U6370 ( .A(n4666), .B(n4465), .Z(n4466) );
  XNOR U6371 ( .A(n4887), .B(n4466), .Z(out[807]) );
  XNOR U6372 ( .A(n4467), .B(in[719]), .Z(n4891) );
  NANDN U6373 ( .A(n4667), .B(n4468), .Z(n4469) );
  XNOR U6374 ( .A(n4891), .B(n4469), .Z(out[808]) );
  XNOR U6375 ( .A(n4470), .B(in[720]), .Z(n4895) );
  NANDN U6376 ( .A(n4668), .B(n4471), .Z(n4472) );
  XNOR U6377 ( .A(n4895), .B(n4472), .Z(out[809]) );
  ANDN U6378 ( .B(n4474), .A(n4473), .Z(n4475) );
  XOR U6379 ( .A(n4476), .B(n4475), .Z(out[80]) );
  XNOR U6380 ( .A(n4477), .B(in[721]), .Z(n4899) );
  NANDN U6381 ( .A(n4669), .B(n4478), .Z(n4479) );
  XNOR U6382 ( .A(n4899), .B(n4479), .Z(out[810]) );
  XNOR U6383 ( .A(n4480), .B(in[722]), .Z(n4903) );
  NAND U6384 ( .A(n4481), .B(n4670), .Z(n4482) );
  XNOR U6385 ( .A(n4903), .B(n4482), .Z(out[811]) );
  XNOR U6386 ( .A(n4483), .B(in[723]), .Z(n4910) );
  NANDN U6387 ( .A(n4672), .B(n4484), .Z(n4485) );
  XNOR U6388 ( .A(n4910), .B(n4485), .Z(out[812]) );
  XNOR U6389 ( .A(in[724]), .B(n4486), .Z(n4914) );
  NANDN U6390 ( .A(n4673), .B(n4487), .Z(n4488) );
  XNOR U6391 ( .A(n4914), .B(n4488), .Z(out[813]) );
  XNOR U6392 ( .A(in[725]), .B(n4489), .Z(n4918) );
  NANDN U6393 ( .A(n4674), .B(n4490), .Z(n4491) );
  XNOR U6394 ( .A(n4918), .B(n4491), .Z(out[814]) );
  XNOR U6395 ( .A(in[726]), .B(n4492), .Z(n4922) );
  NANDN U6396 ( .A(n4675), .B(n4493), .Z(n4494) );
  XNOR U6397 ( .A(n4922), .B(n4494), .Z(out[815]) );
  XNOR U6398 ( .A(in[727]), .B(n4495), .Z(n4926) );
  NANDN U6399 ( .A(n4679), .B(n4496), .Z(n4497) );
  XNOR U6400 ( .A(n4926), .B(n4497), .Z(out[816]) );
  XNOR U6401 ( .A(in[728]), .B(n4498), .Z(n4930) );
  NANDN U6402 ( .A(n4680), .B(n4499), .Z(n4500) );
  XNOR U6403 ( .A(n4930), .B(n4500), .Z(out[817]) );
  XNOR U6404 ( .A(in[729]), .B(n4501), .Z(n4934) );
  NANDN U6405 ( .A(n4681), .B(n4502), .Z(n4503) );
  XNOR U6406 ( .A(n4934), .B(n4503), .Z(out[818]) );
  XNOR U6407 ( .A(in[730]), .B(n4504), .Z(n4938) );
  NANDN U6408 ( .A(n4682), .B(n4505), .Z(n4506) );
  XNOR U6409 ( .A(n4938), .B(n4506), .Z(out[819]) );
  ANDN U6410 ( .B(n4508), .A(n4507), .Z(n4509) );
  XOR U6411 ( .A(n4510), .B(n4509), .Z(out[81]) );
  XOR U6412 ( .A(in[731]), .B(n4511), .Z(n4942) );
  NANDN U6413 ( .A(n4683), .B(n4512), .Z(n4513) );
  XNOR U6414 ( .A(n4942), .B(n4513), .Z(out[820]) );
  XOR U6415 ( .A(in[732]), .B(n4514), .Z(n4946) );
  NANDN U6416 ( .A(n4684), .B(n4515), .Z(n4516) );
  XNOR U6417 ( .A(n4946), .B(n4516), .Z(out[821]) );
  XOR U6418 ( .A(in[733]), .B(n4517), .Z(n4954) );
  NANDN U6419 ( .A(n4685), .B(n4518), .Z(n4519) );
  XNOR U6420 ( .A(n4954), .B(n4519), .Z(out[822]) );
  XNOR U6421 ( .A(in[734]), .B(n4520), .Z(n4958) );
  IV U6422 ( .A(n4521), .Z(n4686) );
  NANDN U6423 ( .A(n4522), .B(n4686), .Z(n4523) );
  XNOR U6424 ( .A(n4958), .B(n4523), .Z(out[823]) );
  XNOR U6425 ( .A(in[735]), .B(n4524), .Z(n4962) );
  IV U6426 ( .A(n4525), .Z(n4688) );
  NANDN U6427 ( .A(n4526), .B(n4688), .Z(n4527) );
  XNOR U6428 ( .A(n4962), .B(n4527), .Z(out[824]) );
  XNOR U6429 ( .A(in[736]), .B(n4528), .Z(n4966) );
  IV U6430 ( .A(n4529), .Z(n4690) );
  NANDN U6431 ( .A(n4530), .B(n4690), .Z(n4531) );
  XNOR U6432 ( .A(n4966), .B(n4531), .Z(out[825]) );
  XNOR U6433 ( .A(in[737]), .B(n4532), .Z(n4970) );
  IV U6434 ( .A(n4533), .Z(n4695) );
  NANDN U6435 ( .A(n4534), .B(n4695), .Z(n4535) );
  XNOR U6436 ( .A(n4970), .B(n4535), .Z(out[826]) );
  XNOR U6437 ( .A(in[738]), .B(n4536), .Z(n4974) );
  IV U6438 ( .A(n4537), .Z(n4697) );
  NANDN U6439 ( .A(n4538), .B(n4697), .Z(n4539) );
  XNOR U6440 ( .A(n4974), .B(n4539), .Z(out[827]) );
  XNOR U6441 ( .A(in[739]), .B(n4540), .Z(n4978) );
  IV U6442 ( .A(n4541), .Z(n4699) );
  NANDN U6443 ( .A(n4542), .B(n4699), .Z(n4543) );
  XNOR U6444 ( .A(n4978), .B(n4543), .Z(out[828]) );
  XOR U6445 ( .A(in[740]), .B(n4544), .Z(n4702) );
  IV U6446 ( .A(n4702), .Z(n4982) );
  ANDN U6447 ( .B(n4547), .A(n4546), .Z(n4548) );
  XOR U6448 ( .A(n4549), .B(n4548), .Z(out[82]) );
  XOR U6449 ( .A(in[741]), .B(n4550), .Z(n4705) );
  IV U6450 ( .A(n4705), .Z(n4986) );
  XOR U6451 ( .A(in[742]), .B(n4552), .Z(n4708) );
  IV U6452 ( .A(n4708), .Z(n4990) );
  NANDN U6453 ( .A(n4555), .B(n4554), .Z(n4556) );
  XOR U6454 ( .A(n4711), .B(n4556), .Z(out[832]) );
  NANDN U6455 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U6456 ( .A(n4715), .B(n4559), .Z(out[833]) );
  NANDN U6457 ( .A(n4561), .B(n4560), .Z(n4562) );
  XOR U6458 ( .A(n4719), .B(n4562), .Z(out[834]) );
  NANDN U6459 ( .A(n4564), .B(n4563), .Z(n4565) );
  XOR U6460 ( .A(n4723), .B(n4565), .Z(out[835]) );
  NANDN U6461 ( .A(n4566), .B(n4734), .Z(n4567) );
  XOR U6462 ( .A(n4735), .B(n4567), .Z(out[836]) );
  NANDN U6463 ( .A(n4568), .B(n4738), .Z(n4569) );
  XOR U6464 ( .A(n4739), .B(n4569), .Z(out[837]) );
  NANDN U6465 ( .A(n4570), .B(n4742), .Z(n4571) );
  XOR U6466 ( .A(n4743), .B(n4571), .Z(out[838]) );
  NANDN U6467 ( .A(n4573), .B(n4572), .Z(n4574) );
  XOR U6468 ( .A(n4747), .B(n4574), .Z(out[839]) );
  ANDN U6469 ( .B(n4576), .A(n4575), .Z(n4577) );
  XOR U6470 ( .A(n4578), .B(n4577), .Z(out[83]) );
  NANDN U6471 ( .A(n4579), .B(n4751), .Z(n4580) );
  XNOR U6472 ( .A(n4750), .B(n4580), .Z(out[840]) );
  NANDN U6473 ( .A(n4581), .B(n4755), .Z(n4582) );
  XNOR U6474 ( .A(n4754), .B(n4582), .Z(out[841]) );
  NANDN U6475 ( .A(n4583), .B(n4759), .Z(n4584) );
  XNOR U6476 ( .A(n4758), .B(n4584), .Z(out[842]) );
  NANDN U6477 ( .A(n4585), .B(n4763), .Z(n4586) );
  XNOR U6478 ( .A(n4762), .B(n4586), .Z(out[843]) );
  NANDN U6479 ( .A(n4587), .B(n4767), .Z(n4588) );
  XNOR U6480 ( .A(n4766), .B(n4588), .Z(out[844]) );
  NANDN U6481 ( .A(n4589), .B(n4771), .Z(n4590) );
  XNOR U6482 ( .A(n4770), .B(n4590), .Z(out[845]) );
  NANDN U6483 ( .A(n4591), .B(n4779), .Z(n4592) );
  XNOR U6484 ( .A(n4778), .B(n4592), .Z(out[846]) );
  NANDN U6485 ( .A(n4593), .B(n4783), .Z(n4594) );
  XNOR U6486 ( .A(n4782), .B(n4594), .Z(out[847]) );
  NANDN U6487 ( .A(n4596), .B(n4595), .Z(n4597) );
  XNOR U6488 ( .A(n4786), .B(n4597), .Z(out[848]) );
  NANDN U6489 ( .A(n4598), .B(n4791), .Z(n4599) );
  XNOR U6490 ( .A(n4790), .B(n4599), .Z(out[849]) );
  ANDN U6491 ( .B(n4601), .A(n4600), .Z(n4602) );
  XOR U6492 ( .A(n4603), .B(n4602), .Z(out[84]) );
  NANDN U6493 ( .A(n4604), .B(n4795), .Z(n4605) );
  XNOR U6494 ( .A(n4794), .B(n4605), .Z(out[850]) );
  NANDN U6495 ( .A(n4606), .B(n4799), .Z(n4607) );
  XNOR U6496 ( .A(n4798), .B(n4607), .Z(out[851]) );
  NANDN U6497 ( .A(n4608), .B(n4803), .Z(n4609) );
  XNOR U6498 ( .A(n4802), .B(n4609), .Z(out[852]) );
  NANDN U6499 ( .A(n4610), .B(n4807), .Z(n4611) );
  XNOR U6500 ( .A(n4806), .B(n4611), .Z(out[853]) );
  NANDN U6501 ( .A(n4613), .B(n4612), .Z(n4614) );
  XNOR U6502 ( .A(n4810), .B(n4614), .Z(out[854]) );
  NANDN U6503 ( .A(n4616), .B(n4615), .Z(n4617) );
  XNOR U6504 ( .A(n4814), .B(n4617), .Z(out[855]) );
  NANDN U6505 ( .A(n4619), .B(n4618), .Z(n4620) );
  XNOR U6506 ( .A(n4822), .B(n4620), .Z(out[856]) );
  NANDN U6507 ( .A(n4622), .B(n4621), .Z(n4623) );
  XNOR U6508 ( .A(n4826), .B(n4623), .Z(out[857]) );
  NANDN U6509 ( .A(n4624), .B(n4831), .Z(n4625) );
  XNOR U6510 ( .A(n4830), .B(n4625), .Z(out[858]) );
  NANDN U6511 ( .A(n4626), .B(n4835), .Z(n4627) );
  XNOR U6512 ( .A(n4834), .B(n4627), .Z(out[859]) );
  NANDN U6513 ( .A(n4632), .B(n4631), .Z(n4633) );
  XNOR U6514 ( .A(n4838), .B(n4633), .Z(out[860]) );
  NANDN U6515 ( .A(n4635), .B(n4634), .Z(n4636) );
  XNOR U6516 ( .A(n4842), .B(n4636), .Z(out[861]) );
  NANDN U6517 ( .A(n4638), .B(n4637), .Z(n4639) );
  XNOR U6518 ( .A(n4846), .B(n4639), .Z(out[862]) );
  NANDN U6519 ( .A(n4642), .B(n4641), .Z(n4643) );
  XNOR U6520 ( .A(n4854), .B(n4643), .Z(out[864]) );
  NANDN U6521 ( .A(n4645), .B(n4644), .Z(n4646) );
  XNOR U6522 ( .A(n4858), .B(n4646), .Z(out[865]) );
  NANDN U6523 ( .A(n4648), .B(n4647), .Z(n4649) );
  XNOR U6524 ( .A(n4866), .B(n4649), .Z(out[866]) );
  NANDN U6525 ( .A(n4651), .B(n4650), .Z(n4652) );
  XNOR U6526 ( .A(n4870), .B(n4652), .Z(out[867]) );
  NANDN U6527 ( .A(n4654), .B(n4653), .Z(n4655) );
  XNOR U6528 ( .A(n4874), .B(n4655), .Z(out[868]) );
  IV U6529 ( .A(n4656), .Z(n4657) );
  OR U6530 ( .A(n4879), .B(n4657), .Z(n4658) );
  XNOR U6531 ( .A(n4878), .B(n4658), .Z(out[869]) );
  ANDN U6532 ( .B(n4660), .A(n4659), .Z(n4661) );
  XOR U6533 ( .A(n4662), .B(n4661), .Z(out[86]) );
  IV U6534 ( .A(n4663), .Z(n4664) );
  OR U6535 ( .A(n4883), .B(n4664), .Z(n4665) );
  XNOR U6536 ( .A(n4882), .B(n4665), .Z(out[870]) );
  OR U6537 ( .A(n4903), .B(n4670), .Z(n4671) );
  XNOR U6538 ( .A(n4902), .B(n4671), .Z(out[875]) );
  OR U6539 ( .A(n4958), .B(n4686), .Z(n4687) );
  XOR U6540 ( .A(n4959), .B(n4687), .Z(out[887]) );
  OR U6541 ( .A(n4962), .B(n4688), .Z(n4689) );
  XOR U6542 ( .A(n4963), .B(n4689), .Z(out[888]) );
  OR U6543 ( .A(n4966), .B(n4690), .Z(n4691) );
  XOR U6544 ( .A(n4967), .B(n4691), .Z(out[889]) );
  OR U6545 ( .A(n4970), .B(n4695), .Z(n4696) );
  XOR U6546 ( .A(n4971), .B(n4696), .Z(out[890]) );
  OR U6547 ( .A(n4974), .B(n4697), .Z(n4698) );
  XOR U6548 ( .A(n4975), .B(n4698), .Z(out[891]) );
  OR U6549 ( .A(n4978), .B(n4699), .Z(n4700) );
  XOR U6550 ( .A(n4979), .B(n4700), .Z(out[892]) );
  NANDN U6551 ( .A(n4702), .B(n4701), .Z(n4703) );
  XOR U6552 ( .A(n4983), .B(n4703), .Z(out[893]) );
  NANDN U6553 ( .A(n4705), .B(n4704), .Z(n4706) );
  XOR U6554 ( .A(n4987), .B(n4706), .Z(out[894]) );
  NANDN U6555 ( .A(n4708), .B(n4707), .Z(n4709) );
  XOR U6556 ( .A(n4991), .B(n4709), .Z(out[895]) );
  ANDN U6557 ( .B(n4711), .A(n4710), .Z(n4712) );
  XOR U6558 ( .A(n4713), .B(n4712), .Z(out[896]) );
  ANDN U6559 ( .B(n4715), .A(n4714), .Z(n4716) );
  XOR U6560 ( .A(n4717), .B(n4716), .Z(out[897]) );
  ANDN U6561 ( .B(n4719), .A(n4718), .Z(n4720) );
  XOR U6562 ( .A(n4721), .B(n4720), .Z(out[898]) );
  ANDN U6563 ( .B(n4723), .A(n4722), .Z(n4724) );
  XOR U6564 ( .A(n4725), .B(n4724), .Z(out[899]) );
  ANDN U6565 ( .B(n4727), .A(n4726), .Z(n4728) );
  XOR U6566 ( .A(n4729), .B(n4728), .Z(out[89]) );
  OR U6567 ( .A(n4731), .B(n4730), .Z(n4732) );
  XNOR U6568 ( .A(n4733), .B(n4732), .Z(out[8]) );
  ANDN U6569 ( .B(n4735), .A(n4734), .Z(n4736) );
  XOR U6570 ( .A(n4737), .B(n4736), .Z(out[900]) );
  ANDN U6571 ( .B(n4739), .A(n4738), .Z(n4740) );
  XOR U6572 ( .A(n4741), .B(n4740), .Z(out[901]) );
  ANDN U6573 ( .B(n4743), .A(n4742), .Z(n4744) );
  XOR U6574 ( .A(n4745), .B(n4744), .Z(out[902]) );
  ANDN U6575 ( .B(n4747), .A(n4746), .Z(n4748) );
  XOR U6576 ( .A(n4749), .B(n4748), .Z(out[903]) );
  NOR U6577 ( .A(n4751), .B(n4750), .Z(n4752) );
  XOR U6578 ( .A(n4753), .B(n4752), .Z(out[904]) );
  NOR U6579 ( .A(n4755), .B(n4754), .Z(n4756) );
  XOR U6580 ( .A(n4757), .B(n4756), .Z(out[905]) );
  NOR U6581 ( .A(n4759), .B(n4758), .Z(n4760) );
  XOR U6582 ( .A(n4761), .B(n4760), .Z(out[906]) );
  NOR U6583 ( .A(n4763), .B(n4762), .Z(n4764) );
  XOR U6584 ( .A(n4765), .B(n4764), .Z(out[907]) );
  NOR U6585 ( .A(n4767), .B(n4766), .Z(n4768) );
  XOR U6586 ( .A(n4769), .B(n4768), .Z(out[908]) );
  NOR U6587 ( .A(n4771), .B(n4770), .Z(n4772) );
  XOR U6588 ( .A(n4773), .B(n4772), .Z(out[909]) );
  ANDN U6589 ( .B(n4775), .A(n4774), .Z(n4776) );
  XOR U6590 ( .A(n4777), .B(n4776), .Z(out[90]) );
  NOR U6591 ( .A(n4779), .B(n4778), .Z(n4780) );
  XOR U6592 ( .A(n4781), .B(n4780), .Z(out[910]) );
  NOR U6593 ( .A(n4783), .B(n4782), .Z(n4784) );
  XOR U6594 ( .A(n4785), .B(n4784), .Z(out[911]) );
  NOR U6595 ( .A(n4787), .B(n4786), .Z(n4788) );
  XOR U6596 ( .A(n4789), .B(n4788), .Z(out[912]) );
  NOR U6597 ( .A(n4791), .B(n4790), .Z(n4792) );
  XOR U6598 ( .A(n4793), .B(n4792), .Z(out[913]) );
  NOR U6599 ( .A(n4795), .B(n4794), .Z(n4796) );
  XOR U6600 ( .A(n4797), .B(n4796), .Z(out[914]) );
  NOR U6601 ( .A(n4799), .B(n4798), .Z(n4800) );
  XOR U6602 ( .A(n4801), .B(n4800), .Z(out[915]) );
  NOR U6603 ( .A(n4803), .B(n4802), .Z(n4804) );
  XOR U6604 ( .A(n4805), .B(n4804), .Z(out[916]) );
  NOR U6605 ( .A(n4807), .B(n4806), .Z(n4808) );
  XOR U6606 ( .A(n4809), .B(n4808), .Z(out[917]) );
  NOR U6607 ( .A(n4811), .B(n4810), .Z(n4812) );
  XOR U6608 ( .A(n4813), .B(n4812), .Z(out[918]) );
  NOR U6609 ( .A(n4815), .B(n4814), .Z(n4816) );
  XOR U6610 ( .A(n4817), .B(n4816), .Z(out[919]) );
  ANDN U6611 ( .B(n4819), .A(n4818), .Z(n4820) );
  XOR U6612 ( .A(n4821), .B(n4820), .Z(out[91]) );
  NOR U6613 ( .A(n4823), .B(n4822), .Z(n4824) );
  XOR U6614 ( .A(n4825), .B(n4824), .Z(out[920]) );
  NOR U6615 ( .A(n4827), .B(n4826), .Z(n4828) );
  XOR U6616 ( .A(n4829), .B(n4828), .Z(out[921]) );
  NOR U6617 ( .A(n4831), .B(n4830), .Z(n4832) );
  XOR U6618 ( .A(n4833), .B(n4832), .Z(out[922]) );
  NOR U6619 ( .A(n4835), .B(n4834), .Z(n4836) );
  XOR U6620 ( .A(n4837), .B(n4836), .Z(out[923]) );
  NOR U6621 ( .A(n4839), .B(n4838), .Z(n4840) );
  XOR U6622 ( .A(n4841), .B(n4840), .Z(out[924]) );
  NOR U6623 ( .A(n4843), .B(n4842), .Z(n4844) );
  XOR U6624 ( .A(n4845), .B(n4844), .Z(out[925]) );
  NOR U6625 ( .A(n4847), .B(n4846), .Z(n4848) );
  XOR U6626 ( .A(n4849), .B(n4848), .Z(out[926]) );
  NOR U6627 ( .A(n4851), .B(n4850), .Z(n4852) );
  XOR U6628 ( .A(n4853), .B(n4852), .Z(out[927]) );
  NOR U6629 ( .A(n4855), .B(n4854), .Z(n4856) );
  XOR U6630 ( .A(n4857), .B(n4856), .Z(out[928]) );
  NOR U6631 ( .A(n4859), .B(n4858), .Z(n4860) );
  XOR U6632 ( .A(n4861), .B(n4860), .Z(out[929]) );
  AND U6633 ( .A(n4863), .B(n4862), .Z(n4864) );
  XNOR U6634 ( .A(n4865), .B(n4864), .Z(out[92]) );
  NOR U6635 ( .A(n4867), .B(n4866), .Z(n4868) );
  XOR U6636 ( .A(n4869), .B(n4868), .Z(out[930]) );
  NOR U6637 ( .A(n4871), .B(n4870), .Z(n4872) );
  XOR U6638 ( .A(n4873), .B(n4872), .Z(out[931]) );
  NOR U6639 ( .A(n4875), .B(n4874), .Z(n4876) );
  XOR U6640 ( .A(n4877), .B(n4876), .Z(out[932]) );
  ANDN U6641 ( .B(n4879), .A(n4878), .Z(n4880) );
  XOR U6642 ( .A(n4881), .B(n4880), .Z(out[933]) );
  ANDN U6643 ( .B(n4883), .A(n4882), .Z(n4884) );
  XOR U6644 ( .A(n4885), .B(n4884), .Z(out[934]) );
  ANDN U6645 ( .B(n4887), .A(n4886), .Z(n4888) );
  XOR U6646 ( .A(n4889), .B(n4888), .Z(out[935]) );
  ANDN U6647 ( .B(n4891), .A(n4890), .Z(n4892) );
  XOR U6648 ( .A(n4893), .B(n4892), .Z(out[936]) );
  ANDN U6649 ( .B(n4895), .A(n4894), .Z(n4896) );
  XOR U6650 ( .A(n4897), .B(n4896), .Z(out[937]) );
  ANDN U6651 ( .B(n4899), .A(n4898), .Z(n4900) );
  XOR U6652 ( .A(n4901), .B(n4900), .Z(out[938]) );
  ANDN U6653 ( .B(n4903), .A(n4902), .Z(n4904) );
  XOR U6654 ( .A(n4905), .B(n4904), .Z(out[939]) );
  AND U6655 ( .A(n4907), .B(n4906), .Z(n4908) );
  XNOR U6656 ( .A(n4909), .B(n4908), .Z(out[93]) );
  AND U6657 ( .A(n4911), .B(n4910), .Z(n4912) );
  XNOR U6658 ( .A(n4913), .B(n4912), .Z(out[940]) );
  AND U6659 ( .A(n4915), .B(n4914), .Z(n4916) );
  XNOR U6660 ( .A(n4917), .B(n4916), .Z(out[941]) );
  AND U6661 ( .A(n4919), .B(n4918), .Z(n4920) );
  XNOR U6662 ( .A(n4921), .B(n4920), .Z(out[942]) );
  AND U6663 ( .A(n4923), .B(n4922), .Z(n4924) );
  XNOR U6664 ( .A(n4925), .B(n4924), .Z(out[943]) );
  AND U6665 ( .A(n4927), .B(n4926), .Z(n4928) );
  XNOR U6666 ( .A(n4929), .B(n4928), .Z(out[944]) );
  AND U6667 ( .A(n4931), .B(n4930), .Z(n4932) );
  XNOR U6668 ( .A(n4933), .B(n4932), .Z(out[945]) );
  AND U6669 ( .A(n4935), .B(n4934), .Z(n4936) );
  XNOR U6670 ( .A(n4937), .B(n4936), .Z(out[946]) );
  AND U6671 ( .A(n4939), .B(n4938), .Z(n4940) );
  XNOR U6672 ( .A(n4941), .B(n4940), .Z(out[947]) );
  AND U6673 ( .A(n4943), .B(n4942), .Z(n4944) );
  XNOR U6674 ( .A(n4945), .B(n4944), .Z(out[948]) );
  AND U6675 ( .A(n4947), .B(n4946), .Z(n4948) );
  XNOR U6676 ( .A(n4949), .B(n4948), .Z(out[949]) );
  AND U6677 ( .A(n4951), .B(n4950), .Z(n4952) );
  XNOR U6678 ( .A(n4953), .B(n4952), .Z(out[94]) );
  AND U6679 ( .A(n4955), .B(n4954), .Z(n4956) );
  XNOR U6680 ( .A(n4957), .B(n4956), .Z(out[950]) );
  AND U6681 ( .A(n4959), .B(n4958), .Z(n4960) );
  XNOR U6682 ( .A(n4961), .B(n4960), .Z(out[951]) );
  AND U6683 ( .A(n4963), .B(n4962), .Z(n4964) );
  XNOR U6684 ( .A(n4965), .B(n4964), .Z(out[952]) );
  AND U6685 ( .A(n4967), .B(n4966), .Z(n4968) );
  XNOR U6686 ( .A(n4969), .B(n4968), .Z(out[953]) );
  AND U6687 ( .A(n4971), .B(n4970), .Z(n4972) );
  XNOR U6688 ( .A(n4973), .B(n4972), .Z(out[954]) );
  AND U6689 ( .A(n4975), .B(n4974), .Z(n4976) );
  XNOR U6690 ( .A(n4977), .B(n4976), .Z(out[955]) );
  AND U6691 ( .A(n4979), .B(n4978), .Z(n4980) );
  XOR U6692 ( .A(n4981), .B(n4980), .Z(out[956]) );
  ANDN U6693 ( .B(n4983), .A(n4982), .Z(n4984) );
  XOR U6694 ( .A(n4985), .B(n4984), .Z(out[957]) );
  ANDN U6695 ( .B(n4987), .A(n4986), .Z(n4988) );
  XOR U6696 ( .A(n4989), .B(n4988), .Z(out[958]) );
  ANDN U6697 ( .B(n4991), .A(n4990), .Z(n4992) );
  XNOR U6698 ( .A(n4993), .B(n4992), .Z(out[959]) );
  AND U6699 ( .A(n4995), .B(n4994), .Z(n4996) );
  XNOR U6700 ( .A(n4997), .B(n4996), .Z(out[95]) );
  ANDN U6701 ( .B(n4999), .A(n4998), .Z(n5000) );
  XOR U6702 ( .A(n5001), .B(n5000), .Z(out[960]) );
  ANDN U6703 ( .B(n5003), .A(n5002), .Z(n5004) );
  XOR U6704 ( .A(n5005), .B(n5004), .Z(out[961]) );
  ANDN U6705 ( .B(n5007), .A(n5006), .Z(n5008) );
  XOR U6706 ( .A(n5009), .B(n5008), .Z(out[962]) );
  ANDN U6707 ( .B(n5011), .A(n5010), .Z(n5012) );
  XOR U6708 ( .A(n5013), .B(n5012), .Z(out[963]) );
  ANDN U6709 ( .B(n5015), .A(n5014), .Z(n5016) );
  XOR U6710 ( .A(n5017), .B(n5016), .Z(out[964]) );
  ANDN U6711 ( .B(n5019), .A(n5018), .Z(n5020) );
  XOR U6712 ( .A(n5021), .B(n5020), .Z(out[965]) );
  ANDN U6713 ( .B(n5023), .A(n5022), .Z(n5024) );
  XOR U6714 ( .A(n5025), .B(n5024), .Z(out[966]) );
  ANDN U6715 ( .B(n5027), .A(n5026), .Z(n5028) );
  XOR U6716 ( .A(n5029), .B(n5028), .Z(out[967]) );
  ANDN U6717 ( .B(n5031), .A(n5030), .Z(n5032) );
  XOR U6718 ( .A(n5033), .B(n5032), .Z(out[968]) );
  ANDN U6719 ( .B(n5035), .A(n5034), .Z(n5036) );
  XOR U6720 ( .A(n5037), .B(n5036), .Z(out[969]) );
  AND U6721 ( .A(n5039), .B(n5038), .Z(n5040) );
  XNOR U6722 ( .A(n5041), .B(n5040), .Z(out[96]) );
  ANDN U6723 ( .B(n5043), .A(n5042), .Z(n5044) );
  XOR U6724 ( .A(n5045), .B(n5044), .Z(out[970]) );
  ANDN U6725 ( .B(n5047), .A(n5046), .Z(n5048) );
  XOR U6726 ( .A(n5049), .B(n5048), .Z(out[971]) );
  ANDN U6727 ( .B(n5051), .A(n5050), .Z(n5052) );
  XOR U6728 ( .A(n5053), .B(n5052), .Z(out[972]) );
  ANDN U6729 ( .B(n5055), .A(n5054), .Z(n5056) );
  XOR U6730 ( .A(n5057), .B(n5056), .Z(out[973]) );
  ANDN U6731 ( .B(n5059), .A(n5058), .Z(n5060) );
  XOR U6732 ( .A(n5061), .B(n5060), .Z(out[974]) );
  ANDN U6733 ( .B(n5063), .A(n5062), .Z(n5064) );
  XOR U6734 ( .A(n5065), .B(n5064), .Z(out[975]) );
  ANDN U6735 ( .B(n5076), .A(n5075), .Z(n5077) );
  XOR U6736 ( .A(n5078), .B(n5077), .Z(out[979]) );
  AND U6737 ( .A(n5080), .B(n5079), .Z(n5081) );
  XNOR U6738 ( .A(n5082), .B(n5081), .Z(out[97]) );
  ANDN U6739 ( .B(n5108), .A(n5107), .Z(n5109) );
  XOR U6740 ( .A(n5110), .B(n5109), .Z(out[988]) );
  ANDN U6741 ( .B(n5115), .A(n5114), .Z(n5116) );
  XNOR U6742 ( .A(n5117), .B(n5116), .Z(out[98]) );
  ANDN U6743 ( .B(n5122), .A(n5121), .Z(n5123) );
  XOR U6744 ( .A(n5124), .B(n5123), .Z(out[991]) );
  ANDN U6745 ( .B(n5126), .A(n5125), .Z(n5127) );
  XOR U6746 ( .A(n5128), .B(n5127), .Z(out[992]) );
  ANDN U6747 ( .B(n5130), .A(n5129), .Z(n5131) );
  XOR U6748 ( .A(n5132), .B(n5131), .Z(out[993]) );
  ANDN U6749 ( .B(n5134), .A(n5133), .Z(n5135) );
  XOR U6750 ( .A(n5136), .B(n5135), .Z(out[994]) );
  ANDN U6751 ( .B(n5138), .A(n5137), .Z(n5139) );
  XNOR U6752 ( .A(n5140), .B(n5139), .Z(out[995]) );
  ANDN U6753 ( .B(n5142), .A(n5141), .Z(n5143) );
  XNOR U6754 ( .A(n5144), .B(n5143), .Z(out[996]) );
  ANDN U6755 ( .B(n5146), .A(n5145), .Z(n5147) );
  XNOR U6756 ( .A(n5148), .B(n5147), .Z(out[997]) );
  AND U6757 ( .A(n5150), .B(n5149), .Z(n5151) );
  XNOR U6758 ( .A(n5152), .B(n5151), .Z(out[998]) );
  ANDN U6759 ( .B(n5154), .A(n5153), .Z(n5155) );
  XNOR U6760 ( .A(n5156), .B(n5155), .Z(out[999]) );
  ANDN U6761 ( .B(n5158), .A(n5157), .Z(n5159) );
  XNOR U6762 ( .A(n5160), .B(n5159), .Z(out[99]) );
  OR U6763 ( .A(n5162), .B(n5161), .Z(n5163) );
  XNOR U6764 ( .A(n5164), .B(n5163), .Z(out[9]) );
endmodule


module sha3_seq_CC6 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N444, N445, N446, N447, N448, N449, N450, N451, N452, N453,
         N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464,
         N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N491, N492, N493, N494, N495, N496, N497,
         N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519,
         N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530,
         N531, N532, N533, N534, N535, N536, N537, N538, N539, N540, N541,
         N542, N543, N544, N545, N546, N547, N548, N549, N550, N551, N552,
         N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563,
         N564, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596,
         N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N614, N615, N616, N617, N618,
         N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629,
         N630, N631, N632, N633, N634, N635, N636, N637, N638, N639, N640,
         N641, N642, N643, N644, N645, N646, N647, N648, N649, N650, N651,
         N652, N653, N654, N655, N656, N657, N658, N659, N660, N661, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N679, N680, N681, N682, N683, N684,
         N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695,
         N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706,
         N707, N708, N709, N710, N711, N712, N713, N714, N715, N716, N717,
         N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183,
         N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193,
         N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203,
         N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213,
         N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223,
         N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233,
         N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243,
         N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253,
         N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273,
         N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283,
         N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293,
         N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303,
         N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313,
         N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333,
         N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343,
         N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353,
         N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361, N1362, N1363,
         N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373,
         N1374, N1375, N1376, N1377, N1378, N1379, N1380, N1381, N1382, N1383,
         N1384, N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393,
         N1394, N1395, N1396, N1397, N1398, N1399, N1400, N1401, N1402, N1403,
         N1404, N1405, N1406, N1407, N1408, N1409, N1410, N1411, N1412, N1413,
         N1414, N1415, N1416, N1417, N1418, N1419, N1420, N1421, N1422, N1423,
         N1424, N1425, N1426, N1427, N1428, N1429, N1430, N1431, N1432, N1433,
         N1434, N1435, N1436, N1437, N1438, N1439, N1440, N1441, N1442, N1443,
         N1444, N1445, N1446, N1447, N1448, N1449, N1450, N1451, N1452, N1453,
         N1454, N1455, N1456, N1457, N1458, N1459, N1460, N1461, N1462, N1463,
         N1464, N1465, N1466, N1467, N1468, N1469, N1470, N1471, N1472, N1473,
         N1474, N1475, N1476, N1477, N1478, N1479, N1480, N1481, N1482, N1483,
         N1484, N1485, N1486, N1487, N1488, N1489, N1490, N1491, N1492, N1493,
         N1494, N1495, N1496, N1497, N1498, N1499, N1500, N1501, N1502, N1503,
         N1504, N1505, N1506, N1507, N1508, N1509, N1510, N1511, N1512, N1513,
         N1514, N1515, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523,
         N1524, N1525, N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533,
         N1534, N1535, N1536, N1537, N1538, N1539, N1540, N1541, N1542, N1543,
         N1544, N1545, N1546, N1547, N1548, N1549, N1550, N1551, N1552, N1553,
         N1554, N1555, N1556, N1557, N1558, N1559, N1560, N1561, N1562, N1563,
         N1564, N1565, N1566, N1567, N1568, N1569, N1570, N1571, N1572, N1573,
         N1574, N1575, N1576, N1577, N1578, N1579, N1580, N1581, N1582, N1583,
         N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593,
         N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602, N1603,
         N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1611,
         \round_in[3][1599] , \round_in[3][1598] , \round_in[3][1597] ,
         \round_in[3][1596] , \round_in[3][1595] , \round_in[3][1594] ,
         \round_in[3][1593] , \round_in[3][1592] , \round_in[3][1591] ,
         \round_in[3][1590] , \round_in[3][1589] , \round_in[3][1588] ,
         \round_in[3][1587] , \round_in[3][1586] , \round_in[3][1585] ,
         \round_in[3][1584] , \round_in[3][1583] , \round_in[3][1582] ,
         \round_in[3][1581] , \round_in[3][1580] , \round_in[3][1579] ,
         \round_in[3][1578] , \round_in[3][1577] , \round_in[3][1576] ,
         \round_in[3][1575] , \round_in[3][1574] , \round_in[3][1573] ,
         \round_in[3][1572] , \round_in[3][1571] , \round_in[3][1570] ,
         \round_in[3][1569] , \round_in[3][1568] , \round_in[3][1567] ,
         \round_in[3][1566] , \round_in[3][1565] , \round_in[3][1564] ,
         \round_in[3][1563] , \round_in[3][1562] , \round_in[3][1561] ,
         \round_in[3][1560] , \round_in[3][1559] , \round_in[3][1558] ,
         \round_in[3][1557] , \round_in[3][1556] , \round_in[3][1555] ,
         \round_in[3][1554] , \round_in[3][1553] , \round_in[3][1552] ,
         \round_in[3][1551] , \round_in[3][1550] , \round_in[3][1549] ,
         \round_in[3][1548] , \round_in[3][1547] , \round_in[3][1546] ,
         \round_in[3][1545] , \round_in[3][1544] , \round_in[3][1543] ,
         \round_in[3][1542] , \round_in[3][1541] , \round_in[3][1540] ,
         \round_in[3][1539] , \round_in[3][1538] , \round_in[3][1537] ,
         \round_in[3][1536] , \round_in[3][1535] , \round_in[3][1534] ,
         \round_in[3][1533] , \round_in[3][1532] , \round_in[3][1531] ,
         \round_in[3][1530] , \round_in[3][1529] , \round_in[3][1528] ,
         \round_in[3][1527] , \round_in[3][1526] , \round_in[3][1525] ,
         \round_in[3][1524] , \round_in[3][1523] , \round_in[3][1522] ,
         \round_in[3][1521] , \round_in[3][1520] , \round_in[3][1519] ,
         \round_in[3][1518] , \round_in[3][1517] , \round_in[3][1516] ,
         \round_in[3][1515] , \round_in[3][1514] , \round_in[3][1513] ,
         \round_in[3][1512] , \round_in[3][1511] , \round_in[3][1510] ,
         \round_in[3][1509] , \round_in[3][1508] , \round_in[3][1507] ,
         \round_in[3][1506] , \round_in[3][1505] , \round_in[3][1504] ,
         \round_in[3][1503] , \round_in[3][1502] , \round_in[3][1501] ,
         \round_in[3][1500] , \round_in[3][1499] , \round_in[3][1498] ,
         \round_in[3][1497] , \round_in[3][1496] , \round_in[3][1495] ,
         \round_in[3][1494] , \round_in[3][1493] , \round_in[3][1492] ,
         \round_in[3][1491] , \round_in[3][1490] , \round_in[3][1489] ,
         \round_in[3][1488] , \round_in[3][1487] , \round_in[3][1486] ,
         \round_in[3][1485] , \round_in[3][1484] , \round_in[3][1483] ,
         \round_in[3][1482] , \round_in[3][1481] , \round_in[3][1480] ,
         \round_in[3][1479] , \round_in[3][1478] , \round_in[3][1477] ,
         \round_in[3][1476] , \round_in[3][1475] , \round_in[3][1474] ,
         \round_in[3][1473] , \round_in[3][1472] , \round_in[3][1471] ,
         \round_in[3][1470] , \round_in[3][1469] , \round_in[3][1468] ,
         \round_in[3][1467] , \round_in[3][1466] , \round_in[3][1465] ,
         \round_in[3][1464] , \round_in[3][1463] , \round_in[3][1462] ,
         \round_in[3][1461] , \round_in[3][1460] , \round_in[3][1459] ,
         \round_in[3][1458] , \round_in[3][1457] , \round_in[3][1456] ,
         \round_in[3][1455] , \round_in[3][1454] , \round_in[3][1453] ,
         \round_in[3][1452] , \round_in[3][1451] , \round_in[3][1450] ,
         \round_in[3][1449] , \round_in[3][1448] , \round_in[3][1447] ,
         \round_in[3][1446] , \round_in[3][1445] , \round_in[3][1444] ,
         \round_in[3][1443] , \round_in[3][1442] , \round_in[3][1441] ,
         \round_in[3][1440] , \round_in[3][1439] , \round_in[3][1438] ,
         \round_in[3][1437] , \round_in[3][1436] , \round_in[3][1435] ,
         \round_in[3][1434] , \round_in[3][1433] , \round_in[3][1432] ,
         \round_in[3][1431] , \round_in[3][1430] , \round_in[3][1429] ,
         \round_in[3][1428] , \round_in[3][1427] , \round_in[3][1426] ,
         \round_in[3][1425] , \round_in[3][1424] , \round_in[3][1423] ,
         \round_in[3][1422] , \round_in[3][1421] , \round_in[3][1420] ,
         \round_in[3][1419] , \round_in[3][1418] , \round_in[3][1417] ,
         \round_in[3][1416] , \round_in[3][1415] , \round_in[3][1414] ,
         \round_in[3][1413] , \round_in[3][1412] , \round_in[3][1411] ,
         \round_in[3][1410] , \round_in[3][1409] , \round_in[3][1408] ,
         \round_in[3][1407] , \round_in[3][1406] , \round_in[3][1405] ,
         \round_in[3][1404] , \round_in[3][1403] , \round_in[3][1402] ,
         \round_in[3][1401] , \round_in[3][1400] , \round_in[3][1399] ,
         \round_in[3][1398] , \round_in[3][1397] , \round_in[3][1396] ,
         \round_in[3][1395] , \round_in[3][1394] , \round_in[3][1393] ,
         \round_in[3][1392] , \round_in[3][1391] , \round_in[3][1390] ,
         \round_in[3][1389] , \round_in[3][1388] , \round_in[3][1387] ,
         \round_in[3][1386] , \round_in[3][1385] , \round_in[3][1384] ,
         \round_in[3][1383] , \round_in[3][1382] , \round_in[3][1381] ,
         \round_in[3][1380] , \round_in[3][1379] , \round_in[3][1378] ,
         \round_in[3][1377] , \round_in[3][1376] , \round_in[3][1375] ,
         \round_in[3][1374] , \round_in[3][1373] , \round_in[3][1372] ,
         \round_in[3][1371] , \round_in[3][1370] , \round_in[3][1369] ,
         \round_in[3][1368] , \round_in[3][1367] , \round_in[3][1366] ,
         \round_in[3][1365] , \round_in[3][1364] , \round_in[3][1363] ,
         \round_in[3][1362] , \round_in[3][1361] , \round_in[3][1360] ,
         \round_in[3][1359] , \round_in[3][1358] , \round_in[3][1357] ,
         \round_in[3][1356] , \round_in[3][1355] , \round_in[3][1354] ,
         \round_in[3][1353] , \round_in[3][1352] , \round_in[3][1351] ,
         \round_in[3][1350] , \round_in[3][1349] , \round_in[3][1348] ,
         \round_in[3][1347] , \round_in[3][1346] , \round_in[3][1345] ,
         \round_in[3][1344] , \round_in[3][1343] , \round_in[3][1342] ,
         \round_in[3][1341] , \round_in[3][1340] , \round_in[3][1339] ,
         \round_in[3][1338] , \round_in[3][1337] , \round_in[3][1336] ,
         \round_in[3][1335] , \round_in[3][1334] , \round_in[3][1333] ,
         \round_in[3][1332] , \round_in[3][1331] , \round_in[3][1330] ,
         \round_in[3][1329] , \round_in[3][1328] , \round_in[3][1327] ,
         \round_in[3][1326] , \round_in[3][1325] , \round_in[3][1324] ,
         \round_in[3][1323] , \round_in[3][1322] , \round_in[3][1321] ,
         \round_in[3][1320] , \round_in[3][1319] , \round_in[3][1318] ,
         \round_in[3][1317] , \round_in[3][1316] , \round_in[3][1315] ,
         \round_in[3][1314] , \round_in[3][1313] , \round_in[3][1312] ,
         \round_in[3][1311] , \round_in[3][1310] , \round_in[3][1309] ,
         \round_in[3][1308] , \round_in[3][1307] , \round_in[3][1306] ,
         \round_in[3][1305] , \round_in[3][1304] , \round_in[3][1303] ,
         \round_in[3][1302] , \round_in[3][1301] , \round_in[3][1300] ,
         \round_in[3][1299] , \round_in[3][1298] , \round_in[3][1297] ,
         \round_in[3][1296] , \round_in[3][1295] , \round_in[3][1294] ,
         \round_in[3][1293] , \round_in[3][1292] , \round_in[3][1291] ,
         \round_in[3][1290] , \round_in[3][1289] , \round_in[3][1288] ,
         \round_in[3][1287] , \round_in[3][1286] , \round_in[3][1285] ,
         \round_in[3][1284] , \round_in[3][1283] , \round_in[3][1282] ,
         \round_in[3][1281] , \round_in[3][1280] , \round_in[3][1279] ,
         \round_in[3][1278] , \round_in[3][1277] , \round_in[3][1276] ,
         \round_in[3][1275] , \round_in[3][1274] , \round_in[3][1273] ,
         \round_in[3][1272] , \round_in[3][1271] , \round_in[3][1270] ,
         \round_in[3][1269] , \round_in[3][1268] , \round_in[3][1267] ,
         \round_in[3][1266] , \round_in[3][1265] , \round_in[3][1264] ,
         \round_in[3][1263] , \round_in[3][1262] , \round_in[3][1261] ,
         \round_in[3][1260] , \round_in[3][1259] , \round_in[3][1258] ,
         \round_in[3][1257] , \round_in[3][1256] , \round_in[3][1255] ,
         \round_in[3][1254] , \round_in[3][1253] , \round_in[3][1252] ,
         \round_in[3][1251] , \round_in[3][1250] , \round_in[3][1249] ,
         \round_in[3][1248] , \round_in[3][1247] , \round_in[3][1246] ,
         \round_in[3][1245] , \round_in[3][1244] , \round_in[3][1243] ,
         \round_in[3][1242] , \round_in[3][1241] , \round_in[3][1240] ,
         \round_in[3][1239] , \round_in[3][1238] , \round_in[3][1237] ,
         \round_in[3][1236] , \round_in[3][1235] , \round_in[3][1234] ,
         \round_in[3][1233] , \round_in[3][1232] , \round_in[3][1231] ,
         \round_in[3][1230] , \round_in[3][1229] , \round_in[3][1228] ,
         \round_in[3][1227] , \round_in[3][1226] , \round_in[3][1225] ,
         \round_in[3][1224] , \round_in[3][1223] , \round_in[3][1222] ,
         \round_in[3][1221] , \round_in[3][1220] , \round_in[3][1219] ,
         \round_in[3][1218] , \round_in[3][1217] , \round_in[3][1216] ,
         \round_in[3][1215] , \round_in[3][1214] , \round_in[3][1213] ,
         \round_in[3][1212] , \round_in[3][1211] , \round_in[3][1210] ,
         \round_in[3][1209] , \round_in[3][1208] , \round_in[3][1207] ,
         \round_in[3][1206] , \round_in[3][1205] , \round_in[3][1204] ,
         \round_in[3][1203] , \round_in[3][1202] , \round_in[3][1201] ,
         \round_in[3][1200] , \round_in[3][1199] , \round_in[3][1198] ,
         \round_in[3][1197] , \round_in[3][1196] , \round_in[3][1195] ,
         \round_in[3][1194] , \round_in[3][1193] , \round_in[3][1192] ,
         \round_in[3][1191] , \round_in[3][1190] , \round_in[3][1189] ,
         \round_in[3][1188] , \round_in[3][1187] , \round_in[3][1186] ,
         \round_in[3][1185] , \round_in[3][1184] , \round_in[3][1183] ,
         \round_in[3][1182] , \round_in[3][1181] , \round_in[3][1180] ,
         \round_in[3][1179] , \round_in[3][1178] , \round_in[3][1177] ,
         \round_in[3][1176] , \round_in[3][1175] , \round_in[3][1174] ,
         \round_in[3][1173] , \round_in[3][1172] , \round_in[3][1171] ,
         \round_in[3][1170] , \round_in[3][1169] , \round_in[3][1168] ,
         \round_in[3][1167] , \round_in[3][1166] , \round_in[3][1165] ,
         \round_in[3][1164] , \round_in[3][1163] , \round_in[3][1162] ,
         \round_in[3][1161] , \round_in[3][1160] , \round_in[3][1159] ,
         \round_in[3][1158] , \round_in[3][1157] , \round_in[3][1156] ,
         \round_in[3][1155] , \round_in[3][1154] , \round_in[3][1153] ,
         \round_in[3][1152] , \round_in[3][1151] , \round_in[3][1150] ,
         \round_in[3][1149] , \round_in[3][1148] , \round_in[3][1147] ,
         \round_in[3][1146] , \round_in[3][1145] , \round_in[3][1144] ,
         \round_in[3][1143] , \round_in[3][1142] , \round_in[3][1141] ,
         \round_in[3][1140] , \round_in[3][1139] , \round_in[3][1138] ,
         \round_in[3][1137] , \round_in[3][1136] , \round_in[3][1135] ,
         \round_in[3][1134] , \round_in[3][1133] , \round_in[3][1132] ,
         \round_in[3][1131] , \round_in[3][1130] , \round_in[3][1129] ,
         \round_in[3][1128] , \round_in[3][1127] , \round_in[3][1126] ,
         \round_in[3][1125] , \round_in[3][1124] , \round_in[3][1123] ,
         \round_in[3][1122] , \round_in[3][1121] , \round_in[3][1120] ,
         \round_in[3][1119] , \round_in[3][1118] , \round_in[3][1117] ,
         \round_in[3][1116] , \round_in[3][1115] , \round_in[3][1114] ,
         \round_in[3][1113] , \round_in[3][1112] , \round_in[3][1111] ,
         \round_in[3][1110] , \round_in[3][1109] , \round_in[3][1108] ,
         \round_in[3][1107] , \round_in[3][1106] , \round_in[3][1105] ,
         \round_in[3][1104] , \round_in[3][1103] , \round_in[3][1102] ,
         \round_in[3][1101] , \round_in[3][1100] , \round_in[3][1099] ,
         \round_in[3][1098] , \round_in[3][1097] , \round_in[3][1096] ,
         \round_in[3][1095] , \round_in[3][1094] , \round_in[3][1093] ,
         \round_in[3][1092] , \round_in[3][1091] , \round_in[3][1090] ,
         \round_in[3][1089] , \round_in[3][1088] , \round_in[3][1087] ,
         \round_in[3][1086] , \round_in[3][1085] , \round_in[3][1084] ,
         \round_in[3][1083] , \round_in[3][1082] , \round_in[3][1081] ,
         \round_in[3][1080] , \round_in[3][1079] , \round_in[3][1078] ,
         \round_in[3][1077] , \round_in[3][1076] , \round_in[3][1075] ,
         \round_in[3][1074] , \round_in[3][1073] , \round_in[3][1072] ,
         \round_in[3][1071] , \round_in[3][1070] , \round_in[3][1069] ,
         \round_in[3][1068] , \round_in[3][1067] , \round_in[3][1066] ,
         \round_in[3][1065] , \round_in[3][1064] , \round_in[3][1063] ,
         \round_in[3][1062] , \round_in[3][1061] , \round_in[3][1060] ,
         \round_in[3][1059] , \round_in[3][1058] , \round_in[3][1057] ,
         \round_in[3][1056] , \round_in[3][1055] , \round_in[3][1054] ,
         \round_in[3][1053] , \round_in[3][1052] , \round_in[3][1051] ,
         \round_in[3][1050] , \round_in[3][1049] , \round_in[3][1048] ,
         \round_in[3][1047] , \round_in[3][1046] , \round_in[3][1045] ,
         \round_in[3][1044] , \round_in[3][1043] , \round_in[3][1042] ,
         \round_in[3][1041] , \round_in[3][1040] , \round_in[3][1039] ,
         \round_in[3][1038] , \round_in[3][1037] , \round_in[3][1036] ,
         \round_in[3][1035] , \round_in[3][1034] , \round_in[3][1033] ,
         \round_in[3][1032] , \round_in[3][1031] , \round_in[3][1030] ,
         \round_in[3][1029] , \round_in[3][1028] , \round_in[3][1027] ,
         \round_in[3][1026] , \round_in[3][1025] , \round_in[3][1024] ,
         \round_in[3][1023] , \round_in[3][1022] , \round_in[3][1021] ,
         \round_in[3][1020] , \round_in[3][1019] , \round_in[3][1018] ,
         \round_in[3][1017] , \round_in[3][1016] , \round_in[3][1015] ,
         \round_in[3][1014] , \round_in[3][1013] , \round_in[3][1012] ,
         \round_in[3][1011] , \round_in[3][1010] , \round_in[3][1009] ,
         \round_in[3][1008] , \round_in[3][1007] , \round_in[3][1006] ,
         \round_in[3][1005] , \round_in[3][1004] , \round_in[3][1003] ,
         \round_in[3][1002] , \round_in[3][1001] , \round_in[3][1000] ,
         \round_in[3][999] , \round_in[3][998] , \round_in[3][997] ,
         \round_in[3][996] , \round_in[3][995] , \round_in[3][994] ,
         \round_in[3][993] , \round_in[3][992] , \round_in[3][991] ,
         \round_in[3][990] , \round_in[3][989] , \round_in[3][988] ,
         \round_in[3][987] , \round_in[3][986] , \round_in[3][985] ,
         \round_in[3][984] , \round_in[3][983] , \round_in[3][982] ,
         \round_in[3][981] , \round_in[3][980] , \round_in[3][979] ,
         \round_in[3][978] , \round_in[3][977] , \round_in[3][976] ,
         \round_in[3][975] , \round_in[3][974] , \round_in[3][973] ,
         \round_in[3][972] , \round_in[3][971] , \round_in[3][970] ,
         \round_in[3][969] , \round_in[3][968] , \round_in[3][967] ,
         \round_in[3][966] , \round_in[3][965] , \round_in[3][964] ,
         \round_in[3][963] , \round_in[3][962] , \round_in[3][961] ,
         \round_in[3][960] , \round_in[3][959] , \round_in[3][958] ,
         \round_in[3][957] , \round_in[3][956] , \round_in[3][955] ,
         \round_in[3][954] , \round_in[3][953] , \round_in[3][952] ,
         \round_in[3][951] , \round_in[3][950] , \round_in[3][949] ,
         \round_in[3][948] , \round_in[3][947] , \round_in[3][946] ,
         \round_in[3][945] , \round_in[3][944] , \round_in[3][943] ,
         \round_in[3][942] , \round_in[3][941] , \round_in[3][940] ,
         \round_in[3][939] , \round_in[3][938] , \round_in[3][937] ,
         \round_in[3][936] , \round_in[3][935] , \round_in[3][934] ,
         \round_in[3][933] , \round_in[3][932] , \round_in[3][931] ,
         \round_in[3][930] , \round_in[3][929] , \round_in[3][928] ,
         \round_in[3][927] , \round_in[3][926] , \round_in[3][925] ,
         \round_in[3][924] , \round_in[3][923] , \round_in[3][922] ,
         \round_in[3][921] , \round_in[3][920] , \round_in[3][919] ,
         \round_in[3][918] , \round_in[3][917] , \round_in[3][916] ,
         \round_in[3][915] , \round_in[3][914] , \round_in[3][913] ,
         \round_in[3][912] , \round_in[3][911] , \round_in[3][910] ,
         \round_in[3][909] , \round_in[3][908] , \round_in[3][907] ,
         \round_in[3][906] , \round_in[3][905] , \round_in[3][904] ,
         \round_in[3][903] , \round_in[3][902] , \round_in[3][901] ,
         \round_in[3][900] , \round_in[3][899] , \round_in[3][898] ,
         \round_in[3][897] , \round_in[3][896] , \round_in[3][895] ,
         \round_in[3][894] , \round_in[3][893] , \round_in[3][892] ,
         \round_in[3][891] , \round_in[3][890] , \round_in[3][889] ,
         \round_in[3][888] , \round_in[3][887] , \round_in[3][886] ,
         \round_in[3][885] , \round_in[3][884] , \round_in[3][883] ,
         \round_in[3][882] , \round_in[3][881] , \round_in[3][880] ,
         \round_in[3][879] , \round_in[3][878] , \round_in[3][877] ,
         \round_in[3][876] , \round_in[3][875] , \round_in[3][874] ,
         \round_in[3][873] , \round_in[3][872] , \round_in[3][871] ,
         \round_in[3][870] , \round_in[3][869] , \round_in[3][868] ,
         \round_in[3][867] , \round_in[3][866] , \round_in[3][865] ,
         \round_in[3][864] , \round_in[3][863] , \round_in[3][862] ,
         \round_in[3][861] , \round_in[3][860] , \round_in[3][859] ,
         \round_in[3][858] , \round_in[3][857] , \round_in[3][856] ,
         \round_in[3][855] , \round_in[3][854] , \round_in[3][853] ,
         \round_in[3][852] , \round_in[3][851] , \round_in[3][850] ,
         \round_in[3][849] , \round_in[3][848] , \round_in[3][847] ,
         \round_in[3][846] , \round_in[3][845] , \round_in[3][844] ,
         \round_in[3][843] , \round_in[3][842] , \round_in[3][841] ,
         \round_in[3][840] , \round_in[3][839] , \round_in[3][838] ,
         \round_in[3][837] , \round_in[3][836] , \round_in[3][835] ,
         \round_in[3][834] , \round_in[3][833] , \round_in[3][832] ,
         \round_in[3][831] , \round_in[3][830] , \round_in[3][829] ,
         \round_in[3][828] , \round_in[3][827] , \round_in[3][826] ,
         \round_in[3][825] , \round_in[3][824] , \round_in[3][823] ,
         \round_in[3][822] , \round_in[3][821] , \round_in[3][820] ,
         \round_in[3][819] , \round_in[3][818] , \round_in[3][817] ,
         \round_in[3][816] , \round_in[3][815] , \round_in[3][814] ,
         \round_in[3][813] , \round_in[3][812] , \round_in[3][811] ,
         \round_in[3][810] , \round_in[3][809] , \round_in[3][808] ,
         \round_in[3][807] , \round_in[3][806] , \round_in[3][805] ,
         \round_in[3][804] , \round_in[3][803] , \round_in[3][802] ,
         \round_in[3][801] , \round_in[3][800] , \round_in[3][799] ,
         \round_in[3][798] , \round_in[3][797] , \round_in[3][796] ,
         \round_in[3][795] , \round_in[3][794] , \round_in[3][793] ,
         \round_in[3][792] , \round_in[3][791] , \round_in[3][790] ,
         \round_in[3][789] , \round_in[3][788] , \round_in[3][787] ,
         \round_in[3][786] , \round_in[3][785] , \round_in[3][784] ,
         \round_in[3][783] , \round_in[3][782] , \round_in[3][781] ,
         \round_in[3][780] , \round_in[3][779] , \round_in[3][778] ,
         \round_in[3][777] , \round_in[3][776] , \round_in[3][775] ,
         \round_in[3][774] , \round_in[3][773] , \round_in[3][772] ,
         \round_in[3][771] , \round_in[3][770] , \round_in[3][769] ,
         \round_in[3][768] , \round_in[3][767] , \round_in[3][766] ,
         \round_in[3][765] , \round_in[3][764] , \round_in[3][763] ,
         \round_in[3][762] , \round_in[3][761] , \round_in[3][760] ,
         \round_in[3][759] , \round_in[3][758] , \round_in[3][757] ,
         \round_in[3][756] , \round_in[3][755] , \round_in[3][754] ,
         \round_in[3][753] , \round_in[3][752] , \round_in[3][751] ,
         \round_in[3][750] , \round_in[3][749] , \round_in[3][748] ,
         \round_in[3][747] , \round_in[3][746] , \round_in[3][745] ,
         \round_in[3][744] , \round_in[3][743] , \round_in[3][742] ,
         \round_in[3][741] , \round_in[3][740] , \round_in[3][739] ,
         \round_in[3][738] , \round_in[3][737] , \round_in[3][736] ,
         \round_in[3][735] , \round_in[3][734] , \round_in[3][733] ,
         \round_in[3][732] , \round_in[3][731] , \round_in[3][730] ,
         \round_in[3][729] , \round_in[3][728] , \round_in[3][727] ,
         \round_in[3][726] , \round_in[3][725] , \round_in[3][724] ,
         \round_in[3][723] , \round_in[3][722] , \round_in[3][721] ,
         \round_in[3][720] , \round_in[3][719] , \round_in[3][718] ,
         \round_in[3][717] , \round_in[3][716] , \round_in[3][715] ,
         \round_in[3][714] , \round_in[3][713] , \round_in[3][712] ,
         \round_in[3][711] , \round_in[3][710] , \round_in[3][709] ,
         \round_in[3][708] , \round_in[3][707] , \round_in[3][706] ,
         \round_in[3][705] , \round_in[3][704] , \round_in[3][703] ,
         \round_in[3][702] , \round_in[3][701] , \round_in[3][700] ,
         \round_in[3][699] , \round_in[3][698] , \round_in[3][697] ,
         \round_in[3][696] , \round_in[3][695] , \round_in[3][694] ,
         \round_in[3][693] , \round_in[3][692] , \round_in[3][691] ,
         \round_in[3][690] , \round_in[3][689] , \round_in[3][688] ,
         \round_in[3][687] , \round_in[3][686] , \round_in[3][685] ,
         \round_in[3][684] , \round_in[3][683] , \round_in[3][682] ,
         \round_in[3][681] , \round_in[3][680] , \round_in[3][679] ,
         \round_in[3][678] , \round_in[3][677] , \round_in[3][676] ,
         \round_in[3][675] , \round_in[3][674] , \round_in[3][673] ,
         \round_in[3][672] , \round_in[3][671] , \round_in[3][670] ,
         \round_in[3][669] , \round_in[3][668] , \round_in[3][667] ,
         \round_in[3][666] , \round_in[3][665] , \round_in[3][664] ,
         \round_in[3][663] , \round_in[3][662] , \round_in[3][661] ,
         \round_in[3][660] , \round_in[3][659] , \round_in[3][658] ,
         \round_in[3][657] , \round_in[3][656] , \round_in[3][655] ,
         \round_in[3][654] , \round_in[3][653] , \round_in[3][652] ,
         \round_in[3][651] , \round_in[3][650] , \round_in[3][649] ,
         \round_in[3][648] , \round_in[3][647] , \round_in[3][646] ,
         \round_in[3][645] , \round_in[3][644] , \round_in[3][643] ,
         \round_in[3][642] , \round_in[3][641] , \round_in[3][640] ,
         \round_in[3][639] , \round_in[3][638] , \round_in[3][637] ,
         \round_in[3][636] , \round_in[3][635] , \round_in[3][634] ,
         \round_in[3][633] , \round_in[3][632] , \round_in[3][631] ,
         \round_in[3][630] , \round_in[3][629] , \round_in[3][628] ,
         \round_in[3][627] , \round_in[3][626] , \round_in[3][625] ,
         \round_in[3][624] , \round_in[3][623] , \round_in[3][622] ,
         \round_in[3][621] , \round_in[3][620] , \round_in[3][619] ,
         \round_in[3][618] , \round_in[3][617] , \round_in[3][616] ,
         \round_in[3][615] , \round_in[3][614] , \round_in[3][613] ,
         \round_in[3][612] , \round_in[3][611] , \round_in[3][610] ,
         \round_in[3][609] , \round_in[3][608] , \round_in[3][607] ,
         \round_in[3][606] , \round_in[3][605] , \round_in[3][604] ,
         \round_in[3][603] , \round_in[3][602] , \round_in[3][601] ,
         \round_in[3][600] , \round_in[3][599] , \round_in[3][598] ,
         \round_in[3][597] , \round_in[3][596] , \round_in[3][595] ,
         \round_in[3][594] , \round_in[3][593] , \round_in[3][592] ,
         \round_in[3][591] , \round_in[3][590] , \round_in[3][589] ,
         \round_in[3][588] , \round_in[3][587] , \round_in[3][586] ,
         \round_in[3][585] , \round_in[3][584] , \round_in[3][583] ,
         \round_in[3][582] , \round_in[3][581] , \round_in[3][580] ,
         \round_in[3][579] , \round_in[3][578] , \round_in[3][577] ,
         \round_in[3][576] , \round_in[3][575] , \round_in[3][574] ,
         \round_in[3][573] , \round_in[3][572] , \round_in[3][571] ,
         \round_in[3][570] , \round_in[3][569] , \round_in[3][568] ,
         \round_in[3][567] , \round_in[3][566] , \round_in[3][565] ,
         \round_in[3][564] , \round_in[3][563] , \round_in[3][562] ,
         \round_in[3][561] , \round_in[3][560] , \round_in[3][559] ,
         \round_in[3][558] , \round_in[3][557] , \round_in[3][556] ,
         \round_in[3][555] , \round_in[3][554] , \round_in[3][553] ,
         \round_in[3][552] , \round_in[3][551] , \round_in[3][550] ,
         \round_in[3][549] , \round_in[3][548] , \round_in[3][547] ,
         \round_in[3][546] , \round_in[3][545] , \round_in[3][544] ,
         \round_in[3][543] , \round_in[3][542] , \round_in[3][541] ,
         \round_in[3][540] , \round_in[3][539] , \round_in[3][538] ,
         \round_in[3][537] , \round_in[3][536] , \round_in[3][535] ,
         \round_in[3][534] , \round_in[3][533] , \round_in[3][532] ,
         \round_in[3][531] , \round_in[3][530] , \round_in[3][529] ,
         \round_in[3][528] , \round_in[3][527] , \round_in[3][526] ,
         \round_in[3][525] , \round_in[3][524] , \round_in[3][523] ,
         \round_in[3][522] , \round_in[3][521] , \round_in[3][520] ,
         \round_in[3][519] , \round_in[3][518] , \round_in[3][517] ,
         \round_in[3][516] , \round_in[3][515] , \round_in[3][514] ,
         \round_in[3][513] , \round_in[3][512] , \round_in[3][511] ,
         \round_in[3][510] , \round_in[3][509] , \round_in[3][508] ,
         \round_in[3][507] , \round_in[3][506] , \round_in[3][505] ,
         \round_in[3][504] , \round_in[3][503] , \round_in[3][502] ,
         \round_in[3][501] , \round_in[3][500] , \round_in[3][499] ,
         \round_in[3][498] , \round_in[3][497] , \round_in[3][496] ,
         \round_in[3][495] , \round_in[3][494] , \round_in[3][493] ,
         \round_in[3][492] , \round_in[3][491] , \round_in[3][490] ,
         \round_in[3][489] , \round_in[3][488] , \round_in[3][487] ,
         \round_in[3][486] , \round_in[3][485] , \round_in[3][484] ,
         \round_in[3][483] , \round_in[3][482] , \round_in[3][481] ,
         \round_in[3][480] , \round_in[3][479] , \round_in[3][478] ,
         \round_in[3][477] , \round_in[3][476] , \round_in[3][475] ,
         \round_in[3][474] , \round_in[3][473] , \round_in[3][472] ,
         \round_in[3][471] , \round_in[3][470] , \round_in[3][469] ,
         \round_in[3][468] , \round_in[3][467] , \round_in[3][466] ,
         \round_in[3][465] , \round_in[3][464] , \round_in[3][463] ,
         \round_in[3][462] , \round_in[3][461] , \round_in[3][460] ,
         \round_in[3][459] , \round_in[3][458] , \round_in[3][457] ,
         \round_in[3][456] , \round_in[3][455] , \round_in[3][454] ,
         \round_in[3][453] , \round_in[3][452] , \round_in[3][451] ,
         \round_in[3][450] , \round_in[3][449] , \round_in[3][448] ,
         \round_in[3][447] , \round_in[3][446] , \round_in[3][445] ,
         \round_in[3][444] , \round_in[3][443] , \round_in[3][442] ,
         \round_in[3][441] , \round_in[3][440] , \round_in[3][439] ,
         \round_in[3][438] , \round_in[3][437] , \round_in[3][436] ,
         \round_in[3][435] , \round_in[3][434] , \round_in[3][433] ,
         \round_in[3][432] , \round_in[3][431] , \round_in[3][430] ,
         \round_in[3][429] , \round_in[3][428] , \round_in[3][427] ,
         \round_in[3][426] , \round_in[3][425] , \round_in[3][424] ,
         \round_in[3][423] , \round_in[3][422] , \round_in[3][421] ,
         \round_in[3][420] , \round_in[3][419] , \round_in[3][418] ,
         \round_in[3][417] , \round_in[3][416] , \round_in[3][415] ,
         \round_in[3][414] , \round_in[3][413] , \round_in[3][412] ,
         \round_in[3][411] , \round_in[3][410] , \round_in[3][409] ,
         \round_in[3][408] , \round_in[3][407] , \round_in[3][406] ,
         \round_in[3][405] , \round_in[3][404] , \round_in[3][403] ,
         \round_in[3][402] , \round_in[3][401] , \round_in[3][400] ,
         \round_in[3][399] , \round_in[3][398] , \round_in[3][397] ,
         \round_in[3][396] , \round_in[3][395] , \round_in[3][394] ,
         \round_in[3][393] , \round_in[3][392] , \round_in[3][391] ,
         \round_in[3][390] , \round_in[3][389] , \round_in[3][388] ,
         \round_in[3][387] , \round_in[3][386] , \round_in[3][385] ,
         \round_in[3][384] , \round_in[3][383] , \round_in[3][382] ,
         \round_in[3][381] , \round_in[3][380] , \round_in[3][379] ,
         \round_in[3][378] , \round_in[3][377] , \round_in[3][376] ,
         \round_in[3][375] , \round_in[3][374] , \round_in[3][373] ,
         \round_in[3][372] , \round_in[3][371] , \round_in[3][370] ,
         \round_in[3][369] , \round_in[3][368] , \round_in[3][367] ,
         \round_in[3][366] , \round_in[3][365] , \round_in[3][364] ,
         \round_in[3][363] , \round_in[3][362] , \round_in[3][361] ,
         \round_in[3][360] , \round_in[3][359] , \round_in[3][358] ,
         \round_in[3][357] , \round_in[3][356] , \round_in[3][355] ,
         \round_in[3][354] , \round_in[3][353] , \round_in[3][352] ,
         \round_in[3][351] , \round_in[3][350] , \round_in[3][349] ,
         \round_in[3][348] , \round_in[3][347] , \round_in[3][346] ,
         \round_in[3][345] , \round_in[3][344] , \round_in[3][343] ,
         \round_in[3][342] , \round_in[3][341] , \round_in[3][340] ,
         \round_in[3][339] , \round_in[3][338] , \round_in[3][337] ,
         \round_in[3][336] , \round_in[3][335] , \round_in[3][334] ,
         \round_in[3][333] , \round_in[3][332] , \round_in[3][331] ,
         \round_in[3][330] , \round_in[3][329] , \round_in[3][328] ,
         \round_in[3][327] , \round_in[3][326] , \round_in[3][325] ,
         \round_in[3][324] , \round_in[3][323] , \round_in[3][322] ,
         \round_in[3][321] , \round_in[3][320] , \round_in[3][319] ,
         \round_in[3][318] , \round_in[3][317] , \round_in[3][316] ,
         \round_in[3][315] , \round_in[3][314] , \round_in[3][313] ,
         \round_in[3][312] , \round_in[3][311] , \round_in[3][310] ,
         \round_in[3][309] , \round_in[3][308] , \round_in[3][307] ,
         \round_in[3][306] , \round_in[3][305] , \round_in[3][304] ,
         \round_in[3][303] , \round_in[3][302] , \round_in[3][301] ,
         \round_in[3][300] , \round_in[3][299] , \round_in[3][298] ,
         \round_in[3][297] , \round_in[3][296] , \round_in[3][295] ,
         \round_in[3][294] , \round_in[3][293] , \round_in[3][292] ,
         \round_in[3][291] , \round_in[3][290] , \round_in[3][289] ,
         \round_in[3][288] , \round_in[3][287] , \round_in[3][286] ,
         \round_in[3][285] , \round_in[3][284] , \round_in[3][283] ,
         \round_in[3][282] , \round_in[3][281] , \round_in[3][280] ,
         \round_in[3][279] , \round_in[3][278] , \round_in[3][277] ,
         \round_in[3][276] , \round_in[3][275] , \round_in[3][274] ,
         \round_in[3][273] , \round_in[3][272] , \round_in[3][271] ,
         \round_in[3][270] , \round_in[3][269] , \round_in[3][268] ,
         \round_in[3][267] , \round_in[3][266] , \round_in[3][265] ,
         \round_in[3][264] , \round_in[3][263] , \round_in[3][262] ,
         \round_in[3][261] , \round_in[3][260] , \round_in[3][259] ,
         \round_in[3][258] , \round_in[3][257] , \round_in[3][256] ,
         \round_in[3][255] , \round_in[3][254] , \round_in[3][253] ,
         \round_in[3][252] , \round_in[3][251] , \round_in[3][250] ,
         \round_in[3][249] , \round_in[3][248] , \round_in[3][247] ,
         \round_in[3][246] , \round_in[3][245] , \round_in[3][244] ,
         \round_in[3][243] , \round_in[3][242] , \round_in[3][241] ,
         \round_in[3][240] , \round_in[3][239] , \round_in[3][238] ,
         \round_in[3][237] , \round_in[3][236] , \round_in[3][235] ,
         \round_in[3][234] , \round_in[3][233] , \round_in[3][232] ,
         \round_in[3][231] , \round_in[3][230] , \round_in[3][229] ,
         \round_in[3][228] , \round_in[3][227] , \round_in[3][226] ,
         \round_in[3][225] , \round_in[3][224] , \round_in[3][223] ,
         \round_in[3][222] , \round_in[3][221] , \round_in[3][220] ,
         \round_in[3][219] , \round_in[3][218] , \round_in[3][217] ,
         \round_in[3][216] , \round_in[3][215] , \round_in[3][214] ,
         \round_in[3][213] , \round_in[3][212] , \round_in[3][211] ,
         \round_in[3][210] , \round_in[3][209] , \round_in[3][208] ,
         \round_in[3][207] , \round_in[3][206] , \round_in[3][205] ,
         \round_in[3][204] , \round_in[3][203] , \round_in[3][202] ,
         \round_in[3][201] , \round_in[3][200] , \round_in[3][199] ,
         \round_in[3][198] , \round_in[3][197] , \round_in[3][196] ,
         \round_in[3][195] , \round_in[3][194] , \round_in[3][193] ,
         \round_in[3][192] , \round_in[3][191] , \round_in[3][190] ,
         \round_in[3][189] , \round_in[3][188] , \round_in[3][187] ,
         \round_in[3][186] , \round_in[3][185] , \round_in[3][184] ,
         \round_in[3][183] , \round_in[3][182] , \round_in[3][181] ,
         \round_in[3][180] , \round_in[3][179] , \round_in[3][178] ,
         \round_in[3][177] , \round_in[3][176] , \round_in[3][175] ,
         \round_in[3][174] , \round_in[3][173] , \round_in[3][172] ,
         \round_in[3][171] , \round_in[3][170] , \round_in[3][169] ,
         \round_in[3][168] , \round_in[3][167] , \round_in[3][166] ,
         \round_in[3][165] , \round_in[3][164] , \round_in[3][163] ,
         \round_in[3][162] , \round_in[3][161] , \round_in[3][160] ,
         \round_in[3][159] , \round_in[3][158] , \round_in[3][157] ,
         \round_in[3][156] , \round_in[3][155] , \round_in[3][154] ,
         \round_in[3][153] , \round_in[3][152] , \round_in[3][151] ,
         \round_in[3][150] , \round_in[3][149] , \round_in[3][148] ,
         \round_in[3][147] , \round_in[3][146] , \round_in[3][145] ,
         \round_in[3][144] , \round_in[3][143] , \round_in[3][142] ,
         \round_in[3][141] , \round_in[3][140] , \round_in[3][139] ,
         \round_in[3][138] , \round_in[3][137] , \round_in[3][136] ,
         \round_in[3][135] , \round_in[3][134] , \round_in[3][133] ,
         \round_in[3][132] , \round_in[3][131] , \round_in[3][130] ,
         \round_in[3][129] , \round_in[3][128] , \round_in[3][127] ,
         \round_in[3][126] , \round_in[3][125] , \round_in[3][124] ,
         \round_in[3][123] , \round_in[3][122] , \round_in[3][121] ,
         \round_in[3][120] , \round_in[3][119] , \round_in[3][118] ,
         \round_in[3][117] , \round_in[3][116] , \round_in[3][115] ,
         \round_in[3][114] , \round_in[3][113] , \round_in[3][112] ,
         \round_in[3][111] , \round_in[3][110] , \round_in[3][109] ,
         \round_in[3][108] , \round_in[3][107] , \round_in[3][106] ,
         \round_in[3][105] , \round_in[3][104] , \round_in[3][103] ,
         \round_in[3][102] , \round_in[3][101] , \round_in[3][100] ,
         \round_in[3][99] , \round_in[3][98] , \round_in[3][97] ,
         \round_in[3][96] , \round_in[3][95] , \round_in[3][94] ,
         \round_in[3][93] , \round_in[3][92] , \round_in[3][91] ,
         \round_in[3][90] , \round_in[3][89] , \round_in[3][88] ,
         \round_in[3][87] , \round_in[3][86] , \round_in[3][85] ,
         \round_in[3][84] , \round_in[3][83] , \round_in[3][82] ,
         \round_in[3][81] , \round_in[3][80] , \round_in[3][79] ,
         \round_in[3][78] , \round_in[3][77] , \round_in[3][76] ,
         \round_in[3][75] , \round_in[3][74] , \round_in[3][73] ,
         \round_in[3][72] , \round_in[3][71] , \round_in[3][70] ,
         \round_in[3][69] , \round_in[3][68] , \round_in[3][67] ,
         \round_in[3][66] , \round_in[3][65] , \round_in[3][64] ,
         \round_in[3][63] , \round_in[3][62] , \round_in[3][61] ,
         \round_in[3][60] , \round_in[3][59] , \round_in[3][58] ,
         \round_in[3][57] , \round_in[3][56] , \round_in[3][55] ,
         \round_in[3][54] , \round_in[3][53] , \round_in[3][52] ,
         \round_in[3][51] , \round_in[3][50] , \round_in[3][49] ,
         \round_in[3][48] , \round_in[3][47] , \round_in[3][46] ,
         \round_in[3][45] , \round_in[3][44] , \round_in[3][43] ,
         \round_in[3][42] , \round_in[3][41] , \round_in[3][40] ,
         \round_in[3][39] , \round_in[3][38] , \round_in[3][37] ,
         \round_in[3][36] , \round_in[3][35] , \round_in[3][34] ,
         \round_in[3][33] , \round_in[3][32] , \round_in[3][31] ,
         \round_in[3][30] , \round_in[3][29] , \round_in[3][28] ,
         \round_in[3][27] , \round_in[3][26] , \round_in[3][25] ,
         \round_in[3][24] , \round_in[3][23] , \round_in[3][22] ,
         \round_in[3][21] , \round_in[3][20] , \round_in[3][19] ,
         \round_in[3][18] , \round_in[3][17] , \round_in[3][16] ,
         \round_in[3][15] , \round_in[3][14] , \round_in[3][13] ,
         \round_in[3][12] , \round_in[3][11] , \round_in[3][10] ,
         \round_in[3][9] , \round_in[3][8] , \round_in[3][7] ,
         \round_in[3][6] , \round_in[3][5] , \round_in[3][4] ,
         \round_in[3][3] , \round_in[3][2] , \round_in[3][1] ,
         \round_in[3][0] , \round_in[2][1599] , \round_in[2][1598] ,
         \round_in[2][1597] , \round_in[2][1596] , \round_in[2][1595] ,
         \round_in[2][1594] , \round_in[2][1593] , \round_in[2][1592] ,
         \round_in[2][1591] , \round_in[2][1590] , \round_in[2][1589] ,
         \round_in[2][1588] , \round_in[2][1587] , \round_in[2][1586] ,
         \round_in[2][1585] , \round_in[2][1584] , \round_in[2][1583] ,
         \round_in[2][1582] , \round_in[2][1581] , \round_in[2][1580] ,
         \round_in[2][1579] , \round_in[2][1578] , \round_in[2][1577] ,
         \round_in[2][1576] , \round_in[2][1575] , \round_in[2][1574] ,
         \round_in[2][1573] , \round_in[2][1572] , \round_in[2][1571] ,
         \round_in[2][1570] , \round_in[2][1569] , \round_in[2][1568] ,
         \round_in[2][1567] , \round_in[2][1566] , \round_in[2][1565] ,
         \round_in[2][1564] , \round_in[2][1563] , \round_in[2][1562] ,
         \round_in[2][1561] , \round_in[2][1560] , \round_in[2][1559] ,
         \round_in[2][1558] , \round_in[2][1557] , \round_in[2][1556] ,
         \round_in[2][1555] , \round_in[2][1554] , \round_in[2][1553] ,
         \round_in[2][1552] , \round_in[2][1551] , \round_in[2][1550] ,
         \round_in[2][1549] , \round_in[2][1548] , \round_in[2][1547] ,
         \round_in[2][1546] , \round_in[2][1545] , \round_in[2][1544] ,
         \round_in[2][1543] , \round_in[2][1542] , \round_in[2][1541] ,
         \round_in[2][1540] , \round_in[2][1539] , \round_in[2][1538] ,
         \round_in[2][1537] , \round_in[2][1536] , \round_in[2][1535] ,
         \round_in[2][1534] , \round_in[2][1533] , \round_in[2][1532] ,
         \round_in[2][1531] , \round_in[2][1530] , \round_in[2][1529] ,
         \round_in[2][1528] , \round_in[2][1527] , \round_in[2][1526] ,
         \round_in[2][1525] , \round_in[2][1524] , \round_in[2][1523] ,
         \round_in[2][1522] , \round_in[2][1521] , \round_in[2][1520] ,
         \round_in[2][1519] , \round_in[2][1518] , \round_in[2][1517] ,
         \round_in[2][1516] , \round_in[2][1515] , \round_in[2][1514] ,
         \round_in[2][1513] , \round_in[2][1512] , \round_in[2][1511] ,
         \round_in[2][1510] , \round_in[2][1509] , \round_in[2][1508] ,
         \round_in[2][1507] , \round_in[2][1506] , \round_in[2][1505] ,
         \round_in[2][1504] , \round_in[2][1503] , \round_in[2][1502] ,
         \round_in[2][1501] , \round_in[2][1500] , \round_in[2][1499] ,
         \round_in[2][1498] , \round_in[2][1497] , \round_in[2][1496] ,
         \round_in[2][1495] , \round_in[2][1494] , \round_in[2][1493] ,
         \round_in[2][1492] , \round_in[2][1491] , \round_in[2][1490] ,
         \round_in[2][1489] , \round_in[2][1488] , \round_in[2][1487] ,
         \round_in[2][1486] , \round_in[2][1485] , \round_in[2][1484] ,
         \round_in[2][1483] , \round_in[2][1482] , \round_in[2][1481] ,
         \round_in[2][1480] , \round_in[2][1479] , \round_in[2][1478] ,
         \round_in[2][1477] , \round_in[2][1476] , \round_in[2][1475] ,
         \round_in[2][1474] , \round_in[2][1473] , \round_in[2][1472] ,
         \round_in[2][1471] , \round_in[2][1470] , \round_in[2][1469] ,
         \round_in[2][1468] , \round_in[2][1467] , \round_in[2][1466] ,
         \round_in[2][1465] , \round_in[2][1464] , \round_in[2][1463] ,
         \round_in[2][1462] , \round_in[2][1461] , \round_in[2][1460] ,
         \round_in[2][1459] , \round_in[2][1458] , \round_in[2][1457] ,
         \round_in[2][1456] , \round_in[2][1455] , \round_in[2][1454] ,
         \round_in[2][1453] , \round_in[2][1452] , \round_in[2][1451] ,
         \round_in[2][1450] , \round_in[2][1449] , \round_in[2][1448] ,
         \round_in[2][1447] , \round_in[2][1446] , \round_in[2][1445] ,
         \round_in[2][1444] , \round_in[2][1443] , \round_in[2][1442] ,
         \round_in[2][1441] , \round_in[2][1440] , \round_in[2][1439] ,
         \round_in[2][1438] , \round_in[2][1437] , \round_in[2][1436] ,
         \round_in[2][1435] , \round_in[2][1434] , \round_in[2][1433] ,
         \round_in[2][1432] , \round_in[2][1431] , \round_in[2][1430] ,
         \round_in[2][1429] , \round_in[2][1428] , \round_in[2][1427] ,
         \round_in[2][1426] , \round_in[2][1425] , \round_in[2][1424] ,
         \round_in[2][1423] , \round_in[2][1422] , \round_in[2][1421] ,
         \round_in[2][1420] , \round_in[2][1419] , \round_in[2][1418] ,
         \round_in[2][1417] , \round_in[2][1416] , \round_in[2][1415] ,
         \round_in[2][1414] , \round_in[2][1413] , \round_in[2][1412] ,
         \round_in[2][1411] , \round_in[2][1410] , \round_in[2][1409] ,
         \round_in[2][1408] , \round_in[2][1407] , \round_in[2][1406] ,
         \round_in[2][1405] , \round_in[2][1404] , \round_in[2][1403] ,
         \round_in[2][1402] , \round_in[2][1401] , \round_in[2][1400] ,
         \round_in[2][1399] , \round_in[2][1398] , \round_in[2][1397] ,
         \round_in[2][1396] , \round_in[2][1395] , \round_in[2][1394] ,
         \round_in[2][1393] , \round_in[2][1392] , \round_in[2][1391] ,
         \round_in[2][1390] , \round_in[2][1389] , \round_in[2][1388] ,
         \round_in[2][1387] , \round_in[2][1386] , \round_in[2][1385] ,
         \round_in[2][1384] , \round_in[2][1383] , \round_in[2][1382] ,
         \round_in[2][1381] , \round_in[2][1380] , \round_in[2][1379] ,
         \round_in[2][1378] , \round_in[2][1377] , \round_in[2][1376] ,
         \round_in[2][1375] , \round_in[2][1374] , \round_in[2][1373] ,
         \round_in[2][1372] , \round_in[2][1371] , \round_in[2][1370] ,
         \round_in[2][1369] , \round_in[2][1368] , \round_in[2][1367] ,
         \round_in[2][1366] , \round_in[2][1365] , \round_in[2][1364] ,
         \round_in[2][1363] , \round_in[2][1362] , \round_in[2][1361] ,
         \round_in[2][1360] , \round_in[2][1359] , \round_in[2][1358] ,
         \round_in[2][1357] , \round_in[2][1356] , \round_in[2][1355] ,
         \round_in[2][1354] , \round_in[2][1353] , \round_in[2][1352] ,
         \round_in[2][1351] , \round_in[2][1350] , \round_in[2][1349] ,
         \round_in[2][1348] , \round_in[2][1347] , \round_in[2][1346] ,
         \round_in[2][1345] , \round_in[2][1344] , \round_in[2][1343] ,
         \round_in[2][1342] , \round_in[2][1341] , \round_in[2][1340] ,
         \round_in[2][1339] , \round_in[2][1338] , \round_in[2][1337] ,
         \round_in[2][1336] , \round_in[2][1335] , \round_in[2][1334] ,
         \round_in[2][1333] , \round_in[2][1332] , \round_in[2][1331] ,
         \round_in[2][1330] , \round_in[2][1329] , \round_in[2][1328] ,
         \round_in[2][1327] , \round_in[2][1326] , \round_in[2][1325] ,
         \round_in[2][1324] , \round_in[2][1323] , \round_in[2][1322] ,
         \round_in[2][1321] , \round_in[2][1320] , \round_in[2][1319] ,
         \round_in[2][1318] , \round_in[2][1317] , \round_in[2][1316] ,
         \round_in[2][1315] , \round_in[2][1314] , \round_in[2][1313] ,
         \round_in[2][1312] , \round_in[2][1311] , \round_in[2][1310] ,
         \round_in[2][1309] , \round_in[2][1308] , \round_in[2][1307] ,
         \round_in[2][1306] , \round_in[2][1305] , \round_in[2][1304] ,
         \round_in[2][1303] , \round_in[2][1302] , \round_in[2][1301] ,
         \round_in[2][1300] , \round_in[2][1299] , \round_in[2][1298] ,
         \round_in[2][1297] , \round_in[2][1296] , \round_in[2][1295] ,
         \round_in[2][1294] , \round_in[2][1293] , \round_in[2][1292] ,
         \round_in[2][1291] , \round_in[2][1290] , \round_in[2][1289] ,
         \round_in[2][1288] , \round_in[2][1287] , \round_in[2][1286] ,
         \round_in[2][1285] , \round_in[2][1284] , \round_in[2][1283] ,
         \round_in[2][1282] , \round_in[2][1281] , \round_in[2][1280] ,
         \round_in[2][1279] , \round_in[2][1278] , \round_in[2][1277] ,
         \round_in[2][1276] , \round_in[2][1275] , \round_in[2][1274] ,
         \round_in[2][1273] , \round_in[2][1272] , \round_in[2][1271] ,
         \round_in[2][1270] , \round_in[2][1269] , \round_in[2][1268] ,
         \round_in[2][1267] , \round_in[2][1266] , \round_in[2][1265] ,
         \round_in[2][1264] , \round_in[2][1263] , \round_in[2][1262] ,
         \round_in[2][1261] , \round_in[2][1260] , \round_in[2][1259] ,
         \round_in[2][1258] , \round_in[2][1257] , \round_in[2][1256] ,
         \round_in[2][1255] , \round_in[2][1254] , \round_in[2][1253] ,
         \round_in[2][1252] , \round_in[2][1251] , \round_in[2][1250] ,
         \round_in[2][1249] , \round_in[2][1248] , \round_in[2][1247] ,
         \round_in[2][1246] , \round_in[2][1245] , \round_in[2][1244] ,
         \round_in[2][1243] , \round_in[2][1242] , \round_in[2][1241] ,
         \round_in[2][1240] , \round_in[2][1239] , \round_in[2][1238] ,
         \round_in[2][1237] , \round_in[2][1236] , \round_in[2][1235] ,
         \round_in[2][1234] , \round_in[2][1233] , \round_in[2][1232] ,
         \round_in[2][1231] , \round_in[2][1230] , \round_in[2][1229] ,
         \round_in[2][1228] , \round_in[2][1227] , \round_in[2][1226] ,
         \round_in[2][1225] , \round_in[2][1224] , \round_in[2][1223] ,
         \round_in[2][1222] , \round_in[2][1221] , \round_in[2][1220] ,
         \round_in[2][1219] , \round_in[2][1218] , \round_in[2][1217] ,
         \round_in[2][1216] , \round_in[2][1215] , \round_in[2][1214] ,
         \round_in[2][1213] , \round_in[2][1212] , \round_in[2][1211] ,
         \round_in[2][1210] , \round_in[2][1209] , \round_in[2][1208] ,
         \round_in[2][1207] , \round_in[2][1206] , \round_in[2][1205] ,
         \round_in[2][1204] , \round_in[2][1203] , \round_in[2][1202] ,
         \round_in[2][1201] , \round_in[2][1200] , \round_in[2][1199] ,
         \round_in[2][1198] , \round_in[2][1197] , \round_in[2][1196] ,
         \round_in[2][1195] , \round_in[2][1194] , \round_in[2][1193] ,
         \round_in[2][1192] , \round_in[2][1191] , \round_in[2][1190] ,
         \round_in[2][1189] , \round_in[2][1188] , \round_in[2][1187] ,
         \round_in[2][1186] , \round_in[2][1185] , \round_in[2][1184] ,
         \round_in[2][1183] , \round_in[2][1182] , \round_in[2][1181] ,
         \round_in[2][1180] , \round_in[2][1179] , \round_in[2][1178] ,
         \round_in[2][1177] , \round_in[2][1176] , \round_in[2][1175] ,
         \round_in[2][1174] , \round_in[2][1173] , \round_in[2][1172] ,
         \round_in[2][1171] , \round_in[2][1170] , \round_in[2][1169] ,
         \round_in[2][1168] , \round_in[2][1167] , \round_in[2][1166] ,
         \round_in[2][1165] , \round_in[2][1164] , \round_in[2][1163] ,
         \round_in[2][1162] , \round_in[2][1161] , \round_in[2][1160] ,
         \round_in[2][1159] , \round_in[2][1158] , \round_in[2][1157] ,
         \round_in[2][1156] , \round_in[2][1155] , \round_in[2][1154] ,
         \round_in[2][1153] , \round_in[2][1152] , \round_in[2][1151] ,
         \round_in[2][1150] , \round_in[2][1149] , \round_in[2][1148] ,
         \round_in[2][1147] , \round_in[2][1146] , \round_in[2][1145] ,
         \round_in[2][1144] , \round_in[2][1143] , \round_in[2][1142] ,
         \round_in[2][1141] , \round_in[2][1140] , \round_in[2][1139] ,
         \round_in[2][1138] , \round_in[2][1137] , \round_in[2][1136] ,
         \round_in[2][1135] , \round_in[2][1134] , \round_in[2][1133] ,
         \round_in[2][1132] , \round_in[2][1131] , \round_in[2][1130] ,
         \round_in[2][1129] , \round_in[2][1128] , \round_in[2][1127] ,
         \round_in[2][1126] , \round_in[2][1125] , \round_in[2][1124] ,
         \round_in[2][1123] , \round_in[2][1122] , \round_in[2][1121] ,
         \round_in[2][1120] , \round_in[2][1119] , \round_in[2][1118] ,
         \round_in[2][1117] , \round_in[2][1116] , \round_in[2][1115] ,
         \round_in[2][1114] , \round_in[2][1113] , \round_in[2][1112] ,
         \round_in[2][1111] , \round_in[2][1110] , \round_in[2][1109] ,
         \round_in[2][1108] , \round_in[2][1107] , \round_in[2][1106] ,
         \round_in[2][1105] , \round_in[2][1104] , \round_in[2][1103] ,
         \round_in[2][1102] , \round_in[2][1101] , \round_in[2][1100] ,
         \round_in[2][1099] , \round_in[2][1098] , \round_in[2][1097] ,
         \round_in[2][1096] , \round_in[2][1095] , \round_in[2][1094] ,
         \round_in[2][1093] , \round_in[2][1092] , \round_in[2][1091] ,
         \round_in[2][1090] , \round_in[2][1089] , \round_in[2][1088] ,
         \round_in[2][1087] , \round_in[2][1086] , \round_in[2][1085] ,
         \round_in[2][1084] , \round_in[2][1083] , \round_in[2][1082] ,
         \round_in[2][1081] , \round_in[2][1080] , \round_in[2][1079] ,
         \round_in[2][1078] , \round_in[2][1077] , \round_in[2][1076] ,
         \round_in[2][1075] , \round_in[2][1074] , \round_in[2][1073] ,
         \round_in[2][1072] , \round_in[2][1071] , \round_in[2][1070] ,
         \round_in[2][1069] , \round_in[2][1068] , \round_in[2][1067] ,
         \round_in[2][1066] , \round_in[2][1065] , \round_in[2][1064] ,
         \round_in[2][1063] , \round_in[2][1062] , \round_in[2][1061] ,
         \round_in[2][1060] , \round_in[2][1059] , \round_in[2][1058] ,
         \round_in[2][1057] , \round_in[2][1056] , \round_in[2][1055] ,
         \round_in[2][1054] , \round_in[2][1053] , \round_in[2][1052] ,
         \round_in[2][1051] , \round_in[2][1050] , \round_in[2][1049] ,
         \round_in[2][1048] , \round_in[2][1047] , \round_in[2][1046] ,
         \round_in[2][1045] , \round_in[2][1044] , \round_in[2][1043] ,
         \round_in[2][1042] , \round_in[2][1041] , \round_in[2][1040] ,
         \round_in[2][1039] , \round_in[2][1038] , \round_in[2][1037] ,
         \round_in[2][1036] , \round_in[2][1035] , \round_in[2][1034] ,
         \round_in[2][1033] , \round_in[2][1032] , \round_in[2][1031] ,
         \round_in[2][1030] , \round_in[2][1029] , \round_in[2][1028] ,
         \round_in[2][1027] , \round_in[2][1026] , \round_in[2][1025] ,
         \round_in[2][1024] , \round_in[2][1023] , \round_in[2][1022] ,
         \round_in[2][1021] , \round_in[2][1020] , \round_in[2][1019] ,
         \round_in[2][1018] , \round_in[2][1017] , \round_in[2][1016] ,
         \round_in[2][1015] , \round_in[2][1014] , \round_in[2][1013] ,
         \round_in[2][1012] , \round_in[2][1011] , \round_in[2][1010] ,
         \round_in[2][1009] , \round_in[2][1008] , \round_in[2][1007] ,
         \round_in[2][1006] , \round_in[2][1005] , \round_in[2][1004] ,
         \round_in[2][1003] , \round_in[2][1002] , \round_in[2][1001] ,
         \round_in[2][1000] , \round_in[2][999] , \round_in[2][998] ,
         \round_in[2][997] , \round_in[2][996] , \round_in[2][995] ,
         \round_in[2][994] , \round_in[2][993] , \round_in[2][992] ,
         \round_in[2][991] , \round_in[2][990] , \round_in[2][989] ,
         \round_in[2][988] , \round_in[2][987] , \round_in[2][986] ,
         \round_in[2][985] , \round_in[2][984] , \round_in[2][983] ,
         \round_in[2][982] , \round_in[2][981] , \round_in[2][980] ,
         \round_in[2][979] , \round_in[2][978] , \round_in[2][977] ,
         \round_in[2][976] , \round_in[2][975] , \round_in[2][974] ,
         \round_in[2][973] , \round_in[2][972] , \round_in[2][971] ,
         \round_in[2][970] , \round_in[2][969] , \round_in[2][968] ,
         \round_in[2][967] , \round_in[2][966] , \round_in[2][965] ,
         \round_in[2][964] , \round_in[2][963] , \round_in[2][962] ,
         \round_in[2][961] , \round_in[2][960] , \round_in[2][959] ,
         \round_in[2][958] , \round_in[2][957] , \round_in[2][956] ,
         \round_in[2][955] , \round_in[2][954] , \round_in[2][953] ,
         \round_in[2][952] , \round_in[2][951] , \round_in[2][950] ,
         \round_in[2][949] , \round_in[2][948] , \round_in[2][947] ,
         \round_in[2][946] , \round_in[2][945] , \round_in[2][944] ,
         \round_in[2][943] , \round_in[2][942] , \round_in[2][941] ,
         \round_in[2][940] , \round_in[2][939] , \round_in[2][938] ,
         \round_in[2][937] , \round_in[2][936] , \round_in[2][935] ,
         \round_in[2][934] , \round_in[2][933] , \round_in[2][932] ,
         \round_in[2][931] , \round_in[2][930] , \round_in[2][929] ,
         \round_in[2][928] , \round_in[2][927] , \round_in[2][926] ,
         \round_in[2][925] , \round_in[2][924] , \round_in[2][923] ,
         \round_in[2][922] , \round_in[2][921] , \round_in[2][920] ,
         \round_in[2][919] , \round_in[2][918] , \round_in[2][917] ,
         \round_in[2][916] , \round_in[2][915] , \round_in[2][914] ,
         \round_in[2][913] , \round_in[2][912] , \round_in[2][911] ,
         \round_in[2][910] , \round_in[2][909] , \round_in[2][908] ,
         \round_in[2][907] , \round_in[2][906] , \round_in[2][905] ,
         \round_in[2][904] , \round_in[2][903] , \round_in[2][902] ,
         \round_in[2][901] , \round_in[2][900] , \round_in[2][899] ,
         \round_in[2][898] , \round_in[2][897] , \round_in[2][896] ,
         \round_in[2][895] , \round_in[2][894] , \round_in[2][893] ,
         \round_in[2][892] , \round_in[2][891] , \round_in[2][890] ,
         \round_in[2][889] , \round_in[2][888] , \round_in[2][887] ,
         \round_in[2][886] , \round_in[2][885] , \round_in[2][884] ,
         \round_in[2][883] , \round_in[2][882] , \round_in[2][881] ,
         \round_in[2][880] , \round_in[2][879] , \round_in[2][878] ,
         \round_in[2][877] , \round_in[2][876] , \round_in[2][875] ,
         \round_in[2][874] , \round_in[2][873] , \round_in[2][872] ,
         \round_in[2][871] , \round_in[2][870] , \round_in[2][869] ,
         \round_in[2][868] , \round_in[2][867] , \round_in[2][866] ,
         \round_in[2][865] , \round_in[2][864] , \round_in[2][863] ,
         \round_in[2][862] , \round_in[2][861] , \round_in[2][860] ,
         \round_in[2][859] , \round_in[2][858] , \round_in[2][857] ,
         \round_in[2][856] , \round_in[2][855] , \round_in[2][854] ,
         \round_in[2][853] , \round_in[2][852] , \round_in[2][851] ,
         \round_in[2][850] , \round_in[2][849] , \round_in[2][848] ,
         \round_in[2][847] , \round_in[2][846] , \round_in[2][845] ,
         \round_in[2][844] , \round_in[2][843] , \round_in[2][842] ,
         \round_in[2][841] , \round_in[2][840] , \round_in[2][839] ,
         \round_in[2][838] , \round_in[2][837] , \round_in[2][836] ,
         \round_in[2][835] , \round_in[2][834] , \round_in[2][833] ,
         \round_in[2][832] , \round_in[2][831] , \round_in[2][830] ,
         \round_in[2][829] , \round_in[2][828] , \round_in[2][827] ,
         \round_in[2][826] , \round_in[2][825] , \round_in[2][824] ,
         \round_in[2][823] , \round_in[2][822] , \round_in[2][821] ,
         \round_in[2][820] , \round_in[2][819] , \round_in[2][818] ,
         \round_in[2][817] , \round_in[2][816] , \round_in[2][815] ,
         \round_in[2][814] , \round_in[2][813] , \round_in[2][812] ,
         \round_in[2][811] , \round_in[2][810] , \round_in[2][809] ,
         \round_in[2][808] , \round_in[2][807] , \round_in[2][806] ,
         \round_in[2][805] , \round_in[2][804] , \round_in[2][803] ,
         \round_in[2][802] , \round_in[2][801] , \round_in[2][800] ,
         \round_in[2][799] , \round_in[2][798] , \round_in[2][797] ,
         \round_in[2][796] , \round_in[2][795] , \round_in[2][794] ,
         \round_in[2][793] , \round_in[2][792] , \round_in[2][791] ,
         \round_in[2][790] , \round_in[2][789] , \round_in[2][788] ,
         \round_in[2][787] , \round_in[2][786] , \round_in[2][785] ,
         \round_in[2][784] , \round_in[2][783] , \round_in[2][782] ,
         \round_in[2][781] , \round_in[2][780] , \round_in[2][779] ,
         \round_in[2][778] , \round_in[2][777] , \round_in[2][776] ,
         \round_in[2][775] , \round_in[2][774] , \round_in[2][773] ,
         \round_in[2][772] , \round_in[2][771] , \round_in[2][770] ,
         \round_in[2][769] , \round_in[2][768] , \round_in[2][767] ,
         \round_in[2][766] , \round_in[2][765] , \round_in[2][764] ,
         \round_in[2][763] , \round_in[2][762] , \round_in[2][761] ,
         \round_in[2][760] , \round_in[2][759] , \round_in[2][758] ,
         \round_in[2][757] , \round_in[2][756] , \round_in[2][755] ,
         \round_in[2][754] , \round_in[2][753] , \round_in[2][752] ,
         \round_in[2][751] , \round_in[2][750] , \round_in[2][749] ,
         \round_in[2][748] , \round_in[2][747] , \round_in[2][746] ,
         \round_in[2][745] , \round_in[2][744] , \round_in[2][743] ,
         \round_in[2][742] , \round_in[2][741] , \round_in[2][740] ,
         \round_in[2][739] , \round_in[2][738] , \round_in[2][737] ,
         \round_in[2][736] , \round_in[2][735] , \round_in[2][734] ,
         \round_in[2][733] , \round_in[2][732] , \round_in[2][731] ,
         \round_in[2][730] , \round_in[2][729] , \round_in[2][728] ,
         \round_in[2][727] , \round_in[2][726] , \round_in[2][725] ,
         \round_in[2][724] , \round_in[2][723] , \round_in[2][722] ,
         \round_in[2][721] , \round_in[2][720] , \round_in[2][719] ,
         \round_in[2][718] , \round_in[2][717] , \round_in[2][716] ,
         \round_in[2][715] , \round_in[2][714] , \round_in[2][713] ,
         \round_in[2][712] , \round_in[2][711] , \round_in[2][710] ,
         \round_in[2][709] , \round_in[2][708] , \round_in[2][707] ,
         \round_in[2][706] , \round_in[2][705] , \round_in[2][704] ,
         \round_in[2][703] , \round_in[2][702] , \round_in[2][701] ,
         \round_in[2][700] , \round_in[2][699] , \round_in[2][698] ,
         \round_in[2][697] , \round_in[2][696] , \round_in[2][695] ,
         \round_in[2][694] , \round_in[2][693] , \round_in[2][692] ,
         \round_in[2][691] , \round_in[2][690] , \round_in[2][689] ,
         \round_in[2][688] , \round_in[2][687] , \round_in[2][686] ,
         \round_in[2][685] , \round_in[2][684] , \round_in[2][683] ,
         \round_in[2][682] , \round_in[2][681] , \round_in[2][680] ,
         \round_in[2][679] , \round_in[2][678] , \round_in[2][677] ,
         \round_in[2][676] , \round_in[2][675] , \round_in[2][674] ,
         \round_in[2][673] , \round_in[2][672] , \round_in[2][671] ,
         \round_in[2][670] , \round_in[2][669] , \round_in[2][668] ,
         \round_in[2][667] , \round_in[2][666] , \round_in[2][665] ,
         \round_in[2][664] , \round_in[2][663] , \round_in[2][662] ,
         \round_in[2][661] , \round_in[2][660] , \round_in[2][659] ,
         \round_in[2][658] , \round_in[2][657] , \round_in[2][656] ,
         \round_in[2][655] , \round_in[2][654] , \round_in[2][653] ,
         \round_in[2][652] , \round_in[2][651] , \round_in[2][650] ,
         \round_in[2][649] , \round_in[2][648] , \round_in[2][647] ,
         \round_in[2][646] , \round_in[2][645] , \round_in[2][644] ,
         \round_in[2][643] , \round_in[2][642] , \round_in[2][641] ,
         \round_in[2][640] , \round_in[2][639] , \round_in[2][638] ,
         \round_in[2][637] , \round_in[2][636] , \round_in[2][635] ,
         \round_in[2][634] , \round_in[2][633] , \round_in[2][632] ,
         \round_in[2][631] , \round_in[2][630] , \round_in[2][629] ,
         \round_in[2][628] , \round_in[2][627] , \round_in[2][626] ,
         \round_in[2][625] , \round_in[2][624] , \round_in[2][623] ,
         \round_in[2][622] , \round_in[2][621] , \round_in[2][620] ,
         \round_in[2][619] , \round_in[2][618] , \round_in[2][617] ,
         \round_in[2][616] , \round_in[2][615] , \round_in[2][614] ,
         \round_in[2][613] , \round_in[2][612] , \round_in[2][611] ,
         \round_in[2][610] , \round_in[2][609] , \round_in[2][608] ,
         \round_in[2][607] , \round_in[2][606] , \round_in[2][605] ,
         \round_in[2][604] , \round_in[2][603] , \round_in[2][602] ,
         \round_in[2][601] , \round_in[2][600] , \round_in[2][599] ,
         \round_in[2][598] , \round_in[2][597] , \round_in[2][596] ,
         \round_in[2][595] , \round_in[2][594] , \round_in[2][593] ,
         \round_in[2][592] , \round_in[2][591] , \round_in[2][590] ,
         \round_in[2][589] , \round_in[2][588] , \round_in[2][587] ,
         \round_in[2][586] , \round_in[2][585] , \round_in[2][584] ,
         \round_in[2][583] , \round_in[2][582] , \round_in[2][581] ,
         \round_in[2][580] , \round_in[2][579] , \round_in[2][578] ,
         \round_in[2][577] , \round_in[2][576] , \round_in[2][575] ,
         \round_in[2][574] , \round_in[2][573] , \round_in[2][572] ,
         \round_in[2][571] , \round_in[2][570] , \round_in[2][569] ,
         \round_in[2][568] , \round_in[2][567] , \round_in[2][566] ,
         \round_in[2][565] , \round_in[2][564] , \round_in[2][563] ,
         \round_in[2][562] , \round_in[2][561] , \round_in[2][560] ,
         \round_in[2][559] , \round_in[2][558] , \round_in[2][557] ,
         \round_in[2][556] , \round_in[2][555] , \round_in[2][554] ,
         \round_in[2][553] , \round_in[2][552] , \round_in[2][551] ,
         \round_in[2][550] , \round_in[2][549] , \round_in[2][548] ,
         \round_in[2][547] , \round_in[2][546] , \round_in[2][545] ,
         \round_in[2][544] , \round_in[2][543] , \round_in[2][542] ,
         \round_in[2][541] , \round_in[2][540] , \round_in[2][539] ,
         \round_in[2][538] , \round_in[2][537] , \round_in[2][536] ,
         \round_in[2][535] , \round_in[2][534] , \round_in[2][533] ,
         \round_in[2][532] , \round_in[2][531] , \round_in[2][530] ,
         \round_in[2][529] , \round_in[2][528] , \round_in[2][527] ,
         \round_in[2][526] , \round_in[2][525] , \round_in[2][524] ,
         \round_in[2][523] , \round_in[2][522] , \round_in[2][521] ,
         \round_in[2][520] , \round_in[2][519] , \round_in[2][518] ,
         \round_in[2][517] , \round_in[2][516] , \round_in[2][515] ,
         \round_in[2][514] , \round_in[2][513] , \round_in[2][512] ,
         \round_in[2][511] , \round_in[2][510] , \round_in[2][509] ,
         \round_in[2][508] , \round_in[2][507] , \round_in[2][506] ,
         \round_in[2][505] , \round_in[2][504] , \round_in[2][503] ,
         \round_in[2][502] , \round_in[2][501] , \round_in[2][500] ,
         \round_in[2][499] , \round_in[2][498] , \round_in[2][497] ,
         \round_in[2][496] , \round_in[2][495] , \round_in[2][494] ,
         \round_in[2][493] , \round_in[2][492] , \round_in[2][491] ,
         \round_in[2][490] , \round_in[2][489] , \round_in[2][488] ,
         \round_in[2][487] , \round_in[2][486] , \round_in[2][485] ,
         \round_in[2][484] , \round_in[2][483] , \round_in[2][482] ,
         \round_in[2][481] , \round_in[2][480] , \round_in[2][479] ,
         \round_in[2][478] , \round_in[2][477] , \round_in[2][476] ,
         \round_in[2][475] , \round_in[2][474] , \round_in[2][473] ,
         \round_in[2][472] , \round_in[2][471] , \round_in[2][470] ,
         \round_in[2][469] , \round_in[2][468] , \round_in[2][467] ,
         \round_in[2][466] , \round_in[2][465] , \round_in[2][464] ,
         \round_in[2][463] , \round_in[2][462] , \round_in[2][461] ,
         \round_in[2][460] , \round_in[2][459] , \round_in[2][458] ,
         \round_in[2][457] , \round_in[2][456] , \round_in[2][455] ,
         \round_in[2][454] , \round_in[2][453] , \round_in[2][452] ,
         \round_in[2][451] , \round_in[2][450] , \round_in[2][449] ,
         \round_in[2][448] , \round_in[2][447] , \round_in[2][446] ,
         \round_in[2][445] , \round_in[2][444] , \round_in[2][443] ,
         \round_in[2][442] , \round_in[2][441] , \round_in[2][440] ,
         \round_in[2][439] , \round_in[2][438] , \round_in[2][437] ,
         \round_in[2][436] , \round_in[2][435] , \round_in[2][434] ,
         \round_in[2][433] , \round_in[2][432] , \round_in[2][431] ,
         \round_in[2][430] , \round_in[2][429] , \round_in[2][428] ,
         \round_in[2][427] , \round_in[2][426] , \round_in[2][425] ,
         \round_in[2][424] , \round_in[2][423] , \round_in[2][422] ,
         \round_in[2][421] , \round_in[2][420] , \round_in[2][419] ,
         \round_in[2][418] , \round_in[2][417] , \round_in[2][416] ,
         \round_in[2][415] , \round_in[2][414] , \round_in[2][413] ,
         \round_in[2][412] , \round_in[2][411] , \round_in[2][410] ,
         \round_in[2][409] , \round_in[2][408] , \round_in[2][407] ,
         \round_in[2][406] , \round_in[2][405] , \round_in[2][404] ,
         \round_in[2][403] , \round_in[2][402] , \round_in[2][401] ,
         \round_in[2][400] , \round_in[2][399] , \round_in[2][398] ,
         \round_in[2][397] , \round_in[2][396] , \round_in[2][395] ,
         \round_in[2][394] , \round_in[2][393] , \round_in[2][392] ,
         \round_in[2][391] , \round_in[2][390] , \round_in[2][389] ,
         \round_in[2][388] , \round_in[2][387] , \round_in[2][386] ,
         \round_in[2][385] , \round_in[2][384] , \round_in[2][383] ,
         \round_in[2][382] , \round_in[2][381] , \round_in[2][380] ,
         \round_in[2][379] , \round_in[2][378] , \round_in[2][377] ,
         \round_in[2][376] , \round_in[2][375] , \round_in[2][374] ,
         \round_in[2][373] , \round_in[2][372] , \round_in[2][371] ,
         \round_in[2][370] , \round_in[2][369] , \round_in[2][368] ,
         \round_in[2][367] , \round_in[2][366] , \round_in[2][365] ,
         \round_in[2][364] , \round_in[2][363] , \round_in[2][362] ,
         \round_in[2][361] , \round_in[2][360] , \round_in[2][359] ,
         \round_in[2][358] , \round_in[2][357] , \round_in[2][356] ,
         \round_in[2][355] , \round_in[2][354] , \round_in[2][353] ,
         \round_in[2][352] , \round_in[2][351] , \round_in[2][350] ,
         \round_in[2][349] , \round_in[2][348] , \round_in[2][347] ,
         \round_in[2][346] , \round_in[2][345] , \round_in[2][344] ,
         \round_in[2][343] , \round_in[2][342] , \round_in[2][341] ,
         \round_in[2][340] , \round_in[2][339] , \round_in[2][338] ,
         \round_in[2][337] , \round_in[2][336] , \round_in[2][335] ,
         \round_in[2][334] , \round_in[2][333] , \round_in[2][332] ,
         \round_in[2][331] , \round_in[2][330] , \round_in[2][329] ,
         \round_in[2][328] , \round_in[2][327] , \round_in[2][326] ,
         \round_in[2][325] , \round_in[2][324] , \round_in[2][323] ,
         \round_in[2][322] , \round_in[2][321] , \round_in[2][320] ,
         \round_in[2][319] , \round_in[2][318] , \round_in[2][317] ,
         \round_in[2][316] , \round_in[2][315] , \round_in[2][314] ,
         \round_in[2][313] , \round_in[2][312] , \round_in[2][311] ,
         \round_in[2][310] , \round_in[2][309] , \round_in[2][308] ,
         \round_in[2][307] , \round_in[2][306] , \round_in[2][305] ,
         \round_in[2][304] , \round_in[2][303] , \round_in[2][302] ,
         \round_in[2][301] , \round_in[2][300] , \round_in[2][299] ,
         \round_in[2][298] , \round_in[2][297] , \round_in[2][296] ,
         \round_in[2][295] , \round_in[2][294] , \round_in[2][293] ,
         \round_in[2][292] , \round_in[2][291] , \round_in[2][290] ,
         \round_in[2][289] , \round_in[2][288] , \round_in[2][287] ,
         \round_in[2][286] , \round_in[2][285] , \round_in[2][284] ,
         \round_in[2][283] , \round_in[2][282] , \round_in[2][281] ,
         \round_in[2][280] , \round_in[2][279] , \round_in[2][278] ,
         \round_in[2][277] , \round_in[2][276] , \round_in[2][275] ,
         \round_in[2][274] , \round_in[2][273] , \round_in[2][272] ,
         \round_in[2][271] , \round_in[2][270] , \round_in[2][269] ,
         \round_in[2][268] , \round_in[2][267] , \round_in[2][266] ,
         \round_in[2][265] , \round_in[2][264] , \round_in[2][263] ,
         \round_in[2][262] , \round_in[2][261] , \round_in[2][260] ,
         \round_in[2][259] , \round_in[2][258] , \round_in[2][257] ,
         \round_in[2][256] , \round_in[2][255] , \round_in[2][254] ,
         \round_in[2][253] , \round_in[2][252] , \round_in[2][251] ,
         \round_in[2][250] , \round_in[2][249] , \round_in[2][248] ,
         \round_in[2][247] , \round_in[2][246] , \round_in[2][245] ,
         \round_in[2][244] , \round_in[2][243] , \round_in[2][242] ,
         \round_in[2][241] , \round_in[2][240] , \round_in[2][239] ,
         \round_in[2][238] , \round_in[2][237] , \round_in[2][236] ,
         \round_in[2][235] , \round_in[2][234] , \round_in[2][233] ,
         \round_in[2][232] , \round_in[2][231] , \round_in[2][230] ,
         \round_in[2][229] , \round_in[2][228] , \round_in[2][227] ,
         \round_in[2][226] , \round_in[2][225] , \round_in[2][224] ,
         \round_in[2][223] , \round_in[2][222] , \round_in[2][221] ,
         \round_in[2][220] , \round_in[2][219] , \round_in[2][218] ,
         \round_in[2][217] , \round_in[2][216] , \round_in[2][215] ,
         \round_in[2][214] , \round_in[2][213] , \round_in[2][212] ,
         \round_in[2][211] , \round_in[2][210] , \round_in[2][209] ,
         \round_in[2][208] , \round_in[2][207] , \round_in[2][206] ,
         \round_in[2][205] , \round_in[2][204] , \round_in[2][203] ,
         \round_in[2][202] , \round_in[2][201] , \round_in[2][200] ,
         \round_in[2][199] , \round_in[2][198] , \round_in[2][197] ,
         \round_in[2][196] , \round_in[2][195] , \round_in[2][194] ,
         \round_in[2][193] , \round_in[2][192] , \round_in[2][191] ,
         \round_in[2][190] , \round_in[2][189] , \round_in[2][188] ,
         \round_in[2][187] , \round_in[2][186] , \round_in[2][185] ,
         \round_in[2][184] , \round_in[2][183] , \round_in[2][182] ,
         \round_in[2][181] , \round_in[2][180] , \round_in[2][179] ,
         \round_in[2][178] , \round_in[2][177] , \round_in[2][176] ,
         \round_in[2][175] , \round_in[2][174] , \round_in[2][173] ,
         \round_in[2][172] , \round_in[2][171] , \round_in[2][170] ,
         \round_in[2][169] , \round_in[2][168] , \round_in[2][167] ,
         \round_in[2][166] , \round_in[2][165] , \round_in[2][164] ,
         \round_in[2][163] , \round_in[2][162] , \round_in[2][161] ,
         \round_in[2][160] , \round_in[2][159] , \round_in[2][158] ,
         \round_in[2][157] , \round_in[2][156] , \round_in[2][155] ,
         \round_in[2][154] , \round_in[2][153] , \round_in[2][152] ,
         \round_in[2][151] , \round_in[2][150] , \round_in[2][149] ,
         \round_in[2][148] , \round_in[2][147] , \round_in[2][146] ,
         \round_in[2][145] , \round_in[2][144] , \round_in[2][143] ,
         \round_in[2][142] , \round_in[2][141] , \round_in[2][140] ,
         \round_in[2][139] , \round_in[2][138] , \round_in[2][137] ,
         \round_in[2][136] , \round_in[2][135] , \round_in[2][134] ,
         \round_in[2][133] , \round_in[2][132] , \round_in[2][131] ,
         \round_in[2][130] , \round_in[2][129] , \round_in[2][128] ,
         \round_in[2][127] , \round_in[2][126] , \round_in[2][125] ,
         \round_in[2][124] , \round_in[2][123] , \round_in[2][122] ,
         \round_in[2][121] , \round_in[2][120] , \round_in[2][119] ,
         \round_in[2][118] , \round_in[2][117] , \round_in[2][116] ,
         \round_in[2][115] , \round_in[2][114] , \round_in[2][113] ,
         \round_in[2][112] , \round_in[2][111] , \round_in[2][110] ,
         \round_in[2][109] , \round_in[2][108] , \round_in[2][107] ,
         \round_in[2][106] , \round_in[2][105] , \round_in[2][104] ,
         \round_in[2][103] , \round_in[2][102] , \round_in[2][101] ,
         \round_in[2][100] , \round_in[2][99] , \round_in[2][98] ,
         \round_in[2][97] , \round_in[2][96] , \round_in[2][95] ,
         \round_in[2][94] , \round_in[2][93] , \round_in[2][92] ,
         \round_in[2][91] , \round_in[2][90] , \round_in[2][89] ,
         \round_in[2][88] , \round_in[2][87] , \round_in[2][86] ,
         \round_in[2][85] , \round_in[2][84] , \round_in[2][83] ,
         \round_in[2][82] , \round_in[2][81] , \round_in[2][80] ,
         \round_in[2][79] , \round_in[2][78] , \round_in[2][77] ,
         \round_in[2][76] , \round_in[2][75] , \round_in[2][74] ,
         \round_in[2][73] , \round_in[2][72] , \round_in[2][71] ,
         \round_in[2][70] , \round_in[2][69] , \round_in[2][68] ,
         \round_in[2][67] , \round_in[2][66] , \round_in[2][65] ,
         \round_in[2][64] , \round_in[2][63] , \round_in[2][62] ,
         \round_in[2][61] , \round_in[2][60] , \round_in[2][59] ,
         \round_in[2][58] , \round_in[2][57] , \round_in[2][56] ,
         \round_in[2][55] , \round_in[2][54] , \round_in[2][53] ,
         \round_in[2][52] , \round_in[2][51] , \round_in[2][50] ,
         \round_in[2][49] , \round_in[2][48] , \round_in[2][47] ,
         \round_in[2][46] , \round_in[2][45] , \round_in[2][44] ,
         \round_in[2][43] , \round_in[2][42] , \round_in[2][41] ,
         \round_in[2][40] , \round_in[2][39] , \round_in[2][38] ,
         \round_in[2][37] , \round_in[2][36] , \round_in[2][35] ,
         \round_in[2][34] , \round_in[2][33] , \round_in[2][32] ,
         \round_in[2][31] , \round_in[2][30] , \round_in[2][29] ,
         \round_in[2][28] , \round_in[2][27] , \round_in[2][26] ,
         \round_in[2][25] , \round_in[2][24] , \round_in[2][23] ,
         \round_in[2][22] , \round_in[2][21] , \round_in[2][20] ,
         \round_in[2][19] , \round_in[2][18] , \round_in[2][17] ,
         \round_in[2][16] , \round_in[2][15] , \round_in[2][14] ,
         \round_in[2][13] , \round_in[2][12] , \round_in[2][11] ,
         \round_in[2][10] , \round_in[2][9] , \round_in[2][8] ,
         \round_in[2][7] , \round_in[2][6] , \round_in[2][5] ,
         \round_in[2][4] , \round_in[2][3] , \round_in[2][2] ,
         \round_in[2][1] , \round_in[2][0] , \round_in[1][1599] ,
         \round_in[1][1598] , \round_in[1][1597] , \round_in[1][1596] ,
         \round_in[1][1595] , \round_in[1][1594] , \round_in[1][1593] ,
         \round_in[1][1592] , \round_in[1][1591] , \round_in[1][1590] ,
         \round_in[1][1589] , \round_in[1][1588] , \round_in[1][1587] ,
         \round_in[1][1586] , \round_in[1][1585] , \round_in[1][1584] ,
         \round_in[1][1583] , \round_in[1][1582] , \round_in[1][1581] ,
         \round_in[1][1580] , \round_in[1][1579] , \round_in[1][1578] ,
         \round_in[1][1577] , \round_in[1][1576] , \round_in[1][1575] ,
         \round_in[1][1574] , \round_in[1][1573] , \round_in[1][1572] ,
         \round_in[1][1571] , \round_in[1][1570] , \round_in[1][1569] ,
         \round_in[1][1568] , \round_in[1][1567] , \round_in[1][1566] ,
         \round_in[1][1565] , \round_in[1][1564] , \round_in[1][1563] ,
         \round_in[1][1562] , \round_in[1][1561] , \round_in[1][1560] ,
         \round_in[1][1559] , \round_in[1][1558] , \round_in[1][1557] ,
         \round_in[1][1556] , \round_in[1][1555] , \round_in[1][1554] ,
         \round_in[1][1553] , \round_in[1][1552] , \round_in[1][1551] ,
         \round_in[1][1550] , \round_in[1][1549] , \round_in[1][1548] ,
         \round_in[1][1547] , \round_in[1][1546] , \round_in[1][1545] ,
         \round_in[1][1544] , \round_in[1][1543] , \round_in[1][1542] ,
         \round_in[1][1541] , \round_in[1][1540] , \round_in[1][1539] ,
         \round_in[1][1538] , \round_in[1][1537] , \round_in[1][1536] ,
         \round_in[1][1535] , \round_in[1][1534] , \round_in[1][1533] ,
         \round_in[1][1532] , \round_in[1][1531] , \round_in[1][1530] ,
         \round_in[1][1529] , \round_in[1][1528] , \round_in[1][1527] ,
         \round_in[1][1526] , \round_in[1][1525] , \round_in[1][1524] ,
         \round_in[1][1523] , \round_in[1][1522] , \round_in[1][1521] ,
         \round_in[1][1520] , \round_in[1][1519] , \round_in[1][1518] ,
         \round_in[1][1517] , \round_in[1][1516] , \round_in[1][1515] ,
         \round_in[1][1514] , \round_in[1][1513] , \round_in[1][1512] ,
         \round_in[1][1511] , \round_in[1][1510] , \round_in[1][1509] ,
         \round_in[1][1508] , \round_in[1][1507] , \round_in[1][1506] ,
         \round_in[1][1505] , \round_in[1][1504] , \round_in[1][1503] ,
         \round_in[1][1502] , \round_in[1][1501] , \round_in[1][1500] ,
         \round_in[1][1499] , \round_in[1][1498] , \round_in[1][1497] ,
         \round_in[1][1496] , \round_in[1][1495] , \round_in[1][1494] ,
         \round_in[1][1493] , \round_in[1][1492] , \round_in[1][1491] ,
         \round_in[1][1490] , \round_in[1][1489] , \round_in[1][1488] ,
         \round_in[1][1487] , \round_in[1][1486] , \round_in[1][1485] ,
         \round_in[1][1484] , \round_in[1][1483] , \round_in[1][1482] ,
         \round_in[1][1481] , \round_in[1][1480] , \round_in[1][1479] ,
         \round_in[1][1478] , \round_in[1][1477] , \round_in[1][1476] ,
         \round_in[1][1475] , \round_in[1][1474] , \round_in[1][1473] ,
         \round_in[1][1472] , \round_in[1][1471] , \round_in[1][1470] ,
         \round_in[1][1469] , \round_in[1][1468] , \round_in[1][1467] ,
         \round_in[1][1466] , \round_in[1][1465] , \round_in[1][1464] ,
         \round_in[1][1463] , \round_in[1][1462] , \round_in[1][1461] ,
         \round_in[1][1460] , \round_in[1][1459] , \round_in[1][1458] ,
         \round_in[1][1457] , \round_in[1][1456] , \round_in[1][1455] ,
         \round_in[1][1454] , \round_in[1][1453] , \round_in[1][1452] ,
         \round_in[1][1451] , \round_in[1][1450] , \round_in[1][1449] ,
         \round_in[1][1448] , \round_in[1][1447] , \round_in[1][1446] ,
         \round_in[1][1445] , \round_in[1][1444] , \round_in[1][1443] ,
         \round_in[1][1442] , \round_in[1][1441] , \round_in[1][1440] ,
         \round_in[1][1439] , \round_in[1][1438] , \round_in[1][1437] ,
         \round_in[1][1436] , \round_in[1][1435] , \round_in[1][1434] ,
         \round_in[1][1433] , \round_in[1][1432] , \round_in[1][1431] ,
         \round_in[1][1430] , \round_in[1][1429] , \round_in[1][1428] ,
         \round_in[1][1427] , \round_in[1][1426] , \round_in[1][1425] ,
         \round_in[1][1424] , \round_in[1][1423] , \round_in[1][1422] ,
         \round_in[1][1421] , \round_in[1][1420] , \round_in[1][1419] ,
         \round_in[1][1418] , \round_in[1][1417] , \round_in[1][1416] ,
         \round_in[1][1415] , \round_in[1][1414] , \round_in[1][1413] ,
         \round_in[1][1412] , \round_in[1][1411] , \round_in[1][1410] ,
         \round_in[1][1409] , \round_in[1][1408] , \round_in[1][1407] ,
         \round_in[1][1406] , \round_in[1][1405] , \round_in[1][1404] ,
         \round_in[1][1403] , \round_in[1][1402] , \round_in[1][1401] ,
         \round_in[1][1400] , \round_in[1][1399] , \round_in[1][1398] ,
         \round_in[1][1397] , \round_in[1][1396] , \round_in[1][1395] ,
         \round_in[1][1394] , \round_in[1][1393] , \round_in[1][1392] ,
         \round_in[1][1391] , \round_in[1][1390] , \round_in[1][1389] ,
         \round_in[1][1388] , \round_in[1][1387] , \round_in[1][1386] ,
         \round_in[1][1385] , \round_in[1][1384] , \round_in[1][1383] ,
         \round_in[1][1382] , \round_in[1][1381] , \round_in[1][1380] ,
         \round_in[1][1379] , \round_in[1][1378] , \round_in[1][1377] ,
         \round_in[1][1376] , \round_in[1][1375] , \round_in[1][1374] ,
         \round_in[1][1373] , \round_in[1][1372] , \round_in[1][1371] ,
         \round_in[1][1370] , \round_in[1][1369] , \round_in[1][1368] ,
         \round_in[1][1367] , \round_in[1][1366] , \round_in[1][1365] ,
         \round_in[1][1364] , \round_in[1][1363] , \round_in[1][1362] ,
         \round_in[1][1361] , \round_in[1][1360] , \round_in[1][1359] ,
         \round_in[1][1358] , \round_in[1][1357] , \round_in[1][1356] ,
         \round_in[1][1355] , \round_in[1][1354] , \round_in[1][1353] ,
         \round_in[1][1352] , \round_in[1][1351] , \round_in[1][1350] ,
         \round_in[1][1349] , \round_in[1][1348] , \round_in[1][1347] ,
         \round_in[1][1346] , \round_in[1][1345] , \round_in[1][1344] ,
         \round_in[1][1343] , \round_in[1][1342] , \round_in[1][1341] ,
         \round_in[1][1340] , \round_in[1][1339] , \round_in[1][1338] ,
         \round_in[1][1337] , \round_in[1][1336] , \round_in[1][1335] ,
         \round_in[1][1334] , \round_in[1][1333] , \round_in[1][1332] ,
         \round_in[1][1331] , \round_in[1][1330] , \round_in[1][1329] ,
         \round_in[1][1328] , \round_in[1][1327] , \round_in[1][1326] ,
         \round_in[1][1325] , \round_in[1][1324] , \round_in[1][1323] ,
         \round_in[1][1322] , \round_in[1][1321] , \round_in[1][1320] ,
         \round_in[1][1319] , \round_in[1][1318] , \round_in[1][1317] ,
         \round_in[1][1316] , \round_in[1][1315] , \round_in[1][1314] ,
         \round_in[1][1313] , \round_in[1][1312] , \round_in[1][1311] ,
         \round_in[1][1310] , \round_in[1][1309] , \round_in[1][1308] ,
         \round_in[1][1307] , \round_in[1][1306] , \round_in[1][1305] ,
         \round_in[1][1304] , \round_in[1][1303] , \round_in[1][1302] ,
         \round_in[1][1301] , \round_in[1][1300] , \round_in[1][1299] ,
         \round_in[1][1298] , \round_in[1][1297] , \round_in[1][1296] ,
         \round_in[1][1295] , \round_in[1][1294] , \round_in[1][1293] ,
         \round_in[1][1292] , \round_in[1][1291] , \round_in[1][1290] ,
         \round_in[1][1289] , \round_in[1][1288] , \round_in[1][1287] ,
         \round_in[1][1286] , \round_in[1][1285] , \round_in[1][1284] ,
         \round_in[1][1283] , \round_in[1][1282] , \round_in[1][1281] ,
         \round_in[1][1280] , \round_in[1][1279] , \round_in[1][1278] ,
         \round_in[1][1277] , \round_in[1][1276] , \round_in[1][1275] ,
         \round_in[1][1274] , \round_in[1][1273] , \round_in[1][1272] ,
         \round_in[1][1271] , \round_in[1][1270] , \round_in[1][1269] ,
         \round_in[1][1268] , \round_in[1][1267] , \round_in[1][1266] ,
         \round_in[1][1265] , \round_in[1][1264] , \round_in[1][1263] ,
         \round_in[1][1262] , \round_in[1][1261] , \round_in[1][1260] ,
         \round_in[1][1259] , \round_in[1][1258] , \round_in[1][1257] ,
         \round_in[1][1256] , \round_in[1][1255] , \round_in[1][1254] ,
         \round_in[1][1253] , \round_in[1][1252] , \round_in[1][1251] ,
         \round_in[1][1250] , \round_in[1][1249] , \round_in[1][1248] ,
         \round_in[1][1247] , \round_in[1][1246] , \round_in[1][1245] ,
         \round_in[1][1244] , \round_in[1][1243] , \round_in[1][1242] ,
         \round_in[1][1241] , \round_in[1][1240] , \round_in[1][1239] ,
         \round_in[1][1238] , \round_in[1][1237] , \round_in[1][1236] ,
         \round_in[1][1235] , \round_in[1][1234] , \round_in[1][1233] ,
         \round_in[1][1232] , \round_in[1][1231] , \round_in[1][1230] ,
         \round_in[1][1229] , \round_in[1][1228] , \round_in[1][1227] ,
         \round_in[1][1226] , \round_in[1][1225] , \round_in[1][1224] ,
         \round_in[1][1223] , \round_in[1][1222] , \round_in[1][1221] ,
         \round_in[1][1220] , \round_in[1][1219] , \round_in[1][1218] ,
         \round_in[1][1217] , \round_in[1][1216] , \round_in[1][1215] ,
         \round_in[1][1214] , \round_in[1][1213] , \round_in[1][1212] ,
         \round_in[1][1211] , \round_in[1][1210] , \round_in[1][1209] ,
         \round_in[1][1208] , \round_in[1][1207] , \round_in[1][1206] ,
         \round_in[1][1205] , \round_in[1][1204] , \round_in[1][1203] ,
         \round_in[1][1202] , \round_in[1][1201] , \round_in[1][1200] ,
         \round_in[1][1199] , \round_in[1][1198] , \round_in[1][1197] ,
         \round_in[1][1196] , \round_in[1][1195] , \round_in[1][1194] ,
         \round_in[1][1193] , \round_in[1][1192] , \round_in[1][1191] ,
         \round_in[1][1190] , \round_in[1][1189] , \round_in[1][1188] ,
         \round_in[1][1187] , \round_in[1][1186] , \round_in[1][1185] ,
         \round_in[1][1184] , \round_in[1][1183] , \round_in[1][1182] ,
         \round_in[1][1181] , \round_in[1][1180] , \round_in[1][1179] ,
         \round_in[1][1178] , \round_in[1][1177] , \round_in[1][1176] ,
         \round_in[1][1175] , \round_in[1][1174] , \round_in[1][1173] ,
         \round_in[1][1172] , \round_in[1][1171] , \round_in[1][1170] ,
         \round_in[1][1169] , \round_in[1][1168] , \round_in[1][1167] ,
         \round_in[1][1166] , \round_in[1][1165] , \round_in[1][1164] ,
         \round_in[1][1163] , \round_in[1][1162] , \round_in[1][1161] ,
         \round_in[1][1160] , \round_in[1][1159] , \round_in[1][1158] ,
         \round_in[1][1157] , \round_in[1][1156] , \round_in[1][1155] ,
         \round_in[1][1154] , \round_in[1][1153] , \round_in[1][1152] ,
         \round_in[1][1151] , \round_in[1][1150] , \round_in[1][1149] ,
         \round_in[1][1148] , \round_in[1][1147] , \round_in[1][1146] ,
         \round_in[1][1145] , \round_in[1][1144] , \round_in[1][1143] ,
         \round_in[1][1142] , \round_in[1][1141] , \round_in[1][1140] ,
         \round_in[1][1139] , \round_in[1][1138] , \round_in[1][1137] ,
         \round_in[1][1136] , \round_in[1][1135] , \round_in[1][1134] ,
         \round_in[1][1133] , \round_in[1][1132] , \round_in[1][1131] ,
         \round_in[1][1130] , \round_in[1][1129] , \round_in[1][1128] ,
         \round_in[1][1127] , \round_in[1][1126] , \round_in[1][1125] ,
         \round_in[1][1124] , \round_in[1][1123] , \round_in[1][1122] ,
         \round_in[1][1121] , \round_in[1][1120] , \round_in[1][1119] ,
         \round_in[1][1118] , \round_in[1][1117] , \round_in[1][1116] ,
         \round_in[1][1115] , \round_in[1][1114] , \round_in[1][1113] ,
         \round_in[1][1112] , \round_in[1][1111] , \round_in[1][1110] ,
         \round_in[1][1109] , \round_in[1][1108] , \round_in[1][1107] ,
         \round_in[1][1106] , \round_in[1][1105] , \round_in[1][1104] ,
         \round_in[1][1103] , \round_in[1][1102] , \round_in[1][1101] ,
         \round_in[1][1100] , \round_in[1][1099] , \round_in[1][1098] ,
         \round_in[1][1097] , \round_in[1][1096] , \round_in[1][1095] ,
         \round_in[1][1094] , \round_in[1][1093] , \round_in[1][1092] ,
         \round_in[1][1091] , \round_in[1][1090] , \round_in[1][1089] ,
         \round_in[1][1088] , \round_in[1][1087] , \round_in[1][1086] ,
         \round_in[1][1085] , \round_in[1][1084] , \round_in[1][1083] ,
         \round_in[1][1082] , \round_in[1][1081] , \round_in[1][1080] ,
         \round_in[1][1079] , \round_in[1][1078] , \round_in[1][1077] ,
         \round_in[1][1076] , \round_in[1][1075] , \round_in[1][1074] ,
         \round_in[1][1073] , \round_in[1][1072] , \round_in[1][1071] ,
         \round_in[1][1070] , \round_in[1][1069] , \round_in[1][1068] ,
         \round_in[1][1067] , \round_in[1][1066] , \round_in[1][1065] ,
         \round_in[1][1064] , \round_in[1][1063] , \round_in[1][1062] ,
         \round_in[1][1061] , \round_in[1][1060] , \round_in[1][1059] ,
         \round_in[1][1058] , \round_in[1][1057] , \round_in[1][1056] ,
         \round_in[1][1055] , \round_in[1][1054] , \round_in[1][1053] ,
         \round_in[1][1052] , \round_in[1][1051] , \round_in[1][1050] ,
         \round_in[1][1049] , \round_in[1][1048] , \round_in[1][1047] ,
         \round_in[1][1046] , \round_in[1][1045] , \round_in[1][1044] ,
         \round_in[1][1043] , \round_in[1][1042] , \round_in[1][1041] ,
         \round_in[1][1040] , \round_in[1][1039] , \round_in[1][1038] ,
         \round_in[1][1037] , \round_in[1][1036] , \round_in[1][1035] ,
         \round_in[1][1034] , \round_in[1][1033] , \round_in[1][1032] ,
         \round_in[1][1031] , \round_in[1][1030] , \round_in[1][1029] ,
         \round_in[1][1028] , \round_in[1][1027] , \round_in[1][1026] ,
         \round_in[1][1025] , \round_in[1][1024] , \round_in[1][1023] ,
         \round_in[1][1022] , \round_in[1][1021] , \round_in[1][1020] ,
         \round_in[1][1019] , \round_in[1][1018] , \round_in[1][1017] ,
         \round_in[1][1016] , \round_in[1][1015] , \round_in[1][1014] ,
         \round_in[1][1013] , \round_in[1][1012] , \round_in[1][1011] ,
         \round_in[1][1010] , \round_in[1][1009] , \round_in[1][1008] ,
         \round_in[1][1007] , \round_in[1][1006] , \round_in[1][1005] ,
         \round_in[1][1004] , \round_in[1][1003] , \round_in[1][1002] ,
         \round_in[1][1001] , \round_in[1][1000] , \round_in[1][999] ,
         \round_in[1][998] , \round_in[1][997] , \round_in[1][996] ,
         \round_in[1][995] , \round_in[1][994] , \round_in[1][993] ,
         \round_in[1][992] , \round_in[1][991] , \round_in[1][990] ,
         \round_in[1][989] , \round_in[1][988] , \round_in[1][987] ,
         \round_in[1][986] , \round_in[1][985] , \round_in[1][984] ,
         \round_in[1][983] , \round_in[1][982] , \round_in[1][981] ,
         \round_in[1][980] , \round_in[1][979] , \round_in[1][978] ,
         \round_in[1][977] , \round_in[1][976] , \round_in[1][975] ,
         \round_in[1][974] , \round_in[1][973] , \round_in[1][972] ,
         \round_in[1][971] , \round_in[1][970] , \round_in[1][969] ,
         \round_in[1][968] , \round_in[1][967] , \round_in[1][966] ,
         \round_in[1][965] , \round_in[1][964] , \round_in[1][963] ,
         \round_in[1][962] , \round_in[1][961] , \round_in[1][960] ,
         \round_in[1][959] , \round_in[1][958] , \round_in[1][957] ,
         \round_in[1][956] , \round_in[1][955] , \round_in[1][954] ,
         \round_in[1][953] , \round_in[1][952] , \round_in[1][951] ,
         \round_in[1][950] , \round_in[1][949] , \round_in[1][948] ,
         \round_in[1][947] , \round_in[1][946] , \round_in[1][945] ,
         \round_in[1][944] , \round_in[1][943] , \round_in[1][942] ,
         \round_in[1][941] , \round_in[1][940] , \round_in[1][939] ,
         \round_in[1][938] , \round_in[1][937] , \round_in[1][936] ,
         \round_in[1][935] , \round_in[1][934] , \round_in[1][933] ,
         \round_in[1][932] , \round_in[1][931] , \round_in[1][930] ,
         \round_in[1][929] , \round_in[1][928] , \round_in[1][927] ,
         \round_in[1][926] , \round_in[1][925] , \round_in[1][924] ,
         \round_in[1][923] , \round_in[1][922] , \round_in[1][921] ,
         \round_in[1][920] , \round_in[1][919] , \round_in[1][918] ,
         \round_in[1][917] , \round_in[1][916] , \round_in[1][915] ,
         \round_in[1][914] , \round_in[1][913] , \round_in[1][912] ,
         \round_in[1][911] , \round_in[1][910] , \round_in[1][909] ,
         \round_in[1][908] , \round_in[1][907] , \round_in[1][906] ,
         \round_in[1][905] , \round_in[1][904] , \round_in[1][903] ,
         \round_in[1][902] , \round_in[1][901] , \round_in[1][900] ,
         \round_in[1][899] , \round_in[1][898] , \round_in[1][897] ,
         \round_in[1][896] , \round_in[1][895] , \round_in[1][894] ,
         \round_in[1][893] , \round_in[1][892] , \round_in[1][891] ,
         \round_in[1][890] , \round_in[1][889] , \round_in[1][888] ,
         \round_in[1][887] , \round_in[1][886] , \round_in[1][885] ,
         \round_in[1][884] , \round_in[1][883] , \round_in[1][882] ,
         \round_in[1][881] , \round_in[1][880] , \round_in[1][879] ,
         \round_in[1][878] , \round_in[1][877] , \round_in[1][876] ,
         \round_in[1][875] , \round_in[1][874] , \round_in[1][873] ,
         \round_in[1][872] , \round_in[1][871] , \round_in[1][870] ,
         \round_in[1][869] , \round_in[1][868] , \round_in[1][867] ,
         \round_in[1][866] , \round_in[1][865] , \round_in[1][864] ,
         \round_in[1][863] , \round_in[1][862] , \round_in[1][861] ,
         \round_in[1][860] , \round_in[1][859] , \round_in[1][858] ,
         \round_in[1][857] , \round_in[1][856] , \round_in[1][855] ,
         \round_in[1][854] , \round_in[1][853] , \round_in[1][852] ,
         \round_in[1][851] , \round_in[1][850] , \round_in[1][849] ,
         \round_in[1][848] , \round_in[1][847] , \round_in[1][846] ,
         \round_in[1][845] , \round_in[1][844] , \round_in[1][843] ,
         \round_in[1][842] , \round_in[1][841] , \round_in[1][840] ,
         \round_in[1][839] , \round_in[1][838] , \round_in[1][837] ,
         \round_in[1][836] , \round_in[1][835] , \round_in[1][834] ,
         \round_in[1][833] , \round_in[1][832] , \round_in[1][831] ,
         \round_in[1][830] , \round_in[1][829] , \round_in[1][828] ,
         \round_in[1][827] , \round_in[1][826] , \round_in[1][825] ,
         \round_in[1][824] , \round_in[1][823] , \round_in[1][822] ,
         \round_in[1][821] , \round_in[1][820] , \round_in[1][819] ,
         \round_in[1][818] , \round_in[1][817] , \round_in[1][816] ,
         \round_in[1][815] , \round_in[1][814] , \round_in[1][813] ,
         \round_in[1][812] , \round_in[1][811] , \round_in[1][810] ,
         \round_in[1][809] , \round_in[1][808] , \round_in[1][807] ,
         \round_in[1][806] , \round_in[1][805] , \round_in[1][804] ,
         \round_in[1][803] , \round_in[1][802] , \round_in[1][801] ,
         \round_in[1][800] , \round_in[1][799] , \round_in[1][798] ,
         \round_in[1][797] , \round_in[1][796] , \round_in[1][795] ,
         \round_in[1][794] , \round_in[1][793] , \round_in[1][792] ,
         \round_in[1][791] , \round_in[1][790] , \round_in[1][789] ,
         \round_in[1][788] , \round_in[1][787] , \round_in[1][786] ,
         \round_in[1][785] , \round_in[1][784] , \round_in[1][783] ,
         \round_in[1][782] , \round_in[1][781] , \round_in[1][780] ,
         \round_in[1][779] , \round_in[1][778] , \round_in[1][777] ,
         \round_in[1][776] , \round_in[1][775] , \round_in[1][774] ,
         \round_in[1][773] , \round_in[1][772] , \round_in[1][771] ,
         \round_in[1][770] , \round_in[1][769] , \round_in[1][768] ,
         \round_in[1][767] , \round_in[1][766] , \round_in[1][765] ,
         \round_in[1][764] , \round_in[1][763] , \round_in[1][762] ,
         \round_in[1][761] , \round_in[1][760] , \round_in[1][759] ,
         \round_in[1][758] , \round_in[1][757] , \round_in[1][756] ,
         \round_in[1][755] , \round_in[1][754] , \round_in[1][753] ,
         \round_in[1][752] , \round_in[1][751] , \round_in[1][750] ,
         \round_in[1][749] , \round_in[1][748] , \round_in[1][747] ,
         \round_in[1][746] , \round_in[1][745] , \round_in[1][744] ,
         \round_in[1][743] , \round_in[1][742] , \round_in[1][741] ,
         \round_in[1][740] , \round_in[1][739] , \round_in[1][738] ,
         \round_in[1][737] , \round_in[1][736] , \round_in[1][735] ,
         \round_in[1][734] , \round_in[1][733] , \round_in[1][732] ,
         \round_in[1][731] , \round_in[1][730] , \round_in[1][729] ,
         \round_in[1][728] , \round_in[1][727] , \round_in[1][726] ,
         \round_in[1][725] , \round_in[1][724] , \round_in[1][723] ,
         \round_in[1][722] , \round_in[1][721] , \round_in[1][720] ,
         \round_in[1][719] , \round_in[1][718] , \round_in[1][717] ,
         \round_in[1][716] , \round_in[1][715] , \round_in[1][714] ,
         \round_in[1][713] , \round_in[1][712] , \round_in[1][711] ,
         \round_in[1][710] , \round_in[1][709] , \round_in[1][708] ,
         \round_in[1][707] , \round_in[1][706] , \round_in[1][705] ,
         \round_in[1][704] , \round_in[1][703] , \round_in[1][702] ,
         \round_in[1][701] , \round_in[1][700] , \round_in[1][699] ,
         \round_in[1][698] , \round_in[1][697] , \round_in[1][696] ,
         \round_in[1][695] , \round_in[1][694] , \round_in[1][693] ,
         \round_in[1][692] , \round_in[1][691] , \round_in[1][690] ,
         \round_in[1][689] , \round_in[1][688] , \round_in[1][687] ,
         \round_in[1][686] , \round_in[1][685] , \round_in[1][684] ,
         \round_in[1][683] , \round_in[1][682] , \round_in[1][681] ,
         \round_in[1][680] , \round_in[1][679] , \round_in[1][678] ,
         \round_in[1][677] , \round_in[1][676] , \round_in[1][675] ,
         \round_in[1][674] , \round_in[1][673] , \round_in[1][672] ,
         \round_in[1][671] , \round_in[1][670] , \round_in[1][669] ,
         \round_in[1][668] , \round_in[1][667] , \round_in[1][666] ,
         \round_in[1][665] , \round_in[1][664] , \round_in[1][663] ,
         \round_in[1][662] , \round_in[1][661] , \round_in[1][660] ,
         \round_in[1][659] , \round_in[1][658] , \round_in[1][657] ,
         \round_in[1][656] , \round_in[1][655] , \round_in[1][654] ,
         \round_in[1][653] , \round_in[1][652] , \round_in[1][651] ,
         \round_in[1][650] , \round_in[1][649] , \round_in[1][648] ,
         \round_in[1][647] , \round_in[1][646] , \round_in[1][645] ,
         \round_in[1][644] , \round_in[1][643] , \round_in[1][642] ,
         \round_in[1][641] , \round_in[1][640] , \round_in[1][639] ,
         \round_in[1][638] , \round_in[1][637] , \round_in[1][636] ,
         \round_in[1][635] , \round_in[1][634] , \round_in[1][633] ,
         \round_in[1][632] , \round_in[1][631] , \round_in[1][630] ,
         \round_in[1][629] , \round_in[1][628] , \round_in[1][627] ,
         \round_in[1][626] , \round_in[1][625] , \round_in[1][624] ,
         \round_in[1][623] , \round_in[1][622] , \round_in[1][621] ,
         \round_in[1][620] , \round_in[1][619] , \round_in[1][618] ,
         \round_in[1][617] , \round_in[1][616] , \round_in[1][615] ,
         \round_in[1][614] , \round_in[1][613] , \round_in[1][612] ,
         \round_in[1][611] , \round_in[1][610] , \round_in[1][609] ,
         \round_in[1][608] , \round_in[1][607] , \round_in[1][606] ,
         \round_in[1][605] , \round_in[1][604] , \round_in[1][603] ,
         \round_in[1][602] , \round_in[1][601] , \round_in[1][600] ,
         \round_in[1][599] , \round_in[1][598] , \round_in[1][597] ,
         \round_in[1][596] , \round_in[1][595] , \round_in[1][594] ,
         \round_in[1][593] , \round_in[1][592] , \round_in[1][591] ,
         \round_in[1][590] , \round_in[1][589] , \round_in[1][588] ,
         \round_in[1][587] , \round_in[1][586] , \round_in[1][585] ,
         \round_in[1][584] , \round_in[1][583] , \round_in[1][582] ,
         \round_in[1][581] , \round_in[1][580] , \round_in[1][579] ,
         \round_in[1][578] , \round_in[1][577] , \round_in[1][576] ,
         \round_in[1][575] , \round_in[1][574] , \round_in[1][573] ,
         \round_in[1][572] , \round_in[1][571] , \round_in[1][570] ,
         \round_in[1][569] , \round_in[1][568] , \round_in[1][567] ,
         \round_in[1][566] , \round_in[1][565] , \round_in[1][564] ,
         \round_in[1][563] , \round_in[1][562] , \round_in[1][561] ,
         \round_in[1][560] , \round_in[1][559] , \round_in[1][558] ,
         \round_in[1][557] , \round_in[1][556] , \round_in[1][555] ,
         \round_in[1][554] , \round_in[1][553] , \round_in[1][552] ,
         \round_in[1][551] , \round_in[1][550] , \round_in[1][549] ,
         \round_in[1][548] , \round_in[1][547] , \round_in[1][546] ,
         \round_in[1][545] , \round_in[1][544] , \round_in[1][543] ,
         \round_in[1][542] , \round_in[1][541] , \round_in[1][540] ,
         \round_in[1][539] , \round_in[1][538] , \round_in[1][537] ,
         \round_in[1][536] , \round_in[1][535] , \round_in[1][534] ,
         \round_in[1][533] , \round_in[1][532] , \round_in[1][531] ,
         \round_in[1][530] , \round_in[1][529] , \round_in[1][528] ,
         \round_in[1][527] , \round_in[1][526] , \round_in[1][525] ,
         \round_in[1][524] , \round_in[1][523] , \round_in[1][522] ,
         \round_in[1][521] , \round_in[1][520] , \round_in[1][519] ,
         \round_in[1][518] , \round_in[1][517] , \round_in[1][516] ,
         \round_in[1][515] , \round_in[1][514] , \round_in[1][513] ,
         \round_in[1][512] , \round_in[1][511] , \round_in[1][510] ,
         \round_in[1][509] , \round_in[1][508] , \round_in[1][507] ,
         \round_in[1][506] , \round_in[1][505] , \round_in[1][504] ,
         \round_in[1][503] , \round_in[1][502] , \round_in[1][501] ,
         \round_in[1][500] , \round_in[1][499] , \round_in[1][498] ,
         \round_in[1][497] , \round_in[1][496] , \round_in[1][495] ,
         \round_in[1][494] , \round_in[1][493] , \round_in[1][492] ,
         \round_in[1][491] , \round_in[1][490] , \round_in[1][489] ,
         \round_in[1][488] , \round_in[1][487] , \round_in[1][486] ,
         \round_in[1][485] , \round_in[1][484] , \round_in[1][483] ,
         \round_in[1][482] , \round_in[1][481] , \round_in[1][480] ,
         \round_in[1][479] , \round_in[1][478] , \round_in[1][477] ,
         \round_in[1][476] , \round_in[1][475] , \round_in[1][474] ,
         \round_in[1][473] , \round_in[1][472] , \round_in[1][471] ,
         \round_in[1][470] , \round_in[1][469] , \round_in[1][468] ,
         \round_in[1][467] , \round_in[1][466] , \round_in[1][465] ,
         \round_in[1][464] , \round_in[1][463] , \round_in[1][462] ,
         \round_in[1][461] , \round_in[1][460] , \round_in[1][459] ,
         \round_in[1][458] , \round_in[1][457] , \round_in[1][456] ,
         \round_in[1][455] , \round_in[1][454] , \round_in[1][453] ,
         \round_in[1][452] , \round_in[1][451] , \round_in[1][450] ,
         \round_in[1][449] , \round_in[1][448] , \round_in[1][447] ,
         \round_in[1][446] , \round_in[1][445] , \round_in[1][444] ,
         \round_in[1][443] , \round_in[1][442] , \round_in[1][441] ,
         \round_in[1][440] , \round_in[1][439] , \round_in[1][438] ,
         \round_in[1][437] , \round_in[1][436] , \round_in[1][435] ,
         \round_in[1][434] , \round_in[1][433] , \round_in[1][432] ,
         \round_in[1][431] , \round_in[1][430] , \round_in[1][429] ,
         \round_in[1][428] , \round_in[1][427] , \round_in[1][426] ,
         \round_in[1][425] , \round_in[1][424] , \round_in[1][423] ,
         \round_in[1][422] , \round_in[1][421] , \round_in[1][420] ,
         \round_in[1][419] , \round_in[1][418] , \round_in[1][417] ,
         \round_in[1][416] , \round_in[1][415] , \round_in[1][414] ,
         \round_in[1][413] , \round_in[1][412] , \round_in[1][411] ,
         \round_in[1][410] , \round_in[1][409] , \round_in[1][408] ,
         \round_in[1][407] , \round_in[1][406] , \round_in[1][405] ,
         \round_in[1][404] , \round_in[1][403] , \round_in[1][402] ,
         \round_in[1][401] , \round_in[1][400] , \round_in[1][399] ,
         \round_in[1][398] , \round_in[1][397] , \round_in[1][396] ,
         \round_in[1][395] , \round_in[1][394] , \round_in[1][393] ,
         \round_in[1][392] , \round_in[1][391] , \round_in[1][390] ,
         \round_in[1][389] , \round_in[1][388] , \round_in[1][387] ,
         \round_in[1][386] , \round_in[1][385] , \round_in[1][384] ,
         \round_in[1][383] , \round_in[1][382] , \round_in[1][381] ,
         \round_in[1][380] , \round_in[1][379] , \round_in[1][378] ,
         \round_in[1][377] , \round_in[1][376] , \round_in[1][375] ,
         \round_in[1][374] , \round_in[1][373] , \round_in[1][372] ,
         \round_in[1][371] , \round_in[1][370] , \round_in[1][369] ,
         \round_in[1][368] , \round_in[1][367] , \round_in[1][366] ,
         \round_in[1][365] , \round_in[1][364] , \round_in[1][363] ,
         \round_in[1][362] , \round_in[1][361] , \round_in[1][360] ,
         \round_in[1][359] , \round_in[1][358] , \round_in[1][357] ,
         \round_in[1][356] , \round_in[1][355] , \round_in[1][354] ,
         \round_in[1][353] , \round_in[1][352] , \round_in[1][351] ,
         \round_in[1][350] , \round_in[1][349] , \round_in[1][348] ,
         \round_in[1][347] , \round_in[1][346] , \round_in[1][345] ,
         \round_in[1][344] , \round_in[1][343] , \round_in[1][342] ,
         \round_in[1][341] , \round_in[1][340] , \round_in[1][339] ,
         \round_in[1][338] , \round_in[1][337] , \round_in[1][336] ,
         \round_in[1][335] , \round_in[1][334] , \round_in[1][333] ,
         \round_in[1][332] , \round_in[1][331] , \round_in[1][330] ,
         \round_in[1][329] , \round_in[1][328] , \round_in[1][327] ,
         \round_in[1][326] , \round_in[1][325] , \round_in[1][324] ,
         \round_in[1][323] , \round_in[1][322] , \round_in[1][321] ,
         \round_in[1][320] , \round_in[1][319] , \round_in[1][318] ,
         \round_in[1][317] , \round_in[1][316] , \round_in[1][315] ,
         \round_in[1][314] , \round_in[1][313] , \round_in[1][312] ,
         \round_in[1][311] , \round_in[1][310] , \round_in[1][309] ,
         \round_in[1][308] , \round_in[1][307] , \round_in[1][306] ,
         \round_in[1][305] , \round_in[1][304] , \round_in[1][303] ,
         \round_in[1][302] , \round_in[1][301] , \round_in[1][300] ,
         \round_in[1][299] , \round_in[1][298] , \round_in[1][297] ,
         \round_in[1][296] , \round_in[1][295] , \round_in[1][294] ,
         \round_in[1][293] , \round_in[1][292] , \round_in[1][291] ,
         \round_in[1][290] , \round_in[1][289] , \round_in[1][288] ,
         \round_in[1][287] , \round_in[1][286] , \round_in[1][285] ,
         \round_in[1][284] , \round_in[1][283] , \round_in[1][282] ,
         \round_in[1][281] , \round_in[1][280] , \round_in[1][279] ,
         \round_in[1][278] , \round_in[1][277] , \round_in[1][276] ,
         \round_in[1][275] , \round_in[1][274] , \round_in[1][273] ,
         \round_in[1][272] , \round_in[1][271] , \round_in[1][270] ,
         \round_in[1][269] , \round_in[1][268] , \round_in[1][267] ,
         \round_in[1][266] , \round_in[1][265] , \round_in[1][264] ,
         \round_in[1][263] , \round_in[1][262] , \round_in[1][261] ,
         \round_in[1][260] , \round_in[1][259] , \round_in[1][258] ,
         \round_in[1][257] , \round_in[1][256] , \round_in[1][255] ,
         \round_in[1][254] , \round_in[1][253] , \round_in[1][252] ,
         \round_in[1][251] , \round_in[1][250] , \round_in[1][249] ,
         \round_in[1][248] , \round_in[1][247] , \round_in[1][246] ,
         \round_in[1][245] , \round_in[1][244] , \round_in[1][243] ,
         \round_in[1][242] , \round_in[1][241] , \round_in[1][240] ,
         \round_in[1][239] , \round_in[1][238] , \round_in[1][237] ,
         \round_in[1][236] , \round_in[1][235] , \round_in[1][234] ,
         \round_in[1][233] , \round_in[1][232] , \round_in[1][231] ,
         \round_in[1][230] , \round_in[1][229] , \round_in[1][228] ,
         \round_in[1][227] , \round_in[1][226] , \round_in[1][225] ,
         \round_in[1][224] , \round_in[1][223] , \round_in[1][222] ,
         \round_in[1][221] , \round_in[1][220] , \round_in[1][219] ,
         \round_in[1][218] , \round_in[1][217] , \round_in[1][216] ,
         \round_in[1][215] , \round_in[1][214] , \round_in[1][213] ,
         \round_in[1][212] , \round_in[1][211] , \round_in[1][210] ,
         \round_in[1][209] , \round_in[1][208] , \round_in[1][207] ,
         \round_in[1][206] , \round_in[1][205] , \round_in[1][204] ,
         \round_in[1][203] , \round_in[1][202] , \round_in[1][201] ,
         \round_in[1][200] , \round_in[1][199] , \round_in[1][198] ,
         \round_in[1][197] , \round_in[1][196] , \round_in[1][195] ,
         \round_in[1][194] , \round_in[1][193] , \round_in[1][192] ,
         \round_in[1][191] , \round_in[1][190] , \round_in[1][189] ,
         \round_in[1][188] , \round_in[1][187] , \round_in[1][186] ,
         \round_in[1][185] , \round_in[1][184] , \round_in[1][183] ,
         \round_in[1][182] , \round_in[1][181] , \round_in[1][180] ,
         \round_in[1][179] , \round_in[1][178] , \round_in[1][177] ,
         \round_in[1][176] , \round_in[1][175] , \round_in[1][174] ,
         \round_in[1][173] , \round_in[1][172] , \round_in[1][171] ,
         \round_in[1][170] , \round_in[1][169] , \round_in[1][168] ,
         \round_in[1][167] , \round_in[1][166] , \round_in[1][165] ,
         \round_in[1][164] , \round_in[1][163] , \round_in[1][162] ,
         \round_in[1][161] , \round_in[1][160] , \round_in[1][159] ,
         \round_in[1][158] , \round_in[1][157] , \round_in[1][156] ,
         \round_in[1][155] , \round_in[1][154] , \round_in[1][153] ,
         \round_in[1][152] , \round_in[1][151] , \round_in[1][150] ,
         \round_in[1][149] , \round_in[1][148] , \round_in[1][147] ,
         \round_in[1][146] , \round_in[1][145] , \round_in[1][144] ,
         \round_in[1][143] , \round_in[1][142] , \round_in[1][141] ,
         \round_in[1][140] , \round_in[1][139] , \round_in[1][138] ,
         \round_in[1][137] , \round_in[1][136] , \round_in[1][135] ,
         \round_in[1][134] , \round_in[1][133] , \round_in[1][132] ,
         \round_in[1][131] , \round_in[1][130] , \round_in[1][129] ,
         \round_in[1][128] , \round_in[1][127] , \round_in[1][126] ,
         \round_in[1][125] , \round_in[1][124] , \round_in[1][123] ,
         \round_in[1][122] , \round_in[1][121] , \round_in[1][120] ,
         \round_in[1][119] , \round_in[1][118] , \round_in[1][117] ,
         \round_in[1][116] , \round_in[1][115] , \round_in[1][114] ,
         \round_in[1][113] , \round_in[1][112] , \round_in[1][111] ,
         \round_in[1][110] , \round_in[1][109] , \round_in[1][108] ,
         \round_in[1][107] , \round_in[1][106] , \round_in[1][105] ,
         \round_in[1][104] , \round_in[1][103] , \round_in[1][102] ,
         \round_in[1][101] , \round_in[1][100] , \round_in[1][99] ,
         \round_in[1][98] , \round_in[1][97] , \round_in[1][96] ,
         \round_in[1][95] , \round_in[1][94] , \round_in[1][93] ,
         \round_in[1][92] , \round_in[1][91] , \round_in[1][90] ,
         \round_in[1][89] , \round_in[1][88] , \round_in[1][87] ,
         \round_in[1][86] , \round_in[1][85] , \round_in[1][84] ,
         \round_in[1][83] , \round_in[1][82] , \round_in[1][81] ,
         \round_in[1][80] , \round_in[1][79] , \round_in[1][78] ,
         \round_in[1][77] , \round_in[1][76] , \round_in[1][75] ,
         \round_in[1][74] , \round_in[1][73] , \round_in[1][72] ,
         \round_in[1][71] , \round_in[1][70] , \round_in[1][69] ,
         \round_in[1][68] , \round_in[1][67] , \round_in[1][66] ,
         \round_in[1][65] , \round_in[1][64] , \round_in[1][63] ,
         \round_in[1][62] , \round_in[1][61] , \round_in[1][60] ,
         \round_in[1][59] , \round_in[1][58] , \round_in[1][57] ,
         \round_in[1][56] , \round_in[1][55] , \round_in[1][54] ,
         \round_in[1][53] , \round_in[1][52] , \round_in[1][51] ,
         \round_in[1][50] , \round_in[1][49] , \round_in[1][48] ,
         \round_in[1][47] , \round_in[1][46] , \round_in[1][45] ,
         \round_in[1][44] , \round_in[1][43] , \round_in[1][42] ,
         \round_in[1][41] , \round_in[1][40] , \round_in[1][39] ,
         \round_in[1][38] , \round_in[1][37] , \round_in[1][36] ,
         \round_in[1][35] , \round_in[1][34] , \round_in[1][33] ,
         \round_in[1][32] , \round_in[1][31] , \round_in[1][30] ,
         \round_in[1][29] , \round_in[1][28] , \round_in[1][27] ,
         \round_in[1][26] , \round_in[1][25] , \round_in[1][24] ,
         \round_in[1][23] , \round_in[1][22] , \round_in[1][21] ,
         \round_in[1][20] , \round_in[1][19] , \round_in[1][18] ,
         \round_in[1][17] , \round_in[1][16] , \round_in[1][15] ,
         \round_in[1][14] , \round_in[1][13] , \round_in[1][12] ,
         \round_in[1][11] , \round_in[1][10] , \round_in[1][9] ,
         \round_in[1][8] , \round_in[1][7] , \round_in[1][6] ,
         \round_in[1][5] , \round_in[1][4] , \round_in[1][3] ,
         \round_in[1][2] , \round_in[1][1] , \round_in[1][0] ,
         \round_in[0][1599] , \round_in[0][1598] , \round_in[0][1597] ,
         \round_in[0][1596] , \round_in[0][1595] , \round_in[0][1594] ,
         \round_in[0][1593] , \round_in[0][1592] , \round_in[0][1591] ,
         \round_in[0][1590] , \round_in[0][1589] , \round_in[0][1588] ,
         \round_in[0][1587] , \round_in[0][1586] , \round_in[0][1585] ,
         \round_in[0][1584] , \round_in[0][1583] , \round_in[0][1582] ,
         \round_in[0][1581] , \round_in[0][1580] , \round_in[0][1579] ,
         \round_in[0][1578] , \round_in[0][1577] , \round_in[0][1576] ,
         \round_in[0][1575] , \round_in[0][1574] , \round_in[0][1573] ,
         \round_in[0][1572] , \round_in[0][1571] , \round_in[0][1570] ,
         \round_in[0][1569] , \round_in[0][1568] , \round_in[0][1567] ,
         \round_in[0][1566] , \round_in[0][1565] , \round_in[0][1564] ,
         \round_in[0][1563] , \round_in[0][1562] , \round_in[0][1561] ,
         \round_in[0][1560] , \round_in[0][1559] , \round_in[0][1558] ,
         \round_in[0][1557] , \round_in[0][1556] , \round_in[0][1555] ,
         \round_in[0][1554] , \round_in[0][1553] , \round_in[0][1552] ,
         \round_in[0][1551] , \round_in[0][1550] , \round_in[0][1549] ,
         \round_in[0][1548] , \round_in[0][1547] , \round_in[0][1546] ,
         \round_in[0][1545] , \round_in[0][1544] , \round_in[0][1543] ,
         \round_in[0][1542] , \round_in[0][1541] , \round_in[0][1540] ,
         \round_in[0][1539] , \round_in[0][1538] , \round_in[0][1537] ,
         \round_in[0][1536] , \round_in[0][1535] , \round_in[0][1534] ,
         \round_in[0][1533] , \round_in[0][1532] , \round_in[0][1531] ,
         \round_in[0][1530] , \round_in[0][1529] , \round_in[0][1528] ,
         \round_in[0][1527] , \round_in[0][1526] , \round_in[0][1525] ,
         \round_in[0][1524] , \round_in[0][1523] , \round_in[0][1522] ,
         \round_in[0][1521] , \round_in[0][1520] , \round_in[0][1519] ,
         \round_in[0][1518] , \round_in[0][1517] , \round_in[0][1516] ,
         \round_in[0][1515] , \round_in[0][1514] , \round_in[0][1513] ,
         \round_in[0][1512] , \round_in[0][1511] , \round_in[0][1510] ,
         \round_in[0][1509] , \round_in[0][1508] , \round_in[0][1507] ,
         \round_in[0][1506] , \round_in[0][1505] , \round_in[0][1504] ,
         \round_in[0][1503] , \round_in[0][1502] , \round_in[0][1501] ,
         \round_in[0][1500] , \round_in[0][1499] , \round_in[0][1498] ,
         \round_in[0][1497] , \round_in[0][1496] , \round_in[0][1495] ,
         \round_in[0][1494] , \round_in[0][1493] , \round_in[0][1492] ,
         \round_in[0][1491] , \round_in[0][1490] , \round_in[0][1489] ,
         \round_in[0][1488] , \round_in[0][1487] , \round_in[0][1486] ,
         \round_in[0][1485] , \round_in[0][1484] , \round_in[0][1483] ,
         \round_in[0][1482] , \round_in[0][1481] , \round_in[0][1480] ,
         \round_in[0][1479] , \round_in[0][1478] , \round_in[0][1477] ,
         \round_in[0][1476] , \round_in[0][1475] , \round_in[0][1474] ,
         \round_in[0][1473] , \round_in[0][1472] , \round_in[0][1471] ,
         \round_in[0][1470] , \round_in[0][1469] , \round_in[0][1468] ,
         \round_in[0][1467] , \round_in[0][1466] , \round_in[0][1465] ,
         \round_in[0][1464] , \round_in[0][1463] , \round_in[0][1462] ,
         \round_in[0][1461] , \round_in[0][1460] , \round_in[0][1459] ,
         \round_in[0][1458] , \round_in[0][1457] , \round_in[0][1456] ,
         \round_in[0][1455] , \round_in[0][1454] , \round_in[0][1453] ,
         \round_in[0][1452] , \round_in[0][1451] , \round_in[0][1450] ,
         \round_in[0][1449] , \round_in[0][1448] , \round_in[0][1447] ,
         \round_in[0][1446] , \round_in[0][1445] , \round_in[0][1444] ,
         \round_in[0][1443] , \round_in[0][1442] , \round_in[0][1441] ,
         \round_in[0][1440] , \round_in[0][1439] , \round_in[0][1438] ,
         \round_in[0][1437] , \round_in[0][1436] , \round_in[0][1435] ,
         \round_in[0][1434] , \round_in[0][1433] , \round_in[0][1432] ,
         \round_in[0][1431] , \round_in[0][1430] , \round_in[0][1429] ,
         \round_in[0][1428] , \round_in[0][1427] , \round_in[0][1426] ,
         \round_in[0][1425] , \round_in[0][1424] , \round_in[0][1423] ,
         \round_in[0][1422] , \round_in[0][1421] , \round_in[0][1420] ,
         \round_in[0][1419] , \round_in[0][1418] , \round_in[0][1417] ,
         \round_in[0][1416] , \round_in[0][1415] , \round_in[0][1414] ,
         \round_in[0][1413] , \round_in[0][1412] , \round_in[0][1411] ,
         \round_in[0][1410] , \round_in[0][1409] , \round_in[0][1408] ,
         \round_in[0][1407] , \round_in[0][1406] , \round_in[0][1405] ,
         \round_in[0][1404] , \round_in[0][1403] , \round_in[0][1402] ,
         \round_in[0][1401] , \round_in[0][1400] , \round_in[0][1399] ,
         \round_in[0][1398] , \round_in[0][1397] , \round_in[0][1396] ,
         \round_in[0][1395] , \round_in[0][1394] , \round_in[0][1393] ,
         \round_in[0][1392] , \round_in[0][1391] , \round_in[0][1390] ,
         \round_in[0][1389] , \round_in[0][1388] , \round_in[0][1387] ,
         \round_in[0][1386] , \round_in[0][1385] , \round_in[0][1384] ,
         \round_in[0][1383] , \round_in[0][1382] , \round_in[0][1381] ,
         \round_in[0][1380] , \round_in[0][1379] , \round_in[0][1378] ,
         \round_in[0][1377] , \round_in[0][1376] , \round_in[0][1375] ,
         \round_in[0][1374] , \round_in[0][1373] , \round_in[0][1372] ,
         \round_in[0][1371] , \round_in[0][1370] , \round_in[0][1369] ,
         \round_in[0][1368] , \round_in[0][1367] , \round_in[0][1366] ,
         \round_in[0][1365] , \round_in[0][1364] , \round_in[0][1363] ,
         \round_in[0][1362] , \round_in[0][1361] , \round_in[0][1360] ,
         \round_in[0][1359] , \round_in[0][1358] , \round_in[0][1357] ,
         \round_in[0][1356] , \round_in[0][1355] , \round_in[0][1354] ,
         \round_in[0][1353] , \round_in[0][1352] , \round_in[0][1351] ,
         \round_in[0][1350] , \round_in[0][1349] , \round_in[0][1348] ,
         \round_in[0][1347] , \round_in[0][1346] , \round_in[0][1345] ,
         \round_in[0][1344] , \round_in[0][1343] , \round_in[0][1342] ,
         \round_in[0][1341] , \round_in[0][1340] , \round_in[0][1339] ,
         \round_in[0][1338] , \round_in[0][1337] , \round_in[0][1336] ,
         \round_in[0][1335] , \round_in[0][1334] , \round_in[0][1333] ,
         \round_in[0][1332] , \round_in[0][1331] , \round_in[0][1330] ,
         \round_in[0][1329] , \round_in[0][1328] , \round_in[0][1327] ,
         \round_in[0][1326] , \round_in[0][1325] , \round_in[0][1324] ,
         \round_in[0][1323] , \round_in[0][1322] , \round_in[0][1321] ,
         \round_in[0][1320] , \round_in[0][1319] , \round_in[0][1318] ,
         \round_in[0][1317] , \round_in[0][1316] , \round_in[0][1315] ,
         \round_in[0][1314] , \round_in[0][1313] , \round_in[0][1312] ,
         \round_in[0][1311] , \round_in[0][1310] , \round_in[0][1309] ,
         \round_in[0][1308] , \round_in[0][1307] , \round_in[0][1306] ,
         \round_in[0][1305] , \round_in[0][1304] , \round_in[0][1303] ,
         \round_in[0][1302] , \round_in[0][1301] , \round_in[0][1300] ,
         \round_in[0][1299] , \round_in[0][1298] , \round_in[0][1297] ,
         \round_in[0][1296] , \round_in[0][1295] , \round_in[0][1294] ,
         \round_in[0][1293] , \round_in[0][1292] , \round_in[0][1291] ,
         \round_in[0][1290] , \round_in[0][1289] , \round_in[0][1288] ,
         \round_in[0][1287] , \round_in[0][1286] , \round_in[0][1285] ,
         \round_in[0][1284] , \round_in[0][1283] , \round_in[0][1282] ,
         \round_in[0][1281] , \round_in[0][1280] , \round_in[0][1279] ,
         \round_in[0][1278] , \round_in[0][1277] , \round_in[0][1276] ,
         \round_in[0][1275] , \round_in[0][1274] , \round_in[0][1273] ,
         \round_in[0][1272] , \round_in[0][1271] , \round_in[0][1270] ,
         \round_in[0][1269] , \round_in[0][1268] , \round_in[0][1267] ,
         \round_in[0][1266] , \round_in[0][1265] , \round_in[0][1264] ,
         \round_in[0][1263] , \round_in[0][1262] , \round_in[0][1261] ,
         \round_in[0][1260] , \round_in[0][1259] , \round_in[0][1258] ,
         \round_in[0][1257] , \round_in[0][1256] , \round_in[0][1255] ,
         \round_in[0][1254] , \round_in[0][1253] , \round_in[0][1252] ,
         \round_in[0][1251] , \round_in[0][1250] , \round_in[0][1249] ,
         \round_in[0][1248] , \round_in[0][1247] , \round_in[0][1246] ,
         \round_in[0][1245] , \round_in[0][1244] , \round_in[0][1243] ,
         \round_in[0][1242] , \round_in[0][1241] , \round_in[0][1240] ,
         \round_in[0][1239] , \round_in[0][1238] , \round_in[0][1237] ,
         \round_in[0][1236] , \round_in[0][1235] , \round_in[0][1234] ,
         \round_in[0][1233] , \round_in[0][1232] , \round_in[0][1231] ,
         \round_in[0][1230] , \round_in[0][1229] , \round_in[0][1228] ,
         \round_in[0][1227] , \round_in[0][1226] , \round_in[0][1225] ,
         \round_in[0][1224] , \round_in[0][1223] , \round_in[0][1222] ,
         \round_in[0][1221] , \round_in[0][1220] , \round_in[0][1219] ,
         \round_in[0][1218] , \round_in[0][1217] , \round_in[0][1216] ,
         \round_in[0][1215] , \round_in[0][1214] , \round_in[0][1213] ,
         \round_in[0][1212] , \round_in[0][1211] , \round_in[0][1210] ,
         \round_in[0][1209] , \round_in[0][1208] , \round_in[0][1207] ,
         \round_in[0][1206] , \round_in[0][1205] , \round_in[0][1204] ,
         \round_in[0][1203] , \round_in[0][1202] , \round_in[0][1201] ,
         \round_in[0][1200] , \round_in[0][1199] , \round_in[0][1198] ,
         \round_in[0][1197] , \round_in[0][1196] , \round_in[0][1195] ,
         \round_in[0][1194] , \round_in[0][1193] , \round_in[0][1192] ,
         \round_in[0][1191] , \round_in[0][1190] , \round_in[0][1189] ,
         \round_in[0][1188] , \round_in[0][1187] , \round_in[0][1186] ,
         \round_in[0][1185] , \round_in[0][1184] , \round_in[0][1183] ,
         \round_in[0][1182] , \round_in[0][1181] , \round_in[0][1180] ,
         \round_in[0][1179] , \round_in[0][1178] , \round_in[0][1177] ,
         \round_in[0][1176] , \round_in[0][1175] , \round_in[0][1174] ,
         \round_in[0][1173] , \round_in[0][1172] , \round_in[0][1171] ,
         \round_in[0][1170] , \round_in[0][1169] , \round_in[0][1168] ,
         \round_in[0][1167] , \round_in[0][1166] , \round_in[0][1165] ,
         \round_in[0][1164] , \round_in[0][1163] , \round_in[0][1162] ,
         \round_in[0][1161] , \round_in[0][1160] , \round_in[0][1159] ,
         \round_in[0][1158] , \round_in[0][1157] , \round_in[0][1156] ,
         \round_in[0][1155] , \round_in[0][1154] , \round_in[0][1153] ,
         \round_in[0][1152] , \round_in[0][1151] , \round_in[0][1150] ,
         \round_in[0][1149] , \round_in[0][1148] , \round_in[0][1147] ,
         \round_in[0][1146] , \round_in[0][1145] , \round_in[0][1144] ,
         \round_in[0][1143] , \round_in[0][1142] , \round_in[0][1141] ,
         \round_in[0][1140] , \round_in[0][1139] , \round_in[0][1138] ,
         \round_in[0][1137] , \round_in[0][1136] , \round_in[0][1135] ,
         \round_in[0][1134] , \round_in[0][1133] , \round_in[0][1132] ,
         \round_in[0][1131] , \round_in[0][1130] , \round_in[0][1129] ,
         \round_in[0][1128] , \round_in[0][1127] , \round_in[0][1126] ,
         \round_in[0][1125] , \round_in[0][1124] , \round_in[0][1123] ,
         \round_in[0][1122] , \round_in[0][1121] , \round_in[0][1120] ,
         \round_in[0][1119] , \round_in[0][1118] , \round_in[0][1117] ,
         \round_in[0][1116] , \round_in[0][1115] , \round_in[0][1114] ,
         \round_in[0][1113] , \round_in[0][1112] , \round_in[0][1111] ,
         \round_in[0][1110] , \round_in[0][1109] , \round_in[0][1108] ,
         \round_in[0][1107] , \round_in[0][1106] , \round_in[0][1105] ,
         \round_in[0][1104] , \round_in[0][1103] , \round_in[0][1102] ,
         \round_in[0][1101] , \round_in[0][1100] , \round_in[0][1099] ,
         \round_in[0][1098] , \round_in[0][1097] , \round_in[0][1096] ,
         \round_in[0][1095] , \round_in[0][1094] , \round_in[0][1093] ,
         \round_in[0][1092] , \round_in[0][1091] , \round_in[0][1090] ,
         \round_in[0][1089] , \round_in[0][1088] , \round_in[0][1087] ,
         \round_in[0][1086] , \round_in[0][1085] , \round_in[0][1084] ,
         \round_in[0][1083] , \round_in[0][1082] , \round_in[0][1081] ,
         \round_in[0][1080] , \round_in[0][1079] , \round_in[0][1078] ,
         \round_in[0][1077] , \round_in[0][1076] , \round_in[0][1075] ,
         \round_in[0][1074] , \round_in[0][1073] , \round_in[0][1072] ,
         \round_in[0][1071] , \round_in[0][1070] , \round_in[0][1069] ,
         \round_in[0][1068] , \round_in[0][1067] , \round_in[0][1066] ,
         \round_in[0][1065] , \round_in[0][1064] , \round_in[0][1063] ,
         \round_in[0][1062] , \round_in[0][1061] , \round_in[0][1060] ,
         \round_in[0][1059] , \round_in[0][1058] , \round_in[0][1057] ,
         \round_in[0][1056] , \round_in[0][1055] , \round_in[0][1054] ,
         \round_in[0][1053] , \round_in[0][1052] , \round_in[0][1051] ,
         \round_in[0][1050] , \round_in[0][1049] , \round_in[0][1048] ,
         \round_in[0][1047] , \round_in[0][1046] , \round_in[0][1045] ,
         \round_in[0][1044] , \round_in[0][1043] , \round_in[0][1042] ,
         \round_in[0][1041] , \round_in[0][1040] , \round_in[0][1039] ,
         \round_in[0][1038] , \round_in[0][1037] , \round_in[0][1036] ,
         \round_in[0][1035] , \round_in[0][1034] , \round_in[0][1033] ,
         \round_in[0][1032] , \round_in[0][1031] , \round_in[0][1030] ,
         \round_in[0][1029] , \round_in[0][1028] , \round_in[0][1027] ,
         \round_in[0][1026] , \round_in[0][1025] , \round_in[0][1024] ,
         \round_in[0][1023] , \round_in[0][1022] , \round_in[0][1021] ,
         \round_in[0][1020] , \round_in[0][1019] , \round_in[0][1018] ,
         \round_in[0][1017] , \round_in[0][1016] , \round_in[0][1015] ,
         \round_in[0][1014] , \round_in[0][1013] , \round_in[0][1012] ,
         \round_in[0][1011] , \round_in[0][1010] , \round_in[0][1009] ,
         \round_in[0][1008] , \round_in[0][1007] , \round_in[0][1006] ,
         \round_in[0][1005] , \round_in[0][1004] , \round_in[0][1003] ,
         \round_in[0][1002] , \round_in[0][1001] , \round_in[0][1000] ,
         \round_in[0][999] , \round_in[0][998] , \round_in[0][997] ,
         \round_in[0][996] , \round_in[0][995] , \round_in[0][994] ,
         \round_in[0][993] , \round_in[0][992] , \round_in[0][991] ,
         \round_in[0][990] , \round_in[0][989] , \round_in[0][988] ,
         \round_in[0][987] , \round_in[0][986] , \round_in[0][985] ,
         \round_in[0][984] , \round_in[0][983] , \round_in[0][982] ,
         \round_in[0][981] , \round_in[0][980] , \round_in[0][979] ,
         \round_in[0][978] , \round_in[0][977] , \round_in[0][976] ,
         \round_in[0][975] , \round_in[0][974] , \round_in[0][973] ,
         \round_in[0][972] , \round_in[0][971] , \round_in[0][970] ,
         \round_in[0][969] , \round_in[0][968] , \round_in[0][967] ,
         \round_in[0][966] , \round_in[0][965] , \round_in[0][964] ,
         \round_in[0][963] , \round_in[0][962] , \round_in[0][961] ,
         \round_in[0][960] , \round_in[0][959] , \round_in[0][958] ,
         \round_in[0][957] , \round_in[0][956] , \round_in[0][955] ,
         \round_in[0][954] , \round_in[0][953] , \round_in[0][952] ,
         \round_in[0][951] , \round_in[0][950] , \round_in[0][949] ,
         \round_in[0][948] , \round_in[0][947] , \round_in[0][946] ,
         \round_in[0][945] , \round_in[0][944] , \round_in[0][943] ,
         \round_in[0][942] , \round_in[0][941] , \round_in[0][940] ,
         \round_in[0][939] , \round_in[0][938] , \round_in[0][937] ,
         \round_in[0][936] , \round_in[0][935] , \round_in[0][934] ,
         \round_in[0][933] , \round_in[0][932] , \round_in[0][931] ,
         \round_in[0][930] , \round_in[0][929] , \round_in[0][928] ,
         \round_in[0][927] , \round_in[0][926] , \round_in[0][925] ,
         \round_in[0][924] , \round_in[0][923] , \round_in[0][922] ,
         \round_in[0][921] , \round_in[0][920] , \round_in[0][919] ,
         \round_in[0][918] , \round_in[0][917] , \round_in[0][916] ,
         \round_in[0][915] , \round_in[0][914] , \round_in[0][913] ,
         \round_in[0][912] , \round_in[0][911] , \round_in[0][910] ,
         \round_in[0][909] , \round_in[0][908] , \round_in[0][907] ,
         \round_in[0][906] , \round_in[0][905] , \round_in[0][904] ,
         \round_in[0][903] , \round_in[0][902] , \round_in[0][901] ,
         \round_in[0][900] , \round_in[0][899] , \round_in[0][898] ,
         \round_in[0][897] , \round_in[0][896] , \round_in[0][895] ,
         \round_in[0][894] , \round_in[0][893] , \round_in[0][892] ,
         \round_in[0][891] , \round_in[0][890] , \round_in[0][889] ,
         \round_in[0][888] , \round_in[0][887] , \round_in[0][886] ,
         \round_in[0][885] , \round_in[0][884] , \round_in[0][883] ,
         \round_in[0][882] , \round_in[0][881] , \round_in[0][880] ,
         \round_in[0][879] , \round_in[0][878] , \round_in[0][877] ,
         \round_in[0][876] , \round_in[0][875] , \round_in[0][874] ,
         \round_in[0][873] , \round_in[0][872] , \round_in[0][871] ,
         \round_in[0][870] , \round_in[0][869] , \round_in[0][868] ,
         \round_in[0][867] , \round_in[0][866] , \round_in[0][865] ,
         \round_in[0][864] , \round_in[0][863] , \round_in[0][862] ,
         \round_in[0][861] , \round_in[0][860] , \round_in[0][859] ,
         \round_in[0][858] , \round_in[0][857] , \round_in[0][856] ,
         \round_in[0][855] , \round_in[0][854] , \round_in[0][853] ,
         \round_in[0][852] , \round_in[0][851] , \round_in[0][850] ,
         \round_in[0][849] , \round_in[0][848] , \round_in[0][847] ,
         \round_in[0][846] , \round_in[0][845] , \round_in[0][844] ,
         \round_in[0][843] , \round_in[0][842] , \round_in[0][841] ,
         \round_in[0][840] , \round_in[0][839] , \round_in[0][838] ,
         \round_in[0][837] , \round_in[0][836] , \round_in[0][835] ,
         \round_in[0][834] , \round_in[0][833] , \round_in[0][832] ,
         \round_in[0][831] , \round_in[0][830] , \round_in[0][829] ,
         \round_in[0][828] , \round_in[0][827] , \round_in[0][826] ,
         \round_in[0][825] , \round_in[0][824] , \round_in[0][823] ,
         \round_in[0][822] , \round_in[0][821] , \round_in[0][820] ,
         \round_in[0][819] , \round_in[0][818] , \round_in[0][817] ,
         \round_in[0][816] , \round_in[0][815] , \round_in[0][814] ,
         \round_in[0][813] , \round_in[0][812] , \round_in[0][811] ,
         \round_in[0][810] , \round_in[0][809] , \round_in[0][808] ,
         \round_in[0][807] , \round_in[0][806] , \round_in[0][805] ,
         \round_in[0][804] , \round_in[0][803] , \round_in[0][802] ,
         \round_in[0][801] , \round_in[0][800] , \round_in[0][799] ,
         \round_in[0][798] , \round_in[0][797] , \round_in[0][796] ,
         \round_in[0][795] , \round_in[0][794] , \round_in[0][793] ,
         \round_in[0][792] , \round_in[0][791] , \round_in[0][790] ,
         \round_in[0][789] , \round_in[0][788] , \round_in[0][787] ,
         \round_in[0][786] , \round_in[0][785] , \round_in[0][784] ,
         \round_in[0][783] , \round_in[0][782] , \round_in[0][781] ,
         \round_in[0][780] , \round_in[0][779] , \round_in[0][778] ,
         \round_in[0][777] , \round_in[0][776] , \round_in[0][775] ,
         \round_in[0][774] , \round_in[0][773] , \round_in[0][772] ,
         \round_in[0][771] , \round_in[0][770] , \round_in[0][769] ,
         \round_in[0][768] , \round_in[0][767] , \round_in[0][766] ,
         \round_in[0][765] , \round_in[0][764] , \round_in[0][763] ,
         \round_in[0][762] , \round_in[0][761] , \round_in[0][760] ,
         \round_in[0][759] , \round_in[0][758] , \round_in[0][757] ,
         \round_in[0][756] , \round_in[0][755] , \round_in[0][754] ,
         \round_in[0][753] , \round_in[0][752] , \round_in[0][751] ,
         \round_in[0][750] , \round_in[0][749] , \round_in[0][748] ,
         \round_in[0][747] , \round_in[0][746] , \round_in[0][745] ,
         \round_in[0][744] , \round_in[0][743] , \round_in[0][742] ,
         \round_in[0][741] , \round_in[0][740] , \round_in[0][739] ,
         \round_in[0][738] , \round_in[0][737] , \round_in[0][736] ,
         \round_in[0][735] , \round_in[0][734] , \round_in[0][733] ,
         \round_in[0][732] , \round_in[0][731] , \round_in[0][730] ,
         \round_in[0][729] , \round_in[0][728] , \round_in[0][727] ,
         \round_in[0][726] , \round_in[0][725] , \round_in[0][724] ,
         \round_in[0][723] , \round_in[0][722] , \round_in[0][721] ,
         \round_in[0][720] , \round_in[0][719] , \round_in[0][718] ,
         \round_in[0][717] , \round_in[0][716] , \round_in[0][715] ,
         \round_in[0][714] , \round_in[0][713] , \round_in[0][712] ,
         \round_in[0][711] , \round_in[0][710] , \round_in[0][709] ,
         \round_in[0][708] , \round_in[0][707] , \round_in[0][706] ,
         \round_in[0][705] , \round_in[0][704] , \round_in[0][703] ,
         \round_in[0][702] , \round_in[0][701] , \round_in[0][700] ,
         \round_in[0][699] , \round_in[0][698] , \round_in[0][697] ,
         \round_in[0][696] , \round_in[0][695] , \round_in[0][694] ,
         \round_in[0][693] , \round_in[0][692] , \round_in[0][691] ,
         \round_in[0][690] , \round_in[0][689] , \round_in[0][688] ,
         \round_in[0][687] , \round_in[0][686] , \round_in[0][685] ,
         \round_in[0][684] , \round_in[0][683] , \round_in[0][682] ,
         \round_in[0][681] , \round_in[0][680] , \round_in[0][679] ,
         \round_in[0][678] , \round_in[0][677] , \round_in[0][676] ,
         \round_in[0][675] , \round_in[0][674] , \round_in[0][673] ,
         \round_in[0][672] , \round_in[0][671] , \round_in[0][670] ,
         \round_in[0][669] , \round_in[0][668] , \round_in[0][667] ,
         \round_in[0][666] , \round_in[0][665] , \round_in[0][664] ,
         \round_in[0][663] , \round_in[0][662] , \round_in[0][661] ,
         \round_in[0][660] , \round_in[0][659] , \round_in[0][658] ,
         \round_in[0][657] , \round_in[0][656] , \round_in[0][655] ,
         \round_in[0][654] , \round_in[0][653] , \round_in[0][652] ,
         \round_in[0][651] , \round_in[0][650] , \round_in[0][649] ,
         \round_in[0][648] , \round_in[0][647] , \round_in[0][646] ,
         \round_in[0][645] , \round_in[0][644] , \round_in[0][643] ,
         \round_in[0][642] , \round_in[0][641] , \round_in[0][640] ,
         \round_in[0][639] , \round_in[0][638] , \round_in[0][637] ,
         \round_in[0][636] , \round_in[0][635] , \round_in[0][634] ,
         \round_in[0][633] , \round_in[0][632] , \round_in[0][631] ,
         \round_in[0][630] , \round_in[0][629] , \round_in[0][628] ,
         \round_in[0][627] , \round_in[0][626] , \round_in[0][625] ,
         \round_in[0][624] , \round_in[0][623] , \round_in[0][622] ,
         \round_in[0][621] , \round_in[0][620] , \round_in[0][619] ,
         \round_in[0][618] , \round_in[0][617] , \round_in[0][616] ,
         \round_in[0][615] , \round_in[0][614] , \round_in[0][613] ,
         \round_in[0][612] , \round_in[0][611] , \round_in[0][610] ,
         \round_in[0][609] , \round_in[0][608] , \round_in[0][607] ,
         \round_in[0][606] , \round_in[0][605] , \round_in[0][604] ,
         \round_in[0][603] , \round_in[0][602] , \round_in[0][601] ,
         \round_in[0][600] , \round_in[0][599] , \round_in[0][598] ,
         \round_in[0][597] , \round_in[0][596] , \round_in[0][595] ,
         \round_in[0][594] , \round_in[0][593] , \round_in[0][592] ,
         \round_in[0][591] , \round_in[0][590] , \round_in[0][589] ,
         \round_in[0][588] , \round_in[0][587] , \round_in[0][586] ,
         \round_in[0][585] , \round_in[0][584] , \round_in[0][583] ,
         \round_in[0][582] , \round_in[0][581] , \round_in[0][580] ,
         \round_in[0][579] , \round_in[0][578] , \round_in[0][577] ,
         \round_in[0][576] , \round_in[0][575] , \round_in[0][574] ,
         \round_in[0][573] , \round_in[0][572] , \round_in[0][571] ,
         \round_in[0][570] , \round_in[0][569] , \round_in[0][568] ,
         \round_in[0][567] , \round_in[0][566] , \round_in[0][565] ,
         \round_in[0][564] , \round_in[0][563] , \round_in[0][562] ,
         \round_in[0][561] , \round_in[0][560] , \round_in[0][559] ,
         \round_in[0][558] , \round_in[0][557] , \round_in[0][556] ,
         \round_in[0][555] , \round_in[0][554] , \round_in[0][553] ,
         \round_in[0][552] , \round_in[0][551] , \round_in[0][550] ,
         \round_in[0][549] , \round_in[0][548] , \round_in[0][547] ,
         \round_in[0][546] , \round_in[0][545] , \round_in[0][544] ,
         \round_in[0][543] , \round_in[0][542] , \round_in[0][541] ,
         \round_in[0][540] , \round_in[0][539] , \round_in[0][538] ,
         \round_in[0][537] , \round_in[0][536] , \round_in[0][535] ,
         \round_in[0][534] , \round_in[0][533] , \round_in[0][532] ,
         \round_in[0][531] , \round_in[0][530] , \round_in[0][529] ,
         \round_in[0][528] , \round_in[0][527] , \round_in[0][526] ,
         \round_in[0][525] , \round_in[0][524] , \round_in[0][523] ,
         \round_in[0][522] , \round_in[0][521] , \round_in[0][520] ,
         \round_in[0][519] , \round_in[0][518] , \round_in[0][517] ,
         \round_in[0][516] , \round_in[0][515] , \round_in[0][514] ,
         \round_in[0][513] , \round_in[0][512] , \round_in[0][511] ,
         \round_in[0][510] , \round_in[0][509] , \round_in[0][508] ,
         \round_in[0][507] , \round_in[0][506] , \round_in[0][505] ,
         \round_in[0][504] , \round_in[0][503] , \round_in[0][502] ,
         \round_in[0][501] , \round_in[0][500] , \round_in[0][499] ,
         \round_in[0][498] , \round_in[0][497] , \round_in[0][496] ,
         \round_in[0][495] , \round_in[0][494] , \round_in[0][493] ,
         \round_in[0][492] , \round_in[0][491] , \round_in[0][490] ,
         \round_in[0][489] , \round_in[0][488] , \round_in[0][487] ,
         \round_in[0][486] , \round_in[0][485] , \round_in[0][484] ,
         \round_in[0][483] , \round_in[0][482] , \round_in[0][481] ,
         \round_in[0][480] , \round_in[0][479] , \round_in[0][478] ,
         \round_in[0][477] , \round_in[0][476] , \round_in[0][475] ,
         \round_in[0][474] , \round_in[0][473] , \round_in[0][472] ,
         \round_in[0][471] , \round_in[0][470] , \round_in[0][469] ,
         \round_in[0][468] , \round_in[0][467] , \round_in[0][466] ,
         \round_in[0][465] , \round_in[0][464] , \round_in[0][463] ,
         \round_in[0][462] , \round_in[0][461] , \round_in[0][460] ,
         \round_in[0][459] , \round_in[0][458] , \round_in[0][457] ,
         \round_in[0][456] , \round_in[0][455] , \round_in[0][454] ,
         \round_in[0][453] , \round_in[0][452] , \round_in[0][451] ,
         \round_in[0][450] , \round_in[0][449] , \round_in[0][448] ,
         \round_in[0][447] , \round_in[0][446] , \round_in[0][445] ,
         \round_in[0][444] , \round_in[0][443] , \round_in[0][442] ,
         \round_in[0][441] , \round_in[0][440] , \round_in[0][439] ,
         \round_in[0][438] , \round_in[0][437] , \round_in[0][436] ,
         \round_in[0][435] , \round_in[0][434] , \round_in[0][433] ,
         \round_in[0][432] , \round_in[0][431] , \round_in[0][430] ,
         \round_in[0][429] , \round_in[0][428] , \round_in[0][427] ,
         \round_in[0][426] , \round_in[0][425] , \round_in[0][424] ,
         \round_in[0][423] , \round_in[0][422] , \round_in[0][421] ,
         \round_in[0][420] , \round_in[0][419] , \round_in[0][418] ,
         \round_in[0][417] , \round_in[0][416] , \round_in[0][415] ,
         \round_in[0][414] , \round_in[0][413] , \round_in[0][412] ,
         \round_in[0][411] , \round_in[0][410] , \round_in[0][409] ,
         \round_in[0][408] , \round_in[0][407] , \round_in[0][406] ,
         \round_in[0][405] , \round_in[0][404] , \round_in[0][403] ,
         \round_in[0][402] , \round_in[0][401] , \round_in[0][400] ,
         \round_in[0][399] , \round_in[0][398] , \round_in[0][397] ,
         \round_in[0][396] , \round_in[0][395] , \round_in[0][394] ,
         \round_in[0][393] , \round_in[0][392] , \round_in[0][391] ,
         \round_in[0][390] , \round_in[0][389] , \round_in[0][388] ,
         \round_in[0][387] , \round_in[0][386] , \round_in[0][385] ,
         \round_in[0][384] , \round_in[0][383] , \round_in[0][382] ,
         \round_in[0][381] , \round_in[0][380] , \round_in[0][379] ,
         \round_in[0][378] , \round_in[0][377] , \round_in[0][376] ,
         \round_in[0][375] , \round_in[0][374] , \round_in[0][373] ,
         \round_in[0][372] , \round_in[0][371] , \round_in[0][370] ,
         \round_in[0][369] , \round_in[0][368] , \round_in[0][367] ,
         \round_in[0][366] , \round_in[0][365] , \round_in[0][364] ,
         \round_in[0][363] , \round_in[0][362] , \round_in[0][361] ,
         \round_in[0][360] , \round_in[0][359] , \round_in[0][358] ,
         \round_in[0][357] , \round_in[0][356] , \round_in[0][355] ,
         \round_in[0][354] , \round_in[0][353] , \round_in[0][352] ,
         \round_in[0][351] , \round_in[0][350] , \round_in[0][349] ,
         \round_in[0][348] , \round_in[0][347] , \round_in[0][346] ,
         \round_in[0][345] , \round_in[0][344] , \round_in[0][343] ,
         \round_in[0][342] , \round_in[0][341] , \round_in[0][340] ,
         \round_in[0][339] , \round_in[0][338] , \round_in[0][337] ,
         \round_in[0][336] , \round_in[0][335] , \round_in[0][334] ,
         \round_in[0][333] , \round_in[0][332] , \round_in[0][331] ,
         \round_in[0][330] , \round_in[0][329] , \round_in[0][328] ,
         \round_in[0][327] , \round_in[0][326] , \round_in[0][325] ,
         \round_in[0][324] , \round_in[0][323] , \round_in[0][322] ,
         \round_in[0][321] , \round_in[0][320] , \round_in[0][319] ,
         \round_in[0][318] , \round_in[0][317] , \round_in[0][316] ,
         \round_in[0][315] , \round_in[0][314] , \round_in[0][313] ,
         \round_in[0][312] , \round_in[0][311] , \round_in[0][310] ,
         \round_in[0][309] , \round_in[0][308] , \round_in[0][307] ,
         \round_in[0][306] , \round_in[0][305] , \round_in[0][304] ,
         \round_in[0][303] , \round_in[0][302] , \round_in[0][301] ,
         \round_in[0][300] , \round_in[0][299] , \round_in[0][298] ,
         \round_in[0][297] , \round_in[0][296] , \round_in[0][295] ,
         \round_in[0][294] , \round_in[0][293] , \round_in[0][292] ,
         \round_in[0][291] , \round_in[0][290] , \round_in[0][289] ,
         \round_in[0][288] , \round_in[0][287] , \round_in[0][286] ,
         \round_in[0][285] , \round_in[0][284] , \round_in[0][283] ,
         \round_in[0][282] , \round_in[0][281] , \round_in[0][280] ,
         \round_in[0][279] , \round_in[0][278] , \round_in[0][277] ,
         \round_in[0][276] , \round_in[0][275] , \round_in[0][274] ,
         \round_in[0][273] , \round_in[0][272] , \round_in[0][271] ,
         \round_in[0][270] , \round_in[0][269] , \round_in[0][268] ,
         \round_in[0][267] , \round_in[0][266] , \round_in[0][265] ,
         \round_in[0][264] , \round_in[0][263] , \round_in[0][262] ,
         \round_in[0][261] , \round_in[0][260] , \round_in[0][259] ,
         \round_in[0][258] , \round_in[0][257] , \round_in[0][256] ,
         \round_in[0][255] , \round_in[0][254] , \round_in[0][253] ,
         \round_in[0][252] , \round_in[0][251] , \round_in[0][250] ,
         \round_in[0][249] , \round_in[0][248] , \round_in[0][247] ,
         \round_in[0][246] , \round_in[0][245] , \round_in[0][244] ,
         \round_in[0][243] , \round_in[0][242] , \round_in[0][241] ,
         \round_in[0][240] , \round_in[0][239] , \round_in[0][238] ,
         \round_in[0][237] , \round_in[0][236] , \round_in[0][235] ,
         \round_in[0][234] , \round_in[0][233] , \round_in[0][232] ,
         \round_in[0][231] , \round_in[0][230] , \round_in[0][229] ,
         \round_in[0][228] , \round_in[0][227] , \round_in[0][226] ,
         \round_in[0][225] , \round_in[0][224] , \round_in[0][223] ,
         \round_in[0][222] , \round_in[0][221] , \round_in[0][220] ,
         \round_in[0][219] , \round_in[0][218] , \round_in[0][217] ,
         \round_in[0][216] , \round_in[0][215] , \round_in[0][214] ,
         \round_in[0][213] , \round_in[0][212] , \round_in[0][211] ,
         \round_in[0][210] , \round_in[0][209] , \round_in[0][208] ,
         \round_in[0][207] , \round_in[0][206] , \round_in[0][205] ,
         \round_in[0][204] , \round_in[0][203] , \round_in[0][202] ,
         \round_in[0][201] , \round_in[0][200] , \round_in[0][199] ,
         \round_in[0][198] , \round_in[0][197] , \round_in[0][196] ,
         \round_in[0][195] , \round_in[0][194] , \round_in[0][193] ,
         \round_in[0][192] , \round_in[0][191] , \round_in[0][190] ,
         \round_in[0][189] , \round_in[0][188] , \round_in[0][187] ,
         \round_in[0][186] , \round_in[0][185] , \round_in[0][184] ,
         \round_in[0][183] , \round_in[0][182] , \round_in[0][181] ,
         \round_in[0][180] , \round_in[0][179] , \round_in[0][178] ,
         \round_in[0][177] , \round_in[0][176] , \round_in[0][175] ,
         \round_in[0][174] , \round_in[0][173] , \round_in[0][172] ,
         \round_in[0][171] , \round_in[0][170] , \round_in[0][169] ,
         \round_in[0][168] , \round_in[0][167] , \round_in[0][166] ,
         \round_in[0][165] , \round_in[0][164] , \round_in[0][163] ,
         \round_in[0][162] , \round_in[0][161] , \round_in[0][160] ,
         \round_in[0][159] , \round_in[0][158] , \round_in[0][157] ,
         \round_in[0][156] , \round_in[0][155] , \round_in[0][154] ,
         \round_in[0][153] , \round_in[0][152] , \round_in[0][151] ,
         \round_in[0][150] , \round_in[0][149] , \round_in[0][148] ,
         \round_in[0][147] , \round_in[0][146] , \round_in[0][145] ,
         \round_in[0][144] , \round_in[0][143] , \round_in[0][142] ,
         \round_in[0][141] , \round_in[0][140] , \round_in[0][139] ,
         \round_in[0][138] , \round_in[0][137] , \round_in[0][136] ,
         \round_in[0][135] , \round_in[0][134] , \round_in[0][133] ,
         \round_in[0][132] , \round_in[0][131] , \round_in[0][130] ,
         \round_in[0][129] , \round_in[0][128] , \round_in[0][127] ,
         \round_in[0][126] , \round_in[0][125] , \round_in[0][124] ,
         \round_in[0][123] , \round_in[0][122] , \round_in[0][121] ,
         \round_in[0][120] , \round_in[0][119] , \round_in[0][118] ,
         \round_in[0][117] , \round_in[0][116] , \round_in[0][115] ,
         \round_in[0][114] , \round_in[0][113] , \round_in[0][112] ,
         \round_in[0][111] , \round_in[0][110] , \round_in[0][109] ,
         \round_in[0][108] , \round_in[0][107] , \round_in[0][106] ,
         \round_in[0][105] , \round_in[0][104] , \round_in[0][103] ,
         \round_in[0][102] , \round_in[0][101] , \round_in[0][100] ,
         \round_in[0][99] , \round_in[0][98] , \round_in[0][97] ,
         \round_in[0][96] , \round_in[0][95] , \round_in[0][94] ,
         \round_in[0][93] , \round_in[0][92] , \round_in[0][91] ,
         \round_in[0][90] , \round_in[0][89] , \round_in[0][88] ,
         \round_in[0][87] , \round_in[0][86] , \round_in[0][85] ,
         \round_in[0][84] , \round_in[0][83] , \round_in[0][82] ,
         \round_in[0][81] , \round_in[0][80] , \round_in[0][79] ,
         \round_in[0][78] , \round_in[0][77] , \round_in[0][76] ,
         \round_in[0][75] , \round_in[0][74] , \round_in[0][73] ,
         \round_in[0][72] , \round_in[0][71] , \round_in[0][70] ,
         \round_in[0][69] , \round_in[0][68] , \round_in[0][67] ,
         \round_in[0][66] , \round_in[0][65] , \round_in[0][64] ,
         \round_in[0][63] , \round_in[0][62] , \round_in[0][61] ,
         \round_in[0][60] , \round_in[0][59] , \round_in[0][58] ,
         \round_in[0][57] , \round_in[0][56] , \round_in[0][55] ,
         \round_in[0][54] , \round_in[0][53] , \round_in[0][52] ,
         \round_in[0][51] , \round_in[0][50] , \round_in[0][49] ,
         \round_in[0][48] , \round_in[0][47] , \round_in[0][46] ,
         \round_in[0][45] , \round_in[0][44] , \round_in[0][43] ,
         \round_in[0][42] , \round_in[0][41] , \round_in[0][40] ,
         \round_in[0][39] , \round_in[0][38] , \round_in[0][37] ,
         \round_in[0][36] , \round_in[0][35] , \round_in[0][34] ,
         \round_in[0][33] , \round_in[0][32] , \round_in[0][31] ,
         \round_in[0][30] , \round_in[0][29] , \round_in[0][28] ,
         \round_in[0][27] , \round_in[0][26] , \round_in[0][25] ,
         \round_in[0][24] , \round_in[0][23] , \round_in[0][22] ,
         \round_in[0][21] , \round_in[0][20] , \round_in[0][19] ,
         \round_in[0][18] , \round_in[0][17] , \round_in[0][16] ,
         \round_in[0][15] , \round_in[0][14] , \round_in[0][13] ,
         \round_in[0][12] , \round_in[0][11] , \round_in[0][10] ,
         \round_in[0][9] , \round_in[0][8] , \round_in[0][7] ,
         \round_in[0][6] , \round_in[0][5] , \round_in[0][4] ,
         \round_in[0][3] , \round_in[0][2] , \round_in[0][1] ,
         \round_in[0][0] , \rc[3][63] , \rc[3][31] , \rc[3][15] , \rc[3][3] ,
         \rc[3][1] , \rc[2][0] , \rc[1][7] , \RCONST[0].rconst_/N67 ,
         \RCONST[0].rconst_/N56 , \RCONST[0].rconst_/N48 ,
         \RCONST[0].rconst_/N25 , \RCONST[0].rconst_/N17 ,
         \RCONST[1].rconst_/N68 , \RCONST[1].rconst_/N49 ,
         \RCONST[1].rconst_/N26 , \RCONST[1].rconst_/N15 ,
         \RCONST[2].rconst_/N57 , \RCONST[2].rconst_/N47 ,
         \RCONST[2].rconst_/N28 , \RCONST[2].rconst_/N18 ,
         \RCONST[3].rconst_/N10 , n1610, n1614, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008;
  wire   [5:0] rc_i;
  wire   [1599:0] round_reg;

  round_2 \ROUND[0].round_  ( .in({\round_in[0][1599] , \round_in[0][1598] , 
        \round_in[0][1597] , \round_in[0][1596] , \round_in[0][1595] , 
        \round_in[0][1594] , \round_in[0][1593] , \round_in[0][1592] , 
        \round_in[0][1591] , \round_in[0][1590] , \round_in[0][1589] , 
        \round_in[0][1588] , \round_in[0][1587] , \round_in[0][1586] , 
        \round_in[0][1585] , \round_in[0][1584] , \round_in[0][1583] , 
        \round_in[0][1582] , \round_in[0][1581] , \round_in[0][1580] , 
        \round_in[0][1579] , \round_in[0][1578] , \round_in[0][1577] , 
        \round_in[0][1576] , \round_in[0][1575] , \round_in[0][1574] , 
        \round_in[0][1573] , \round_in[0][1572] , \round_in[0][1571] , 
        \round_in[0][1570] , \round_in[0][1569] , \round_in[0][1568] , 
        \round_in[0][1567] , \round_in[0][1566] , \round_in[0][1565] , 
        \round_in[0][1564] , \round_in[0][1563] , \round_in[0][1562] , 
        \round_in[0][1561] , \round_in[0][1560] , \round_in[0][1559] , 
        \round_in[0][1558] , \round_in[0][1557] , \round_in[0][1556] , 
        \round_in[0][1555] , \round_in[0][1554] , \round_in[0][1553] , 
        \round_in[0][1552] , \round_in[0][1551] , \round_in[0][1550] , 
        \round_in[0][1549] , \round_in[0][1548] , \round_in[0][1547] , 
        \round_in[0][1546] , \round_in[0][1545] , \round_in[0][1544] , 
        \round_in[0][1543] , \round_in[0][1542] , \round_in[0][1541] , 
        \round_in[0][1540] , \round_in[0][1539] , \round_in[0][1538] , 
        \round_in[0][1537] , \round_in[0][1536] , \round_in[0][1535] , 
        \round_in[0][1534] , \round_in[0][1533] , \round_in[0][1532] , 
        \round_in[0][1531] , \round_in[0][1530] , \round_in[0][1529] , 
        \round_in[0][1528] , \round_in[0][1527] , \round_in[0][1526] , 
        \round_in[0][1525] , \round_in[0][1524] , \round_in[0][1523] , 
        \round_in[0][1522] , \round_in[0][1521] , \round_in[0][1520] , 
        \round_in[0][1519] , \round_in[0][1518] , \round_in[0][1517] , 
        \round_in[0][1516] , \round_in[0][1515] , \round_in[0][1514] , 
        \round_in[0][1513] , \round_in[0][1512] , \round_in[0][1511] , 
        \round_in[0][1510] , \round_in[0][1509] , \round_in[0][1508] , 
        \round_in[0][1507] , \round_in[0][1506] , \round_in[0][1505] , 
        \round_in[0][1504] , \round_in[0][1503] , \round_in[0][1502] , 
        \round_in[0][1501] , \round_in[0][1500] , \round_in[0][1499] , 
        \round_in[0][1498] , \round_in[0][1497] , \round_in[0][1496] , 
        \round_in[0][1495] , \round_in[0][1494] , \round_in[0][1493] , 
        \round_in[0][1492] , \round_in[0][1491] , \round_in[0][1490] , 
        \round_in[0][1489] , \round_in[0][1488] , \round_in[0][1487] , 
        \round_in[0][1486] , \round_in[0][1485] , \round_in[0][1484] , 
        \round_in[0][1483] , \round_in[0][1482] , \round_in[0][1481] , 
        \round_in[0][1480] , \round_in[0][1479] , \round_in[0][1478] , 
        \round_in[0][1477] , \round_in[0][1476] , \round_in[0][1475] , 
        \round_in[0][1474] , \round_in[0][1473] , \round_in[0][1472] , 
        \round_in[0][1471] , \round_in[0][1470] , \round_in[0][1469] , 
        \round_in[0][1468] , \round_in[0][1467] , \round_in[0][1466] , 
        \round_in[0][1465] , \round_in[0][1464] , \round_in[0][1463] , 
        \round_in[0][1462] , \round_in[0][1461] , \round_in[0][1460] , 
        \round_in[0][1459] , \round_in[0][1458] , \round_in[0][1457] , 
        \round_in[0][1456] , \round_in[0][1455] , \round_in[0][1454] , 
        \round_in[0][1453] , \round_in[0][1452] , \round_in[0][1451] , 
        \round_in[0][1450] , \round_in[0][1449] , \round_in[0][1448] , 
        \round_in[0][1447] , \round_in[0][1446] , \round_in[0][1445] , 
        \round_in[0][1444] , \round_in[0][1443] , \round_in[0][1442] , 
        \round_in[0][1441] , \round_in[0][1440] , \round_in[0][1439] , 
        \round_in[0][1438] , \round_in[0][1437] , \round_in[0][1436] , 
        \round_in[0][1435] , \round_in[0][1434] , \round_in[0][1433] , 
        \round_in[0][1432] , \round_in[0][1431] , \round_in[0][1430] , 
        \round_in[0][1429] , \round_in[0][1428] , \round_in[0][1427] , 
        \round_in[0][1426] , \round_in[0][1425] , \round_in[0][1424] , 
        \round_in[0][1423] , \round_in[0][1422] , \round_in[0][1421] , 
        \round_in[0][1420] , \round_in[0][1419] , \round_in[0][1418] , 
        \round_in[0][1417] , \round_in[0][1416] , \round_in[0][1415] , 
        \round_in[0][1414] , \round_in[0][1413] , \round_in[0][1412] , 
        \round_in[0][1411] , \round_in[0][1410] , \round_in[0][1409] , 
        \round_in[0][1408] , \round_in[0][1407] , \round_in[0][1406] , 
        \round_in[0][1405] , \round_in[0][1404] , \round_in[0][1403] , 
        \round_in[0][1402] , \round_in[0][1401] , \round_in[0][1400] , 
        \round_in[0][1399] , \round_in[0][1398] , \round_in[0][1397] , 
        \round_in[0][1396] , \round_in[0][1395] , \round_in[0][1394] , 
        \round_in[0][1393] , \round_in[0][1392] , \round_in[0][1391] , 
        \round_in[0][1390] , \round_in[0][1389] , \round_in[0][1388] , 
        \round_in[0][1387] , \round_in[0][1386] , \round_in[0][1385] , 
        \round_in[0][1384] , \round_in[0][1383] , \round_in[0][1382] , 
        \round_in[0][1381] , \round_in[0][1380] , \round_in[0][1379] , 
        \round_in[0][1378] , \round_in[0][1377] , \round_in[0][1376] , 
        \round_in[0][1375] , \round_in[0][1374] , \round_in[0][1373] , 
        \round_in[0][1372] , \round_in[0][1371] , \round_in[0][1370] , 
        \round_in[0][1369] , \round_in[0][1368] , \round_in[0][1367] , 
        \round_in[0][1366] , \round_in[0][1365] , \round_in[0][1364] , 
        \round_in[0][1363] , \round_in[0][1362] , \round_in[0][1361] , 
        \round_in[0][1360] , \round_in[0][1359] , \round_in[0][1358] , 
        \round_in[0][1357] , \round_in[0][1356] , \round_in[0][1355] , 
        \round_in[0][1354] , \round_in[0][1353] , \round_in[0][1352] , 
        \round_in[0][1351] , \round_in[0][1350] , \round_in[0][1349] , 
        \round_in[0][1348] , \round_in[0][1347] , \round_in[0][1346] , 
        \round_in[0][1345] , \round_in[0][1344] , \round_in[0][1343] , 
        \round_in[0][1342] , \round_in[0][1341] , \round_in[0][1340] , 
        \round_in[0][1339] , \round_in[0][1338] , \round_in[0][1337] , 
        \round_in[0][1336] , \round_in[0][1335] , \round_in[0][1334] , 
        \round_in[0][1333] , \round_in[0][1332] , \round_in[0][1331] , 
        \round_in[0][1330] , \round_in[0][1329] , \round_in[0][1328] , 
        \round_in[0][1327] , \round_in[0][1326] , \round_in[0][1325] , 
        \round_in[0][1324] , \round_in[0][1323] , \round_in[0][1322] , 
        \round_in[0][1321] , \round_in[0][1320] , \round_in[0][1319] , 
        \round_in[0][1318] , \round_in[0][1317] , \round_in[0][1316] , 
        \round_in[0][1315] , \round_in[0][1314] , \round_in[0][1313] , 
        \round_in[0][1312] , \round_in[0][1311] , \round_in[0][1310] , 
        \round_in[0][1309] , \round_in[0][1308] , \round_in[0][1307] , 
        \round_in[0][1306] , \round_in[0][1305] , \round_in[0][1304] , 
        \round_in[0][1303] , \round_in[0][1302] , \round_in[0][1301] , 
        \round_in[0][1300] , \round_in[0][1299] , \round_in[0][1298] , 
        \round_in[0][1297] , \round_in[0][1296] , \round_in[0][1295] , 
        \round_in[0][1294] , \round_in[0][1293] , \round_in[0][1292] , 
        \round_in[0][1291] , \round_in[0][1290] , \round_in[0][1289] , 
        \round_in[0][1288] , \round_in[0][1287] , \round_in[0][1286] , 
        \round_in[0][1285] , \round_in[0][1284] , \round_in[0][1283] , 
        \round_in[0][1282] , \round_in[0][1281] , \round_in[0][1280] , 
        \round_in[0][1279] , \round_in[0][1278] , \round_in[0][1277] , 
        \round_in[0][1276] , \round_in[0][1275] , \round_in[0][1274] , 
        \round_in[0][1273] , \round_in[0][1272] , \round_in[0][1271] , 
        \round_in[0][1270] , \round_in[0][1269] , \round_in[0][1268] , 
        \round_in[0][1267] , \round_in[0][1266] , \round_in[0][1265] , 
        \round_in[0][1264] , \round_in[0][1263] , \round_in[0][1262] , 
        \round_in[0][1261] , \round_in[0][1260] , \round_in[0][1259] , 
        \round_in[0][1258] , \round_in[0][1257] , \round_in[0][1256] , 
        \round_in[0][1255] , \round_in[0][1254] , \round_in[0][1253] , 
        \round_in[0][1252] , \round_in[0][1251] , \round_in[0][1250] , 
        \round_in[0][1249] , \round_in[0][1248] , \round_in[0][1247] , 
        \round_in[0][1246] , \round_in[0][1245] , \round_in[0][1244] , 
        \round_in[0][1243] , \round_in[0][1242] , \round_in[0][1241] , 
        \round_in[0][1240] , \round_in[0][1239] , \round_in[0][1238] , 
        \round_in[0][1237] , \round_in[0][1236] , \round_in[0][1235] , 
        \round_in[0][1234] , \round_in[0][1233] , \round_in[0][1232] , 
        \round_in[0][1231] , \round_in[0][1230] , \round_in[0][1229] , 
        \round_in[0][1228] , \round_in[0][1227] , \round_in[0][1226] , 
        \round_in[0][1225] , \round_in[0][1224] , \round_in[0][1223] , 
        \round_in[0][1222] , \round_in[0][1221] , \round_in[0][1220] , 
        \round_in[0][1219] , \round_in[0][1218] , \round_in[0][1217] , 
        \round_in[0][1216] , \round_in[0][1215] , \round_in[0][1214] , 
        \round_in[0][1213] , \round_in[0][1212] , \round_in[0][1211] , 
        \round_in[0][1210] , \round_in[0][1209] , \round_in[0][1208] , 
        \round_in[0][1207] , \round_in[0][1206] , \round_in[0][1205] , 
        \round_in[0][1204] , \round_in[0][1203] , \round_in[0][1202] , 
        \round_in[0][1201] , \round_in[0][1200] , \round_in[0][1199] , 
        \round_in[0][1198] , \round_in[0][1197] , \round_in[0][1196] , 
        \round_in[0][1195] , \round_in[0][1194] , \round_in[0][1193] , 
        \round_in[0][1192] , \round_in[0][1191] , \round_in[0][1190] , 
        \round_in[0][1189] , \round_in[0][1188] , \round_in[0][1187] , 
        \round_in[0][1186] , \round_in[0][1185] , \round_in[0][1184] , 
        \round_in[0][1183] , \round_in[0][1182] , \round_in[0][1181] , 
        \round_in[0][1180] , \round_in[0][1179] , \round_in[0][1178] , 
        \round_in[0][1177] , \round_in[0][1176] , \round_in[0][1175] , 
        \round_in[0][1174] , \round_in[0][1173] , \round_in[0][1172] , 
        \round_in[0][1171] , \round_in[0][1170] , \round_in[0][1169] , 
        \round_in[0][1168] , \round_in[0][1167] , \round_in[0][1166] , 
        \round_in[0][1165] , \round_in[0][1164] , \round_in[0][1163] , 
        \round_in[0][1162] , \round_in[0][1161] , \round_in[0][1160] , 
        \round_in[0][1159] , \round_in[0][1158] , \round_in[0][1157] , 
        \round_in[0][1156] , \round_in[0][1155] , \round_in[0][1154] , 
        \round_in[0][1153] , \round_in[0][1152] , \round_in[0][1151] , 
        \round_in[0][1150] , \round_in[0][1149] , \round_in[0][1148] , 
        \round_in[0][1147] , \round_in[0][1146] , \round_in[0][1145] , 
        \round_in[0][1144] , \round_in[0][1143] , \round_in[0][1142] , 
        \round_in[0][1141] , \round_in[0][1140] , \round_in[0][1139] , 
        \round_in[0][1138] , \round_in[0][1137] , \round_in[0][1136] , 
        \round_in[0][1135] , \round_in[0][1134] , \round_in[0][1133] , 
        \round_in[0][1132] , \round_in[0][1131] , \round_in[0][1130] , 
        \round_in[0][1129] , \round_in[0][1128] , \round_in[0][1127] , 
        \round_in[0][1126] , \round_in[0][1125] , \round_in[0][1124] , 
        \round_in[0][1123] , \round_in[0][1122] , \round_in[0][1121] , 
        \round_in[0][1120] , \round_in[0][1119] , \round_in[0][1118] , 
        \round_in[0][1117] , \round_in[0][1116] , \round_in[0][1115] , 
        \round_in[0][1114] , \round_in[0][1113] , \round_in[0][1112] , 
        \round_in[0][1111] , \round_in[0][1110] , \round_in[0][1109] , 
        \round_in[0][1108] , \round_in[0][1107] , \round_in[0][1106] , 
        \round_in[0][1105] , \round_in[0][1104] , \round_in[0][1103] , 
        \round_in[0][1102] , \round_in[0][1101] , \round_in[0][1100] , 
        \round_in[0][1099] , \round_in[0][1098] , \round_in[0][1097] , 
        \round_in[0][1096] , \round_in[0][1095] , \round_in[0][1094] , 
        \round_in[0][1093] , \round_in[0][1092] , \round_in[0][1091] , 
        \round_in[0][1090] , \round_in[0][1089] , \round_in[0][1088] , 
        \round_in[0][1087] , \round_in[0][1086] , \round_in[0][1085] , 
        \round_in[0][1084] , \round_in[0][1083] , \round_in[0][1082] , 
        \round_in[0][1081] , \round_in[0][1080] , \round_in[0][1079] , 
        \round_in[0][1078] , \round_in[0][1077] , \round_in[0][1076] , 
        \round_in[0][1075] , \round_in[0][1074] , \round_in[0][1073] , 
        \round_in[0][1072] , \round_in[0][1071] , \round_in[0][1070] , 
        \round_in[0][1069] , \round_in[0][1068] , \round_in[0][1067] , 
        \round_in[0][1066] , \round_in[0][1065] , \round_in[0][1064] , 
        \round_in[0][1063] , \round_in[0][1062] , \round_in[0][1061] , 
        \round_in[0][1060] , \round_in[0][1059] , \round_in[0][1058] , 
        \round_in[0][1057] , \round_in[0][1056] , \round_in[0][1055] , 
        \round_in[0][1054] , \round_in[0][1053] , \round_in[0][1052] , 
        \round_in[0][1051] , \round_in[0][1050] , \round_in[0][1049] , 
        \round_in[0][1048] , \round_in[0][1047] , \round_in[0][1046] , 
        \round_in[0][1045] , \round_in[0][1044] , \round_in[0][1043] , 
        \round_in[0][1042] , \round_in[0][1041] , \round_in[0][1040] , 
        \round_in[0][1039] , \round_in[0][1038] , \round_in[0][1037] , 
        \round_in[0][1036] , \round_in[0][1035] , \round_in[0][1034] , 
        \round_in[0][1033] , \round_in[0][1032] , \round_in[0][1031] , 
        \round_in[0][1030] , \round_in[0][1029] , \round_in[0][1028] , 
        \round_in[0][1027] , \round_in[0][1026] , \round_in[0][1025] , 
        \round_in[0][1024] , \round_in[0][1023] , \round_in[0][1022] , 
        \round_in[0][1021] , \round_in[0][1020] , \round_in[0][1019] , 
        \round_in[0][1018] , \round_in[0][1017] , \round_in[0][1016] , 
        \round_in[0][1015] , \round_in[0][1014] , \round_in[0][1013] , 
        \round_in[0][1012] , \round_in[0][1011] , \round_in[0][1010] , 
        \round_in[0][1009] , \round_in[0][1008] , \round_in[0][1007] , 
        \round_in[0][1006] , \round_in[0][1005] , \round_in[0][1004] , 
        \round_in[0][1003] , \round_in[0][1002] , \round_in[0][1001] , 
        \round_in[0][1000] , \round_in[0][999] , \round_in[0][998] , 
        \round_in[0][997] , \round_in[0][996] , \round_in[0][995] , 
        \round_in[0][994] , \round_in[0][993] , \round_in[0][992] , 
        \round_in[0][991] , \round_in[0][990] , \round_in[0][989] , 
        \round_in[0][988] , \round_in[0][987] , \round_in[0][986] , 
        \round_in[0][985] , \round_in[0][984] , \round_in[0][983] , 
        \round_in[0][982] , \round_in[0][981] , \round_in[0][980] , 
        \round_in[0][979] , \round_in[0][978] , \round_in[0][977] , 
        \round_in[0][976] , \round_in[0][975] , \round_in[0][974] , 
        \round_in[0][973] , \round_in[0][972] , \round_in[0][971] , 
        \round_in[0][970] , \round_in[0][969] , \round_in[0][968] , 
        \round_in[0][967] , \round_in[0][966] , \round_in[0][965] , 
        \round_in[0][964] , \round_in[0][963] , \round_in[0][962] , 
        \round_in[0][961] , \round_in[0][960] , \round_in[0][959] , 
        \round_in[0][958] , \round_in[0][957] , \round_in[0][956] , 
        \round_in[0][955] , \round_in[0][954] , \round_in[0][953] , 
        \round_in[0][952] , \round_in[0][951] , \round_in[0][950] , 
        \round_in[0][949] , \round_in[0][948] , \round_in[0][947] , 
        \round_in[0][946] , \round_in[0][945] , \round_in[0][944] , 
        \round_in[0][943] , \round_in[0][942] , \round_in[0][941] , 
        \round_in[0][940] , \round_in[0][939] , \round_in[0][938] , 
        \round_in[0][937] , \round_in[0][936] , \round_in[0][935] , 
        \round_in[0][934] , \round_in[0][933] , \round_in[0][932] , 
        \round_in[0][931] , \round_in[0][930] , \round_in[0][929] , 
        \round_in[0][928] , \round_in[0][927] , \round_in[0][926] , 
        \round_in[0][925] , \round_in[0][924] , \round_in[0][923] , 
        \round_in[0][922] , \round_in[0][921] , \round_in[0][920] , 
        \round_in[0][919] , \round_in[0][918] , \round_in[0][917] , 
        \round_in[0][916] , \round_in[0][915] , \round_in[0][914] , 
        \round_in[0][913] , \round_in[0][912] , \round_in[0][911] , 
        \round_in[0][910] , \round_in[0][909] , \round_in[0][908] , 
        \round_in[0][907] , \round_in[0][906] , \round_in[0][905] , 
        \round_in[0][904] , \round_in[0][903] , \round_in[0][902] , 
        \round_in[0][901] , \round_in[0][900] , \round_in[0][899] , 
        \round_in[0][898] , \round_in[0][897] , \round_in[0][896] , 
        \round_in[0][895] , \round_in[0][894] , \round_in[0][893] , 
        \round_in[0][892] , \round_in[0][891] , \round_in[0][890] , 
        \round_in[0][889] , \round_in[0][888] , \round_in[0][887] , 
        \round_in[0][886] , \round_in[0][885] , \round_in[0][884] , 
        \round_in[0][883] , \round_in[0][882] , \round_in[0][881] , 
        \round_in[0][880] , \round_in[0][879] , \round_in[0][878] , 
        \round_in[0][877] , \round_in[0][876] , \round_in[0][875] , 
        \round_in[0][874] , \round_in[0][873] , \round_in[0][872] , 
        \round_in[0][871] , \round_in[0][870] , \round_in[0][869] , 
        \round_in[0][868] , \round_in[0][867] , \round_in[0][866] , 
        \round_in[0][865] , \round_in[0][864] , \round_in[0][863] , 
        \round_in[0][862] , \round_in[0][861] , \round_in[0][860] , 
        \round_in[0][859] , \round_in[0][858] , \round_in[0][857] , 
        \round_in[0][856] , \round_in[0][855] , \round_in[0][854] , 
        \round_in[0][853] , \round_in[0][852] , \round_in[0][851] , 
        \round_in[0][850] , \round_in[0][849] , \round_in[0][848] , 
        \round_in[0][847] , \round_in[0][846] , \round_in[0][845] , 
        \round_in[0][844] , \round_in[0][843] , \round_in[0][842] , 
        \round_in[0][841] , \round_in[0][840] , \round_in[0][839] , 
        \round_in[0][838] , \round_in[0][837] , \round_in[0][836] , 
        \round_in[0][835] , \round_in[0][834] , \round_in[0][833] , 
        \round_in[0][832] , \round_in[0][831] , \round_in[0][830] , 
        \round_in[0][829] , \round_in[0][828] , \round_in[0][827] , 
        \round_in[0][826] , \round_in[0][825] , \round_in[0][824] , 
        \round_in[0][823] , \round_in[0][822] , \round_in[0][821] , 
        \round_in[0][820] , \round_in[0][819] , \round_in[0][818] , 
        \round_in[0][817] , \round_in[0][816] , \round_in[0][815] , 
        \round_in[0][814] , \round_in[0][813] , \round_in[0][812] , 
        \round_in[0][811] , \round_in[0][810] , \round_in[0][809] , 
        \round_in[0][808] , \round_in[0][807] , \round_in[0][806] , 
        \round_in[0][805] , \round_in[0][804] , \round_in[0][803] , 
        \round_in[0][802] , \round_in[0][801] , \round_in[0][800] , 
        \round_in[0][799] , \round_in[0][798] , \round_in[0][797] , 
        \round_in[0][796] , \round_in[0][795] , \round_in[0][794] , 
        \round_in[0][793] , \round_in[0][792] , \round_in[0][791] , 
        \round_in[0][790] , \round_in[0][789] , \round_in[0][788] , 
        \round_in[0][787] , \round_in[0][786] , \round_in[0][785] , 
        \round_in[0][784] , \round_in[0][783] , \round_in[0][782] , 
        \round_in[0][781] , \round_in[0][780] , \round_in[0][779] , 
        \round_in[0][778] , \round_in[0][777] , \round_in[0][776] , 
        \round_in[0][775] , \round_in[0][774] , \round_in[0][773] , 
        \round_in[0][772] , \round_in[0][771] , \round_in[0][770] , 
        \round_in[0][769] , \round_in[0][768] , \round_in[0][767] , 
        \round_in[0][766] , \round_in[0][765] , \round_in[0][764] , 
        \round_in[0][763] , \round_in[0][762] , \round_in[0][761] , 
        \round_in[0][760] , \round_in[0][759] , \round_in[0][758] , 
        \round_in[0][757] , \round_in[0][756] , \round_in[0][755] , 
        \round_in[0][754] , \round_in[0][753] , \round_in[0][752] , 
        \round_in[0][751] , \round_in[0][750] , \round_in[0][749] , 
        \round_in[0][748] , \round_in[0][747] , \round_in[0][746] , 
        \round_in[0][745] , \round_in[0][744] , \round_in[0][743] , 
        \round_in[0][742] , \round_in[0][741] , \round_in[0][740] , 
        \round_in[0][739] , \round_in[0][738] , \round_in[0][737] , 
        \round_in[0][736] , \round_in[0][735] , \round_in[0][734] , 
        \round_in[0][733] , \round_in[0][732] , \round_in[0][731] , 
        \round_in[0][730] , \round_in[0][729] , \round_in[0][728] , 
        \round_in[0][727] , \round_in[0][726] , \round_in[0][725] , 
        \round_in[0][724] , \round_in[0][723] , \round_in[0][722] , 
        \round_in[0][721] , \round_in[0][720] , \round_in[0][719] , 
        \round_in[0][718] , \round_in[0][717] , \round_in[0][716] , 
        \round_in[0][715] , \round_in[0][714] , \round_in[0][713] , 
        \round_in[0][712] , \round_in[0][711] , \round_in[0][710] , 
        \round_in[0][709] , \round_in[0][708] , \round_in[0][707] , 
        \round_in[0][706] , \round_in[0][705] , \round_in[0][704] , 
        \round_in[0][703] , \round_in[0][702] , \round_in[0][701] , 
        \round_in[0][700] , \round_in[0][699] , \round_in[0][698] , 
        \round_in[0][697] , \round_in[0][696] , \round_in[0][695] , 
        \round_in[0][694] , \round_in[0][693] , \round_in[0][692] , 
        \round_in[0][691] , \round_in[0][690] , \round_in[0][689] , 
        \round_in[0][688] , \round_in[0][687] , \round_in[0][686] , 
        \round_in[0][685] , \round_in[0][684] , \round_in[0][683] , 
        \round_in[0][682] , \round_in[0][681] , \round_in[0][680] , 
        \round_in[0][679] , \round_in[0][678] , \round_in[0][677] , 
        \round_in[0][676] , \round_in[0][675] , \round_in[0][674] , 
        \round_in[0][673] , \round_in[0][672] , \round_in[0][671] , 
        \round_in[0][670] , \round_in[0][669] , \round_in[0][668] , 
        \round_in[0][667] , \round_in[0][666] , \round_in[0][665] , 
        \round_in[0][664] , \round_in[0][663] , \round_in[0][662] , 
        \round_in[0][661] , \round_in[0][660] , \round_in[0][659] , 
        \round_in[0][658] , \round_in[0][657] , \round_in[0][656] , 
        \round_in[0][655] , \round_in[0][654] , \round_in[0][653] , 
        \round_in[0][652] , \round_in[0][651] , \round_in[0][650] , 
        \round_in[0][649] , \round_in[0][648] , \round_in[0][647] , 
        \round_in[0][646] , \round_in[0][645] , \round_in[0][644] , 
        \round_in[0][643] , \round_in[0][642] , \round_in[0][641] , 
        \round_in[0][640] , \round_in[0][639] , \round_in[0][638] , 
        \round_in[0][637] , \round_in[0][636] , \round_in[0][635] , 
        \round_in[0][634] , \round_in[0][633] , \round_in[0][632] , 
        \round_in[0][631] , \round_in[0][630] , \round_in[0][629] , 
        \round_in[0][628] , \round_in[0][627] , \round_in[0][626] , 
        \round_in[0][625] , \round_in[0][624] , \round_in[0][623] , 
        \round_in[0][622] , \round_in[0][621] , \round_in[0][620] , 
        \round_in[0][619] , \round_in[0][618] , \round_in[0][617] , 
        \round_in[0][616] , \round_in[0][615] , \round_in[0][614] , 
        \round_in[0][613] , \round_in[0][612] , \round_in[0][611] , 
        \round_in[0][610] , \round_in[0][609] , \round_in[0][608] , 
        \round_in[0][607] , \round_in[0][606] , \round_in[0][605] , 
        \round_in[0][604] , \round_in[0][603] , \round_in[0][602] , 
        \round_in[0][601] , \round_in[0][600] , \round_in[0][599] , 
        \round_in[0][598] , \round_in[0][597] , \round_in[0][596] , 
        \round_in[0][595] , \round_in[0][594] , \round_in[0][593] , 
        \round_in[0][592] , \round_in[0][591] , \round_in[0][590] , 
        \round_in[0][589] , \round_in[0][588] , \round_in[0][587] , 
        \round_in[0][586] , \round_in[0][585] , \round_in[0][584] , 
        \round_in[0][583] , \round_in[0][582] , \round_in[0][581] , 
        \round_in[0][580] , \round_in[0][579] , \round_in[0][578] , 
        \round_in[0][577] , \round_in[0][576] , \round_in[0][575] , 
        \round_in[0][574] , \round_in[0][573] , \round_in[0][572] , 
        \round_in[0][571] , \round_in[0][570] , \round_in[0][569] , 
        \round_in[0][568] , \round_in[0][567] , \round_in[0][566] , 
        \round_in[0][565] , \round_in[0][564] , \round_in[0][563] , 
        \round_in[0][562] , \round_in[0][561] , \round_in[0][560] , 
        \round_in[0][559] , \round_in[0][558] , \round_in[0][557] , 
        \round_in[0][556] , \round_in[0][555] , \round_in[0][554] , 
        \round_in[0][553] , \round_in[0][552] , \round_in[0][551] , 
        \round_in[0][550] , \round_in[0][549] , \round_in[0][548] , 
        \round_in[0][547] , \round_in[0][546] , \round_in[0][545] , 
        \round_in[0][544] , \round_in[0][543] , \round_in[0][542] , 
        \round_in[0][541] , \round_in[0][540] , \round_in[0][539] , 
        \round_in[0][538] , \round_in[0][537] , \round_in[0][536] , 
        \round_in[0][535] , \round_in[0][534] , \round_in[0][533] , 
        \round_in[0][532] , \round_in[0][531] , \round_in[0][530] , 
        \round_in[0][529] , \round_in[0][528] , \round_in[0][527] , 
        \round_in[0][526] , \round_in[0][525] , \round_in[0][524] , 
        \round_in[0][523] , \round_in[0][522] , \round_in[0][521] , 
        \round_in[0][520] , \round_in[0][519] , \round_in[0][518] , 
        \round_in[0][517] , \round_in[0][516] , \round_in[0][515] , 
        \round_in[0][514] , \round_in[0][513] , \round_in[0][512] , 
        \round_in[0][511] , \round_in[0][510] , \round_in[0][509] , 
        \round_in[0][508] , \round_in[0][507] , \round_in[0][506] , 
        \round_in[0][505] , \round_in[0][504] , \round_in[0][503] , 
        \round_in[0][502] , \round_in[0][501] , \round_in[0][500] , 
        \round_in[0][499] , \round_in[0][498] , \round_in[0][497] , 
        \round_in[0][496] , \round_in[0][495] , \round_in[0][494] , 
        \round_in[0][493] , \round_in[0][492] , \round_in[0][491] , 
        \round_in[0][490] , \round_in[0][489] , \round_in[0][488] , 
        \round_in[0][487] , \round_in[0][486] , \round_in[0][485] , 
        \round_in[0][484] , \round_in[0][483] , \round_in[0][482] , 
        \round_in[0][481] , \round_in[0][480] , \round_in[0][479] , 
        \round_in[0][478] , \round_in[0][477] , \round_in[0][476] , 
        \round_in[0][475] , \round_in[0][474] , \round_in[0][473] , 
        \round_in[0][472] , \round_in[0][471] , \round_in[0][470] , 
        \round_in[0][469] , \round_in[0][468] , \round_in[0][467] , 
        \round_in[0][466] , \round_in[0][465] , \round_in[0][464] , 
        \round_in[0][463] , \round_in[0][462] , \round_in[0][461] , 
        \round_in[0][460] , \round_in[0][459] , \round_in[0][458] , 
        \round_in[0][457] , \round_in[0][456] , \round_in[0][455] , 
        \round_in[0][454] , \round_in[0][453] , \round_in[0][452] , 
        \round_in[0][451] , \round_in[0][450] , \round_in[0][449] , 
        \round_in[0][448] , \round_in[0][447] , \round_in[0][446] , 
        \round_in[0][445] , \round_in[0][444] , \round_in[0][443] , 
        \round_in[0][442] , \round_in[0][441] , \round_in[0][440] , 
        \round_in[0][439] , \round_in[0][438] , \round_in[0][437] , 
        \round_in[0][436] , \round_in[0][435] , \round_in[0][434] , 
        \round_in[0][433] , \round_in[0][432] , \round_in[0][431] , 
        \round_in[0][430] , \round_in[0][429] , \round_in[0][428] , 
        \round_in[0][427] , \round_in[0][426] , \round_in[0][425] , 
        \round_in[0][424] , \round_in[0][423] , \round_in[0][422] , 
        \round_in[0][421] , \round_in[0][420] , \round_in[0][419] , 
        \round_in[0][418] , \round_in[0][417] , \round_in[0][416] , 
        \round_in[0][415] , \round_in[0][414] , \round_in[0][413] , 
        \round_in[0][412] , \round_in[0][411] , \round_in[0][410] , 
        \round_in[0][409] , \round_in[0][408] , \round_in[0][407] , 
        \round_in[0][406] , \round_in[0][405] , \round_in[0][404] , 
        \round_in[0][403] , \round_in[0][402] , \round_in[0][401] , 
        \round_in[0][400] , \round_in[0][399] , \round_in[0][398] , 
        \round_in[0][397] , \round_in[0][396] , \round_in[0][395] , 
        \round_in[0][394] , \round_in[0][393] , \round_in[0][392] , 
        \round_in[0][391] , \round_in[0][390] , \round_in[0][389] , 
        \round_in[0][388] , \round_in[0][387] , \round_in[0][386] , 
        \round_in[0][385] , \round_in[0][384] , \round_in[0][383] , 
        \round_in[0][382] , \round_in[0][381] , \round_in[0][380] , 
        \round_in[0][379] , \round_in[0][378] , \round_in[0][377] , 
        \round_in[0][376] , \round_in[0][375] , \round_in[0][374] , 
        \round_in[0][373] , \round_in[0][372] , \round_in[0][371] , 
        \round_in[0][370] , \round_in[0][369] , \round_in[0][368] , 
        \round_in[0][367] , \round_in[0][366] , \round_in[0][365] , 
        \round_in[0][364] , \round_in[0][363] , \round_in[0][362] , 
        \round_in[0][361] , \round_in[0][360] , \round_in[0][359] , 
        \round_in[0][358] , \round_in[0][357] , \round_in[0][356] , 
        \round_in[0][355] , \round_in[0][354] , \round_in[0][353] , 
        \round_in[0][352] , \round_in[0][351] , \round_in[0][350] , 
        \round_in[0][349] , \round_in[0][348] , \round_in[0][347] , 
        \round_in[0][346] , \round_in[0][345] , \round_in[0][344] , 
        \round_in[0][343] , \round_in[0][342] , \round_in[0][341] , 
        \round_in[0][340] , \round_in[0][339] , \round_in[0][338] , 
        \round_in[0][337] , \round_in[0][336] , \round_in[0][335] , 
        \round_in[0][334] , \round_in[0][333] , \round_in[0][332] , 
        \round_in[0][331] , \round_in[0][330] , \round_in[0][329] , 
        \round_in[0][328] , \round_in[0][327] , \round_in[0][326] , 
        \round_in[0][325] , \round_in[0][324] , \round_in[0][323] , 
        \round_in[0][322] , \round_in[0][321] , \round_in[0][320] , 
        \round_in[0][319] , \round_in[0][318] , \round_in[0][317] , 
        \round_in[0][316] , \round_in[0][315] , \round_in[0][314] , 
        \round_in[0][313] , \round_in[0][312] , \round_in[0][311] , 
        \round_in[0][310] , \round_in[0][309] , \round_in[0][308] , 
        \round_in[0][307] , \round_in[0][306] , \round_in[0][305] , 
        \round_in[0][304] , \round_in[0][303] , \round_in[0][302] , 
        \round_in[0][301] , \round_in[0][300] , \round_in[0][299] , 
        \round_in[0][298] , \round_in[0][297] , \round_in[0][296] , 
        \round_in[0][295] , \round_in[0][294] , \round_in[0][293] , 
        \round_in[0][292] , \round_in[0][291] , \round_in[0][290] , 
        \round_in[0][289] , \round_in[0][288] , \round_in[0][287] , 
        \round_in[0][286] , \round_in[0][285] , \round_in[0][284] , 
        \round_in[0][283] , \round_in[0][282] , \round_in[0][281] , 
        \round_in[0][280] , \round_in[0][279] , \round_in[0][278] , 
        \round_in[0][277] , \round_in[0][276] , \round_in[0][275] , 
        \round_in[0][274] , \round_in[0][273] , \round_in[0][272] , 
        \round_in[0][271] , \round_in[0][270] , \round_in[0][269] , 
        \round_in[0][268] , \round_in[0][267] , \round_in[0][266] , 
        \round_in[0][265] , \round_in[0][264] , \round_in[0][263] , 
        \round_in[0][262] , \round_in[0][261] , \round_in[0][260] , 
        \round_in[0][259] , \round_in[0][258] , \round_in[0][257] , 
        \round_in[0][256] , \round_in[0][255] , \round_in[0][254] , 
        \round_in[0][253] , \round_in[0][252] , \round_in[0][251] , 
        \round_in[0][250] , \round_in[0][249] , \round_in[0][248] , 
        \round_in[0][247] , \round_in[0][246] , \round_in[0][245] , 
        \round_in[0][244] , \round_in[0][243] , \round_in[0][242] , 
        \round_in[0][241] , \round_in[0][240] , \round_in[0][239] , 
        \round_in[0][238] , \round_in[0][237] , \round_in[0][236] , 
        \round_in[0][235] , \round_in[0][234] , \round_in[0][233] , 
        \round_in[0][232] , \round_in[0][231] , \round_in[0][230] , 
        \round_in[0][229] , \round_in[0][228] , \round_in[0][227] , 
        \round_in[0][226] , \round_in[0][225] , \round_in[0][224] , 
        \round_in[0][223] , \round_in[0][222] , \round_in[0][221] , 
        \round_in[0][220] , \round_in[0][219] , \round_in[0][218] , 
        \round_in[0][217] , \round_in[0][216] , \round_in[0][215] , 
        \round_in[0][214] , \round_in[0][213] , \round_in[0][212] , 
        \round_in[0][211] , \round_in[0][210] , \round_in[0][209] , 
        \round_in[0][208] , \round_in[0][207] , \round_in[0][206] , 
        \round_in[0][205] , \round_in[0][204] , \round_in[0][203] , 
        \round_in[0][202] , \round_in[0][201] , \round_in[0][200] , 
        \round_in[0][199] , \round_in[0][198] , \round_in[0][197] , 
        \round_in[0][196] , \round_in[0][195] , \round_in[0][194] , 
        \round_in[0][193] , \round_in[0][192] , \round_in[0][191] , 
        \round_in[0][190] , \round_in[0][189] , \round_in[0][188] , 
        \round_in[0][187] , \round_in[0][186] , \round_in[0][185] , 
        \round_in[0][184] , \round_in[0][183] , \round_in[0][182] , 
        \round_in[0][181] , \round_in[0][180] , \round_in[0][179] , 
        \round_in[0][178] , \round_in[0][177] , \round_in[0][176] , 
        \round_in[0][175] , \round_in[0][174] , \round_in[0][173] , 
        \round_in[0][172] , \round_in[0][171] , \round_in[0][170] , 
        \round_in[0][169] , \round_in[0][168] , \round_in[0][167] , 
        \round_in[0][166] , \round_in[0][165] , \round_in[0][164] , 
        \round_in[0][163] , \round_in[0][162] , \round_in[0][161] , 
        \round_in[0][160] , \round_in[0][159] , \round_in[0][158] , 
        \round_in[0][157] , \round_in[0][156] , \round_in[0][155] , 
        \round_in[0][154] , \round_in[0][153] , \round_in[0][152] , 
        \round_in[0][151] , \round_in[0][150] , \round_in[0][149] , 
        \round_in[0][148] , \round_in[0][147] , \round_in[0][146] , 
        \round_in[0][145] , \round_in[0][144] , \round_in[0][143] , 
        \round_in[0][142] , \round_in[0][141] , \round_in[0][140] , 
        \round_in[0][139] , \round_in[0][138] , \round_in[0][137] , 
        \round_in[0][136] , \round_in[0][135] , \round_in[0][134] , 
        \round_in[0][133] , \round_in[0][132] , \round_in[0][131] , 
        \round_in[0][130] , \round_in[0][129] , \round_in[0][128] , 
        \round_in[0][127] , \round_in[0][126] , \round_in[0][125] , 
        \round_in[0][124] , \round_in[0][123] , \round_in[0][122] , 
        \round_in[0][121] , \round_in[0][120] , \round_in[0][119] , 
        \round_in[0][118] , \round_in[0][117] , \round_in[0][116] , 
        \round_in[0][115] , \round_in[0][114] , \round_in[0][113] , 
        \round_in[0][112] , \round_in[0][111] , \round_in[0][110] , 
        \round_in[0][109] , \round_in[0][108] , \round_in[0][107] , 
        \round_in[0][106] , \round_in[0][105] , \round_in[0][104] , 
        \round_in[0][103] , \round_in[0][102] , \round_in[0][101] , 
        \round_in[0][100] , \round_in[0][99] , \round_in[0][98] , 
        \round_in[0][97] , \round_in[0][96] , \round_in[0][95] , 
        \round_in[0][94] , \round_in[0][93] , \round_in[0][92] , 
        \round_in[0][91] , \round_in[0][90] , \round_in[0][89] , 
        \round_in[0][88] , \round_in[0][87] , \round_in[0][86] , 
        \round_in[0][85] , \round_in[0][84] , \round_in[0][83] , 
        \round_in[0][82] , \round_in[0][81] , \round_in[0][80] , 
        \round_in[0][79] , \round_in[0][78] , \round_in[0][77] , 
        \round_in[0][76] , \round_in[0][75] , \round_in[0][74] , 
        \round_in[0][73] , \round_in[0][72] , \round_in[0][71] , 
        \round_in[0][70] , \round_in[0][69] , \round_in[0][68] , 
        \round_in[0][67] , \round_in[0][66] , \round_in[0][65] , 
        \round_in[0][64] , \round_in[0][63] , \round_in[0][62] , 
        \round_in[0][61] , \round_in[0][60] , \round_in[0][59] , 
        \round_in[0][58] , \round_in[0][57] , \round_in[0][56] , 
        \round_in[0][55] , \round_in[0][54] , \round_in[0][53] , 
        \round_in[0][52] , \round_in[0][51] , \round_in[0][50] , 
        \round_in[0][49] , \round_in[0][48] , \round_in[0][47] , 
        \round_in[0][46] , \round_in[0][45] , \round_in[0][44] , 
        \round_in[0][43] , \round_in[0][42] , \round_in[0][41] , 
        \round_in[0][40] , \round_in[0][39] , \round_in[0][38] , 
        \round_in[0][37] , \round_in[0][36] , \round_in[0][35] , 
        \round_in[0][34] , \round_in[0][33] , \round_in[0][32] , 
        \round_in[0][31] , \round_in[0][30] , \round_in[0][29] , 
        \round_in[0][28] , \round_in[0][27] , \round_in[0][26] , 
        \round_in[0][25] , \round_in[0][24] , \round_in[0][23] , 
        \round_in[0][22] , \round_in[0][21] , \round_in[0][20] , 
        \round_in[0][19] , \round_in[0][18] , \round_in[0][17] , 
        \round_in[0][16] , \round_in[0][15] , \round_in[0][14] , 
        \round_in[0][13] , \round_in[0][12] , \round_in[0][11] , 
        \round_in[0][10] , \round_in[0][9] , \round_in[0][8] , 
        \round_in[0][7] , \round_in[0][6] , \round_in[0][5] , \round_in[0][4] , 
        \round_in[0][3] , \round_in[0][2] , \round_in[0][1] , \round_in[0][0] }), .round_const({\RCONST[0].rconst_/N67 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, \RCONST[0].rconst_/N56 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[0].rconst_/N48 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \rc[2][0] , 1'b0, 1'b0, 1'b0, \RCONST[0].rconst_/N25 , 1'b0, 
        \RCONST[0].rconst_/N17 , \rc[3][15] }), .out({\round_in[1][1599] , 
        \round_in[1][1598] , \round_in[1][1597] , \round_in[1][1596] , 
        \round_in[1][1595] , \round_in[1][1594] , \round_in[1][1593] , 
        \round_in[1][1592] , \round_in[1][1591] , \round_in[1][1590] , 
        \round_in[1][1589] , \round_in[1][1588] , \round_in[1][1587] , 
        \round_in[1][1586] , \round_in[1][1585] , \round_in[1][1584] , 
        \round_in[1][1583] , \round_in[1][1582] , \round_in[1][1581] , 
        \round_in[1][1580] , \round_in[1][1579] , \round_in[1][1578] , 
        \round_in[1][1577] , \round_in[1][1576] , \round_in[1][1575] , 
        \round_in[1][1574] , \round_in[1][1573] , \round_in[1][1572] , 
        \round_in[1][1571] , \round_in[1][1570] , \round_in[1][1569] , 
        \round_in[1][1568] , \round_in[1][1567] , \round_in[1][1566] , 
        \round_in[1][1565] , \round_in[1][1564] , \round_in[1][1563] , 
        \round_in[1][1562] , \round_in[1][1561] , \round_in[1][1560] , 
        \round_in[1][1559] , \round_in[1][1558] , \round_in[1][1557] , 
        \round_in[1][1556] , \round_in[1][1555] , \round_in[1][1554] , 
        \round_in[1][1553] , \round_in[1][1552] , \round_in[1][1551] , 
        \round_in[1][1550] , \round_in[1][1549] , \round_in[1][1548] , 
        \round_in[1][1547] , \round_in[1][1546] , \round_in[1][1545] , 
        \round_in[1][1544] , \round_in[1][1543] , \round_in[1][1542] , 
        \round_in[1][1541] , \round_in[1][1540] , \round_in[1][1539] , 
        \round_in[1][1538] , \round_in[1][1537] , \round_in[1][1536] , 
        \round_in[1][1535] , \round_in[1][1534] , \round_in[1][1533] , 
        \round_in[1][1532] , \round_in[1][1531] , \round_in[1][1530] , 
        \round_in[1][1529] , \round_in[1][1528] , \round_in[1][1527] , 
        \round_in[1][1526] , \round_in[1][1525] , \round_in[1][1524] , 
        \round_in[1][1523] , \round_in[1][1522] , \round_in[1][1521] , 
        \round_in[1][1520] , \round_in[1][1519] , \round_in[1][1518] , 
        \round_in[1][1517] , \round_in[1][1516] , \round_in[1][1515] , 
        \round_in[1][1514] , \round_in[1][1513] , \round_in[1][1512] , 
        \round_in[1][1511] , \round_in[1][1510] , \round_in[1][1509] , 
        \round_in[1][1508] , \round_in[1][1507] , \round_in[1][1506] , 
        \round_in[1][1505] , \round_in[1][1504] , \round_in[1][1503] , 
        \round_in[1][1502] , \round_in[1][1501] , \round_in[1][1500] , 
        \round_in[1][1499] , \round_in[1][1498] , \round_in[1][1497] , 
        \round_in[1][1496] , \round_in[1][1495] , \round_in[1][1494] , 
        \round_in[1][1493] , \round_in[1][1492] , \round_in[1][1491] , 
        \round_in[1][1490] , \round_in[1][1489] , \round_in[1][1488] , 
        \round_in[1][1487] , \round_in[1][1486] , \round_in[1][1485] , 
        \round_in[1][1484] , \round_in[1][1483] , \round_in[1][1482] , 
        \round_in[1][1481] , \round_in[1][1480] , \round_in[1][1479] , 
        \round_in[1][1478] , \round_in[1][1477] , \round_in[1][1476] , 
        \round_in[1][1475] , \round_in[1][1474] , \round_in[1][1473] , 
        \round_in[1][1472] , \round_in[1][1471] , \round_in[1][1470] , 
        \round_in[1][1469] , \round_in[1][1468] , \round_in[1][1467] , 
        \round_in[1][1466] , \round_in[1][1465] , \round_in[1][1464] , 
        \round_in[1][1463] , \round_in[1][1462] , \round_in[1][1461] , 
        \round_in[1][1460] , \round_in[1][1459] , \round_in[1][1458] , 
        \round_in[1][1457] , \round_in[1][1456] , \round_in[1][1455] , 
        \round_in[1][1454] , \round_in[1][1453] , \round_in[1][1452] , 
        \round_in[1][1451] , \round_in[1][1450] , \round_in[1][1449] , 
        \round_in[1][1448] , \round_in[1][1447] , \round_in[1][1446] , 
        \round_in[1][1445] , \round_in[1][1444] , \round_in[1][1443] , 
        \round_in[1][1442] , \round_in[1][1441] , \round_in[1][1440] , 
        \round_in[1][1439] , \round_in[1][1438] , \round_in[1][1437] , 
        \round_in[1][1436] , \round_in[1][1435] , \round_in[1][1434] , 
        \round_in[1][1433] , \round_in[1][1432] , \round_in[1][1431] , 
        \round_in[1][1430] , \round_in[1][1429] , \round_in[1][1428] , 
        \round_in[1][1427] , \round_in[1][1426] , \round_in[1][1425] , 
        \round_in[1][1424] , \round_in[1][1423] , \round_in[1][1422] , 
        \round_in[1][1421] , \round_in[1][1420] , \round_in[1][1419] , 
        \round_in[1][1418] , \round_in[1][1417] , \round_in[1][1416] , 
        \round_in[1][1415] , \round_in[1][1414] , \round_in[1][1413] , 
        \round_in[1][1412] , \round_in[1][1411] , \round_in[1][1410] , 
        \round_in[1][1409] , \round_in[1][1408] , \round_in[1][1407] , 
        \round_in[1][1406] , \round_in[1][1405] , \round_in[1][1404] , 
        \round_in[1][1403] , \round_in[1][1402] , \round_in[1][1401] , 
        \round_in[1][1400] , \round_in[1][1399] , \round_in[1][1398] , 
        \round_in[1][1397] , \round_in[1][1396] , \round_in[1][1395] , 
        \round_in[1][1394] , \round_in[1][1393] , \round_in[1][1392] , 
        \round_in[1][1391] , \round_in[1][1390] , \round_in[1][1389] , 
        \round_in[1][1388] , \round_in[1][1387] , \round_in[1][1386] , 
        \round_in[1][1385] , \round_in[1][1384] , \round_in[1][1383] , 
        \round_in[1][1382] , \round_in[1][1381] , \round_in[1][1380] , 
        \round_in[1][1379] , \round_in[1][1378] , \round_in[1][1377] , 
        \round_in[1][1376] , \round_in[1][1375] , \round_in[1][1374] , 
        \round_in[1][1373] , \round_in[1][1372] , \round_in[1][1371] , 
        \round_in[1][1370] , \round_in[1][1369] , \round_in[1][1368] , 
        \round_in[1][1367] , \round_in[1][1366] , \round_in[1][1365] , 
        \round_in[1][1364] , \round_in[1][1363] , \round_in[1][1362] , 
        \round_in[1][1361] , \round_in[1][1360] , \round_in[1][1359] , 
        \round_in[1][1358] , \round_in[1][1357] , \round_in[1][1356] , 
        \round_in[1][1355] , \round_in[1][1354] , \round_in[1][1353] , 
        \round_in[1][1352] , \round_in[1][1351] , \round_in[1][1350] , 
        \round_in[1][1349] , \round_in[1][1348] , \round_in[1][1347] , 
        \round_in[1][1346] , \round_in[1][1345] , \round_in[1][1344] , 
        \round_in[1][1343] , \round_in[1][1342] , \round_in[1][1341] , 
        \round_in[1][1340] , \round_in[1][1339] , \round_in[1][1338] , 
        \round_in[1][1337] , \round_in[1][1336] , \round_in[1][1335] , 
        \round_in[1][1334] , \round_in[1][1333] , \round_in[1][1332] , 
        \round_in[1][1331] , \round_in[1][1330] , \round_in[1][1329] , 
        \round_in[1][1328] , \round_in[1][1327] , \round_in[1][1326] , 
        \round_in[1][1325] , \round_in[1][1324] , \round_in[1][1323] , 
        \round_in[1][1322] , \round_in[1][1321] , \round_in[1][1320] , 
        \round_in[1][1319] , \round_in[1][1318] , \round_in[1][1317] , 
        \round_in[1][1316] , \round_in[1][1315] , \round_in[1][1314] , 
        \round_in[1][1313] , \round_in[1][1312] , \round_in[1][1311] , 
        \round_in[1][1310] , \round_in[1][1309] , \round_in[1][1308] , 
        \round_in[1][1307] , \round_in[1][1306] , \round_in[1][1305] , 
        \round_in[1][1304] , \round_in[1][1303] , \round_in[1][1302] , 
        \round_in[1][1301] , \round_in[1][1300] , \round_in[1][1299] , 
        \round_in[1][1298] , \round_in[1][1297] , \round_in[1][1296] , 
        \round_in[1][1295] , \round_in[1][1294] , \round_in[1][1293] , 
        \round_in[1][1292] , \round_in[1][1291] , \round_in[1][1290] , 
        \round_in[1][1289] , \round_in[1][1288] , \round_in[1][1287] , 
        \round_in[1][1286] , \round_in[1][1285] , \round_in[1][1284] , 
        \round_in[1][1283] , \round_in[1][1282] , \round_in[1][1281] , 
        \round_in[1][1280] , \round_in[1][1279] , \round_in[1][1278] , 
        \round_in[1][1277] , \round_in[1][1276] , \round_in[1][1275] , 
        \round_in[1][1274] , \round_in[1][1273] , \round_in[1][1272] , 
        \round_in[1][1271] , \round_in[1][1270] , \round_in[1][1269] , 
        \round_in[1][1268] , \round_in[1][1267] , \round_in[1][1266] , 
        \round_in[1][1265] , \round_in[1][1264] , \round_in[1][1263] , 
        \round_in[1][1262] , \round_in[1][1261] , \round_in[1][1260] , 
        \round_in[1][1259] , \round_in[1][1258] , \round_in[1][1257] , 
        \round_in[1][1256] , \round_in[1][1255] , \round_in[1][1254] , 
        \round_in[1][1253] , \round_in[1][1252] , \round_in[1][1251] , 
        \round_in[1][1250] , \round_in[1][1249] , \round_in[1][1248] , 
        \round_in[1][1247] , \round_in[1][1246] , \round_in[1][1245] , 
        \round_in[1][1244] , \round_in[1][1243] , \round_in[1][1242] , 
        \round_in[1][1241] , \round_in[1][1240] , \round_in[1][1239] , 
        \round_in[1][1238] , \round_in[1][1237] , \round_in[1][1236] , 
        \round_in[1][1235] , \round_in[1][1234] , \round_in[1][1233] , 
        \round_in[1][1232] , \round_in[1][1231] , \round_in[1][1230] , 
        \round_in[1][1229] , \round_in[1][1228] , \round_in[1][1227] , 
        \round_in[1][1226] , \round_in[1][1225] , \round_in[1][1224] , 
        \round_in[1][1223] , \round_in[1][1222] , \round_in[1][1221] , 
        \round_in[1][1220] , \round_in[1][1219] , \round_in[1][1218] , 
        \round_in[1][1217] , \round_in[1][1216] , \round_in[1][1215] , 
        \round_in[1][1214] , \round_in[1][1213] , \round_in[1][1212] , 
        \round_in[1][1211] , \round_in[1][1210] , \round_in[1][1209] , 
        \round_in[1][1208] , \round_in[1][1207] , \round_in[1][1206] , 
        \round_in[1][1205] , \round_in[1][1204] , \round_in[1][1203] , 
        \round_in[1][1202] , \round_in[1][1201] , \round_in[1][1200] , 
        \round_in[1][1199] , \round_in[1][1198] , \round_in[1][1197] , 
        \round_in[1][1196] , \round_in[1][1195] , \round_in[1][1194] , 
        \round_in[1][1193] , \round_in[1][1192] , \round_in[1][1191] , 
        \round_in[1][1190] , \round_in[1][1189] , \round_in[1][1188] , 
        \round_in[1][1187] , \round_in[1][1186] , \round_in[1][1185] , 
        \round_in[1][1184] , \round_in[1][1183] , \round_in[1][1182] , 
        \round_in[1][1181] , \round_in[1][1180] , \round_in[1][1179] , 
        \round_in[1][1178] , \round_in[1][1177] , \round_in[1][1176] , 
        \round_in[1][1175] , \round_in[1][1174] , \round_in[1][1173] , 
        \round_in[1][1172] , \round_in[1][1171] , \round_in[1][1170] , 
        \round_in[1][1169] , \round_in[1][1168] , \round_in[1][1167] , 
        \round_in[1][1166] , \round_in[1][1165] , \round_in[1][1164] , 
        \round_in[1][1163] , \round_in[1][1162] , \round_in[1][1161] , 
        \round_in[1][1160] , \round_in[1][1159] , \round_in[1][1158] , 
        \round_in[1][1157] , \round_in[1][1156] , \round_in[1][1155] , 
        \round_in[1][1154] , \round_in[1][1153] , \round_in[1][1152] , 
        \round_in[1][1151] , \round_in[1][1150] , \round_in[1][1149] , 
        \round_in[1][1148] , \round_in[1][1147] , \round_in[1][1146] , 
        \round_in[1][1145] , \round_in[1][1144] , \round_in[1][1143] , 
        \round_in[1][1142] , \round_in[1][1141] , \round_in[1][1140] , 
        \round_in[1][1139] , \round_in[1][1138] , \round_in[1][1137] , 
        \round_in[1][1136] , \round_in[1][1135] , \round_in[1][1134] , 
        \round_in[1][1133] , \round_in[1][1132] , \round_in[1][1131] , 
        \round_in[1][1130] , \round_in[1][1129] , \round_in[1][1128] , 
        \round_in[1][1127] , \round_in[1][1126] , \round_in[1][1125] , 
        \round_in[1][1124] , \round_in[1][1123] , \round_in[1][1122] , 
        \round_in[1][1121] , \round_in[1][1120] , \round_in[1][1119] , 
        \round_in[1][1118] , \round_in[1][1117] , \round_in[1][1116] , 
        \round_in[1][1115] , \round_in[1][1114] , \round_in[1][1113] , 
        \round_in[1][1112] , \round_in[1][1111] , \round_in[1][1110] , 
        \round_in[1][1109] , \round_in[1][1108] , \round_in[1][1107] , 
        \round_in[1][1106] , \round_in[1][1105] , \round_in[1][1104] , 
        \round_in[1][1103] , \round_in[1][1102] , \round_in[1][1101] , 
        \round_in[1][1100] , \round_in[1][1099] , \round_in[1][1098] , 
        \round_in[1][1097] , \round_in[1][1096] , \round_in[1][1095] , 
        \round_in[1][1094] , \round_in[1][1093] , \round_in[1][1092] , 
        \round_in[1][1091] , \round_in[1][1090] , \round_in[1][1089] , 
        \round_in[1][1088] , \round_in[1][1087] , \round_in[1][1086] , 
        \round_in[1][1085] , \round_in[1][1084] , \round_in[1][1083] , 
        \round_in[1][1082] , \round_in[1][1081] , \round_in[1][1080] , 
        \round_in[1][1079] , \round_in[1][1078] , \round_in[1][1077] , 
        \round_in[1][1076] , \round_in[1][1075] , \round_in[1][1074] , 
        \round_in[1][1073] , \round_in[1][1072] , \round_in[1][1071] , 
        \round_in[1][1070] , \round_in[1][1069] , \round_in[1][1068] , 
        \round_in[1][1067] , \round_in[1][1066] , \round_in[1][1065] , 
        \round_in[1][1064] , \round_in[1][1063] , \round_in[1][1062] , 
        \round_in[1][1061] , \round_in[1][1060] , \round_in[1][1059] , 
        \round_in[1][1058] , \round_in[1][1057] , \round_in[1][1056] , 
        \round_in[1][1055] , \round_in[1][1054] , \round_in[1][1053] , 
        \round_in[1][1052] , \round_in[1][1051] , \round_in[1][1050] , 
        \round_in[1][1049] , \round_in[1][1048] , \round_in[1][1047] , 
        \round_in[1][1046] , \round_in[1][1045] , \round_in[1][1044] , 
        \round_in[1][1043] , \round_in[1][1042] , \round_in[1][1041] , 
        \round_in[1][1040] , \round_in[1][1039] , \round_in[1][1038] , 
        \round_in[1][1037] , \round_in[1][1036] , \round_in[1][1035] , 
        \round_in[1][1034] , \round_in[1][1033] , \round_in[1][1032] , 
        \round_in[1][1031] , \round_in[1][1030] , \round_in[1][1029] , 
        \round_in[1][1028] , \round_in[1][1027] , \round_in[1][1026] , 
        \round_in[1][1025] , \round_in[1][1024] , \round_in[1][1023] , 
        \round_in[1][1022] , \round_in[1][1021] , \round_in[1][1020] , 
        \round_in[1][1019] , \round_in[1][1018] , \round_in[1][1017] , 
        \round_in[1][1016] , \round_in[1][1015] , \round_in[1][1014] , 
        \round_in[1][1013] , \round_in[1][1012] , \round_in[1][1011] , 
        \round_in[1][1010] , \round_in[1][1009] , \round_in[1][1008] , 
        \round_in[1][1007] , \round_in[1][1006] , \round_in[1][1005] , 
        \round_in[1][1004] , \round_in[1][1003] , \round_in[1][1002] , 
        \round_in[1][1001] , \round_in[1][1000] , \round_in[1][999] , 
        \round_in[1][998] , \round_in[1][997] , \round_in[1][996] , 
        \round_in[1][995] , \round_in[1][994] , \round_in[1][993] , 
        \round_in[1][992] , \round_in[1][991] , \round_in[1][990] , 
        \round_in[1][989] , \round_in[1][988] , \round_in[1][987] , 
        \round_in[1][986] , \round_in[1][985] , \round_in[1][984] , 
        \round_in[1][983] , \round_in[1][982] , \round_in[1][981] , 
        \round_in[1][980] , \round_in[1][979] , \round_in[1][978] , 
        \round_in[1][977] , \round_in[1][976] , \round_in[1][975] , 
        \round_in[1][974] , \round_in[1][973] , \round_in[1][972] , 
        \round_in[1][971] , \round_in[1][970] , \round_in[1][969] , 
        \round_in[1][968] , \round_in[1][967] , \round_in[1][966] , 
        \round_in[1][965] , \round_in[1][964] , \round_in[1][963] , 
        \round_in[1][962] , \round_in[1][961] , \round_in[1][960] , 
        \round_in[1][959] , \round_in[1][958] , \round_in[1][957] , 
        \round_in[1][956] , \round_in[1][955] , \round_in[1][954] , 
        \round_in[1][953] , \round_in[1][952] , \round_in[1][951] , 
        \round_in[1][950] , \round_in[1][949] , \round_in[1][948] , 
        \round_in[1][947] , \round_in[1][946] , \round_in[1][945] , 
        \round_in[1][944] , \round_in[1][943] , \round_in[1][942] , 
        \round_in[1][941] , \round_in[1][940] , \round_in[1][939] , 
        \round_in[1][938] , \round_in[1][937] , \round_in[1][936] , 
        \round_in[1][935] , \round_in[1][934] , \round_in[1][933] , 
        \round_in[1][932] , \round_in[1][931] , \round_in[1][930] , 
        \round_in[1][929] , \round_in[1][928] , \round_in[1][927] , 
        \round_in[1][926] , \round_in[1][925] , \round_in[1][924] , 
        \round_in[1][923] , \round_in[1][922] , \round_in[1][921] , 
        \round_in[1][920] , \round_in[1][919] , \round_in[1][918] , 
        \round_in[1][917] , \round_in[1][916] , \round_in[1][915] , 
        \round_in[1][914] , \round_in[1][913] , \round_in[1][912] , 
        \round_in[1][911] , \round_in[1][910] , \round_in[1][909] , 
        \round_in[1][908] , \round_in[1][907] , \round_in[1][906] , 
        \round_in[1][905] , \round_in[1][904] , \round_in[1][903] , 
        \round_in[1][902] , \round_in[1][901] , \round_in[1][900] , 
        \round_in[1][899] , \round_in[1][898] , \round_in[1][897] , 
        \round_in[1][896] , \round_in[1][895] , \round_in[1][894] , 
        \round_in[1][893] , \round_in[1][892] , \round_in[1][891] , 
        \round_in[1][890] , \round_in[1][889] , \round_in[1][888] , 
        \round_in[1][887] , \round_in[1][886] , \round_in[1][885] , 
        \round_in[1][884] , \round_in[1][883] , \round_in[1][882] , 
        \round_in[1][881] , \round_in[1][880] , \round_in[1][879] , 
        \round_in[1][878] , \round_in[1][877] , \round_in[1][876] , 
        \round_in[1][875] , \round_in[1][874] , \round_in[1][873] , 
        \round_in[1][872] , \round_in[1][871] , \round_in[1][870] , 
        \round_in[1][869] , \round_in[1][868] , \round_in[1][867] , 
        \round_in[1][866] , \round_in[1][865] , \round_in[1][864] , 
        \round_in[1][863] , \round_in[1][862] , \round_in[1][861] , 
        \round_in[1][860] , \round_in[1][859] , \round_in[1][858] , 
        \round_in[1][857] , \round_in[1][856] , \round_in[1][855] , 
        \round_in[1][854] , \round_in[1][853] , \round_in[1][852] , 
        \round_in[1][851] , \round_in[1][850] , \round_in[1][849] , 
        \round_in[1][848] , \round_in[1][847] , \round_in[1][846] , 
        \round_in[1][845] , \round_in[1][844] , \round_in[1][843] , 
        \round_in[1][842] , \round_in[1][841] , \round_in[1][840] , 
        \round_in[1][839] , \round_in[1][838] , \round_in[1][837] , 
        \round_in[1][836] , \round_in[1][835] , \round_in[1][834] , 
        \round_in[1][833] , \round_in[1][832] , \round_in[1][831] , 
        \round_in[1][830] , \round_in[1][829] , \round_in[1][828] , 
        \round_in[1][827] , \round_in[1][826] , \round_in[1][825] , 
        \round_in[1][824] , \round_in[1][823] , \round_in[1][822] , 
        \round_in[1][821] , \round_in[1][820] , \round_in[1][819] , 
        \round_in[1][818] , \round_in[1][817] , \round_in[1][816] , 
        \round_in[1][815] , \round_in[1][814] , \round_in[1][813] , 
        \round_in[1][812] , \round_in[1][811] , \round_in[1][810] , 
        \round_in[1][809] , \round_in[1][808] , \round_in[1][807] , 
        \round_in[1][806] , \round_in[1][805] , \round_in[1][804] , 
        \round_in[1][803] , \round_in[1][802] , \round_in[1][801] , 
        \round_in[1][800] , \round_in[1][799] , \round_in[1][798] , 
        \round_in[1][797] , \round_in[1][796] , \round_in[1][795] , 
        \round_in[1][794] , \round_in[1][793] , \round_in[1][792] , 
        \round_in[1][791] , \round_in[1][790] , \round_in[1][789] , 
        \round_in[1][788] , \round_in[1][787] , \round_in[1][786] , 
        \round_in[1][785] , \round_in[1][784] , \round_in[1][783] , 
        \round_in[1][782] , \round_in[1][781] , \round_in[1][780] , 
        \round_in[1][779] , \round_in[1][778] , \round_in[1][777] , 
        \round_in[1][776] , \round_in[1][775] , \round_in[1][774] , 
        \round_in[1][773] , \round_in[1][772] , \round_in[1][771] , 
        \round_in[1][770] , \round_in[1][769] , \round_in[1][768] , 
        \round_in[1][767] , \round_in[1][766] , \round_in[1][765] , 
        \round_in[1][764] , \round_in[1][763] , \round_in[1][762] , 
        \round_in[1][761] , \round_in[1][760] , \round_in[1][759] , 
        \round_in[1][758] , \round_in[1][757] , \round_in[1][756] , 
        \round_in[1][755] , \round_in[1][754] , \round_in[1][753] , 
        \round_in[1][752] , \round_in[1][751] , \round_in[1][750] , 
        \round_in[1][749] , \round_in[1][748] , \round_in[1][747] , 
        \round_in[1][746] , \round_in[1][745] , \round_in[1][744] , 
        \round_in[1][743] , \round_in[1][742] , \round_in[1][741] , 
        \round_in[1][740] , \round_in[1][739] , \round_in[1][738] , 
        \round_in[1][737] , \round_in[1][736] , \round_in[1][735] , 
        \round_in[1][734] , \round_in[1][733] , \round_in[1][732] , 
        \round_in[1][731] , \round_in[1][730] , \round_in[1][729] , 
        \round_in[1][728] , \round_in[1][727] , \round_in[1][726] , 
        \round_in[1][725] , \round_in[1][724] , \round_in[1][723] , 
        \round_in[1][722] , \round_in[1][721] , \round_in[1][720] , 
        \round_in[1][719] , \round_in[1][718] , \round_in[1][717] , 
        \round_in[1][716] , \round_in[1][715] , \round_in[1][714] , 
        \round_in[1][713] , \round_in[1][712] , \round_in[1][711] , 
        \round_in[1][710] , \round_in[1][709] , \round_in[1][708] , 
        \round_in[1][707] , \round_in[1][706] , \round_in[1][705] , 
        \round_in[1][704] , \round_in[1][703] , \round_in[1][702] , 
        \round_in[1][701] , \round_in[1][700] , \round_in[1][699] , 
        \round_in[1][698] , \round_in[1][697] , \round_in[1][696] , 
        \round_in[1][695] , \round_in[1][694] , \round_in[1][693] , 
        \round_in[1][692] , \round_in[1][691] , \round_in[1][690] , 
        \round_in[1][689] , \round_in[1][688] , \round_in[1][687] , 
        \round_in[1][686] , \round_in[1][685] , \round_in[1][684] , 
        \round_in[1][683] , \round_in[1][682] , \round_in[1][681] , 
        \round_in[1][680] , \round_in[1][679] , \round_in[1][678] , 
        \round_in[1][677] , \round_in[1][676] , \round_in[1][675] , 
        \round_in[1][674] , \round_in[1][673] , \round_in[1][672] , 
        \round_in[1][671] , \round_in[1][670] , \round_in[1][669] , 
        \round_in[1][668] , \round_in[1][667] , \round_in[1][666] , 
        \round_in[1][665] , \round_in[1][664] , \round_in[1][663] , 
        \round_in[1][662] , \round_in[1][661] , \round_in[1][660] , 
        \round_in[1][659] , \round_in[1][658] , \round_in[1][657] , 
        \round_in[1][656] , \round_in[1][655] , \round_in[1][654] , 
        \round_in[1][653] , \round_in[1][652] , \round_in[1][651] , 
        \round_in[1][650] , \round_in[1][649] , \round_in[1][648] , 
        \round_in[1][647] , \round_in[1][646] , \round_in[1][645] , 
        \round_in[1][644] , \round_in[1][643] , \round_in[1][642] , 
        \round_in[1][641] , \round_in[1][640] , \round_in[1][639] , 
        \round_in[1][638] , \round_in[1][637] , \round_in[1][636] , 
        \round_in[1][635] , \round_in[1][634] , \round_in[1][633] , 
        \round_in[1][632] , \round_in[1][631] , \round_in[1][630] , 
        \round_in[1][629] , \round_in[1][628] , \round_in[1][627] , 
        \round_in[1][626] , \round_in[1][625] , \round_in[1][624] , 
        \round_in[1][623] , \round_in[1][622] , \round_in[1][621] , 
        \round_in[1][620] , \round_in[1][619] , \round_in[1][618] , 
        \round_in[1][617] , \round_in[1][616] , \round_in[1][615] , 
        \round_in[1][614] , \round_in[1][613] , \round_in[1][612] , 
        \round_in[1][611] , \round_in[1][610] , \round_in[1][609] , 
        \round_in[1][608] , \round_in[1][607] , \round_in[1][606] , 
        \round_in[1][605] , \round_in[1][604] , \round_in[1][603] , 
        \round_in[1][602] , \round_in[1][601] , \round_in[1][600] , 
        \round_in[1][599] , \round_in[1][598] , \round_in[1][597] , 
        \round_in[1][596] , \round_in[1][595] , \round_in[1][594] , 
        \round_in[1][593] , \round_in[1][592] , \round_in[1][591] , 
        \round_in[1][590] , \round_in[1][589] , \round_in[1][588] , 
        \round_in[1][587] , \round_in[1][586] , \round_in[1][585] , 
        \round_in[1][584] , \round_in[1][583] , \round_in[1][582] , 
        \round_in[1][581] , \round_in[1][580] , \round_in[1][579] , 
        \round_in[1][578] , \round_in[1][577] , \round_in[1][576] , 
        \round_in[1][575] , \round_in[1][574] , \round_in[1][573] , 
        \round_in[1][572] , \round_in[1][571] , \round_in[1][570] , 
        \round_in[1][569] , \round_in[1][568] , \round_in[1][567] , 
        \round_in[1][566] , \round_in[1][565] , \round_in[1][564] , 
        \round_in[1][563] , \round_in[1][562] , \round_in[1][561] , 
        \round_in[1][560] , \round_in[1][559] , \round_in[1][558] , 
        \round_in[1][557] , \round_in[1][556] , \round_in[1][555] , 
        \round_in[1][554] , \round_in[1][553] , \round_in[1][552] , 
        \round_in[1][551] , \round_in[1][550] , \round_in[1][549] , 
        \round_in[1][548] , \round_in[1][547] , \round_in[1][546] , 
        \round_in[1][545] , \round_in[1][544] , \round_in[1][543] , 
        \round_in[1][542] , \round_in[1][541] , \round_in[1][540] , 
        \round_in[1][539] , \round_in[1][538] , \round_in[1][537] , 
        \round_in[1][536] , \round_in[1][535] , \round_in[1][534] , 
        \round_in[1][533] , \round_in[1][532] , \round_in[1][531] , 
        \round_in[1][530] , \round_in[1][529] , \round_in[1][528] , 
        \round_in[1][527] , \round_in[1][526] , \round_in[1][525] , 
        \round_in[1][524] , \round_in[1][523] , \round_in[1][522] , 
        \round_in[1][521] , \round_in[1][520] , \round_in[1][519] , 
        \round_in[1][518] , \round_in[1][517] , \round_in[1][516] , 
        \round_in[1][515] , \round_in[1][514] , \round_in[1][513] , 
        \round_in[1][512] , \round_in[1][511] , \round_in[1][510] , 
        \round_in[1][509] , \round_in[1][508] , \round_in[1][507] , 
        \round_in[1][506] , \round_in[1][505] , \round_in[1][504] , 
        \round_in[1][503] , \round_in[1][502] , \round_in[1][501] , 
        \round_in[1][500] , \round_in[1][499] , \round_in[1][498] , 
        \round_in[1][497] , \round_in[1][496] , \round_in[1][495] , 
        \round_in[1][494] , \round_in[1][493] , \round_in[1][492] , 
        \round_in[1][491] , \round_in[1][490] , \round_in[1][489] , 
        \round_in[1][488] , \round_in[1][487] , \round_in[1][486] , 
        \round_in[1][485] , \round_in[1][484] , \round_in[1][483] , 
        \round_in[1][482] , \round_in[1][481] , \round_in[1][480] , 
        \round_in[1][479] , \round_in[1][478] , \round_in[1][477] , 
        \round_in[1][476] , \round_in[1][475] , \round_in[1][474] , 
        \round_in[1][473] , \round_in[1][472] , \round_in[1][471] , 
        \round_in[1][470] , \round_in[1][469] , \round_in[1][468] , 
        \round_in[1][467] , \round_in[1][466] , \round_in[1][465] , 
        \round_in[1][464] , \round_in[1][463] , \round_in[1][462] , 
        \round_in[1][461] , \round_in[1][460] , \round_in[1][459] , 
        \round_in[1][458] , \round_in[1][457] , \round_in[1][456] , 
        \round_in[1][455] , \round_in[1][454] , \round_in[1][453] , 
        \round_in[1][452] , \round_in[1][451] , \round_in[1][450] , 
        \round_in[1][449] , \round_in[1][448] , \round_in[1][447] , 
        \round_in[1][446] , \round_in[1][445] , \round_in[1][444] , 
        \round_in[1][443] , \round_in[1][442] , \round_in[1][441] , 
        \round_in[1][440] , \round_in[1][439] , \round_in[1][438] , 
        \round_in[1][437] , \round_in[1][436] , \round_in[1][435] , 
        \round_in[1][434] , \round_in[1][433] , \round_in[1][432] , 
        \round_in[1][431] , \round_in[1][430] , \round_in[1][429] , 
        \round_in[1][428] , \round_in[1][427] , \round_in[1][426] , 
        \round_in[1][425] , \round_in[1][424] , \round_in[1][423] , 
        \round_in[1][422] , \round_in[1][421] , \round_in[1][420] , 
        \round_in[1][419] , \round_in[1][418] , \round_in[1][417] , 
        \round_in[1][416] , \round_in[1][415] , \round_in[1][414] , 
        \round_in[1][413] , \round_in[1][412] , \round_in[1][411] , 
        \round_in[1][410] , \round_in[1][409] , \round_in[1][408] , 
        \round_in[1][407] , \round_in[1][406] , \round_in[1][405] , 
        \round_in[1][404] , \round_in[1][403] , \round_in[1][402] , 
        \round_in[1][401] , \round_in[1][400] , \round_in[1][399] , 
        \round_in[1][398] , \round_in[1][397] , \round_in[1][396] , 
        \round_in[1][395] , \round_in[1][394] , \round_in[1][393] , 
        \round_in[1][392] , \round_in[1][391] , \round_in[1][390] , 
        \round_in[1][389] , \round_in[1][388] , \round_in[1][387] , 
        \round_in[1][386] , \round_in[1][385] , \round_in[1][384] , 
        \round_in[1][383] , \round_in[1][382] , \round_in[1][381] , 
        \round_in[1][380] , \round_in[1][379] , \round_in[1][378] , 
        \round_in[1][377] , \round_in[1][376] , \round_in[1][375] , 
        \round_in[1][374] , \round_in[1][373] , \round_in[1][372] , 
        \round_in[1][371] , \round_in[1][370] , \round_in[1][369] , 
        \round_in[1][368] , \round_in[1][367] , \round_in[1][366] , 
        \round_in[1][365] , \round_in[1][364] , \round_in[1][363] , 
        \round_in[1][362] , \round_in[1][361] , \round_in[1][360] , 
        \round_in[1][359] , \round_in[1][358] , \round_in[1][357] , 
        \round_in[1][356] , \round_in[1][355] , \round_in[1][354] , 
        \round_in[1][353] , \round_in[1][352] , \round_in[1][351] , 
        \round_in[1][350] , \round_in[1][349] , \round_in[1][348] , 
        \round_in[1][347] , \round_in[1][346] , \round_in[1][345] , 
        \round_in[1][344] , \round_in[1][343] , \round_in[1][342] , 
        \round_in[1][341] , \round_in[1][340] , \round_in[1][339] , 
        \round_in[1][338] , \round_in[1][337] , \round_in[1][336] , 
        \round_in[1][335] , \round_in[1][334] , \round_in[1][333] , 
        \round_in[1][332] , \round_in[1][331] , \round_in[1][330] , 
        \round_in[1][329] , \round_in[1][328] , \round_in[1][327] , 
        \round_in[1][326] , \round_in[1][325] , \round_in[1][324] , 
        \round_in[1][323] , \round_in[1][322] , \round_in[1][321] , 
        \round_in[1][320] , \round_in[1][319] , \round_in[1][318] , 
        \round_in[1][317] , \round_in[1][316] , \round_in[1][315] , 
        \round_in[1][314] , \round_in[1][313] , \round_in[1][312] , 
        \round_in[1][311] , \round_in[1][310] , \round_in[1][309] , 
        \round_in[1][308] , \round_in[1][307] , \round_in[1][306] , 
        \round_in[1][305] , \round_in[1][304] , \round_in[1][303] , 
        \round_in[1][302] , \round_in[1][301] , \round_in[1][300] , 
        \round_in[1][299] , \round_in[1][298] , \round_in[1][297] , 
        \round_in[1][296] , \round_in[1][295] , \round_in[1][294] , 
        \round_in[1][293] , \round_in[1][292] , \round_in[1][291] , 
        \round_in[1][290] , \round_in[1][289] , \round_in[1][288] , 
        \round_in[1][287] , \round_in[1][286] , \round_in[1][285] , 
        \round_in[1][284] , \round_in[1][283] , \round_in[1][282] , 
        \round_in[1][281] , \round_in[1][280] , \round_in[1][279] , 
        \round_in[1][278] , \round_in[1][277] , \round_in[1][276] , 
        \round_in[1][275] , \round_in[1][274] , \round_in[1][273] , 
        \round_in[1][272] , \round_in[1][271] , \round_in[1][270] , 
        \round_in[1][269] , \round_in[1][268] , \round_in[1][267] , 
        \round_in[1][266] , \round_in[1][265] , \round_in[1][264] , 
        \round_in[1][263] , \round_in[1][262] , \round_in[1][261] , 
        \round_in[1][260] , \round_in[1][259] , \round_in[1][258] , 
        \round_in[1][257] , \round_in[1][256] , \round_in[1][255] , 
        \round_in[1][254] , \round_in[1][253] , \round_in[1][252] , 
        \round_in[1][251] , \round_in[1][250] , \round_in[1][249] , 
        \round_in[1][248] , \round_in[1][247] , \round_in[1][246] , 
        \round_in[1][245] , \round_in[1][244] , \round_in[1][243] , 
        \round_in[1][242] , \round_in[1][241] , \round_in[1][240] , 
        \round_in[1][239] , \round_in[1][238] , \round_in[1][237] , 
        \round_in[1][236] , \round_in[1][235] , \round_in[1][234] , 
        \round_in[1][233] , \round_in[1][232] , \round_in[1][231] , 
        \round_in[1][230] , \round_in[1][229] , \round_in[1][228] , 
        \round_in[1][227] , \round_in[1][226] , \round_in[1][225] , 
        \round_in[1][224] , \round_in[1][223] , \round_in[1][222] , 
        \round_in[1][221] , \round_in[1][220] , \round_in[1][219] , 
        \round_in[1][218] , \round_in[1][217] , \round_in[1][216] , 
        \round_in[1][215] , \round_in[1][214] , \round_in[1][213] , 
        \round_in[1][212] , \round_in[1][211] , \round_in[1][210] , 
        \round_in[1][209] , \round_in[1][208] , \round_in[1][207] , 
        \round_in[1][206] , \round_in[1][205] , \round_in[1][204] , 
        \round_in[1][203] , \round_in[1][202] , \round_in[1][201] , 
        \round_in[1][200] , \round_in[1][199] , \round_in[1][198] , 
        \round_in[1][197] , \round_in[1][196] , \round_in[1][195] , 
        \round_in[1][194] , \round_in[1][193] , \round_in[1][192] , 
        \round_in[1][191] , \round_in[1][190] , \round_in[1][189] , 
        \round_in[1][188] , \round_in[1][187] , \round_in[1][186] , 
        \round_in[1][185] , \round_in[1][184] , \round_in[1][183] , 
        \round_in[1][182] , \round_in[1][181] , \round_in[1][180] , 
        \round_in[1][179] , \round_in[1][178] , \round_in[1][177] , 
        \round_in[1][176] , \round_in[1][175] , \round_in[1][174] , 
        \round_in[1][173] , \round_in[1][172] , \round_in[1][171] , 
        \round_in[1][170] , \round_in[1][169] , \round_in[1][168] , 
        \round_in[1][167] , \round_in[1][166] , \round_in[1][165] , 
        \round_in[1][164] , \round_in[1][163] , \round_in[1][162] , 
        \round_in[1][161] , \round_in[1][160] , \round_in[1][159] , 
        \round_in[1][158] , \round_in[1][157] , \round_in[1][156] , 
        \round_in[1][155] , \round_in[1][154] , \round_in[1][153] , 
        \round_in[1][152] , \round_in[1][151] , \round_in[1][150] , 
        \round_in[1][149] , \round_in[1][148] , \round_in[1][147] , 
        \round_in[1][146] , \round_in[1][145] , \round_in[1][144] , 
        \round_in[1][143] , \round_in[1][142] , \round_in[1][141] , 
        \round_in[1][140] , \round_in[1][139] , \round_in[1][138] , 
        \round_in[1][137] , \round_in[1][136] , \round_in[1][135] , 
        \round_in[1][134] , \round_in[1][133] , \round_in[1][132] , 
        \round_in[1][131] , \round_in[1][130] , \round_in[1][129] , 
        \round_in[1][128] , \round_in[1][127] , \round_in[1][126] , 
        \round_in[1][125] , \round_in[1][124] , \round_in[1][123] , 
        \round_in[1][122] , \round_in[1][121] , \round_in[1][120] , 
        \round_in[1][119] , \round_in[1][118] , \round_in[1][117] , 
        \round_in[1][116] , \round_in[1][115] , \round_in[1][114] , 
        \round_in[1][113] , \round_in[1][112] , \round_in[1][111] , 
        \round_in[1][110] , \round_in[1][109] , \round_in[1][108] , 
        \round_in[1][107] , \round_in[1][106] , \round_in[1][105] , 
        \round_in[1][104] , \round_in[1][103] , \round_in[1][102] , 
        \round_in[1][101] , \round_in[1][100] , \round_in[1][99] , 
        \round_in[1][98] , \round_in[1][97] , \round_in[1][96] , 
        \round_in[1][95] , \round_in[1][94] , \round_in[1][93] , 
        \round_in[1][92] , \round_in[1][91] , \round_in[1][90] , 
        \round_in[1][89] , \round_in[1][88] , \round_in[1][87] , 
        \round_in[1][86] , \round_in[1][85] , \round_in[1][84] , 
        \round_in[1][83] , \round_in[1][82] , \round_in[1][81] , 
        \round_in[1][80] , \round_in[1][79] , \round_in[1][78] , 
        \round_in[1][77] , \round_in[1][76] , \round_in[1][75] , 
        \round_in[1][74] , \round_in[1][73] , \round_in[1][72] , 
        \round_in[1][71] , \round_in[1][70] , \round_in[1][69] , 
        \round_in[1][68] , \round_in[1][67] , \round_in[1][66] , 
        \round_in[1][65] , \round_in[1][64] , \round_in[1][63] , 
        \round_in[1][62] , \round_in[1][61] , \round_in[1][60] , 
        \round_in[1][59] , \round_in[1][58] , \round_in[1][57] , 
        \round_in[1][56] , \round_in[1][55] , \round_in[1][54] , 
        \round_in[1][53] , \round_in[1][52] , \round_in[1][51] , 
        \round_in[1][50] , \round_in[1][49] , \round_in[1][48] , 
        \round_in[1][47] , \round_in[1][46] , \round_in[1][45] , 
        \round_in[1][44] , \round_in[1][43] , \round_in[1][42] , 
        \round_in[1][41] , \round_in[1][40] , \round_in[1][39] , 
        \round_in[1][38] , \round_in[1][37] , \round_in[1][36] , 
        \round_in[1][35] , \round_in[1][34] , \round_in[1][33] , 
        \round_in[1][32] , \round_in[1][31] , \round_in[1][30] , 
        \round_in[1][29] , \round_in[1][28] , \round_in[1][27] , 
        \round_in[1][26] , \round_in[1][25] , \round_in[1][24] , 
        \round_in[1][23] , \round_in[1][22] , \round_in[1][21] , 
        \round_in[1][20] , \round_in[1][19] , \round_in[1][18] , 
        \round_in[1][17] , \round_in[1][16] , \round_in[1][15] , 
        \round_in[1][14] , \round_in[1][13] , \round_in[1][12] , 
        \round_in[1][11] , \round_in[1][10] , \round_in[1][9] , 
        \round_in[1][8] , \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , 
        \round_in[1][4] , \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , 
        \round_in[1][0] }) );
  round_5 \ROUND[1].round_  ( .in({\round_in[1][1599] , \round_in[1][1598] , 
        \round_in[1][1597] , \round_in[1][1596] , \round_in[1][1595] , 
        \round_in[1][1594] , \round_in[1][1593] , \round_in[1][1592] , 
        \round_in[1][1591] , \round_in[1][1590] , \round_in[1][1589] , 
        \round_in[1][1588] , \round_in[1][1587] , \round_in[1][1586] , 
        \round_in[1][1585] , \round_in[1][1584] , \round_in[1][1583] , 
        \round_in[1][1582] , \round_in[1][1581] , \round_in[1][1580] , 
        \round_in[1][1579] , \round_in[1][1578] , \round_in[1][1577] , 
        \round_in[1][1576] , \round_in[1][1575] , \round_in[1][1574] , 
        \round_in[1][1573] , \round_in[1][1572] , \round_in[1][1571] , 
        \round_in[1][1570] , \round_in[1][1569] , \round_in[1][1568] , 
        \round_in[1][1567] , \round_in[1][1566] , \round_in[1][1565] , 
        \round_in[1][1564] , \round_in[1][1563] , \round_in[1][1562] , 
        \round_in[1][1561] , \round_in[1][1560] , \round_in[1][1559] , 
        \round_in[1][1558] , \round_in[1][1557] , \round_in[1][1556] , 
        \round_in[1][1555] , \round_in[1][1554] , \round_in[1][1553] , 
        \round_in[1][1552] , \round_in[1][1551] , \round_in[1][1550] , 
        \round_in[1][1549] , \round_in[1][1548] , \round_in[1][1547] , 
        \round_in[1][1546] , \round_in[1][1545] , \round_in[1][1544] , 
        \round_in[1][1543] , \round_in[1][1542] , \round_in[1][1541] , 
        \round_in[1][1540] , \round_in[1][1539] , \round_in[1][1538] , 
        \round_in[1][1537] , \round_in[1][1536] , \round_in[1][1535] , 
        \round_in[1][1534] , \round_in[1][1533] , \round_in[1][1532] , 
        \round_in[1][1531] , \round_in[1][1530] , \round_in[1][1529] , 
        \round_in[1][1528] , \round_in[1][1527] , \round_in[1][1526] , 
        \round_in[1][1525] , \round_in[1][1524] , \round_in[1][1523] , 
        \round_in[1][1522] , \round_in[1][1521] , \round_in[1][1520] , 
        \round_in[1][1519] , \round_in[1][1518] , \round_in[1][1517] , 
        \round_in[1][1516] , \round_in[1][1515] , \round_in[1][1514] , 
        \round_in[1][1513] , \round_in[1][1512] , \round_in[1][1511] , 
        \round_in[1][1510] , \round_in[1][1509] , \round_in[1][1508] , 
        \round_in[1][1507] , \round_in[1][1506] , \round_in[1][1505] , 
        \round_in[1][1504] , \round_in[1][1503] , \round_in[1][1502] , 
        \round_in[1][1501] , \round_in[1][1500] , \round_in[1][1499] , 
        \round_in[1][1498] , \round_in[1][1497] , \round_in[1][1496] , 
        \round_in[1][1495] , \round_in[1][1494] , \round_in[1][1493] , 
        \round_in[1][1492] , \round_in[1][1491] , \round_in[1][1490] , 
        \round_in[1][1489] , \round_in[1][1488] , \round_in[1][1487] , 
        \round_in[1][1486] , \round_in[1][1485] , \round_in[1][1484] , 
        \round_in[1][1483] , \round_in[1][1482] , \round_in[1][1481] , 
        \round_in[1][1480] , \round_in[1][1479] , \round_in[1][1478] , 
        \round_in[1][1477] , \round_in[1][1476] , \round_in[1][1475] , 
        \round_in[1][1474] , \round_in[1][1473] , \round_in[1][1472] , 
        \round_in[1][1471] , \round_in[1][1470] , \round_in[1][1469] , 
        \round_in[1][1468] , \round_in[1][1467] , \round_in[1][1466] , 
        \round_in[1][1465] , \round_in[1][1464] , \round_in[1][1463] , 
        \round_in[1][1462] , \round_in[1][1461] , \round_in[1][1460] , 
        \round_in[1][1459] , \round_in[1][1458] , \round_in[1][1457] , 
        \round_in[1][1456] , \round_in[1][1455] , \round_in[1][1454] , 
        \round_in[1][1453] , \round_in[1][1452] , \round_in[1][1451] , 
        \round_in[1][1450] , \round_in[1][1449] , \round_in[1][1448] , 
        \round_in[1][1447] , \round_in[1][1446] , \round_in[1][1445] , 
        \round_in[1][1444] , \round_in[1][1443] , \round_in[1][1442] , 
        \round_in[1][1441] , \round_in[1][1440] , \round_in[1][1439] , 
        \round_in[1][1438] , \round_in[1][1437] , \round_in[1][1436] , 
        \round_in[1][1435] , \round_in[1][1434] , \round_in[1][1433] , 
        \round_in[1][1432] , \round_in[1][1431] , \round_in[1][1430] , 
        \round_in[1][1429] , \round_in[1][1428] , \round_in[1][1427] , 
        \round_in[1][1426] , \round_in[1][1425] , \round_in[1][1424] , 
        \round_in[1][1423] , \round_in[1][1422] , \round_in[1][1421] , 
        \round_in[1][1420] , \round_in[1][1419] , \round_in[1][1418] , 
        \round_in[1][1417] , \round_in[1][1416] , \round_in[1][1415] , 
        \round_in[1][1414] , \round_in[1][1413] , \round_in[1][1412] , 
        \round_in[1][1411] , \round_in[1][1410] , \round_in[1][1409] , 
        \round_in[1][1408] , \round_in[1][1407] , \round_in[1][1406] , 
        \round_in[1][1405] , \round_in[1][1404] , \round_in[1][1403] , 
        \round_in[1][1402] , \round_in[1][1401] , \round_in[1][1400] , 
        \round_in[1][1399] , \round_in[1][1398] , \round_in[1][1397] , 
        \round_in[1][1396] , \round_in[1][1395] , \round_in[1][1394] , 
        \round_in[1][1393] , \round_in[1][1392] , \round_in[1][1391] , 
        \round_in[1][1390] , \round_in[1][1389] , \round_in[1][1388] , 
        \round_in[1][1387] , \round_in[1][1386] , \round_in[1][1385] , 
        \round_in[1][1384] , \round_in[1][1383] , \round_in[1][1382] , 
        \round_in[1][1381] , \round_in[1][1380] , \round_in[1][1379] , 
        \round_in[1][1378] , \round_in[1][1377] , \round_in[1][1376] , 
        \round_in[1][1375] , \round_in[1][1374] , \round_in[1][1373] , 
        \round_in[1][1372] , \round_in[1][1371] , \round_in[1][1370] , 
        \round_in[1][1369] , \round_in[1][1368] , \round_in[1][1367] , 
        \round_in[1][1366] , \round_in[1][1365] , \round_in[1][1364] , 
        \round_in[1][1363] , \round_in[1][1362] , \round_in[1][1361] , 
        \round_in[1][1360] , \round_in[1][1359] , \round_in[1][1358] , 
        \round_in[1][1357] , \round_in[1][1356] , \round_in[1][1355] , 
        \round_in[1][1354] , \round_in[1][1353] , \round_in[1][1352] , 
        \round_in[1][1351] , \round_in[1][1350] , \round_in[1][1349] , 
        \round_in[1][1348] , \round_in[1][1347] , \round_in[1][1346] , 
        \round_in[1][1345] , \round_in[1][1344] , \round_in[1][1343] , 
        \round_in[1][1342] , \round_in[1][1341] , \round_in[1][1340] , 
        \round_in[1][1339] , \round_in[1][1338] , \round_in[1][1337] , 
        \round_in[1][1336] , \round_in[1][1335] , \round_in[1][1334] , 
        \round_in[1][1333] , \round_in[1][1332] , \round_in[1][1331] , 
        \round_in[1][1330] , \round_in[1][1329] , \round_in[1][1328] , 
        \round_in[1][1327] , \round_in[1][1326] , \round_in[1][1325] , 
        \round_in[1][1324] , \round_in[1][1323] , \round_in[1][1322] , 
        \round_in[1][1321] , \round_in[1][1320] , \round_in[1][1319] , 
        \round_in[1][1318] , \round_in[1][1317] , \round_in[1][1316] , 
        \round_in[1][1315] , \round_in[1][1314] , \round_in[1][1313] , 
        \round_in[1][1312] , \round_in[1][1311] , \round_in[1][1310] , 
        \round_in[1][1309] , \round_in[1][1308] , \round_in[1][1307] , 
        \round_in[1][1306] , \round_in[1][1305] , \round_in[1][1304] , 
        \round_in[1][1303] , \round_in[1][1302] , \round_in[1][1301] , 
        \round_in[1][1300] , \round_in[1][1299] , \round_in[1][1298] , 
        \round_in[1][1297] , \round_in[1][1296] , \round_in[1][1295] , 
        \round_in[1][1294] , \round_in[1][1293] , \round_in[1][1292] , 
        \round_in[1][1291] , \round_in[1][1290] , \round_in[1][1289] , 
        \round_in[1][1288] , \round_in[1][1287] , \round_in[1][1286] , 
        \round_in[1][1285] , \round_in[1][1284] , \round_in[1][1283] , 
        \round_in[1][1282] , \round_in[1][1281] , \round_in[1][1280] , 
        \round_in[1][1279] , \round_in[1][1278] , \round_in[1][1277] , 
        \round_in[1][1276] , \round_in[1][1275] , \round_in[1][1274] , 
        \round_in[1][1273] , \round_in[1][1272] , \round_in[1][1271] , 
        \round_in[1][1270] , \round_in[1][1269] , \round_in[1][1268] , 
        \round_in[1][1267] , \round_in[1][1266] , \round_in[1][1265] , 
        \round_in[1][1264] , \round_in[1][1263] , \round_in[1][1262] , 
        \round_in[1][1261] , \round_in[1][1260] , \round_in[1][1259] , 
        \round_in[1][1258] , \round_in[1][1257] , \round_in[1][1256] , 
        \round_in[1][1255] , \round_in[1][1254] , \round_in[1][1253] , 
        \round_in[1][1252] , \round_in[1][1251] , \round_in[1][1250] , 
        \round_in[1][1249] , \round_in[1][1248] , \round_in[1][1247] , 
        \round_in[1][1246] , \round_in[1][1245] , \round_in[1][1244] , 
        \round_in[1][1243] , \round_in[1][1242] , \round_in[1][1241] , 
        \round_in[1][1240] , \round_in[1][1239] , \round_in[1][1238] , 
        \round_in[1][1237] , \round_in[1][1236] , \round_in[1][1235] , 
        \round_in[1][1234] , \round_in[1][1233] , \round_in[1][1232] , 
        \round_in[1][1231] , \round_in[1][1230] , \round_in[1][1229] , 
        \round_in[1][1228] , \round_in[1][1227] , \round_in[1][1226] , 
        \round_in[1][1225] , \round_in[1][1224] , \round_in[1][1223] , 
        \round_in[1][1222] , \round_in[1][1221] , \round_in[1][1220] , 
        \round_in[1][1219] , \round_in[1][1218] , \round_in[1][1217] , 
        \round_in[1][1216] , \round_in[1][1215] , \round_in[1][1214] , 
        \round_in[1][1213] , \round_in[1][1212] , \round_in[1][1211] , 
        \round_in[1][1210] , \round_in[1][1209] , \round_in[1][1208] , 
        \round_in[1][1207] , \round_in[1][1206] , \round_in[1][1205] , 
        \round_in[1][1204] , \round_in[1][1203] , \round_in[1][1202] , 
        \round_in[1][1201] , \round_in[1][1200] , \round_in[1][1199] , 
        \round_in[1][1198] , \round_in[1][1197] , \round_in[1][1196] , 
        \round_in[1][1195] , \round_in[1][1194] , \round_in[1][1193] , 
        \round_in[1][1192] , \round_in[1][1191] , \round_in[1][1190] , 
        \round_in[1][1189] , \round_in[1][1188] , \round_in[1][1187] , 
        \round_in[1][1186] , \round_in[1][1185] , \round_in[1][1184] , 
        \round_in[1][1183] , \round_in[1][1182] , \round_in[1][1181] , 
        \round_in[1][1180] , \round_in[1][1179] , \round_in[1][1178] , 
        \round_in[1][1177] , \round_in[1][1176] , \round_in[1][1175] , 
        \round_in[1][1174] , \round_in[1][1173] , \round_in[1][1172] , 
        \round_in[1][1171] , \round_in[1][1170] , \round_in[1][1169] , 
        \round_in[1][1168] , \round_in[1][1167] , \round_in[1][1166] , 
        \round_in[1][1165] , \round_in[1][1164] , \round_in[1][1163] , 
        \round_in[1][1162] , \round_in[1][1161] , \round_in[1][1160] , 
        \round_in[1][1159] , \round_in[1][1158] , \round_in[1][1157] , 
        \round_in[1][1156] , \round_in[1][1155] , \round_in[1][1154] , 
        \round_in[1][1153] , \round_in[1][1152] , \round_in[1][1151] , 
        \round_in[1][1150] , \round_in[1][1149] , \round_in[1][1148] , 
        \round_in[1][1147] , \round_in[1][1146] , \round_in[1][1145] , 
        \round_in[1][1144] , \round_in[1][1143] , \round_in[1][1142] , 
        \round_in[1][1141] , \round_in[1][1140] , \round_in[1][1139] , 
        \round_in[1][1138] , \round_in[1][1137] , \round_in[1][1136] , 
        \round_in[1][1135] , \round_in[1][1134] , \round_in[1][1133] , 
        \round_in[1][1132] , \round_in[1][1131] , \round_in[1][1130] , 
        \round_in[1][1129] , \round_in[1][1128] , \round_in[1][1127] , 
        \round_in[1][1126] , \round_in[1][1125] , \round_in[1][1124] , 
        \round_in[1][1123] , \round_in[1][1122] , \round_in[1][1121] , 
        \round_in[1][1120] , \round_in[1][1119] , \round_in[1][1118] , 
        \round_in[1][1117] , \round_in[1][1116] , \round_in[1][1115] , 
        \round_in[1][1114] , \round_in[1][1113] , \round_in[1][1112] , 
        \round_in[1][1111] , \round_in[1][1110] , \round_in[1][1109] , 
        \round_in[1][1108] , \round_in[1][1107] , \round_in[1][1106] , 
        \round_in[1][1105] , \round_in[1][1104] , \round_in[1][1103] , 
        \round_in[1][1102] , \round_in[1][1101] , \round_in[1][1100] , 
        \round_in[1][1099] , \round_in[1][1098] , \round_in[1][1097] , 
        \round_in[1][1096] , \round_in[1][1095] , \round_in[1][1094] , 
        \round_in[1][1093] , \round_in[1][1092] , \round_in[1][1091] , 
        \round_in[1][1090] , \round_in[1][1089] , \round_in[1][1088] , 
        \round_in[1][1087] , \round_in[1][1086] , \round_in[1][1085] , 
        \round_in[1][1084] , \round_in[1][1083] , \round_in[1][1082] , 
        \round_in[1][1081] , \round_in[1][1080] , \round_in[1][1079] , 
        \round_in[1][1078] , \round_in[1][1077] , \round_in[1][1076] , 
        \round_in[1][1075] , \round_in[1][1074] , \round_in[1][1073] , 
        \round_in[1][1072] , \round_in[1][1071] , \round_in[1][1070] , 
        \round_in[1][1069] , \round_in[1][1068] , \round_in[1][1067] , 
        \round_in[1][1066] , \round_in[1][1065] , \round_in[1][1064] , 
        \round_in[1][1063] , \round_in[1][1062] , \round_in[1][1061] , 
        \round_in[1][1060] , \round_in[1][1059] , \round_in[1][1058] , 
        \round_in[1][1057] , \round_in[1][1056] , \round_in[1][1055] , 
        \round_in[1][1054] , \round_in[1][1053] , \round_in[1][1052] , 
        \round_in[1][1051] , \round_in[1][1050] , \round_in[1][1049] , 
        \round_in[1][1048] , \round_in[1][1047] , \round_in[1][1046] , 
        \round_in[1][1045] , \round_in[1][1044] , \round_in[1][1043] , 
        \round_in[1][1042] , \round_in[1][1041] , \round_in[1][1040] , 
        \round_in[1][1039] , \round_in[1][1038] , \round_in[1][1037] , 
        \round_in[1][1036] , \round_in[1][1035] , \round_in[1][1034] , 
        \round_in[1][1033] , \round_in[1][1032] , \round_in[1][1031] , 
        \round_in[1][1030] , \round_in[1][1029] , \round_in[1][1028] , 
        \round_in[1][1027] , \round_in[1][1026] , \round_in[1][1025] , 
        \round_in[1][1024] , \round_in[1][1023] , \round_in[1][1022] , 
        \round_in[1][1021] , \round_in[1][1020] , \round_in[1][1019] , 
        \round_in[1][1018] , \round_in[1][1017] , \round_in[1][1016] , 
        \round_in[1][1015] , \round_in[1][1014] , \round_in[1][1013] , 
        \round_in[1][1012] , \round_in[1][1011] , \round_in[1][1010] , 
        \round_in[1][1009] , \round_in[1][1008] , \round_in[1][1007] , 
        \round_in[1][1006] , \round_in[1][1005] , \round_in[1][1004] , 
        \round_in[1][1003] , \round_in[1][1002] , \round_in[1][1001] , 
        \round_in[1][1000] , \round_in[1][999] , \round_in[1][998] , 
        \round_in[1][997] , \round_in[1][996] , \round_in[1][995] , 
        \round_in[1][994] , \round_in[1][993] , \round_in[1][992] , 
        \round_in[1][991] , \round_in[1][990] , \round_in[1][989] , 
        \round_in[1][988] , \round_in[1][987] , \round_in[1][986] , 
        \round_in[1][985] , \round_in[1][984] , \round_in[1][983] , 
        \round_in[1][982] , \round_in[1][981] , \round_in[1][980] , 
        \round_in[1][979] , \round_in[1][978] , \round_in[1][977] , 
        \round_in[1][976] , \round_in[1][975] , \round_in[1][974] , 
        \round_in[1][973] , \round_in[1][972] , \round_in[1][971] , 
        \round_in[1][970] , \round_in[1][969] , \round_in[1][968] , 
        \round_in[1][967] , \round_in[1][966] , \round_in[1][965] , 
        \round_in[1][964] , \round_in[1][963] , \round_in[1][962] , 
        \round_in[1][961] , \round_in[1][960] , \round_in[1][959] , 
        \round_in[1][958] , \round_in[1][957] , \round_in[1][956] , 
        \round_in[1][955] , \round_in[1][954] , \round_in[1][953] , 
        \round_in[1][952] , \round_in[1][951] , \round_in[1][950] , 
        \round_in[1][949] , \round_in[1][948] , \round_in[1][947] , 
        \round_in[1][946] , \round_in[1][945] , \round_in[1][944] , 
        \round_in[1][943] , \round_in[1][942] , \round_in[1][941] , 
        \round_in[1][940] , \round_in[1][939] , \round_in[1][938] , 
        \round_in[1][937] , \round_in[1][936] , \round_in[1][935] , 
        \round_in[1][934] , \round_in[1][933] , \round_in[1][932] , 
        \round_in[1][931] , \round_in[1][930] , \round_in[1][929] , 
        \round_in[1][928] , \round_in[1][927] , \round_in[1][926] , 
        \round_in[1][925] , \round_in[1][924] , \round_in[1][923] , 
        \round_in[1][922] , \round_in[1][921] , \round_in[1][920] , 
        \round_in[1][919] , \round_in[1][918] , \round_in[1][917] , 
        \round_in[1][916] , \round_in[1][915] , \round_in[1][914] , 
        \round_in[1][913] , \round_in[1][912] , \round_in[1][911] , 
        \round_in[1][910] , \round_in[1][909] , \round_in[1][908] , 
        \round_in[1][907] , \round_in[1][906] , \round_in[1][905] , 
        \round_in[1][904] , \round_in[1][903] , \round_in[1][902] , 
        \round_in[1][901] , \round_in[1][900] , \round_in[1][899] , 
        \round_in[1][898] , \round_in[1][897] , \round_in[1][896] , 
        \round_in[1][895] , \round_in[1][894] , \round_in[1][893] , 
        \round_in[1][892] , \round_in[1][891] , \round_in[1][890] , 
        \round_in[1][889] , \round_in[1][888] , \round_in[1][887] , 
        \round_in[1][886] , \round_in[1][885] , \round_in[1][884] , 
        \round_in[1][883] , \round_in[1][882] , \round_in[1][881] , 
        \round_in[1][880] , \round_in[1][879] , \round_in[1][878] , 
        \round_in[1][877] , \round_in[1][876] , \round_in[1][875] , 
        \round_in[1][874] , \round_in[1][873] , \round_in[1][872] , 
        \round_in[1][871] , \round_in[1][870] , \round_in[1][869] , 
        \round_in[1][868] , \round_in[1][867] , \round_in[1][866] , 
        \round_in[1][865] , \round_in[1][864] , \round_in[1][863] , 
        \round_in[1][862] , \round_in[1][861] , \round_in[1][860] , 
        \round_in[1][859] , \round_in[1][858] , \round_in[1][857] , 
        \round_in[1][856] , \round_in[1][855] , \round_in[1][854] , 
        \round_in[1][853] , \round_in[1][852] , \round_in[1][851] , 
        \round_in[1][850] , \round_in[1][849] , \round_in[1][848] , 
        \round_in[1][847] , \round_in[1][846] , \round_in[1][845] , 
        \round_in[1][844] , \round_in[1][843] , \round_in[1][842] , 
        \round_in[1][841] , \round_in[1][840] , \round_in[1][839] , 
        \round_in[1][838] , \round_in[1][837] , \round_in[1][836] , 
        \round_in[1][835] , \round_in[1][834] , \round_in[1][833] , 
        \round_in[1][832] , \round_in[1][831] , \round_in[1][830] , 
        \round_in[1][829] , \round_in[1][828] , \round_in[1][827] , 
        \round_in[1][826] , \round_in[1][825] , \round_in[1][824] , 
        \round_in[1][823] , \round_in[1][822] , \round_in[1][821] , 
        \round_in[1][820] , \round_in[1][819] , \round_in[1][818] , 
        \round_in[1][817] , \round_in[1][816] , \round_in[1][815] , 
        \round_in[1][814] , \round_in[1][813] , \round_in[1][812] , 
        \round_in[1][811] , \round_in[1][810] , \round_in[1][809] , 
        \round_in[1][808] , \round_in[1][807] , \round_in[1][806] , 
        \round_in[1][805] , \round_in[1][804] , \round_in[1][803] , 
        \round_in[1][802] , \round_in[1][801] , \round_in[1][800] , 
        \round_in[1][799] , \round_in[1][798] , \round_in[1][797] , 
        \round_in[1][796] , \round_in[1][795] , \round_in[1][794] , 
        \round_in[1][793] , \round_in[1][792] , \round_in[1][791] , 
        \round_in[1][790] , \round_in[1][789] , \round_in[1][788] , 
        \round_in[1][787] , \round_in[1][786] , \round_in[1][785] , 
        \round_in[1][784] , \round_in[1][783] , \round_in[1][782] , 
        \round_in[1][781] , \round_in[1][780] , \round_in[1][779] , 
        \round_in[1][778] , \round_in[1][777] , \round_in[1][776] , 
        \round_in[1][775] , \round_in[1][774] , \round_in[1][773] , 
        \round_in[1][772] , \round_in[1][771] , \round_in[1][770] , 
        \round_in[1][769] , \round_in[1][768] , \round_in[1][767] , 
        \round_in[1][766] , \round_in[1][765] , \round_in[1][764] , 
        \round_in[1][763] , \round_in[1][762] , \round_in[1][761] , 
        \round_in[1][760] , \round_in[1][759] , \round_in[1][758] , 
        \round_in[1][757] , \round_in[1][756] , \round_in[1][755] , 
        \round_in[1][754] , \round_in[1][753] , \round_in[1][752] , 
        \round_in[1][751] , \round_in[1][750] , \round_in[1][749] , 
        \round_in[1][748] , \round_in[1][747] , \round_in[1][746] , 
        \round_in[1][745] , \round_in[1][744] , \round_in[1][743] , 
        \round_in[1][742] , \round_in[1][741] , \round_in[1][740] , 
        \round_in[1][739] , \round_in[1][738] , \round_in[1][737] , 
        \round_in[1][736] , \round_in[1][735] , \round_in[1][734] , 
        \round_in[1][733] , \round_in[1][732] , \round_in[1][731] , 
        \round_in[1][730] , \round_in[1][729] , \round_in[1][728] , 
        \round_in[1][727] , \round_in[1][726] , \round_in[1][725] , 
        \round_in[1][724] , \round_in[1][723] , \round_in[1][722] , 
        \round_in[1][721] , \round_in[1][720] , \round_in[1][719] , 
        \round_in[1][718] , \round_in[1][717] , \round_in[1][716] , 
        \round_in[1][715] , \round_in[1][714] , \round_in[1][713] , 
        \round_in[1][712] , \round_in[1][711] , \round_in[1][710] , 
        \round_in[1][709] , \round_in[1][708] , \round_in[1][707] , 
        \round_in[1][706] , \round_in[1][705] , \round_in[1][704] , 
        \round_in[1][703] , \round_in[1][702] , \round_in[1][701] , 
        \round_in[1][700] , \round_in[1][699] , \round_in[1][698] , 
        \round_in[1][697] , \round_in[1][696] , \round_in[1][695] , 
        \round_in[1][694] , \round_in[1][693] , \round_in[1][692] , 
        \round_in[1][691] , \round_in[1][690] , \round_in[1][689] , 
        \round_in[1][688] , \round_in[1][687] , \round_in[1][686] , 
        \round_in[1][685] , \round_in[1][684] , \round_in[1][683] , 
        \round_in[1][682] , \round_in[1][681] , \round_in[1][680] , 
        \round_in[1][679] , \round_in[1][678] , \round_in[1][677] , 
        \round_in[1][676] , \round_in[1][675] , \round_in[1][674] , 
        \round_in[1][673] , \round_in[1][672] , \round_in[1][671] , 
        \round_in[1][670] , \round_in[1][669] , \round_in[1][668] , 
        \round_in[1][667] , \round_in[1][666] , \round_in[1][665] , 
        \round_in[1][664] , \round_in[1][663] , \round_in[1][662] , 
        \round_in[1][661] , \round_in[1][660] , \round_in[1][659] , 
        \round_in[1][658] , \round_in[1][657] , \round_in[1][656] , 
        \round_in[1][655] , \round_in[1][654] , \round_in[1][653] , 
        \round_in[1][652] , \round_in[1][651] , \round_in[1][650] , 
        \round_in[1][649] , \round_in[1][648] , \round_in[1][647] , 
        \round_in[1][646] , \round_in[1][645] , \round_in[1][644] , 
        \round_in[1][643] , \round_in[1][642] , \round_in[1][641] , 
        \round_in[1][640] , \round_in[1][639] , \round_in[1][638] , 
        \round_in[1][637] , \round_in[1][636] , \round_in[1][635] , 
        \round_in[1][634] , \round_in[1][633] , \round_in[1][632] , 
        \round_in[1][631] , \round_in[1][630] , \round_in[1][629] , 
        \round_in[1][628] , \round_in[1][627] , \round_in[1][626] , 
        \round_in[1][625] , \round_in[1][624] , \round_in[1][623] , 
        \round_in[1][622] , \round_in[1][621] , \round_in[1][620] , 
        \round_in[1][619] , \round_in[1][618] , \round_in[1][617] , 
        \round_in[1][616] , \round_in[1][615] , \round_in[1][614] , 
        \round_in[1][613] , \round_in[1][612] , \round_in[1][611] , 
        \round_in[1][610] , \round_in[1][609] , \round_in[1][608] , 
        \round_in[1][607] , \round_in[1][606] , \round_in[1][605] , 
        \round_in[1][604] , \round_in[1][603] , \round_in[1][602] , 
        \round_in[1][601] , \round_in[1][600] , \round_in[1][599] , 
        \round_in[1][598] , \round_in[1][597] , \round_in[1][596] , 
        \round_in[1][595] , \round_in[1][594] , \round_in[1][593] , 
        \round_in[1][592] , \round_in[1][591] , \round_in[1][590] , 
        \round_in[1][589] , \round_in[1][588] , \round_in[1][587] , 
        \round_in[1][586] , \round_in[1][585] , \round_in[1][584] , 
        \round_in[1][583] , \round_in[1][582] , \round_in[1][581] , 
        \round_in[1][580] , \round_in[1][579] , \round_in[1][578] , 
        \round_in[1][577] , \round_in[1][576] , \round_in[1][575] , 
        \round_in[1][574] , \round_in[1][573] , \round_in[1][572] , 
        \round_in[1][571] , \round_in[1][570] , \round_in[1][569] , 
        \round_in[1][568] , \round_in[1][567] , \round_in[1][566] , 
        \round_in[1][565] , \round_in[1][564] , \round_in[1][563] , 
        \round_in[1][562] , \round_in[1][561] , \round_in[1][560] , 
        \round_in[1][559] , \round_in[1][558] , \round_in[1][557] , 
        \round_in[1][556] , \round_in[1][555] , \round_in[1][554] , 
        \round_in[1][553] , \round_in[1][552] , \round_in[1][551] , 
        \round_in[1][550] , \round_in[1][549] , \round_in[1][548] , 
        \round_in[1][547] , \round_in[1][546] , \round_in[1][545] , 
        \round_in[1][544] , \round_in[1][543] , \round_in[1][542] , 
        \round_in[1][541] , \round_in[1][540] , \round_in[1][539] , 
        \round_in[1][538] , \round_in[1][537] , \round_in[1][536] , 
        \round_in[1][535] , \round_in[1][534] , \round_in[1][533] , 
        \round_in[1][532] , \round_in[1][531] , \round_in[1][530] , 
        \round_in[1][529] , \round_in[1][528] , \round_in[1][527] , 
        \round_in[1][526] , \round_in[1][525] , \round_in[1][524] , 
        \round_in[1][523] , \round_in[1][522] , \round_in[1][521] , 
        \round_in[1][520] , \round_in[1][519] , \round_in[1][518] , 
        \round_in[1][517] , \round_in[1][516] , \round_in[1][515] , 
        \round_in[1][514] , \round_in[1][513] , \round_in[1][512] , 
        \round_in[1][511] , \round_in[1][510] , \round_in[1][509] , 
        \round_in[1][508] , \round_in[1][507] , \round_in[1][506] , 
        \round_in[1][505] , \round_in[1][504] , \round_in[1][503] , 
        \round_in[1][502] , \round_in[1][501] , \round_in[1][500] , 
        \round_in[1][499] , \round_in[1][498] , \round_in[1][497] , 
        \round_in[1][496] , \round_in[1][495] , \round_in[1][494] , 
        \round_in[1][493] , \round_in[1][492] , \round_in[1][491] , 
        \round_in[1][490] , \round_in[1][489] , \round_in[1][488] , 
        \round_in[1][487] , \round_in[1][486] , \round_in[1][485] , 
        \round_in[1][484] , \round_in[1][483] , \round_in[1][482] , 
        \round_in[1][481] , \round_in[1][480] , \round_in[1][479] , 
        \round_in[1][478] , \round_in[1][477] , \round_in[1][476] , 
        \round_in[1][475] , \round_in[1][474] , \round_in[1][473] , 
        \round_in[1][472] , \round_in[1][471] , \round_in[1][470] , 
        \round_in[1][469] , \round_in[1][468] , \round_in[1][467] , 
        \round_in[1][466] , \round_in[1][465] , \round_in[1][464] , 
        \round_in[1][463] , \round_in[1][462] , \round_in[1][461] , 
        \round_in[1][460] , \round_in[1][459] , \round_in[1][458] , 
        \round_in[1][457] , \round_in[1][456] , \round_in[1][455] , 
        \round_in[1][454] , \round_in[1][453] , \round_in[1][452] , 
        \round_in[1][451] , \round_in[1][450] , \round_in[1][449] , 
        \round_in[1][448] , \round_in[1][447] , \round_in[1][446] , 
        \round_in[1][445] , \round_in[1][444] , \round_in[1][443] , 
        \round_in[1][442] , \round_in[1][441] , \round_in[1][440] , 
        \round_in[1][439] , \round_in[1][438] , \round_in[1][437] , 
        \round_in[1][436] , \round_in[1][435] , \round_in[1][434] , 
        \round_in[1][433] , \round_in[1][432] , \round_in[1][431] , 
        \round_in[1][430] , \round_in[1][429] , \round_in[1][428] , 
        \round_in[1][427] , \round_in[1][426] , \round_in[1][425] , 
        \round_in[1][424] , \round_in[1][423] , \round_in[1][422] , 
        \round_in[1][421] , \round_in[1][420] , \round_in[1][419] , 
        \round_in[1][418] , \round_in[1][417] , \round_in[1][416] , 
        \round_in[1][415] , \round_in[1][414] , \round_in[1][413] , 
        \round_in[1][412] , \round_in[1][411] , \round_in[1][410] , 
        \round_in[1][409] , \round_in[1][408] , \round_in[1][407] , 
        \round_in[1][406] , \round_in[1][405] , \round_in[1][404] , 
        \round_in[1][403] , \round_in[1][402] , \round_in[1][401] , 
        \round_in[1][400] , \round_in[1][399] , \round_in[1][398] , 
        \round_in[1][397] , \round_in[1][396] , \round_in[1][395] , 
        \round_in[1][394] , \round_in[1][393] , \round_in[1][392] , 
        \round_in[1][391] , \round_in[1][390] , \round_in[1][389] , 
        \round_in[1][388] , \round_in[1][387] , \round_in[1][386] , 
        \round_in[1][385] , \round_in[1][384] , \round_in[1][383] , 
        \round_in[1][382] , \round_in[1][381] , \round_in[1][380] , 
        \round_in[1][379] , \round_in[1][378] , \round_in[1][377] , 
        \round_in[1][376] , \round_in[1][375] , \round_in[1][374] , 
        \round_in[1][373] , \round_in[1][372] , \round_in[1][371] , 
        \round_in[1][370] , \round_in[1][369] , \round_in[1][368] , 
        \round_in[1][367] , \round_in[1][366] , \round_in[1][365] , 
        \round_in[1][364] , \round_in[1][363] , \round_in[1][362] , 
        \round_in[1][361] , \round_in[1][360] , \round_in[1][359] , 
        \round_in[1][358] , \round_in[1][357] , \round_in[1][356] , 
        \round_in[1][355] , \round_in[1][354] , \round_in[1][353] , 
        \round_in[1][352] , \round_in[1][351] , \round_in[1][350] , 
        \round_in[1][349] , \round_in[1][348] , \round_in[1][347] , 
        \round_in[1][346] , \round_in[1][345] , \round_in[1][344] , 
        \round_in[1][343] , \round_in[1][342] , \round_in[1][341] , 
        \round_in[1][340] , \round_in[1][339] , \round_in[1][338] , 
        \round_in[1][337] , \round_in[1][336] , \round_in[1][335] , 
        \round_in[1][334] , \round_in[1][333] , \round_in[1][332] , 
        \round_in[1][331] , \round_in[1][330] , \round_in[1][329] , 
        \round_in[1][328] , \round_in[1][327] , \round_in[1][326] , 
        \round_in[1][325] , \round_in[1][324] , \round_in[1][323] , 
        \round_in[1][322] , \round_in[1][321] , \round_in[1][320] , 
        \round_in[1][319] , \round_in[1][318] , \round_in[1][317] , 
        \round_in[1][316] , \round_in[1][315] , \round_in[1][314] , 
        \round_in[1][313] , \round_in[1][312] , \round_in[1][311] , 
        \round_in[1][310] , \round_in[1][309] , \round_in[1][308] , 
        \round_in[1][307] , \round_in[1][306] , \round_in[1][305] , 
        \round_in[1][304] , \round_in[1][303] , \round_in[1][302] , 
        \round_in[1][301] , \round_in[1][300] , \round_in[1][299] , 
        \round_in[1][298] , \round_in[1][297] , \round_in[1][296] , 
        \round_in[1][295] , \round_in[1][294] , \round_in[1][293] , 
        \round_in[1][292] , \round_in[1][291] , \round_in[1][290] , 
        \round_in[1][289] , \round_in[1][288] , \round_in[1][287] , 
        \round_in[1][286] , \round_in[1][285] , \round_in[1][284] , 
        \round_in[1][283] , \round_in[1][282] , \round_in[1][281] , 
        \round_in[1][280] , \round_in[1][279] , \round_in[1][278] , 
        \round_in[1][277] , \round_in[1][276] , \round_in[1][275] , 
        \round_in[1][274] , \round_in[1][273] , \round_in[1][272] , 
        \round_in[1][271] , \round_in[1][270] , \round_in[1][269] , 
        \round_in[1][268] , \round_in[1][267] , \round_in[1][266] , 
        \round_in[1][265] , \round_in[1][264] , \round_in[1][263] , 
        \round_in[1][262] , \round_in[1][261] , \round_in[1][260] , 
        \round_in[1][259] , \round_in[1][258] , \round_in[1][257] , 
        \round_in[1][256] , \round_in[1][255] , \round_in[1][254] , 
        \round_in[1][253] , \round_in[1][252] , \round_in[1][251] , 
        \round_in[1][250] , \round_in[1][249] , \round_in[1][248] , 
        \round_in[1][247] , \round_in[1][246] , \round_in[1][245] , 
        \round_in[1][244] , \round_in[1][243] , \round_in[1][242] , 
        \round_in[1][241] , \round_in[1][240] , \round_in[1][239] , 
        \round_in[1][238] , \round_in[1][237] , \round_in[1][236] , 
        \round_in[1][235] , \round_in[1][234] , \round_in[1][233] , 
        \round_in[1][232] , \round_in[1][231] , \round_in[1][230] , 
        \round_in[1][229] , \round_in[1][228] , \round_in[1][227] , 
        \round_in[1][226] , \round_in[1][225] , \round_in[1][224] , 
        \round_in[1][223] , \round_in[1][222] , \round_in[1][221] , 
        \round_in[1][220] , \round_in[1][219] , \round_in[1][218] , 
        \round_in[1][217] , \round_in[1][216] , \round_in[1][215] , 
        \round_in[1][214] , \round_in[1][213] , \round_in[1][212] , 
        \round_in[1][211] , \round_in[1][210] , \round_in[1][209] , 
        \round_in[1][208] , \round_in[1][207] , \round_in[1][206] , 
        \round_in[1][205] , \round_in[1][204] , \round_in[1][203] , 
        \round_in[1][202] , \round_in[1][201] , \round_in[1][200] , 
        \round_in[1][199] , \round_in[1][198] , \round_in[1][197] , 
        \round_in[1][196] , \round_in[1][195] , \round_in[1][194] , 
        \round_in[1][193] , \round_in[1][192] , \round_in[1][191] , 
        \round_in[1][190] , \round_in[1][189] , \round_in[1][188] , 
        \round_in[1][187] , \round_in[1][186] , \round_in[1][185] , 
        \round_in[1][184] , \round_in[1][183] , \round_in[1][182] , 
        \round_in[1][181] , \round_in[1][180] , \round_in[1][179] , 
        \round_in[1][178] , \round_in[1][177] , \round_in[1][176] , 
        \round_in[1][175] , \round_in[1][174] , \round_in[1][173] , 
        \round_in[1][172] , \round_in[1][171] , \round_in[1][170] , 
        \round_in[1][169] , \round_in[1][168] , \round_in[1][167] , 
        \round_in[1][166] , \round_in[1][165] , \round_in[1][164] , 
        \round_in[1][163] , \round_in[1][162] , \round_in[1][161] , 
        \round_in[1][160] , \round_in[1][159] , \round_in[1][158] , 
        \round_in[1][157] , \round_in[1][156] , \round_in[1][155] , 
        \round_in[1][154] , \round_in[1][153] , \round_in[1][152] , 
        \round_in[1][151] , \round_in[1][150] , \round_in[1][149] , 
        \round_in[1][148] , \round_in[1][147] , \round_in[1][146] , 
        \round_in[1][145] , \round_in[1][144] , \round_in[1][143] , 
        \round_in[1][142] , \round_in[1][141] , \round_in[1][140] , 
        \round_in[1][139] , \round_in[1][138] , \round_in[1][137] , 
        \round_in[1][136] , \round_in[1][135] , \round_in[1][134] , 
        \round_in[1][133] , \round_in[1][132] , \round_in[1][131] , 
        \round_in[1][130] , \round_in[1][129] , \round_in[1][128] , 
        \round_in[1][127] , \round_in[1][126] , \round_in[1][125] , 
        \round_in[1][124] , \round_in[1][123] , \round_in[1][122] , 
        \round_in[1][121] , \round_in[1][120] , \round_in[1][119] , 
        \round_in[1][118] , \round_in[1][117] , \round_in[1][116] , 
        \round_in[1][115] , \round_in[1][114] , \round_in[1][113] , 
        \round_in[1][112] , \round_in[1][111] , \round_in[1][110] , 
        \round_in[1][109] , \round_in[1][108] , \round_in[1][107] , 
        \round_in[1][106] , \round_in[1][105] , \round_in[1][104] , 
        \round_in[1][103] , \round_in[1][102] , \round_in[1][101] , 
        \round_in[1][100] , \round_in[1][99] , \round_in[1][98] , 
        \round_in[1][97] , \round_in[1][96] , \round_in[1][95] , 
        \round_in[1][94] , \round_in[1][93] , \round_in[1][92] , 
        \round_in[1][91] , \round_in[1][90] , \round_in[1][89] , 
        \round_in[1][88] , \round_in[1][87] , \round_in[1][86] , 
        \round_in[1][85] , \round_in[1][84] , \round_in[1][83] , 
        \round_in[1][82] , \round_in[1][81] , \round_in[1][80] , 
        \round_in[1][79] , \round_in[1][78] , \round_in[1][77] , 
        \round_in[1][76] , \round_in[1][75] , \round_in[1][74] , 
        \round_in[1][73] , \round_in[1][72] , \round_in[1][71] , 
        \round_in[1][70] , \round_in[1][69] , \round_in[1][68] , 
        \round_in[1][67] , \round_in[1][66] , \round_in[1][65] , 
        \round_in[1][64] , \round_in[1][63] , \round_in[1][62] , 
        \round_in[1][61] , \round_in[1][60] , \round_in[1][59] , 
        \round_in[1][58] , \round_in[1][57] , \round_in[1][56] , 
        \round_in[1][55] , \round_in[1][54] , \round_in[1][53] , 
        \round_in[1][52] , \round_in[1][51] , \round_in[1][50] , 
        \round_in[1][49] , \round_in[1][48] , \round_in[1][47] , 
        \round_in[1][46] , \round_in[1][45] , \round_in[1][44] , 
        \round_in[1][43] , \round_in[1][42] , \round_in[1][41] , 
        \round_in[1][40] , \round_in[1][39] , \round_in[1][38] , 
        \round_in[1][37] , \round_in[1][36] , \round_in[1][35] , 
        \round_in[1][34] , \round_in[1][33] , \round_in[1][32] , 
        \round_in[1][31] , \round_in[1][30] , \round_in[1][29] , 
        \round_in[1][28] , \round_in[1][27] , \round_in[1][26] , 
        \round_in[1][25] , \round_in[1][24] , \round_in[1][23] , 
        \round_in[1][22] , \round_in[1][21] , \round_in[1][20] , 
        \round_in[1][19] , \round_in[1][18] , \round_in[1][17] , 
        \round_in[1][16] , \round_in[1][15] , \round_in[1][14] , 
        \round_in[1][13] , \round_in[1][12] , \round_in[1][11] , 
        \round_in[1][10] , \round_in[1][9] , \round_in[1][8] , 
        \round_in[1][7] , \round_in[1][6] , \round_in[1][5] , \round_in[1][4] , 
        \round_in[1][3] , \round_in[1][2] , \round_in[1][1] , \round_in[1][0] }), .round_const({\RCONST[1].rconst_/N68 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, rc_i[1], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \RCONST[1].rconst_/N49 , 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[1][7] , 1'b0, 1'b0, 1'b0, 
        \RCONST[1].rconst_/N26 , 1'b0, \RCONST[1].rconst_/N15 , 
        \RCONST[3].rconst_/N10 }), .out({\round_in[2][1599] , 
        \round_in[2][1598] , \round_in[2][1597] , \round_in[2][1596] , 
        \round_in[2][1595] , \round_in[2][1594] , \round_in[2][1593] , 
        \round_in[2][1592] , \round_in[2][1591] , \round_in[2][1590] , 
        \round_in[2][1589] , \round_in[2][1588] , \round_in[2][1587] , 
        \round_in[2][1586] , \round_in[2][1585] , \round_in[2][1584] , 
        \round_in[2][1583] , \round_in[2][1582] , \round_in[2][1581] , 
        \round_in[2][1580] , \round_in[2][1579] , \round_in[2][1578] , 
        \round_in[2][1577] , \round_in[2][1576] , \round_in[2][1575] , 
        \round_in[2][1574] , \round_in[2][1573] , \round_in[2][1572] , 
        \round_in[2][1571] , \round_in[2][1570] , \round_in[2][1569] , 
        \round_in[2][1568] , \round_in[2][1567] , \round_in[2][1566] , 
        \round_in[2][1565] , \round_in[2][1564] , \round_in[2][1563] , 
        \round_in[2][1562] , \round_in[2][1561] , \round_in[2][1560] , 
        \round_in[2][1559] , \round_in[2][1558] , \round_in[2][1557] , 
        \round_in[2][1556] , \round_in[2][1555] , \round_in[2][1554] , 
        \round_in[2][1553] , \round_in[2][1552] , \round_in[2][1551] , 
        \round_in[2][1550] , \round_in[2][1549] , \round_in[2][1548] , 
        \round_in[2][1547] , \round_in[2][1546] , \round_in[2][1545] , 
        \round_in[2][1544] , \round_in[2][1543] , \round_in[2][1542] , 
        \round_in[2][1541] , \round_in[2][1540] , \round_in[2][1539] , 
        \round_in[2][1538] , \round_in[2][1537] , \round_in[2][1536] , 
        \round_in[2][1535] , \round_in[2][1534] , \round_in[2][1533] , 
        \round_in[2][1532] , \round_in[2][1531] , \round_in[2][1530] , 
        \round_in[2][1529] , \round_in[2][1528] , \round_in[2][1527] , 
        \round_in[2][1526] , \round_in[2][1525] , \round_in[2][1524] , 
        \round_in[2][1523] , \round_in[2][1522] , \round_in[2][1521] , 
        \round_in[2][1520] , \round_in[2][1519] , \round_in[2][1518] , 
        \round_in[2][1517] , \round_in[2][1516] , \round_in[2][1515] , 
        \round_in[2][1514] , \round_in[2][1513] , \round_in[2][1512] , 
        \round_in[2][1511] , \round_in[2][1510] , \round_in[2][1509] , 
        \round_in[2][1508] , \round_in[2][1507] , \round_in[2][1506] , 
        \round_in[2][1505] , \round_in[2][1504] , \round_in[2][1503] , 
        \round_in[2][1502] , \round_in[2][1501] , \round_in[2][1500] , 
        \round_in[2][1499] , \round_in[2][1498] , \round_in[2][1497] , 
        \round_in[2][1496] , \round_in[2][1495] , \round_in[2][1494] , 
        \round_in[2][1493] , \round_in[2][1492] , \round_in[2][1491] , 
        \round_in[2][1490] , \round_in[2][1489] , \round_in[2][1488] , 
        \round_in[2][1487] , \round_in[2][1486] , \round_in[2][1485] , 
        \round_in[2][1484] , \round_in[2][1483] , \round_in[2][1482] , 
        \round_in[2][1481] , \round_in[2][1480] , \round_in[2][1479] , 
        \round_in[2][1478] , \round_in[2][1477] , \round_in[2][1476] , 
        \round_in[2][1475] , \round_in[2][1474] , \round_in[2][1473] , 
        \round_in[2][1472] , \round_in[2][1471] , \round_in[2][1470] , 
        \round_in[2][1469] , \round_in[2][1468] , \round_in[2][1467] , 
        \round_in[2][1466] , \round_in[2][1465] , \round_in[2][1464] , 
        \round_in[2][1463] , \round_in[2][1462] , \round_in[2][1461] , 
        \round_in[2][1460] , \round_in[2][1459] , \round_in[2][1458] , 
        \round_in[2][1457] , \round_in[2][1456] , \round_in[2][1455] , 
        \round_in[2][1454] , \round_in[2][1453] , \round_in[2][1452] , 
        \round_in[2][1451] , \round_in[2][1450] , \round_in[2][1449] , 
        \round_in[2][1448] , \round_in[2][1447] , \round_in[2][1446] , 
        \round_in[2][1445] , \round_in[2][1444] , \round_in[2][1443] , 
        \round_in[2][1442] , \round_in[2][1441] , \round_in[2][1440] , 
        \round_in[2][1439] , \round_in[2][1438] , \round_in[2][1437] , 
        \round_in[2][1436] , \round_in[2][1435] , \round_in[2][1434] , 
        \round_in[2][1433] , \round_in[2][1432] , \round_in[2][1431] , 
        \round_in[2][1430] , \round_in[2][1429] , \round_in[2][1428] , 
        \round_in[2][1427] , \round_in[2][1426] , \round_in[2][1425] , 
        \round_in[2][1424] , \round_in[2][1423] , \round_in[2][1422] , 
        \round_in[2][1421] , \round_in[2][1420] , \round_in[2][1419] , 
        \round_in[2][1418] , \round_in[2][1417] , \round_in[2][1416] , 
        \round_in[2][1415] , \round_in[2][1414] , \round_in[2][1413] , 
        \round_in[2][1412] , \round_in[2][1411] , \round_in[2][1410] , 
        \round_in[2][1409] , \round_in[2][1408] , \round_in[2][1407] , 
        \round_in[2][1406] , \round_in[2][1405] , \round_in[2][1404] , 
        \round_in[2][1403] , \round_in[2][1402] , \round_in[2][1401] , 
        \round_in[2][1400] , \round_in[2][1399] , \round_in[2][1398] , 
        \round_in[2][1397] , \round_in[2][1396] , \round_in[2][1395] , 
        \round_in[2][1394] , \round_in[2][1393] , \round_in[2][1392] , 
        \round_in[2][1391] , \round_in[2][1390] , \round_in[2][1389] , 
        \round_in[2][1388] , \round_in[2][1387] , \round_in[2][1386] , 
        \round_in[2][1385] , \round_in[2][1384] , \round_in[2][1383] , 
        \round_in[2][1382] , \round_in[2][1381] , \round_in[2][1380] , 
        \round_in[2][1379] , \round_in[2][1378] , \round_in[2][1377] , 
        \round_in[2][1376] , \round_in[2][1375] , \round_in[2][1374] , 
        \round_in[2][1373] , \round_in[2][1372] , \round_in[2][1371] , 
        \round_in[2][1370] , \round_in[2][1369] , \round_in[2][1368] , 
        \round_in[2][1367] , \round_in[2][1366] , \round_in[2][1365] , 
        \round_in[2][1364] , \round_in[2][1363] , \round_in[2][1362] , 
        \round_in[2][1361] , \round_in[2][1360] , \round_in[2][1359] , 
        \round_in[2][1358] , \round_in[2][1357] , \round_in[2][1356] , 
        \round_in[2][1355] , \round_in[2][1354] , \round_in[2][1353] , 
        \round_in[2][1352] , \round_in[2][1351] , \round_in[2][1350] , 
        \round_in[2][1349] , \round_in[2][1348] , \round_in[2][1347] , 
        \round_in[2][1346] , \round_in[2][1345] , \round_in[2][1344] , 
        \round_in[2][1343] , \round_in[2][1342] , \round_in[2][1341] , 
        \round_in[2][1340] , \round_in[2][1339] , \round_in[2][1338] , 
        \round_in[2][1337] , \round_in[2][1336] , \round_in[2][1335] , 
        \round_in[2][1334] , \round_in[2][1333] , \round_in[2][1332] , 
        \round_in[2][1331] , \round_in[2][1330] , \round_in[2][1329] , 
        \round_in[2][1328] , \round_in[2][1327] , \round_in[2][1326] , 
        \round_in[2][1325] , \round_in[2][1324] , \round_in[2][1323] , 
        \round_in[2][1322] , \round_in[2][1321] , \round_in[2][1320] , 
        \round_in[2][1319] , \round_in[2][1318] , \round_in[2][1317] , 
        \round_in[2][1316] , \round_in[2][1315] , \round_in[2][1314] , 
        \round_in[2][1313] , \round_in[2][1312] , \round_in[2][1311] , 
        \round_in[2][1310] , \round_in[2][1309] , \round_in[2][1308] , 
        \round_in[2][1307] , \round_in[2][1306] , \round_in[2][1305] , 
        \round_in[2][1304] , \round_in[2][1303] , \round_in[2][1302] , 
        \round_in[2][1301] , \round_in[2][1300] , \round_in[2][1299] , 
        \round_in[2][1298] , \round_in[2][1297] , \round_in[2][1296] , 
        \round_in[2][1295] , \round_in[2][1294] , \round_in[2][1293] , 
        \round_in[2][1292] , \round_in[2][1291] , \round_in[2][1290] , 
        \round_in[2][1289] , \round_in[2][1288] , \round_in[2][1287] , 
        \round_in[2][1286] , \round_in[2][1285] , \round_in[2][1284] , 
        \round_in[2][1283] , \round_in[2][1282] , \round_in[2][1281] , 
        \round_in[2][1280] , \round_in[2][1279] , \round_in[2][1278] , 
        \round_in[2][1277] , \round_in[2][1276] , \round_in[2][1275] , 
        \round_in[2][1274] , \round_in[2][1273] , \round_in[2][1272] , 
        \round_in[2][1271] , \round_in[2][1270] , \round_in[2][1269] , 
        \round_in[2][1268] , \round_in[2][1267] , \round_in[2][1266] , 
        \round_in[2][1265] , \round_in[2][1264] , \round_in[2][1263] , 
        \round_in[2][1262] , \round_in[2][1261] , \round_in[2][1260] , 
        \round_in[2][1259] , \round_in[2][1258] , \round_in[2][1257] , 
        \round_in[2][1256] , \round_in[2][1255] , \round_in[2][1254] , 
        \round_in[2][1253] , \round_in[2][1252] , \round_in[2][1251] , 
        \round_in[2][1250] , \round_in[2][1249] , \round_in[2][1248] , 
        \round_in[2][1247] , \round_in[2][1246] , \round_in[2][1245] , 
        \round_in[2][1244] , \round_in[2][1243] , \round_in[2][1242] , 
        \round_in[2][1241] , \round_in[2][1240] , \round_in[2][1239] , 
        \round_in[2][1238] , \round_in[2][1237] , \round_in[2][1236] , 
        \round_in[2][1235] , \round_in[2][1234] , \round_in[2][1233] , 
        \round_in[2][1232] , \round_in[2][1231] , \round_in[2][1230] , 
        \round_in[2][1229] , \round_in[2][1228] , \round_in[2][1227] , 
        \round_in[2][1226] , \round_in[2][1225] , \round_in[2][1224] , 
        \round_in[2][1223] , \round_in[2][1222] , \round_in[2][1221] , 
        \round_in[2][1220] , \round_in[2][1219] , \round_in[2][1218] , 
        \round_in[2][1217] , \round_in[2][1216] , \round_in[2][1215] , 
        \round_in[2][1214] , \round_in[2][1213] , \round_in[2][1212] , 
        \round_in[2][1211] , \round_in[2][1210] , \round_in[2][1209] , 
        \round_in[2][1208] , \round_in[2][1207] , \round_in[2][1206] , 
        \round_in[2][1205] , \round_in[2][1204] , \round_in[2][1203] , 
        \round_in[2][1202] , \round_in[2][1201] , \round_in[2][1200] , 
        \round_in[2][1199] , \round_in[2][1198] , \round_in[2][1197] , 
        \round_in[2][1196] , \round_in[2][1195] , \round_in[2][1194] , 
        \round_in[2][1193] , \round_in[2][1192] , \round_in[2][1191] , 
        \round_in[2][1190] , \round_in[2][1189] , \round_in[2][1188] , 
        \round_in[2][1187] , \round_in[2][1186] , \round_in[2][1185] , 
        \round_in[2][1184] , \round_in[2][1183] , \round_in[2][1182] , 
        \round_in[2][1181] , \round_in[2][1180] , \round_in[2][1179] , 
        \round_in[2][1178] , \round_in[2][1177] , \round_in[2][1176] , 
        \round_in[2][1175] , \round_in[2][1174] , \round_in[2][1173] , 
        \round_in[2][1172] , \round_in[2][1171] , \round_in[2][1170] , 
        \round_in[2][1169] , \round_in[2][1168] , \round_in[2][1167] , 
        \round_in[2][1166] , \round_in[2][1165] , \round_in[2][1164] , 
        \round_in[2][1163] , \round_in[2][1162] , \round_in[2][1161] , 
        \round_in[2][1160] , \round_in[2][1159] , \round_in[2][1158] , 
        \round_in[2][1157] , \round_in[2][1156] , \round_in[2][1155] , 
        \round_in[2][1154] , \round_in[2][1153] , \round_in[2][1152] , 
        \round_in[2][1151] , \round_in[2][1150] , \round_in[2][1149] , 
        \round_in[2][1148] , \round_in[2][1147] , \round_in[2][1146] , 
        \round_in[2][1145] , \round_in[2][1144] , \round_in[2][1143] , 
        \round_in[2][1142] , \round_in[2][1141] , \round_in[2][1140] , 
        \round_in[2][1139] , \round_in[2][1138] , \round_in[2][1137] , 
        \round_in[2][1136] , \round_in[2][1135] , \round_in[2][1134] , 
        \round_in[2][1133] , \round_in[2][1132] , \round_in[2][1131] , 
        \round_in[2][1130] , \round_in[2][1129] , \round_in[2][1128] , 
        \round_in[2][1127] , \round_in[2][1126] , \round_in[2][1125] , 
        \round_in[2][1124] , \round_in[2][1123] , \round_in[2][1122] , 
        \round_in[2][1121] , \round_in[2][1120] , \round_in[2][1119] , 
        \round_in[2][1118] , \round_in[2][1117] , \round_in[2][1116] , 
        \round_in[2][1115] , \round_in[2][1114] , \round_in[2][1113] , 
        \round_in[2][1112] , \round_in[2][1111] , \round_in[2][1110] , 
        \round_in[2][1109] , \round_in[2][1108] , \round_in[2][1107] , 
        \round_in[2][1106] , \round_in[2][1105] , \round_in[2][1104] , 
        \round_in[2][1103] , \round_in[2][1102] , \round_in[2][1101] , 
        \round_in[2][1100] , \round_in[2][1099] , \round_in[2][1098] , 
        \round_in[2][1097] , \round_in[2][1096] , \round_in[2][1095] , 
        \round_in[2][1094] , \round_in[2][1093] , \round_in[2][1092] , 
        \round_in[2][1091] , \round_in[2][1090] , \round_in[2][1089] , 
        \round_in[2][1088] , \round_in[2][1087] , \round_in[2][1086] , 
        \round_in[2][1085] , \round_in[2][1084] , \round_in[2][1083] , 
        \round_in[2][1082] , \round_in[2][1081] , \round_in[2][1080] , 
        \round_in[2][1079] , \round_in[2][1078] , \round_in[2][1077] , 
        \round_in[2][1076] , \round_in[2][1075] , \round_in[2][1074] , 
        \round_in[2][1073] , \round_in[2][1072] , \round_in[2][1071] , 
        \round_in[2][1070] , \round_in[2][1069] , \round_in[2][1068] , 
        \round_in[2][1067] , \round_in[2][1066] , \round_in[2][1065] , 
        \round_in[2][1064] , \round_in[2][1063] , \round_in[2][1062] , 
        \round_in[2][1061] , \round_in[2][1060] , \round_in[2][1059] , 
        \round_in[2][1058] , \round_in[2][1057] , \round_in[2][1056] , 
        \round_in[2][1055] , \round_in[2][1054] , \round_in[2][1053] , 
        \round_in[2][1052] , \round_in[2][1051] , \round_in[2][1050] , 
        \round_in[2][1049] , \round_in[2][1048] , \round_in[2][1047] , 
        \round_in[2][1046] , \round_in[2][1045] , \round_in[2][1044] , 
        \round_in[2][1043] , \round_in[2][1042] , \round_in[2][1041] , 
        \round_in[2][1040] , \round_in[2][1039] , \round_in[2][1038] , 
        \round_in[2][1037] , \round_in[2][1036] , \round_in[2][1035] , 
        \round_in[2][1034] , \round_in[2][1033] , \round_in[2][1032] , 
        \round_in[2][1031] , \round_in[2][1030] , \round_in[2][1029] , 
        \round_in[2][1028] , \round_in[2][1027] , \round_in[2][1026] , 
        \round_in[2][1025] , \round_in[2][1024] , \round_in[2][1023] , 
        \round_in[2][1022] , \round_in[2][1021] , \round_in[2][1020] , 
        \round_in[2][1019] , \round_in[2][1018] , \round_in[2][1017] , 
        \round_in[2][1016] , \round_in[2][1015] , \round_in[2][1014] , 
        \round_in[2][1013] , \round_in[2][1012] , \round_in[2][1011] , 
        \round_in[2][1010] , \round_in[2][1009] , \round_in[2][1008] , 
        \round_in[2][1007] , \round_in[2][1006] , \round_in[2][1005] , 
        \round_in[2][1004] , \round_in[2][1003] , \round_in[2][1002] , 
        \round_in[2][1001] , \round_in[2][1000] , \round_in[2][999] , 
        \round_in[2][998] , \round_in[2][997] , \round_in[2][996] , 
        \round_in[2][995] , \round_in[2][994] , \round_in[2][993] , 
        \round_in[2][992] , \round_in[2][991] , \round_in[2][990] , 
        \round_in[2][989] , \round_in[2][988] , \round_in[2][987] , 
        \round_in[2][986] , \round_in[2][985] , \round_in[2][984] , 
        \round_in[2][983] , \round_in[2][982] , \round_in[2][981] , 
        \round_in[2][980] , \round_in[2][979] , \round_in[2][978] , 
        \round_in[2][977] , \round_in[2][976] , \round_in[2][975] , 
        \round_in[2][974] , \round_in[2][973] , \round_in[2][972] , 
        \round_in[2][971] , \round_in[2][970] , \round_in[2][969] , 
        \round_in[2][968] , \round_in[2][967] , \round_in[2][966] , 
        \round_in[2][965] , \round_in[2][964] , \round_in[2][963] , 
        \round_in[2][962] , \round_in[2][961] , \round_in[2][960] , 
        \round_in[2][959] , \round_in[2][958] , \round_in[2][957] , 
        \round_in[2][956] , \round_in[2][955] , \round_in[2][954] , 
        \round_in[2][953] , \round_in[2][952] , \round_in[2][951] , 
        \round_in[2][950] , \round_in[2][949] , \round_in[2][948] , 
        \round_in[2][947] , \round_in[2][946] , \round_in[2][945] , 
        \round_in[2][944] , \round_in[2][943] , \round_in[2][942] , 
        \round_in[2][941] , \round_in[2][940] , \round_in[2][939] , 
        \round_in[2][938] , \round_in[2][937] , \round_in[2][936] , 
        \round_in[2][935] , \round_in[2][934] , \round_in[2][933] , 
        \round_in[2][932] , \round_in[2][931] , \round_in[2][930] , 
        \round_in[2][929] , \round_in[2][928] , \round_in[2][927] , 
        \round_in[2][926] , \round_in[2][925] , \round_in[2][924] , 
        \round_in[2][923] , \round_in[2][922] , \round_in[2][921] , 
        \round_in[2][920] , \round_in[2][919] , \round_in[2][918] , 
        \round_in[2][917] , \round_in[2][916] , \round_in[2][915] , 
        \round_in[2][914] , \round_in[2][913] , \round_in[2][912] , 
        \round_in[2][911] , \round_in[2][910] , \round_in[2][909] , 
        \round_in[2][908] , \round_in[2][907] , \round_in[2][906] , 
        \round_in[2][905] , \round_in[2][904] , \round_in[2][903] , 
        \round_in[2][902] , \round_in[2][901] , \round_in[2][900] , 
        \round_in[2][899] , \round_in[2][898] , \round_in[2][897] , 
        \round_in[2][896] , \round_in[2][895] , \round_in[2][894] , 
        \round_in[2][893] , \round_in[2][892] , \round_in[2][891] , 
        \round_in[2][890] , \round_in[2][889] , \round_in[2][888] , 
        \round_in[2][887] , \round_in[2][886] , \round_in[2][885] , 
        \round_in[2][884] , \round_in[2][883] , \round_in[2][882] , 
        \round_in[2][881] , \round_in[2][880] , \round_in[2][879] , 
        \round_in[2][878] , \round_in[2][877] , \round_in[2][876] , 
        \round_in[2][875] , \round_in[2][874] , \round_in[2][873] , 
        \round_in[2][872] , \round_in[2][871] , \round_in[2][870] , 
        \round_in[2][869] , \round_in[2][868] , \round_in[2][867] , 
        \round_in[2][866] , \round_in[2][865] , \round_in[2][864] , 
        \round_in[2][863] , \round_in[2][862] , \round_in[2][861] , 
        \round_in[2][860] , \round_in[2][859] , \round_in[2][858] , 
        \round_in[2][857] , \round_in[2][856] , \round_in[2][855] , 
        \round_in[2][854] , \round_in[2][853] , \round_in[2][852] , 
        \round_in[2][851] , \round_in[2][850] , \round_in[2][849] , 
        \round_in[2][848] , \round_in[2][847] , \round_in[2][846] , 
        \round_in[2][845] , \round_in[2][844] , \round_in[2][843] , 
        \round_in[2][842] , \round_in[2][841] , \round_in[2][840] , 
        \round_in[2][839] , \round_in[2][838] , \round_in[2][837] , 
        \round_in[2][836] , \round_in[2][835] , \round_in[2][834] , 
        \round_in[2][833] , \round_in[2][832] , \round_in[2][831] , 
        \round_in[2][830] , \round_in[2][829] , \round_in[2][828] , 
        \round_in[2][827] , \round_in[2][826] , \round_in[2][825] , 
        \round_in[2][824] , \round_in[2][823] , \round_in[2][822] , 
        \round_in[2][821] , \round_in[2][820] , \round_in[2][819] , 
        \round_in[2][818] , \round_in[2][817] , \round_in[2][816] , 
        \round_in[2][815] , \round_in[2][814] , \round_in[2][813] , 
        \round_in[2][812] , \round_in[2][811] , \round_in[2][810] , 
        \round_in[2][809] , \round_in[2][808] , \round_in[2][807] , 
        \round_in[2][806] , \round_in[2][805] , \round_in[2][804] , 
        \round_in[2][803] , \round_in[2][802] , \round_in[2][801] , 
        \round_in[2][800] , \round_in[2][799] , \round_in[2][798] , 
        \round_in[2][797] , \round_in[2][796] , \round_in[2][795] , 
        \round_in[2][794] , \round_in[2][793] , \round_in[2][792] , 
        \round_in[2][791] , \round_in[2][790] , \round_in[2][789] , 
        \round_in[2][788] , \round_in[2][787] , \round_in[2][786] , 
        \round_in[2][785] , \round_in[2][784] , \round_in[2][783] , 
        \round_in[2][782] , \round_in[2][781] , \round_in[2][780] , 
        \round_in[2][779] , \round_in[2][778] , \round_in[2][777] , 
        \round_in[2][776] , \round_in[2][775] , \round_in[2][774] , 
        \round_in[2][773] , \round_in[2][772] , \round_in[2][771] , 
        \round_in[2][770] , \round_in[2][769] , \round_in[2][768] , 
        \round_in[2][767] , \round_in[2][766] , \round_in[2][765] , 
        \round_in[2][764] , \round_in[2][763] , \round_in[2][762] , 
        \round_in[2][761] , \round_in[2][760] , \round_in[2][759] , 
        \round_in[2][758] , \round_in[2][757] , \round_in[2][756] , 
        \round_in[2][755] , \round_in[2][754] , \round_in[2][753] , 
        \round_in[2][752] , \round_in[2][751] , \round_in[2][750] , 
        \round_in[2][749] , \round_in[2][748] , \round_in[2][747] , 
        \round_in[2][746] , \round_in[2][745] , \round_in[2][744] , 
        \round_in[2][743] , \round_in[2][742] , \round_in[2][741] , 
        \round_in[2][740] , \round_in[2][739] , \round_in[2][738] , 
        \round_in[2][737] , \round_in[2][736] , \round_in[2][735] , 
        \round_in[2][734] , \round_in[2][733] , \round_in[2][732] , 
        \round_in[2][731] , \round_in[2][730] , \round_in[2][729] , 
        \round_in[2][728] , \round_in[2][727] , \round_in[2][726] , 
        \round_in[2][725] , \round_in[2][724] , \round_in[2][723] , 
        \round_in[2][722] , \round_in[2][721] , \round_in[2][720] , 
        \round_in[2][719] , \round_in[2][718] , \round_in[2][717] , 
        \round_in[2][716] , \round_in[2][715] , \round_in[2][714] , 
        \round_in[2][713] , \round_in[2][712] , \round_in[2][711] , 
        \round_in[2][710] , \round_in[2][709] , \round_in[2][708] , 
        \round_in[2][707] , \round_in[2][706] , \round_in[2][705] , 
        \round_in[2][704] , \round_in[2][703] , \round_in[2][702] , 
        \round_in[2][701] , \round_in[2][700] , \round_in[2][699] , 
        \round_in[2][698] , \round_in[2][697] , \round_in[2][696] , 
        \round_in[2][695] , \round_in[2][694] , \round_in[2][693] , 
        \round_in[2][692] , \round_in[2][691] , \round_in[2][690] , 
        \round_in[2][689] , \round_in[2][688] , \round_in[2][687] , 
        \round_in[2][686] , \round_in[2][685] , \round_in[2][684] , 
        \round_in[2][683] , \round_in[2][682] , \round_in[2][681] , 
        \round_in[2][680] , \round_in[2][679] , \round_in[2][678] , 
        \round_in[2][677] , \round_in[2][676] , \round_in[2][675] , 
        \round_in[2][674] , \round_in[2][673] , \round_in[2][672] , 
        \round_in[2][671] , \round_in[2][670] , \round_in[2][669] , 
        \round_in[2][668] , \round_in[2][667] , \round_in[2][666] , 
        \round_in[2][665] , \round_in[2][664] , \round_in[2][663] , 
        \round_in[2][662] , \round_in[2][661] , \round_in[2][660] , 
        \round_in[2][659] , \round_in[2][658] , \round_in[2][657] , 
        \round_in[2][656] , \round_in[2][655] , \round_in[2][654] , 
        \round_in[2][653] , \round_in[2][652] , \round_in[2][651] , 
        \round_in[2][650] , \round_in[2][649] , \round_in[2][648] , 
        \round_in[2][647] , \round_in[2][646] , \round_in[2][645] , 
        \round_in[2][644] , \round_in[2][643] , \round_in[2][642] , 
        \round_in[2][641] , \round_in[2][640] , \round_in[2][639] , 
        \round_in[2][638] , \round_in[2][637] , \round_in[2][636] , 
        \round_in[2][635] , \round_in[2][634] , \round_in[2][633] , 
        \round_in[2][632] , \round_in[2][631] , \round_in[2][630] , 
        \round_in[2][629] , \round_in[2][628] , \round_in[2][627] , 
        \round_in[2][626] , \round_in[2][625] , \round_in[2][624] , 
        \round_in[2][623] , \round_in[2][622] , \round_in[2][621] , 
        \round_in[2][620] , \round_in[2][619] , \round_in[2][618] , 
        \round_in[2][617] , \round_in[2][616] , \round_in[2][615] , 
        \round_in[2][614] , \round_in[2][613] , \round_in[2][612] , 
        \round_in[2][611] , \round_in[2][610] , \round_in[2][609] , 
        \round_in[2][608] , \round_in[2][607] , \round_in[2][606] , 
        \round_in[2][605] , \round_in[2][604] , \round_in[2][603] , 
        \round_in[2][602] , \round_in[2][601] , \round_in[2][600] , 
        \round_in[2][599] , \round_in[2][598] , \round_in[2][597] , 
        \round_in[2][596] , \round_in[2][595] , \round_in[2][594] , 
        \round_in[2][593] , \round_in[2][592] , \round_in[2][591] , 
        \round_in[2][590] , \round_in[2][589] , \round_in[2][588] , 
        \round_in[2][587] , \round_in[2][586] , \round_in[2][585] , 
        \round_in[2][584] , \round_in[2][583] , \round_in[2][582] , 
        \round_in[2][581] , \round_in[2][580] , \round_in[2][579] , 
        \round_in[2][578] , \round_in[2][577] , \round_in[2][576] , 
        \round_in[2][575] , \round_in[2][574] , \round_in[2][573] , 
        \round_in[2][572] , \round_in[2][571] , \round_in[2][570] , 
        \round_in[2][569] , \round_in[2][568] , \round_in[2][567] , 
        \round_in[2][566] , \round_in[2][565] , \round_in[2][564] , 
        \round_in[2][563] , \round_in[2][562] , \round_in[2][561] , 
        \round_in[2][560] , \round_in[2][559] , \round_in[2][558] , 
        \round_in[2][557] , \round_in[2][556] , \round_in[2][555] , 
        \round_in[2][554] , \round_in[2][553] , \round_in[2][552] , 
        \round_in[2][551] , \round_in[2][550] , \round_in[2][549] , 
        \round_in[2][548] , \round_in[2][547] , \round_in[2][546] , 
        \round_in[2][545] , \round_in[2][544] , \round_in[2][543] , 
        \round_in[2][542] , \round_in[2][541] , \round_in[2][540] , 
        \round_in[2][539] , \round_in[2][538] , \round_in[2][537] , 
        \round_in[2][536] , \round_in[2][535] , \round_in[2][534] , 
        \round_in[2][533] , \round_in[2][532] , \round_in[2][531] , 
        \round_in[2][530] , \round_in[2][529] , \round_in[2][528] , 
        \round_in[2][527] , \round_in[2][526] , \round_in[2][525] , 
        \round_in[2][524] , \round_in[2][523] , \round_in[2][522] , 
        \round_in[2][521] , \round_in[2][520] , \round_in[2][519] , 
        \round_in[2][518] , \round_in[2][517] , \round_in[2][516] , 
        \round_in[2][515] , \round_in[2][514] , \round_in[2][513] , 
        \round_in[2][512] , \round_in[2][511] , \round_in[2][510] , 
        \round_in[2][509] , \round_in[2][508] , \round_in[2][507] , 
        \round_in[2][506] , \round_in[2][505] , \round_in[2][504] , 
        \round_in[2][503] , \round_in[2][502] , \round_in[2][501] , 
        \round_in[2][500] , \round_in[2][499] , \round_in[2][498] , 
        \round_in[2][497] , \round_in[2][496] , \round_in[2][495] , 
        \round_in[2][494] , \round_in[2][493] , \round_in[2][492] , 
        \round_in[2][491] , \round_in[2][490] , \round_in[2][489] , 
        \round_in[2][488] , \round_in[2][487] , \round_in[2][486] , 
        \round_in[2][485] , \round_in[2][484] , \round_in[2][483] , 
        \round_in[2][482] , \round_in[2][481] , \round_in[2][480] , 
        \round_in[2][479] , \round_in[2][478] , \round_in[2][477] , 
        \round_in[2][476] , \round_in[2][475] , \round_in[2][474] , 
        \round_in[2][473] , \round_in[2][472] , \round_in[2][471] , 
        \round_in[2][470] , \round_in[2][469] , \round_in[2][468] , 
        \round_in[2][467] , \round_in[2][466] , \round_in[2][465] , 
        \round_in[2][464] , \round_in[2][463] , \round_in[2][462] , 
        \round_in[2][461] , \round_in[2][460] , \round_in[2][459] , 
        \round_in[2][458] , \round_in[2][457] , \round_in[2][456] , 
        \round_in[2][455] , \round_in[2][454] , \round_in[2][453] , 
        \round_in[2][452] , \round_in[2][451] , \round_in[2][450] , 
        \round_in[2][449] , \round_in[2][448] , \round_in[2][447] , 
        \round_in[2][446] , \round_in[2][445] , \round_in[2][444] , 
        \round_in[2][443] , \round_in[2][442] , \round_in[2][441] , 
        \round_in[2][440] , \round_in[2][439] , \round_in[2][438] , 
        \round_in[2][437] , \round_in[2][436] , \round_in[2][435] , 
        \round_in[2][434] , \round_in[2][433] , \round_in[2][432] , 
        \round_in[2][431] , \round_in[2][430] , \round_in[2][429] , 
        \round_in[2][428] , \round_in[2][427] , \round_in[2][426] , 
        \round_in[2][425] , \round_in[2][424] , \round_in[2][423] , 
        \round_in[2][422] , \round_in[2][421] , \round_in[2][420] , 
        \round_in[2][419] , \round_in[2][418] , \round_in[2][417] , 
        \round_in[2][416] , \round_in[2][415] , \round_in[2][414] , 
        \round_in[2][413] , \round_in[2][412] , \round_in[2][411] , 
        \round_in[2][410] , \round_in[2][409] , \round_in[2][408] , 
        \round_in[2][407] , \round_in[2][406] , \round_in[2][405] , 
        \round_in[2][404] , \round_in[2][403] , \round_in[2][402] , 
        \round_in[2][401] , \round_in[2][400] , \round_in[2][399] , 
        \round_in[2][398] , \round_in[2][397] , \round_in[2][396] , 
        \round_in[2][395] , \round_in[2][394] , \round_in[2][393] , 
        \round_in[2][392] , \round_in[2][391] , \round_in[2][390] , 
        \round_in[2][389] , \round_in[2][388] , \round_in[2][387] , 
        \round_in[2][386] , \round_in[2][385] , \round_in[2][384] , 
        \round_in[2][383] , \round_in[2][382] , \round_in[2][381] , 
        \round_in[2][380] , \round_in[2][379] , \round_in[2][378] , 
        \round_in[2][377] , \round_in[2][376] , \round_in[2][375] , 
        \round_in[2][374] , \round_in[2][373] , \round_in[2][372] , 
        \round_in[2][371] , \round_in[2][370] , \round_in[2][369] , 
        \round_in[2][368] , \round_in[2][367] , \round_in[2][366] , 
        \round_in[2][365] , \round_in[2][364] , \round_in[2][363] , 
        \round_in[2][362] , \round_in[2][361] , \round_in[2][360] , 
        \round_in[2][359] , \round_in[2][358] , \round_in[2][357] , 
        \round_in[2][356] , \round_in[2][355] , \round_in[2][354] , 
        \round_in[2][353] , \round_in[2][352] , \round_in[2][351] , 
        \round_in[2][350] , \round_in[2][349] , \round_in[2][348] , 
        \round_in[2][347] , \round_in[2][346] , \round_in[2][345] , 
        \round_in[2][344] , \round_in[2][343] , \round_in[2][342] , 
        \round_in[2][341] , \round_in[2][340] , \round_in[2][339] , 
        \round_in[2][338] , \round_in[2][337] , \round_in[2][336] , 
        \round_in[2][335] , \round_in[2][334] , \round_in[2][333] , 
        \round_in[2][332] , \round_in[2][331] , \round_in[2][330] , 
        \round_in[2][329] , \round_in[2][328] , \round_in[2][327] , 
        \round_in[2][326] , \round_in[2][325] , \round_in[2][324] , 
        \round_in[2][323] , \round_in[2][322] , \round_in[2][321] , 
        \round_in[2][320] , \round_in[2][319] , \round_in[2][318] , 
        \round_in[2][317] , \round_in[2][316] , \round_in[2][315] , 
        \round_in[2][314] , \round_in[2][313] , \round_in[2][312] , 
        \round_in[2][311] , \round_in[2][310] , \round_in[2][309] , 
        \round_in[2][308] , \round_in[2][307] , \round_in[2][306] , 
        \round_in[2][305] , \round_in[2][304] , \round_in[2][303] , 
        \round_in[2][302] , \round_in[2][301] , \round_in[2][300] , 
        \round_in[2][299] , \round_in[2][298] , \round_in[2][297] , 
        \round_in[2][296] , \round_in[2][295] , \round_in[2][294] , 
        \round_in[2][293] , \round_in[2][292] , \round_in[2][291] , 
        \round_in[2][290] , \round_in[2][289] , \round_in[2][288] , 
        \round_in[2][287] , \round_in[2][286] , \round_in[2][285] , 
        \round_in[2][284] , \round_in[2][283] , \round_in[2][282] , 
        \round_in[2][281] , \round_in[2][280] , \round_in[2][279] , 
        \round_in[2][278] , \round_in[2][277] , \round_in[2][276] , 
        \round_in[2][275] , \round_in[2][274] , \round_in[2][273] , 
        \round_in[2][272] , \round_in[2][271] , \round_in[2][270] , 
        \round_in[2][269] , \round_in[2][268] , \round_in[2][267] , 
        \round_in[2][266] , \round_in[2][265] , \round_in[2][264] , 
        \round_in[2][263] , \round_in[2][262] , \round_in[2][261] , 
        \round_in[2][260] , \round_in[2][259] , \round_in[2][258] , 
        \round_in[2][257] , \round_in[2][256] , \round_in[2][255] , 
        \round_in[2][254] , \round_in[2][253] , \round_in[2][252] , 
        \round_in[2][251] , \round_in[2][250] , \round_in[2][249] , 
        \round_in[2][248] , \round_in[2][247] , \round_in[2][246] , 
        \round_in[2][245] , \round_in[2][244] , \round_in[2][243] , 
        \round_in[2][242] , \round_in[2][241] , \round_in[2][240] , 
        \round_in[2][239] , \round_in[2][238] , \round_in[2][237] , 
        \round_in[2][236] , \round_in[2][235] , \round_in[2][234] , 
        \round_in[2][233] , \round_in[2][232] , \round_in[2][231] , 
        \round_in[2][230] , \round_in[2][229] , \round_in[2][228] , 
        \round_in[2][227] , \round_in[2][226] , \round_in[2][225] , 
        \round_in[2][224] , \round_in[2][223] , \round_in[2][222] , 
        \round_in[2][221] , \round_in[2][220] , \round_in[2][219] , 
        \round_in[2][218] , \round_in[2][217] , \round_in[2][216] , 
        \round_in[2][215] , \round_in[2][214] , \round_in[2][213] , 
        \round_in[2][212] , \round_in[2][211] , \round_in[2][210] , 
        \round_in[2][209] , \round_in[2][208] , \round_in[2][207] , 
        \round_in[2][206] , \round_in[2][205] , \round_in[2][204] , 
        \round_in[2][203] , \round_in[2][202] , \round_in[2][201] , 
        \round_in[2][200] , \round_in[2][199] , \round_in[2][198] , 
        \round_in[2][197] , \round_in[2][196] , \round_in[2][195] , 
        \round_in[2][194] , \round_in[2][193] , \round_in[2][192] , 
        \round_in[2][191] , \round_in[2][190] , \round_in[2][189] , 
        \round_in[2][188] , \round_in[2][187] , \round_in[2][186] , 
        \round_in[2][185] , \round_in[2][184] , \round_in[2][183] , 
        \round_in[2][182] , \round_in[2][181] , \round_in[2][180] , 
        \round_in[2][179] , \round_in[2][178] , \round_in[2][177] , 
        \round_in[2][176] , \round_in[2][175] , \round_in[2][174] , 
        \round_in[2][173] , \round_in[2][172] , \round_in[2][171] , 
        \round_in[2][170] , \round_in[2][169] , \round_in[2][168] , 
        \round_in[2][167] , \round_in[2][166] , \round_in[2][165] , 
        \round_in[2][164] , \round_in[2][163] , \round_in[2][162] , 
        \round_in[2][161] , \round_in[2][160] , \round_in[2][159] , 
        \round_in[2][158] , \round_in[2][157] , \round_in[2][156] , 
        \round_in[2][155] , \round_in[2][154] , \round_in[2][153] , 
        \round_in[2][152] , \round_in[2][151] , \round_in[2][150] , 
        \round_in[2][149] , \round_in[2][148] , \round_in[2][147] , 
        \round_in[2][146] , \round_in[2][145] , \round_in[2][144] , 
        \round_in[2][143] , \round_in[2][142] , \round_in[2][141] , 
        \round_in[2][140] , \round_in[2][139] , \round_in[2][138] , 
        \round_in[2][137] , \round_in[2][136] , \round_in[2][135] , 
        \round_in[2][134] , \round_in[2][133] , \round_in[2][132] , 
        \round_in[2][131] , \round_in[2][130] , \round_in[2][129] , 
        \round_in[2][128] , \round_in[2][127] , \round_in[2][126] , 
        \round_in[2][125] , \round_in[2][124] , \round_in[2][123] , 
        \round_in[2][122] , \round_in[2][121] , \round_in[2][120] , 
        \round_in[2][119] , \round_in[2][118] , \round_in[2][117] , 
        \round_in[2][116] , \round_in[2][115] , \round_in[2][114] , 
        \round_in[2][113] , \round_in[2][112] , \round_in[2][111] , 
        \round_in[2][110] , \round_in[2][109] , \round_in[2][108] , 
        \round_in[2][107] , \round_in[2][106] , \round_in[2][105] , 
        \round_in[2][104] , \round_in[2][103] , \round_in[2][102] , 
        \round_in[2][101] , \round_in[2][100] , \round_in[2][99] , 
        \round_in[2][98] , \round_in[2][97] , \round_in[2][96] , 
        \round_in[2][95] , \round_in[2][94] , \round_in[2][93] , 
        \round_in[2][92] , \round_in[2][91] , \round_in[2][90] , 
        \round_in[2][89] , \round_in[2][88] , \round_in[2][87] , 
        \round_in[2][86] , \round_in[2][85] , \round_in[2][84] , 
        \round_in[2][83] , \round_in[2][82] , \round_in[2][81] , 
        \round_in[2][80] , \round_in[2][79] , \round_in[2][78] , 
        \round_in[2][77] , \round_in[2][76] , \round_in[2][75] , 
        \round_in[2][74] , \round_in[2][73] , \round_in[2][72] , 
        \round_in[2][71] , \round_in[2][70] , \round_in[2][69] , 
        \round_in[2][68] , \round_in[2][67] , \round_in[2][66] , 
        \round_in[2][65] , \round_in[2][64] , \round_in[2][63] , 
        \round_in[2][62] , \round_in[2][61] , \round_in[2][60] , 
        \round_in[2][59] , \round_in[2][58] , \round_in[2][57] , 
        \round_in[2][56] , \round_in[2][55] , \round_in[2][54] , 
        \round_in[2][53] , \round_in[2][52] , \round_in[2][51] , 
        \round_in[2][50] , \round_in[2][49] , \round_in[2][48] , 
        \round_in[2][47] , \round_in[2][46] , \round_in[2][45] , 
        \round_in[2][44] , \round_in[2][43] , \round_in[2][42] , 
        \round_in[2][41] , \round_in[2][40] , \round_in[2][39] , 
        \round_in[2][38] , \round_in[2][37] , \round_in[2][36] , 
        \round_in[2][35] , \round_in[2][34] , \round_in[2][33] , 
        \round_in[2][32] , \round_in[2][31] , \round_in[2][30] , 
        \round_in[2][29] , \round_in[2][28] , \round_in[2][27] , 
        \round_in[2][26] , \round_in[2][25] , \round_in[2][24] , 
        \round_in[2][23] , \round_in[2][22] , \round_in[2][21] , 
        \round_in[2][20] , \round_in[2][19] , \round_in[2][18] , 
        \round_in[2][17] , \round_in[2][16] , \round_in[2][15] , 
        \round_in[2][14] , \round_in[2][13] , \round_in[2][12] , 
        \round_in[2][11] , \round_in[2][10] , \round_in[2][9] , 
        \round_in[2][8] , \round_in[2][7] , \round_in[2][6] , \round_in[2][5] , 
        \round_in[2][4] , \round_in[2][3] , \round_in[2][2] , \round_in[2][1] , 
        \round_in[2][0] }) );
  round_4 \ROUND[2].round_  ( .in({\round_in[2][1599] , \round_in[2][1598] , 
        \round_in[2][1597] , \round_in[2][1596] , \round_in[2][1595] , 
        \round_in[2][1594] , \round_in[2][1593] , \round_in[2][1592] , 
        \round_in[2][1591] , \round_in[2][1590] , \round_in[2][1589] , 
        \round_in[2][1588] , \round_in[2][1587] , \round_in[2][1586] , 
        \round_in[2][1585] , \round_in[2][1584] , \round_in[2][1583] , 
        \round_in[2][1582] , \round_in[2][1581] , \round_in[2][1580] , 
        \round_in[2][1579] , \round_in[2][1578] , \round_in[2][1577] , 
        \round_in[2][1576] , \round_in[2][1575] , \round_in[2][1574] , 
        \round_in[2][1573] , \round_in[2][1572] , \round_in[2][1571] , 
        \round_in[2][1570] , \round_in[2][1569] , \round_in[2][1568] , 
        \round_in[2][1567] , \round_in[2][1566] , \round_in[2][1565] , 
        \round_in[2][1564] , \round_in[2][1563] , \round_in[2][1562] , 
        \round_in[2][1561] , \round_in[2][1560] , \round_in[2][1559] , 
        \round_in[2][1558] , \round_in[2][1557] , \round_in[2][1556] , 
        \round_in[2][1555] , \round_in[2][1554] , \round_in[2][1553] , 
        \round_in[2][1552] , \round_in[2][1551] , \round_in[2][1550] , 
        \round_in[2][1549] , \round_in[2][1548] , \round_in[2][1547] , 
        \round_in[2][1546] , \round_in[2][1545] , \round_in[2][1544] , 
        \round_in[2][1543] , \round_in[2][1542] , \round_in[2][1541] , 
        \round_in[2][1540] , \round_in[2][1539] , \round_in[2][1538] , 
        \round_in[2][1537] , \round_in[2][1536] , \round_in[2][1535] , 
        \round_in[2][1534] , \round_in[2][1533] , \round_in[2][1532] , 
        \round_in[2][1531] , \round_in[2][1530] , \round_in[2][1529] , 
        \round_in[2][1528] , \round_in[2][1527] , \round_in[2][1526] , 
        \round_in[2][1525] , \round_in[2][1524] , \round_in[2][1523] , 
        \round_in[2][1522] , \round_in[2][1521] , \round_in[2][1520] , 
        \round_in[2][1519] , \round_in[2][1518] , \round_in[2][1517] , 
        \round_in[2][1516] , \round_in[2][1515] , \round_in[2][1514] , 
        \round_in[2][1513] , \round_in[2][1512] , \round_in[2][1511] , 
        \round_in[2][1510] , \round_in[2][1509] , \round_in[2][1508] , 
        \round_in[2][1507] , \round_in[2][1506] , \round_in[2][1505] , 
        \round_in[2][1504] , \round_in[2][1503] , \round_in[2][1502] , 
        \round_in[2][1501] , \round_in[2][1500] , \round_in[2][1499] , 
        \round_in[2][1498] , \round_in[2][1497] , \round_in[2][1496] , 
        \round_in[2][1495] , \round_in[2][1494] , \round_in[2][1493] , 
        \round_in[2][1492] , \round_in[2][1491] , \round_in[2][1490] , 
        \round_in[2][1489] , \round_in[2][1488] , \round_in[2][1487] , 
        \round_in[2][1486] , \round_in[2][1485] , \round_in[2][1484] , 
        \round_in[2][1483] , \round_in[2][1482] , \round_in[2][1481] , 
        \round_in[2][1480] , \round_in[2][1479] , \round_in[2][1478] , 
        \round_in[2][1477] , \round_in[2][1476] , \round_in[2][1475] , 
        \round_in[2][1474] , \round_in[2][1473] , \round_in[2][1472] , 
        \round_in[2][1471] , \round_in[2][1470] , \round_in[2][1469] , 
        \round_in[2][1468] , \round_in[2][1467] , \round_in[2][1466] , 
        \round_in[2][1465] , \round_in[2][1464] , \round_in[2][1463] , 
        \round_in[2][1462] , \round_in[2][1461] , \round_in[2][1460] , 
        \round_in[2][1459] , \round_in[2][1458] , \round_in[2][1457] , 
        \round_in[2][1456] , \round_in[2][1455] , \round_in[2][1454] , 
        \round_in[2][1453] , \round_in[2][1452] , \round_in[2][1451] , 
        \round_in[2][1450] , \round_in[2][1449] , \round_in[2][1448] , 
        \round_in[2][1447] , \round_in[2][1446] , \round_in[2][1445] , 
        \round_in[2][1444] , \round_in[2][1443] , \round_in[2][1442] , 
        \round_in[2][1441] , \round_in[2][1440] , \round_in[2][1439] , 
        \round_in[2][1438] , \round_in[2][1437] , \round_in[2][1436] , 
        \round_in[2][1435] , \round_in[2][1434] , \round_in[2][1433] , 
        \round_in[2][1432] , \round_in[2][1431] , \round_in[2][1430] , 
        \round_in[2][1429] , \round_in[2][1428] , \round_in[2][1427] , 
        \round_in[2][1426] , \round_in[2][1425] , \round_in[2][1424] , 
        \round_in[2][1423] , \round_in[2][1422] , \round_in[2][1421] , 
        \round_in[2][1420] , \round_in[2][1419] , \round_in[2][1418] , 
        \round_in[2][1417] , \round_in[2][1416] , \round_in[2][1415] , 
        \round_in[2][1414] , \round_in[2][1413] , \round_in[2][1412] , 
        \round_in[2][1411] , \round_in[2][1410] , \round_in[2][1409] , 
        \round_in[2][1408] , \round_in[2][1407] , \round_in[2][1406] , 
        \round_in[2][1405] , \round_in[2][1404] , \round_in[2][1403] , 
        \round_in[2][1402] , \round_in[2][1401] , \round_in[2][1400] , 
        \round_in[2][1399] , \round_in[2][1398] , \round_in[2][1397] , 
        \round_in[2][1396] , \round_in[2][1395] , \round_in[2][1394] , 
        \round_in[2][1393] , \round_in[2][1392] , \round_in[2][1391] , 
        \round_in[2][1390] , \round_in[2][1389] , \round_in[2][1388] , 
        \round_in[2][1387] , \round_in[2][1386] , \round_in[2][1385] , 
        \round_in[2][1384] , \round_in[2][1383] , \round_in[2][1382] , 
        \round_in[2][1381] , \round_in[2][1380] , \round_in[2][1379] , 
        \round_in[2][1378] , \round_in[2][1377] , \round_in[2][1376] , 
        \round_in[2][1375] , \round_in[2][1374] , \round_in[2][1373] , 
        \round_in[2][1372] , \round_in[2][1371] , \round_in[2][1370] , 
        \round_in[2][1369] , \round_in[2][1368] , \round_in[2][1367] , 
        \round_in[2][1366] , \round_in[2][1365] , \round_in[2][1364] , 
        \round_in[2][1363] , \round_in[2][1362] , \round_in[2][1361] , 
        \round_in[2][1360] , \round_in[2][1359] , \round_in[2][1358] , 
        \round_in[2][1357] , \round_in[2][1356] , \round_in[2][1355] , 
        \round_in[2][1354] , \round_in[2][1353] , \round_in[2][1352] , 
        \round_in[2][1351] , \round_in[2][1350] , \round_in[2][1349] , 
        \round_in[2][1348] , \round_in[2][1347] , \round_in[2][1346] , 
        \round_in[2][1345] , \round_in[2][1344] , \round_in[2][1343] , 
        \round_in[2][1342] , \round_in[2][1341] , \round_in[2][1340] , 
        \round_in[2][1339] , \round_in[2][1338] , \round_in[2][1337] , 
        \round_in[2][1336] , \round_in[2][1335] , \round_in[2][1334] , 
        \round_in[2][1333] , \round_in[2][1332] , \round_in[2][1331] , 
        \round_in[2][1330] , \round_in[2][1329] , \round_in[2][1328] , 
        \round_in[2][1327] , \round_in[2][1326] , \round_in[2][1325] , 
        \round_in[2][1324] , \round_in[2][1323] , \round_in[2][1322] , 
        \round_in[2][1321] , \round_in[2][1320] , \round_in[2][1319] , 
        \round_in[2][1318] , \round_in[2][1317] , \round_in[2][1316] , 
        \round_in[2][1315] , \round_in[2][1314] , \round_in[2][1313] , 
        \round_in[2][1312] , \round_in[2][1311] , \round_in[2][1310] , 
        \round_in[2][1309] , \round_in[2][1308] , \round_in[2][1307] , 
        \round_in[2][1306] , \round_in[2][1305] , \round_in[2][1304] , 
        \round_in[2][1303] , \round_in[2][1302] , \round_in[2][1301] , 
        \round_in[2][1300] , \round_in[2][1299] , \round_in[2][1298] , 
        \round_in[2][1297] , \round_in[2][1296] , \round_in[2][1295] , 
        \round_in[2][1294] , \round_in[2][1293] , \round_in[2][1292] , 
        \round_in[2][1291] , \round_in[2][1290] , \round_in[2][1289] , 
        \round_in[2][1288] , \round_in[2][1287] , \round_in[2][1286] , 
        \round_in[2][1285] , \round_in[2][1284] , \round_in[2][1283] , 
        \round_in[2][1282] , \round_in[2][1281] , \round_in[2][1280] , 
        \round_in[2][1279] , \round_in[2][1278] , \round_in[2][1277] , 
        \round_in[2][1276] , \round_in[2][1275] , \round_in[2][1274] , 
        \round_in[2][1273] , \round_in[2][1272] , \round_in[2][1271] , 
        \round_in[2][1270] , \round_in[2][1269] , \round_in[2][1268] , 
        \round_in[2][1267] , \round_in[2][1266] , \round_in[2][1265] , 
        \round_in[2][1264] , \round_in[2][1263] , \round_in[2][1262] , 
        \round_in[2][1261] , \round_in[2][1260] , \round_in[2][1259] , 
        \round_in[2][1258] , \round_in[2][1257] , \round_in[2][1256] , 
        \round_in[2][1255] , \round_in[2][1254] , \round_in[2][1253] , 
        \round_in[2][1252] , \round_in[2][1251] , \round_in[2][1250] , 
        \round_in[2][1249] , \round_in[2][1248] , \round_in[2][1247] , 
        \round_in[2][1246] , \round_in[2][1245] , \round_in[2][1244] , 
        \round_in[2][1243] , \round_in[2][1242] , \round_in[2][1241] , 
        \round_in[2][1240] , \round_in[2][1239] , \round_in[2][1238] , 
        \round_in[2][1237] , \round_in[2][1236] , \round_in[2][1235] , 
        \round_in[2][1234] , \round_in[2][1233] , \round_in[2][1232] , 
        \round_in[2][1231] , \round_in[2][1230] , \round_in[2][1229] , 
        \round_in[2][1228] , \round_in[2][1227] , \round_in[2][1226] , 
        \round_in[2][1225] , \round_in[2][1224] , \round_in[2][1223] , 
        \round_in[2][1222] , \round_in[2][1221] , \round_in[2][1220] , 
        \round_in[2][1219] , \round_in[2][1218] , \round_in[2][1217] , 
        \round_in[2][1216] , \round_in[2][1215] , \round_in[2][1214] , 
        \round_in[2][1213] , \round_in[2][1212] , \round_in[2][1211] , 
        \round_in[2][1210] , \round_in[2][1209] , \round_in[2][1208] , 
        \round_in[2][1207] , \round_in[2][1206] , \round_in[2][1205] , 
        \round_in[2][1204] , \round_in[2][1203] , \round_in[2][1202] , 
        \round_in[2][1201] , \round_in[2][1200] , \round_in[2][1199] , 
        \round_in[2][1198] , \round_in[2][1197] , \round_in[2][1196] , 
        \round_in[2][1195] , \round_in[2][1194] , \round_in[2][1193] , 
        \round_in[2][1192] , \round_in[2][1191] , \round_in[2][1190] , 
        \round_in[2][1189] , \round_in[2][1188] , \round_in[2][1187] , 
        \round_in[2][1186] , \round_in[2][1185] , \round_in[2][1184] , 
        \round_in[2][1183] , \round_in[2][1182] , \round_in[2][1181] , 
        \round_in[2][1180] , \round_in[2][1179] , \round_in[2][1178] , 
        \round_in[2][1177] , \round_in[2][1176] , \round_in[2][1175] , 
        \round_in[2][1174] , \round_in[2][1173] , \round_in[2][1172] , 
        \round_in[2][1171] , \round_in[2][1170] , \round_in[2][1169] , 
        \round_in[2][1168] , \round_in[2][1167] , \round_in[2][1166] , 
        \round_in[2][1165] , \round_in[2][1164] , \round_in[2][1163] , 
        \round_in[2][1162] , \round_in[2][1161] , \round_in[2][1160] , 
        \round_in[2][1159] , \round_in[2][1158] , \round_in[2][1157] , 
        \round_in[2][1156] , \round_in[2][1155] , \round_in[2][1154] , 
        \round_in[2][1153] , \round_in[2][1152] , \round_in[2][1151] , 
        \round_in[2][1150] , \round_in[2][1149] , \round_in[2][1148] , 
        \round_in[2][1147] , \round_in[2][1146] , \round_in[2][1145] , 
        \round_in[2][1144] , \round_in[2][1143] , \round_in[2][1142] , 
        \round_in[2][1141] , \round_in[2][1140] , \round_in[2][1139] , 
        \round_in[2][1138] , \round_in[2][1137] , \round_in[2][1136] , 
        \round_in[2][1135] , \round_in[2][1134] , \round_in[2][1133] , 
        \round_in[2][1132] , \round_in[2][1131] , \round_in[2][1130] , 
        \round_in[2][1129] , \round_in[2][1128] , \round_in[2][1127] , 
        \round_in[2][1126] , \round_in[2][1125] , \round_in[2][1124] , 
        \round_in[2][1123] , \round_in[2][1122] , \round_in[2][1121] , 
        \round_in[2][1120] , \round_in[2][1119] , \round_in[2][1118] , 
        \round_in[2][1117] , \round_in[2][1116] , \round_in[2][1115] , 
        \round_in[2][1114] , \round_in[2][1113] , \round_in[2][1112] , 
        \round_in[2][1111] , \round_in[2][1110] , \round_in[2][1109] , 
        \round_in[2][1108] , \round_in[2][1107] , \round_in[2][1106] , 
        \round_in[2][1105] , \round_in[2][1104] , \round_in[2][1103] , 
        \round_in[2][1102] , \round_in[2][1101] , \round_in[2][1100] , 
        \round_in[2][1099] , \round_in[2][1098] , \round_in[2][1097] , 
        \round_in[2][1096] , \round_in[2][1095] , \round_in[2][1094] , 
        \round_in[2][1093] , \round_in[2][1092] , \round_in[2][1091] , 
        \round_in[2][1090] , \round_in[2][1089] , \round_in[2][1088] , 
        \round_in[2][1087] , \round_in[2][1086] , \round_in[2][1085] , 
        \round_in[2][1084] , \round_in[2][1083] , \round_in[2][1082] , 
        \round_in[2][1081] , \round_in[2][1080] , \round_in[2][1079] , 
        \round_in[2][1078] , \round_in[2][1077] , \round_in[2][1076] , 
        \round_in[2][1075] , \round_in[2][1074] , \round_in[2][1073] , 
        \round_in[2][1072] , \round_in[2][1071] , \round_in[2][1070] , 
        \round_in[2][1069] , \round_in[2][1068] , \round_in[2][1067] , 
        \round_in[2][1066] , \round_in[2][1065] , \round_in[2][1064] , 
        \round_in[2][1063] , \round_in[2][1062] , \round_in[2][1061] , 
        \round_in[2][1060] , \round_in[2][1059] , \round_in[2][1058] , 
        \round_in[2][1057] , \round_in[2][1056] , \round_in[2][1055] , 
        \round_in[2][1054] , \round_in[2][1053] , \round_in[2][1052] , 
        \round_in[2][1051] , \round_in[2][1050] , \round_in[2][1049] , 
        \round_in[2][1048] , \round_in[2][1047] , \round_in[2][1046] , 
        \round_in[2][1045] , \round_in[2][1044] , \round_in[2][1043] , 
        \round_in[2][1042] , \round_in[2][1041] , \round_in[2][1040] , 
        \round_in[2][1039] , \round_in[2][1038] , \round_in[2][1037] , 
        \round_in[2][1036] , \round_in[2][1035] , \round_in[2][1034] , 
        \round_in[2][1033] , \round_in[2][1032] , \round_in[2][1031] , 
        \round_in[2][1030] , \round_in[2][1029] , \round_in[2][1028] , 
        \round_in[2][1027] , \round_in[2][1026] , \round_in[2][1025] , 
        \round_in[2][1024] , \round_in[2][1023] , \round_in[2][1022] , 
        \round_in[2][1021] , \round_in[2][1020] , \round_in[2][1019] , 
        \round_in[2][1018] , \round_in[2][1017] , \round_in[2][1016] , 
        \round_in[2][1015] , \round_in[2][1014] , \round_in[2][1013] , 
        \round_in[2][1012] , \round_in[2][1011] , \round_in[2][1010] , 
        \round_in[2][1009] , \round_in[2][1008] , \round_in[2][1007] , 
        \round_in[2][1006] , \round_in[2][1005] , \round_in[2][1004] , 
        \round_in[2][1003] , \round_in[2][1002] , \round_in[2][1001] , 
        \round_in[2][1000] , \round_in[2][999] , \round_in[2][998] , 
        \round_in[2][997] , \round_in[2][996] , \round_in[2][995] , 
        \round_in[2][994] , \round_in[2][993] , \round_in[2][992] , 
        \round_in[2][991] , \round_in[2][990] , \round_in[2][989] , 
        \round_in[2][988] , \round_in[2][987] , \round_in[2][986] , 
        \round_in[2][985] , \round_in[2][984] , \round_in[2][983] , 
        \round_in[2][982] , \round_in[2][981] , \round_in[2][980] , 
        \round_in[2][979] , \round_in[2][978] , \round_in[2][977] , 
        \round_in[2][976] , \round_in[2][975] , \round_in[2][974] , 
        \round_in[2][973] , \round_in[2][972] , \round_in[2][971] , 
        \round_in[2][970] , \round_in[2][969] , \round_in[2][968] , 
        \round_in[2][967] , \round_in[2][966] , \round_in[2][965] , 
        \round_in[2][964] , \round_in[2][963] , \round_in[2][962] , 
        \round_in[2][961] , \round_in[2][960] , \round_in[2][959] , 
        \round_in[2][958] , \round_in[2][957] , \round_in[2][956] , 
        \round_in[2][955] , \round_in[2][954] , \round_in[2][953] , 
        \round_in[2][952] , \round_in[2][951] , \round_in[2][950] , 
        \round_in[2][949] , \round_in[2][948] , \round_in[2][947] , 
        \round_in[2][946] , \round_in[2][945] , \round_in[2][944] , 
        \round_in[2][943] , \round_in[2][942] , \round_in[2][941] , 
        \round_in[2][940] , \round_in[2][939] , \round_in[2][938] , 
        \round_in[2][937] , \round_in[2][936] , \round_in[2][935] , 
        \round_in[2][934] , \round_in[2][933] , \round_in[2][932] , 
        \round_in[2][931] , \round_in[2][930] , \round_in[2][929] , 
        \round_in[2][928] , \round_in[2][927] , \round_in[2][926] , 
        \round_in[2][925] , \round_in[2][924] , \round_in[2][923] , 
        \round_in[2][922] , \round_in[2][921] , \round_in[2][920] , 
        \round_in[2][919] , \round_in[2][918] , \round_in[2][917] , 
        \round_in[2][916] , \round_in[2][915] , \round_in[2][914] , 
        \round_in[2][913] , \round_in[2][912] , \round_in[2][911] , 
        \round_in[2][910] , \round_in[2][909] , \round_in[2][908] , 
        \round_in[2][907] , \round_in[2][906] , \round_in[2][905] , 
        \round_in[2][904] , \round_in[2][903] , \round_in[2][902] , 
        \round_in[2][901] , \round_in[2][900] , \round_in[2][899] , 
        \round_in[2][898] , \round_in[2][897] , \round_in[2][896] , 
        \round_in[2][895] , \round_in[2][894] , \round_in[2][893] , 
        \round_in[2][892] , \round_in[2][891] , \round_in[2][890] , 
        \round_in[2][889] , \round_in[2][888] , \round_in[2][887] , 
        \round_in[2][886] , \round_in[2][885] , \round_in[2][884] , 
        \round_in[2][883] , \round_in[2][882] , \round_in[2][881] , 
        \round_in[2][880] , \round_in[2][879] , \round_in[2][878] , 
        \round_in[2][877] , \round_in[2][876] , \round_in[2][875] , 
        \round_in[2][874] , \round_in[2][873] , \round_in[2][872] , 
        \round_in[2][871] , \round_in[2][870] , \round_in[2][869] , 
        \round_in[2][868] , \round_in[2][867] , \round_in[2][866] , 
        \round_in[2][865] , \round_in[2][864] , \round_in[2][863] , 
        \round_in[2][862] , \round_in[2][861] , \round_in[2][860] , 
        \round_in[2][859] , \round_in[2][858] , \round_in[2][857] , 
        \round_in[2][856] , \round_in[2][855] , \round_in[2][854] , 
        \round_in[2][853] , \round_in[2][852] , \round_in[2][851] , 
        \round_in[2][850] , \round_in[2][849] , \round_in[2][848] , 
        \round_in[2][847] , \round_in[2][846] , \round_in[2][845] , 
        \round_in[2][844] , \round_in[2][843] , \round_in[2][842] , 
        \round_in[2][841] , \round_in[2][840] , \round_in[2][839] , 
        \round_in[2][838] , \round_in[2][837] , \round_in[2][836] , 
        \round_in[2][835] , \round_in[2][834] , \round_in[2][833] , 
        \round_in[2][832] , \round_in[2][831] , \round_in[2][830] , 
        \round_in[2][829] , \round_in[2][828] , \round_in[2][827] , 
        \round_in[2][826] , \round_in[2][825] , \round_in[2][824] , 
        \round_in[2][823] , \round_in[2][822] , \round_in[2][821] , 
        \round_in[2][820] , \round_in[2][819] , \round_in[2][818] , 
        \round_in[2][817] , \round_in[2][816] , \round_in[2][815] , 
        \round_in[2][814] , \round_in[2][813] , \round_in[2][812] , 
        \round_in[2][811] , \round_in[2][810] , \round_in[2][809] , 
        \round_in[2][808] , \round_in[2][807] , \round_in[2][806] , 
        \round_in[2][805] , \round_in[2][804] , \round_in[2][803] , 
        \round_in[2][802] , \round_in[2][801] , \round_in[2][800] , 
        \round_in[2][799] , \round_in[2][798] , \round_in[2][797] , 
        \round_in[2][796] , \round_in[2][795] , \round_in[2][794] , 
        \round_in[2][793] , \round_in[2][792] , \round_in[2][791] , 
        \round_in[2][790] , \round_in[2][789] , \round_in[2][788] , 
        \round_in[2][787] , \round_in[2][786] , \round_in[2][785] , 
        \round_in[2][784] , \round_in[2][783] , \round_in[2][782] , 
        \round_in[2][781] , \round_in[2][780] , \round_in[2][779] , 
        \round_in[2][778] , \round_in[2][777] , \round_in[2][776] , 
        \round_in[2][775] , \round_in[2][774] , \round_in[2][773] , 
        \round_in[2][772] , \round_in[2][771] , \round_in[2][770] , 
        \round_in[2][769] , \round_in[2][768] , \round_in[2][767] , 
        \round_in[2][766] , \round_in[2][765] , \round_in[2][764] , 
        \round_in[2][763] , \round_in[2][762] , \round_in[2][761] , 
        \round_in[2][760] , \round_in[2][759] , \round_in[2][758] , 
        \round_in[2][757] , \round_in[2][756] , \round_in[2][755] , 
        \round_in[2][754] , \round_in[2][753] , \round_in[2][752] , 
        \round_in[2][751] , \round_in[2][750] , \round_in[2][749] , 
        \round_in[2][748] , \round_in[2][747] , \round_in[2][746] , 
        \round_in[2][745] , \round_in[2][744] , \round_in[2][743] , 
        \round_in[2][742] , \round_in[2][741] , \round_in[2][740] , 
        \round_in[2][739] , \round_in[2][738] , \round_in[2][737] , 
        \round_in[2][736] , \round_in[2][735] , \round_in[2][734] , 
        \round_in[2][733] , \round_in[2][732] , \round_in[2][731] , 
        \round_in[2][730] , \round_in[2][729] , \round_in[2][728] , 
        \round_in[2][727] , \round_in[2][726] , \round_in[2][725] , 
        \round_in[2][724] , \round_in[2][723] , \round_in[2][722] , 
        \round_in[2][721] , \round_in[2][720] , \round_in[2][719] , 
        \round_in[2][718] , \round_in[2][717] , \round_in[2][716] , 
        \round_in[2][715] , \round_in[2][714] , \round_in[2][713] , 
        \round_in[2][712] , \round_in[2][711] , \round_in[2][710] , 
        \round_in[2][709] , \round_in[2][708] , \round_in[2][707] , 
        \round_in[2][706] , \round_in[2][705] , \round_in[2][704] , 
        \round_in[2][703] , \round_in[2][702] , \round_in[2][701] , 
        \round_in[2][700] , \round_in[2][699] , \round_in[2][698] , 
        \round_in[2][697] , \round_in[2][696] , \round_in[2][695] , 
        \round_in[2][694] , \round_in[2][693] , \round_in[2][692] , 
        \round_in[2][691] , \round_in[2][690] , \round_in[2][689] , 
        \round_in[2][688] , \round_in[2][687] , \round_in[2][686] , 
        \round_in[2][685] , \round_in[2][684] , \round_in[2][683] , 
        \round_in[2][682] , \round_in[2][681] , \round_in[2][680] , 
        \round_in[2][679] , \round_in[2][678] , \round_in[2][677] , 
        \round_in[2][676] , \round_in[2][675] , \round_in[2][674] , 
        \round_in[2][673] , \round_in[2][672] , \round_in[2][671] , 
        \round_in[2][670] , \round_in[2][669] , \round_in[2][668] , 
        \round_in[2][667] , \round_in[2][666] , \round_in[2][665] , 
        \round_in[2][664] , \round_in[2][663] , \round_in[2][662] , 
        \round_in[2][661] , \round_in[2][660] , \round_in[2][659] , 
        \round_in[2][658] , \round_in[2][657] , \round_in[2][656] , 
        \round_in[2][655] , \round_in[2][654] , \round_in[2][653] , 
        \round_in[2][652] , \round_in[2][651] , \round_in[2][650] , 
        \round_in[2][649] , \round_in[2][648] , \round_in[2][647] , 
        \round_in[2][646] , \round_in[2][645] , \round_in[2][644] , 
        \round_in[2][643] , \round_in[2][642] , \round_in[2][641] , 
        \round_in[2][640] , \round_in[2][639] , \round_in[2][638] , 
        \round_in[2][637] , \round_in[2][636] , \round_in[2][635] , 
        \round_in[2][634] , \round_in[2][633] , \round_in[2][632] , 
        \round_in[2][631] , \round_in[2][630] , \round_in[2][629] , 
        \round_in[2][628] , \round_in[2][627] , \round_in[2][626] , 
        \round_in[2][625] , \round_in[2][624] , \round_in[2][623] , 
        \round_in[2][622] , \round_in[2][621] , \round_in[2][620] , 
        \round_in[2][619] , \round_in[2][618] , \round_in[2][617] , 
        \round_in[2][616] , \round_in[2][615] , \round_in[2][614] , 
        \round_in[2][613] , \round_in[2][612] , \round_in[2][611] , 
        \round_in[2][610] , \round_in[2][609] , \round_in[2][608] , 
        \round_in[2][607] , \round_in[2][606] , \round_in[2][605] , 
        \round_in[2][604] , \round_in[2][603] , \round_in[2][602] , 
        \round_in[2][601] , \round_in[2][600] , \round_in[2][599] , 
        \round_in[2][598] , \round_in[2][597] , \round_in[2][596] , 
        \round_in[2][595] , \round_in[2][594] , \round_in[2][593] , 
        \round_in[2][592] , \round_in[2][591] , \round_in[2][590] , 
        \round_in[2][589] , \round_in[2][588] , \round_in[2][587] , 
        \round_in[2][586] , \round_in[2][585] , \round_in[2][584] , 
        \round_in[2][583] , \round_in[2][582] , \round_in[2][581] , 
        \round_in[2][580] , \round_in[2][579] , \round_in[2][578] , 
        \round_in[2][577] , \round_in[2][576] , \round_in[2][575] , 
        \round_in[2][574] , \round_in[2][573] , \round_in[2][572] , 
        \round_in[2][571] , \round_in[2][570] , \round_in[2][569] , 
        \round_in[2][568] , \round_in[2][567] , \round_in[2][566] , 
        \round_in[2][565] , \round_in[2][564] , \round_in[2][563] , 
        \round_in[2][562] , \round_in[2][561] , \round_in[2][560] , 
        \round_in[2][559] , \round_in[2][558] , \round_in[2][557] , 
        \round_in[2][556] , \round_in[2][555] , \round_in[2][554] , 
        \round_in[2][553] , \round_in[2][552] , \round_in[2][551] , 
        \round_in[2][550] , \round_in[2][549] , \round_in[2][548] , 
        \round_in[2][547] , \round_in[2][546] , \round_in[2][545] , 
        \round_in[2][544] , \round_in[2][543] , \round_in[2][542] , 
        \round_in[2][541] , \round_in[2][540] , \round_in[2][539] , 
        \round_in[2][538] , \round_in[2][537] , \round_in[2][536] , 
        \round_in[2][535] , \round_in[2][534] , \round_in[2][533] , 
        \round_in[2][532] , \round_in[2][531] , \round_in[2][530] , 
        \round_in[2][529] , \round_in[2][528] , \round_in[2][527] , 
        \round_in[2][526] , \round_in[2][525] , \round_in[2][524] , 
        \round_in[2][523] , \round_in[2][522] , \round_in[2][521] , 
        \round_in[2][520] , \round_in[2][519] , \round_in[2][518] , 
        \round_in[2][517] , \round_in[2][516] , \round_in[2][515] , 
        \round_in[2][514] , \round_in[2][513] , \round_in[2][512] , 
        \round_in[2][511] , \round_in[2][510] , \round_in[2][509] , 
        \round_in[2][508] , \round_in[2][507] , \round_in[2][506] , 
        \round_in[2][505] , \round_in[2][504] , \round_in[2][503] , 
        \round_in[2][502] , \round_in[2][501] , \round_in[2][500] , 
        \round_in[2][499] , \round_in[2][498] , \round_in[2][497] , 
        \round_in[2][496] , \round_in[2][495] , \round_in[2][494] , 
        \round_in[2][493] , \round_in[2][492] , \round_in[2][491] , 
        \round_in[2][490] , \round_in[2][489] , \round_in[2][488] , 
        \round_in[2][487] , \round_in[2][486] , \round_in[2][485] , 
        \round_in[2][484] , \round_in[2][483] , \round_in[2][482] , 
        \round_in[2][481] , \round_in[2][480] , \round_in[2][479] , 
        \round_in[2][478] , \round_in[2][477] , \round_in[2][476] , 
        \round_in[2][475] , \round_in[2][474] , \round_in[2][473] , 
        \round_in[2][472] , \round_in[2][471] , \round_in[2][470] , 
        \round_in[2][469] , \round_in[2][468] , \round_in[2][467] , 
        \round_in[2][466] , \round_in[2][465] , \round_in[2][464] , 
        \round_in[2][463] , \round_in[2][462] , \round_in[2][461] , 
        \round_in[2][460] , \round_in[2][459] , \round_in[2][458] , 
        \round_in[2][457] , \round_in[2][456] , \round_in[2][455] , 
        \round_in[2][454] , \round_in[2][453] , \round_in[2][452] , 
        \round_in[2][451] , \round_in[2][450] , \round_in[2][449] , 
        \round_in[2][448] , \round_in[2][447] , \round_in[2][446] , 
        \round_in[2][445] , \round_in[2][444] , \round_in[2][443] , 
        \round_in[2][442] , \round_in[2][441] , \round_in[2][440] , 
        \round_in[2][439] , \round_in[2][438] , \round_in[2][437] , 
        \round_in[2][436] , \round_in[2][435] , \round_in[2][434] , 
        \round_in[2][433] , \round_in[2][432] , \round_in[2][431] , 
        \round_in[2][430] , \round_in[2][429] , \round_in[2][428] , 
        \round_in[2][427] , \round_in[2][426] , \round_in[2][425] , 
        \round_in[2][424] , \round_in[2][423] , \round_in[2][422] , 
        \round_in[2][421] , \round_in[2][420] , \round_in[2][419] , 
        \round_in[2][418] , \round_in[2][417] , \round_in[2][416] , 
        \round_in[2][415] , \round_in[2][414] , \round_in[2][413] , 
        \round_in[2][412] , \round_in[2][411] , \round_in[2][410] , 
        \round_in[2][409] , \round_in[2][408] , \round_in[2][407] , 
        \round_in[2][406] , \round_in[2][405] , \round_in[2][404] , 
        \round_in[2][403] , \round_in[2][402] , \round_in[2][401] , 
        \round_in[2][400] , \round_in[2][399] , \round_in[2][398] , 
        \round_in[2][397] , \round_in[2][396] , \round_in[2][395] , 
        \round_in[2][394] , \round_in[2][393] , \round_in[2][392] , 
        \round_in[2][391] , \round_in[2][390] , \round_in[2][389] , 
        \round_in[2][388] , \round_in[2][387] , \round_in[2][386] , 
        \round_in[2][385] , \round_in[2][384] , \round_in[2][383] , 
        \round_in[2][382] , \round_in[2][381] , \round_in[2][380] , 
        \round_in[2][379] , \round_in[2][378] , \round_in[2][377] , 
        \round_in[2][376] , \round_in[2][375] , \round_in[2][374] , 
        \round_in[2][373] , \round_in[2][372] , \round_in[2][371] , 
        \round_in[2][370] , \round_in[2][369] , \round_in[2][368] , 
        \round_in[2][367] , \round_in[2][366] , \round_in[2][365] , 
        \round_in[2][364] , \round_in[2][363] , \round_in[2][362] , 
        \round_in[2][361] , \round_in[2][360] , \round_in[2][359] , 
        \round_in[2][358] , \round_in[2][357] , \round_in[2][356] , 
        \round_in[2][355] , \round_in[2][354] , \round_in[2][353] , 
        \round_in[2][352] , \round_in[2][351] , \round_in[2][350] , 
        \round_in[2][349] , \round_in[2][348] , \round_in[2][347] , 
        \round_in[2][346] , \round_in[2][345] , \round_in[2][344] , 
        \round_in[2][343] , \round_in[2][342] , \round_in[2][341] , 
        \round_in[2][340] , \round_in[2][339] , \round_in[2][338] , 
        \round_in[2][337] , \round_in[2][336] , \round_in[2][335] , 
        \round_in[2][334] , \round_in[2][333] , \round_in[2][332] , 
        \round_in[2][331] , \round_in[2][330] , \round_in[2][329] , 
        \round_in[2][328] , \round_in[2][327] , \round_in[2][326] , 
        \round_in[2][325] , \round_in[2][324] , \round_in[2][323] , 
        \round_in[2][322] , \round_in[2][321] , \round_in[2][320] , 
        \round_in[2][319] , \round_in[2][318] , \round_in[2][317] , 
        \round_in[2][316] , \round_in[2][315] , \round_in[2][314] , 
        \round_in[2][313] , \round_in[2][312] , \round_in[2][311] , 
        \round_in[2][310] , \round_in[2][309] , \round_in[2][308] , 
        \round_in[2][307] , \round_in[2][306] , \round_in[2][305] , 
        \round_in[2][304] , \round_in[2][303] , \round_in[2][302] , 
        \round_in[2][301] , \round_in[2][300] , \round_in[2][299] , 
        \round_in[2][298] , \round_in[2][297] , \round_in[2][296] , 
        \round_in[2][295] , \round_in[2][294] , \round_in[2][293] , 
        \round_in[2][292] , \round_in[2][291] , \round_in[2][290] , 
        \round_in[2][289] , \round_in[2][288] , \round_in[2][287] , 
        \round_in[2][286] , \round_in[2][285] , \round_in[2][284] , 
        \round_in[2][283] , \round_in[2][282] , \round_in[2][281] , 
        \round_in[2][280] , \round_in[2][279] , \round_in[2][278] , 
        \round_in[2][277] , \round_in[2][276] , \round_in[2][275] , 
        \round_in[2][274] , \round_in[2][273] , \round_in[2][272] , 
        \round_in[2][271] , \round_in[2][270] , \round_in[2][269] , 
        \round_in[2][268] , \round_in[2][267] , \round_in[2][266] , 
        \round_in[2][265] , \round_in[2][264] , \round_in[2][263] , 
        \round_in[2][262] , \round_in[2][261] , \round_in[2][260] , 
        \round_in[2][259] , \round_in[2][258] , \round_in[2][257] , 
        \round_in[2][256] , \round_in[2][255] , \round_in[2][254] , 
        \round_in[2][253] , \round_in[2][252] , \round_in[2][251] , 
        \round_in[2][250] , \round_in[2][249] , \round_in[2][248] , 
        \round_in[2][247] , \round_in[2][246] , \round_in[2][245] , 
        \round_in[2][244] , \round_in[2][243] , \round_in[2][242] , 
        \round_in[2][241] , \round_in[2][240] , \round_in[2][239] , 
        \round_in[2][238] , \round_in[2][237] , \round_in[2][236] , 
        \round_in[2][235] , \round_in[2][234] , \round_in[2][233] , 
        \round_in[2][232] , \round_in[2][231] , \round_in[2][230] , 
        \round_in[2][229] , \round_in[2][228] , \round_in[2][227] , 
        \round_in[2][226] , \round_in[2][225] , \round_in[2][224] , 
        \round_in[2][223] , \round_in[2][222] , \round_in[2][221] , 
        \round_in[2][220] , \round_in[2][219] , \round_in[2][218] , 
        \round_in[2][217] , \round_in[2][216] , \round_in[2][215] , 
        \round_in[2][214] , \round_in[2][213] , \round_in[2][212] , 
        \round_in[2][211] , \round_in[2][210] , \round_in[2][209] , 
        \round_in[2][208] , \round_in[2][207] , \round_in[2][206] , 
        \round_in[2][205] , \round_in[2][204] , \round_in[2][203] , 
        \round_in[2][202] , \round_in[2][201] , \round_in[2][200] , 
        \round_in[2][199] , \round_in[2][198] , \round_in[2][197] , 
        \round_in[2][196] , \round_in[2][195] , \round_in[2][194] , 
        \round_in[2][193] , \round_in[2][192] , \round_in[2][191] , 
        \round_in[2][190] , \round_in[2][189] , \round_in[2][188] , 
        \round_in[2][187] , \round_in[2][186] , \round_in[2][185] , 
        \round_in[2][184] , \round_in[2][183] , \round_in[2][182] , 
        \round_in[2][181] , \round_in[2][180] , \round_in[2][179] , 
        \round_in[2][178] , \round_in[2][177] , \round_in[2][176] , 
        \round_in[2][175] , \round_in[2][174] , \round_in[2][173] , 
        \round_in[2][172] , \round_in[2][171] , \round_in[2][170] , 
        \round_in[2][169] , \round_in[2][168] , \round_in[2][167] , 
        \round_in[2][166] , \round_in[2][165] , \round_in[2][164] , 
        \round_in[2][163] , \round_in[2][162] , \round_in[2][161] , 
        \round_in[2][160] , \round_in[2][159] , \round_in[2][158] , 
        \round_in[2][157] , \round_in[2][156] , \round_in[2][155] , 
        \round_in[2][154] , \round_in[2][153] , \round_in[2][152] , 
        \round_in[2][151] , \round_in[2][150] , \round_in[2][149] , 
        \round_in[2][148] , \round_in[2][147] , \round_in[2][146] , 
        \round_in[2][145] , \round_in[2][144] , \round_in[2][143] , 
        \round_in[2][142] , \round_in[2][141] , \round_in[2][140] , 
        \round_in[2][139] , \round_in[2][138] , \round_in[2][137] , 
        \round_in[2][136] , \round_in[2][135] , \round_in[2][134] , 
        \round_in[2][133] , \round_in[2][132] , \round_in[2][131] , 
        \round_in[2][130] , \round_in[2][129] , \round_in[2][128] , 
        \round_in[2][127] , \round_in[2][126] , \round_in[2][125] , 
        \round_in[2][124] , \round_in[2][123] , \round_in[2][122] , 
        \round_in[2][121] , \round_in[2][120] , \round_in[2][119] , 
        \round_in[2][118] , \round_in[2][117] , \round_in[2][116] , 
        \round_in[2][115] , \round_in[2][114] , \round_in[2][113] , 
        \round_in[2][112] , \round_in[2][111] , \round_in[2][110] , 
        \round_in[2][109] , \round_in[2][108] , \round_in[2][107] , 
        \round_in[2][106] , \round_in[2][105] , \round_in[2][104] , 
        \round_in[2][103] , \round_in[2][102] , \round_in[2][101] , 
        \round_in[2][100] , \round_in[2][99] , \round_in[2][98] , 
        \round_in[2][97] , \round_in[2][96] , \round_in[2][95] , 
        \round_in[2][94] , \round_in[2][93] , \round_in[2][92] , 
        \round_in[2][91] , \round_in[2][90] , \round_in[2][89] , 
        \round_in[2][88] , \round_in[2][87] , \round_in[2][86] , 
        \round_in[2][85] , \round_in[2][84] , \round_in[2][83] , 
        \round_in[2][82] , \round_in[2][81] , \round_in[2][80] , 
        \round_in[2][79] , \round_in[2][78] , \round_in[2][77] , 
        \round_in[2][76] , \round_in[2][75] , \round_in[2][74] , 
        \round_in[2][73] , \round_in[2][72] , \round_in[2][71] , 
        \round_in[2][70] , \round_in[2][69] , \round_in[2][68] , 
        \round_in[2][67] , \round_in[2][66] , \round_in[2][65] , 
        \round_in[2][64] , \round_in[2][63] , \round_in[2][62] , 
        \round_in[2][61] , \round_in[2][60] , \round_in[2][59] , 
        \round_in[2][58] , \round_in[2][57] , \round_in[2][56] , 
        \round_in[2][55] , \round_in[2][54] , \round_in[2][53] , 
        \round_in[2][52] , \round_in[2][51] , \round_in[2][50] , 
        \round_in[2][49] , \round_in[2][48] , \round_in[2][47] , 
        \round_in[2][46] , \round_in[2][45] , \round_in[2][44] , 
        \round_in[2][43] , \round_in[2][42] , \round_in[2][41] , 
        \round_in[2][40] , \round_in[2][39] , \round_in[2][38] , 
        \round_in[2][37] , \round_in[2][36] , \round_in[2][35] , 
        \round_in[2][34] , \round_in[2][33] , \round_in[2][32] , 
        \round_in[2][31] , \round_in[2][30] , \round_in[2][29] , 
        \round_in[2][28] , \round_in[2][27] , \round_in[2][26] , 
        \round_in[2][25] , \round_in[2][24] , \round_in[2][23] , 
        \round_in[2][22] , \round_in[2][21] , \round_in[2][20] , 
        \round_in[2][19] , \round_in[2][18] , \round_in[2][17] , 
        \round_in[2][16] , \round_in[2][15] , \round_in[2][14] , 
        \round_in[2][13] , \round_in[2][12] , \round_in[2][11] , 
        \round_in[2][10] , \round_in[2][9] , \round_in[2][8] , 
        \round_in[2][7] , \round_in[2][6] , \round_in[2][5] , \round_in[2][4] , 
        \round_in[2][3] , \round_in[2][2] , \round_in[2][1] , \round_in[2][0] }), .round_const({n1610, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[2].rconst_/N57 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \RCONST[2].rconst_/N47 , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        n1610, 1'b0, 1'b0, 1'b0, \RCONST[2].rconst_/N28 , 1'b0, 
        \RCONST[2].rconst_/N18 , \rc[2][0] }), .out({\round_in[3][1599] , 
        \round_in[3][1598] , \round_in[3][1597] , \round_in[3][1596] , 
        \round_in[3][1595] , \round_in[3][1594] , \round_in[3][1593] , 
        \round_in[3][1592] , \round_in[3][1591] , \round_in[3][1590] , 
        \round_in[3][1589] , \round_in[3][1588] , \round_in[3][1587] , 
        \round_in[3][1586] , \round_in[3][1585] , \round_in[3][1584] , 
        \round_in[3][1583] , \round_in[3][1582] , \round_in[3][1581] , 
        \round_in[3][1580] , \round_in[3][1579] , \round_in[3][1578] , 
        \round_in[3][1577] , \round_in[3][1576] , \round_in[3][1575] , 
        \round_in[3][1574] , \round_in[3][1573] , \round_in[3][1572] , 
        \round_in[3][1571] , \round_in[3][1570] , \round_in[3][1569] , 
        \round_in[3][1568] , \round_in[3][1567] , \round_in[3][1566] , 
        \round_in[3][1565] , \round_in[3][1564] , \round_in[3][1563] , 
        \round_in[3][1562] , \round_in[3][1561] , \round_in[3][1560] , 
        \round_in[3][1559] , \round_in[3][1558] , \round_in[3][1557] , 
        \round_in[3][1556] , \round_in[3][1555] , \round_in[3][1554] , 
        \round_in[3][1553] , \round_in[3][1552] , \round_in[3][1551] , 
        \round_in[3][1550] , \round_in[3][1549] , \round_in[3][1548] , 
        \round_in[3][1547] , \round_in[3][1546] , \round_in[3][1545] , 
        \round_in[3][1544] , \round_in[3][1543] , \round_in[3][1542] , 
        \round_in[3][1541] , \round_in[3][1540] , \round_in[3][1539] , 
        \round_in[3][1538] , \round_in[3][1537] , \round_in[3][1536] , 
        \round_in[3][1535] , \round_in[3][1534] , \round_in[3][1533] , 
        \round_in[3][1532] , \round_in[3][1531] , \round_in[3][1530] , 
        \round_in[3][1529] , \round_in[3][1528] , \round_in[3][1527] , 
        \round_in[3][1526] , \round_in[3][1525] , \round_in[3][1524] , 
        \round_in[3][1523] , \round_in[3][1522] , \round_in[3][1521] , 
        \round_in[3][1520] , \round_in[3][1519] , \round_in[3][1518] , 
        \round_in[3][1517] , \round_in[3][1516] , \round_in[3][1515] , 
        \round_in[3][1514] , \round_in[3][1513] , \round_in[3][1512] , 
        \round_in[3][1511] , \round_in[3][1510] , \round_in[3][1509] , 
        \round_in[3][1508] , \round_in[3][1507] , \round_in[3][1506] , 
        \round_in[3][1505] , \round_in[3][1504] , \round_in[3][1503] , 
        \round_in[3][1502] , \round_in[3][1501] , \round_in[3][1500] , 
        \round_in[3][1499] , \round_in[3][1498] , \round_in[3][1497] , 
        \round_in[3][1496] , \round_in[3][1495] , \round_in[3][1494] , 
        \round_in[3][1493] , \round_in[3][1492] , \round_in[3][1491] , 
        \round_in[3][1490] , \round_in[3][1489] , \round_in[3][1488] , 
        \round_in[3][1487] , \round_in[3][1486] , \round_in[3][1485] , 
        \round_in[3][1484] , \round_in[3][1483] , \round_in[3][1482] , 
        \round_in[3][1481] , \round_in[3][1480] , \round_in[3][1479] , 
        \round_in[3][1478] , \round_in[3][1477] , \round_in[3][1476] , 
        \round_in[3][1475] , \round_in[3][1474] , \round_in[3][1473] , 
        \round_in[3][1472] , \round_in[3][1471] , \round_in[3][1470] , 
        \round_in[3][1469] , \round_in[3][1468] , \round_in[3][1467] , 
        \round_in[3][1466] , \round_in[3][1465] , \round_in[3][1464] , 
        \round_in[3][1463] , \round_in[3][1462] , \round_in[3][1461] , 
        \round_in[3][1460] , \round_in[3][1459] , \round_in[3][1458] , 
        \round_in[3][1457] , \round_in[3][1456] , \round_in[3][1455] , 
        \round_in[3][1454] , \round_in[3][1453] , \round_in[3][1452] , 
        \round_in[3][1451] , \round_in[3][1450] , \round_in[3][1449] , 
        \round_in[3][1448] , \round_in[3][1447] , \round_in[3][1446] , 
        \round_in[3][1445] , \round_in[3][1444] , \round_in[3][1443] , 
        \round_in[3][1442] , \round_in[3][1441] , \round_in[3][1440] , 
        \round_in[3][1439] , \round_in[3][1438] , \round_in[3][1437] , 
        \round_in[3][1436] , \round_in[3][1435] , \round_in[3][1434] , 
        \round_in[3][1433] , \round_in[3][1432] , \round_in[3][1431] , 
        \round_in[3][1430] , \round_in[3][1429] , \round_in[3][1428] , 
        \round_in[3][1427] , \round_in[3][1426] , \round_in[3][1425] , 
        \round_in[3][1424] , \round_in[3][1423] , \round_in[3][1422] , 
        \round_in[3][1421] , \round_in[3][1420] , \round_in[3][1419] , 
        \round_in[3][1418] , \round_in[3][1417] , \round_in[3][1416] , 
        \round_in[3][1415] , \round_in[3][1414] , \round_in[3][1413] , 
        \round_in[3][1412] , \round_in[3][1411] , \round_in[3][1410] , 
        \round_in[3][1409] , \round_in[3][1408] , \round_in[3][1407] , 
        \round_in[3][1406] , \round_in[3][1405] , \round_in[3][1404] , 
        \round_in[3][1403] , \round_in[3][1402] , \round_in[3][1401] , 
        \round_in[3][1400] , \round_in[3][1399] , \round_in[3][1398] , 
        \round_in[3][1397] , \round_in[3][1396] , \round_in[3][1395] , 
        \round_in[3][1394] , \round_in[3][1393] , \round_in[3][1392] , 
        \round_in[3][1391] , \round_in[3][1390] , \round_in[3][1389] , 
        \round_in[3][1388] , \round_in[3][1387] , \round_in[3][1386] , 
        \round_in[3][1385] , \round_in[3][1384] , \round_in[3][1383] , 
        \round_in[3][1382] , \round_in[3][1381] , \round_in[3][1380] , 
        \round_in[3][1379] , \round_in[3][1378] , \round_in[3][1377] , 
        \round_in[3][1376] , \round_in[3][1375] , \round_in[3][1374] , 
        \round_in[3][1373] , \round_in[3][1372] , \round_in[3][1371] , 
        \round_in[3][1370] , \round_in[3][1369] , \round_in[3][1368] , 
        \round_in[3][1367] , \round_in[3][1366] , \round_in[3][1365] , 
        \round_in[3][1364] , \round_in[3][1363] , \round_in[3][1362] , 
        \round_in[3][1361] , \round_in[3][1360] , \round_in[3][1359] , 
        \round_in[3][1358] , \round_in[3][1357] , \round_in[3][1356] , 
        \round_in[3][1355] , \round_in[3][1354] , \round_in[3][1353] , 
        \round_in[3][1352] , \round_in[3][1351] , \round_in[3][1350] , 
        \round_in[3][1349] , \round_in[3][1348] , \round_in[3][1347] , 
        \round_in[3][1346] , \round_in[3][1345] , \round_in[3][1344] , 
        \round_in[3][1343] , \round_in[3][1342] , \round_in[3][1341] , 
        \round_in[3][1340] , \round_in[3][1339] , \round_in[3][1338] , 
        \round_in[3][1337] , \round_in[3][1336] , \round_in[3][1335] , 
        \round_in[3][1334] , \round_in[3][1333] , \round_in[3][1332] , 
        \round_in[3][1331] , \round_in[3][1330] , \round_in[3][1329] , 
        \round_in[3][1328] , \round_in[3][1327] , \round_in[3][1326] , 
        \round_in[3][1325] , \round_in[3][1324] , \round_in[3][1323] , 
        \round_in[3][1322] , \round_in[3][1321] , \round_in[3][1320] , 
        \round_in[3][1319] , \round_in[3][1318] , \round_in[3][1317] , 
        \round_in[3][1316] , \round_in[3][1315] , \round_in[3][1314] , 
        \round_in[3][1313] , \round_in[3][1312] , \round_in[3][1311] , 
        \round_in[3][1310] , \round_in[3][1309] , \round_in[3][1308] , 
        \round_in[3][1307] , \round_in[3][1306] , \round_in[3][1305] , 
        \round_in[3][1304] , \round_in[3][1303] , \round_in[3][1302] , 
        \round_in[3][1301] , \round_in[3][1300] , \round_in[3][1299] , 
        \round_in[3][1298] , \round_in[3][1297] , \round_in[3][1296] , 
        \round_in[3][1295] , \round_in[3][1294] , \round_in[3][1293] , 
        \round_in[3][1292] , \round_in[3][1291] , \round_in[3][1290] , 
        \round_in[3][1289] , \round_in[3][1288] , \round_in[3][1287] , 
        \round_in[3][1286] , \round_in[3][1285] , \round_in[3][1284] , 
        \round_in[3][1283] , \round_in[3][1282] , \round_in[3][1281] , 
        \round_in[3][1280] , \round_in[3][1279] , \round_in[3][1278] , 
        \round_in[3][1277] , \round_in[3][1276] , \round_in[3][1275] , 
        \round_in[3][1274] , \round_in[3][1273] , \round_in[3][1272] , 
        \round_in[3][1271] , \round_in[3][1270] , \round_in[3][1269] , 
        \round_in[3][1268] , \round_in[3][1267] , \round_in[3][1266] , 
        \round_in[3][1265] , \round_in[3][1264] , \round_in[3][1263] , 
        \round_in[3][1262] , \round_in[3][1261] , \round_in[3][1260] , 
        \round_in[3][1259] , \round_in[3][1258] , \round_in[3][1257] , 
        \round_in[3][1256] , \round_in[3][1255] , \round_in[3][1254] , 
        \round_in[3][1253] , \round_in[3][1252] , \round_in[3][1251] , 
        \round_in[3][1250] , \round_in[3][1249] , \round_in[3][1248] , 
        \round_in[3][1247] , \round_in[3][1246] , \round_in[3][1245] , 
        \round_in[3][1244] , \round_in[3][1243] , \round_in[3][1242] , 
        \round_in[3][1241] , \round_in[3][1240] , \round_in[3][1239] , 
        \round_in[3][1238] , \round_in[3][1237] , \round_in[3][1236] , 
        \round_in[3][1235] , \round_in[3][1234] , \round_in[3][1233] , 
        \round_in[3][1232] , \round_in[3][1231] , \round_in[3][1230] , 
        \round_in[3][1229] , \round_in[3][1228] , \round_in[3][1227] , 
        \round_in[3][1226] , \round_in[3][1225] , \round_in[3][1224] , 
        \round_in[3][1223] , \round_in[3][1222] , \round_in[3][1221] , 
        \round_in[3][1220] , \round_in[3][1219] , \round_in[3][1218] , 
        \round_in[3][1217] , \round_in[3][1216] , \round_in[3][1215] , 
        \round_in[3][1214] , \round_in[3][1213] , \round_in[3][1212] , 
        \round_in[3][1211] , \round_in[3][1210] , \round_in[3][1209] , 
        \round_in[3][1208] , \round_in[3][1207] , \round_in[3][1206] , 
        \round_in[3][1205] , \round_in[3][1204] , \round_in[3][1203] , 
        \round_in[3][1202] , \round_in[3][1201] , \round_in[3][1200] , 
        \round_in[3][1199] , \round_in[3][1198] , \round_in[3][1197] , 
        \round_in[3][1196] , \round_in[3][1195] , \round_in[3][1194] , 
        \round_in[3][1193] , \round_in[3][1192] , \round_in[3][1191] , 
        \round_in[3][1190] , \round_in[3][1189] , \round_in[3][1188] , 
        \round_in[3][1187] , \round_in[3][1186] , \round_in[3][1185] , 
        \round_in[3][1184] , \round_in[3][1183] , \round_in[3][1182] , 
        \round_in[3][1181] , \round_in[3][1180] , \round_in[3][1179] , 
        \round_in[3][1178] , \round_in[3][1177] , \round_in[3][1176] , 
        \round_in[3][1175] , \round_in[3][1174] , \round_in[3][1173] , 
        \round_in[3][1172] , \round_in[3][1171] , \round_in[3][1170] , 
        \round_in[3][1169] , \round_in[3][1168] , \round_in[3][1167] , 
        \round_in[3][1166] , \round_in[3][1165] , \round_in[3][1164] , 
        \round_in[3][1163] , \round_in[3][1162] , \round_in[3][1161] , 
        \round_in[3][1160] , \round_in[3][1159] , \round_in[3][1158] , 
        \round_in[3][1157] , \round_in[3][1156] , \round_in[3][1155] , 
        \round_in[3][1154] , \round_in[3][1153] , \round_in[3][1152] , 
        \round_in[3][1151] , \round_in[3][1150] , \round_in[3][1149] , 
        \round_in[3][1148] , \round_in[3][1147] , \round_in[3][1146] , 
        \round_in[3][1145] , \round_in[3][1144] , \round_in[3][1143] , 
        \round_in[3][1142] , \round_in[3][1141] , \round_in[3][1140] , 
        \round_in[3][1139] , \round_in[3][1138] , \round_in[3][1137] , 
        \round_in[3][1136] , \round_in[3][1135] , \round_in[3][1134] , 
        \round_in[3][1133] , \round_in[3][1132] , \round_in[3][1131] , 
        \round_in[3][1130] , \round_in[3][1129] , \round_in[3][1128] , 
        \round_in[3][1127] , \round_in[3][1126] , \round_in[3][1125] , 
        \round_in[3][1124] , \round_in[3][1123] , \round_in[3][1122] , 
        \round_in[3][1121] , \round_in[3][1120] , \round_in[3][1119] , 
        \round_in[3][1118] , \round_in[3][1117] , \round_in[3][1116] , 
        \round_in[3][1115] , \round_in[3][1114] , \round_in[3][1113] , 
        \round_in[3][1112] , \round_in[3][1111] , \round_in[3][1110] , 
        \round_in[3][1109] , \round_in[3][1108] , \round_in[3][1107] , 
        \round_in[3][1106] , \round_in[3][1105] , \round_in[3][1104] , 
        \round_in[3][1103] , \round_in[3][1102] , \round_in[3][1101] , 
        \round_in[3][1100] , \round_in[3][1099] , \round_in[3][1098] , 
        \round_in[3][1097] , \round_in[3][1096] , \round_in[3][1095] , 
        \round_in[3][1094] , \round_in[3][1093] , \round_in[3][1092] , 
        \round_in[3][1091] , \round_in[3][1090] , \round_in[3][1089] , 
        \round_in[3][1088] , \round_in[3][1087] , \round_in[3][1086] , 
        \round_in[3][1085] , \round_in[3][1084] , \round_in[3][1083] , 
        \round_in[3][1082] , \round_in[3][1081] , \round_in[3][1080] , 
        \round_in[3][1079] , \round_in[3][1078] , \round_in[3][1077] , 
        \round_in[3][1076] , \round_in[3][1075] , \round_in[3][1074] , 
        \round_in[3][1073] , \round_in[3][1072] , \round_in[3][1071] , 
        \round_in[3][1070] , \round_in[3][1069] , \round_in[3][1068] , 
        \round_in[3][1067] , \round_in[3][1066] , \round_in[3][1065] , 
        \round_in[3][1064] , \round_in[3][1063] , \round_in[3][1062] , 
        \round_in[3][1061] , \round_in[3][1060] , \round_in[3][1059] , 
        \round_in[3][1058] , \round_in[3][1057] , \round_in[3][1056] , 
        \round_in[3][1055] , \round_in[3][1054] , \round_in[3][1053] , 
        \round_in[3][1052] , \round_in[3][1051] , \round_in[3][1050] , 
        \round_in[3][1049] , \round_in[3][1048] , \round_in[3][1047] , 
        \round_in[3][1046] , \round_in[3][1045] , \round_in[3][1044] , 
        \round_in[3][1043] , \round_in[3][1042] , \round_in[3][1041] , 
        \round_in[3][1040] , \round_in[3][1039] , \round_in[3][1038] , 
        \round_in[3][1037] , \round_in[3][1036] , \round_in[3][1035] , 
        \round_in[3][1034] , \round_in[3][1033] , \round_in[3][1032] , 
        \round_in[3][1031] , \round_in[3][1030] , \round_in[3][1029] , 
        \round_in[3][1028] , \round_in[3][1027] , \round_in[3][1026] , 
        \round_in[3][1025] , \round_in[3][1024] , \round_in[3][1023] , 
        \round_in[3][1022] , \round_in[3][1021] , \round_in[3][1020] , 
        \round_in[3][1019] , \round_in[3][1018] , \round_in[3][1017] , 
        \round_in[3][1016] , \round_in[3][1015] , \round_in[3][1014] , 
        \round_in[3][1013] , \round_in[3][1012] , \round_in[3][1011] , 
        \round_in[3][1010] , \round_in[3][1009] , \round_in[3][1008] , 
        \round_in[3][1007] , \round_in[3][1006] , \round_in[3][1005] , 
        \round_in[3][1004] , \round_in[3][1003] , \round_in[3][1002] , 
        \round_in[3][1001] , \round_in[3][1000] , \round_in[3][999] , 
        \round_in[3][998] , \round_in[3][997] , \round_in[3][996] , 
        \round_in[3][995] , \round_in[3][994] , \round_in[3][993] , 
        \round_in[3][992] , \round_in[3][991] , \round_in[3][990] , 
        \round_in[3][989] , \round_in[3][988] , \round_in[3][987] , 
        \round_in[3][986] , \round_in[3][985] , \round_in[3][984] , 
        \round_in[3][983] , \round_in[3][982] , \round_in[3][981] , 
        \round_in[3][980] , \round_in[3][979] , \round_in[3][978] , 
        \round_in[3][977] , \round_in[3][976] , \round_in[3][975] , 
        \round_in[3][974] , \round_in[3][973] , \round_in[3][972] , 
        \round_in[3][971] , \round_in[3][970] , \round_in[3][969] , 
        \round_in[3][968] , \round_in[3][967] , \round_in[3][966] , 
        \round_in[3][965] , \round_in[3][964] , \round_in[3][963] , 
        \round_in[3][962] , \round_in[3][961] , \round_in[3][960] , 
        \round_in[3][959] , \round_in[3][958] , \round_in[3][957] , 
        \round_in[3][956] , \round_in[3][955] , \round_in[3][954] , 
        \round_in[3][953] , \round_in[3][952] , \round_in[3][951] , 
        \round_in[3][950] , \round_in[3][949] , \round_in[3][948] , 
        \round_in[3][947] , \round_in[3][946] , \round_in[3][945] , 
        \round_in[3][944] , \round_in[3][943] , \round_in[3][942] , 
        \round_in[3][941] , \round_in[3][940] , \round_in[3][939] , 
        \round_in[3][938] , \round_in[3][937] , \round_in[3][936] , 
        \round_in[3][935] , \round_in[3][934] , \round_in[3][933] , 
        \round_in[3][932] , \round_in[3][931] , \round_in[3][930] , 
        \round_in[3][929] , \round_in[3][928] , \round_in[3][927] , 
        \round_in[3][926] , \round_in[3][925] , \round_in[3][924] , 
        \round_in[3][923] , \round_in[3][922] , \round_in[3][921] , 
        \round_in[3][920] , \round_in[3][919] , \round_in[3][918] , 
        \round_in[3][917] , \round_in[3][916] , \round_in[3][915] , 
        \round_in[3][914] , \round_in[3][913] , \round_in[3][912] , 
        \round_in[3][911] , \round_in[3][910] , \round_in[3][909] , 
        \round_in[3][908] , \round_in[3][907] , \round_in[3][906] , 
        \round_in[3][905] , \round_in[3][904] , \round_in[3][903] , 
        \round_in[3][902] , \round_in[3][901] , \round_in[3][900] , 
        \round_in[3][899] , \round_in[3][898] , \round_in[3][897] , 
        \round_in[3][896] , \round_in[3][895] , \round_in[3][894] , 
        \round_in[3][893] , \round_in[3][892] , \round_in[3][891] , 
        \round_in[3][890] , \round_in[3][889] , \round_in[3][888] , 
        \round_in[3][887] , \round_in[3][886] , \round_in[3][885] , 
        \round_in[3][884] , \round_in[3][883] , \round_in[3][882] , 
        \round_in[3][881] , \round_in[3][880] , \round_in[3][879] , 
        \round_in[3][878] , \round_in[3][877] , \round_in[3][876] , 
        \round_in[3][875] , \round_in[3][874] , \round_in[3][873] , 
        \round_in[3][872] , \round_in[3][871] , \round_in[3][870] , 
        \round_in[3][869] , \round_in[3][868] , \round_in[3][867] , 
        \round_in[3][866] , \round_in[3][865] , \round_in[3][864] , 
        \round_in[3][863] , \round_in[3][862] , \round_in[3][861] , 
        \round_in[3][860] , \round_in[3][859] , \round_in[3][858] , 
        \round_in[3][857] , \round_in[3][856] , \round_in[3][855] , 
        \round_in[3][854] , \round_in[3][853] , \round_in[3][852] , 
        \round_in[3][851] , \round_in[3][850] , \round_in[3][849] , 
        \round_in[3][848] , \round_in[3][847] , \round_in[3][846] , 
        \round_in[3][845] , \round_in[3][844] , \round_in[3][843] , 
        \round_in[3][842] , \round_in[3][841] , \round_in[3][840] , 
        \round_in[3][839] , \round_in[3][838] , \round_in[3][837] , 
        \round_in[3][836] , \round_in[3][835] , \round_in[3][834] , 
        \round_in[3][833] , \round_in[3][832] , \round_in[3][831] , 
        \round_in[3][830] , \round_in[3][829] , \round_in[3][828] , 
        \round_in[3][827] , \round_in[3][826] , \round_in[3][825] , 
        \round_in[3][824] , \round_in[3][823] , \round_in[3][822] , 
        \round_in[3][821] , \round_in[3][820] , \round_in[3][819] , 
        \round_in[3][818] , \round_in[3][817] , \round_in[3][816] , 
        \round_in[3][815] , \round_in[3][814] , \round_in[3][813] , 
        \round_in[3][812] , \round_in[3][811] , \round_in[3][810] , 
        \round_in[3][809] , \round_in[3][808] , \round_in[3][807] , 
        \round_in[3][806] , \round_in[3][805] , \round_in[3][804] , 
        \round_in[3][803] , \round_in[3][802] , \round_in[3][801] , 
        \round_in[3][800] , \round_in[3][799] , \round_in[3][798] , 
        \round_in[3][797] , \round_in[3][796] , \round_in[3][795] , 
        \round_in[3][794] , \round_in[3][793] , \round_in[3][792] , 
        \round_in[3][791] , \round_in[3][790] , \round_in[3][789] , 
        \round_in[3][788] , \round_in[3][787] , \round_in[3][786] , 
        \round_in[3][785] , \round_in[3][784] , \round_in[3][783] , 
        \round_in[3][782] , \round_in[3][781] , \round_in[3][780] , 
        \round_in[3][779] , \round_in[3][778] , \round_in[3][777] , 
        \round_in[3][776] , \round_in[3][775] , \round_in[3][774] , 
        \round_in[3][773] , \round_in[3][772] , \round_in[3][771] , 
        \round_in[3][770] , \round_in[3][769] , \round_in[3][768] , 
        \round_in[3][767] , \round_in[3][766] , \round_in[3][765] , 
        \round_in[3][764] , \round_in[3][763] , \round_in[3][762] , 
        \round_in[3][761] , \round_in[3][760] , \round_in[3][759] , 
        \round_in[3][758] , \round_in[3][757] , \round_in[3][756] , 
        \round_in[3][755] , \round_in[3][754] , \round_in[3][753] , 
        \round_in[3][752] , \round_in[3][751] , \round_in[3][750] , 
        \round_in[3][749] , \round_in[3][748] , \round_in[3][747] , 
        \round_in[3][746] , \round_in[3][745] , \round_in[3][744] , 
        \round_in[3][743] , \round_in[3][742] , \round_in[3][741] , 
        \round_in[3][740] , \round_in[3][739] , \round_in[3][738] , 
        \round_in[3][737] , \round_in[3][736] , \round_in[3][735] , 
        \round_in[3][734] , \round_in[3][733] , \round_in[3][732] , 
        \round_in[3][731] , \round_in[3][730] , \round_in[3][729] , 
        \round_in[3][728] , \round_in[3][727] , \round_in[3][726] , 
        \round_in[3][725] , \round_in[3][724] , \round_in[3][723] , 
        \round_in[3][722] , \round_in[3][721] , \round_in[3][720] , 
        \round_in[3][719] , \round_in[3][718] , \round_in[3][717] , 
        \round_in[3][716] , \round_in[3][715] , \round_in[3][714] , 
        \round_in[3][713] , \round_in[3][712] , \round_in[3][711] , 
        \round_in[3][710] , \round_in[3][709] , \round_in[3][708] , 
        \round_in[3][707] , \round_in[3][706] , \round_in[3][705] , 
        \round_in[3][704] , \round_in[3][703] , \round_in[3][702] , 
        \round_in[3][701] , \round_in[3][700] , \round_in[3][699] , 
        \round_in[3][698] , \round_in[3][697] , \round_in[3][696] , 
        \round_in[3][695] , \round_in[3][694] , \round_in[3][693] , 
        \round_in[3][692] , \round_in[3][691] , \round_in[3][690] , 
        \round_in[3][689] , \round_in[3][688] , \round_in[3][687] , 
        \round_in[3][686] , \round_in[3][685] , \round_in[3][684] , 
        \round_in[3][683] , \round_in[3][682] , \round_in[3][681] , 
        \round_in[3][680] , \round_in[3][679] , \round_in[3][678] , 
        \round_in[3][677] , \round_in[3][676] , \round_in[3][675] , 
        \round_in[3][674] , \round_in[3][673] , \round_in[3][672] , 
        \round_in[3][671] , \round_in[3][670] , \round_in[3][669] , 
        \round_in[3][668] , \round_in[3][667] , \round_in[3][666] , 
        \round_in[3][665] , \round_in[3][664] , \round_in[3][663] , 
        \round_in[3][662] , \round_in[3][661] , \round_in[3][660] , 
        \round_in[3][659] , \round_in[3][658] , \round_in[3][657] , 
        \round_in[3][656] , \round_in[3][655] , \round_in[3][654] , 
        \round_in[3][653] , \round_in[3][652] , \round_in[3][651] , 
        \round_in[3][650] , \round_in[3][649] , \round_in[3][648] , 
        \round_in[3][647] , \round_in[3][646] , \round_in[3][645] , 
        \round_in[3][644] , \round_in[3][643] , \round_in[3][642] , 
        \round_in[3][641] , \round_in[3][640] , \round_in[3][639] , 
        \round_in[3][638] , \round_in[3][637] , \round_in[3][636] , 
        \round_in[3][635] , \round_in[3][634] , \round_in[3][633] , 
        \round_in[3][632] , \round_in[3][631] , \round_in[3][630] , 
        \round_in[3][629] , \round_in[3][628] , \round_in[3][627] , 
        \round_in[3][626] , \round_in[3][625] , \round_in[3][624] , 
        \round_in[3][623] , \round_in[3][622] , \round_in[3][621] , 
        \round_in[3][620] , \round_in[3][619] , \round_in[3][618] , 
        \round_in[3][617] , \round_in[3][616] , \round_in[3][615] , 
        \round_in[3][614] , \round_in[3][613] , \round_in[3][612] , 
        \round_in[3][611] , \round_in[3][610] , \round_in[3][609] , 
        \round_in[3][608] , \round_in[3][607] , \round_in[3][606] , 
        \round_in[3][605] , \round_in[3][604] , \round_in[3][603] , 
        \round_in[3][602] , \round_in[3][601] , \round_in[3][600] , 
        \round_in[3][599] , \round_in[3][598] , \round_in[3][597] , 
        \round_in[3][596] , \round_in[3][595] , \round_in[3][594] , 
        \round_in[3][593] , \round_in[3][592] , \round_in[3][591] , 
        \round_in[3][590] , \round_in[3][589] , \round_in[3][588] , 
        \round_in[3][587] , \round_in[3][586] , \round_in[3][585] , 
        \round_in[3][584] , \round_in[3][583] , \round_in[3][582] , 
        \round_in[3][581] , \round_in[3][580] , \round_in[3][579] , 
        \round_in[3][578] , \round_in[3][577] , \round_in[3][576] , 
        \round_in[3][575] , \round_in[3][574] , \round_in[3][573] , 
        \round_in[3][572] , \round_in[3][571] , \round_in[3][570] , 
        \round_in[3][569] , \round_in[3][568] , \round_in[3][567] , 
        \round_in[3][566] , \round_in[3][565] , \round_in[3][564] , 
        \round_in[3][563] , \round_in[3][562] , \round_in[3][561] , 
        \round_in[3][560] , \round_in[3][559] , \round_in[3][558] , 
        \round_in[3][557] , \round_in[3][556] , \round_in[3][555] , 
        \round_in[3][554] , \round_in[3][553] , \round_in[3][552] , 
        \round_in[3][551] , \round_in[3][550] , \round_in[3][549] , 
        \round_in[3][548] , \round_in[3][547] , \round_in[3][546] , 
        \round_in[3][545] , \round_in[3][544] , \round_in[3][543] , 
        \round_in[3][542] , \round_in[3][541] , \round_in[3][540] , 
        \round_in[3][539] , \round_in[3][538] , \round_in[3][537] , 
        \round_in[3][536] , \round_in[3][535] , \round_in[3][534] , 
        \round_in[3][533] , \round_in[3][532] , \round_in[3][531] , 
        \round_in[3][530] , \round_in[3][529] , \round_in[3][528] , 
        \round_in[3][527] , \round_in[3][526] , \round_in[3][525] , 
        \round_in[3][524] , \round_in[3][523] , \round_in[3][522] , 
        \round_in[3][521] , \round_in[3][520] , \round_in[3][519] , 
        \round_in[3][518] , \round_in[3][517] , \round_in[3][516] , 
        \round_in[3][515] , \round_in[3][514] , \round_in[3][513] , 
        \round_in[3][512] , \round_in[3][511] , \round_in[3][510] , 
        \round_in[3][509] , \round_in[3][508] , \round_in[3][507] , 
        \round_in[3][506] , \round_in[3][505] , \round_in[3][504] , 
        \round_in[3][503] , \round_in[3][502] , \round_in[3][501] , 
        \round_in[3][500] , \round_in[3][499] , \round_in[3][498] , 
        \round_in[3][497] , \round_in[3][496] , \round_in[3][495] , 
        \round_in[3][494] , \round_in[3][493] , \round_in[3][492] , 
        \round_in[3][491] , \round_in[3][490] , \round_in[3][489] , 
        \round_in[3][488] , \round_in[3][487] , \round_in[3][486] , 
        \round_in[3][485] , \round_in[3][484] , \round_in[3][483] , 
        \round_in[3][482] , \round_in[3][481] , \round_in[3][480] , 
        \round_in[3][479] , \round_in[3][478] , \round_in[3][477] , 
        \round_in[3][476] , \round_in[3][475] , \round_in[3][474] , 
        \round_in[3][473] , \round_in[3][472] , \round_in[3][471] , 
        \round_in[3][470] , \round_in[3][469] , \round_in[3][468] , 
        \round_in[3][467] , \round_in[3][466] , \round_in[3][465] , 
        \round_in[3][464] , \round_in[3][463] , \round_in[3][462] , 
        \round_in[3][461] , \round_in[3][460] , \round_in[3][459] , 
        \round_in[3][458] , \round_in[3][457] , \round_in[3][456] , 
        \round_in[3][455] , \round_in[3][454] , \round_in[3][453] , 
        \round_in[3][452] , \round_in[3][451] , \round_in[3][450] , 
        \round_in[3][449] , \round_in[3][448] , \round_in[3][447] , 
        \round_in[3][446] , \round_in[3][445] , \round_in[3][444] , 
        \round_in[3][443] , \round_in[3][442] , \round_in[3][441] , 
        \round_in[3][440] , \round_in[3][439] , \round_in[3][438] , 
        \round_in[3][437] , \round_in[3][436] , \round_in[3][435] , 
        \round_in[3][434] , \round_in[3][433] , \round_in[3][432] , 
        \round_in[3][431] , \round_in[3][430] , \round_in[3][429] , 
        \round_in[3][428] , \round_in[3][427] , \round_in[3][426] , 
        \round_in[3][425] , \round_in[3][424] , \round_in[3][423] , 
        \round_in[3][422] , \round_in[3][421] , \round_in[3][420] , 
        \round_in[3][419] , \round_in[3][418] , \round_in[3][417] , 
        \round_in[3][416] , \round_in[3][415] , \round_in[3][414] , 
        \round_in[3][413] , \round_in[3][412] , \round_in[3][411] , 
        \round_in[3][410] , \round_in[3][409] , \round_in[3][408] , 
        \round_in[3][407] , \round_in[3][406] , \round_in[3][405] , 
        \round_in[3][404] , \round_in[3][403] , \round_in[3][402] , 
        \round_in[3][401] , \round_in[3][400] , \round_in[3][399] , 
        \round_in[3][398] , \round_in[3][397] , \round_in[3][396] , 
        \round_in[3][395] , \round_in[3][394] , \round_in[3][393] , 
        \round_in[3][392] , \round_in[3][391] , \round_in[3][390] , 
        \round_in[3][389] , \round_in[3][388] , \round_in[3][387] , 
        \round_in[3][386] , \round_in[3][385] , \round_in[3][384] , 
        \round_in[3][383] , \round_in[3][382] , \round_in[3][381] , 
        \round_in[3][380] , \round_in[3][379] , \round_in[3][378] , 
        \round_in[3][377] , \round_in[3][376] , \round_in[3][375] , 
        \round_in[3][374] , \round_in[3][373] , \round_in[3][372] , 
        \round_in[3][371] , \round_in[3][370] , \round_in[3][369] , 
        \round_in[3][368] , \round_in[3][367] , \round_in[3][366] , 
        \round_in[3][365] , \round_in[3][364] , \round_in[3][363] , 
        \round_in[3][362] , \round_in[3][361] , \round_in[3][360] , 
        \round_in[3][359] , \round_in[3][358] , \round_in[3][357] , 
        \round_in[3][356] , \round_in[3][355] , \round_in[3][354] , 
        \round_in[3][353] , \round_in[3][352] , \round_in[3][351] , 
        \round_in[3][350] , \round_in[3][349] , \round_in[3][348] , 
        \round_in[3][347] , \round_in[3][346] , \round_in[3][345] , 
        \round_in[3][344] , \round_in[3][343] , \round_in[3][342] , 
        \round_in[3][341] , \round_in[3][340] , \round_in[3][339] , 
        \round_in[3][338] , \round_in[3][337] , \round_in[3][336] , 
        \round_in[3][335] , \round_in[3][334] , \round_in[3][333] , 
        \round_in[3][332] , \round_in[3][331] , \round_in[3][330] , 
        \round_in[3][329] , \round_in[3][328] , \round_in[3][327] , 
        \round_in[3][326] , \round_in[3][325] , \round_in[3][324] , 
        \round_in[3][323] , \round_in[3][322] , \round_in[3][321] , 
        \round_in[3][320] , \round_in[3][319] , \round_in[3][318] , 
        \round_in[3][317] , \round_in[3][316] , \round_in[3][315] , 
        \round_in[3][314] , \round_in[3][313] , \round_in[3][312] , 
        \round_in[3][311] , \round_in[3][310] , \round_in[3][309] , 
        \round_in[3][308] , \round_in[3][307] , \round_in[3][306] , 
        \round_in[3][305] , \round_in[3][304] , \round_in[3][303] , 
        \round_in[3][302] , \round_in[3][301] , \round_in[3][300] , 
        \round_in[3][299] , \round_in[3][298] , \round_in[3][297] , 
        \round_in[3][296] , \round_in[3][295] , \round_in[3][294] , 
        \round_in[3][293] , \round_in[3][292] , \round_in[3][291] , 
        \round_in[3][290] , \round_in[3][289] , \round_in[3][288] , 
        \round_in[3][287] , \round_in[3][286] , \round_in[3][285] , 
        \round_in[3][284] , \round_in[3][283] , \round_in[3][282] , 
        \round_in[3][281] , \round_in[3][280] , \round_in[3][279] , 
        \round_in[3][278] , \round_in[3][277] , \round_in[3][276] , 
        \round_in[3][275] , \round_in[3][274] , \round_in[3][273] , 
        \round_in[3][272] , \round_in[3][271] , \round_in[3][270] , 
        \round_in[3][269] , \round_in[3][268] , \round_in[3][267] , 
        \round_in[3][266] , \round_in[3][265] , \round_in[3][264] , 
        \round_in[3][263] , \round_in[3][262] , \round_in[3][261] , 
        \round_in[3][260] , \round_in[3][259] , \round_in[3][258] , 
        \round_in[3][257] , \round_in[3][256] , \round_in[3][255] , 
        \round_in[3][254] , \round_in[3][253] , \round_in[3][252] , 
        \round_in[3][251] , \round_in[3][250] , \round_in[3][249] , 
        \round_in[3][248] , \round_in[3][247] , \round_in[3][246] , 
        \round_in[3][245] , \round_in[3][244] , \round_in[3][243] , 
        \round_in[3][242] , \round_in[3][241] , \round_in[3][240] , 
        \round_in[3][239] , \round_in[3][238] , \round_in[3][237] , 
        \round_in[3][236] , \round_in[3][235] , \round_in[3][234] , 
        \round_in[3][233] , \round_in[3][232] , \round_in[3][231] , 
        \round_in[3][230] , \round_in[3][229] , \round_in[3][228] , 
        \round_in[3][227] , \round_in[3][226] , \round_in[3][225] , 
        \round_in[3][224] , \round_in[3][223] , \round_in[3][222] , 
        \round_in[3][221] , \round_in[3][220] , \round_in[3][219] , 
        \round_in[3][218] , \round_in[3][217] , \round_in[3][216] , 
        \round_in[3][215] , \round_in[3][214] , \round_in[3][213] , 
        \round_in[3][212] , \round_in[3][211] , \round_in[3][210] , 
        \round_in[3][209] , \round_in[3][208] , \round_in[3][207] , 
        \round_in[3][206] , \round_in[3][205] , \round_in[3][204] , 
        \round_in[3][203] , \round_in[3][202] , \round_in[3][201] , 
        \round_in[3][200] , \round_in[3][199] , \round_in[3][198] , 
        \round_in[3][197] , \round_in[3][196] , \round_in[3][195] , 
        \round_in[3][194] , \round_in[3][193] , \round_in[3][192] , 
        \round_in[3][191] , \round_in[3][190] , \round_in[3][189] , 
        \round_in[3][188] , \round_in[3][187] , \round_in[3][186] , 
        \round_in[3][185] , \round_in[3][184] , \round_in[3][183] , 
        \round_in[3][182] , \round_in[3][181] , \round_in[3][180] , 
        \round_in[3][179] , \round_in[3][178] , \round_in[3][177] , 
        \round_in[3][176] , \round_in[3][175] , \round_in[3][174] , 
        \round_in[3][173] , \round_in[3][172] , \round_in[3][171] , 
        \round_in[3][170] , \round_in[3][169] , \round_in[3][168] , 
        \round_in[3][167] , \round_in[3][166] , \round_in[3][165] , 
        \round_in[3][164] , \round_in[3][163] , \round_in[3][162] , 
        \round_in[3][161] , \round_in[3][160] , \round_in[3][159] , 
        \round_in[3][158] , \round_in[3][157] , \round_in[3][156] , 
        \round_in[3][155] , \round_in[3][154] , \round_in[3][153] , 
        \round_in[3][152] , \round_in[3][151] , \round_in[3][150] , 
        \round_in[3][149] , \round_in[3][148] , \round_in[3][147] , 
        \round_in[3][146] , \round_in[3][145] , \round_in[3][144] , 
        \round_in[3][143] , \round_in[3][142] , \round_in[3][141] , 
        \round_in[3][140] , \round_in[3][139] , \round_in[3][138] , 
        \round_in[3][137] , \round_in[3][136] , \round_in[3][135] , 
        \round_in[3][134] , \round_in[3][133] , \round_in[3][132] , 
        \round_in[3][131] , \round_in[3][130] , \round_in[3][129] , 
        \round_in[3][128] , \round_in[3][127] , \round_in[3][126] , 
        \round_in[3][125] , \round_in[3][124] , \round_in[3][123] , 
        \round_in[3][122] , \round_in[3][121] , \round_in[3][120] , 
        \round_in[3][119] , \round_in[3][118] , \round_in[3][117] , 
        \round_in[3][116] , \round_in[3][115] , \round_in[3][114] , 
        \round_in[3][113] , \round_in[3][112] , \round_in[3][111] , 
        \round_in[3][110] , \round_in[3][109] , \round_in[3][108] , 
        \round_in[3][107] , \round_in[3][106] , \round_in[3][105] , 
        \round_in[3][104] , \round_in[3][103] , \round_in[3][102] , 
        \round_in[3][101] , \round_in[3][100] , \round_in[3][99] , 
        \round_in[3][98] , \round_in[3][97] , \round_in[3][96] , 
        \round_in[3][95] , \round_in[3][94] , \round_in[3][93] , 
        \round_in[3][92] , \round_in[3][91] , \round_in[3][90] , 
        \round_in[3][89] , \round_in[3][88] , \round_in[3][87] , 
        \round_in[3][86] , \round_in[3][85] , \round_in[3][84] , 
        \round_in[3][83] , \round_in[3][82] , \round_in[3][81] , 
        \round_in[3][80] , \round_in[3][79] , \round_in[3][78] , 
        \round_in[3][77] , \round_in[3][76] , \round_in[3][75] , 
        \round_in[3][74] , \round_in[3][73] , \round_in[3][72] , 
        \round_in[3][71] , \round_in[3][70] , \round_in[3][69] , 
        \round_in[3][68] , \round_in[3][67] , \round_in[3][66] , 
        \round_in[3][65] , \round_in[3][64] , \round_in[3][63] , 
        \round_in[3][62] , \round_in[3][61] , \round_in[3][60] , 
        \round_in[3][59] , \round_in[3][58] , \round_in[3][57] , 
        \round_in[3][56] , \round_in[3][55] , \round_in[3][54] , 
        \round_in[3][53] , \round_in[3][52] , \round_in[3][51] , 
        \round_in[3][50] , \round_in[3][49] , \round_in[3][48] , 
        \round_in[3][47] , \round_in[3][46] , \round_in[3][45] , 
        \round_in[3][44] , \round_in[3][43] , \round_in[3][42] , 
        \round_in[3][41] , \round_in[3][40] , \round_in[3][39] , 
        \round_in[3][38] , \round_in[3][37] , \round_in[3][36] , 
        \round_in[3][35] , \round_in[3][34] , \round_in[3][33] , 
        \round_in[3][32] , \round_in[3][31] , \round_in[3][30] , 
        \round_in[3][29] , \round_in[3][28] , \round_in[3][27] , 
        \round_in[3][26] , \round_in[3][25] , \round_in[3][24] , 
        \round_in[3][23] , \round_in[3][22] , \round_in[3][21] , 
        \round_in[3][20] , \round_in[3][19] , \round_in[3][18] , 
        \round_in[3][17] , \round_in[3][16] , \round_in[3][15] , 
        \round_in[3][14] , \round_in[3][13] , \round_in[3][12] , 
        \round_in[3][11] , \round_in[3][10] , \round_in[3][9] , 
        \round_in[3][8] , \round_in[3][7] , \round_in[3][6] , \round_in[3][5] , 
        \round_in[3][4] , \round_in[3][3] , \round_in[3][2] , \round_in[3][1] , 
        \round_in[3][0] }) );
  round_3 \ROUND[3].round_  ( .in({\round_in[3][1599] , \round_in[3][1598] , 
        \round_in[3][1597] , \round_in[3][1596] , \round_in[3][1595] , 
        \round_in[3][1594] , \round_in[3][1593] , \round_in[3][1592] , 
        \round_in[3][1591] , \round_in[3][1590] , \round_in[3][1589] , 
        \round_in[3][1588] , \round_in[3][1587] , \round_in[3][1586] , 
        \round_in[3][1585] , \round_in[3][1584] , \round_in[3][1583] , 
        \round_in[3][1582] , \round_in[3][1581] , \round_in[3][1580] , 
        \round_in[3][1579] , \round_in[3][1578] , \round_in[3][1577] , 
        \round_in[3][1576] , \round_in[3][1575] , \round_in[3][1574] , 
        \round_in[3][1573] , \round_in[3][1572] , \round_in[3][1571] , 
        \round_in[3][1570] , \round_in[3][1569] , \round_in[3][1568] , 
        \round_in[3][1567] , \round_in[3][1566] , \round_in[3][1565] , 
        \round_in[3][1564] , \round_in[3][1563] , \round_in[3][1562] , 
        \round_in[3][1561] , \round_in[3][1560] , \round_in[3][1559] , 
        \round_in[3][1558] , \round_in[3][1557] , \round_in[3][1556] , 
        \round_in[3][1555] , \round_in[3][1554] , \round_in[3][1553] , 
        \round_in[3][1552] , \round_in[3][1551] , \round_in[3][1550] , 
        \round_in[3][1549] , \round_in[3][1548] , \round_in[3][1547] , 
        \round_in[3][1546] , \round_in[3][1545] , \round_in[3][1544] , 
        \round_in[3][1543] , \round_in[3][1542] , \round_in[3][1541] , 
        \round_in[3][1540] , \round_in[3][1539] , \round_in[3][1538] , 
        \round_in[3][1537] , \round_in[3][1536] , \round_in[3][1535] , 
        \round_in[3][1534] , \round_in[3][1533] , \round_in[3][1532] , 
        \round_in[3][1531] , \round_in[3][1530] , \round_in[3][1529] , 
        \round_in[3][1528] , \round_in[3][1527] , \round_in[3][1526] , 
        \round_in[3][1525] , \round_in[3][1524] , \round_in[3][1523] , 
        \round_in[3][1522] , \round_in[3][1521] , \round_in[3][1520] , 
        \round_in[3][1519] , \round_in[3][1518] , \round_in[3][1517] , 
        \round_in[3][1516] , \round_in[3][1515] , \round_in[3][1514] , 
        \round_in[3][1513] , \round_in[3][1512] , \round_in[3][1511] , 
        \round_in[3][1510] , \round_in[3][1509] , \round_in[3][1508] , 
        \round_in[3][1507] , \round_in[3][1506] , \round_in[3][1505] , 
        \round_in[3][1504] , \round_in[3][1503] , \round_in[3][1502] , 
        \round_in[3][1501] , \round_in[3][1500] , \round_in[3][1499] , 
        \round_in[3][1498] , \round_in[3][1497] , \round_in[3][1496] , 
        \round_in[3][1495] , \round_in[3][1494] , \round_in[3][1493] , 
        \round_in[3][1492] , \round_in[3][1491] , \round_in[3][1490] , 
        \round_in[3][1489] , \round_in[3][1488] , \round_in[3][1487] , 
        \round_in[3][1486] , \round_in[3][1485] , \round_in[3][1484] , 
        \round_in[3][1483] , \round_in[3][1482] , \round_in[3][1481] , 
        \round_in[3][1480] , \round_in[3][1479] , \round_in[3][1478] , 
        \round_in[3][1477] , \round_in[3][1476] , \round_in[3][1475] , 
        \round_in[3][1474] , \round_in[3][1473] , \round_in[3][1472] , 
        \round_in[3][1471] , \round_in[3][1470] , \round_in[3][1469] , 
        \round_in[3][1468] , \round_in[3][1467] , \round_in[3][1466] , 
        \round_in[3][1465] , \round_in[3][1464] , \round_in[3][1463] , 
        \round_in[3][1462] , \round_in[3][1461] , \round_in[3][1460] , 
        \round_in[3][1459] , \round_in[3][1458] , \round_in[3][1457] , 
        \round_in[3][1456] , \round_in[3][1455] , \round_in[3][1454] , 
        \round_in[3][1453] , \round_in[3][1452] , \round_in[3][1451] , 
        \round_in[3][1450] , \round_in[3][1449] , \round_in[3][1448] , 
        \round_in[3][1447] , \round_in[3][1446] , \round_in[3][1445] , 
        \round_in[3][1444] , \round_in[3][1443] , \round_in[3][1442] , 
        \round_in[3][1441] , \round_in[3][1440] , \round_in[3][1439] , 
        \round_in[3][1438] , \round_in[3][1437] , \round_in[3][1436] , 
        \round_in[3][1435] , \round_in[3][1434] , \round_in[3][1433] , 
        \round_in[3][1432] , \round_in[3][1431] , \round_in[3][1430] , 
        \round_in[3][1429] , \round_in[3][1428] , \round_in[3][1427] , 
        \round_in[3][1426] , \round_in[3][1425] , \round_in[3][1424] , 
        \round_in[3][1423] , \round_in[3][1422] , \round_in[3][1421] , 
        \round_in[3][1420] , \round_in[3][1419] , \round_in[3][1418] , 
        \round_in[3][1417] , \round_in[3][1416] , \round_in[3][1415] , 
        \round_in[3][1414] , \round_in[3][1413] , \round_in[3][1412] , 
        \round_in[3][1411] , \round_in[3][1410] , \round_in[3][1409] , 
        \round_in[3][1408] , \round_in[3][1407] , \round_in[3][1406] , 
        \round_in[3][1405] , \round_in[3][1404] , \round_in[3][1403] , 
        \round_in[3][1402] , \round_in[3][1401] , \round_in[3][1400] , 
        \round_in[3][1399] , \round_in[3][1398] , \round_in[3][1397] , 
        \round_in[3][1396] , \round_in[3][1395] , \round_in[3][1394] , 
        \round_in[3][1393] , \round_in[3][1392] , \round_in[3][1391] , 
        \round_in[3][1390] , \round_in[3][1389] , \round_in[3][1388] , 
        \round_in[3][1387] , \round_in[3][1386] , \round_in[3][1385] , 
        \round_in[3][1384] , \round_in[3][1383] , \round_in[3][1382] , 
        \round_in[3][1381] , \round_in[3][1380] , \round_in[3][1379] , 
        \round_in[3][1378] , \round_in[3][1377] , \round_in[3][1376] , 
        \round_in[3][1375] , \round_in[3][1374] , \round_in[3][1373] , 
        \round_in[3][1372] , \round_in[3][1371] , \round_in[3][1370] , 
        \round_in[3][1369] , \round_in[3][1368] , \round_in[3][1367] , 
        \round_in[3][1366] , \round_in[3][1365] , \round_in[3][1364] , 
        \round_in[3][1363] , \round_in[3][1362] , \round_in[3][1361] , 
        \round_in[3][1360] , \round_in[3][1359] , \round_in[3][1358] , 
        \round_in[3][1357] , \round_in[3][1356] , \round_in[3][1355] , 
        \round_in[3][1354] , \round_in[3][1353] , \round_in[3][1352] , 
        \round_in[3][1351] , \round_in[3][1350] , \round_in[3][1349] , 
        \round_in[3][1348] , \round_in[3][1347] , \round_in[3][1346] , 
        \round_in[3][1345] , \round_in[3][1344] , \round_in[3][1343] , 
        \round_in[3][1342] , \round_in[3][1341] , \round_in[3][1340] , 
        \round_in[3][1339] , \round_in[3][1338] , \round_in[3][1337] , 
        \round_in[3][1336] , \round_in[3][1335] , \round_in[3][1334] , 
        \round_in[3][1333] , \round_in[3][1332] , \round_in[3][1331] , 
        \round_in[3][1330] , \round_in[3][1329] , \round_in[3][1328] , 
        \round_in[3][1327] , \round_in[3][1326] , \round_in[3][1325] , 
        \round_in[3][1324] , \round_in[3][1323] , \round_in[3][1322] , 
        \round_in[3][1321] , \round_in[3][1320] , \round_in[3][1319] , 
        \round_in[3][1318] , \round_in[3][1317] , \round_in[3][1316] , 
        \round_in[3][1315] , \round_in[3][1314] , \round_in[3][1313] , 
        \round_in[3][1312] , \round_in[3][1311] , \round_in[3][1310] , 
        \round_in[3][1309] , \round_in[3][1308] , \round_in[3][1307] , 
        \round_in[3][1306] , \round_in[3][1305] , \round_in[3][1304] , 
        \round_in[3][1303] , \round_in[3][1302] , \round_in[3][1301] , 
        \round_in[3][1300] , \round_in[3][1299] , \round_in[3][1298] , 
        \round_in[3][1297] , \round_in[3][1296] , \round_in[3][1295] , 
        \round_in[3][1294] , \round_in[3][1293] , \round_in[3][1292] , 
        \round_in[3][1291] , \round_in[3][1290] , \round_in[3][1289] , 
        \round_in[3][1288] , \round_in[3][1287] , \round_in[3][1286] , 
        \round_in[3][1285] , \round_in[3][1284] , \round_in[3][1283] , 
        \round_in[3][1282] , \round_in[3][1281] , \round_in[3][1280] , 
        \round_in[3][1279] , \round_in[3][1278] , \round_in[3][1277] , 
        \round_in[3][1276] , \round_in[3][1275] , \round_in[3][1274] , 
        \round_in[3][1273] , \round_in[3][1272] , \round_in[3][1271] , 
        \round_in[3][1270] , \round_in[3][1269] , \round_in[3][1268] , 
        \round_in[3][1267] , \round_in[3][1266] , \round_in[3][1265] , 
        \round_in[3][1264] , \round_in[3][1263] , \round_in[3][1262] , 
        \round_in[3][1261] , \round_in[3][1260] , \round_in[3][1259] , 
        \round_in[3][1258] , \round_in[3][1257] , \round_in[3][1256] , 
        \round_in[3][1255] , \round_in[3][1254] , \round_in[3][1253] , 
        \round_in[3][1252] , \round_in[3][1251] , \round_in[3][1250] , 
        \round_in[3][1249] , \round_in[3][1248] , \round_in[3][1247] , 
        \round_in[3][1246] , \round_in[3][1245] , \round_in[3][1244] , 
        \round_in[3][1243] , \round_in[3][1242] , \round_in[3][1241] , 
        \round_in[3][1240] , \round_in[3][1239] , \round_in[3][1238] , 
        \round_in[3][1237] , \round_in[3][1236] , \round_in[3][1235] , 
        \round_in[3][1234] , \round_in[3][1233] , \round_in[3][1232] , 
        \round_in[3][1231] , \round_in[3][1230] , \round_in[3][1229] , 
        \round_in[3][1228] , \round_in[3][1227] , \round_in[3][1226] , 
        \round_in[3][1225] , \round_in[3][1224] , \round_in[3][1223] , 
        \round_in[3][1222] , \round_in[3][1221] , \round_in[3][1220] , 
        \round_in[3][1219] , \round_in[3][1218] , \round_in[3][1217] , 
        \round_in[3][1216] , \round_in[3][1215] , \round_in[3][1214] , 
        \round_in[3][1213] , \round_in[3][1212] , \round_in[3][1211] , 
        \round_in[3][1210] , \round_in[3][1209] , \round_in[3][1208] , 
        \round_in[3][1207] , \round_in[3][1206] , \round_in[3][1205] , 
        \round_in[3][1204] , \round_in[3][1203] , \round_in[3][1202] , 
        \round_in[3][1201] , \round_in[3][1200] , \round_in[3][1199] , 
        \round_in[3][1198] , \round_in[3][1197] , \round_in[3][1196] , 
        \round_in[3][1195] , \round_in[3][1194] , \round_in[3][1193] , 
        \round_in[3][1192] , \round_in[3][1191] , \round_in[3][1190] , 
        \round_in[3][1189] , \round_in[3][1188] , \round_in[3][1187] , 
        \round_in[3][1186] , \round_in[3][1185] , \round_in[3][1184] , 
        \round_in[3][1183] , \round_in[3][1182] , \round_in[3][1181] , 
        \round_in[3][1180] , \round_in[3][1179] , \round_in[3][1178] , 
        \round_in[3][1177] , \round_in[3][1176] , \round_in[3][1175] , 
        \round_in[3][1174] , \round_in[3][1173] , \round_in[3][1172] , 
        \round_in[3][1171] , \round_in[3][1170] , \round_in[3][1169] , 
        \round_in[3][1168] , \round_in[3][1167] , \round_in[3][1166] , 
        \round_in[3][1165] , \round_in[3][1164] , \round_in[3][1163] , 
        \round_in[3][1162] , \round_in[3][1161] , \round_in[3][1160] , 
        \round_in[3][1159] , \round_in[3][1158] , \round_in[3][1157] , 
        \round_in[3][1156] , \round_in[3][1155] , \round_in[3][1154] , 
        \round_in[3][1153] , \round_in[3][1152] , \round_in[3][1151] , 
        \round_in[3][1150] , \round_in[3][1149] , \round_in[3][1148] , 
        \round_in[3][1147] , \round_in[3][1146] , \round_in[3][1145] , 
        \round_in[3][1144] , \round_in[3][1143] , \round_in[3][1142] , 
        \round_in[3][1141] , \round_in[3][1140] , \round_in[3][1139] , 
        \round_in[3][1138] , \round_in[3][1137] , \round_in[3][1136] , 
        \round_in[3][1135] , \round_in[3][1134] , \round_in[3][1133] , 
        \round_in[3][1132] , \round_in[3][1131] , \round_in[3][1130] , 
        \round_in[3][1129] , \round_in[3][1128] , \round_in[3][1127] , 
        \round_in[3][1126] , \round_in[3][1125] , \round_in[3][1124] , 
        \round_in[3][1123] , \round_in[3][1122] , \round_in[3][1121] , 
        \round_in[3][1120] , \round_in[3][1119] , \round_in[3][1118] , 
        \round_in[3][1117] , \round_in[3][1116] , \round_in[3][1115] , 
        \round_in[3][1114] , \round_in[3][1113] , \round_in[3][1112] , 
        \round_in[3][1111] , \round_in[3][1110] , \round_in[3][1109] , 
        \round_in[3][1108] , \round_in[3][1107] , \round_in[3][1106] , 
        \round_in[3][1105] , \round_in[3][1104] , \round_in[3][1103] , 
        \round_in[3][1102] , \round_in[3][1101] , \round_in[3][1100] , 
        \round_in[3][1099] , \round_in[3][1098] , \round_in[3][1097] , 
        \round_in[3][1096] , \round_in[3][1095] , \round_in[3][1094] , 
        \round_in[3][1093] , \round_in[3][1092] , \round_in[3][1091] , 
        \round_in[3][1090] , \round_in[3][1089] , \round_in[3][1088] , 
        \round_in[3][1087] , \round_in[3][1086] , \round_in[3][1085] , 
        \round_in[3][1084] , \round_in[3][1083] , \round_in[3][1082] , 
        \round_in[3][1081] , \round_in[3][1080] , \round_in[3][1079] , 
        \round_in[3][1078] , \round_in[3][1077] , \round_in[3][1076] , 
        \round_in[3][1075] , \round_in[3][1074] , \round_in[3][1073] , 
        \round_in[3][1072] , \round_in[3][1071] , \round_in[3][1070] , 
        \round_in[3][1069] , \round_in[3][1068] , \round_in[3][1067] , 
        \round_in[3][1066] , \round_in[3][1065] , \round_in[3][1064] , 
        \round_in[3][1063] , \round_in[3][1062] , \round_in[3][1061] , 
        \round_in[3][1060] , \round_in[3][1059] , \round_in[3][1058] , 
        \round_in[3][1057] , \round_in[3][1056] , \round_in[3][1055] , 
        \round_in[3][1054] , \round_in[3][1053] , \round_in[3][1052] , 
        \round_in[3][1051] , \round_in[3][1050] , \round_in[3][1049] , 
        \round_in[3][1048] , \round_in[3][1047] , \round_in[3][1046] , 
        \round_in[3][1045] , \round_in[3][1044] , \round_in[3][1043] , 
        \round_in[3][1042] , \round_in[3][1041] , \round_in[3][1040] , 
        \round_in[3][1039] , \round_in[3][1038] , \round_in[3][1037] , 
        \round_in[3][1036] , \round_in[3][1035] , \round_in[3][1034] , 
        \round_in[3][1033] , \round_in[3][1032] , \round_in[3][1031] , 
        \round_in[3][1030] , \round_in[3][1029] , \round_in[3][1028] , 
        \round_in[3][1027] , \round_in[3][1026] , \round_in[3][1025] , 
        \round_in[3][1024] , \round_in[3][1023] , \round_in[3][1022] , 
        \round_in[3][1021] , \round_in[3][1020] , \round_in[3][1019] , 
        \round_in[3][1018] , \round_in[3][1017] , \round_in[3][1016] , 
        \round_in[3][1015] , \round_in[3][1014] , \round_in[3][1013] , 
        \round_in[3][1012] , \round_in[3][1011] , \round_in[3][1010] , 
        \round_in[3][1009] , \round_in[3][1008] , \round_in[3][1007] , 
        \round_in[3][1006] , \round_in[3][1005] , \round_in[3][1004] , 
        \round_in[3][1003] , \round_in[3][1002] , \round_in[3][1001] , 
        \round_in[3][1000] , \round_in[3][999] , \round_in[3][998] , 
        \round_in[3][997] , \round_in[3][996] , \round_in[3][995] , 
        \round_in[3][994] , \round_in[3][993] , \round_in[3][992] , 
        \round_in[3][991] , \round_in[3][990] , \round_in[3][989] , 
        \round_in[3][988] , \round_in[3][987] , \round_in[3][986] , 
        \round_in[3][985] , \round_in[3][984] , \round_in[3][983] , 
        \round_in[3][982] , \round_in[3][981] , \round_in[3][980] , 
        \round_in[3][979] , \round_in[3][978] , \round_in[3][977] , 
        \round_in[3][976] , \round_in[3][975] , \round_in[3][974] , 
        \round_in[3][973] , \round_in[3][972] , \round_in[3][971] , 
        \round_in[3][970] , \round_in[3][969] , \round_in[3][968] , 
        \round_in[3][967] , \round_in[3][966] , \round_in[3][965] , 
        \round_in[3][964] , \round_in[3][963] , \round_in[3][962] , 
        \round_in[3][961] , \round_in[3][960] , \round_in[3][959] , 
        \round_in[3][958] , \round_in[3][957] , \round_in[3][956] , 
        \round_in[3][955] , \round_in[3][954] , \round_in[3][953] , 
        \round_in[3][952] , \round_in[3][951] , \round_in[3][950] , 
        \round_in[3][949] , \round_in[3][948] , \round_in[3][947] , 
        \round_in[3][946] , \round_in[3][945] , \round_in[3][944] , 
        \round_in[3][943] , \round_in[3][942] , \round_in[3][941] , 
        \round_in[3][940] , \round_in[3][939] , \round_in[3][938] , 
        \round_in[3][937] , \round_in[3][936] , \round_in[3][935] , 
        \round_in[3][934] , \round_in[3][933] , \round_in[3][932] , 
        \round_in[3][931] , \round_in[3][930] , \round_in[3][929] , 
        \round_in[3][928] , \round_in[3][927] , \round_in[3][926] , 
        \round_in[3][925] , \round_in[3][924] , \round_in[3][923] , 
        \round_in[3][922] , \round_in[3][921] , \round_in[3][920] , 
        \round_in[3][919] , \round_in[3][918] , \round_in[3][917] , 
        \round_in[3][916] , \round_in[3][915] , \round_in[3][914] , 
        \round_in[3][913] , \round_in[3][912] , \round_in[3][911] , 
        \round_in[3][910] , \round_in[3][909] , \round_in[3][908] , 
        \round_in[3][907] , \round_in[3][906] , \round_in[3][905] , 
        \round_in[3][904] , \round_in[3][903] , \round_in[3][902] , 
        \round_in[3][901] , \round_in[3][900] , \round_in[3][899] , 
        \round_in[3][898] , \round_in[3][897] , \round_in[3][896] , 
        \round_in[3][895] , \round_in[3][894] , \round_in[3][893] , 
        \round_in[3][892] , \round_in[3][891] , \round_in[3][890] , 
        \round_in[3][889] , \round_in[3][888] , \round_in[3][887] , 
        \round_in[3][886] , \round_in[3][885] , \round_in[3][884] , 
        \round_in[3][883] , \round_in[3][882] , \round_in[3][881] , 
        \round_in[3][880] , \round_in[3][879] , \round_in[3][878] , 
        \round_in[3][877] , \round_in[3][876] , \round_in[3][875] , 
        \round_in[3][874] , \round_in[3][873] , \round_in[3][872] , 
        \round_in[3][871] , \round_in[3][870] , \round_in[3][869] , 
        \round_in[3][868] , \round_in[3][867] , \round_in[3][866] , 
        \round_in[3][865] , \round_in[3][864] , \round_in[3][863] , 
        \round_in[3][862] , \round_in[3][861] , \round_in[3][860] , 
        \round_in[3][859] , \round_in[3][858] , \round_in[3][857] , 
        \round_in[3][856] , \round_in[3][855] , \round_in[3][854] , 
        \round_in[3][853] , \round_in[3][852] , \round_in[3][851] , 
        \round_in[3][850] , \round_in[3][849] , \round_in[3][848] , 
        \round_in[3][847] , \round_in[3][846] , \round_in[3][845] , 
        \round_in[3][844] , \round_in[3][843] , \round_in[3][842] , 
        \round_in[3][841] , \round_in[3][840] , \round_in[3][839] , 
        \round_in[3][838] , \round_in[3][837] , \round_in[3][836] , 
        \round_in[3][835] , \round_in[3][834] , \round_in[3][833] , 
        \round_in[3][832] , \round_in[3][831] , \round_in[3][830] , 
        \round_in[3][829] , \round_in[3][828] , \round_in[3][827] , 
        \round_in[3][826] , \round_in[3][825] , \round_in[3][824] , 
        \round_in[3][823] , \round_in[3][822] , \round_in[3][821] , 
        \round_in[3][820] , \round_in[3][819] , \round_in[3][818] , 
        \round_in[3][817] , \round_in[3][816] , \round_in[3][815] , 
        \round_in[3][814] , \round_in[3][813] , \round_in[3][812] , 
        \round_in[3][811] , \round_in[3][810] , \round_in[3][809] , 
        \round_in[3][808] , \round_in[3][807] , \round_in[3][806] , 
        \round_in[3][805] , \round_in[3][804] , \round_in[3][803] , 
        \round_in[3][802] , \round_in[3][801] , \round_in[3][800] , 
        \round_in[3][799] , \round_in[3][798] , \round_in[3][797] , 
        \round_in[3][796] , \round_in[3][795] , \round_in[3][794] , 
        \round_in[3][793] , \round_in[3][792] , \round_in[3][791] , 
        \round_in[3][790] , \round_in[3][789] , \round_in[3][788] , 
        \round_in[3][787] , \round_in[3][786] , \round_in[3][785] , 
        \round_in[3][784] , \round_in[3][783] , \round_in[3][782] , 
        \round_in[3][781] , \round_in[3][780] , \round_in[3][779] , 
        \round_in[3][778] , \round_in[3][777] , \round_in[3][776] , 
        \round_in[3][775] , \round_in[3][774] , \round_in[3][773] , 
        \round_in[3][772] , \round_in[3][771] , \round_in[3][770] , 
        \round_in[3][769] , \round_in[3][768] , \round_in[3][767] , 
        \round_in[3][766] , \round_in[3][765] , \round_in[3][764] , 
        \round_in[3][763] , \round_in[3][762] , \round_in[3][761] , 
        \round_in[3][760] , \round_in[3][759] , \round_in[3][758] , 
        \round_in[3][757] , \round_in[3][756] , \round_in[3][755] , 
        \round_in[3][754] , \round_in[3][753] , \round_in[3][752] , 
        \round_in[3][751] , \round_in[3][750] , \round_in[3][749] , 
        \round_in[3][748] , \round_in[3][747] , \round_in[3][746] , 
        \round_in[3][745] , \round_in[3][744] , \round_in[3][743] , 
        \round_in[3][742] , \round_in[3][741] , \round_in[3][740] , 
        \round_in[3][739] , \round_in[3][738] , \round_in[3][737] , 
        \round_in[3][736] , \round_in[3][735] , \round_in[3][734] , 
        \round_in[3][733] , \round_in[3][732] , \round_in[3][731] , 
        \round_in[3][730] , \round_in[3][729] , \round_in[3][728] , 
        \round_in[3][727] , \round_in[3][726] , \round_in[3][725] , 
        \round_in[3][724] , \round_in[3][723] , \round_in[3][722] , 
        \round_in[3][721] , \round_in[3][720] , \round_in[3][719] , 
        \round_in[3][718] , \round_in[3][717] , \round_in[3][716] , 
        \round_in[3][715] , \round_in[3][714] , \round_in[3][713] , 
        \round_in[3][712] , \round_in[3][711] , \round_in[3][710] , 
        \round_in[3][709] , \round_in[3][708] , \round_in[3][707] , 
        \round_in[3][706] , \round_in[3][705] , \round_in[3][704] , 
        \round_in[3][703] , \round_in[3][702] , \round_in[3][701] , 
        \round_in[3][700] , \round_in[3][699] , \round_in[3][698] , 
        \round_in[3][697] , \round_in[3][696] , \round_in[3][695] , 
        \round_in[3][694] , \round_in[3][693] , \round_in[3][692] , 
        \round_in[3][691] , \round_in[3][690] , \round_in[3][689] , 
        \round_in[3][688] , \round_in[3][687] , \round_in[3][686] , 
        \round_in[3][685] , \round_in[3][684] , \round_in[3][683] , 
        \round_in[3][682] , \round_in[3][681] , \round_in[3][680] , 
        \round_in[3][679] , \round_in[3][678] , \round_in[3][677] , 
        \round_in[3][676] , \round_in[3][675] , \round_in[3][674] , 
        \round_in[3][673] , \round_in[3][672] , \round_in[3][671] , 
        \round_in[3][670] , \round_in[3][669] , \round_in[3][668] , 
        \round_in[3][667] , \round_in[3][666] , \round_in[3][665] , 
        \round_in[3][664] , \round_in[3][663] , \round_in[3][662] , 
        \round_in[3][661] , \round_in[3][660] , \round_in[3][659] , 
        \round_in[3][658] , \round_in[3][657] , \round_in[3][656] , 
        \round_in[3][655] , \round_in[3][654] , \round_in[3][653] , 
        \round_in[3][652] , \round_in[3][651] , \round_in[3][650] , 
        \round_in[3][649] , \round_in[3][648] , \round_in[3][647] , 
        \round_in[3][646] , \round_in[3][645] , \round_in[3][644] , 
        \round_in[3][643] , \round_in[3][642] , \round_in[3][641] , 
        \round_in[3][640] , \round_in[3][639] , \round_in[3][638] , 
        \round_in[3][637] , \round_in[3][636] , \round_in[3][635] , 
        \round_in[3][634] , \round_in[3][633] , \round_in[3][632] , 
        \round_in[3][631] , \round_in[3][630] , \round_in[3][629] , 
        \round_in[3][628] , \round_in[3][627] , \round_in[3][626] , 
        \round_in[3][625] , \round_in[3][624] , \round_in[3][623] , 
        \round_in[3][622] , \round_in[3][621] , \round_in[3][620] , 
        \round_in[3][619] , \round_in[3][618] , \round_in[3][617] , 
        \round_in[3][616] , \round_in[3][615] , \round_in[3][614] , 
        \round_in[3][613] , \round_in[3][612] , \round_in[3][611] , 
        \round_in[3][610] , \round_in[3][609] , \round_in[3][608] , 
        \round_in[3][607] , \round_in[3][606] , \round_in[3][605] , 
        \round_in[3][604] , \round_in[3][603] , \round_in[3][602] , 
        \round_in[3][601] , \round_in[3][600] , \round_in[3][599] , 
        \round_in[3][598] , \round_in[3][597] , \round_in[3][596] , 
        \round_in[3][595] , \round_in[3][594] , \round_in[3][593] , 
        \round_in[3][592] , \round_in[3][591] , \round_in[3][590] , 
        \round_in[3][589] , \round_in[3][588] , \round_in[3][587] , 
        \round_in[3][586] , \round_in[3][585] , \round_in[3][584] , 
        \round_in[3][583] , \round_in[3][582] , \round_in[3][581] , 
        \round_in[3][580] , \round_in[3][579] , \round_in[3][578] , 
        \round_in[3][577] , \round_in[3][576] , \round_in[3][575] , 
        \round_in[3][574] , \round_in[3][573] , \round_in[3][572] , 
        \round_in[3][571] , \round_in[3][570] , \round_in[3][569] , 
        \round_in[3][568] , \round_in[3][567] , \round_in[3][566] , 
        \round_in[3][565] , \round_in[3][564] , \round_in[3][563] , 
        \round_in[3][562] , \round_in[3][561] , \round_in[3][560] , 
        \round_in[3][559] , \round_in[3][558] , \round_in[3][557] , 
        \round_in[3][556] , \round_in[3][555] , \round_in[3][554] , 
        \round_in[3][553] , \round_in[3][552] , \round_in[3][551] , 
        \round_in[3][550] , \round_in[3][549] , \round_in[3][548] , 
        \round_in[3][547] , \round_in[3][546] , \round_in[3][545] , 
        \round_in[3][544] , \round_in[3][543] , \round_in[3][542] , 
        \round_in[3][541] , \round_in[3][540] , \round_in[3][539] , 
        \round_in[3][538] , \round_in[3][537] , \round_in[3][536] , 
        \round_in[3][535] , \round_in[3][534] , \round_in[3][533] , 
        \round_in[3][532] , \round_in[3][531] , \round_in[3][530] , 
        \round_in[3][529] , \round_in[3][528] , \round_in[3][527] , 
        \round_in[3][526] , \round_in[3][525] , \round_in[3][524] , 
        \round_in[3][523] , \round_in[3][522] , \round_in[3][521] , 
        \round_in[3][520] , \round_in[3][519] , \round_in[3][518] , 
        \round_in[3][517] , \round_in[3][516] , \round_in[3][515] , 
        \round_in[3][514] , \round_in[3][513] , \round_in[3][512] , 
        \round_in[3][511] , \round_in[3][510] , \round_in[3][509] , 
        \round_in[3][508] , \round_in[3][507] , \round_in[3][506] , 
        \round_in[3][505] , \round_in[3][504] , \round_in[3][503] , 
        \round_in[3][502] , \round_in[3][501] , \round_in[3][500] , 
        \round_in[3][499] , \round_in[3][498] , \round_in[3][497] , 
        \round_in[3][496] , \round_in[3][495] , \round_in[3][494] , 
        \round_in[3][493] , \round_in[3][492] , \round_in[3][491] , 
        \round_in[3][490] , \round_in[3][489] , \round_in[3][488] , 
        \round_in[3][487] , \round_in[3][486] , \round_in[3][485] , 
        \round_in[3][484] , \round_in[3][483] , \round_in[3][482] , 
        \round_in[3][481] , \round_in[3][480] , \round_in[3][479] , 
        \round_in[3][478] , \round_in[3][477] , \round_in[3][476] , 
        \round_in[3][475] , \round_in[3][474] , \round_in[3][473] , 
        \round_in[3][472] , \round_in[3][471] , \round_in[3][470] , 
        \round_in[3][469] , \round_in[3][468] , \round_in[3][467] , 
        \round_in[3][466] , \round_in[3][465] , \round_in[3][464] , 
        \round_in[3][463] , \round_in[3][462] , \round_in[3][461] , 
        \round_in[3][460] , \round_in[3][459] , \round_in[3][458] , 
        \round_in[3][457] , \round_in[3][456] , \round_in[3][455] , 
        \round_in[3][454] , \round_in[3][453] , \round_in[3][452] , 
        \round_in[3][451] , \round_in[3][450] , \round_in[3][449] , 
        \round_in[3][448] , \round_in[3][447] , \round_in[3][446] , 
        \round_in[3][445] , \round_in[3][444] , \round_in[3][443] , 
        \round_in[3][442] , \round_in[3][441] , \round_in[3][440] , 
        \round_in[3][439] , \round_in[3][438] , \round_in[3][437] , 
        \round_in[3][436] , \round_in[3][435] , \round_in[3][434] , 
        \round_in[3][433] , \round_in[3][432] , \round_in[3][431] , 
        \round_in[3][430] , \round_in[3][429] , \round_in[3][428] , 
        \round_in[3][427] , \round_in[3][426] , \round_in[3][425] , 
        \round_in[3][424] , \round_in[3][423] , \round_in[3][422] , 
        \round_in[3][421] , \round_in[3][420] , \round_in[3][419] , 
        \round_in[3][418] , \round_in[3][417] , \round_in[3][416] , 
        \round_in[3][415] , \round_in[3][414] , \round_in[3][413] , 
        \round_in[3][412] , \round_in[3][411] , \round_in[3][410] , 
        \round_in[3][409] , \round_in[3][408] , \round_in[3][407] , 
        \round_in[3][406] , \round_in[3][405] , \round_in[3][404] , 
        \round_in[3][403] , \round_in[3][402] , \round_in[3][401] , 
        \round_in[3][400] , \round_in[3][399] , \round_in[3][398] , 
        \round_in[3][397] , \round_in[3][396] , \round_in[3][395] , 
        \round_in[3][394] , \round_in[3][393] , \round_in[3][392] , 
        \round_in[3][391] , \round_in[3][390] , \round_in[3][389] , 
        \round_in[3][388] , \round_in[3][387] , \round_in[3][386] , 
        \round_in[3][385] , \round_in[3][384] , \round_in[3][383] , 
        \round_in[3][382] , \round_in[3][381] , \round_in[3][380] , 
        \round_in[3][379] , \round_in[3][378] , \round_in[3][377] , 
        \round_in[3][376] , \round_in[3][375] , \round_in[3][374] , 
        \round_in[3][373] , \round_in[3][372] , \round_in[3][371] , 
        \round_in[3][370] , \round_in[3][369] , \round_in[3][368] , 
        \round_in[3][367] , \round_in[3][366] , \round_in[3][365] , 
        \round_in[3][364] , \round_in[3][363] , \round_in[3][362] , 
        \round_in[3][361] , \round_in[3][360] , \round_in[3][359] , 
        \round_in[3][358] , \round_in[3][357] , \round_in[3][356] , 
        \round_in[3][355] , \round_in[3][354] , \round_in[3][353] , 
        \round_in[3][352] , \round_in[3][351] , \round_in[3][350] , 
        \round_in[3][349] , \round_in[3][348] , \round_in[3][347] , 
        \round_in[3][346] , \round_in[3][345] , \round_in[3][344] , 
        \round_in[3][343] , \round_in[3][342] , \round_in[3][341] , 
        \round_in[3][340] , \round_in[3][339] , \round_in[3][338] , 
        \round_in[3][337] , \round_in[3][336] , \round_in[3][335] , 
        \round_in[3][334] , \round_in[3][333] , \round_in[3][332] , 
        \round_in[3][331] , \round_in[3][330] , \round_in[3][329] , 
        \round_in[3][328] , \round_in[3][327] , \round_in[3][326] , 
        \round_in[3][325] , \round_in[3][324] , \round_in[3][323] , 
        \round_in[3][322] , \round_in[3][321] , \round_in[3][320] , 
        \round_in[3][319] , \round_in[3][318] , \round_in[3][317] , 
        \round_in[3][316] , \round_in[3][315] , \round_in[3][314] , 
        \round_in[3][313] , \round_in[3][312] , \round_in[3][311] , 
        \round_in[3][310] , \round_in[3][309] , \round_in[3][308] , 
        \round_in[3][307] , \round_in[3][306] , \round_in[3][305] , 
        \round_in[3][304] , \round_in[3][303] , \round_in[3][302] , 
        \round_in[3][301] , \round_in[3][300] , \round_in[3][299] , 
        \round_in[3][298] , \round_in[3][297] , \round_in[3][296] , 
        \round_in[3][295] , \round_in[3][294] , \round_in[3][293] , 
        \round_in[3][292] , \round_in[3][291] , \round_in[3][290] , 
        \round_in[3][289] , \round_in[3][288] , \round_in[3][287] , 
        \round_in[3][286] , \round_in[3][285] , \round_in[3][284] , 
        \round_in[3][283] , \round_in[3][282] , \round_in[3][281] , 
        \round_in[3][280] , \round_in[3][279] , \round_in[3][278] , 
        \round_in[3][277] , \round_in[3][276] , \round_in[3][275] , 
        \round_in[3][274] , \round_in[3][273] , \round_in[3][272] , 
        \round_in[3][271] , \round_in[3][270] , \round_in[3][269] , 
        \round_in[3][268] , \round_in[3][267] , \round_in[3][266] , 
        \round_in[3][265] , \round_in[3][264] , \round_in[3][263] , 
        \round_in[3][262] , \round_in[3][261] , \round_in[3][260] , 
        \round_in[3][259] , \round_in[3][258] , \round_in[3][257] , 
        \round_in[3][256] , \round_in[3][255] , \round_in[3][254] , 
        \round_in[3][253] , \round_in[3][252] , \round_in[3][251] , 
        \round_in[3][250] , \round_in[3][249] , \round_in[3][248] , 
        \round_in[3][247] , \round_in[3][246] , \round_in[3][245] , 
        \round_in[3][244] , \round_in[3][243] , \round_in[3][242] , 
        \round_in[3][241] , \round_in[3][240] , \round_in[3][239] , 
        \round_in[3][238] , \round_in[3][237] , \round_in[3][236] , 
        \round_in[3][235] , \round_in[3][234] , \round_in[3][233] , 
        \round_in[3][232] , \round_in[3][231] , \round_in[3][230] , 
        \round_in[3][229] , \round_in[3][228] , \round_in[3][227] , 
        \round_in[3][226] , \round_in[3][225] , \round_in[3][224] , 
        \round_in[3][223] , \round_in[3][222] , \round_in[3][221] , 
        \round_in[3][220] , \round_in[3][219] , \round_in[3][218] , 
        \round_in[3][217] , \round_in[3][216] , \round_in[3][215] , 
        \round_in[3][214] , \round_in[3][213] , \round_in[3][212] , 
        \round_in[3][211] , \round_in[3][210] , \round_in[3][209] , 
        \round_in[3][208] , \round_in[3][207] , \round_in[3][206] , 
        \round_in[3][205] , \round_in[3][204] , \round_in[3][203] , 
        \round_in[3][202] , \round_in[3][201] , \round_in[3][200] , 
        \round_in[3][199] , \round_in[3][198] , \round_in[3][197] , 
        \round_in[3][196] , \round_in[3][195] , \round_in[3][194] , 
        \round_in[3][193] , \round_in[3][192] , \round_in[3][191] , 
        \round_in[3][190] , \round_in[3][189] , \round_in[3][188] , 
        \round_in[3][187] , \round_in[3][186] , \round_in[3][185] , 
        \round_in[3][184] , \round_in[3][183] , \round_in[3][182] , 
        \round_in[3][181] , \round_in[3][180] , \round_in[3][179] , 
        \round_in[3][178] , \round_in[3][177] , \round_in[3][176] , 
        \round_in[3][175] , \round_in[3][174] , \round_in[3][173] , 
        \round_in[3][172] , \round_in[3][171] , \round_in[3][170] , 
        \round_in[3][169] , \round_in[3][168] , \round_in[3][167] , 
        \round_in[3][166] , \round_in[3][165] , \round_in[3][164] , 
        \round_in[3][163] , \round_in[3][162] , \round_in[3][161] , 
        \round_in[3][160] , \round_in[3][159] , \round_in[3][158] , 
        \round_in[3][157] , \round_in[3][156] , \round_in[3][155] , 
        \round_in[3][154] , \round_in[3][153] , \round_in[3][152] , 
        \round_in[3][151] , \round_in[3][150] , \round_in[3][149] , 
        \round_in[3][148] , \round_in[3][147] , \round_in[3][146] , 
        \round_in[3][145] , \round_in[3][144] , \round_in[3][143] , 
        \round_in[3][142] , \round_in[3][141] , \round_in[3][140] , 
        \round_in[3][139] , \round_in[3][138] , \round_in[3][137] , 
        \round_in[3][136] , \round_in[3][135] , \round_in[3][134] , 
        \round_in[3][133] , \round_in[3][132] , \round_in[3][131] , 
        \round_in[3][130] , \round_in[3][129] , \round_in[3][128] , 
        \round_in[3][127] , \round_in[3][126] , \round_in[3][125] , 
        \round_in[3][124] , \round_in[3][123] , \round_in[3][122] , 
        \round_in[3][121] , \round_in[3][120] , \round_in[3][119] , 
        \round_in[3][118] , \round_in[3][117] , \round_in[3][116] , 
        \round_in[3][115] , \round_in[3][114] , \round_in[3][113] , 
        \round_in[3][112] , \round_in[3][111] , \round_in[3][110] , 
        \round_in[3][109] , \round_in[3][108] , \round_in[3][107] , 
        \round_in[3][106] , \round_in[3][105] , \round_in[3][104] , 
        \round_in[3][103] , \round_in[3][102] , \round_in[3][101] , 
        \round_in[3][100] , \round_in[3][99] , \round_in[3][98] , 
        \round_in[3][97] , \round_in[3][96] , \round_in[3][95] , 
        \round_in[3][94] , \round_in[3][93] , \round_in[3][92] , 
        \round_in[3][91] , \round_in[3][90] , \round_in[3][89] , 
        \round_in[3][88] , \round_in[3][87] , \round_in[3][86] , 
        \round_in[3][85] , \round_in[3][84] , \round_in[3][83] , 
        \round_in[3][82] , \round_in[3][81] , \round_in[3][80] , 
        \round_in[3][79] , \round_in[3][78] , \round_in[3][77] , 
        \round_in[3][76] , \round_in[3][75] , \round_in[3][74] , 
        \round_in[3][73] , \round_in[3][72] , \round_in[3][71] , 
        \round_in[3][70] , \round_in[3][69] , \round_in[3][68] , 
        \round_in[3][67] , \round_in[3][66] , \round_in[3][65] , 
        \round_in[3][64] , \round_in[3][63] , \round_in[3][62] , 
        \round_in[3][61] , \round_in[3][60] , \round_in[3][59] , 
        \round_in[3][58] , \round_in[3][57] , \round_in[3][56] , 
        \round_in[3][55] , \round_in[3][54] , \round_in[3][53] , 
        \round_in[3][52] , \round_in[3][51] , \round_in[3][50] , 
        \round_in[3][49] , \round_in[3][48] , \round_in[3][47] , 
        \round_in[3][46] , \round_in[3][45] , \round_in[3][44] , 
        \round_in[3][43] , \round_in[3][42] , \round_in[3][41] , 
        \round_in[3][40] , \round_in[3][39] , \round_in[3][38] , 
        \round_in[3][37] , \round_in[3][36] , \round_in[3][35] , 
        \round_in[3][34] , \round_in[3][33] , \round_in[3][32] , 
        \round_in[3][31] , \round_in[3][30] , \round_in[3][29] , 
        \round_in[3][28] , \round_in[3][27] , \round_in[3][26] , 
        \round_in[3][25] , \round_in[3][24] , \round_in[3][23] , 
        \round_in[3][22] , \round_in[3][21] , \round_in[3][20] , 
        \round_in[3][19] , \round_in[3][18] , \round_in[3][17] , 
        \round_in[3][16] , \round_in[3][15] , \round_in[3][14] , 
        \round_in[3][13] , \round_in[3][12] , \round_in[3][11] , 
        \round_in[3][10] , \round_in[3][9] , \round_in[3][8] , 
        \round_in[3][7] , \round_in[3][6] , \round_in[3][5] , \round_in[3][4] , 
        \round_in[3][3] , \round_in[3][2] , \round_in[3][1] , \round_in[3][0] }), .round_const({\rc[3][63] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        \rc[3][31] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[3][15] , 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \rc[3][3] , 1'b0, 
        \rc[3][1] , \RCONST[3].rconst_/N10 }), .out(out) );
  DFF init_reg ( .D(n1614), .CLK(clk), .RST(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(N6), .CLK(clk), .RST(1'b0), .Q(rc_i[0]) );
  DFF \rc_i_reg[1]  ( .D(N7), .CLK(clk), .RST(1'b0), .Q(rc_i[1]) );
  DFF \rc_i_reg[2]  ( .D(N8), .CLK(clk), .RST(1'b0), .Q(rc_i[2]) );
  DFF \rc_i_reg[3]  ( .D(N9), .CLK(clk), .RST(1'b0), .Q(rc_i[3]) );
  DFF \rc_i_reg[4]  ( .D(N10), .CLK(clk), .RST(1'b0), .Q(rc_i[4]) );
  DFF \rc_i_reg[5]  ( .D(N11), .CLK(clk), .RST(1'b0), .Q(rc_i[5]) );
  DFF \round_reg_reg[0]  ( .D(N12), .CLK(clk), .RST(1'b0), .Q(round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(N13), .CLK(clk), .RST(1'b0), .Q(round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(N14), .CLK(clk), .RST(1'b0), .Q(round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(N15), .CLK(clk), .RST(1'b0), .Q(round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(N16), .CLK(clk), .RST(1'b0), .Q(round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(N17), .CLK(clk), .RST(1'b0), .Q(round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(N18), .CLK(clk), .RST(1'b0), .Q(round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(N19), .CLK(clk), .RST(1'b0), .Q(round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(N20), .CLK(clk), .RST(1'b0), .Q(round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(N21), .CLK(clk), .RST(1'b0), .Q(round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(N22), .CLK(clk), .RST(1'b0), .Q(round_reg[10])
         );
  DFF \round_reg_reg[11]  ( .D(N23), .CLK(clk), .RST(1'b0), .Q(round_reg[11])
         );
  DFF \round_reg_reg[12]  ( .D(N24), .CLK(clk), .RST(1'b0), .Q(round_reg[12])
         );
  DFF \round_reg_reg[13]  ( .D(N25), .CLK(clk), .RST(1'b0), .Q(round_reg[13])
         );
  DFF \round_reg_reg[14]  ( .D(N26), .CLK(clk), .RST(1'b0), .Q(round_reg[14])
         );
  DFF \round_reg_reg[15]  ( .D(N27), .CLK(clk), .RST(1'b0), .Q(round_reg[15])
         );
  DFF \round_reg_reg[16]  ( .D(N28), .CLK(clk), .RST(1'b0), .Q(round_reg[16])
         );
  DFF \round_reg_reg[17]  ( .D(N29), .CLK(clk), .RST(1'b0), .Q(round_reg[17])
         );
  DFF \round_reg_reg[18]  ( .D(N30), .CLK(clk), .RST(1'b0), .Q(round_reg[18])
         );
  DFF \round_reg_reg[19]  ( .D(N31), .CLK(clk), .RST(1'b0), .Q(round_reg[19])
         );
  DFF \round_reg_reg[20]  ( .D(N32), .CLK(clk), .RST(1'b0), .Q(round_reg[20])
         );
  DFF \round_reg_reg[21]  ( .D(N33), .CLK(clk), .RST(1'b0), .Q(round_reg[21])
         );
  DFF \round_reg_reg[22]  ( .D(N34), .CLK(clk), .RST(1'b0), .Q(round_reg[22])
         );
  DFF \round_reg_reg[23]  ( .D(N35), .CLK(clk), .RST(1'b0), .Q(round_reg[23])
         );
  DFF \round_reg_reg[24]  ( .D(N36), .CLK(clk), .RST(1'b0), .Q(round_reg[24])
         );
  DFF \round_reg_reg[25]  ( .D(N37), .CLK(clk), .RST(1'b0), .Q(round_reg[25])
         );
  DFF \round_reg_reg[26]  ( .D(N38), .CLK(clk), .RST(1'b0), .Q(round_reg[26])
         );
  DFF \round_reg_reg[27]  ( .D(N39), .CLK(clk), .RST(1'b0), .Q(round_reg[27])
         );
  DFF \round_reg_reg[28]  ( .D(N40), .CLK(clk), .RST(1'b0), .Q(round_reg[28])
         );
  DFF \round_reg_reg[29]  ( .D(N41), .CLK(clk), .RST(1'b0), .Q(round_reg[29])
         );
  DFF \round_reg_reg[30]  ( .D(N42), .CLK(clk), .RST(1'b0), .Q(round_reg[30])
         );
  DFF \round_reg_reg[31]  ( .D(N43), .CLK(clk), .RST(1'b0), .Q(round_reg[31])
         );
  DFF \round_reg_reg[32]  ( .D(N44), .CLK(clk), .RST(1'b0), .Q(round_reg[32])
         );
  DFF \round_reg_reg[33]  ( .D(N45), .CLK(clk), .RST(1'b0), .Q(round_reg[33])
         );
  DFF \round_reg_reg[34]  ( .D(N46), .CLK(clk), .RST(1'b0), .Q(round_reg[34])
         );
  DFF \round_reg_reg[35]  ( .D(N47), .CLK(clk), .RST(1'b0), .Q(round_reg[35])
         );
  DFF \round_reg_reg[36]  ( .D(N48), .CLK(clk), .RST(1'b0), .Q(round_reg[36])
         );
  DFF \round_reg_reg[37]  ( .D(N49), .CLK(clk), .RST(1'b0), .Q(round_reg[37])
         );
  DFF \round_reg_reg[38]  ( .D(N50), .CLK(clk), .RST(1'b0), .Q(round_reg[38])
         );
  DFF \round_reg_reg[39]  ( .D(N51), .CLK(clk), .RST(1'b0), .Q(round_reg[39])
         );
  DFF \round_reg_reg[40]  ( .D(N52), .CLK(clk), .RST(1'b0), .Q(round_reg[40])
         );
  DFF \round_reg_reg[41]  ( .D(N53), .CLK(clk), .RST(1'b0), .Q(round_reg[41])
         );
  DFF \round_reg_reg[42]  ( .D(N54), .CLK(clk), .RST(1'b0), .Q(round_reg[42])
         );
  DFF \round_reg_reg[43]  ( .D(N55), .CLK(clk), .RST(1'b0), .Q(round_reg[43])
         );
  DFF \round_reg_reg[44]  ( .D(N56), .CLK(clk), .RST(1'b0), .Q(round_reg[44])
         );
  DFF \round_reg_reg[45]  ( .D(N57), .CLK(clk), .RST(1'b0), .Q(round_reg[45])
         );
  DFF \round_reg_reg[46]  ( .D(N58), .CLK(clk), .RST(1'b0), .Q(round_reg[46])
         );
  DFF \round_reg_reg[47]  ( .D(N59), .CLK(clk), .RST(1'b0), .Q(round_reg[47])
         );
  DFF \round_reg_reg[48]  ( .D(N60), .CLK(clk), .RST(1'b0), .Q(round_reg[48])
         );
  DFF \round_reg_reg[49]  ( .D(N61), .CLK(clk), .RST(1'b0), .Q(round_reg[49])
         );
  DFF \round_reg_reg[50]  ( .D(N62), .CLK(clk), .RST(1'b0), .Q(round_reg[50])
         );
  DFF \round_reg_reg[51]  ( .D(N63), .CLK(clk), .RST(1'b0), .Q(round_reg[51])
         );
  DFF \round_reg_reg[52]  ( .D(N64), .CLK(clk), .RST(1'b0), .Q(round_reg[52])
         );
  DFF \round_reg_reg[53]  ( .D(N65), .CLK(clk), .RST(1'b0), .Q(round_reg[53])
         );
  DFF \round_reg_reg[54]  ( .D(N66), .CLK(clk), .RST(1'b0), .Q(round_reg[54])
         );
  DFF \round_reg_reg[55]  ( .D(N67), .CLK(clk), .RST(1'b0), .Q(round_reg[55])
         );
  DFF \round_reg_reg[56]  ( .D(N68), .CLK(clk), .RST(1'b0), .Q(round_reg[56])
         );
  DFF \round_reg_reg[57]  ( .D(N69), .CLK(clk), .RST(1'b0), .Q(round_reg[57])
         );
  DFF \round_reg_reg[58]  ( .D(N70), .CLK(clk), .RST(1'b0), .Q(round_reg[58])
         );
  DFF \round_reg_reg[59]  ( .D(N71), .CLK(clk), .RST(1'b0), .Q(round_reg[59])
         );
  DFF \round_reg_reg[60]  ( .D(N72), .CLK(clk), .RST(1'b0), .Q(round_reg[60])
         );
  DFF \round_reg_reg[61]  ( .D(N73), .CLK(clk), .RST(1'b0), .Q(round_reg[61])
         );
  DFF \round_reg_reg[62]  ( .D(N74), .CLK(clk), .RST(1'b0), .Q(round_reg[62])
         );
  DFF \round_reg_reg[63]  ( .D(N75), .CLK(clk), .RST(1'b0), .Q(round_reg[63])
         );
  DFF \round_reg_reg[64]  ( .D(N76), .CLK(clk), .RST(1'b0), .Q(round_reg[64])
         );
  DFF \round_reg_reg[65]  ( .D(N77), .CLK(clk), .RST(1'b0), .Q(round_reg[65])
         );
  DFF \round_reg_reg[66]  ( .D(N78), .CLK(clk), .RST(1'b0), .Q(round_reg[66])
         );
  DFF \round_reg_reg[67]  ( .D(N79), .CLK(clk), .RST(1'b0), .Q(round_reg[67])
         );
  DFF \round_reg_reg[68]  ( .D(N80), .CLK(clk), .RST(1'b0), .Q(round_reg[68])
         );
  DFF \round_reg_reg[69]  ( .D(N81), .CLK(clk), .RST(1'b0), .Q(round_reg[69])
         );
  DFF \round_reg_reg[70]  ( .D(N82), .CLK(clk), .RST(1'b0), .Q(round_reg[70])
         );
  DFF \round_reg_reg[71]  ( .D(N83), .CLK(clk), .RST(1'b0), .Q(round_reg[71])
         );
  DFF \round_reg_reg[72]  ( .D(N84), .CLK(clk), .RST(1'b0), .Q(round_reg[72])
         );
  DFF \round_reg_reg[73]  ( .D(N85), .CLK(clk), .RST(1'b0), .Q(round_reg[73])
         );
  DFF \round_reg_reg[74]  ( .D(N86), .CLK(clk), .RST(1'b0), .Q(round_reg[74])
         );
  DFF \round_reg_reg[75]  ( .D(N87), .CLK(clk), .RST(1'b0), .Q(round_reg[75])
         );
  DFF \round_reg_reg[76]  ( .D(N88), .CLK(clk), .RST(1'b0), .Q(round_reg[76])
         );
  DFF \round_reg_reg[77]  ( .D(N89), .CLK(clk), .RST(1'b0), .Q(round_reg[77])
         );
  DFF \round_reg_reg[78]  ( .D(N90), .CLK(clk), .RST(1'b0), .Q(round_reg[78])
         );
  DFF \round_reg_reg[79]  ( .D(N91), .CLK(clk), .RST(1'b0), .Q(round_reg[79])
         );
  DFF \round_reg_reg[80]  ( .D(N92), .CLK(clk), .RST(1'b0), .Q(round_reg[80])
         );
  DFF \round_reg_reg[81]  ( .D(N93), .CLK(clk), .RST(1'b0), .Q(round_reg[81])
         );
  DFF \round_reg_reg[82]  ( .D(N94), .CLK(clk), .RST(1'b0), .Q(round_reg[82])
         );
  DFF \round_reg_reg[83]  ( .D(N95), .CLK(clk), .RST(1'b0), .Q(round_reg[83])
         );
  DFF \round_reg_reg[84]  ( .D(N96), .CLK(clk), .RST(1'b0), .Q(round_reg[84])
         );
  DFF \round_reg_reg[85]  ( .D(N97), .CLK(clk), .RST(1'b0), .Q(round_reg[85])
         );
  DFF \round_reg_reg[86]  ( .D(N98), .CLK(clk), .RST(1'b0), .Q(round_reg[86])
         );
  DFF \round_reg_reg[87]  ( .D(N99), .CLK(clk), .RST(1'b0), .Q(round_reg[87])
         );
  DFF \round_reg_reg[88]  ( .D(N100), .CLK(clk), .RST(1'b0), .Q(round_reg[88])
         );
  DFF \round_reg_reg[89]  ( .D(N101), .CLK(clk), .RST(1'b0), .Q(round_reg[89])
         );
  DFF \round_reg_reg[90]  ( .D(N102), .CLK(clk), .RST(1'b0), .Q(round_reg[90])
         );
  DFF \round_reg_reg[91]  ( .D(N103), .CLK(clk), .RST(1'b0), .Q(round_reg[91])
         );
  DFF \round_reg_reg[92]  ( .D(N104), .CLK(clk), .RST(1'b0), .Q(round_reg[92])
         );
  DFF \round_reg_reg[93]  ( .D(N105), .CLK(clk), .RST(1'b0), .Q(round_reg[93])
         );
  DFF \round_reg_reg[94]  ( .D(N106), .CLK(clk), .RST(1'b0), .Q(round_reg[94])
         );
  DFF \round_reg_reg[95]  ( .D(N107), .CLK(clk), .RST(1'b0), .Q(round_reg[95])
         );
  DFF \round_reg_reg[96]  ( .D(N108), .CLK(clk), .RST(1'b0), .Q(round_reg[96])
         );
  DFF \round_reg_reg[97]  ( .D(N109), .CLK(clk), .RST(1'b0), .Q(round_reg[97])
         );
  DFF \round_reg_reg[98]  ( .D(N110), .CLK(clk), .RST(1'b0), .Q(round_reg[98])
         );
  DFF \round_reg_reg[99]  ( .D(N111), .CLK(clk), .RST(1'b0), .Q(round_reg[99])
         );
  DFF \round_reg_reg[100]  ( .D(N112), .CLK(clk), .RST(1'b0), .Q(
        round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(N113), .CLK(clk), .RST(1'b0), .Q(
        round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(N114), .CLK(clk), .RST(1'b0), .Q(
        round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(N115), .CLK(clk), .RST(1'b0), .Q(
        round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(N116), .CLK(clk), .RST(1'b0), .Q(
        round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(N117), .CLK(clk), .RST(1'b0), .Q(
        round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(N118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(N119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(N120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(N121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(N122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(N123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(N124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(N125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(N126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(N127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(N128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(N129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(N130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(N131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(N132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(N133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(N134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(N135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(N136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(N137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(N138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(N139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(N140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(N141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(N142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(N143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(N144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(N145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(N146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(N147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(N148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(N149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(N150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(N151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(N152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(N153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(N154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(N155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(N156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(N157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(N158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(N159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(N160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(N161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(N162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(N163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(N164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(N165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(N166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(N167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(N168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(N169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(N170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(N171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(N172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(N173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(N174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(N175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(N176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(N177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(N178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(N179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(N180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(N181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(N182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(N183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(N184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(N185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(N186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(N187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(N188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(N189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(N190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(N191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(N192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(N193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(N194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(N195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(N196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(N197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(N198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(N199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(N200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(N201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(N202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(N203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(N204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(N205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(N206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(N207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(N208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(N209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(N210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(N211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(N212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(N213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(N214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(N215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(N216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(N217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(N218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(N219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(N220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(N221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(N222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(N223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(N224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(N225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(N226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(N227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(N228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(N229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(N230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(N231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(N232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(N233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(N234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(N235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(N236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(N237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(N238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(N239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(N240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(N241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(N242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(N243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(N244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(N245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(N246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(N247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(N248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(N249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(N250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(N251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(N252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(N253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(N254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(N255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(N256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(N257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(N258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(N259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(N260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(N261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(N262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(N263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(N264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(N265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(N266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(N267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(N268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(N269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(N270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(N271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(N272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(N273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(N274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(N275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(N276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(N277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(N278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(N279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(N280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(N281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(N282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(N283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(N284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(N285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(N286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(N287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(N288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(N289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(N290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(N291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(N292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(N293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(N294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(N295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(N296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(N297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(N298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(N299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(N300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(N301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(N302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(N303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(N304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(N305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(N306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(N307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(N308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(N309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(N310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(N311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(N312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(N313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(N314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(N315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(N316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(N317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(N318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(N319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(N320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(N321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(N322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(N323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(N324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(N325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(N326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(N327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(N328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(N329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(N330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(N331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(N332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(N333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(N334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(N335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(N336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(N337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(N338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(N339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(N340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(N341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(N342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(N343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(N344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(N345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(N346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(N347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(N348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(N349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(N350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(N351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(N352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(N353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(N354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(N355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(N356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(N357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(N358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(N359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(N360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(N361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(N362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(N363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(N364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(N365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(N366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(N367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(N368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(N369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(N370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(N371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(N372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(N373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(N374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(N375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(N376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(N377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(N378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(N379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(N380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(N381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(N382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(N383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(N384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(N385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(N386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(N387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(N388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(N389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(N390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(N391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(N392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(N393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(N394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(N395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(N396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(N397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(N398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(N399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(N400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(N401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(N402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(N403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(N404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(N405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(N406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(N407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(N408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(N409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(N410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(N411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(N412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(N413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(N414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(N415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(N416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(N417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(N418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(N419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(N420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(N421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(N422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(N423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(N424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(N425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(N426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(N427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(N428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(N429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(N430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(N431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(N432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(N433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(N434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(N435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(N436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(N437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(N438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(N439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(N440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(N441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(N442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(N443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(N444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(N445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(N446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(N447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(N448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(N449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(N450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(N451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(N452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(N453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(N454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(N455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(N456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(N457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(N458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(N459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(N460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(N461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(N462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(N463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(N464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(N465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(N466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(N467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(N468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(N469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(N470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(N471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(N472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(N473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(N474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(N475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(N476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(N477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(N478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(N479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(N480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(N481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(N482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(N483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(N484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(N485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(N486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(N487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(N488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(N489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(N490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(N491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(N492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(N493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(N494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(N495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(N496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(N497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(N498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(N499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(N500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(N501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(N502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(N503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(N504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(N505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(N506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(N507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(N508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(N509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(N510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(N511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(N512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(N513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(N514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(N515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(N516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(N517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(N518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(N519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(N520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(N521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(N522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(N523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(N524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(N525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(N526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(N527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(N528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(N529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(N530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(N531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(N532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(N533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(N534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(N535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(N536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(N537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(N538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(N539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(N540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(N541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(N542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(N543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(N544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(N545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(N546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(N547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(N548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(N549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(N550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(N551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(N552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(N553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(N554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(N555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(N556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(N557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(N558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(N559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(N560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(N561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(N562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(N563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(N564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(N565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(N566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(N567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(N568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(N569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(N570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(N571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(N572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(N573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(N574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(N575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(N576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(N577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(N578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(N579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(N580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(N581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(N582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(N583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(N584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(N585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(N586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(N587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(N588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(N589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(N590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(N591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(N592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(N593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(N594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(N595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(N596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(N597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(N598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(N599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(N600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(N601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(N602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(N603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(N604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(N605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(N606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(N607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(N608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(N609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(N610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(N611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(N612), .CLK(clk), .RST(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(N613), .CLK(clk), .RST(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(N614), .CLK(clk), .RST(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(N615), .CLK(clk), .RST(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(N616), .CLK(clk), .RST(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(N617), .CLK(clk), .RST(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(N618), .CLK(clk), .RST(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(N619), .CLK(clk), .RST(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(N620), .CLK(clk), .RST(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(N621), .CLK(clk), .RST(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(N622), .CLK(clk), .RST(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(N623), .CLK(clk), .RST(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(N624), .CLK(clk), .RST(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(N625), .CLK(clk), .RST(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(N626), .CLK(clk), .RST(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(N627), .CLK(clk), .RST(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(N628), .CLK(clk), .RST(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(N629), .CLK(clk), .RST(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(N630), .CLK(clk), .RST(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(N631), .CLK(clk), .RST(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(N632), .CLK(clk), .RST(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(N633), .CLK(clk), .RST(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(N634), .CLK(clk), .RST(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(N635), .CLK(clk), .RST(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(N636), .CLK(clk), .RST(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(N637), .CLK(clk), .RST(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(N638), .CLK(clk), .RST(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(N639), .CLK(clk), .RST(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(N640), .CLK(clk), .RST(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(N641), .CLK(clk), .RST(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(N642), .CLK(clk), .RST(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(N643), .CLK(clk), .RST(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(N644), .CLK(clk), .RST(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(N645), .CLK(clk), .RST(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(N646), .CLK(clk), .RST(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(N647), .CLK(clk), .RST(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(N648), .CLK(clk), .RST(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(N649), .CLK(clk), .RST(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(N650), .CLK(clk), .RST(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(N651), .CLK(clk), .RST(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(N652), .CLK(clk), .RST(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(N653), .CLK(clk), .RST(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(N654), .CLK(clk), .RST(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(N655), .CLK(clk), .RST(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(N656), .CLK(clk), .RST(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(N657), .CLK(clk), .RST(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(N658), .CLK(clk), .RST(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(N659), .CLK(clk), .RST(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(N660), .CLK(clk), .RST(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(N661), .CLK(clk), .RST(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(N662), .CLK(clk), .RST(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(N663), .CLK(clk), .RST(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(N664), .CLK(clk), .RST(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(N665), .CLK(clk), .RST(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(N666), .CLK(clk), .RST(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(N667), .CLK(clk), .RST(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(N668), .CLK(clk), .RST(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(N669), .CLK(clk), .RST(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(N670), .CLK(clk), .RST(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(N671), .CLK(clk), .RST(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(N672), .CLK(clk), .RST(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(N673), .CLK(clk), .RST(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(N674), .CLK(clk), .RST(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(N675), .CLK(clk), .RST(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(N676), .CLK(clk), .RST(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(N677), .CLK(clk), .RST(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(N678), .CLK(clk), .RST(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(N679), .CLK(clk), .RST(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(N680), .CLK(clk), .RST(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(N681), .CLK(clk), .RST(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(N682), .CLK(clk), .RST(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(N683), .CLK(clk), .RST(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(N684), .CLK(clk), .RST(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(N685), .CLK(clk), .RST(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(N686), .CLK(clk), .RST(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(N687), .CLK(clk), .RST(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(N688), .CLK(clk), .RST(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(N689), .CLK(clk), .RST(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(N690), .CLK(clk), .RST(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(N691), .CLK(clk), .RST(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(N692), .CLK(clk), .RST(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(N693), .CLK(clk), .RST(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(N694), .CLK(clk), .RST(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(N695), .CLK(clk), .RST(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(N696), .CLK(clk), .RST(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(N697), .CLK(clk), .RST(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(N698), .CLK(clk), .RST(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(N699), .CLK(clk), .RST(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(N700), .CLK(clk), .RST(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(N701), .CLK(clk), .RST(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(N702), .CLK(clk), .RST(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(N703), .CLK(clk), .RST(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(N704), .CLK(clk), .RST(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(N705), .CLK(clk), .RST(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(N706), .CLK(clk), .RST(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(N707), .CLK(clk), .RST(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(N708), .CLK(clk), .RST(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(N709), .CLK(clk), .RST(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(N710), .CLK(clk), .RST(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(N711), .CLK(clk), .RST(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(N712), .CLK(clk), .RST(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(N713), .CLK(clk), .RST(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(N714), .CLK(clk), .RST(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(N715), .CLK(clk), .RST(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(N716), .CLK(clk), .RST(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(N717), .CLK(clk), .RST(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(N718), .CLK(clk), .RST(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(N719), .CLK(clk), .RST(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(N720), .CLK(clk), .RST(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(N721), .CLK(clk), .RST(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(N722), .CLK(clk), .RST(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(N723), .CLK(clk), .RST(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(N724), .CLK(clk), .RST(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(N725), .CLK(clk), .RST(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(N726), .CLK(clk), .RST(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(N727), .CLK(clk), .RST(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(N728), .CLK(clk), .RST(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(N729), .CLK(clk), .RST(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(N730), .CLK(clk), .RST(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(N731), .CLK(clk), .RST(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(N732), .CLK(clk), .RST(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(N733), .CLK(clk), .RST(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(N734), .CLK(clk), .RST(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(N735), .CLK(clk), .RST(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(N736), .CLK(clk), .RST(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(N737), .CLK(clk), .RST(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(N738), .CLK(clk), .RST(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(N739), .CLK(clk), .RST(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(N740), .CLK(clk), .RST(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(N741), .CLK(clk), .RST(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(N742), .CLK(clk), .RST(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(N743), .CLK(clk), .RST(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(N744), .CLK(clk), .RST(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(N745), .CLK(clk), .RST(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(N746), .CLK(clk), .RST(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(N747), .CLK(clk), .RST(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(N748), .CLK(clk), .RST(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(N749), .CLK(clk), .RST(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(N750), .CLK(clk), .RST(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(N751), .CLK(clk), .RST(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(N752), .CLK(clk), .RST(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(N753), .CLK(clk), .RST(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(N754), .CLK(clk), .RST(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(N755), .CLK(clk), .RST(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(N756), .CLK(clk), .RST(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(N757), .CLK(clk), .RST(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(N758), .CLK(clk), .RST(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(N759), .CLK(clk), .RST(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(N760), .CLK(clk), .RST(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(N761), .CLK(clk), .RST(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(N762), .CLK(clk), .RST(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(N763), .CLK(clk), .RST(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(N764), .CLK(clk), .RST(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(N765), .CLK(clk), .RST(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(N766), .CLK(clk), .RST(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(N767), .CLK(clk), .RST(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(N768), .CLK(clk), .RST(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(N769), .CLK(clk), .RST(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(N770), .CLK(clk), .RST(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(N771), .CLK(clk), .RST(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(N772), .CLK(clk), .RST(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(N773), .CLK(clk), .RST(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(N774), .CLK(clk), .RST(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(N775), .CLK(clk), .RST(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(N776), .CLK(clk), .RST(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(N777), .CLK(clk), .RST(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(N778), .CLK(clk), .RST(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(N779), .CLK(clk), .RST(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(N780), .CLK(clk), .RST(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(N781), .CLK(clk), .RST(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(N782), .CLK(clk), .RST(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(N783), .CLK(clk), .RST(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(N784), .CLK(clk), .RST(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(N785), .CLK(clk), .RST(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(N786), .CLK(clk), .RST(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(N787), .CLK(clk), .RST(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(N788), .CLK(clk), .RST(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(N789), .CLK(clk), .RST(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(N790), .CLK(clk), .RST(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(N791), .CLK(clk), .RST(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(N792), .CLK(clk), .RST(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(N793), .CLK(clk), .RST(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(N794), .CLK(clk), .RST(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(N795), .CLK(clk), .RST(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(N796), .CLK(clk), .RST(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(N797), .CLK(clk), .RST(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(N798), .CLK(clk), .RST(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(N799), .CLK(clk), .RST(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(N800), .CLK(clk), .RST(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(N801), .CLK(clk), .RST(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(N802), .CLK(clk), .RST(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(N803), .CLK(clk), .RST(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(N804), .CLK(clk), .RST(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(N805), .CLK(clk), .RST(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(N806), .CLK(clk), .RST(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(N807), .CLK(clk), .RST(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(N808), .CLK(clk), .RST(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(N809), .CLK(clk), .RST(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(N810), .CLK(clk), .RST(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(N811), .CLK(clk), .RST(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(N812), .CLK(clk), .RST(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(N813), .CLK(clk), .RST(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(N814), .CLK(clk), .RST(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(N815), .CLK(clk), .RST(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(N816), .CLK(clk), .RST(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(N817), .CLK(clk), .RST(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(N818), .CLK(clk), .RST(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(N819), .CLK(clk), .RST(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(N820), .CLK(clk), .RST(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(N821), .CLK(clk), .RST(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(N822), .CLK(clk), .RST(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(N823), .CLK(clk), .RST(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(N824), .CLK(clk), .RST(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(N825), .CLK(clk), .RST(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(N826), .CLK(clk), .RST(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(N827), .CLK(clk), .RST(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(N828), .CLK(clk), .RST(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(N829), .CLK(clk), .RST(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(N830), .CLK(clk), .RST(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(N831), .CLK(clk), .RST(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(N832), .CLK(clk), .RST(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(N833), .CLK(clk), .RST(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(N834), .CLK(clk), .RST(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(N835), .CLK(clk), .RST(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(N836), .CLK(clk), .RST(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(N837), .CLK(clk), .RST(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(N838), .CLK(clk), .RST(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(N839), .CLK(clk), .RST(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(N840), .CLK(clk), .RST(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(N841), .CLK(clk), .RST(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(N842), .CLK(clk), .RST(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(N843), .CLK(clk), .RST(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(N844), .CLK(clk), .RST(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(N845), .CLK(clk), .RST(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(N846), .CLK(clk), .RST(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(N847), .CLK(clk), .RST(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(N848), .CLK(clk), .RST(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(N849), .CLK(clk), .RST(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(N850), .CLK(clk), .RST(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(N851), .CLK(clk), .RST(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(N852), .CLK(clk), .RST(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(N853), .CLK(clk), .RST(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(N854), .CLK(clk), .RST(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(N855), .CLK(clk), .RST(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(N856), .CLK(clk), .RST(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(N857), .CLK(clk), .RST(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(N858), .CLK(clk), .RST(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(N859), .CLK(clk), .RST(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(N860), .CLK(clk), .RST(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(N861), .CLK(clk), .RST(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(N862), .CLK(clk), .RST(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(N863), .CLK(clk), .RST(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(N864), .CLK(clk), .RST(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(N865), .CLK(clk), .RST(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(N866), .CLK(clk), .RST(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(N867), .CLK(clk), .RST(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(N868), .CLK(clk), .RST(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(N869), .CLK(clk), .RST(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(N870), .CLK(clk), .RST(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(N871), .CLK(clk), .RST(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(N872), .CLK(clk), .RST(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(N873), .CLK(clk), .RST(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(N874), .CLK(clk), .RST(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(N875), .CLK(clk), .RST(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(N876), .CLK(clk), .RST(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(N877), .CLK(clk), .RST(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(N878), .CLK(clk), .RST(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(N879), .CLK(clk), .RST(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(N880), .CLK(clk), .RST(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(N881), .CLK(clk), .RST(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(N882), .CLK(clk), .RST(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(N883), .CLK(clk), .RST(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(N884), .CLK(clk), .RST(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(N885), .CLK(clk), .RST(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(N886), .CLK(clk), .RST(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(N887), .CLK(clk), .RST(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(N888), .CLK(clk), .RST(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(N889), .CLK(clk), .RST(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(N890), .CLK(clk), .RST(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(N891), .CLK(clk), .RST(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(N892), .CLK(clk), .RST(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(N893), .CLK(clk), .RST(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(N894), .CLK(clk), .RST(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(N895), .CLK(clk), .RST(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(N896), .CLK(clk), .RST(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(N897), .CLK(clk), .RST(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(N898), .CLK(clk), .RST(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(N899), .CLK(clk), .RST(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(N900), .CLK(clk), .RST(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(N901), .CLK(clk), .RST(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(N902), .CLK(clk), .RST(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(N903), .CLK(clk), .RST(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(N904), .CLK(clk), .RST(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(N905), .CLK(clk), .RST(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(N906), .CLK(clk), .RST(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(N907), .CLK(clk), .RST(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(N908), .CLK(clk), .RST(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(N909), .CLK(clk), .RST(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(N910), .CLK(clk), .RST(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(N911), .CLK(clk), .RST(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(N912), .CLK(clk), .RST(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(N913), .CLK(clk), .RST(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(N914), .CLK(clk), .RST(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(N915), .CLK(clk), .RST(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(N916), .CLK(clk), .RST(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(N917), .CLK(clk), .RST(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(N918), .CLK(clk), .RST(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(N919), .CLK(clk), .RST(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(N920), .CLK(clk), .RST(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(N921), .CLK(clk), .RST(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(N922), .CLK(clk), .RST(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(N923), .CLK(clk), .RST(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(N924), .CLK(clk), .RST(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(N925), .CLK(clk), .RST(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(N926), .CLK(clk), .RST(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(N927), .CLK(clk), .RST(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(N928), .CLK(clk), .RST(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(N929), .CLK(clk), .RST(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(N930), .CLK(clk), .RST(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(N931), .CLK(clk), .RST(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(N932), .CLK(clk), .RST(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(N933), .CLK(clk), .RST(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(N934), .CLK(clk), .RST(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(N935), .CLK(clk), .RST(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(N936), .CLK(clk), .RST(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(N937), .CLK(clk), .RST(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(N938), .CLK(clk), .RST(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(N939), .CLK(clk), .RST(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(N940), .CLK(clk), .RST(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(N941), .CLK(clk), .RST(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(N942), .CLK(clk), .RST(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(N943), .CLK(clk), .RST(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(N944), .CLK(clk), .RST(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(N945), .CLK(clk), .RST(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(N946), .CLK(clk), .RST(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(N947), .CLK(clk), .RST(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(N948), .CLK(clk), .RST(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(N949), .CLK(clk), .RST(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(N950), .CLK(clk), .RST(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(N951), .CLK(clk), .RST(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(N952), .CLK(clk), .RST(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(N953), .CLK(clk), .RST(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(N954), .CLK(clk), .RST(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(N955), .CLK(clk), .RST(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(N956), .CLK(clk), .RST(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(N957), .CLK(clk), .RST(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(N958), .CLK(clk), .RST(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(N959), .CLK(clk), .RST(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(N960), .CLK(clk), .RST(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(N961), .CLK(clk), .RST(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(N962), .CLK(clk), .RST(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(N963), .CLK(clk), .RST(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(N964), .CLK(clk), .RST(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(N965), .CLK(clk), .RST(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(N966), .CLK(clk), .RST(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(N967), .CLK(clk), .RST(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(N968), .CLK(clk), .RST(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(N969), .CLK(clk), .RST(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(N970), .CLK(clk), .RST(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(N971), .CLK(clk), .RST(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(N972), .CLK(clk), .RST(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(N973), .CLK(clk), .RST(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(N974), .CLK(clk), .RST(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(N975), .CLK(clk), .RST(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(N976), .CLK(clk), .RST(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(N977), .CLK(clk), .RST(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(N978), .CLK(clk), .RST(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(N979), .CLK(clk), .RST(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(N980), .CLK(clk), .RST(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(N981), .CLK(clk), .RST(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(N982), .CLK(clk), .RST(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(N983), .CLK(clk), .RST(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(N984), .CLK(clk), .RST(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(N985), .CLK(clk), .RST(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(N986), .CLK(clk), .RST(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(N987), .CLK(clk), .RST(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(N988), .CLK(clk), .RST(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(N989), .CLK(clk), .RST(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(N990), .CLK(clk), .RST(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(N991), .CLK(clk), .RST(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(N992), .CLK(clk), .RST(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(N993), .CLK(clk), .RST(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(N994), .CLK(clk), .RST(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(N995), .CLK(clk), .RST(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(N996), .CLK(clk), .RST(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(N997), .CLK(clk), .RST(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(N998), .CLK(clk), .RST(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(N999), .CLK(clk), .RST(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(N1000), .CLK(clk), .RST(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(N1001), .CLK(clk), .RST(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(N1002), .CLK(clk), .RST(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(N1003), .CLK(clk), .RST(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(N1004), .CLK(clk), .RST(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(N1005), .CLK(clk), .RST(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(N1006), .CLK(clk), .RST(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(N1007), .CLK(clk), .RST(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(N1008), .CLK(clk), .RST(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(N1009), .CLK(clk), .RST(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(N1010), .CLK(clk), .RST(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(N1011), .CLK(clk), .RST(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(N1012), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(N1013), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(N1014), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(N1015), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(N1016), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(N1017), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(N1018), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(N1019), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(N1020), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(N1021), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(N1022), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(N1023), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(N1024), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(N1025), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(N1026), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(N1027), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(N1028), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(N1029), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(N1030), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(N1031), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(N1032), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(N1033), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(N1034), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(N1035), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(N1036), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(N1037), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(N1038), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(N1039), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(N1040), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(N1041), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(N1042), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(N1043), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(N1044), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(N1045), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(N1046), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(N1047), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(N1048), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(N1049), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(N1050), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(N1051), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(N1052), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(N1053), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(N1054), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(N1055), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(N1056), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(N1057), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(N1058), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(N1059), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(N1060), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(N1061), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(N1062), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(N1063), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(N1064), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(N1065), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(N1066), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(N1067), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(N1068), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(N1069), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(N1070), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(N1071), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(N1072), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(N1073), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(N1074), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(N1075), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(N1076), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(N1077), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(N1078), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(N1079), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(N1080), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(N1081), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(N1082), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(N1083), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(N1084), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(N1085), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(N1086), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(N1087), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(N1088), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(N1089), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(N1090), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(N1091), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(N1092), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(N1093), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(N1094), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(N1095), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(N1096), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(N1097), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(N1098), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(N1099), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(N1100), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(N1101), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(N1102), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(N1103), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(N1104), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(N1105), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(N1106), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(N1107), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(N1108), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(N1109), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(N1110), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(N1111), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(N1112), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(N1113), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(N1114), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(N1115), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(N1116), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(N1117), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(N1118), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(N1119), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(N1120), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(N1121), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(N1122), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(N1123), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(N1124), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(N1125), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(N1126), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(N1127), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(N1128), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(N1129), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(N1130), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(N1131), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(N1132), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(N1133), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(N1134), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(N1135), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(N1136), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(N1137), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(N1138), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(N1139), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(N1140), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(N1141), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(N1142), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(N1143), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(N1144), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(N1145), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(N1146), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(N1147), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(N1148), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(N1149), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(N1150), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(N1151), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(N1152), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(N1153), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(N1154), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(N1155), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(N1156), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(N1157), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(N1158), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(N1159), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(N1160), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(N1161), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(N1162), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(N1163), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(N1164), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(N1165), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(N1166), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(N1167), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(N1168), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(N1169), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(N1170), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(N1171), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(N1172), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(N1173), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(N1174), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(N1175), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(N1176), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(N1177), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(N1178), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(N1179), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(N1180), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(N1181), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(N1182), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(N1183), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(N1184), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(N1185), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(N1186), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(N1187), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(N1188), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(N1189), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(N1190), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(N1191), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(N1192), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(N1193), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(N1194), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(N1195), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(N1196), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(N1197), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(N1198), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(N1199), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(N1200), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(N1201), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(N1202), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(N1203), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(N1204), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(N1205), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(N1206), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(N1207), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(N1208), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(N1209), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(N1210), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(N1211), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(N1212), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(N1213), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(N1214), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(N1215), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(N1216), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(N1217), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(N1218), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(N1219), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(N1220), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(N1221), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(N1222), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(N1223), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(N1224), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(N1225), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(N1226), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(N1227), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(N1228), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(N1229), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(N1230), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(N1231), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(N1232), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(N1233), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(N1234), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(N1235), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(N1236), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(N1237), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(N1238), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(N1239), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(N1240), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(N1241), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(N1242), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(N1243), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(N1244), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(N1245), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(N1246), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(N1247), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(N1248), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(N1249), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(N1250), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(N1251), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(N1252), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(N1253), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(N1254), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(N1255), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(N1256), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(N1257), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(N1258), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(N1259), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(N1260), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(N1261), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(N1262), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(N1263), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(N1264), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(N1265), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(N1266), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(N1267), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(N1268), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(N1269), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(N1270), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(N1271), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(N1272), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(N1273), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(N1274), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(N1275), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(N1276), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(N1277), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(N1278), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(N1279), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(N1280), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(N1281), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(N1282), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(N1283), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(N1284), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(N1285), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(N1286), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(N1287), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(N1288), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(N1289), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(N1290), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(N1291), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(N1292), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(N1293), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(N1294), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(N1295), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(N1296), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(N1297), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(N1298), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(N1299), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(N1300), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(N1301), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(N1302), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(N1303), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(N1304), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(N1305), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(N1306), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(N1307), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(N1308), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(N1309), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(N1310), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(N1311), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(N1312), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(N1313), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(N1314), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(N1315), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(N1316), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(N1317), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(N1318), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(N1319), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(N1320), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(N1321), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(N1322), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(N1323), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(N1324), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(N1325), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(N1326), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(N1327), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(N1328), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(N1329), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(N1330), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(N1331), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(N1332), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(N1333), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(N1334), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(N1335), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(N1336), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(N1337), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(N1338), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(N1339), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(N1340), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(N1341), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(N1342), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(N1343), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(N1344), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(N1345), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(N1346), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(N1347), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(N1348), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(N1349), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(N1350), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(N1351), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(N1352), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(N1353), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(N1354), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(N1355), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(N1356), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(N1357), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(N1358), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(N1359), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(N1360), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(N1361), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(N1362), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(N1363), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(N1364), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(N1365), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(N1366), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(N1367), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(N1368), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(N1369), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(N1370), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(N1371), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(N1372), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(N1373), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(N1374), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(N1375), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(N1376), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(N1377), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(N1378), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(N1379), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(N1380), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(N1381), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(N1382), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(N1383), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(N1384), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(N1385), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(N1386), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(N1387), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(N1388), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(N1389), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(N1390), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(N1391), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(N1392), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(N1393), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(N1394), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(N1395), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(N1396), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(N1397), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(N1398), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(N1399), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(N1400), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(N1401), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(N1402), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(N1403), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(N1404), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(N1405), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(N1406), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(N1407), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(N1408), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(N1409), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(N1410), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(N1411), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(N1412), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(N1413), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(N1414), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(N1415), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(N1416), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(N1417), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(N1418), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(N1419), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(N1420), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(N1421), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(N1422), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(N1423), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(N1424), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(N1425), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(N1426), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(N1427), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(N1428), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(N1429), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(N1430), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(N1431), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(N1432), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(N1433), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(N1434), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(N1435), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(N1436), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(N1437), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(N1438), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(N1439), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(N1440), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(N1441), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(N1442), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(N1443), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(N1444), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(N1445), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(N1446), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(N1447), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(N1448), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(N1449), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(N1450), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(N1451), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(N1452), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(N1453), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(N1454), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(N1455), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(N1456), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(N1457), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(N1458), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(N1459), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(N1460), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(N1461), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(N1462), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(N1463), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(N1464), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(N1465), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(N1466), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(N1467), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(N1468), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(N1469), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(N1470), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(N1471), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(N1472), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(N1473), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(N1474), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(N1475), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(N1476), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(N1477), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(N1478), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(N1479), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(N1480), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(N1481), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(N1482), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(N1483), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(N1484), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(N1485), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(N1486), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(N1487), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(N1488), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(N1489), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(N1490), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(N1491), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(N1492), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(N1493), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(N1494), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(N1495), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(N1496), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(N1497), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(N1498), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(N1499), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(N1500), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(N1501), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(N1502), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(N1503), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(N1504), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(N1505), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(N1506), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(N1507), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(N1508), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(N1509), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(N1510), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(N1511), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(N1512), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(N1513), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(N1514), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(N1515), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(N1516), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(N1517), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(N1518), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(N1519), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(N1520), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(N1521), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(N1522), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(N1523), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(N1524), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(N1525), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(N1526), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(N1527), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(N1528), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(N1529), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(N1530), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(N1531), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(N1532), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(N1533), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(N1534), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(N1535), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(N1536), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(N1537), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(N1538), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(N1539), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(N1540), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(N1541), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(N1542), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(N1543), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(N1544), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(N1545), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(N1546), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(N1547), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(N1548), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(N1549), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(N1550), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(N1551), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(N1552), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(N1553), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(N1554), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(N1555), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(N1556), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(N1557), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(N1558), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(N1559), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(N1560), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(N1561), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(N1562), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(N1563), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(N1564), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(N1565), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(N1566), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(N1567), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(N1568), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(N1569), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(N1570), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(N1571), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(N1572), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(N1573), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(N1574), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(N1575), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(N1576), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(N1577), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(N1578), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(N1579), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(N1580), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(N1581), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(N1582), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(N1583), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(N1584), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(N1585), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(N1586), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(N1587), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(N1588), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(N1589), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(N1590), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(N1591), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(N1592), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(N1593), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(N1594), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(N1595), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(N1596), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(N1597), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(N1598), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(N1599), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(N1600), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(N1601), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(N1602), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(N1603), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(N1604), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(N1605), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(N1606), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(N1607), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(N1608), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(N1609), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(N1610), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(N1611), .CLK(clk), .RST(1'b0), .Q(
        round_reg[1599]) );
  NANDN U5999 ( .A(rc_i[0]), .B(n2856), .Z(\RCONST[2].rconst_/N18 ) );
  NANDN U6000 ( .A(\rc[3][15] ), .B(n2856), .Z(\rc[3][63] ) );
  IV U6001 ( .A(init), .Z(n2770) );
  IV U6002 ( .A(init), .Z(n2771) );
  IV U6003 ( .A(init), .Z(n2772) );
  IV U6004 ( .A(init), .Z(n2773) );
  IV U6005 ( .A(init), .Z(n2774) );
  IV U6006 ( .A(init), .Z(n2775) );
  IV U6007 ( .A(init), .Z(n2776) );
  IV U6008 ( .A(init), .Z(n2777) );
  IV U6009 ( .A(init), .Z(n2778) );
  IV U6010 ( .A(init), .Z(n2779) );
  IV U6011 ( .A(init), .Z(n2780) );
  IV U6012 ( .A(init), .Z(n2781) );
  IV U6013 ( .A(init), .Z(n2782) );
  IV U6014 ( .A(init), .Z(n2783) );
  IV U6015 ( .A(init), .Z(n2784) );
  IV U6016 ( .A(init), .Z(n2785) );
  IV U6017 ( .A(init), .Z(n2786) );
  IV U6018 ( .A(init), .Z(n2787) );
  IV U6019 ( .A(init), .Z(n2788) );
  IV U6020 ( .A(init), .Z(n2789) );
  IV U6021 ( .A(init), .Z(n2790) );
  IV U6022 ( .A(init), .Z(n2791) );
  IV U6023 ( .A(init), .Z(n2792) );
  IV U6024 ( .A(init), .Z(n2793) );
  IV U6025 ( .A(init), .Z(n2794) );
  IV U6026 ( .A(init), .Z(n2795) );
  IV U6027 ( .A(init), .Z(n2796) );
  IV U6028 ( .A(init), .Z(n2797) );
  IV U6029 ( .A(init), .Z(n2798) );
  IV U6030 ( .A(init), .Z(n2799) );
  IV U6031 ( .A(init), .Z(n2800) );
  IV U6032 ( .A(init), .Z(n2801) );
  IV U6033 ( .A(init), .Z(n2802) );
  IV U6034 ( .A(init), .Z(n2803) );
  IV U6035 ( .A(init), .Z(n2804) );
  IV U6036 ( .A(init), .Z(n2805) );
  IV U6037 ( .A(init), .Z(n2806) );
  IV U6038 ( .A(init), .Z(n2807) );
  IV U6039 ( .A(init), .Z(n2808) );
  IV U6040 ( .A(init), .Z(n2809) );
  IV U6041 ( .A(init), .Z(n2810) );
  IV U6042 ( .A(init), .Z(n2811) );
  IV U6043 ( .A(init), .Z(n2812) );
  IV U6044 ( .A(init), .Z(n2813) );
  IV U6045 ( .A(init), .Z(n2814) );
  IV U6046 ( .A(init), .Z(n2815) );
  IV U6047 ( .A(init), .Z(n2816) );
  IV U6048 ( .A(init), .Z(n2817) );
  IV U6049 ( .A(init), .Z(n2818) );
  IV U6050 ( .A(init), .Z(n2819) );
  IV U6051 ( .A(init), .Z(n2820) );
  IV U6052 ( .A(init), .Z(n2821) );
  IV U6053 ( .A(init), .Z(n2822) );
  IV U6054 ( .A(init), .Z(n2823) );
  IV U6055 ( .A(init), .Z(n2824) );
  IV U6056 ( .A(init), .Z(n2825) );
  IV U6057 ( .A(init), .Z(n2826) );
  IV U6058 ( .A(init), .Z(n2827) );
  IV U6059 ( .A(init), .Z(n2828) );
  IV U6060 ( .A(init), .Z(n2829) );
  IV U6061 ( .A(init), .Z(n2830) );
  IV U6062 ( .A(init), .Z(n2831) );
  IV U6063 ( .A(init), .Z(n2832) );
  IV U6064 ( .A(init), .Z(n2833) );
  IV U6065 ( .A(init), .Z(n2834) );
  IV U6066 ( .A(init), .Z(n2835) );
  IV U6067 ( .A(init), .Z(n2836) );
  IV U6068 ( .A(init), .Z(n2837) );
  IV U6069 ( .A(init), .Z(n2838) );
  IV U6070 ( .A(init), .Z(n2839) );
  IV U6071 ( .A(init), .Z(n2840) );
  IV U6072 ( .A(init), .Z(n2841) );
  IV U6073 ( .A(init), .Z(n2842) );
  IV U6074 ( .A(init), .Z(n2843) );
  IV U6075 ( .A(init), .Z(n2844) );
  IV U6076 ( .A(init), .Z(n2845) );
  IV U6077 ( .A(init), .Z(n2846) );
  IV U6078 ( .A(init), .Z(n2847) );
  IV U6079 ( .A(init), .Z(n2848) );
  IV U6080 ( .A(init), .Z(n2849) );
  IV U6081 ( .A(init), .Z(n2850) );
  IV U6082 ( .A(init), .Z(n2851) );
  IV U6083 ( .A(init), .Z(n2852) );
  IV U6085 ( .A(rst), .Z(n1614) );
  AND U6086 ( .A(rc_i[3]), .B(n1614), .Z(N10) );
  AND U6087 ( .A(out[88]), .B(n1614), .Z(N100) );
  AND U6088 ( .A(out[988]), .B(n1614), .Z(N1000) );
  AND U6089 ( .A(out[989]), .B(n1614), .Z(N1001) );
  AND U6090 ( .A(out[990]), .B(n1614), .Z(N1002) );
  AND U6091 ( .A(out[991]), .B(n1614), .Z(N1003) );
  AND U6092 ( .A(out[992]), .B(n1614), .Z(N1004) );
  AND U6093 ( .A(out[993]), .B(n1614), .Z(N1005) );
  AND U6094 ( .A(out[994]), .B(n1614), .Z(N1006) );
  AND U6095 ( .A(out[995]), .B(n1614), .Z(N1007) );
  AND U6096 ( .A(out[996]), .B(n1614), .Z(N1008) );
  AND U6097 ( .A(out[997]), .B(n1614), .Z(N1009) );
  AND U6098 ( .A(out[89]), .B(n1614), .Z(N101) );
  AND U6099 ( .A(out[998]), .B(n1614), .Z(N1010) );
  AND U6100 ( .A(out[999]), .B(n1614), .Z(N1011) );
  AND U6101 ( .A(out[1000]), .B(n1614), .Z(N1012) );
  AND U6102 ( .A(out[1001]), .B(n1614), .Z(N1013) );
  AND U6103 ( .A(out[1002]), .B(n1614), .Z(N1014) );
  AND U6104 ( .A(out[1003]), .B(n1614), .Z(N1015) );
  AND U6105 ( .A(out[1004]), .B(n1614), .Z(N1016) );
  AND U6106 ( .A(out[1005]), .B(n1614), .Z(N1017) );
  AND U6107 ( .A(out[1006]), .B(n1614), .Z(N1018) );
  AND U6108 ( .A(out[1007]), .B(n1614), .Z(N1019) );
  AND U6109 ( .A(out[90]), .B(n1614), .Z(N102) );
  AND U6110 ( .A(out[1008]), .B(n1614), .Z(N1020) );
  AND U6111 ( .A(out[1009]), .B(n1614), .Z(N1021) );
  AND U6112 ( .A(out[1010]), .B(n1614), .Z(N1022) );
  AND U6113 ( .A(out[1011]), .B(n1614), .Z(N1023) );
  AND U6114 ( .A(out[1012]), .B(n1614), .Z(N1024) );
  AND U6115 ( .A(out[1013]), .B(n1614), .Z(N1025) );
  AND U6116 ( .A(out[1014]), .B(n1614), .Z(N1026) );
  AND U6117 ( .A(out[1015]), .B(n1614), .Z(N1027) );
  AND U6118 ( .A(out[1016]), .B(n1614), .Z(N1028) );
  AND U6119 ( .A(out[1017]), .B(n1614), .Z(N1029) );
  AND U6120 ( .A(out[91]), .B(n1614), .Z(N103) );
  AND U6121 ( .A(out[1018]), .B(n1614), .Z(N1030) );
  AND U6122 ( .A(out[1019]), .B(n1614), .Z(N1031) );
  AND U6123 ( .A(out[1020]), .B(n1614), .Z(N1032) );
  AND U6124 ( .A(out[1021]), .B(n1614), .Z(N1033) );
  AND U6125 ( .A(out[1022]), .B(n1614), .Z(N1034) );
  AND U6126 ( .A(out[1023]), .B(n1614), .Z(N1035) );
  AND U6127 ( .A(out[1024]), .B(n1614), .Z(N1036) );
  AND U6128 ( .A(out[1025]), .B(n1614), .Z(N1037) );
  AND U6129 ( .A(out[1026]), .B(n1614), .Z(N1038) );
  AND U6130 ( .A(out[1027]), .B(n1614), .Z(N1039) );
  AND U6131 ( .A(out[92]), .B(n1614), .Z(N104) );
  AND U6132 ( .A(out[1028]), .B(n1614), .Z(N1040) );
  AND U6133 ( .A(out[1029]), .B(n1614), .Z(N1041) );
  AND U6134 ( .A(out[1030]), .B(n1614), .Z(N1042) );
  AND U6135 ( .A(out[1031]), .B(n1614), .Z(N1043) );
  AND U6136 ( .A(out[1032]), .B(n1614), .Z(N1044) );
  AND U6137 ( .A(out[1033]), .B(n1614), .Z(N1045) );
  AND U6138 ( .A(out[1034]), .B(n1614), .Z(N1046) );
  AND U6139 ( .A(out[1035]), .B(n1614), .Z(N1047) );
  AND U6140 ( .A(out[1036]), .B(n1614), .Z(N1048) );
  AND U6141 ( .A(out[1037]), .B(n1614), .Z(N1049) );
  AND U6142 ( .A(out[93]), .B(n1614), .Z(N105) );
  AND U6143 ( .A(out[1038]), .B(n1614), .Z(N1050) );
  AND U6144 ( .A(out[1039]), .B(n1614), .Z(N1051) );
  AND U6145 ( .A(out[1040]), .B(n1614), .Z(N1052) );
  AND U6146 ( .A(out[1041]), .B(n1614), .Z(N1053) );
  AND U6147 ( .A(out[1042]), .B(n1614), .Z(N1054) );
  AND U6148 ( .A(out[1043]), .B(n1614), .Z(N1055) );
  AND U6149 ( .A(out[1044]), .B(n1614), .Z(N1056) );
  AND U6150 ( .A(out[1045]), .B(n1614), .Z(N1057) );
  AND U6151 ( .A(out[1046]), .B(n1614), .Z(N1058) );
  AND U6152 ( .A(out[1047]), .B(n1614), .Z(N1059) );
  AND U6153 ( .A(out[94]), .B(n1614), .Z(N106) );
  AND U6154 ( .A(out[1048]), .B(n1614), .Z(N1060) );
  AND U6155 ( .A(out[1049]), .B(n1614), .Z(N1061) );
  AND U6156 ( .A(out[1050]), .B(n1614), .Z(N1062) );
  AND U6157 ( .A(out[1051]), .B(n1614), .Z(N1063) );
  AND U6158 ( .A(out[1052]), .B(n1614), .Z(N1064) );
  AND U6159 ( .A(out[1053]), .B(n1614), .Z(N1065) );
  AND U6160 ( .A(out[1054]), .B(n1614), .Z(N1066) );
  AND U6161 ( .A(out[1055]), .B(n1614), .Z(N1067) );
  AND U6162 ( .A(out[1056]), .B(n1614), .Z(N1068) );
  AND U6163 ( .A(out[1057]), .B(n1614), .Z(N1069) );
  AND U6164 ( .A(out[95]), .B(n1614), .Z(N107) );
  AND U6165 ( .A(out[1058]), .B(n1614), .Z(N1070) );
  AND U6166 ( .A(out[1059]), .B(n1614), .Z(N1071) );
  AND U6167 ( .A(out[1060]), .B(n1614), .Z(N1072) );
  AND U6168 ( .A(out[1061]), .B(n1614), .Z(N1073) );
  AND U6169 ( .A(out[1062]), .B(n1614), .Z(N1074) );
  AND U6170 ( .A(out[1063]), .B(n1614), .Z(N1075) );
  AND U6171 ( .A(out[1064]), .B(n1614), .Z(N1076) );
  AND U6172 ( .A(out[1065]), .B(n1614), .Z(N1077) );
  AND U6173 ( .A(out[1066]), .B(n1614), .Z(N1078) );
  AND U6174 ( .A(out[1067]), .B(n1614), .Z(N1079) );
  AND U6175 ( .A(out[96]), .B(n1614), .Z(N108) );
  AND U6176 ( .A(out[1068]), .B(n1614), .Z(N1080) );
  AND U6177 ( .A(out[1069]), .B(n1614), .Z(N1081) );
  AND U6178 ( .A(out[1070]), .B(n1614), .Z(N1082) );
  AND U6179 ( .A(out[1071]), .B(n1614), .Z(N1083) );
  AND U6180 ( .A(out[1072]), .B(n1614), .Z(N1084) );
  AND U6181 ( .A(out[1073]), .B(n1614), .Z(N1085) );
  AND U6182 ( .A(out[1074]), .B(n1614), .Z(N1086) );
  AND U6183 ( .A(out[1075]), .B(n1614), .Z(N1087) );
  AND U6184 ( .A(out[1076]), .B(n1614), .Z(N1088) );
  AND U6185 ( .A(out[1077]), .B(n1614), .Z(N1089) );
  AND U6186 ( .A(out[97]), .B(n1614), .Z(N109) );
  AND U6187 ( .A(out[1078]), .B(n1614), .Z(N1090) );
  AND U6188 ( .A(out[1079]), .B(n1614), .Z(N1091) );
  AND U6189 ( .A(out[1080]), .B(n1614), .Z(N1092) );
  AND U6190 ( .A(out[1081]), .B(n1614), .Z(N1093) );
  AND U6191 ( .A(out[1082]), .B(n1614), .Z(N1094) );
  AND U6192 ( .A(out[1083]), .B(n1614), .Z(N1095) );
  AND U6193 ( .A(out[1084]), .B(n1614), .Z(N1096) );
  AND U6194 ( .A(out[1085]), .B(n1614), .Z(N1097) );
  AND U6195 ( .A(out[1086]), .B(n1614), .Z(N1098) );
  AND U6196 ( .A(out[1087]), .B(n1614), .Z(N1099) );
  AND U6197 ( .A(rc_i[4]), .B(n1614), .Z(N11) );
  AND U6198 ( .A(out[98]), .B(n1614), .Z(N110) );
  AND U6199 ( .A(out[1088]), .B(n1614), .Z(N1100) );
  AND U6200 ( .A(out[1089]), .B(n1614), .Z(N1101) );
  AND U6201 ( .A(out[1090]), .B(n1614), .Z(N1102) );
  AND U6202 ( .A(out[1091]), .B(n1614), .Z(N1103) );
  AND U6203 ( .A(out[1092]), .B(n1614), .Z(N1104) );
  AND U6204 ( .A(out[1093]), .B(n1614), .Z(N1105) );
  AND U6205 ( .A(out[1094]), .B(n1614), .Z(N1106) );
  AND U6206 ( .A(out[1095]), .B(n1614), .Z(N1107) );
  AND U6207 ( .A(out[1096]), .B(n1614), .Z(N1108) );
  AND U6208 ( .A(out[1097]), .B(n1614), .Z(N1109) );
  AND U6209 ( .A(out[99]), .B(n1614), .Z(N111) );
  AND U6210 ( .A(out[1098]), .B(n1614), .Z(N1110) );
  AND U6211 ( .A(out[1099]), .B(n1614), .Z(N1111) );
  AND U6212 ( .A(out[1100]), .B(n1614), .Z(N1112) );
  AND U6213 ( .A(out[1101]), .B(n1614), .Z(N1113) );
  AND U6214 ( .A(out[1102]), .B(n1614), .Z(N1114) );
  AND U6215 ( .A(out[1103]), .B(n1614), .Z(N1115) );
  AND U6216 ( .A(out[1104]), .B(n1614), .Z(N1116) );
  AND U6217 ( .A(out[1105]), .B(n1614), .Z(N1117) );
  AND U6218 ( .A(out[1106]), .B(n1614), .Z(N1118) );
  AND U6219 ( .A(out[1107]), .B(n1614), .Z(N1119) );
  AND U6220 ( .A(out[100]), .B(n1614), .Z(N112) );
  AND U6221 ( .A(out[1108]), .B(n1614), .Z(N1120) );
  AND U6222 ( .A(out[1109]), .B(n1614), .Z(N1121) );
  AND U6223 ( .A(out[1110]), .B(n1614), .Z(N1122) );
  AND U6224 ( .A(out[1111]), .B(n1614), .Z(N1123) );
  AND U6225 ( .A(out[1112]), .B(n1614), .Z(N1124) );
  AND U6226 ( .A(out[1113]), .B(n1614), .Z(N1125) );
  AND U6227 ( .A(out[1114]), .B(n1614), .Z(N1126) );
  AND U6228 ( .A(out[1115]), .B(n1614), .Z(N1127) );
  AND U6229 ( .A(out[1116]), .B(n1614), .Z(N1128) );
  AND U6230 ( .A(out[1117]), .B(n1614), .Z(N1129) );
  AND U6231 ( .A(out[101]), .B(n1614), .Z(N113) );
  AND U6232 ( .A(out[1118]), .B(n1614), .Z(N1130) );
  AND U6233 ( .A(out[1119]), .B(n1614), .Z(N1131) );
  AND U6234 ( .A(out[1120]), .B(n1614), .Z(N1132) );
  AND U6235 ( .A(out[1121]), .B(n1614), .Z(N1133) );
  AND U6236 ( .A(out[1122]), .B(n1614), .Z(N1134) );
  AND U6237 ( .A(out[1123]), .B(n1614), .Z(N1135) );
  AND U6238 ( .A(out[1124]), .B(n1614), .Z(N1136) );
  AND U6239 ( .A(out[1125]), .B(n1614), .Z(N1137) );
  AND U6240 ( .A(out[1126]), .B(n1614), .Z(N1138) );
  AND U6241 ( .A(out[1127]), .B(n1614), .Z(N1139) );
  AND U6242 ( .A(out[102]), .B(n1614), .Z(N114) );
  AND U6243 ( .A(out[1128]), .B(n1614), .Z(N1140) );
  AND U6244 ( .A(out[1129]), .B(n1614), .Z(N1141) );
  AND U6245 ( .A(out[1130]), .B(n1614), .Z(N1142) );
  AND U6246 ( .A(out[1131]), .B(n1614), .Z(N1143) );
  AND U6247 ( .A(out[1132]), .B(n1614), .Z(N1144) );
  AND U6248 ( .A(out[1133]), .B(n1614), .Z(N1145) );
  AND U6249 ( .A(out[1134]), .B(n1614), .Z(N1146) );
  AND U6250 ( .A(out[1135]), .B(n1614), .Z(N1147) );
  AND U6251 ( .A(out[1136]), .B(n1614), .Z(N1148) );
  AND U6252 ( .A(out[1137]), .B(n1614), .Z(N1149) );
  AND U6253 ( .A(out[103]), .B(n1614), .Z(N115) );
  AND U6254 ( .A(out[1138]), .B(n1614), .Z(N1150) );
  AND U6255 ( .A(out[1139]), .B(n1614), .Z(N1151) );
  AND U6256 ( .A(out[1140]), .B(n1614), .Z(N1152) );
  AND U6257 ( .A(out[1141]), .B(n1614), .Z(N1153) );
  AND U6258 ( .A(out[1142]), .B(n1614), .Z(N1154) );
  AND U6259 ( .A(out[1143]), .B(n1614), .Z(N1155) );
  AND U6260 ( .A(out[1144]), .B(n1614), .Z(N1156) );
  AND U6261 ( .A(out[1145]), .B(n1614), .Z(N1157) );
  AND U6262 ( .A(out[1146]), .B(n1614), .Z(N1158) );
  AND U6263 ( .A(out[1147]), .B(n1614), .Z(N1159) );
  AND U6264 ( .A(out[104]), .B(n1614), .Z(N116) );
  AND U6265 ( .A(out[1148]), .B(n1614), .Z(N1160) );
  AND U6266 ( .A(out[1149]), .B(n1614), .Z(N1161) );
  AND U6267 ( .A(out[1150]), .B(n1614), .Z(N1162) );
  AND U6268 ( .A(out[1151]), .B(n1614), .Z(N1163) );
  AND U6269 ( .A(out[1152]), .B(n1614), .Z(N1164) );
  AND U6270 ( .A(out[1153]), .B(n1614), .Z(N1165) );
  AND U6271 ( .A(out[1154]), .B(n1614), .Z(N1166) );
  AND U6272 ( .A(out[1155]), .B(n1614), .Z(N1167) );
  AND U6273 ( .A(out[1156]), .B(n1614), .Z(N1168) );
  AND U6274 ( .A(out[1157]), .B(n1614), .Z(N1169) );
  AND U6275 ( .A(out[105]), .B(n1614), .Z(N117) );
  AND U6276 ( .A(out[1158]), .B(n1614), .Z(N1170) );
  AND U6277 ( .A(out[1159]), .B(n1614), .Z(N1171) );
  AND U6278 ( .A(out[1160]), .B(n1614), .Z(N1172) );
  AND U6279 ( .A(out[1161]), .B(n1614), .Z(N1173) );
  AND U6280 ( .A(out[1162]), .B(n1614), .Z(N1174) );
  AND U6281 ( .A(out[1163]), .B(n1614), .Z(N1175) );
  AND U6282 ( .A(out[1164]), .B(n1614), .Z(N1176) );
  AND U6283 ( .A(out[1165]), .B(n1614), .Z(N1177) );
  AND U6284 ( .A(out[1166]), .B(n1614), .Z(N1178) );
  AND U6285 ( .A(out[1167]), .B(n1614), .Z(N1179) );
  AND U6286 ( .A(out[106]), .B(n1614), .Z(N118) );
  AND U6287 ( .A(out[1168]), .B(n1614), .Z(N1180) );
  AND U6288 ( .A(out[1169]), .B(n1614), .Z(N1181) );
  AND U6289 ( .A(out[1170]), .B(n1614), .Z(N1182) );
  AND U6290 ( .A(out[1171]), .B(n1614), .Z(N1183) );
  AND U6291 ( .A(out[1172]), .B(n1614), .Z(N1184) );
  AND U6292 ( .A(out[1173]), .B(n1614), .Z(N1185) );
  AND U6293 ( .A(out[1174]), .B(n1614), .Z(N1186) );
  AND U6294 ( .A(out[1175]), .B(n1614), .Z(N1187) );
  AND U6295 ( .A(out[1176]), .B(n1614), .Z(N1188) );
  AND U6296 ( .A(out[1177]), .B(n1614), .Z(N1189) );
  AND U6297 ( .A(out[107]), .B(n1614), .Z(N119) );
  AND U6298 ( .A(out[1178]), .B(n1614), .Z(N1190) );
  AND U6299 ( .A(out[1179]), .B(n1614), .Z(N1191) );
  AND U6300 ( .A(out[1180]), .B(n1614), .Z(N1192) );
  AND U6301 ( .A(out[1181]), .B(n1614), .Z(N1193) );
  AND U6302 ( .A(out[1182]), .B(n1614), .Z(N1194) );
  AND U6303 ( .A(out[1183]), .B(n1614), .Z(N1195) );
  AND U6304 ( .A(out[1184]), .B(n1614), .Z(N1196) );
  AND U6305 ( .A(out[1185]), .B(n1614), .Z(N1197) );
  AND U6306 ( .A(out[1186]), .B(n1614), .Z(N1198) );
  AND U6307 ( .A(out[1187]), .B(n1614), .Z(N1199) );
  AND U6308 ( .A(out[0]), .B(n1614), .Z(N12) );
  AND U6309 ( .A(out[108]), .B(n1614), .Z(N120) );
  AND U6310 ( .A(out[1188]), .B(n1614), .Z(N1200) );
  AND U6311 ( .A(out[1189]), .B(n1614), .Z(N1201) );
  AND U6312 ( .A(out[1190]), .B(n1614), .Z(N1202) );
  AND U6313 ( .A(out[1191]), .B(n1614), .Z(N1203) );
  AND U6314 ( .A(out[1192]), .B(n1614), .Z(N1204) );
  AND U6315 ( .A(out[1193]), .B(n1614), .Z(N1205) );
  AND U6316 ( .A(out[1194]), .B(n1614), .Z(N1206) );
  AND U6317 ( .A(out[1195]), .B(n1614), .Z(N1207) );
  AND U6318 ( .A(out[1196]), .B(n1614), .Z(N1208) );
  AND U6319 ( .A(out[1197]), .B(n1614), .Z(N1209) );
  AND U6320 ( .A(out[109]), .B(n1614), .Z(N121) );
  AND U6321 ( .A(out[1198]), .B(n1614), .Z(N1210) );
  AND U6322 ( .A(out[1199]), .B(n1614), .Z(N1211) );
  AND U6323 ( .A(out[1200]), .B(n1614), .Z(N1212) );
  AND U6324 ( .A(out[1201]), .B(n1614), .Z(N1213) );
  AND U6325 ( .A(out[1202]), .B(n1614), .Z(N1214) );
  AND U6326 ( .A(out[1203]), .B(n1614), .Z(N1215) );
  AND U6327 ( .A(out[1204]), .B(n1614), .Z(N1216) );
  AND U6328 ( .A(out[1205]), .B(n1614), .Z(N1217) );
  AND U6329 ( .A(out[1206]), .B(n1614), .Z(N1218) );
  AND U6330 ( .A(out[1207]), .B(n1614), .Z(N1219) );
  AND U6331 ( .A(out[110]), .B(n1614), .Z(N122) );
  AND U6332 ( .A(out[1208]), .B(n1614), .Z(N1220) );
  AND U6333 ( .A(out[1209]), .B(n1614), .Z(N1221) );
  AND U6334 ( .A(out[1210]), .B(n1614), .Z(N1222) );
  AND U6335 ( .A(out[1211]), .B(n1614), .Z(N1223) );
  AND U6336 ( .A(out[1212]), .B(n1614), .Z(N1224) );
  AND U6337 ( .A(out[1213]), .B(n1614), .Z(N1225) );
  AND U6338 ( .A(out[1214]), .B(n1614), .Z(N1226) );
  AND U6339 ( .A(out[1215]), .B(n1614), .Z(N1227) );
  AND U6340 ( .A(out[1216]), .B(n1614), .Z(N1228) );
  AND U6341 ( .A(out[1217]), .B(n1614), .Z(N1229) );
  AND U6342 ( .A(out[111]), .B(n1614), .Z(N123) );
  AND U6343 ( .A(out[1218]), .B(n1614), .Z(N1230) );
  AND U6344 ( .A(out[1219]), .B(n1614), .Z(N1231) );
  AND U6345 ( .A(out[1220]), .B(n1614), .Z(N1232) );
  AND U6346 ( .A(out[1221]), .B(n1614), .Z(N1233) );
  AND U6347 ( .A(out[1222]), .B(n1614), .Z(N1234) );
  AND U6348 ( .A(out[1223]), .B(n1614), .Z(N1235) );
  AND U6349 ( .A(out[1224]), .B(n1614), .Z(N1236) );
  AND U6350 ( .A(out[1225]), .B(n1614), .Z(N1237) );
  AND U6351 ( .A(out[1226]), .B(n1614), .Z(N1238) );
  AND U6352 ( .A(out[1227]), .B(n1614), .Z(N1239) );
  AND U6353 ( .A(out[112]), .B(n1614), .Z(N124) );
  AND U6354 ( .A(out[1228]), .B(n1614), .Z(N1240) );
  AND U6355 ( .A(out[1229]), .B(n1614), .Z(N1241) );
  AND U6356 ( .A(out[1230]), .B(n1614), .Z(N1242) );
  AND U6357 ( .A(out[1231]), .B(n1614), .Z(N1243) );
  AND U6358 ( .A(out[1232]), .B(n1614), .Z(N1244) );
  AND U6359 ( .A(out[1233]), .B(n1614), .Z(N1245) );
  AND U6360 ( .A(out[1234]), .B(n1614), .Z(N1246) );
  AND U6361 ( .A(out[1235]), .B(n1614), .Z(N1247) );
  AND U6362 ( .A(out[1236]), .B(n1614), .Z(N1248) );
  AND U6363 ( .A(out[1237]), .B(n1614), .Z(N1249) );
  AND U6364 ( .A(out[113]), .B(n1614), .Z(N125) );
  AND U6365 ( .A(out[1238]), .B(n1614), .Z(N1250) );
  AND U6366 ( .A(out[1239]), .B(n1614), .Z(N1251) );
  AND U6367 ( .A(out[1240]), .B(n1614), .Z(N1252) );
  AND U6368 ( .A(out[1241]), .B(n1614), .Z(N1253) );
  AND U6369 ( .A(out[1242]), .B(n1614), .Z(N1254) );
  AND U6370 ( .A(out[1243]), .B(n1614), .Z(N1255) );
  AND U6371 ( .A(out[1244]), .B(n1614), .Z(N1256) );
  AND U6372 ( .A(out[1245]), .B(n1614), .Z(N1257) );
  AND U6373 ( .A(out[1246]), .B(n1614), .Z(N1258) );
  AND U6374 ( .A(out[1247]), .B(n1614), .Z(N1259) );
  AND U6375 ( .A(out[114]), .B(n1614), .Z(N126) );
  AND U6376 ( .A(out[1248]), .B(n1614), .Z(N1260) );
  AND U6377 ( .A(out[1249]), .B(n1614), .Z(N1261) );
  AND U6378 ( .A(out[1250]), .B(n1614), .Z(N1262) );
  AND U6379 ( .A(out[1251]), .B(n1614), .Z(N1263) );
  AND U6380 ( .A(out[1252]), .B(n1614), .Z(N1264) );
  AND U6381 ( .A(out[1253]), .B(n1614), .Z(N1265) );
  AND U6382 ( .A(out[1254]), .B(n1614), .Z(N1266) );
  AND U6383 ( .A(out[1255]), .B(n1614), .Z(N1267) );
  AND U6384 ( .A(out[1256]), .B(n1614), .Z(N1268) );
  AND U6385 ( .A(out[1257]), .B(n1614), .Z(N1269) );
  AND U6386 ( .A(out[115]), .B(n1614), .Z(N127) );
  AND U6387 ( .A(out[1258]), .B(n1614), .Z(N1270) );
  AND U6388 ( .A(out[1259]), .B(n1614), .Z(N1271) );
  AND U6389 ( .A(out[1260]), .B(n1614), .Z(N1272) );
  AND U6390 ( .A(out[1261]), .B(n1614), .Z(N1273) );
  AND U6391 ( .A(out[1262]), .B(n1614), .Z(N1274) );
  AND U6392 ( .A(out[1263]), .B(n1614), .Z(N1275) );
  AND U6393 ( .A(out[1264]), .B(n1614), .Z(N1276) );
  AND U6394 ( .A(out[1265]), .B(n1614), .Z(N1277) );
  AND U6395 ( .A(out[1266]), .B(n1614), .Z(N1278) );
  AND U6396 ( .A(out[1267]), .B(n1614), .Z(N1279) );
  AND U6397 ( .A(out[116]), .B(n1614), .Z(N128) );
  AND U6398 ( .A(out[1268]), .B(n1614), .Z(N1280) );
  AND U6399 ( .A(out[1269]), .B(n1614), .Z(N1281) );
  AND U6400 ( .A(out[1270]), .B(n1614), .Z(N1282) );
  AND U6401 ( .A(out[1271]), .B(n1614), .Z(N1283) );
  AND U6402 ( .A(out[1272]), .B(n1614), .Z(N1284) );
  AND U6403 ( .A(out[1273]), .B(n1614), .Z(N1285) );
  AND U6404 ( .A(out[1274]), .B(n1614), .Z(N1286) );
  AND U6405 ( .A(out[1275]), .B(n1614), .Z(N1287) );
  AND U6406 ( .A(out[1276]), .B(n1614), .Z(N1288) );
  AND U6407 ( .A(out[1277]), .B(n1614), .Z(N1289) );
  AND U6408 ( .A(out[117]), .B(n1614), .Z(N129) );
  AND U6409 ( .A(out[1278]), .B(n1614), .Z(N1290) );
  AND U6410 ( .A(out[1279]), .B(n1614), .Z(N1291) );
  AND U6411 ( .A(out[1280]), .B(n1614), .Z(N1292) );
  AND U6412 ( .A(out[1281]), .B(n1614), .Z(N1293) );
  AND U6413 ( .A(out[1282]), .B(n1614), .Z(N1294) );
  AND U6414 ( .A(out[1283]), .B(n1614), .Z(N1295) );
  AND U6415 ( .A(out[1284]), .B(n1614), .Z(N1296) );
  AND U6416 ( .A(out[1285]), .B(n1614), .Z(N1297) );
  AND U6417 ( .A(out[1286]), .B(n1614), .Z(N1298) );
  AND U6418 ( .A(out[1287]), .B(n1614), .Z(N1299) );
  AND U6419 ( .A(out[1]), .B(n1614), .Z(N13) );
  AND U6420 ( .A(out[118]), .B(n1614), .Z(N130) );
  AND U6421 ( .A(out[1288]), .B(n1614), .Z(N1300) );
  AND U6422 ( .A(out[1289]), .B(n1614), .Z(N1301) );
  AND U6423 ( .A(out[1290]), .B(n1614), .Z(N1302) );
  AND U6424 ( .A(out[1291]), .B(n1614), .Z(N1303) );
  AND U6425 ( .A(out[1292]), .B(n1614), .Z(N1304) );
  AND U6426 ( .A(out[1293]), .B(n1614), .Z(N1305) );
  AND U6427 ( .A(out[1294]), .B(n1614), .Z(N1306) );
  AND U6428 ( .A(out[1295]), .B(n1614), .Z(N1307) );
  AND U6429 ( .A(out[1296]), .B(n1614), .Z(N1308) );
  AND U6430 ( .A(out[1297]), .B(n1614), .Z(N1309) );
  AND U6431 ( .A(out[119]), .B(n1614), .Z(N131) );
  AND U6432 ( .A(out[1298]), .B(n1614), .Z(N1310) );
  AND U6433 ( .A(out[1299]), .B(n1614), .Z(N1311) );
  AND U6434 ( .A(out[1300]), .B(n1614), .Z(N1312) );
  AND U6435 ( .A(out[1301]), .B(n1614), .Z(N1313) );
  AND U6436 ( .A(out[1302]), .B(n1614), .Z(N1314) );
  AND U6437 ( .A(out[1303]), .B(n1614), .Z(N1315) );
  AND U6438 ( .A(out[1304]), .B(n1614), .Z(N1316) );
  AND U6439 ( .A(out[1305]), .B(n1614), .Z(N1317) );
  AND U6440 ( .A(out[1306]), .B(n1614), .Z(N1318) );
  AND U6441 ( .A(out[1307]), .B(n1614), .Z(N1319) );
  AND U6442 ( .A(out[120]), .B(n1614), .Z(N132) );
  AND U6443 ( .A(out[1308]), .B(n1614), .Z(N1320) );
  AND U6444 ( .A(out[1309]), .B(n1614), .Z(N1321) );
  AND U6445 ( .A(out[1310]), .B(n1614), .Z(N1322) );
  AND U6446 ( .A(out[1311]), .B(n1614), .Z(N1323) );
  AND U6447 ( .A(out[1312]), .B(n1614), .Z(N1324) );
  AND U6448 ( .A(out[1313]), .B(n1614), .Z(N1325) );
  AND U6449 ( .A(out[1314]), .B(n1614), .Z(N1326) );
  AND U6450 ( .A(out[1315]), .B(n1614), .Z(N1327) );
  AND U6451 ( .A(out[1316]), .B(n1614), .Z(N1328) );
  AND U6452 ( .A(out[1317]), .B(n1614), .Z(N1329) );
  AND U6453 ( .A(out[121]), .B(n1614), .Z(N133) );
  AND U6454 ( .A(out[1318]), .B(n1614), .Z(N1330) );
  AND U6455 ( .A(out[1319]), .B(n1614), .Z(N1331) );
  AND U6456 ( .A(out[1320]), .B(n1614), .Z(N1332) );
  AND U6457 ( .A(out[1321]), .B(n1614), .Z(N1333) );
  AND U6458 ( .A(out[1322]), .B(n1614), .Z(N1334) );
  AND U6459 ( .A(out[1323]), .B(n1614), .Z(N1335) );
  AND U6460 ( .A(out[1324]), .B(n1614), .Z(N1336) );
  AND U6461 ( .A(out[1325]), .B(n1614), .Z(N1337) );
  AND U6462 ( .A(out[1326]), .B(n1614), .Z(N1338) );
  AND U6463 ( .A(out[1327]), .B(n1614), .Z(N1339) );
  AND U6464 ( .A(out[122]), .B(n1614), .Z(N134) );
  AND U6465 ( .A(out[1328]), .B(n1614), .Z(N1340) );
  AND U6466 ( .A(out[1329]), .B(n1614), .Z(N1341) );
  AND U6467 ( .A(out[1330]), .B(n1614), .Z(N1342) );
  AND U6468 ( .A(out[1331]), .B(n1614), .Z(N1343) );
  AND U6469 ( .A(out[1332]), .B(n1614), .Z(N1344) );
  AND U6470 ( .A(out[1333]), .B(n1614), .Z(N1345) );
  AND U6471 ( .A(out[1334]), .B(n1614), .Z(N1346) );
  AND U6472 ( .A(out[1335]), .B(n1614), .Z(N1347) );
  AND U6473 ( .A(out[1336]), .B(n1614), .Z(N1348) );
  AND U6474 ( .A(out[1337]), .B(n1614), .Z(N1349) );
  AND U6475 ( .A(out[123]), .B(n1614), .Z(N135) );
  AND U6476 ( .A(out[1338]), .B(n1614), .Z(N1350) );
  AND U6477 ( .A(out[1339]), .B(n1614), .Z(N1351) );
  AND U6478 ( .A(out[1340]), .B(n1614), .Z(N1352) );
  AND U6479 ( .A(out[1341]), .B(n1614), .Z(N1353) );
  AND U6480 ( .A(out[1342]), .B(n1614), .Z(N1354) );
  AND U6481 ( .A(out[1343]), .B(n1614), .Z(N1355) );
  AND U6482 ( .A(out[1344]), .B(n1614), .Z(N1356) );
  AND U6483 ( .A(out[1345]), .B(n1614), .Z(N1357) );
  AND U6484 ( .A(out[1346]), .B(n1614), .Z(N1358) );
  AND U6485 ( .A(out[1347]), .B(n1614), .Z(N1359) );
  AND U6486 ( .A(out[124]), .B(n1614), .Z(N136) );
  AND U6487 ( .A(out[1348]), .B(n1614), .Z(N1360) );
  AND U6488 ( .A(out[1349]), .B(n1614), .Z(N1361) );
  AND U6489 ( .A(out[1350]), .B(n1614), .Z(N1362) );
  AND U6490 ( .A(out[1351]), .B(n1614), .Z(N1363) );
  AND U6491 ( .A(out[1352]), .B(n1614), .Z(N1364) );
  AND U6492 ( .A(out[1353]), .B(n1614), .Z(N1365) );
  AND U6493 ( .A(out[1354]), .B(n1614), .Z(N1366) );
  AND U6494 ( .A(out[1355]), .B(n1614), .Z(N1367) );
  AND U6495 ( .A(out[1356]), .B(n1614), .Z(N1368) );
  AND U6496 ( .A(out[1357]), .B(n1614), .Z(N1369) );
  AND U6497 ( .A(out[125]), .B(n1614), .Z(N137) );
  AND U6498 ( .A(out[1358]), .B(n1614), .Z(N1370) );
  AND U6499 ( .A(out[1359]), .B(n1614), .Z(N1371) );
  AND U6500 ( .A(out[1360]), .B(n1614), .Z(N1372) );
  AND U6501 ( .A(out[1361]), .B(n1614), .Z(N1373) );
  AND U6502 ( .A(out[1362]), .B(n1614), .Z(N1374) );
  AND U6503 ( .A(out[1363]), .B(n1614), .Z(N1375) );
  AND U6504 ( .A(out[1364]), .B(n1614), .Z(N1376) );
  AND U6505 ( .A(out[1365]), .B(n1614), .Z(N1377) );
  AND U6506 ( .A(out[1366]), .B(n1614), .Z(N1378) );
  AND U6507 ( .A(out[1367]), .B(n1614), .Z(N1379) );
  AND U6508 ( .A(out[126]), .B(n1614), .Z(N138) );
  AND U6509 ( .A(out[1368]), .B(n1614), .Z(N1380) );
  AND U6510 ( .A(out[1369]), .B(n1614), .Z(N1381) );
  AND U6511 ( .A(out[1370]), .B(n1614), .Z(N1382) );
  AND U6512 ( .A(out[1371]), .B(n1614), .Z(N1383) );
  AND U6513 ( .A(out[1372]), .B(n1614), .Z(N1384) );
  AND U6514 ( .A(out[1373]), .B(n1614), .Z(N1385) );
  AND U6515 ( .A(out[1374]), .B(n1614), .Z(N1386) );
  AND U6516 ( .A(out[1375]), .B(n1614), .Z(N1387) );
  AND U6517 ( .A(out[1376]), .B(n1614), .Z(N1388) );
  AND U6518 ( .A(out[1377]), .B(n1614), .Z(N1389) );
  AND U6519 ( .A(out[127]), .B(n1614), .Z(N139) );
  AND U6520 ( .A(out[1378]), .B(n1614), .Z(N1390) );
  AND U6521 ( .A(out[1379]), .B(n1614), .Z(N1391) );
  AND U6522 ( .A(out[1380]), .B(n1614), .Z(N1392) );
  AND U6523 ( .A(out[1381]), .B(n1614), .Z(N1393) );
  AND U6524 ( .A(out[1382]), .B(n1614), .Z(N1394) );
  AND U6525 ( .A(out[1383]), .B(n1614), .Z(N1395) );
  AND U6526 ( .A(out[1384]), .B(n1614), .Z(N1396) );
  AND U6527 ( .A(out[1385]), .B(n1614), .Z(N1397) );
  AND U6528 ( .A(out[1386]), .B(n1614), .Z(N1398) );
  AND U6529 ( .A(out[1387]), .B(n1614), .Z(N1399) );
  AND U6530 ( .A(out[2]), .B(n1614), .Z(N14) );
  AND U6531 ( .A(out[128]), .B(n1614), .Z(N140) );
  AND U6532 ( .A(out[1388]), .B(n1614), .Z(N1400) );
  AND U6533 ( .A(out[1389]), .B(n1614), .Z(N1401) );
  AND U6534 ( .A(out[1390]), .B(n1614), .Z(N1402) );
  AND U6535 ( .A(out[1391]), .B(n1614), .Z(N1403) );
  AND U6536 ( .A(out[1392]), .B(n1614), .Z(N1404) );
  AND U6537 ( .A(out[1393]), .B(n1614), .Z(N1405) );
  AND U6538 ( .A(out[1394]), .B(n1614), .Z(N1406) );
  AND U6539 ( .A(out[1395]), .B(n1614), .Z(N1407) );
  AND U6540 ( .A(out[1396]), .B(n1614), .Z(N1408) );
  AND U6541 ( .A(out[1397]), .B(n1614), .Z(N1409) );
  AND U6542 ( .A(out[129]), .B(n1614), .Z(N141) );
  AND U6543 ( .A(out[1398]), .B(n1614), .Z(N1410) );
  AND U6544 ( .A(out[1399]), .B(n1614), .Z(N1411) );
  AND U6545 ( .A(out[1400]), .B(n1614), .Z(N1412) );
  AND U6546 ( .A(out[1401]), .B(n1614), .Z(N1413) );
  AND U6547 ( .A(out[1402]), .B(n1614), .Z(N1414) );
  AND U6548 ( .A(out[1403]), .B(n1614), .Z(N1415) );
  AND U6549 ( .A(out[1404]), .B(n1614), .Z(N1416) );
  AND U6550 ( .A(out[1405]), .B(n1614), .Z(N1417) );
  AND U6551 ( .A(out[1406]), .B(n1614), .Z(N1418) );
  AND U6552 ( .A(out[1407]), .B(n1614), .Z(N1419) );
  AND U6553 ( .A(out[130]), .B(n1614), .Z(N142) );
  AND U6554 ( .A(out[1408]), .B(n1614), .Z(N1420) );
  AND U6555 ( .A(out[1409]), .B(n1614), .Z(N1421) );
  AND U6556 ( .A(out[1410]), .B(n1614), .Z(N1422) );
  AND U6557 ( .A(out[1411]), .B(n1614), .Z(N1423) );
  AND U6558 ( .A(out[1412]), .B(n1614), .Z(N1424) );
  AND U6559 ( .A(out[1413]), .B(n1614), .Z(N1425) );
  AND U6560 ( .A(out[1414]), .B(n1614), .Z(N1426) );
  AND U6561 ( .A(out[1415]), .B(n1614), .Z(N1427) );
  AND U6562 ( .A(out[1416]), .B(n1614), .Z(N1428) );
  AND U6563 ( .A(out[1417]), .B(n1614), .Z(N1429) );
  AND U6564 ( .A(out[131]), .B(n1614), .Z(N143) );
  AND U6565 ( .A(out[1418]), .B(n1614), .Z(N1430) );
  AND U6566 ( .A(out[1419]), .B(n1614), .Z(N1431) );
  AND U6567 ( .A(out[1420]), .B(n1614), .Z(N1432) );
  AND U6568 ( .A(out[1421]), .B(n1614), .Z(N1433) );
  AND U6569 ( .A(out[1422]), .B(n1614), .Z(N1434) );
  AND U6570 ( .A(out[1423]), .B(n1614), .Z(N1435) );
  AND U6571 ( .A(out[1424]), .B(n1614), .Z(N1436) );
  AND U6572 ( .A(out[1425]), .B(n1614), .Z(N1437) );
  AND U6573 ( .A(out[1426]), .B(n1614), .Z(N1438) );
  AND U6574 ( .A(out[1427]), .B(n1614), .Z(N1439) );
  AND U6575 ( .A(out[132]), .B(n1614), .Z(N144) );
  AND U6576 ( .A(out[1428]), .B(n1614), .Z(N1440) );
  AND U6577 ( .A(out[1429]), .B(n1614), .Z(N1441) );
  AND U6578 ( .A(out[1430]), .B(n1614), .Z(N1442) );
  AND U6579 ( .A(out[1431]), .B(n1614), .Z(N1443) );
  AND U6580 ( .A(out[1432]), .B(n1614), .Z(N1444) );
  AND U6581 ( .A(out[1433]), .B(n1614), .Z(N1445) );
  AND U6582 ( .A(out[1434]), .B(n1614), .Z(N1446) );
  AND U6583 ( .A(out[1435]), .B(n1614), .Z(N1447) );
  AND U6584 ( .A(out[1436]), .B(n1614), .Z(N1448) );
  AND U6585 ( .A(out[1437]), .B(n1614), .Z(N1449) );
  AND U6586 ( .A(out[133]), .B(n1614), .Z(N145) );
  AND U6587 ( .A(out[1438]), .B(n1614), .Z(N1450) );
  AND U6588 ( .A(out[1439]), .B(n1614), .Z(N1451) );
  AND U6589 ( .A(out[1440]), .B(n1614), .Z(N1452) );
  AND U6590 ( .A(out[1441]), .B(n1614), .Z(N1453) );
  AND U6591 ( .A(out[1442]), .B(n1614), .Z(N1454) );
  AND U6592 ( .A(out[1443]), .B(n1614), .Z(N1455) );
  AND U6593 ( .A(out[1444]), .B(n1614), .Z(N1456) );
  AND U6594 ( .A(out[1445]), .B(n1614), .Z(N1457) );
  AND U6595 ( .A(out[1446]), .B(n1614), .Z(N1458) );
  AND U6596 ( .A(out[1447]), .B(n1614), .Z(N1459) );
  AND U6597 ( .A(out[134]), .B(n1614), .Z(N146) );
  AND U6598 ( .A(out[1448]), .B(n1614), .Z(N1460) );
  AND U6599 ( .A(out[1449]), .B(n1614), .Z(N1461) );
  AND U6600 ( .A(out[1450]), .B(n1614), .Z(N1462) );
  AND U6601 ( .A(out[1451]), .B(n1614), .Z(N1463) );
  AND U6602 ( .A(out[1452]), .B(n1614), .Z(N1464) );
  AND U6603 ( .A(out[1453]), .B(n1614), .Z(N1465) );
  AND U6604 ( .A(out[1454]), .B(n1614), .Z(N1466) );
  AND U6605 ( .A(out[1455]), .B(n1614), .Z(N1467) );
  AND U6606 ( .A(out[1456]), .B(n1614), .Z(N1468) );
  AND U6607 ( .A(out[1457]), .B(n1614), .Z(N1469) );
  AND U6608 ( .A(out[135]), .B(n1614), .Z(N147) );
  AND U6609 ( .A(out[1458]), .B(n1614), .Z(N1470) );
  AND U6610 ( .A(out[1459]), .B(n1614), .Z(N1471) );
  AND U6611 ( .A(out[1460]), .B(n1614), .Z(N1472) );
  AND U6612 ( .A(out[1461]), .B(n1614), .Z(N1473) );
  AND U6613 ( .A(out[1462]), .B(n1614), .Z(N1474) );
  AND U6614 ( .A(out[1463]), .B(n1614), .Z(N1475) );
  AND U6615 ( .A(out[1464]), .B(n1614), .Z(N1476) );
  AND U6616 ( .A(out[1465]), .B(n1614), .Z(N1477) );
  AND U6617 ( .A(out[1466]), .B(n1614), .Z(N1478) );
  AND U6618 ( .A(out[1467]), .B(n1614), .Z(N1479) );
  AND U6619 ( .A(out[136]), .B(n1614), .Z(N148) );
  AND U6620 ( .A(out[1468]), .B(n1614), .Z(N1480) );
  AND U6621 ( .A(out[1469]), .B(n1614), .Z(N1481) );
  AND U6622 ( .A(out[1470]), .B(n1614), .Z(N1482) );
  AND U6623 ( .A(out[1471]), .B(n1614), .Z(N1483) );
  AND U6624 ( .A(out[1472]), .B(n1614), .Z(N1484) );
  AND U6625 ( .A(out[1473]), .B(n1614), .Z(N1485) );
  AND U6626 ( .A(out[1474]), .B(n1614), .Z(N1486) );
  AND U6627 ( .A(out[1475]), .B(n1614), .Z(N1487) );
  AND U6628 ( .A(out[1476]), .B(n1614), .Z(N1488) );
  AND U6629 ( .A(out[1477]), .B(n1614), .Z(N1489) );
  AND U6630 ( .A(out[137]), .B(n1614), .Z(N149) );
  AND U6631 ( .A(out[1478]), .B(n1614), .Z(N1490) );
  AND U6632 ( .A(out[1479]), .B(n1614), .Z(N1491) );
  AND U6633 ( .A(out[1480]), .B(n1614), .Z(N1492) );
  AND U6634 ( .A(out[1481]), .B(n1614), .Z(N1493) );
  AND U6635 ( .A(out[1482]), .B(n1614), .Z(N1494) );
  AND U6636 ( .A(out[1483]), .B(n1614), .Z(N1495) );
  AND U6637 ( .A(out[1484]), .B(n1614), .Z(N1496) );
  AND U6638 ( .A(out[1485]), .B(n1614), .Z(N1497) );
  AND U6639 ( .A(out[1486]), .B(n1614), .Z(N1498) );
  AND U6640 ( .A(out[1487]), .B(n1614), .Z(N1499) );
  AND U6641 ( .A(out[3]), .B(n1614), .Z(N15) );
  AND U6642 ( .A(out[138]), .B(n1614), .Z(N150) );
  AND U6643 ( .A(out[1488]), .B(n1614), .Z(N1500) );
  AND U6644 ( .A(out[1489]), .B(n1614), .Z(N1501) );
  AND U6645 ( .A(out[1490]), .B(n1614), .Z(N1502) );
  AND U6646 ( .A(out[1491]), .B(n1614), .Z(N1503) );
  AND U6647 ( .A(out[1492]), .B(n1614), .Z(N1504) );
  AND U6648 ( .A(out[1493]), .B(n1614), .Z(N1505) );
  AND U6649 ( .A(out[1494]), .B(n1614), .Z(N1506) );
  AND U6650 ( .A(out[1495]), .B(n1614), .Z(N1507) );
  AND U6651 ( .A(out[1496]), .B(n1614), .Z(N1508) );
  AND U6652 ( .A(out[1497]), .B(n1614), .Z(N1509) );
  AND U6653 ( .A(out[139]), .B(n1614), .Z(N151) );
  AND U6654 ( .A(out[1498]), .B(n1614), .Z(N1510) );
  AND U6655 ( .A(out[1499]), .B(n1614), .Z(N1511) );
  AND U6656 ( .A(out[1500]), .B(n1614), .Z(N1512) );
  AND U6657 ( .A(out[1501]), .B(n1614), .Z(N1513) );
  AND U6658 ( .A(out[1502]), .B(n1614), .Z(N1514) );
  AND U6659 ( .A(out[1503]), .B(n1614), .Z(N1515) );
  AND U6660 ( .A(out[1504]), .B(n1614), .Z(N1516) );
  AND U6661 ( .A(out[1505]), .B(n1614), .Z(N1517) );
  AND U6662 ( .A(out[1506]), .B(n1614), .Z(N1518) );
  AND U6663 ( .A(out[1507]), .B(n1614), .Z(N1519) );
  AND U6664 ( .A(out[140]), .B(n1614), .Z(N152) );
  AND U6665 ( .A(out[1508]), .B(n1614), .Z(N1520) );
  AND U6666 ( .A(out[1509]), .B(n1614), .Z(N1521) );
  AND U6667 ( .A(out[1510]), .B(n1614), .Z(N1522) );
  AND U6668 ( .A(out[1511]), .B(n1614), .Z(N1523) );
  AND U6669 ( .A(out[1512]), .B(n1614), .Z(N1524) );
  AND U6670 ( .A(out[1513]), .B(n1614), .Z(N1525) );
  AND U6671 ( .A(out[1514]), .B(n1614), .Z(N1526) );
  AND U6672 ( .A(out[1515]), .B(n1614), .Z(N1527) );
  AND U6673 ( .A(out[1516]), .B(n1614), .Z(N1528) );
  AND U6674 ( .A(out[1517]), .B(n1614), .Z(N1529) );
  AND U6675 ( .A(out[141]), .B(n1614), .Z(N153) );
  AND U6676 ( .A(out[1518]), .B(n1614), .Z(N1530) );
  AND U6677 ( .A(out[1519]), .B(n1614), .Z(N1531) );
  AND U6678 ( .A(out[1520]), .B(n1614), .Z(N1532) );
  AND U6679 ( .A(out[1521]), .B(n1614), .Z(N1533) );
  AND U6680 ( .A(out[1522]), .B(n1614), .Z(N1534) );
  AND U6681 ( .A(out[1523]), .B(n1614), .Z(N1535) );
  AND U6682 ( .A(out[1524]), .B(n1614), .Z(N1536) );
  AND U6683 ( .A(out[1525]), .B(n1614), .Z(N1537) );
  AND U6684 ( .A(out[1526]), .B(n1614), .Z(N1538) );
  AND U6685 ( .A(out[1527]), .B(n1614), .Z(N1539) );
  AND U6686 ( .A(out[142]), .B(n1614), .Z(N154) );
  AND U6687 ( .A(out[1528]), .B(n1614), .Z(N1540) );
  AND U6688 ( .A(out[1529]), .B(n1614), .Z(N1541) );
  AND U6689 ( .A(out[1530]), .B(n1614), .Z(N1542) );
  AND U6690 ( .A(out[1531]), .B(n1614), .Z(N1543) );
  AND U6691 ( .A(out[1532]), .B(n1614), .Z(N1544) );
  AND U6692 ( .A(out[1533]), .B(n1614), .Z(N1545) );
  AND U6693 ( .A(out[1534]), .B(n1614), .Z(N1546) );
  AND U6694 ( .A(out[1535]), .B(n1614), .Z(N1547) );
  AND U6695 ( .A(out[1536]), .B(n1614), .Z(N1548) );
  AND U6696 ( .A(out[1537]), .B(n1614), .Z(N1549) );
  AND U6697 ( .A(out[143]), .B(n1614), .Z(N155) );
  AND U6698 ( .A(out[1538]), .B(n1614), .Z(N1550) );
  AND U6699 ( .A(out[1539]), .B(n1614), .Z(N1551) );
  AND U6700 ( .A(out[1540]), .B(n1614), .Z(N1552) );
  AND U6701 ( .A(out[1541]), .B(n1614), .Z(N1553) );
  AND U6702 ( .A(out[1542]), .B(n1614), .Z(N1554) );
  AND U6703 ( .A(out[1543]), .B(n1614), .Z(N1555) );
  AND U6704 ( .A(out[1544]), .B(n1614), .Z(N1556) );
  AND U6705 ( .A(out[1545]), .B(n1614), .Z(N1557) );
  AND U6706 ( .A(out[1546]), .B(n1614), .Z(N1558) );
  AND U6707 ( .A(out[1547]), .B(n1614), .Z(N1559) );
  AND U6708 ( .A(out[144]), .B(n1614), .Z(N156) );
  AND U6709 ( .A(out[1548]), .B(n1614), .Z(N1560) );
  AND U6710 ( .A(out[1549]), .B(n1614), .Z(N1561) );
  AND U6711 ( .A(out[1550]), .B(n1614), .Z(N1562) );
  AND U6712 ( .A(out[1551]), .B(n1614), .Z(N1563) );
  AND U6713 ( .A(out[1552]), .B(n1614), .Z(N1564) );
  AND U6714 ( .A(out[1553]), .B(n1614), .Z(N1565) );
  AND U6715 ( .A(out[1554]), .B(n1614), .Z(N1566) );
  AND U6716 ( .A(out[1555]), .B(n1614), .Z(N1567) );
  AND U6717 ( .A(out[1556]), .B(n1614), .Z(N1568) );
  AND U6718 ( .A(out[1557]), .B(n1614), .Z(N1569) );
  AND U6719 ( .A(out[145]), .B(n1614), .Z(N157) );
  AND U6720 ( .A(out[1558]), .B(n1614), .Z(N1570) );
  AND U6721 ( .A(out[1559]), .B(n1614), .Z(N1571) );
  AND U6722 ( .A(out[1560]), .B(n1614), .Z(N1572) );
  AND U6723 ( .A(out[1561]), .B(n1614), .Z(N1573) );
  AND U6724 ( .A(out[1562]), .B(n1614), .Z(N1574) );
  AND U6725 ( .A(out[1563]), .B(n1614), .Z(N1575) );
  AND U6726 ( .A(out[1564]), .B(n1614), .Z(N1576) );
  AND U6727 ( .A(out[1565]), .B(n1614), .Z(N1577) );
  AND U6728 ( .A(out[1566]), .B(n1614), .Z(N1578) );
  AND U6729 ( .A(out[1567]), .B(n1614), .Z(N1579) );
  AND U6730 ( .A(out[146]), .B(n1614), .Z(N158) );
  AND U6731 ( .A(out[1568]), .B(n1614), .Z(N1580) );
  AND U6732 ( .A(out[1569]), .B(n1614), .Z(N1581) );
  AND U6733 ( .A(out[1570]), .B(n1614), .Z(N1582) );
  AND U6734 ( .A(out[1571]), .B(n1614), .Z(N1583) );
  AND U6735 ( .A(out[1572]), .B(n1614), .Z(N1584) );
  AND U6736 ( .A(out[1573]), .B(n1614), .Z(N1585) );
  AND U6737 ( .A(out[1574]), .B(n1614), .Z(N1586) );
  AND U6738 ( .A(out[1575]), .B(n1614), .Z(N1587) );
  AND U6739 ( .A(out[1576]), .B(n1614), .Z(N1588) );
  AND U6740 ( .A(out[1577]), .B(n1614), .Z(N1589) );
  AND U6741 ( .A(out[147]), .B(n1614), .Z(N159) );
  AND U6742 ( .A(out[1578]), .B(n1614), .Z(N1590) );
  AND U6743 ( .A(out[1579]), .B(n1614), .Z(N1591) );
  AND U6744 ( .A(out[1580]), .B(n1614), .Z(N1592) );
  AND U6745 ( .A(out[1581]), .B(n1614), .Z(N1593) );
  AND U6746 ( .A(out[1582]), .B(n1614), .Z(N1594) );
  AND U6747 ( .A(out[1583]), .B(n1614), .Z(N1595) );
  AND U6748 ( .A(out[1584]), .B(n1614), .Z(N1596) );
  AND U6749 ( .A(out[1585]), .B(n1614), .Z(N1597) );
  AND U6750 ( .A(out[1586]), .B(n1614), .Z(N1598) );
  AND U6751 ( .A(out[1587]), .B(n1614), .Z(N1599) );
  AND U6752 ( .A(out[4]), .B(n1614), .Z(N16) );
  AND U6753 ( .A(out[148]), .B(n1614), .Z(N160) );
  AND U6754 ( .A(out[1588]), .B(n1614), .Z(N1600) );
  AND U6755 ( .A(out[1589]), .B(n1614), .Z(N1601) );
  AND U6756 ( .A(out[1590]), .B(n1614), .Z(N1602) );
  AND U6757 ( .A(out[1591]), .B(n1614), .Z(N1603) );
  AND U6758 ( .A(out[1592]), .B(n1614), .Z(N1604) );
  AND U6759 ( .A(out[1593]), .B(n1614), .Z(N1605) );
  AND U6760 ( .A(out[1594]), .B(n1614), .Z(N1606) );
  AND U6761 ( .A(out[1595]), .B(n1614), .Z(N1607) );
  AND U6762 ( .A(out[1596]), .B(n1614), .Z(N1608) );
  AND U6763 ( .A(out[1597]), .B(n1614), .Z(N1609) );
  AND U6764 ( .A(out[149]), .B(n1614), .Z(N161) );
  AND U6765 ( .A(out[1598]), .B(n1614), .Z(N1610) );
  AND U6766 ( .A(out[1599]), .B(n1614), .Z(N1611) );
  AND U6767 ( .A(out[150]), .B(n1614), .Z(N162) );
  AND U6768 ( .A(out[151]), .B(n1614), .Z(N163) );
  AND U6769 ( .A(out[152]), .B(n1614), .Z(N164) );
  AND U6770 ( .A(out[153]), .B(n1614), .Z(N165) );
  AND U6771 ( .A(out[154]), .B(n1614), .Z(N166) );
  AND U6772 ( .A(out[155]), .B(n1614), .Z(N167) );
  AND U6773 ( .A(out[156]), .B(n1614), .Z(N168) );
  AND U6774 ( .A(out[157]), .B(n1614), .Z(N169) );
  AND U6775 ( .A(out[5]), .B(n1614), .Z(N17) );
  AND U6776 ( .A(out[158]), .B(n1614), .Z(N170) );
  AND U6777 ( .A(out[159]), .B(n1614), .Z(N171) );
  AND U6778 ( .A(out[160]), .B(n1614), .Z(N172) );
  AND U6779 ( .A(out[161]), .B(n1614), .Z(N173) );
  AND U6780 ( .A(out[162]), .B(n1614), .Z(N174) );
  AND U6781 ( .A(out[163]), .B(n1614), .Z(N175) );
  AND U6782 ( .A(out[164]), .B(n1614), .Z(N176) );
  AND U6783 ( .A(out[165]), .B(n1614), .Z(N177) );
  AND U6784 ( .A(out[166]), .B(n1614), .Z(N178) );
  AND U6785 ( .A(out[167]), .B(n1614), .Z(N179) );
  AND U6786 ( .A(out[6]), .B(n1614), .Z(N18) );
  AND U6787 ( .A(out[168]), .B(n1614), .Z(N180) );
  AND U6788 ( .A(out[169]), .B(n1614), .Z(N181) );
  AND U6789 ( .A(out[170]), .B(n1614), .Z(N182) );
  AND U6790 ( .A(out[171]), .B(n1614), .Z(N183) );
  AND U6791 ( .A(out[172]), .B(n1614), .Z(N184) );
  AND U6792 ( .A(out[173]), .B(n1614), .Z(N185) );
  AND U6793 ( .A(out[174]), .B(n1614), .Z(N186) );
  AND U6794 ( .A(out[175]), .B(n1614), .Z(N187) );
  AND U6795 ( .A(out[176]), .B(n1614), .Z(N188) );
  AND U6796 ( .A(out[177]), .B(n1614), .Z(N189) );
  AND U6797 ( .A(out[7]), .B(n1614), .Z(N19) );
  AND U6798 ( .A(out[178]), .B(n1614), .Z(N190) );
  AND U6799 ( .A(out[179]), .B(n1614), .Z(N191) );
  AND U6800 ( .A(out[180]), .B(n1614), .Z(N192) );
  AND U6801 ( .A(out[181]), .B(n1614), .Z(N193) );
  AND U6802 ( .A(out[182]), .B(n1614), .Z(N194) );
  AND U6803 ( .A(out[183]), .B(n1614), .Z(N195) );
  AND U6804 ( .A(out[184]), .B(n1614), .Z(N196) );
  AND U6805 ( .A(out[185]), .B(n1614), .Z(N197) );
  AND U6806 ( .A(out[186]), .B(n1614), .Z(N198) );
  AND U6807 ( .A(out[187]), .B(n1614), .Z(N199) );
  AND U6808 ( .A(out[8]), .B(n1614), .Z(N20) );
  AND U6809 ( .A(out[188]), .B(n1614), .Z(N200) );
  AND U6810 ( .A(out[189]), .B(n1614), .Z(N201) );
  AND U6811 ( .A(out[190]), .B(n1614), .Z(N202) );
  AND U6812 ( .A(out[191]), .B(n1614), .Z(N203) );
  AND U6813 ( .A(out[192]), .B(n1614), .Z(N204) );
  AND U6814 ( .A(out[193]), .B(n1614), .Z(N205) );
  AND U6815 ( .A(out[194]), .B(n1614), .Z(N206) );
  AND U6816 ( .A(out[195]), .B(n1614), .Z(N207) );
  AND U6817 ( .A(out[196]), .B(n1614), .Z(N208) );
  AND U6818 ( .A(out[197]), .B(n1614), .Z(N209) );
  AND U6819 ( .A(out[9]), .B(n1614), .Z(N21) );
  AND U6820 ( .A(out[198]), .B(n1614), .Z(N210) );
  AND U6821 ( .A(out[199]), .B(n1614), .Z(N211) );
  AND U6822 ( .A(out[200]), .B(n1614), .Z(N212) );
  AND U6823 ( .A(out[201]), .B(n1614), .Z(N213) );
  AND U6824 ( .A(out[202]), .B(n1614), .Z(N214) );
  AND U6825 ( .A(out[203]), .B(n1614), .Z(N215) );
  AND U6826 ( .A(out[204]), .B(n1614), .Z(N216) );
  AND U6827 ( .A(out[205]), .B(n1614), .Z(N217) );
  AND U6828 ( .A(out[206]), .B(n1614), .Z(N218) );
  AND U6829 ( .A(out[207]), .B(n1614), .Z(N219) );
  AND U6830 ( .A(out[10]), .B(n1614), .Z(N22) );
  AND U6831 ( .A(out[208]), .B(n1614), .Z(N220) );
  AND U6832 ( .A(out[209]), .B(n1614), .Z(N221) );
  AND U6833 ( .A(out[210]), .B(n1614), .Z(N222) );
  AND U6834 ( .A(out[211]), .B(n1614), .Z(N223) );
  AND U6835 ( .A(out[212]), .B(n1614), .Z(N224) );
  AND U6836 ( .A(out[213]), .B(n1614), .Z(N225) );
  AND U6837 ( .A(out[214]), .B(n1614), .Z(N226) );
  AND U6838 ( .A(out[215]), .B(n1614), .Z(N227) );
  AND U6839 ( .A(out[216]), .B(n1614), .Z(N228) );
  AND U6840 ( .A(out[217]), .B(n1614), .Z(N229) );
  AND U6841 ( .A(out[11]), .B(n1614), .Z(N23) );
  AND U6842 ( .A(out[218]), .B(n1614), .Z(N230) );
  AND U6843 ( .A(out[219]), .B(n1614), .Z(N231) );
  AND U6844 ( .A(out[220]), .B(n1614), .Z(N232) );
  AND U6845 ( .A(out[221]), .B(n1614), .Z(N233) );
  AND U6846 ( .A(out[222]), .B(n1614), .Z(N234) );
  AND U6847 ( .A(out[223]), .B(n1614), .Z(N235) );
  AND U6848 ( .A(out[224]), .B(n1614), .Z(N236) );
  AND U6849 ( .A(out[225]), .B(n1614), .Z(N237) );
  AND U6850 ( .A(out[226]), .B(n1614), .Z(N238) );
  AND U6851 ( .A(out[227]), .B(n1614), .Z(N239) );
  AND U6852 ( .A(out[12]), .B(n1614), .Z(N24) );
  AND U6853 ( .A(out[228]), .B(n1614), .Z(N240) );
  AND U6854 ( .A(out[229]), .B(n1614), .Z(N241) );
  AND U6855 ( .A(out[230]), .B(n1614), .Z(N242) );
  AND U6856 ( .A(out[231]), .B(n1614), .Z(N243) );
  AND U6857 ( .A(out[232]), .B(n1614), .Z(N244) );
  AND U6858 ( .A(out[233]), .B(n1614), .Z(N245) );
  AND U6859 ( .A(out[234]), .B(n1614), .Z(N246) );
  AND U6860 ( .A(out[235]), .B(n1614), .Z(N247) );
  AND U6861 ( .A(out[236]), .B(n1614), .Z(N248) );
  AND U6862 ( .A(out[237]), .B(n1614), .Z(N249) );
  AND U6863 ( .A(out[13]), .B(n1614), .Z(N25) );
  AND U6864 ( .A(out[238]), .B(n1614), .Z(N250) );
  AND U6865 ( .A(out[239]), .B(n1614), .Z(N251) );
  AND U6866 ( .A(out[240]), .B(n1614), .Z(N252) );
  AND U6867 ( .A(out[241]), .B(n1614), .Z(N253) );
  AND U6868 ( .A(out[242]), .B(n1614), .Z(N254) );
  AND U6869 ( .A(out[243]), .B(n1614), .Z(N255) );
  AND U6870 ( .A(out[244]), .B(n1614), .Z(N256) );
  AND U6871 ( .A(out[245]), .B(n1614), .Z(N257) );
  AND U6872 ( .A(out[246]), .B(n1614), .Z(N258) );
  AND U6873 ( .A(out[247]), .B(n1614), .Z(N259) );
  AND U6874 ( .A(out[14]), .B(n1614), .Z(N26) );
  AND U6875 ( .A(out[248]), .B(n1614), .Z(N260) );
  AND U6876 ( .A(out[249]), .B(n1614), .Z(N261) );
  AND U6877 ( .A(out[250]), .B(n1614), .Z(N262) );
  AND U6878 ( .A(out[251]), .B(n1614), .Z(N263) );
  AND U6879 ( .A(out[252]), .B(n1614), .Z(N264) );
  AND U6880 ( .A(out[253]), .B(n1614), .Z(N265) );
  AND U6881 ( .A(out[254]), .B(n1614), .Z(N266) );
  AND U6882 ( .A(out[255]), .B(n1614), .Z(N267) );
  AND U6883 ( .A(out[256]), .B(n1614), .Z(N268) );
  AND U6884 ( .A(out[257]), .B(n1614), .Z(N269) );
  AND U6885 ( .A(out[15]), .B(n1614), .Z(N27) );
  AND U6886 ( .A(out[258]), .B(n1614), .Z(N270) );
  AND U6887 ( .A(out[259]), .B(n1614), .Z(N271) );
  AND U6888 ( .A(out[260]), .B(n1614), .Z(N272) );
  AND U6889 ( .A(out[261]), .B(n1614), .Z(N273) );
  AND U6890 ( .A(out[262]), .B(n1614), .Z(N274) );
  AND U6891 ( .A(out[263]), .B(n1614), .Z(N275) );
  AND U6892 ( .A(out[264]), .B(n1614), .Z(N276) );
  AND U6893 ( .A(out[265]), .B(n1614), .Z(N277) );
  AND U6894 ( .A(out[266]), .B(n1614), .Z(N278) );
  AND U6895 ( .A(out[267]), .B(n1614), .Z(N279) );
  AND U6896 ( .A(out[16]), .B(n1614), .Z(N28) );
  AND U6897 ( .A(out[268]), .B(n1614), .Z(N280) );
  AND U6898 ( .A(out[269]), .B(n1614), .Z(N281) );
  AND U6899 ( .A(out[270]), .B(n1614), .Z(N282) );
  AND U6900 ( .A(out[271]), .B(n1614), .Z(N283) );
  AND U6901 ( .A(out[272]), .B(n1614), .Z(N284) );
  AND U6902 ( .A(out[273]), .B(n1614), .Z(N285) );
  AND U6903 ( .A(out[274]), .B(n1614), .Z(N286) );
  AND U6904 ( .A(out[275]), .B(n1614), .Z(N287) );
  AND U6905 ( .A(out[276]), .B(n1614), .Z(N288) );
  AND U6906 ( .A(out[277]), .B(n1614), .Z(N289) );
  AND U6907 ( .A(out[17]), .B(n1614), .Z(N29) );
  AND U6908 ( .A(out[278]), .B(n1614), .Z(N290) );
  AND U6909 ( .A(out[279]), .B(n1614), .Z(N291) );
  AND U6910 ( .A(out[280]), .B(n1614), .Z(N292) );
  AND U6911 ( .A(out[281]), .B(n1614), .Z(N293) );
  AND U6912 ( .A(out[282]), .B(n1614), .Z(N294) );
  AND U6913 ( .A(out[283]), .B(n1614), .Z(N295) );
  AND U6914 ( .A(out[284]), .B(n1614), .Z(N296) );
  AND U6915 ( .A(out[285]), .B(n1614), .Z(N297) );
  AND U6916 ( .A(out[286]), .B(n1614), .Z(N298) );
  AND U6917 ( .A(out[287]), .B(n1614), .Z(N299) );
  AND U6918 ( .A(out[18]), .B(n1614), .Z(N30) );
  AND U6919 ( .A(out[288]), .B(n1614), .Z(N300) );
  AND U6920 ( .A(out[289]), .B(n1614), .Z(N301) );
  AND U6921 ( .A(out[290]), .B(n1614), .Z(N302) );
  AND U6922 ( .A(out[291]), .B(n1614), .Z(N303) );
  AND U6923 ( .A(out[292]), .B(n1614), .Z(N304) );
  AND U6924 ( .A(out[293]), .B(n1614), .Z(N305) );
  AND U6925 ( .A(out[294]), .B(n1614), .Z(N306) );
  AND U6926 ( .A(out[295]), .B(n1614), .Z(N307) );
  AND U6927 ( .A(out[296]), .B(n1614), .Z(N308) );
  AND U6928 ( .A(out[297]), .B(n1614), .Z(N309) );
  AND U6929 ( .A(out[19]), .B(n1614), .Z(N31) );
  AND U6930 ( .A(out[298]), .B(n1614), .Z(N310) );
  AND U6931 ( .A(out[299]), .B(n1614), .Z(N311) );
  AND U6932 ( .A(out[300]), .B(n1614), .Z(N312) );
  AND U6933 ( .A(out[301]), .B(n1614), .Z(N313) );
  AND U6934 ( .A(out[302]), .B(n1614), .Z(N314) );
  AND U6935 ( .A(out[303]), .B(n1614), .Z(N315) );
  AND U6936 ( .A(out[304]), .B(n1614), .Z(N316) );
  AND U6937 ( .A(out[305]), .B(n1614), .Z(N317) );
  AND U6938 ( .A(out[306]), .B(n1614), .Z(N318) );
  AND U6939 ( .A(out[307]), .B(n1614), .Z(N319) );
  AND U6940 ( .A(out[20]), .B(n1614), .Z(N32) );
  AND U6941 ( .A(out[308]), .B(n1614), .Z(N320) );
  AND U6942 ( .A(out[309]), .B(n1614), .Z(N321) );
  AND U6943 ( .A(out[310]), .B(n1614), .Z(N322) );
  AND U6944 ( .A(out[311]), .B(n1614), .Z(N323) );
  AND U6945 ( .A(out[312]), .B(n1614), .Z(N324) );
  AND U6946 ( .A(out[313]), .B(n1614), .Z(N325) );
  AND U6947 ( .A(out[314]), .B(n1614), .Z(N326) );
  AND U6948 ( .A(out[315]), .B(n1614), .Z(N327) );
  AND U6949 ( .A(out[316]), .B(n1614), .Z(N328) );
  AND U6950 ( .A(out[317]), .B(n1614), .Z(N329) );
  AND U6951 ( .A(out[21]), .B(n1614), .Z(N33) );
  AND U6952 ( .A(out[318]), .B(n1614), .Z(N330) );
  AND U6953 ( .A(out[319]), .B(n1614), .Z(N331) );
  AND U6954 ( .A(out[320]), .B(n1614), .Z(N332) );
  AND U6955 ( .A(out[321]), .B(n1614), .Z(N333) );
  AND U6956 ( .A(out[322]), .B(n1614), .Z(N334) );
  AND U6957 ( .A(out[323]), .B(n1614), .Z(N335) );
  AND U6958 ( .A(out[324]), .B(n1614), .Z(N336) );
  AND U6959 ( .A(out[325]), .B(n1614), .Z(N337) );
  AND U6960 ( .A(out[326]), .B(n1614), .Z(N338) );
  AND U6961 ( .A(out[327]), .B(n1614), .Z(N339) );
  AND U6962 ( .A(out[22]), .B(n1614), .Z(N34) );
  AND U6963 ( .A(out[328]), .B(n1614), .Z(N340) );
  AND U6964 ( .A(out[329]), .B(n1614), .Z(N341) );
  AND U6965 ( .A(out[330]), .B(n1614), .Z(N342) );
  AND U6966 ( .A(out[331]), .B(n1614), .Z(N343) );
  AND U6967 ( .A(out[332]), .B(n1614), .Z(N344) );
  AND U6968 ( .A(out[333]), .B(n1614), .Z(N345) );
  AND U6969 ( .A(out[334]), .B(n1614), .Z(N346) );
  AND U6970 ( .A(out[335]), .B(n1614), .Z(N347) );
  AND U6971 ( .A(out[336]), .B(n1614), .Z(N348) );
  AND U6972 ( .A(out[337]), .B(n1614), .Z(N349) );
  AND U6973 ( .A(out[23]), .B(n1614), .Z(N35) );
  AND U6974 ( .A(out[338]), .B(n1614), .Z(N350) );
  AND U6975 ( .A(out[339]), .B(n1614), .Z(N351) );
  AND U6976 ( .A(out[340]), .B(n1614), .Z(N352) );
  AND U6977 ( .A(out[341]), .B(n1614), .Z(N353) );
  AND U6978 ( .A(out[342]), .B(n1614), .Z(N354) );
  AND U6979 ( .A(out[343]), .B(n1614), .Z(N355) );
  AND U6980 ( .A(out[344]), .B(n1614), .Z(N356) );
  AND U6981 ( .A(out[345]), .B(n1614), .Z(N357) );
  AND U6982 ( .A(out[346]), .B(n1614), .Z(N358) );
  AND U6983 ( .A(out[347]), .B(n1614), .Z(N359) );
  AND U6984 ( .A(out[24]), .B(n1614), .Z(N36) );
  AND U6985 ( .A(out[348]), .B(n1614), .Z(N360) );
  AND U6986 ( .A(out[349]), .B(n1614), .Z(N361) );
  AND U6987 ( .A(out[350]), .B(n1614), .Z(N362) );
  AND U6988 ( .A(out[351]), .B(n1614), .Z(N363) );
  AND U6989 ( .A(out[352]), .B(n1614), .Z(N364) );
  AND U6990 ( .A(out[353]), .B(n1614), .Z(N365) );
  AND U6991 ( .A(out[354]), .B(n1614), .Z(N366) );
  AND U6992 ( .A(out[355]), .B(n1614), .Z(N367) );
  AND U6993 ( .A(out[356]), .B(n1614), .Z(N368) );
  AND U6994 ( .A(out[357]), .B(n1614), .Z(N369) );
  AND U6995 ( .A(out[25]), .B(n1614), .Z(N37) );
  AND U6996 ( .A(out[358]), .B(n1614), .Z(N370) );
  AND U6997 ( .A(out[359]), .B(n1614), .Z(N371) );
  AND U6998 ( .A(out[360]), .B(n1614), .Z(N372) );
  AND U6999 ( .A(out[361]), .B(n1614), .Z(N373) );
  AND U7000 ( .A(out[362]), .B(n1614), .Z(N374) );
  AND U7001 ( .A(out[363]), .B(n1614), .Z(N375) );
  AND U7002 ( .A(out[364]), .B(n1614), .Z(N376) );
  AND U7003 ( .A(out[365]), .B(n1614), .Z(N377) );
  AND U7004 ( .A(out[366]), .B(n1614), .Z(N378) );
  AND U7005 ( .A(out[367]), .B(n1614), .Z(N379) );
  AND U7006 ( .A(out[26]), .B(n1614), .Z(N38) );
  AND U7007 ( .A(out[368]), .B(n1614), .Z(N380) );
  AND U7008 ( .A(out[369]), .B(n1614), .Z(N381) );
  AND U7009 ( .A(out[370]), .B(n1614), .Z(N382) );
  AND U7010 ( .A(out[371]), .B(n1614), .Z(N383) );
  AND U7011 ( .A(out[372]), .B(n1614), .Z(N384) );
  AND U7012 ( .A(out[373]), .B(n1614), .Z(N385) );
  AND U7013 ( .A(out[374]), .B(n1614), .Z(N386) );
  AND U7014 ( .A(out[375]), .B(n1614), .Z(N387) );
  AND U7015 ( .A(out[376]), .B(n1614), .Z(N388) );
  AND U7016 ( .A(out[377]), .B(n1614), .Z(N389) );
  AND U7017 ( .A(out[27]), .B(n1614), .Z(N39) );
  AND U7018 ( .A(out[378]), .B(n1614), .Z(N390) );
  AND U7019 ( .A(out[379]), .B(n1614), .Z(N391) );
  AND U7020 ( .A(out[380]), .B(n1614), .Z(N392) );
  AND U7021 ( .A(out[381]), .B(n1614), .Z(N393) );
  AND U7022 ( .A(out[382]), .B(n1614), .Z(N394) );
  AND U7023 ( .A(out[383]), .B(n1614), .Z(N395) );
  AND U7024 ( .A(out[384]), .B(n1614), .Z(N396) );
  AND U7025 ( .A(out[385]), .B(n1614), .Z(N397) );
  AND U7026 ( .A(out[386]), .B(n1614), .Z(N398) );
  AND U7027 ( .A(out[387]), .B(n1614), .Z(N399) );
  AND U7028 ( .A(out[28]), .B(n1614), .Z(N40) );
  AND U7029 ( .A(out[388]), .B(n1614), .Z(N400) );
  AND U7030 ( .A(out[389]), .B(n1614), .Z(N401) );
  AND U7031 ( .A(out[390]), .B(n1614), .Z(N402) );
  AND U7032 ( .A(out[391]), .B(n1614), .Z(N403) );
  AND U7033 ( .A(out[392]), .B(n1614), .Z(N404) );
  AND U7034 ( .A(out[393]), .B(n1614), .Z(N405) );
  AND U7035 ( .A(out[394]), .B(n1614), .Z(N406) );
  AND U7036 ( .A(out[395]), .B(n1614), .Z(N407) );
  AND U7037 ( .A(out[396]), .B(n1614), .Z(N408) );
  AND U7038 ( .A(out[397]), .B(n1614), .Z(N409) );
  AND U7039 ( .A(out[29]), .B(n1614), .Z(N41) );
  AND U7040 ( .A(out[398]), .B(n1614), .Z(N410) );
  AND U7041 ( .A(out[399]), .B(n1614), .Z(N411) );
  AND U7042 ( .A(out[400]), .B(n1614), .Z(N412) );
  AND U7043 ( .A(out[401]), .B(n1614), .Z(N413) );
  AND U7044 ( .A(out[402]), .B(n1614), .Z(N414) );
  AND U7045 ( .A(out[403]), .B(n1614), .Z(N415) );
  AND U7046 ( .A(out[404]), .B(n1614), .Z(N416) );
  AND U7047 ( .A(out[405]), .B(n1614), .Z(N417) );
  AND U7048 ( .A(out[406]), .B(n1614), .Z(N418) );
  AND U7049 ( .A(out[407]), .B(n1614), .Z(N419) );
  AND U7050 ( .A(out[30]), .B(n1614), .Z(N42) );
  AND U7051 ( .A(out[408]), .B(n1614), .Z(N420) );
  AND U7052 ( .A(out[409]), .B(n1614), .Z(N421) );
  AND U7053 ( .A(out[410]), .B(n1614), .Z(N422) );
  AND U7054 ( .A(out[411]), .B(n1614), .Z(N423) );
  AND U7055 ( .A(out[412]), .B(n1614), .Z(N424) );
  AND U7056 ( .A(out[413]), .B(n1614), .Z(N425) );
  AND U7057 ( .A(out[414]), .B(n1614), .Z(N426) );
  AND U7058 ( .A(out[415]), .B(n1614), .Z(N427) );
  AND U7059 ( .A(out[416]), .B(n1614), .Z(N428) );
  AND U7060 ( .A(out[417]), .B(n1614), .Z(N429) );
  AND U7061 ( .A(out[31]), .B(n1614), .Z(N43) );
  AND U7062 ( .A(out[418]), .B(n1614), .Z(N430) );
  AND U7063 ( .A(out[419]), .B(n1614), .Z(N431) );
  AND U7064 ( .A(out[420]), .B(n1614), .Z(N432) );
  AND U7065 ( .A(out[421]), .B(n1614), .Z(N433) );
  AND U7066 ( .A(out[422]), .B(n1614), .Z(N434) );
  AND U7067 ( .A(out[423]), .B(n1614), .Z(N435) );
  AND U7068 ( .A(out[424]), .B(n1614), .Z(N436) );
  AND U7069 ( .A(out[425]), .B(n1614), .Z(N437) );
  AND U7070 ( .A(out[426]), .B(n1614), .Z(N438) );
  AND U7071 ( .A(out[427]), .B(n1614), .Z(N439) );
  AND U7072 ( .A(out[32]), .B(n1614), .Z(N44) );
  AND U7073 ( .A(out[428]), .B(n1614), .Z(N440) );
  AND U7074 ( .A(out[429]), .B(n1614), .Z(N441) );
  AND U7075 ( .A(out[430]), .B(n1614), .Z(N442) );
  AND U7076 ( .A(out[431]), .B(n1614), .Z(N443) );
  AND U7077 ( .A(out[432]), .B(n1614), .Z(N444) );
  AND U7078 ( .A(out[433]), .B(n1614), .Z(N445) );
  AND U7079 ( .A(out[434]), .B(n1614), .Z(N446) );
  AND U7080 ( .A(out[435]), .B(n1614), .Z(N447) );
  AND U7081 ( .A(out[436]), .B(n1614), .Z(N448) );
  AND U7082 ( .A(out[437]), .B(n1614), .Z(N449) );
  AND U7083 ( .A(out[33]), .B(n1614), .Z(N45) );
  AND U7084 ( .A(out[438]), .B(n1614), .Z(N450) );
  AND U7085 ( .A(out[439]), .B(n1614), .Z(N451) );
  AND U7086 ( .A(out[440]), .B(n1614), .Z(N452) );
  AND U7087 ( .A(out[441]), .B(n1614), .Z(N453) );
  AND U7088 ( .A(out[442]), .B(n1614), .Z(N454) );
  AND U7089 ( .A(out[443]), .B(n1614), .Z(N455) );
  AND U7090 ( .A(out[444]), .B(n1614), .Z(N456) );
  AND U7091 ( .A(out[445]), .B(n1614), .Z(N457) );
  AND U7092 ( .A(out[446]), .B(n1614), .Z(N458) );
  AND U7093 ( .A(out[447]), .B(n1614), .Z(N459) );
  AND U7094 ( .A(out[34]), .B(n1614), .Z(N46) );
  AND U7095 ( .A(out[448]), .B(n1614), .Z(N460) );
  AND U7096 ( .A(out[449]), .B(n1614), .Z(N461) );
  AND U7097 ( .A(out[450]), .B(n1614), .Z(N462) );
  AND U7098 ( .A(out[451]), .B(n1614), .Z(N463) );
  AND U7099 ( .A(out[452]), .B(n1614), .Z(N464) );
  AND U7100 ( .A(out[453]), .B(n1614), .Z(N465) );
  AND U7101 ( .A(out[454]), .B(n1614), .Z(N466) );
  AND U7102 ( .A(out[455]), .B(n1614), .Z(N467) );
  AND U7103 ( .A(out[456]), .B(n1614), .Z(N468) );
  AND U7104 ( .A(out[457]), .B(n1614), .Z(N469) );
  AND U7105 ( .A(out[35]), .B(n1614), .Z(N47) );
  AND U7106 ( .A(out[458]), .B(n1614), .Z(N470) );
  AND U7107 ( .A(out[459]), .B(n1614), .Z(N471) );
  AND U7108 ( .A(out[460]), .B(n1614), .Z(N472) );
  AND U7109 ( .A(out[461]), .B(n1614), .Z(N473) );
  AND U7110 ( .A(out[462]), .B(n1614), .Z(N474) );
  AND U7111 ( .A(out[463]), .B(n1614), .Z(N475) );
  AND U7112 ( .A(out[464]), .B(n1614), .Z(N476) );
  AND U7113 ( .A(out[465]), .B(n1614), .Z(N477) );
  AND U7114 ( .A(out[466]), .B(n1614), .Z(N478) );
  AND U7115 ( .A(out[467]), .B(n1614), .Z(N479) );
  AND U7116 ( .A(out[36]), .B(n1614), .Z(N48) );
  AND U7117 ( .A(out[468]), .B(n1614), .Z(N480) );
  AND U7118 ( .A(out[469]), .B(n1614), .Z(N481) );
  AND U7119 ( .A(out[470]), .B(n1614), .Z(N482) );
  AND U7120 ( .A(out[471]), .B(n1614), .Z(N483) );
  AND U7121 ( .A(out[472]), .B(n1614), .Z(N484) );
  AND U7122 ( .A(out[473]), .B(n1614), .Z(N485) );
  AND U7123 ( .A(out[474]), .B(n1614), .Z(N486) );
  AND U7124 ( .A(out[475]), .B(n1614), .Z(N487) );
  AND U7125 ( .A(out[476]), .B(n1614), .Z(N488) );
  AND U7126 ( .A(out[477]), .B(n1614), .Z(N489) );
  AND U7127 ( .A(out[37]), .B(n1614), .Z(N49) );
  AND U7128 ( .A(out[478]), .B(n1614), .Z(N490) );
  AND U7129 ( .A(out[479]), .B(n1614), .Z(N491) );
  AND U7130 ( .A(out[480]), .B(n1614), .Z(N492) );
  AND U7131 ( .A(out[481]), .B(n1614), .Z(N493) );
  AND U7132 ( .A(out[482]), .B(n1614), .Z(N494) );
  AND U7133 ( .A(out[483]), .B(n1614), .Z(N495) );
  AND U7134 ( .A(out[484]), .B(n1614), .Z(N496) );
  AND U7135 ( .A(out[485]), .B(n1614), .Z(N497) );
  AND U7136 ( .A(out[486]), .B(n1614), .Z(N498) );
  AND U7137 ( .A(out[487]), .B(n1614), .Z(N499) );
  AND U7138 ( .A(out[38]), .B(n1614), .Z(N50) );
  AND U7139 ( .A(out[488]), .B(n1614), .Z(N500) );
  AND U7140 ( .A(out[489]), .B(n1614), .Z(N501) );
  AND U7141 ( .A(out[490]), .B(n1614), .Z(N502) );
  AND U7142 ( .A(out[491]), .B(n1614), .Z(N503) );
  AND U7143 ( .A(out[492]), .B(n1614), .Z(N504) );
  AND U7144 ( .A(out[493]), .B(n1614), .Z(N505) );
  AND U7145 ( .A(out[494]), .B(n1614), .Z(N506) );
  AND U7146 ( .A(out[495]), .B(n1614), .Z(N507) );
  AND U7147 ( .A(out[496]), .B(n1614), .Z(N508) );
  AND U7148 ( .A(out[497]), .B(n1614), .Z(N509) );
  AND U7149 ( .A(out[39]), .B(n1614), .Z(N51) );
  AND U7150 ( .A(out[498]), .B(n1614), .Z(N510) );
  AND U7151 ( .A(out[499]), .B(n1614), .Z(N511) );
  AND U7152 ( .A(out[500]), .B(n1614), .Z(N512) );
  AND U7153 ( .A(out[501]), .B(n1614), .Z(N513) );
  AND U7154 ( .A(out[502]), .B(n1614), .Z(N514) );
  AND U7155 ( .A(out[503]), .B(n1614), .Z(N515) );
  AND U7156 ( .A(out[504]), .B(n1614), .Z(N516) );
  AND U7157 ( .A(out[505]), .B(n1614), .Z(N517) );
  AND U7158 ( .A(out[506]), .B(n1614), .Z(N518) );
  AND U7159 ( .A(out[507]), .B(n1614), .Z(N519) );
  AND U7160 ( .A(out[40]), .B(n1614), .Z(N52) );
  AND U7161 ( .A(out[508]), .B(n1614), .Z(N520) );
  AND U7162 ( .A(out[509]), .B(n1614), .Z(N521) );
  AND U7163 ( .A(out[510]), .B(n1614), .Z(N522) );
  AND U7164 ( .A(out[511]), .B(n1614), .Z(N523) );
  AND U7165 ( .A(out[512]), .B(n1614), .Z(N524) );
  AND U7166 ( .A(out[513]), .B(n1614), .Z(N525) );
  AND U7167 ( .A(out[514]), .B(n1614), .Z(N526) );
  AND U7168 ( .A(out[515]), .B(n1614), .Z(N527) );
  AND U7169 ( .A(out[516]), .B(n1614), .Z(N528) );
  AND U7170 ( .A(out[517]), .B(n1614), .Z(N529) );
  AND U7171 ( .A(out[41]), .B(n1614), .Z(N53) );
  AND U7172 ( .A(out[518]), .B(n1614), .Z(N530) );
  AND U7173 ( .A(out[519]), .B(n1614), .Z(N531) );
  AND U7174 ( .A(out[520]), .B(n1614), .Z(N532) );
  AND U7175 ( .A(out[521]), .B(n1614), .Z(N533) );
  AND U7176 ( .A(out[522]), .B(n1614), .Z(N534) );
  AND U7177 ( .A(out[523]), .B(n1614), .Z(N535) );
  AND U7178 ( .A(out[524]), .B(n1614), .Z(N536) );
  AND U7179 ( .A(out[525]), .B(n1614), .Z(N537) );
  AND U7180 ( .A(out[526]), .B(n1614), .Z(N538) );
  AND U7181 ( .A(out[527]), .B(n1614), .Z(N539) );
  AND U7182 ( .A(out[42]), .B(n1614), .Z(N54) );
  AND U7183 ( .A(out[528]), .B(n1614), .Z(N540) );
  AND U7184 ( .A(out[529]), .B(n1614), .Z(N541) );
  AND U7185 ( .A(out[530]), .B(n1614), .Z(N542) );
  AND U7186 ( .A(out[531]), .B(n1614), .Z(N543) );
  AND U7187 ( .A(out[532]), .B(n1614), .Z(N544) );
  AND U7188 ( .A(out[533]), .B(n1614), .Z(N545) );
  AND U7189 ( .A(out[534]), .B(n1614), .Z(N546) );
  AND U7190 ( .A(out[535]), .B(n1614), .Z(N547) );
  AND U7191 ( .A(out[536]), .B(n1614), .Z(N548) );
  AND U7192 ( .A(out[537]), .B(n1614), .Z(N549) );
  AND U7193 ( .A(out[43]), .B(n1614), .Z(N55) );
  AND U7194 ( .A(out[538]), .B(n1614), .Z(N550) );
  AND U7195 ( .A(out[539]), .B(n1614), .Z(N551) );
  AND U7196 ( .A(out[540]), .B(n1614), .Z(N552) );
  AND U7197 ( .A(out[541]), .B(n1614), .Z(N553) );
  AND U7198 ( .A(out[542]), .B(n1614), .Z(N554) );
  AND U7199 ( .A(out[543]), .B(n1614), .Z(N555) );
  AND U7200 ( .A(out[544]), .B(n1614), .Z(N556) );
  AND U7201 ( .A(out[545]), .B(n1614), .Z(N557) );
  AND U7202 ( .A(out[546]), .B(n1614), .Z(N558) );
  AND U7203 ( .A(out[547]), .B(n1614), .Z(N559) );
  AND U7204 ( .A(out[44]), .B(n1614), .Z(N56) );
  AND U7205 ( .A(out[548]), .B(n1614), .Z(N560) );
  AND U7206 ( .A(out[549]), .B(n1614), .Z(N561) );
  AND U7207 ( .A(out[550]), .B(n1614), .Z(N562) );
  AND U7208 ( .A(out[551]), .B(n1614), .Z(N563) );
  AND U7209 ( .A(out[552]), .B(n1614), .Z(N564) );
  AND U7210 ( .A(out[553]), .B(n1614), .Z(N565) );
  AND U7211 ( .A(out[554]), .B(n1614), .Z(N566) );
  AND U7212 ( .A(out[555]), .B(n1614), .Z(N567) );
  AND U7213 ( .A(out[556]), .B(n1614), .Z(N568) );
  AND U7214 ( .A(out[557]), .B(n1614), .Z(N569) );
  AND U7215 ( .A(out[45]), .B(n1614), .Z(N57) );
  AND U7216 ( .A(out[558]), .B(n1614), .Z(N570) );
  AND U7217 ( .A(out[559]), .B(n1614), .Z(N571) );
  AND U7218 ( .A(out[560]), .B(n1614), .Z(N572) );
  AND U7219 ( .A(out[561]), .B(n1614), .Z(N573) );
  AND U7220 ( .A(out[562]), .B(n1614), .Z(N574) );
  AND U7221 ( .A(out[563]), .B(n1614), .Z(N575) );
  AND U7222 ( .A(out[564]), .B(n1614), .Z(N576) );
  AND U7223 ( .A(out[565]), .B(n1614), .Z(N577) );
  AND U7224 ( .A(out[566]), .B(n1614), .Z(N578) );
  AND U7225 ( .A(out[567]), .B(n1614), .Z(N579) );
  AND U7226 ( .A(out[46]), .B(n1614), .Z(N58) );
  AND U7227 ( .A(out[568]), .B(n1614), .Z(N580) );
  AND U7228 ( .A(out[569]), .B(n1614), .Z(N581) );
  AND U7229 ( .A(out[570]), .B(n1614), .Z(N582) );
  AND U7230 ( .A(out[571]), .B(n1614), .Z(N583) );
  AND U7231 ( .A(out[572]), .B(n1614), .Z(N584) );
  AND U7232 ( .A(out[573]), .B(n1614), .Z(N585) );
  AND U7233 ( .A(out[574]), .B(n1614), .Z(N586) );
  AND U7234 ( .A(out[575]), .B(n1614), .Z(N587) );
  AND U7235 ( .A(out[576]), .B(n1614), .Z(N588) );
  AND U7236 ( .A(out[577]), .B(n1614), .Z(N589) );
  AND U7237 ( .A(out[47]), .B(n1614), .Z(N59) );
  AND U7238 ( .A(out[578]), .B(n1614), .Z(N590) );
  AND U7239 ( .A(out[579]), .B(n1614), .Z(N591) );
  AND U7240 ( .A(out[580]), .B(n1614), .Z(N592) );
  AND U7241 ( .A(out[581]), .B(n1614), .Z(N593) );
  AND U7242 ( .A(out[582]), .B(n1614), .Z(N594) );
  AND U7243 ( .A(out[583]), .B(n1614), .Z(N595) );
  AND U7244 ( .A(out[584]), .B(n1614), .Z(N596) );
  AND U7245 ( .A(out[585]), .B(n1614), .Z(N597) );
  AND U7246 ( .A(out[586]), .B(n1614), .Z(N598) );
  AND U7247 ( .A(out[587]), .B(n1614), .Z(N599) );
  AND U7248 ( .A(n1614), .B(n2770), .Z(N6) );
  AND U7249 ( .A(out[48]), .B(n1614), .Z(N60) );
  AND U7250 ( .A(out[588]), .B(n1614), .Z(N600) );
  AND U7251 ( .A(out[589]), .B(n1614), .Z(N601) );
  AND U7252 ( .A(out[590]), .B(n1614), .Z(N602) );
  AND U7253 ( .A(out[591]), .B(n1614), .Z(N603) );
  AND U7254 ( .A(out[592]), .B(n1614), .Z(N604) );
  AND U7255 ( .A(out[593]), .B(n1614), .Z(N605) );
  AND U7256 ( .A(out[594]), .B(n1614), .Z(N606) );
  AND U7257 ( .A(out[595]), .B(n1614), .Z(N607) );
  AND U7258 ( .A(out[596]), .B(n1614), .Z(N608) );
  AND U7259 ( .A(out[597]), .B(n1614), .Z(N609) );
  AND U7260 ( .A(out[49]), .B(n1614), .Z(N61) );
  AND U7261 ( .A(out[598]), .B(n1614), .Z(N610) );
  AND U7262 ( .A(out[599]), .B(n1614), .Z(N611) );
  AND U7263 ( .A(out[600]), .B(n1614), .Z(N612) );
  AND U7264 ( .A(out[601]), .B(n1614), .Z(N613) );
  AND U7265 ( .A(out[602]), .B(n1614), .Z(N614) );
  AND U7266 ( .A(out[603]), .B(n1614), .Z(N615) );
  AND U7267 ( .A(out[604]), .B(n1614), .Z(N616) );
  AND U7268 ( .A(out[605]), .B(n1614), .Z(N617) );
  AND U7269 ( .A(out[606]), .B(n1614), .Z(N618) );
  AND U7270 ( .A(out[607]), .B(n1614), .Z(N619) );
  AND U7271 ( .A(out[50]), .B(n1614), .Z(N62) );
  AND U7272 ( .A(out[608]), .B(n1614), .Z(N620) );
  AND U7273 ( .A(out[609]), .B(n1614), .Z(N621) );
  AND U7274 ( .A(out[610]), .B(n1614), .Z(N622) );
  AND U7275 ( .A(out[611]), .B(n1614), .Z(N623) );
  AND U7276 ( .A(out[612]), .B(n1614), .Z(N624) );
  AND U7277 ( .A(out[613]), .B(n1614), .Z(N625) );
  AND U7278 ( .A(out[614]), .B(n1614), .Z(N626) );
  AND U7279 ( .A(out[615]), .B(n1614), .Z(N627) );
  AND U7280 ( .A(out[616]), .B(n1614), .Z(N628) );
  AND U7281 ( .A(out[617]), .B(n1614), .Z(N629) );
  AND U7282 ( .A(out[51]), .B(n1614), .Z(N63) );
  AND U7283 ( .A(out[618]), .B(n1614), .Z(N630) );
  AND U7284 ( .A(out[619]), .B(n1614), .Z(N631) );
  AND U7285 ( .A(out[620]), .B(n1614), .Z(N632) );
  AND U7286 ( .A(out[621]), .B(n1614), .Z(N633) );
  AND U7287 ( .A(out[622]), .B(n1614), .Z(N634) );
  AND U7288 ( .A(out[623]), .B(n1614), .Z(N635) );
  AND U7289 ( .A(out[624]), .B(n1614), .Z(N636) );
  AND U7290 ( .A(out[625]), .B(n1614), .Z(N637) );
  AND U7291 ( .A(out[626]), .B(n1614), .Z(N638) );
  AND U7292 ( .A(out[627]), .B(n1614), .Z(N639) );
  AND U7293 ( .A(out[52]), .B(n1614), .Z(N64) );
  AND U7294 ( .A(out[628]), .B(n1614), .Z(N640) );
  AND U7295 ( .A(out[629]), .B(n1614), .Z(N641) );
  AND U7296 ( .A(out[630]), .B(n1614), .Z(N642) );
  AND U7297 ( .A(out[631]), .B(n1614), .Z(N643) );
  AND U7298 ( .A(out[632]), .B(n1614), .Z(N644) );
  AND U7299 ( .A(out[633]), .B(n1614), .Z(N645) );
  AND U7300 ( .A(out[634]), .B(n1614), .Z(N646) );
  AND U7301 ( .A(out[635]), .B(n1614), .Z(N647) );
  AND U7302 ( .A(out[636]), .B(n1614), .Z(N648) );
  AND U7303 ( .A(out[637]), .B(n1614), .Z(N649) );
  AND U7304 ( .A(out[53]), .B(n1614), .Z(N65) );
  AND U7305 ( .A(out[638]), .B(n1614), .Z(N650) );
  AND U7306 ( .A(out[639]), .B(n1614), .Z(N651) );
  AND U7307 ( .A(out[640]), .B(n1614), .Z(N652) );
  AND U7308 ( .A(out[641]), .B(n1614), .Z(N653) );
  AND U7309 ( .A(out[642]), .B(n1614), .Z(N654) );
  AND U7310 ( .A(out[643]), .B(n1614), .Z(N655) );
  AND U7311 ( .A(out[644]), .B(n1614), .Z(N656) );
  AND U7312 ( .A(out[645]), .B(n1614), .Z(N657) );
  AND U7313 ( .A(out[646]), .B(n1614), .Z(N658) );
  AND U7314 ( .A(out[647]), .B(n1614), .Z(N659) );
  AND U7315 ( .A(out[54]), .B(n1614), .Z(N66) );
  AND U7316 ( .A(out[648]), .B(n1614), .Z(N660) );
  AND U7317 ( .A(out[649]), .B(n1614), .Z(N661) );
  AND U7318 ( .A(out[650]), .B(n1614), .Z(N662) );
  AND U7319 ( .A(out[651]), .B(n1614), .Z(N663) );
  AND U7320 ( .A(out[652]), .B(n1614), .Z(N664) );
  AND U7321 ( .A(out[653]), .B(n1614), .Z(N665) );
  AND U7322 ( .A(out[654]), .B(n1614), .Z(N666) );
  AND U7323 ( .A(out[655]), .B(n1614), .Z(N667) );
  AND U7324 ( .A(out[656]), .B(n1614), .Z(N668) );
  AND U7325 ( .A(out[657]), .B(n1614), .Z(N669) );
  AND U7326 ( .A(out[55]), .B(n1614), .Z(N67) );
  AND U7327 ( .A(out[658]), .B(n1614), .Z(N670) );
  AND U7328 ( .A(out[659]), .B(n1614), .Z(N671) );
  AND U7329 ( .A(out[660]), .B(n1614), .Z(N672) );
  AND U7330 ( .A(out[661]), .B(n1614), .Z(N673) );
  AND U7331 ( .A(out[662]), .B(n1614), .Z(N674) );
  AND U7332 ( .A(out[663]), .B(n1614), .Z(N675) );
  AND U7333 ( .A(out[664]), .B(n1614), .Z(N676) );
  AND U7334 ( .A(out[665]), .B(n1614), .Z(N677) );
  AND U7335 ( .A(out[666]), .B(n1614), .Z(N678) );
  AND U7336 ( .A(out[667]), .B(n1614), .Z(N679) );
  AND U7337 ( .A(out[56]), .B(n1614), .Z(N68) );
  AND U7338 ( .A(out[668]), .B(n1614), .Z(N680) );
  AND U7339 ( .A(out[669]), .B(n1614), .Z(N681) );
  AND U7340 ( .A(out[670]), .B(n1614), .Z(N682) );
  AND U7341 ( .A(out[671]), .B(n1614), .Z(N683) );
  AND U7342 ( .A(out[672]), .B(n1614), .Z(N684) );
  AND U7343 ( .A(out[673]), .B(n1614), .Z(N685) );
  AND U7344 ( .A(out[674]), .B(n1614), .Z(N686) );
  AND U7345 ( .A(out[675]), .B(n1614), .Z(N687) );
  AND U7346 ( .A(out[676]), .B(n1614), .Z(N688) );
  AND U7347 ( .A(out[677]), .B(n1614), .Z(N689) );
  AND U7348 ( .A(out[57]), .B(n1614), .Z(N69) );
  AND U7349 ( .A(out[678]), .B(n1614), .Z(N690) );
  AND U7350 ( .A(out[679]), .B(n1614), .Z(N691) );
  AND U7351 ( .A(out[680]), .B(n1614), .Z(N692) );
  AND U7352 ( .A(out[681]), .B(n1614), .Z(N693) );
  AND U7353 ( .A(out[682]), .B(n1614), .Z(N694) );
  AND U7354 ( .A(out[683]), .B(n1614), .Z(N695) );
  AND U7355 ( .A(out[684]), .B(n1614), .Z(N696) );
  AND U7356 ( .A(out[685]), .B(n1614), .Z(N697) );
  AND U7357 ( .A(out[686]), .B(n1614), .Z(N698) );
  AND U7358 ( .A(out[687]), .B(n1614), .Z(N699) );
  AND U7359 ( .A(n1614), .B(rc_i[0]), .Z(N7) );
  AND U7360 ( .A(out[58]), .B(n1614), .Z(N70) );
  AND U7361 ( .A(out[688]), .B(n1614), .Z(N700) );
  AND U7362 ( .A(out[689]), .B(n1614), .Z(N701) );
  AND U7363 ( .A(out[690]), .B(n1614), .Z(N702) );
  AND U7364 ( .A(out[691]), .B(n1614), .Z(N703) );
  AND U7365 ( .A(out[692]), .B(n1614), .Z(N704) );
  AND U7366 ( .A(out[693]), .B(n1614), .Z(N705) );
  AND U7367 ( .A(out[694]), .B(n1614), .Z(N706) );
  AND U7368 ( .A(out[695]), .B(n1614), .Z(N707) );
  AND U7369 ( .A(out[696]), .B(n1614), .Z(N708) );
  AND U7370 ( .A(out[697]), .B(n1614), .Z(N709) );
  AND U7371 ( .A(out[59]), .B(n1614), .Z(N71) );
  AND U7372 ( .A(out[698]), .B(n1614), .Z(N710) );
  AND U7373 ( .A(out[699]), .B(n1614), .Z(N711) );
  AND U7374 ( .A(out[700]), .B(n1614), .Z(N712) );
  AND U7375 ( .A(out[701]), .B(n1614), .Z(N713) );
  AND U7376 ( .A(out[702]), .B(n1614), .Z(N714) );
  AND U7377 ( .A(out[703]), .B(n1614), .Z(N715) );
  AND U7378 ( .A(out[704]), .B(n1614), .Z(N716) );
  AND U7379 ( .A(out[705]), .B(n1614), .Z(N717) );
  AND U7380 ( .A(out[706]), .B(n1614), .Z(N718) );
  AND U7381 ( .A(out[707]), .B(n1614), .Z(N719) );
  AND U7382 ( .A(out[60]), .B(n1614), .Z(N72) );
  AND U7383 ( .A(out[708]), .B(n1614), .Z(N720) );
  AND U7384 ( .A(out[709]), .B(n1614), .Z(N721) );
  AND U7385 ( .A(out[710]), .B(n1614), .Z(N722) );
  AND U7386 ( .A(out[711]), .B(n1614), .Z(N723) );
  AND U7387 ( .A(out[712]), .B(n1614), .Z(N724) );
  AND U7388 ( .A(out[713]), .B(n1614), .Z(N725) );
  AND U7389 ( .A(out[714]), .B(n1614), .Z(N726) );
  AND U7390 ( .A(out[715]), .B(n1614), .Z(N727) );
  AND U7391 ( .A(out[716]), .B(n1614), .Z(N728) );
  AND U7392 ( .A(out[717]), .B(n1614), .Z(N729) );
  AND U7393 ( .A(out[61]), .B(n1614), .Z(N73) );
  AND U7394 ( .A(out[718]), .B(n1614), .Z(N730) );
  AND U7395 ( .A(out[719]), .B(n1614), .Z(N731) );
  AND U7396 ( .A(out[720]), .B(n1614), .Z(N732) );
  AND U7397 ( .A(out[721]), .B(n1614), .Z(N733) );
  AND U7398 ( .A(out[722]), .B(n1614), .Z(N734) );
  AND U7399 ( .A(out[723]), .B(n1614), .Z(N735) );
  AND U7400 ( .A(out[724]), .B(n1614), .Z(N736) );
  AND U7401 ( .A(out[725]), .B(n1614), .Z(N737) );
  AND U7402 ( .A(out[726]), .B(n1614), .Z(N738) );
  AND U7403 ( .A(out[727]), .B(n1614), .Z(N739) );
  AND U7404 ( .A(out[62]), .B(n1614), .Z(N74) );
  AND U7405 ( .A(out[728]), .B(n1614), .Z(N740) );
  AND U7406 ( .A(out[729]), .B(n1614), .Z(N741) );
  AND U7407 ( .A(out[730]), .B(n1614), .Z(N742) );
  AND U7408 ( .A(out[731]), .B(n1614), .Z(N743) );
  AND U7409 ( .A(out[732]), .B(n1614), .Z(N744) );
  AND U7410 ( .A(out[733]), .B(n1614), .Z(N745) );
  AND U7411 ( .A(out[734]), .B(n1614), .Z(N746) );
  AND U7412 ( .A(out[735]), .B(n1614), .Z(N747) );
  AND U7413 ( .A(out[736]), .B(n1614), .Z(N748) );
  AND U7414 ( .A(out[737]), .B(n1614), .Z(N749) );
  AND U7415 ( .A(out[63]), .B(n1614), .Z(N75) );
  AND U7416 ( .A(out[738]), .B(n1614), .Z(N750) );
  AND U7417 ( .A(out[739]), .B(n1614), .Z(N751) );
  AND U7418 ( .A(out[740]), .B(n1614), .Z(N752) );
  AND U7419 ( .A(out[741]), .B(n1614), .Z(N753) );
  AND U7420 ( .A(out[742]), .B(n1614), .Z(N754) );
  AND U7421 ( .A(out[743]), .B(n1614), .Z(N755) );
  AND U7422 ( .A(out[744]), .B(n1614), .Z(N756) );
  AND U7423 ( .A(out[745]), .B(n1614), .Z(N757) );
  AND U7424 ( .A(out[746]), .B(n1614), .Z(N758) );
  AND U7425 ( .A(out[747]), .B(n1614), .Z(N759) );
  AND U7426 ( .A(out[64]), .B(n1614), .Z(N76) );
  AND U7427 ( .A(out[748]), .B(n1614), .Z(N760) );
  AND U7428 ( .A(out[749]), .B(n1614), .Z(N761) );
  AND U7429 ( .A(out[750]), .B(n1614), .Z(N762) );
  AND U7430 ( .A(out[751]), .B(n1614), .Z(N763) );
  AND U7431 ( .A(out[752]), .B(n1614), .Z(N764) );
  AND U7432 ( .A(out[753]), .B(n1614), .Z(N765) );
  AND U7433 ( .A(out[754]), .B(n1614), .Z(N766) );
  AND U7434 ( .A(out[755]), .B(n1614), .Z(N767) );
  AND U7435 ( .A(out[756]), .B(n1614), .Z(N768) );
  AND U7436 ( .A(out[757]), .B(n1614), .Z(N769) );
  AND U7437 ( .A(out[65]), .B(n1614), .Z(N77) );
  AND U7438 ( .A(out[758]), .B(n1614), .Z(N770) );
  AND U7439 ( .A(out[759]), .B(n1614), .Z(N771) );
  AND U7440 ( .A(out[760]), .B(n1614), .Z(N772) );
  AND U7441 ( .A(out[761]), .B(n1614), .Z(N773) );
  AND U7442 ( .A(out[762]), .B(n1614), .Z(N774) );
  AND U7443 ( .A(out[763]), .B(n1614), .Z(N775) );
  AND U7444 ( .A(out[764]), .B(n1614), .Z(N776) );
  AND U7445 ( .A(out[765]), .B(n1614), .Z(N777) );
  AND U7446 ( .A(out[766]), .B(n1614), .Z(N778) );
  AND U7447 ( .A(out[767]), .B(n1614), .Z(N779) );
  AND U7448 ( .A(out[66]), .B(n1614), .Z(N78) );
  AND U7449 ( .A(out[768]), .B(n1614), .Z(N780) );
  AND U7450 ( .A(out[769]), .B(n1614), .Z(N781) );
  AND U7451 ( .A(out[770]), .B(n1614), .Z(N782) );
  AND U7452 ( .A(out[771]), .B(n1614), .Z(N783) );
  AND U7453 ( .A(out[772]), .B(n1614), .Z(N784) );
  AND U7454 ( .A(out[773]), .B(n1614), .Z(N785) );
  AND U7455 ( .A(out[774]), .B(n1614), .Z(N786) );
  AND U7456 ( .A(out[775]), .B(n1614), .Z(N787) );
  AND U7457 ( .A(out[776]), .B(n1614), .Z(N788) );
  AND U7458 ( .A(out[777]), .B(n1614), .Z(N789) );
  AND U7459 ( .A(out[67]), .B(n1614), .Z(N79) );
  AND U7460 ( .A(out[778]), .B(n1614), .Z(N790) );
  AND U7461 ( .A(out[779]), .B(n1614), .Z(N791) );
  AND U7462 ( .A(out[780]), .B(n1614), .Z(N792) );
  AND U7463 ( .A(out[781]), .B(n1614), .Z(N793) );
  AND U7464 ( .A(out[782]), .B(n1614), .Z(N794) );
  AND U7465 ( .A(out[783]), .B(n1614), .Z(N795) );
  AND U7466 ( .A(out[784]), .B(n1614), .Z(N796) );
  AND U7467 ( .A(out[785]), .B(n1614), .Z(N797) );
  AND U7468 ( .A(out[786]), .B(n1614), .Z(N798) );
  AND U7469 ( .A(out[787]), .B(n1614), .Z(N799) );
  AND U7470 ( .A(rc_i[1]), .B(n1614), .Z(N8) );
  AND U7471 ( .A(out[68]), .B(n1614), .Z(N80) );
  AND U7472 ( .A(out[788]), .B(n1614), .Z(N800) );
  AND U7473 ( .A(out[789]), .B(n1614), .Z(N801) );
  AND U7474 ( .A(out[790]), .B(n1614), .Z(N802) );
  AND U7475 ( .A(out[791]), .B(n1614), .Z(N803) );
  AND U7476 ( .A(out[792]), .B(n1614), .Z(N804) );
  AND U7477 ( .A(out[793]), .B(n1614), .Z(N805) );
  AND U7478 ( .A(out[794]), .B(n1614), .Z(N806) );
  AND U7479 ( .A(out[795]), .B(n1614), .Z(N807) );
  AND U7480 ( .A(out[796]), .B(n1614), .Z(N808) );
  AND U7481 ( .A(out[797]), .B(n1614), .Z(N809) );
  AND U7482 ( .A(out[69]), .B(n1614), .Z(N81) );
  AND U7483 ( .A(out[798]), .B(n1614), .Z(N810) );
  AND U7484 ( .A(out[799]), .B(n1614), .Z(N811) );
  AND U7485 ( .A(out[800]), .B(n1614), .Z(N812) );
  AND U7486 ( .A(out[801]), .B(n1614), .Z(N813) );
  AND U7487 ( .A(out[802]), .B(n1614), .Z(N814) );
  AND U7488 ( .A(out[803]), .B(n1614), .Z(N815) );
  AND U7489 ( .A(out[804]), .B(n1614), .Z(N816) );
  AND U7490 ( .A(out[805]), .B(n1614), .Z(N817) );
  AND U7491 ( .A(out[806]), .B(n1614), .Z(N818) );
  AND U7492 ( .A(out[807]), .B(n1614), .Z(N819) );
  AND U7493 ( .A(out[70]), .B(n1614), .Z(N82) );
  AND U7494 ( .A(out[808]), .B(n1614), .Z(N820) );
  AND U7495 ( .A(out[809]), .B(n1614), .Z(N821) );
  AND U7496 ( .A(out[810]), .B(n1614), .Z(N822) );
  AND U7497 ( .A(out[811]), .B(n1614), .Z(N823) );
  AND U7498 ( .A(out[812]), .B(n1614), .Z(N824) );
  AND U7499 ( .A(out[813]), .B(n1614), .Z(N825) );
  AND U7500 ( .A(out[814]), .B(n1614), .Z(N826) );
  AND U7501 ( .A(out[815]), .B(n1614), .Z(N827) );
  AND U7502 ( .A(out[816]), .B(n1614), .Z(N828) );
  AND U7503 ( .A(out[817]), .B(n1614), .Z(N829) );
  AND U7504 ( .A(out[71]), .B(n1614), .Z(N83) );
  AND U7505 ( .A(out[818]), .B(n1614), .Z(N830) );
  AND U7506 ( .A(out[819]), .B(n1614), .Z(N831) );
  AND U7507 ( .A(out[820]), .B(n1614), .Z(N832) );
  AND U7508 ( .A(out[821]), .B(n1614), .Z(N833) );
  AND U7509 ( .A(out[822]), .B(n1614), .Z(N834) );
  AND U7510 ( .A(out[823]), .B(n1614), .Z(N835) );
  AND U7511 ( .A(out[824]), .B(n1614), .Z(N836) );
  AND U7512 ( .A(out[825]), .B(n1614), .Z(N837) );
  AND U7513 ( .A(out[826]), .B(n1614), .Z(N838) );
  AND U7514 ( .A(out[827]), .B(n1614), .Z(N839) );
  AND U7515 ( .A(out[72]), .B(n1614), .Z(N84) );
  AND U7516 ( .A(out[828]), .B(n1614), .Z(N840) );
  AND U7517 ( .A(out[829]), .B(n1614), .Z(N841) );
  AND U7518 ( .A(out[830]), .B(n1614), .Z(N842) );
  AND U7519 ( .A(out[831]), .B(n1614), .Z(N843) );
  AND U7520 ( .A(out[832]), .B(n1614), .Z(N844) );
  AND U7521 ( .A(out[833]), .B(n1614), .Z(N845) );
  AND U7522 ( .A(out[834]), .B(n1614), .Z(N846) );
  AND U7523 ( .A(out[835]), .B(n1614), .Z(N847) );
  AND U7524 ( .A(out[836]), .B(n1614), .Z(N848) );
  AND U7525 ( .A(out[837]), .B(n1614), .Z(N849) );
  AND U7526 ( .A(out[73]), .B(n1614), .Z(N85) );
  AND U7527 ( .A(out[838]), .B(n1614), .Z(N850) );
  AND U7528 ( .A(out[839]), .B(n1614), .Z(N851) );
  AND U7529 ( .A(out[840]), .B(n1614), .Z(N852) );
  AND U7530 ( .A(out[841]), .B(n1614), .Z(N853) );
  AND U7531 ( .A(out[842]), .B(n1614), .Z(N854) );
  AND U7532 ( .A(out[843]), .B(n1614), .Z(N855) );
  AND U7533 ( .A(out[844]), .B(n1614), .Z(N856) );
  AND U7534 ( .A(out[845]), .B(n1614), .Z(N857) );
  AND U7535 ( .A(out[846]), .B(n1614), .Z(N858) );
  AND U7536 ( .A(out[847]), .B(n1614), .Z(N859) );
  AND U7537 ( .A(out[74]), .B(n1614), .Z(N86) );
  AND U7538 ( .A(out[848]), .B(n1614), .Z(N860) );
  AND U7539 ( .A(out[849]), .B(n1614), .Z(N861) );
  AND U7540 ( .A(out[850]), .B(n1614), .Z(N862) );
  AND U7541 ( .A(out[851]), .B(n1614), .Z(N863) );
  AND U7542 ( .A(out[852]), .B(n1614), .Z(N864) );
  AND U7543 ( .A(out[853]), .B(n1614), .Z(N865) );
  AND U7544 ( .A(out[854]), .B(n1614), .Z(N866) );
  AND U7545 ( .A(out[855]), .B(n1614), .Z(N867) );
  AND U7546 ( .A(out[856]), .B(n1614), .Z(N868) );
  AND U7547 ( .A(out[857]), .B(n1614), .Z(N869) );
  AND U7548 ( .A(out[75]), .B(n1614), .Z(N87) );
  AND U7549 ( .A(out[858]), .B(n1614), .Z(N870) );
  AND U7550 ( .A(out[859]), .B(n1614), .Z(N871) );
  AND U7551 ( .A(out[860]), .B(n1614), .Z(N872) );
  AND U7552 ( .A(out[861]), .B(n1614), .Z(N873) );
  AND U7553 ( .A(out[862]), .B(n1614), .Z(N874) );
  AND U7554 ( .A(out[863]), .B(n1614), .Z(N875) );
  AND U7555 ( .A(out[864]), .B(n1614), .Z(N876) );
  AND U7556 ( .A(out[865]), .B(n1614), .Z(N877) );
  AND U7557 ( .A(out[866]), .B(n1614), .Z(N878) );
  AND U7558 ( .A(out[867]), .B(n1614), .Z(N879) );
  AND U7559 ( .A(out[76]), .B(n1614), .Z(N88) );
  AND U7560 ( .A(out[868]), .B(n1614), .Z(N880) );
  AND U7561 ( .A(out[869]), .B(n1614), .Z(N881) );
  AND U7562 ( .A(out[870]), .B(n1614), .Z(N882) );
  AND U7563 ( .A(out[871]), .B(n1614), .Z(N883) );
  AND U7564 ( .A(out[872]), .B(n1614), .Z(N884) );
  AND U7565 ( .A(out[873]), .B(n1614), .Z(N885) );
  AND U7566 ( .A(out[874]), .B(n1614), .Z(N886) );
  AND U7567 ( .A(out[875]), .B(n1614), .Z(N887) );
  AND U7568 ( .A(out[876]), .B(n1614), .Z(N888) );
  AND U7569 ( .A(out[877]), .B(n1614), .Z(N889) );
  AND U7570 ( .A(out[77]), .B(n1614), .Z(N89) );
  AND U7571 ( .A(out[878]), .B(n1614), .Z(N890) );
  AND U7572 ( .A(out[879]), .B(n1614), .Z(N891) );
  AND U7573 ( .A(out[880]), .B(n1614), .Z(N892) );
  AND U7574 ( .A(out[881]), .B(n1614), .Z(N893) );
  AND U7575 ( .A(out[882]), .B(n1614), .Z(N894) );
  AND U7576 ( .A(out[883]), .B(n1614), .Z(N895) );
  AND U7577 ( .A(out[884]), .B(n1614), .Z(N896) );
  AND U7578 ( .A(out[885]), .B(n1614), .Z(N897) );
  AND U7579 ( .A(out[886]), .B(n1614), .Z(N898) );
  AND U7580 ( .A(out[887]), .B(n1614), .Z(N899) );
  AND U7581 ( .A(rc_i[2]), .B(n1614), .Z(N9) );
  AND U7582 ( .A(out[78]), .B(n1614), .Z(N90) );
  AND U7583 ( .A(out[888]), .B(n1614), .Z(N900) );
  AND U7584 ( .A(out[889]), .B(n1614), .Z(N901) );
  AND U7585 ( .A(out[890]), .B(n1614), .Z(N902) );
  AND U7586 ( .A(out[891]), .B(n1614), .Z(N903) );
  AND U7587 ( .A(out[892]), .B(n1614), .Z(N904) );
  AND U7588 ( .A(out[893]), .B(n1614), .Z(N905) );
  AND U7589 ( .A(out[894]), .B(n1614), .Z(N906) );
  AND U7590 ( .A(out[895]), .B(n1614), .Z(N907) );
  AND U7591 ( .A(out[896]), .B(n1614), .Z(N908) );
  AND U7592 ( .A(out[897]), .B(n1614), .Z(N909) );
  AND U7593 ( .A(out[79]), .B(n1614), .Z(N91) );
  AND U7594 ( .A(out[898]), .B(n1614), .Z(N910) );
  AND U7595 ( .A(out[899]), .B(n1614), .Z(N911) );
  AND U7596 ( .A(out[900]), .B(n1614), .Z(N912) );
  AND U7597 ( .A(out[901]), .B(n1614), .Z(N913) );
  AND U7598 ( .A(out[902]), .B(n1614), .Z(N914) );
  AND U7599 ( .A(out[903]), .B(n1614), .Z(N915) );
  AND U7600 ( .A(out[904]), .B(n1614), .Z(N916) );
  AND U7601 ( .A(out[905]), .B(n1614), .Z(N917) );
  AND U7602 ( .A(out[906]), .B(n1614), .Z(N918) );
  AND U7603 ( .A(out[907]), .B(n1614), .Z(N919) );
  AND U7604 ( .A(out[80]), .B(n1614), .Z(N92) );
  AND U7605 ( .A(out[908]), .B(n1614), .Z(N920) );
  AND U7606 ( .A(out[909]), .B(n1614), .Z(N921) );
  AND U7607 ( .A(out[910]), .B(n1614), .Z(N922) );
  AND U7608 ( .A(out[911]), .B(n1614), .Z(N923) );
  AND U7609 ( .A(out[912]), .B(n1614), .Z(N924) );
  AND U7610 ( .A(out[913]), .B(n1614), .Z(N925) );
  AND U7611 ( .A(out[914]), .B(n1614), .Z(N926) );
  AND U7612 ( .A(out[915]), .B(n1614), .Z(N927) );
  AND U7613 ( .A(out[916]), .B(n1614), .Z(N928) );
  AND U7614 ( .A(out[917]), .B(n1614), .Z(N929) );
  AND U7615 ( .A(out[81]), .B(n1614), .Z(N93) );
  AND U7616 ( .A(out[918]), .B(n1614), .Z(N930) );
  AND U7617 ( .A(out[919]), .B(n1614), .Z(N931) );
  AND U7618 ( .A(out[920]), .B(n1614), .Z(N932) );
  AND U7619 ( .A(out[921]), .B(n1614), .Z(N933) );
  AND U7620 ( .A(out[922]), .B(n1614), .Z(N934) );
  AND U7621 ( .A(out[923]), .B(n1614), .Z(N935) );
  AND U7622 ( .A(out[924]), .B(n1614), .Z(N936) );
  AND U7623 ( .A(out[925]), .B(n1614), .Z(N937) );
  AND U7624 ( .A(out[926]), .B(n1614), .Z(N938) );
  AND U7625 ( .A(out[927]), .B(n1614), .Z(N939) );
  AND U7626 ( .A(out[82]), .B(n1614), .Z(N94) );
  AND U7627 ( .A(out[928]), .B(n1614), .Z(N940) );
  AND U7628 ( .A(out[929]), .B(n1614), .Z(N941) );
  AND U7629 ( .A(out[930]), .B(n1614), .Z(N942) );
  AND U7630 ( .A(out[931]), .B(n1614), .Z(N943) );
  AND U7631 ( .A(out[932]), .B(n1614), .Z(N944) );
  AND U7632 ( .A(out[933]), .B(n1614), .Z(N945) );
  AND U7633 ( .A(out[934]), .B(n1614), .Z(N946) );
  AND U7634 ( .A(out[935]), .B(n1614), .Z(N947) );
  AND U7635 ( .A(out[936]), .B(n1614), .Z(N948) );
  AND U7636 ( .A(out[937]), .B(n1614), .Z(N949) );
  AND U7637 ( .A(out[83]), .B(n1614), .Z(N95) );
  AND U7638 ( .A(out[938]), .B(n1614), .Z(N950) );
  AND U7639 ( .A(out[939]), .B(n1614), .Z(N951) );
  AND U7640 ( .A(out[940]), .B(n1614), .Z(N952) );
  AND U7641 ( .A(out[941]), .B(n1614), .Z(N953) );
  AND U7642 ( .A(out[942]), .B(n1614), .Z(N954) );
  AND U7643 ( .A(out[943]), .B(n1614), .Z(N955) );
  AND U7644 ( .A(out[944]), .B(n1614), .Z(N956) );
  AND U7645 ( .A(out[945]), .B(n1614), .Z(N957) );
  AND U7646 ( .A(out[946]), .B(n1614), .Z(N958) );
  AND U7647 ( .A(out[947]), .B(n1614), .Z(N959) );
  AND U7648 ( .A(out[84]), .B(n1614), .Z(N96) );
  AND U7649 ( .A(out[948]), .B(n1614), .Z(N960) );
  AND U7650 ( .A(out[949]), .B(n1614), .Z(N961) );
  AND U7651 ( .A(out[950]), .B(n1614), .Z(N962) );
  AND U7652 ( .A(out[951]), .B(n1614), .Z(N963) );
  AND U7653 ( .A(out[952]), .B(n1614), .Z(N964) );
  AND U7654 ( .A(out[953]), .B(n1614), .Z(N965) );
  AND U7655 ( .A(out[954]), .B(n1614), .Z(N966) );
  AND U7656 ( .A(out[955]), .B(n1614), .Z(N967) );
  AND U7657 ( .A(out[956]), .B(n1614), .Z(N968) );
  AND U7658 ( .A(out[957]), .B(n1614), .Z(N969) );
  AND U7659 ( .A(out[85]), .B(n1614), .Z(N97) );
  AND U7660 ( .A(out[958]), .B(n1614), .Z(N970) );
  AND U7661 ( .A(out[959]), .B(n1614), .Z(N971) );
  AND U7662 ( .A(out[960]), .B(n1614), .Z(N972) );
  AND U7663 ( .A(out[961]), .B(n1614), .Z(N973) );
  AND U7664 ( .A(out[962]), .B(n1614), .Z(N974) );
  AND U7665 ( .A(out[963]), .B(n1614), .Z(N975) );
  AND U7666 ( .A(out[964]), .B(n1614), .Z(N976) );
  AND U7667 ( .A(out[965]), .B(n1614), .Z(N977) );
  AND U7668 ( .A(out[966]), .B(n1614), .Z(N978) );
  AND U7669 ( .A(out[967]), .B(n1614), .Z(N979) );
  AND U7670 ( .A(out[86]), .B(n1614), .Z(N98) );
  AND U7671 ( .A(out[968]), .B(n1614), .Z(N980) );
  AND U7672 ( .A(out[969]), .B(n1614), .Z(N981) );
  AND U7673 ( .A(out[970]), .B(n1614), .Z(N982) );
  AND U7674 ( .A(out[971]), .B(n1614), .Z(N983) );
  AND U7675 ( .A(out[972]), .B(n1614), .Z(N984) );
  AND U7676 ( .A(out[973]), .B(n1614), .Z(N985) );
  AND U7677 ( .A(out[974]), .B(n1614), .Z(N986) );
  AND U7678 ( .A(out[975]), .B(n1614), .Z(N987) );
  AND U7679 ( .A(out[976]), .B(n1614), .Z(N988) );
  AND U7680 ( .A(out[977]), .B(n1614), .Z(N989) );
  AND U7681 ( .A(out[87]), .B(n1614), .Z(N99) );
  AND U7682 ( .A(out[978]), .B(n1614), .Z(N990) );
  AND U7683 ( .A(out[979]), .B(n1614), .Z(N991) );
  AND U7684 ( .A(out[980]), .B(n1614), .Z(N992) );
  AND U7685 ( .A(out[981]), .B(n1614), .Z(N993) );
  AND U7686 ( .A(out[982]), .B(n1614), .Z(N994) );
  AND U7687 ( .A(out[983]), .B(n1614), .Z(N995) );
  AND U7688 ( .A(out[984]), .B(n1614), .Z(N996) );
  AND U7689 ( .A(out[985]), .B(n1614), .Z(N997) );
  AND U7690 ( .A(out[986]), .B(n1614), .Z(N998) );
  AND U7691 ( .A(out[987]), .B(n1614), .Z(N999) );
  NOR U7692 ( .A(rc_i[3]), .B(rc_i[1]), .Z(n2854) );
  IV U7693 ( .A(n2854), .Z(\RCONST[3].rconst_/N10 ) );
  OR U7694 ( .A(rc_i[5]), .B(rc_i[0]), .Z(\RCONST[1].rconst_/N49 ) );
  NANDN U7695 ( .A(\RCONST[1].rconst_/N49 ), .B(n2854), .Z(\rc[3][15] ) );
  OR U7696 ( .A(rc_i[2]), .B(rc_i[3]), .Z(\RCONST[1].rconst_/N26 ) );
  OR U7697 ( .A(\RCONST[1].rconst_/N26 ), .B(rc_i[4]), .Z(\rc[3][1] ) );
  NOR U7698 ( .A(\RCONST[1].rconst_/N26 ), .B(rc_i[1]), .Z(n2853) );
  IV U7699 ( .A(rc_i[4]), .Z(n2856) );
  NAND U7700 ( .A(n2853), .B(n2856), .Z(\RCONST[0].rconst_/N17 ) );
  IV U7701 ( .A(n2853), .Z(\RCONST[0].rconst_/N25 ) );
  NOR U7702 ( .A(rc_i[2]), .B(rc_i[5]), .Z(n2855) );
  NANDN U7703 ( .A(rc_i[1]), .B(n2855), .Z(\RCONST[2].rconst_/N57 ) );
  NAND U7704 ( .A(n2854), .B(n2855), .Z(\rc[2][0] ) );
  NANDN U7705 ( .A(rc_i[5]), .B(n2856), .Z(\RCONST[0].rconst_/N67 ) );
  OR U7706 ( .A(rc_i[5]), .B(rc_i[3]), .Z(\RCONST[0].rconst_/N56 ) );
  OR U7707 ( .A(\RCONST[0].rconst_/N56 ), .B(rc_i[4]), .Z(
        \RCONST[1].rconst_/N68 ) );
  OR U7708 ( .A(\RCONST[0].rconst_/N67 ), .B(\RCONST[3].rconst_/N10 ), .Z(
        \RCONST[0].rconst_/N48 ) );
  OR U7709 ( .A(rc_i[3]), .B(rc_i[0]), .Z(\RCONST[1].rconst_/N15 ) );
  OR U7710 ( .A(\RCONST[2].rconst_/N18 ), .B(\RCONST[1].rconst_/N26 ), .Z(
        \RCONST[2].rconst_/N28 ) );
  OR U7711 ( .A(\RCONST[2].rconst_/N18 ), .B(\RCONST[0].rconst_/N25 ), .Z(
        \RCONST[2].rconst_/N47 ) );
  NANDN U7712 ( .A(\RCONST[2].rconst_/N18 ), .B(n2855), .Z(\rc[3][31] ) );
  OR U7713 ( .A(\RCONST[1].rconst_/N49 ), .B(\rc[3][1] ), .Z(\rc[1][7] ) );
  OR U7714 ( .A(\RCONST[2].rconst_/N57 ), .B(rc_i[4]), .Z(\rc[3][3] ) );
  NAND U7715 ( .A(init), .B(round_reg[0]), .Z(n2858) );
  NAND U7716 ( .A(n2770), .B(in[0]), .Z(n2857) );
  NAND U7717 ( .A(n2858), .B(n2857), .Z(\round_in[0][0] ) );
  AND U7718 ( .A(round_reg[1000]), .B(init), .Z(\round_in[0][1000] ) );
  AND U7719 ( .A(round_reg[1001]), .B(init), .Z(\round_in[0][1001] ) );
  AND U7720 ( .A(round_reg[1002]), .B(init), .Z(\round_in[0][1002] ) );
  AND U7721 ( .A(round_reg[1003]), .B(init), .Z(\round_in[0][1003] ) );
  AND U7722 ( .A(round_reg[1004]), .B(init), .Z(\round_in[0][1004] ) );
  AND U7723 ( .A(round_reg[1005]), .B(init), .Z(\round_in[0][1005] ) );
  AND U7724 ( .A(round_reg[1006]), .B(init), .Z(\round_in[0][1006] ) );
  AND U7725 ( .A(round_reg[1007]), .B(init), .Z(\round_in[0][1007] ) );
  AND U7726 ( .A(round_reg[1008]), .B(init), .Z(\round_in[0][1008] ) );
  AND U7727 ( .A(round_reg[1009]), .B(init), .Z(\round_in[0][1009] ) );
  NAND U7728 ( .A(init), .B(round_reg[100]), .Z(n2860) );
  NAND U7729 ( .A(n2770), .B(in[100]), .Z(n2859) );
  NAND U7730 ( .A(n2860), .B(n2859), .Z(\round_in[0][100] ) );
  AND U7731 ( .A(round_reg[1010]), .B(init), .Z(\round_in[0][1010] ) );
  AND U7732 ( .A(round_reg[1011]), .B(init), .Z(\round_in[0][1011] ) );
  AND U7733 ( .A(round_reg[1012]), .B(init), .Z(\round_in[0][1012] ) );
  AND U7734 ( .A(round_reg[1013]), .B(init), .Z(\round_in[0][1013] ) );
  AND U7735 ( .A(round_reg[1014]), .B(init), .Z(\round_in[0][1014] ) );
  AND U7736 ( .A(round_reg[1015]), .B(init), .Z(\round_in[0][1015] ) );
  AND U7737 ( .A(round_reg[1016]), .B(init), .Z(\round_in[0][1016] ) );
  AND U7738 ( .A(round_reg[1017]), .B(init), .Z(\round_in[0][1017] ) );
  AND U7739 ( .A(round_reg[1018]), .B(init), .Z(\round_in[0][1018] ) );
  AND U7740 ( .A(round_reg[1019]), .B(init), .Z(\round_in[0][1019] ) );
  NAND U7741 ( .A(init), .B(round_reg[101]), .Z(n2862) );
  NAND U7742 ( .A(n2770), .B(in[101]), .Z(n2861) );
  NAND U7743 ( .A(n2862), .B(n2861), .Z(\round_in[0][101] ) );
  AND U7744 ( .A(round_reg[1020]), .B(init), .Z(\round_in[0][1020] ) );
  AND U7745 ( .A(round_reg[1021]), .B(init), .Z(\round_in[0][1021] ) );
  AND U7746 ( .A(round_reg[1022]), .B(init), .Z(\round_in[0][1022] ) );
  AND U7747 ( .A(round_reg[1023]), .B(init), .Z(\round_in[0][1023] ) );
  AND U7748 ( .A(round_reg[1024]), .B(init), .Z(\round_in[0][1024] ) );
  AND U7749 ( .A(round_reg[1025]), .B(init), .Z(\round_in[0][1025] ) );
  AND U7750 ( .A(round_reg[1026]), .B(init), .Z(\round_in[0][1026] ) );
  AND U7751 ( .A(round_reg[1027]), .B(init), .Z(\round_in[0][1027] ) );
  AND U7752 ( .A(round_reg[1028]), .B(init), .Z(\round_in[0][1028] ) );
  AND U7753 ( .A(round_reg[1029]), .B(init), .Z(\round_in[0][1029] ) );
  NAND U7754 ( .A(init), .B(round_reg[102]), .Z(n2864) );
  NAND U7755 ( .A(n2770), .B(in[102]), .Z(n2863) );
  NAND U7756 ( .A(n2864), .B(n2863), .Z(\round_in[0][102] ) );
  AND U7757 ( .A(round_reg[1030]), .B(init), .Z(\round_in[0][1030] ) );
  AND U7758 ( .A(round_reg[1031]), .B(init), .Z(\round_in[0][1031] ) );
  AND U7759 ( .A(round_reg[1032]), .B(init), .Z(\round_in[0][1032] ) );
  AND U7760 ( .A(round_reg[1033]), .B(init), .Z(\round_in[0][1033] ) );
  AND U7761 ( .A(round_reg[1034]), .B(init), .Z(\round_in[0][1034] ) );
  AND U7762 ( .A(round_reg[1035]), .B(init), .Z(\round_in[0][1035] ) );
  AND U7763 ( .A(round_reg[1036]), .B(init), .Z(\round_in[0][1036] ) );
  AND U7764 ( .A(round_reg[1037]), .B(init), .Z(\round_in[0][1037] ) );
  AND U7765 ( .A(round_reg[1038]), .B(init), .Z(\round_in[0][1038] ) );
  AND U7766 ( .A(round_reg[1039]), .B(init), .Z(\round_in[0][1039] ) );
  NAND U7767 ( .A(init), .B(round_reg[103]), .Z(n2866) );
  NAND U7768 ( .A(n2770), .B(in[103]), .Z(n2865) );
  NAND U7769 ( .A(n2866), .B(n2865), .Z(\round_in[0][103] ) );
  AND U7770 ( .A(round_reg[1040]), .B(init), .Z(\round_in[0][1040] ) );
  AND U7771 ( .A(round_reg[1041]), .B(init), .Z(\round_in[0][1041] ) );
  AND U7772 ( .A(round_reg[1042]), .B(init), .Z(\round_in[0][1042] ) );
  AND U7773 ( .A(round_reg[1043]), .B(init), .Z(\round_in[0][1043] ) );
  AND U7774 ( .A(round_reg[1044]), .B(init), .Z(\round_in[0][1044] ) );
  AND U7775 ( .A(round_reg[1045]), .B(init), .Z(\round_in[0][1045] ) );
  AND U7776 ( .A(round_reg[1046]), .B(init), .Z(\round_in[0][1046] ) );
  AND U7777 ( .A(round_reg[1047]), .B(init), .Z(\round_in[0][1047] ) );
  AND U7778 ( .A(round_reg[1048]), .B(init), .Z(\round_in[0][1048] ) );
  AND U7779 ( .A(round_reg[1049]), .B(init), .Z(\round_in[0][1049] ) );
  NAND U7780 ( .A(init), .B(round_reg[104]), .Z(n2868) );
  NAND U7781 ( .A(n2771), .B(in[104]), .Z(n2867) );
  NAND U7782 ( .A(n2868), .B(n2867), .Z(\round_in[0][104] ) );
  AND U7783 ( .A(round_reg[1050]), .B(init), .Z(\round_in[0][1050] ) );
  AND U7784 ( .A(round_reg[1051]), .B(init), .Z(\round_in[0][1051] ) );
  AND U7785 ( .A(round_reg[1052]), .B(init), .Z(\round_in[0][1052] ) );
  AND U7786 ( .A(round_reg[1053]), .B(init), .Z(\round_in[0][1053] ) );
  AND U7787 ( .A(round_reg[1054]), .B(init), .Z(\round_in[0][1054] ) );
  AND U7788 ( .A(round_reg[1055]), .B(init), .Z(\round_in[0][1055] ) );
  AND U7789 ( .A(round_reg[1056]), .B(init), .Z(\round_in[0][1056] ) );
  AND U7790 ( .A(round_reg[1057]), .B(init), .Z(\round_in[0][1057] ) );
  AND U7791 ( .A(round_reg[1058]), .B(init), .Z(\round_in[0][1058] ) );
  AND U7792 ( .A(round_reg[1059]), .B(init), .Z(\round_in[0][1059] ) );
  NAND U7793 ( .A(init), .B(round_reg[105]), .Z(n2870) );
  NAND U7794 ( .A(n2771), .B(in[105]), .Z(n2869) );
  NAND U7795 ( .A(n2870), .B(n2869), .Z(\round_in[0][105] ) );
  AND U7796 ( .A(round_reg[1060]), .B(init), .Z(\round_in[0][1060] ) );
  AND U7797 ( .A(round_reg[1061]), .B(init), .Z(\round_in[0][1061] ) );
  AND U7798 ( .A(round_reg[1062]), .B(init), .Z(\round_in[0][1062] ) );
  AND U7799 ( .A(round_reg[1063]), .B(init), .Z(\round_in[0][1063] ) );
  AND U7800 ( .A(round_reg[1064]), .B(init), .Z(\round_in[0][1064] ) );
  AND U7801 ( .A(round_reg[1065]), .B(init), .Z(\round_in[0][1065] ) );
  AND U7802 ( .A(round_reg[1066]), .B(init), .Z(\round_in[0][1066] ) );
  AND U7803 ( .A(round_reg[1067]), .B(init), .Z(\round_in[0][1067] ) );
  AND U7804 ( .A(round_reg[1068]), .B(init), .Z(\round_in[0][1068] ) );
  AND U7805 ( .A(round_reg[1069]), .B(init), .Z(\round_in[0][1069] ) );
  NAND U7806 ( .A(init), .B(round_reg[106]), .Z(n2872) );
  NAND U7807 ( .A(n2771), .B(in[106]), .Z(n2871) );
  NAND U7808 ( .A(n2872), .B(n2871), .Z(\round_in[0][106] ) );
  AND U7809 ( .A(round_reg[1070]), .B(init), .Z(\round_in[0][1070] ) );
  AND U7810 ( .A(round_reg[1071]), .B(init), .Z(\round_in[0][1071] ) );
  AND U7811 ( .A(round_reg[1072]), .B(init), .Z(\round_in[0][1072] ) );
  AND U7812 ( .A(round_reg[1073]), .B(init), .Z(\round_in[0][1073] ) );
  AND U7813 ( .A(round_reg[1074]), .B(init), .Z(\round_in[0][1074] ) );
  AND U7814 ( .A(round_reg[1075]), .B(init), .Z(\round_in[0][1075] ) );
  AND U7815 ( .A(round_reg[1076]), .B(init), .Z(\round_in[0][1076] ) );
  AND U7816 ( .A(round_reg[1077]), .B(init), .Z(\round_in[0][1077] ) );
  AND U7817 ( .A(round_reg[1078]), .B(init), .Z(\round_in[0][1078] ) );
  AND U7818 ( .A(round_reg[1079]), .B(init), .Z(\round_in[0][1079] ) );
  NAND U7819 ( .A(init), .B(round_reg[107]), .Z(n2874) );
  NAND U7820 ( .A(n2771), .B(in[107]), .Z(n2873) );
  NAND U7821 ( .A(n2874), .B(n2873), .Z(\round_in[0][107] ) );
  AND U7822 ( .A(round_reg[1080]), .B(init), .Z(\round_in[0][1080] ) );
  AND U7823 ( .A(round_reg[1081]), .B(init), .Z(\round_in[0][1081] ) );
  AND U7824 ( .A(round_reg[1082]), .B(init), .Z(\round_in[0][1082] ) );
  AND U7825 ( .A(round_reg[1083]), .B(init), .Z(\round_in[0][1083] ) );
  AND U7826 ( .A(round_reg[1084]), .B(init), .Z(\round_in[0][1084] ) );
  AND U7827 ( .A(round_reg[1085]), .B(init), .Z(\round_in[0][1085] ) );
  AND U7828 ( .A(round_reg[1086]), .B(init), .Z(\round_in[0][1086] ) );
  AND U7829 ( .A(round_reg[1087]), .B(init), .Z(\round_in[0][1087] ) );
  AND U7830 ( .A(round_reg[1088]), .B(init), .Z(\round_in[0][1088] ) );
  AND U7831 ( .A(round_reg[1089]), .B(init), .Z(\round_in[0][1089] ) );
  NAND U7832 ( .A(init), .B(round_reg[108]), .Z(n2876) );
  NAND U7833 ( .A(n2771), .B(in[108]), .Z(n2875) );
  NAND U7834 ( .A(n2876), .B(n2875), .Z(\round_in[0][108] ) );
  AND U7835 ( .A(round_reg[1090]), .B(init), .Z(\round_in[0][1090] ) );
  AND U7836 ( .A(round_reg[1091]), .B(init), .Z(\round_in[0][1091] ) );
  AND U7837 ( .A(round_reg[1092]), .B(init), .Z(\round_in[0][1092] ) );
  AND U7838 ( .A(round_reg[1093]), .B(init), .Z(\round_in[0][1093] ) );
  AND U7839 ( .A(round_reg[1094]), .B(init), .Z(\round_in[0][1094] ) );
  AND U7840 ( .A(round_reg[1095]), .B(init), .Z(\round_in[0][1095] ) );
  AND U7841 ( .A(round_reg[1096]), .B(init), .Z(\round_in[0][1096] ) );
  AND U7842 ( .A(round_reg[1097]), .B(init), .Z(\round_in[0][1097] ) );
  AND U7843 ( .A(round_reg[1098]), .B(init), .Z(\round_in[0][1098] ) );
  AND U7844 ( .A(round_reg[1099]), .B(init), .Z(\round_in[0][1099] ) );
  NAND U7845 ( .A(init), .B(round_reg[109]), .Z(n2878) );
  NAND U7846 ( .A(n2771), .B(in[109]), .Z(n2877) );
  NAND U7847 ( .A(n2878), .B(n2877), .Z(\round_in[0][109] ) );
  NAND U7848 ( .A(init), .B(round_reg[10]), .Z(n2880) );
  NAND U7849 ( .A(n2771), .B(in[10]), .Z(n2879) );
  NAND U7850 ( .A(n2880), .B(n2879), .Z(\round_in[0][10] ) );
  AND U7851 ( .A(round_reg[1100]), .B(init), .Z(\round_in[0][1100] ) );
  AND U7852 ( .A(round_reg[1101]), .B(init), .Z(\round_in[0][1101] ) );
  AND U7853 ( .A(round_reg[1102]), .B(init), .Z(\round_in[0][1102] ) );
  AND U7854 ( .A(round_reg[1103]), .B(init), .Z(\round_in[0][1103] ) );
  AND U7855 ( .A(round_reg[1104]), .B(init), .Z(\round_in[0][1104] ) );
  AND U7856 ( .A(round_reg[1105]), .B(init), .Z(\round_in[0][1105] ) );
  AND U7857 ( .A(round_reg[1106]), .B(init), .Z(\round_in[0][1106] ) );
  AND U7858 ( .A(round_reg[1107]), .B(init), .Z(\round_in[0][1107] ) );
  AND U7859 ( .A(round_reg[1108]), .B(init), .Z(\round_in[0][1108] ) );
  AND U7860 ( .A(round_reg[1109]), .B(init), .Z(\round_in[0][1109] ) );
  NAND U7861 ( .A(init), .B(round_reg[110]), .Z(n2882) );
  NAND U7862 ( .A(n2772), .B(in[110]), .Z(n2881) );
  NAND U7863 ( .A(n2882), .B(n2881), .Z(\round_in[0][110] ) );
  AND U7864 ( .A(round_reg[1110]), .B(init), .Z(\round_in[0][1110] ) );
  AND U7865 ( .A(round_reg[1111]), .B(init), .Z(\round_in[0][1111] ) );
  AND U7866 ( .A(round_reg[1112]), .B(init), .Z(\round_in[0][1112] ) );
  AND U7867 ( .A(round_reg[1113]), .B(init), .Z(\round_in[0][1113] ) );
  AND U7868 ( .A(round_reg[1114]), .B(init), .Z(\round_in[0][1114] ) );
  AND U7869 ( .A(round_reg[1115]), .B(init), .Z(\round_in[0][1115] ) );
  AND U7870 ( .A(round_reg[1116]), .B(init), .Z(\round_in[0][1116] ) );
  AND U7871 ( .A(round_reg[1117]), .B(init), .Z(\round_in[0][1117] ) );
  AND U7872 ( .A(round_reg[1118]), .B(init), .Z(\round_in[0][1118] ) );
  AND U7873 ( .A(round_reg[1119]), .B(init), .Z(\round_in[0][1119] ) );
  NAND U7874 ( .A(init), .B(round_reg[111]), .Z(n2884) );
  NAND U7875 ( .A(n2772), .B(in[111]), .Z(n2883) );
  NAND U7876 ( .A(n2884), .B(n2883), .Z(\round_in[0][111] ) );
  AND U7877 ( .A(round_reg[1120]), .B(init), .Z(\round_in[0][1120] ) );
  AND U7878 ( .A(round_reg[1121]), .B(init), .Z(\round_in[0][1121] ) );
  AND U7879 ( .A(round_reg[1122]), .B(init), .Z(\round_in[0][1122] ) );
  AND U7880 ( .A(round_reg[1123]), .B(init), .Z(\round_in[0][1123] ) );
  AND U7881 ( .A(round_reg[1124]), .B(init), .Z(\round_in[0][1124] ) );
  AND U7882 ( .A(round_reg[1125]), .B(init), .Z(\round_in[0][1125] ) );
  AND U7883 ( .A(round_reg[1126]), .B(init), .Z(\round_in[0][1126] ) );
  AND U7884 ( .A(round_reg[1127]), .B(init), .Z(\round_in[0][1127] ) );
  AND U7885 ( .A(round_reg[1128]), .B(init), .Z(\round_in[0][1128] ) );
  AND U7886 ( .A(round_reg[1129]), .B(init), .Z(\round_in[0][1129] ) );
  NAND U7887 ( .A(init), .B(round_reg[112]), .Z(n2886) );
  NAND U7888 ( .A(n2772), .B(in[112]), .Z(n2885) );
  NAND U7889 ( .A(n2886), .B(n2885), .Z(\round_in[0][112] ) );
  AND U7890 ( .A(round_reg[1130]), .B(init), .Z(\round_in[0][1130] ) );
  AND U7891 ( .A(round_reg[1131]), .B(init), .Z(\round_in[0][1131] ) );
  AND U7892 ( .A(round_reg[1132]), .B(init), .Z(\round_in[0][1132] ) );
  AND U7893 ( .A(round_reg[1133]), .B(init), .Z(\round_in[0][1133] ) );
  AND U7894 ( .A(round_reg[1134]), .B(init), .Z(\round_in[0][1134] ) );
  AND U7895 ( .A(round_reg[1135]), .B(init), .Z(\round_in[0][1135] ) );
  AND U7896 ( .A(round_reg[1136]), .B(init), .Z(\round_in[0][1136] ) );
  AND U7897 ( .A(round_reg[1137]), .B(init), .Z(\round_in[0][1137] ) );
  AND U7898 ( .A(round_reg[1138]), .B(init), .Z(\round_in[0][1138] ) );
  AND U7899 ( .A(round_reg[1139]), .B(init), .Z(\round_in[0][1139] ) );
  NAND U7900 ( .A(init), .B(round_reg[113]), .Z(n2888) );
  NAND U7901 ( .A(n2772), .B(in[113]), .Z(n2887) );
  NAND U7902 ( .A(n2888), .B(n2887), .Z(\round_in[0][113] ) );
  AND U7903 ( .A(round_reg[1140]), .B(init), .Z(\round_in[0][1140] ) );
  AND U7904 ( .A(round_reg[1141]), .B(init), .Z(\round_in[0][1141] ) );
  AND U7905 ( .A(round_reg[1142]), .B(init), .Z(\round_in[0][1142] ) );
  AND U7906 ( .A(round_reg[1143]), .B(init), .Z(\round_in[0][1143] ) );
  AND U7907 ( .A(round_reg[1144]), .B(init), .Z(\round_in[0][1144] ) );
  AND U7908 ( .A(round_reg[1145]), .B(init), .Z(\round_in[0][1145] ) );
  AND U7909 ( .A(round_reg[1146]), .B(init), .Z(\round_in[0][1146] ) );
  AND U7910 ( .A(round_reg[1147]), .B(init), .Z(\round_in[0][1147] ) );
  AND U7911 ( .A(round_reg[1148]), .B(init), .Z(\round_in[0][1148] ) );
  AND U7912 ( .A(round_reg[1149]), .B(init), .Z(\round_in[0][1149] ) );
  NAND U7913 ( .A(init), .B(round_reg[114]), .Z(n2890) );
  NAND U7914 ( .A(n2772), .B(in[114]), .Z(n2889) );
  NAND U7915 ( .A(n2890), .B(n2889), .Z(\round_in[0][114] ) );
  AND U7916 ( .A(round_reg[1150]), .B(init), .Z(\round_in[0][1150] ) );
  AND U7917 ( .A(round_reg[1151]), .B(init), .Z(\round_in[0][1151] ) );
  AND U7918 ( .A(round_reg[1152]), .B(init), .Z(\round_in[0][1152] ) );
  AND U7919 ( .A(round_reg[1153]), .B(init), .Z(\round_in[0][1153] ) );
  AND U7920 ( .A(round_reg[1154]), .B(init), .Z(\round_in[0][1154] ) );
  AND U7921 ( .A(round_reg[1155]), .B(init), .Z(\round_in[0][1155] ) );
  AND U7922 ( .A(round_reg[1156]), .B(init), .Z(\round_in[0][1156] ) );
  AND U7923 ( .A(round_reg[1157]), .B(init), .Z(\round_in[0][1157] ) );
  AND U7924 ( .A(round_reg[1158]), .B(init), .Z(\round_in[0][1158] ) );
  AND U7925 ( .A(round_reg[1159]), .B(init), .Z(\round_in[0][1159] ) );
  NAND U7926 ( .A(init), .B(round_reg[115]), .Z(n2892) );
  NAND U7927 ( .A(n2772), .B(in[115]), .Z(n2891) );
  NAND U7928 ( .A(n2892), .B(n2891), .Z(\round_in[0][115] ) );
  AND U7929 ( .A(round_reg[1160]), .B(init), .Z(\round_in[0][1160] ) );
  AND U7930 ( .A(round_reg[1161]), .B(init), .Z(\round_in[0][1161] ) );
  AND U7931 ( .A(round_reg[1162]), .B(init), .Z(\round_in[0][1162] ) );
  AND U7932 ( .A(round_reg[1163]), .B(init), .Z(\round_in[0][1163] ) );
  AND U7933 ( .A(round_reg[1164]), .B(init), .Z(\round_in[0][1164] ) );
  AND U7934 ( .A(round_reg[1165]), .B(init), .Z(\round_in[0][1165] ) );
  AND U7935 ( .A(round_reg[1166]), .B(init), .Z(\round_in[0][1166] ) );
  AND U7936 ( .A(round_reg[1167]), .B(init), .Z(\round_in[0][1167] ) );
  AND U7937 ( .A(round_reg[1168]), .B(init), .Z(\round_in[0][1168] ) );
  AND U7938 ( .A(round_reg[1169]), .B(init), .Z(\round_in[0][1169] ) );
  NAND U7939 ( .A(init), .B(round_reg[116]), .Z(n2894) );
  NAND U7940 ( .A(n2772), .B(in[116]), .Z(n2893) );
  NAND U7941 ( .A(n2894), .B(n2893), .Z(\round_in[0][116] ) );
  AND U7942 ( .A(round_reg[1170]), .B(init), .Z(\round_in[0][1170] ) );
  AND U7943 ( .A(round_reg[1171]), .B(init), .Z(\round_in[0][1171] ) );
  AND U7944 ( .A(round_reg[1172]), .B(init), .Z(\round_in[0][1172] ) );
  AND U7945 ( .A(round_reg[1173]), .B(init), .Z(\round_in[0][1173] ) );
  AND U7946 ( .A(round_reg[1174]), .B(init), .Z(\round_in[0][1174] ) );
  AND U7947 ( .A(round_reg[1175]), .B(init), .Z(\round_in[0][1175] ) );
  AND U7948 ( .A(round_reg[1176]), .B(init), .Z(\round_in[0][1176] ) );
  AND U7949 ( .A(round_reg[1177]), .B(init), .Z(\round_in[0][1177] ) );
  AND U7950 ( .A(round_reg[1178]), .B(init), .Z(\round_in[0][1178] ) );
  AND U7951 ( .A(round_reg[1179]), .B(init), .Z(\round_in[0][1179] ) );
  NAND U7952 ( .A(init), .B(round_reg[117]), .Z(n2896) );
  NAND U7953 ( .A(n2773), .B(in[117]), .Z(n2895) );
  NAND U7954 ( .A(n2896), .B(n2895), .Z(\round_in[0][117] ) );
  AND U7955 ( .A(round_reg[1180]), .B(init), .Z(\round_in[0][1180] ) );
  AND U7956 ( .A(round_reg[1181]), .B(init), .Z(\round_in[0][1181] ) );
  AND U7957 ( .A(round_reg[1182]), .B(init), .Z(\round_in[0][1182] ) );
  AND U7958 ( .A(round_reg[1183]), .B(init), .Z(\round_in[0][1183] ) );
  AND U7959 ( .A(round_reg[1184]), .B(init), .Z(\round_in[0][1184] ) );
  AND U7960 ( .A(round_reg[1185]), .B(init), .Z(\round_in[0][1185] ) );
  AND U7961 ( .A(round_reg[1186]), .B(init), .Z(\round_in[0][1186] ) );
  AND U7962 ( .A(round_reg[1187]), .B(init), .Z(\round_in[0][1187] ) );
  AND U7963 ( .A(round_reg[1188]), .B(init), .Z(\round_in[0][1188] ) );
  AND U7964 ( .A(round_reg[1189]), .B(init), .Z(\round_in[0][1189] ) );
  NAND U7965 ( .A(init), .B(round_reg[118]), .Z(n2898) );
  NAND U7966 ( .A(n2773), .B(in[118]), .Z(n2897) );
  NAND U7967 ( .A(n2898), .B(n2897), .Z(\round_in[0][118] ) );
  AND U7968 ( .A(round_reg[1190]), .B(init), .Z(\round_in[0][1190] ) );
  AND U7969 ( .A(round_reg[1191]), .B(init), .Z(\round_in[0][1191] ) );
  AND U7970 ( .A(round_reg[1192]), .B(init), .Z(\round_in[0][1192] ) );
  AND U7971 ( .A(round_reg[1193]), .B(init), .Z(\round_in[0][1193] ) );
  AND U7972 ( .A(round_reg[1194]), .B(init), .Z(\round_in[0][1194] ) );
  AND U7973 ( .A(round_reg[1195]), .B(init), .Z(\round_in[0][1195] ) );
  AND U7974 ( .A(round_reg[1196]), .B(init), .Z(\round_in[0][1196] ) );
  AND U7975 ( .A(round_reg[1197]), .B(init), .Z(\round_in[0][1197] ) );
  AND U7976 ( .A(round_reg[1198]), .B(init), .Z(\round_in[0][1198] ) );
  AND U7977 ( .A(round_reg[1199]), .B(init), .Z(\round_in[0][1199] ) );
  NAND U7978 ( .A(init), .B(round_reg[119]), .Z(n2900) );
  NAND U7979 ( .A(n2773), .B(in[119]), .Z(n2899) );
  NAND U7980 ( .A(n2900), .B(n2899), .Z(\round_in[0][119] ) );
  NAND U7981 ( .A(init), .B(round_reg[11]), .Z(n2902) );
  NAND U7982 ( .A(n2773), .B(in[11]), .Z(n2901) );
  NAND U7983 ( .A(n2902), .B(n2901), .Z(\round_in[0][11] ) );
  AND U7984 ( .A(round_reg[1200]), .B(init), .Z(\round_in[0][1200] ) );
  AND U7985 ( .A(round_reg[1201]), .B(init), .Z(\round_in[0][1201] ) );
  AND U7986 ( .A(round_reg[1202]), .B(init), .Z(\round_in[0][1202] ) );
  AND U7987 ( .A(round_reg[1203]), .B(init), .Z(\round_in[0][1203] ) );
  AND U7988 ( .A(round_reg[1204]), .B(init), .Z(\round_in[0][1204] ) );
  AND U7989 ( .A(round_reg[1205]), .B(init), .Z(\round_in[0][1205] ) );
  AND U7990 ( .A(round_reg[1206]), .B(init), .Z(\round_in[0][1206] ) );
  AND U7991 ( .A(round_reg[1207]), .B(init), .Z(\round_in[0][1207] ) );
  AND U7992 ( .A(round_reg[1208]), .B(init), .Z(\round_in[0][1208] ) );
  AND U7993 ( .A(round_reg[1209]), .B(init), .Z(\round_in[0][1209] ) );
  NAND U7994 ( .A(init), .B(round_reg[120]), .Z(n2904) );
  NAND U7995 ( .A(n2773), .B(in[120]), .Z(n2903) );
  NAND U7996 ( .A(n2904), .B(n2903), .Z(\round_in[0][120] ) );
  AND U7997 ( .A(round_reg[1210]), .B(init), .Z(\round_in[0][1210] ) );
  AND U7998 ( .A(round_reg[1211]), .B(init), .Z(\round_in[0][1211] ) );
  AND U7999 ( .A(round_reg[1212]), .B(init), .Z(\round_in[0][1212] ) );
  AND U8000 ( .A(round_reg[1213]), .B(init), .Z(\round_in[0][1213] ) );
  AND U8001 ( .A(round_reg[1214]), .B(init), .Z(\round_in[0][1214] ) );
  AND U8002 ( .A(round_reg[1215]), .B(init), .Z(\round_in[0][1215] ) );
  AND U8003 ( .A(round_reg[1216]), .B(init), .Z(\round_in[0][1216] ) );
  AND U8004 ( .A(round_reg[1217]), .B(init), .Z(\round_in[0][1217] ) );
  AND U8005 ( .A(round_reg[1218]), .B(init), .Z(\round_in[0][1218] ) );
  AND U8006 ( .A(round_reg[1219]), .B(init), .Z(\round_in[0][1219] ) );
  NAND U8007 ( .A(init), .B(round_reg[121]), .Z(n2906) );
  NAND U8008 ( .A(n2773), .B(in[121]), .Z(n2905) );
  NAND U8009 ( .A(n2906), .B(n2905), .Z(\round_in[0][121] ) );
  AND U8010 ( .A(round_reg[1220]), .B(init), .Z(\round_in[0][1220] ) );
  AND U8011 ( .A(round_reg[1221]), .B(init), .Z(\round_in[0][1221] ) );
  AND U8012 ( .A(round_reg[1222]), .B(init), .Z(\round_in[0][1222] ) );
  AND U8013 ( .A(round_reg[1223]), .B(init), .Z(\round_in[0][1223] ) );
  AND U8014 ( .A(round_reg[1224]), .B(init), .Z(\round_in[0][1224] ) );
  AND U8015 ( .A(round_reg[1225]), .B(init), .Z(\round_in[0][1225] ) );
  AND U8016 ( .A(round_reg[1226]), .B(init), .Z(\round_in[0][1226] ) );
  AND U8017 ( .A(round_reg[1227]), .B(init), .Z(\round_in[0][1227] ) );
  AND U8018 ( .A(round_reg[1228]), .B(init), .Z(\round_in[0][1228] ) );
  AND U8019 ( .A(round_reg[1229]), .B(init), .Z(\round_in[0][1229] ) );
  NAND U8020 ( .A(init), .B(round_reg[122]), .Z(n2908) );
  NAND U8021 ( .A(n2773), .B(in[122]), .Z(n2907) );
  NAND U8022 ( .A(n2908), .B(n2907), .Z(\round_in[0][122] ) );
  AND U8023 ( .A(round_reg[1230]), .B(init), .Z(\round_in[0][1230] ) );
  AND U8024 ( .A(round_reg[1231]), .B(init), .Z(\round_in[0][1231] ) );
  AND U8025 ( .A(round_reg[1232]), .B(init), .Z(\round_in[0][1232] ) );
  AND U8026 ( .A(round_reg[1233]), .B(init), .Z(\round_in[0][1233] ) );
  AND U8027 ( .A(round_reg[1234]), .B(init), .Z(\round_in[0][1234] ) );
  AND U8028 ( .A(round_reg[1235]), .B(init), .Z(\round_in[0][1235] ) );
  AND U8029 ( .A(round_reg[1236]), .B(init), .Z(\round_in[0][1236] ) );
  AND U8030 ( .A(round_reg[1237]), .B(init), .Z(\round_in[0][1237] ) );
  AND U8031 ( .A(round_reg[1238]), .B(init), .Z(\round_in[0][1238] ) );
  AND U8032 ( .A(round_reg[1239]), .B(init), .Z(\round_in[0][1239] ) );
  NAND U8033 ( .A(init), .B(round_reg[123]), .Z(n2910) );
  NAND U8034 ( .A(n2774), .B(in[123]), .Z(n2909) );
  NAND U8035 ( .A(n2910), .B(n2909), .Z(\round_in[0][123] ) );
  AND U8036 ( .A(round_reg[1240]), .B(init), .Z(\round_in[0][1240] ) );
  AND U8037 ( .A(round_reg[1241]), .B(init), .Z(\round_in[0][1241] ) );
  AND U8038 ( .A(round_reg[1242]), .B(init), .Z(\round_in[0][1242] ) );
  AND U8039 ( .A(round_reg[1243]), .B(init), .Z(\round_in[0][1243] ) );
  AND U8040 ( .A(round_reg[1244]), .B(init), .Z(\round_in[0][1244] ) );
  AND U8041 ( .A(round_reg[1245]), .B(init), .Z(\round_in[0][1245] ) );
  AND U8042 ( .A(round_reg[1246]), .B(init), .Z(\round_in[0][1246] ) );
  AND U8043 ( .A(round_reg[1247]), .B(init), .Z(\round_in[0][1247] ) );
  AND U8044 ( .A(round_reg[1248]), .B(init), .Z(\round_in[0][1248] ) );
  AND U8045 ( .A(round_reg[1249]), .B(init), .Z(\round_in[0][1249] ) );
  NAND U8046 ( .A(init), .B(round_reg[124]), .Z(n2912) );
  NAND U8047 ( .A(n2774), .B(in[124]), .Z(n2911) );
  NAND U8048 ( .A(n2912), .B(n2911), .Z(\round_in[0][124] ) );
  AND U8049 ( .A(round_reg[1250]), .B(init), .Z(\round_in[0][1250] ) );
  AND U8050 ( .A(round_reg[1251]), .B(init), .Z(\round_in[0][1251] ) );
  AND U8051 ( .A(round_reg[1252]), .B(init), .Z(\round_in[0][1252] ) );
  AND U8052 ( .A(round_reg[1253]), .B(init), .Z(\round_in[0][1253] ) );
  AND U8053 ( .A(round_reg[1254]), .B(init), .Z(\round_in[0][1254] ) );
  AND U8054 ( .A(round_reg[1255]), .B(init), .Z(\round_in[0][1255] ) );
  AND U8055 ( .A(round_reg[1256]), .B(init), .Z(\round_in[0][1256] ) );
  AND U8056 ( .A(round_reg[1257]), .B(init), .Z(\round_in[0][1257] ) );
  AND U8057 ( .A(round_reg[1258]), .B(init), .Z(\round_in[0][1258] ) );
  AND U8058 ( .A(round_reg[1259]), .B(init), .Z(\round_in[0][1259] ) );
  NAND U8059 ( .A(init), .B(round_reg[125]), .Z(n2914) );
  NAND U8060 ( .A(n2774), .B(in[125]), .Z(n2913) );
  NAND U8061 ( .A(n2914), .B(n2913), .Z(\round_in[0][125] ) );
  AND U8062 ( .A(round_reg[1260]), .B(init), .Z(\round_in[0][1260] ) );
  AND U8063 ( .A(round_reg[1261]), .B(init), .Z(\round_in[0][1261] ) );
  AND U8064 ( .A(round_reg[1262]), .B(init), .Z(\round_in[0][1262] ) );
  AND U8065 ( .A(round_reg[1263]), .B(init), .Z(\round_in[0][1263] ) );
  AND U8066 ( .A(round_reg[1264]), .B(init), .Z(\round_in[0][1264] ) );
  AND U8067 ( .A(round_reg[1265]), .B(init), .Z(\round_in[0][1265] ) );
  AND U8068 ( .A(round_reg[1266]), .B(init), .Z(\round_in[0][1266] ) );
  AND U8069 ( .A(round_reg[1267]), .B(init), .Z(\round_in[0][1267] ) );
  AND U8070 ( .A(round_reg[1268]), .B(init), .Z(\round_in[0][1268] ) );
  AND U8071 ( .A(round_reg[1269]), .B(init), .Z(\round_in[0][1269] ) );
  NAND U8072 ( .A(init), .B(round_reg[126]), .Z(n2916) );
  NAND U8073 ( .A(n2774), .B(in[126]), .Z(n2915) );
  NAND U8074 ( .A(n2916), .B(n2915), .Z(\round_in[0][126] ) );
  AND U8075 ( .A(round_reg[1270]), .B(init), .Z(\round_in[0][1270] ) );
  AND U8076 ( .A(round_reg[1271]), .B(init), .Z(\round_in[0][1271] ) );
  AND U8077 ( .A(round_reg[1272]), .B(init), .Z(\round_in[0][1272] ) );
  AND U8078 ( .A(round_reg[1273]), .B(init), .Z(\round_in[0][1273] ) );
  AND U8079 ( .A(round_reg[1274]), .B(init), .Z(\round_in[0][1274] ) );
  AND U8080 ( .A(round_reg[1275]), .B(init), .Z(\round_in[0][1275] ) );
  AND U8081 ( .A(round_reg[1276]), .B(init), .Z(\round_in[0][1276] ) );
  AND U8082 ( .A(round_reg[1277]), .B(init), .Z(\round_in[0][1277] ) );
  AND U8083 ( .A(round_reg[1278]), .B(init), .Z(\round_in[0][1278] ) );
  AND U8084 ( .A(round_reg[1279]), .B(init), .Z(\round_in[0][1279] ) );
  NAND U8085 ( .A(init), .B(round_reg[127]), .Z(n2918) );
  NAND U8086 ( .A(n2774), .B(in[127]), .Z(n2917) );
  NAND U8087 ( .A(n2918), .B(n2917), .Z(\round_in[0][127] ) );
  AND U8088 ( .A(round_reg[1280]), .B(init), .Z(\round_in[0][1280] ) );
  AND U8089 ( .A(round_reg[1281]), .B(init), .Z(\round_in[0][1281] ) );
  AND U8090 ( .A(round_reg[1282]), .B(init), .Z(\round_in[0][1282] ) );
  AND U8091 ( .A(round_reg[1283]), .B(init), .Z(\round_in[0][1283] ) );
  AND U8092 ( .A(round_reg[1284]), .B(init), .Z(\round_in[0][1284] ) );
  AND U8093 ( .A(round_reg[1285]), .B(init), .Z(\round_in[0][1285] ) );
  AND U8094 ( .A(round_reg[1286]), .B(init), .Z(\round_in[0][1286] ) );
  AND U8095 ( .A(round_reg[1287]), .B(init), .Z(\round_in[0][1287] ) );
  AND U8096 ( .A(round_reg[1288]), .B(init), .Z(\round_in[0][1288] ) );
  AND U8097 ( .A(round_reg[1289]), .B(init), .Z(\round_in[0][1289] ) );
  NAND U8098 ( .A(init), .B(round_reg[128]), .Z(n2920) );
  NAND U8099 ( .A(n2774), .B(in[128]), .Z(n2919) );
  NAND U8100 ( .A(n2920), .B(n2919), .Z(\round_in[0][128] ) );
  AND U8101 ( .A(round_reg[1290]), .B(init), .Z(\round_in[0][1290] ) );
  AND U8102 ( .A(round_reg[1291]), .B(init), .Z(\round_in[0][1291] ) );
  AND U8103 ( .A(round_reg[1292]), .B(init), .Z(\round_in[0][1292] ) );
  AND U8104 ( .A(round_reg[1293]), .B(init), .Z(\round_in[0][1293] ) );
  AND U8105 ( .A(round_reg[1294]), .B(init), .Z(\round_in[0][1294] ) );
  AND U8106 ( .A(round_reg[1295]), .B(init), .Z(\round_in[0][1295] ) );
  AND U8107 ( .A(round_reg[1296]), .B(init), .Z(\round_in[0][1296] ) );
  AND U8108 ( .A(round_reg[1297]), .B(init), .Z(\round_in[0][1297] ) );
  AND U8109 ( .A(round_reg[1298]), .B(init), .Z(\round_in[0][1298] ) );
  AND U8110 ( .A(round_reg[1299]), .B(init), .Z(\round_in[0][1299] ) );
  NAND U8111 ( .A(init), .B(round_reg[129]), .Z(n2922) );
  NAND U8112 ( .A(n2774), .B(in[129]), .Z(n2921) );
  NAND U8113 ( .A(n2922), .B(n2921), .Z(\round_in[0][129] ) );
  NAND U8114 ( .A(init), .B(round_reg[12]), .Z(n2924) );
  NAND U8115 ( .A(n2775), .B(in[12]), .Z(n2923) );
  NAND U8116 ( .A(n2924), .B(n2923), .Z(\round_in[0][12] ) );
  AND U8117 ( .A(round_reg[1300]), .B(init), .Z(\round_in[0][1300] ) );
  AND U8118 ( .A(round_reg[1301]), .B(init), .Z(\round_in[0][1301] ) );
  AND U8119 ( .A(round_reg[1302]), .B(init), .Z(\round_in[0][1302] ) );
  AND U8120 ( .A(round_reg[1303]), .B(init), .Z(\round_in[0][1303] ) );
  AND U8121 ( .A(round_reg[1304]), .B(init), .Z(\round_in[0][1304] ) );
  AND U8122 ( .A(round_reg[1305]), .B(init), .Z(\round_in[0][1305] ) );
  AND U8123 ( .A(round_reg[1306]), .B(init), .Z(\round_in[0][1306] ) );
  AND U8124 ( .A(round_reg[1307]), .B(init), .Z(\round_in[0][1307] ) );
  AND U8125 ( .A(round_reg[1308]), .B(init), .Z(\round_in[0][1308] ) );
  AND U8126 ( .A(round_reg[1309]), .B(init), .Z(\round_in[0][1309] ) );
  NAND U8127 ( .A(init), .B(round_reg[130]), .Z(n2926) );
  NAND U8128 ( .A(n2775), .B(in[130]), .Z(n2925) );
  NAND U8129 ( .A(n2926), .B(n2925), .Z(\round_in[0][130] ) );
  AND U8130 ( .A(round_reg[1310]), .B(init), .Z(\round_in[0][1310] ) );
  AND U8131 ( .A(round_reg[1311]), .B(init), .Z(\round_in[0][1311] ) );
  AND U8132 ( .A(round_reg[1312]), .B(init), .Z(\round_in[0][1312] ) );
  AND U8133 ( .A(round_reg[1313]), .B(init), .Z(\round_in[0][1313] ) );
  AND U8134 ( .A(round_reg[1314]), .B(init), .Z(\round_in[0][1314] ) );
  AND U8135 ( .A(round_reg[1315]), .B(init), .Z(\round_in[0][1315] ) );
  AND U8136 ( .A(round_reg[1316]), .B(init), .Z(\round_in[0][1316] ) );
  AND U8137 ( .A(round_reg[1317]), .B(init), .Z(\round_in[0][1317] ) );
  AND U8138 ( .A(round_reg[1318]), .B(init), .Z(\round_in[0][1318] ) );
  AND U8139 ( .A(round_reg[1319]), .B(init), .Z(\round_in[0][1319] ) );
  NAND U8140 ( .A(init), .B(round_reg[131]), .Z(n2928) );
  NAND U8141 ( .A(n2775), .B(in[131]), .Z(n2927) );
  NAND U8142 ( .A(n2928), .B(n2927), .Z(\round_in[0][131] ) );
  AND U8143 ( .A(round_reg[1320]), .B(init), .Z(\round_in[0][1320] ) );
  AND U8144 ( .A(round_reg[1321]), .B(init), .Z(\round_in[0][1321] ) );
  AND U8145 ( .A(round_reg[1322]), .B(init), .Z(\round_in[0][1322] ) );
  AND U8146 ( .A(round_reg[1323]), .B(init), .Z(\round_in[0][1323] ) );
  AND U8147 ( .A(round_reg[1324]), .B(init), .Z(\round_in[0][1324] ) );
  AND U8148 ( .A(round_reg[1325]), .B(init), .Z(\round_in[0][1325] ) );
  AND U8149 ( .A(round_reg[1326]), .B(init), .Z(\round_in[0][1326] ) );
  AND U8150 ( .A(round_reg[1327]), .B(init), .Z(\round_in[0][1327] ) );
  AND U8151 ( .A(round_reg[1328]), .B(init), .Z(\round_in[0][1328] ) );
  AND U8152 ( .A(round_reg[1329]), .B(init), .Z(\round_in[0][1329] ) );
  NAND U8153 ( .A(init), .B(round_reg[132]), .Z(n2930) );
  NAND U8154 ( .A(n2775), .B(in[132]), .Z(n2929) );
  NAND U8155 ( .A(n2930), .B(n2929), .Z(\round_in[0][132] ) );
  AND U8156 ( .A(round_reg[1330]), .B(init), .Z(\round_in[0][1330] ) );
  AND U8157 ( .A(round_reg[1331]), .B(init), .Z(\round_in[0][1331] ) );
  AND U8158 ( .A(round_reg[1332]), .B(init), .Z(\round_in[0][1332] ) );
  AND U8159 ( .A(round_reg[1333]), .B(init), .Z(\round_in[0][1333] ) );
  AND U8160 ( .A(round_reg[1334]), .B(init), .Z(\round_in[0][1334] ) );
  AND U8161 ( .A(round_reg[1335]), .B(init), .Z(\round_in[0][1335] ) );
  AND U8162 ( .A(round_reg[1336]), .B(init), .Z(\round_in[0][1336] ) );
  AND U8163 ( .A(round_reg[1337]), .B(init), .Z(\round_in[0][1337] ) );
  AND U8164 ( .A(round_reg[1338]), .B(init), .Z(\round_in[0][1338] ) );
  AND U8165 ( .A(round_reg[1339]), .B(init), .Z(\round_in[0][1339] ) );
  NAND U8166 ( .A(init), .B(round_reg[133]), .Z(n2932) );
  NAND U8167 ( .A(n2775), .B(in[133]), .Z(n2931) );
  NAND U8168 ( .A(n2932), .B(n2931), .Z(\round_in[0][133] ) );
  AND U8169 ( .A(round_reg[1340]), .B(init), .Z(\round_in[0][1340] ) );
  AND U8170 ( .A(round_reg[1341]), .B(init), .Z(\round_in[0][1341] ) );
  AND U8171 ( .A(round_reg[1342]), .B(init), .Z(\round_in[0][1342] ) );
  AND U8172 ( .A(round_reg[1343]), .B(init), .Z(\round_in[0][1343] ) );
  AND U8173 ( .A(round_reg[1344]), .B(init), .Z(\round_in[0][1344] ) );
  AND U8174 ( .A(round_reg[1345]), .B(init), .Z(\round_in[0][1345] ) );
  AND U8175 ( .A(round_reg[1346]), .B(init), .Z(\round_in[0][1346] ) );
  AND U8176 ( .A(round_reg[1347]), .B(init), .Z(\round_in[0][1347] ) );
  AND U8177 ( .A(round_reg[1348]), .B(init), .Z(\round_in[0][1348] ) );
  AND U8178 ( .A(round_reg[1349]), .B(init), .Z(\round_in[0][1349] ) );
  NAND U8179 ( .A(init), .B(round_reg[134]), .Z(n2934) );
  NAND U8180 ( .A(n2775), .B(in[134]), .Z(n2933) );
  NAND U8181 ( .A(n2934), .B(n2933), .Z(\round_in[0][134] ) );
  AND U8182 ( .A(round_reg[1350]), .B(init), .Z(\round_in[0][1350] ) );
  AND U8183 ( .A(round_reg[1351]), .B(init), .Z(\round_in[0][1351] ) );
  AND U8184 ( .A(round_reg[1352]), .B(init), .Z(\round_in[0][1352] ) );
  AND U8185 ( .A(round_reg[1353]), .B(init), .Z(\round_in[0][1353] ) );
  AND U8186 ( .A(round_reg[1354]), .B(init), .Z(\round_in[0][1354] ) );
  AND U8187 ( .A(round_reg[1355]), .B(init), .Z(\round_in[0][1355] ) );
  AND U8188 ( .A(round_reg[1356]), .B(init), .Z(\round_in[0][1356] ) );
  AND U8189 ( .A(round_reg[1357]), .B(init), .Z(\round_in[0][1357] ) );
  AND U8190 ( .A(round_reg[1358]), .B(init), .Z(\round_in[0][1358] ) );
  AND U8191 ( .A(round_reg[1359]), .B(init), .Z(\round_in[0][1359] ) );
  NAND U8192 ( .A(init), .B(round_reg[135]), .Z(n2936) );
  NAND U8193 ( .A(n2775), .B(in[135]), .Z(n2935) );
  NAND U8194 ( .A(n2936), .B(n2935), .Z(\round_in[0][135] ) );
  AND U8195 ( .A(round_reg[1360]), .B(init), .Z(\round_in[0][1360] ) );
  AND U8196 ( .A(round_reg[1361]), .B(init), .Z(\round_in[0][1361] ) );
  AND U8197 ( .A(round_reg[1362]), .B(init), .Z(\round_in[0][1362] ) );
  AND U8198 ( .A(round_reg[1363]), .B(init), .Z(\round_in[0][1363] ) );
  AND U8199 ( .A(round_reg[1364]), .B(init), .Z(\round_in[0][1364] ) );
  AND U8200 ( .A(round_reg[1365]), .B(init), .Z(\round_in[0][1365] ) );
  AND U8201 ( .A(round_reg[1366]), .B(init), .Z(\round_in[0][1366] ) );
  AND U8202 ( .A(round_reg[1367]), .B(init), .Z(\round_in[0][1367] ) );
  AND U8203 ( .A(round_reg[1368]), .B(init), .Z(\round_in[0][1368] ) );
  AND U8204 ( .A(round_reg[1369]), .B(init), .Z(\round_in[0][1369] ) );
  NAND U8205 ( .A(init), .B(round_reg[136]), .Z(n2938) );
  NAND U8206 ( .A(n2776), .B(in[136]), .Z(n2937) );
  NAND U8207 ( .A(n2938), .B(n2937), .Z(\round_in[0][136] ) );
  AND U8208 ( .A(round_reg[1370]), .B(init), .Z(\round_in[0][1370] ) );
  AND U8209 ( .A(round_reg[1371]), .B(init), .Z(\round_in[0][1371] ) );
  AND U8210 ( .A(round_reg[1372]), .B(init), .Z(\round_in[0][1372] ) );
  AND U8211 ( .A(round_reg[1373]), .B(init), .Z(\round_in[0][1373] ) );
  AND U8212 ( .A(round_reg[1374]), .B(init), .Z(\round_in[0][1374] ) );
  AND U8213 ( .A(round_reg[1375]), .B(init), .Z(\round_in[0][1375] ) );
  AND U8214 ( .A(round_reg[1376]), .B(init), .Z(\round_in[0][1376] ) );
  AND U8215 ( .A(round_reg[1377]), .B(init), .Z(\round_in[0][1377] ) );
  AND U8216 ( .A(round_reg[1378]), .B(init), .Z(\round_in[0][1378] ) );
  AND U8217 ( .A(round_reg[1379]), .B(init), .Z(\round_in[0][1379] ) );
  NAND U8218 ( .A(init), .B(round_reg[137]), .Z(n2940) );
  NAND U8219 ( .A(n2776), .B(in[137]), .Z(n2939) );
  NAND U8220 ( .A(n2940), .B(n2939), .Z(\round_in[0][137] ) );
  AND U8221 ( .A(round_reg[1380]), .B(init), .Z(\round_in[0][1380] ) );
  AND U8222 ( .A(round_reg[1381]), .B(init), .Z(\round_in[0][1381] ) );
  AND U8223 ( .A(round_reg[1382]), .B(init), .Z(\round_in[0][1382] ) );
  AND U8224 ( .A(round_reg[1383]), .B(init), .Z(\round_in[0][1383] ) );
  AND U8225 ( .A(round_reg[1384]), .B(init), .Z(\round_in[0][1384] ) );
  AND U8226 ( .A(round_reg[1385]), .B(init), .Z(\round_in[0][1385] ) );
  AND U8227 ( .A(round_reg[1386]), .B(init), .Z(\round_in[0][1386] ) );
  AND U8228 ( .A(round_reg[1387]), .B(init), .Z(\round_in[0][1387] ) );
  AND U8229 ( .A(round_reg[1388]), .B(init), .Z(\round_in[0][1388] ) );
  AND U8230 ( .A(round_reg[1389]), .B(init), .Z(\round_in[0][1389] ) );
  NAND U8231 ( .A(init), .B(round_reg[138]), .Z(n2942) );
  NAND U8232 ( .A(n2776), .B(in[138]), .Z(n2941) );
  NAND U8233 ( .A(n2942), .B(n2941), .Z(\round_in[0][138] ) );
  AND U8234 ( .A(round_reg[1390]), .B(init), .Z(\round_in[0][1390] ) );
  AND U8235 ( .A(round_reg[1391]), .B(init), .Z(\round_in[0][1391] ) );
  AND U8236 ( .A(round_reg[1392]), .B(init), .Z(\round_in[0][1392] ) );
  AND U8237 ( .A(round_reg[1393]), .B(init), .Z(\round_in[0][1393] ) );
  AND U8238 ( .A(round_reg[1394]), .B(init), .Z(\round_in[0][1394] ) );
  AND U8239 ( .A(round_reg[1395]), .B(init), .Z(\round_in[0][1395] ) );
  AND U8240 ( .A(round_reg[1396]), .B(init), .Z(\round_in[0][1396] ) );
  AND U8241 ( .A(round_reg[1397]), .B(init), .Z(\round_in[0][1397] ) );
  AND U8242 ( .A(round_reg[1398]), .B(init), .Z(\round_in[0][1398] ) );
  AND U8243 ( .A(round_reg[1399]), .B(init), .Z(\round_in[0][1399] ) );
  NAND U8244 ( .A(init), .B(round_reg[139]), .Z(n2944) );
  NAND U8245 ( .A(n2776), .B(in[139]), .Z(n2943) );
  NAND U8246 ( .A(n2944), .B(n2943), .Z(\round_in[0][139] ) );
  NAND U8247 ( .A(init), .B(round_reg[13]), .Z(n2946) );
  NAND U8248 ( .A(n2776), .B(in[13]), .Z(n2945) );
  NAND U8249 ( .A(n2946), .B(n2945), .Z(\round_in[0][13] ) );
  AND U8250 ( .A(round_reg[1400]), .B(init), .Z(\round_in[0][1400] ) );
  AND U8251 ( .A(round_reg[1401]), .B(init), .Z(\round_in[0][1401] ) );
  AND U8252 ( .A(round_reg[1402]), .B(init), .Z(\round_in[0][1402] ) );
  AND U8253 ( .A(round_reg[1403]), .B(init), .Z(\round_in[0][1403] ) );
  AND U8254 ( .A(round_reg[1404]), .B(init), .Z(\round_in[0][1404] ) );
  AND U8255 ( .A(round_reg[1405]), .B(init), .Z(\round_in[0][1405] ) );
  AND U8256 ( .A(round_reg[1406]), .B(init), .Z(\round_in[0][1406] ) );
  AND U8257 ( .A(round_reg[1407]), .B(init), .Z(\round_in[0][1407] ) );
  AND U8258 ( .A(round_reg[1408]), .B(init), .Z(\round_in[0][1408] ) );
  AND U8259 ( .A(round_reg[1409]), .B(init), .Z(\round_in[0][1409] ) );
  NAND U8260 ( .A(init), .B(round_reg[140]), .Z(n2948) );
  NAND U8261 ( .A(n2776), .B(in[140]), .Z(n2947) );
  NAND U8262 ( .A(n2948), .B(n2947), .Z(\round_in[0][140] ) );
  AND U8263 ( .A(round_reg[1410]), .B(init), .Z(\round_in[0][1410] ) );
  AND U8264 ( .A(round_reg[1411]), .B(init), .Z(\round_in[0][1411] ) );
  AND U8265 ( .A(round_reg[1412]), .B(init), .Z(\round_in[0][1412] ) );
  AND U8266 ( .A(round_reg[1413]), .B(init), .Z(\round_in[0][1413] ) );
  AND U8267 ( .A(round_reg[1414]), .B(init), .Z(\round_in[0][1414] ) );
  AND U8268 ( .A(round_reg[1415]), .B(init), .Z(\round_in[0][1415] ) );
  AND U8269 ( .A(round_reg[1416]), .B(init), .Z(\round_in[0][1416] ) );
  AND U8270 ( .A(round_reg[1417]), .B(init), .Z(\round_in[0][1417] ) );
  AND U8271 ( .A(round_reg[1418]), .B(init), .Z(\round_in[0][1418] ) );
  AND U8272 ( .A(round_reg[1419]), .B(init), .Z(\round_in[0][1419] ) );
  NAND U8273 ( .A(init), .B(round_reg[141]), .Z(n2950) );
  NAND U8274 ( .A(n2776), .B(in[141]), .Z(n2949) );
  NAND U8275 ( .A(n2950), .B(n2949), .Z(\round_in[0][141] ) );
  AND U8276 ( .A(round_reg[1420]), .B(init), .Z(\round_in[0][1420] ) );
  AND U8277 ( .A(round_reg[1421]), .B(init), .Z(\round_in[0][1421] ) );
  AND U8278 ( .A(round_reg[1422]), .B(init), .Z(\round_in[0][1422] ) );
  AND U8279 ( .A(round_reg[1423]), .B(init), .Z(\round_in[0][1423] ) );
  AND U8280 ( .A(round_reg[1424]), .B(init), .Z(\round_in[0][1424] ) );
  AND U8281 ( .A(round_reg[1425]), .B(init), .Z(\round_in[0][1425] ) );
  AND U8282 ( .A(round_reg[1426]), .B(init), .Z(\round_in[0][1426] ) );
  AND U8283 ( .A(round_reg[1427]), .B(init), .Z(\round_in[0][1427] ) );
  AND U8284 ( .A(round_reg[1428]), .B(init), .Z(\round_in[0][1428] ) );
  AND U8285 ( .A(round_reg[1429]), .B(init), .Z(\round_in[0][1429] ) );
  NAND U8286 ( .A(init), .B(round_reg[142]), .Z(n2952) );
  NAND U8287 ( .A(n2777), .B(in[142]), .Z(n2951) );
  NAND U8288 ( .A(n2952), .B(n2951), .Z(\round_in[0][142] ) );
  AND U8289 ( .A(round_reg[1430]), .B(init), .Z(\round_in[0][1430] ) );
  AND U8290 ( .A(round_reg[1431]), .B(init), .Z(\round_in[0][1431] ) );
  AND U8291 ( .A(round_reg[1432]), .B(init), .Z(\round_in[0][1432] ) );
  AND U8292 ( .A(round_reg[1433]), .B(init), .Z(\round_in[0][1433] ) );
  AND U8293 ( .A(round_reg[1434]), .B(init), .Z(\round_in[0][1434] ) );
  AND U8294 ( .A(round_reg[1435]), .B(init), .Z(\round_in[0][1435] ) );
  AND U8295 ( .A(round_reg[1436]), .B(init), .Z(\round_in[0][1436] ) );
  AND U8296 ( .A(round_reg[1437]), .B(init), .Z(\round_in[0][1437] ) );
  AND U8297 ( .A(round_reg[1438]), .B(init), .Z(\round_in[0][1438] ) );
  AND U8298 ( .A(round_reg[1439]), .B(init), .Z(\round_in[0][1439] ) );
  NAND U8299 ( .A(init), .B(round_reg[143]), .Z(n2954) );
  NAND U8300 ( .A(n2777), .B(in[143]), .Z(n2953) );
  NAND U8301 ( .A(n2954), .B(n2953), .Z(\round_in[0][143] ) );
  AND U8302 ( .A(round_reg[1440]), .B(init), .Z(\round_in[0][1440] ) );
  AND U8303 ( .A(round_reg[1441]), .B(init), .Z(\round_in[0][1441] ) );
  AND U8304 ( .A(round_reg[1442]), .B(init), .Z(\round_in[0][1442] ) );
  AND U8305 ( .A(round_reg[1443]), .B(init), .Z(\round_in[0][1443] ) );
  AND U8306 ( .A(round_reg[1444]), .B(init), .Z(\round_in[0][1444] ) );
  AND U8307 ( .A(round_reg[1445]), .B(init), .Z(\round_in[0][1445] ) );
  AND U8308 ( .A(round_reg[1446]), .B(init), .Z(\round_in[0][1446] ) );
  AND U8309 ( .A(round_reg[1447]), .B(init), .Z(\round_in[0][1447] ) );
  AND U8310 ( .A(round_reg[1448]), .B(init), .Z(\round_in[0][1448] ) );
  AND U8311 ( .A(round_reg[1449]), .B(init), .Z(\round_in[0][1449] ) );
  NAND U8312 ( .A(init), .B(round_reg[144]), .Z(n2956) );
  NAND U8313 ( .A(n2777), .B(in[144]), .Z(n2955) );
  NAND U8314 ( .A(n2956), .B(n2955), .Z(\round_in[0][144] ) );
  AND U8315 ( .A(round_reg[1450]), .B(init), .Z(\round_in[0][1450] ) );
  AND U8316 ( .A(round_reg[1451]), .B(init), .Z(\round_in[0][1451] ) );
  AND U8317 ( .A(round_reg[1452]), .B(init), .Z(\round_in[0][1452] ) );
  AND U8318 ( .A(round_reg[1453]), .B(init), .Z(\round_in[0][1453] ) );
  AND U8319 ( .A(round_reg[1454]), .B(init), .Z(\round_in[0][1454] ) );
  AND U8320 ( .A(round_reg[1455]), .B(init), .Z(\round_in[0][1455] ) );
  AND U8321 ( .A(round_reg[1456]), .B(init), .Z(\round_in[0][1456] ) );
  AND U8322 ( .A(round_reg[1457]), .B(init), .Z(\round_in[0][1457] ) );
  AND U8323 ( .A(round_reg[1458]), .B(init), .Z(\round_in[0][1458] ) );
  AND U8324 ( .A(round_reg[1459]), .B(init), .Z(\round_in[0][1459] ) );
  NAND U8325 ( .A(init), .B(round_reg[145]), .Z(n2958) );
  NAND U8326 ( .A(n2777), .B(in[145]), .Z(n2957) );
  NAND U8327 ( .A(n2958), .B(n2957), .Z(\round_in[0][145] ) );
  AND U8328 ( .A(round_reg[1460]), .B(init), .Z(\round_in[0][1460] ) );
  AND U8329 ( .A(round_reg[1461]), .B(init), .Z(\round_in[0][1461] ) );
  AND U8330 ( .A(round_reg[1462]), .B(init), .Z(\round_in[0][1462] ) );
  AND U8331 ( .A(round_reg[1463]), .B(init), .Z(\round_in[0][1463] ) );
  AND U8332 ( .A(round_reg[1464]), .B(init), .Z(\round_in[0][1464] ) );
  AND U8333 ( .A(round_reg[1465]), .B(init), .Z(\round_in[0][1465] ) );
  AND U8334 ( .A(round_reg[1466]), .B(init), .Z(\round_in[0][1466] ) );
  AND U8335 ( .A(round_reg[1467]), .B(init), .Z(\round_in[0][1467] ) );
  AND U8336 ( .A(round_reg[1468]), .B(init), .Z(\round_in[0][1468] ) );
  AND U8337 ( .A(round_reg[1469]), .B(init), .Z(\round_in[0][1469] ) );
  NAND U8338 ( .A(init), .B(round_reg[146]), .Z(n2960) );
  NAND U8339 ( .A(n2777), .B(in[146]), .Z(n2959) );
  NAND U8340 ( .A(n2960), .B(n2959), .Z(\round_in[0][146] ) );
  AND U8341 ( .A(round_reg[1470]), .B(init), .Z(\round_in[0][1470] ) );
  AND U8342 ( .A(round_reg[1471]), .B(init), .Z(\round_in[0][1471] ) );
  AND U8343 ( .A(round_reg[1472]), .B(init), .Z(\round_in[0][1472] ) );
  AND U8344 ( .A(round_reg[1473]), .B(init), .Z(\round_in[0][1473] ) );
  AND U8345 ( .A(round_reg[1474]), .B(init), .Z(\round_in[0][1474] ) );
  AND U8346 ( .A(round_reg[1475]), .B(init), .Z(\round_in[0][1475] ) );
  AND U8347 ( .A(round_reg[1476]), .B(init), .Z(\round_in[0][1476] ) );
  AND U8348 ( .A(round_reg[1477]), .B(init), .Z(\round_in[0][1477] ) );
  AND U8349 ( .A(round_reg[1478]), .B(init), .Z(\round_in[0][1478] ) );
  AND U8350 ( .A(round_reg[1479]), .B(init), .Z(\round_in[0][1479] ) );
  NAND U8351 ( .A(init), .B(round_reg[147]), .Z(n2962) );
  NAND U8352 ( .A(n2777), .B(in[147]), .Z(n2961) );
  NAND U8353 ( .A(n2962), .B(n2961), .Z(\round_in[0][147] ) );
  AND U8354 ( .A(round_reg[1480]), .B(init), .Z(\round_in[0][1480] ) );
  AND U8355 ( .A(round_reg[1481]), .B(init), .Z(\round_in[0][1481] ) );
  AND U8356 ( .A(round_reg[1482]), .B(init), .Z(\round_in[0][1482] ) );
  AND U8357 ( .A(round_reg[1483]), .B(init), .Z(\round_in[0][1483] ) );
  AND U8358 ( .A(round_reg[1484]), .B(init), .Z(\round_in[0][1484] ) );
  AND U8359 ( .A(round_reg[1485]), .B(init), .Z(\round_in[0][1485] ) );
  AND U8360 ( .A(round_reg[1486]), .B(init), .Z(\round_in[0][1486] ) );
  AND U8361 ( .A(round_reg[1487]), .B(init), .Z(\round_in[0][1487] ) );
  AND U8362 ( .A(round_reg[1488]), .B(init), .Z(\round_in[0][1488] ) );
  AND U8363 ( .A(round_reg[1489]), .B(init), .Z(\round_in[0][1489] ) );
  NAND U8364 ( .A(init), .B(round_reg[148]), .Z(n2964) );
  NAND U8365 ( .A(n2777), .B(in[148]), .Z(n2963) );
  NAND U8366 ( .A(n2964), .B(n2963), .Z(\round_in[0][148] ) );
  AND U8367 ( .A(round_reg[1490]), .B(init), .Z(\round_in[0][1490] ) );
  AND U8368 ( .A(round_reg[1491]), .B(init), .Z(\round_in[0][1491] ) );
  AND U8369 ( .A(round_reg[1492]), .B(init), .Z(\round_in[0][1492] ) );
  AND U8370 ( .A(round_reg[1493]), .B(init), .Z(\round_in[0][1493] ) );
  AND U8371 ( .A(round_reg[1494]), .B(init), .Z(\round_in[0][1494] ) );
  AND U8372 ( .A(round_reg[1495]), .B(init), .Z(\round_in[0][1495] ) );
  AND U8373 ( .A(round_reg[1496]), .B(init), .Z(\round_in[0][1496] ) );
  AND U8374 ( .A(round_reg[1497]), .B(init), .Z(\round_in[0][1497] ) );
  AND U8375 ( .A(round_reg[1498]), .B(init), .Z(\round_in[0][1498] ) );
  AND U8376 ( .A(round_reg[1499]), .B(init), .Z(\round_in[0][1499] ) );
  NAND U8377 ( .A(init), .B(round_reg[149]), .Z(n2966) );
  NAND U8378 ( .A(n2778), .B(in[149]), .Z(n2965) );
  NAND U8379 ( .A(n2966), .B(n2965), .Z(\round_in[0][149] ) );
  NAND U8380 ( .A(init), .B(round_reg[14]), .Z(n2968) );
  NAND U8381 ( .A(n2778), .B(in[14]), .Z(n2967) );
  NAND U8382 ( .A(n2968), .B(n2967), .Z(\round_in[0][14] ) );
  AND U8383 ( .A(round_reg[1500]), .B(init), .Z(\round_in[0][1500] ) );
  AND U8384 ( .A(round_reg[1501]), .B(init), .Z(\round_in[0][1501] ) );
  AND U8385 ( .A(round_reg[1502]), .B(init), .Z(\round_in[0][1502] ) );
  AND U8386 ( .A(round_reg[1503]), .B(init), .Z(\round_in[0][1503] ) );
  AND U8387 ( .A(round_reg[1504]), .B(init), .Z(\round_in[0][1504] ) );
  AND U8388 ( .A(round_reg[1505]), .B(init), .Z(\round_in[0][1505] ) );
  AND U8389 ( .A(round_reg[1506]), .B(init), .Z(\round_in[0][1506] ) );
  AND U8390 ( .A(round_reg[1507]), .B(init), .Z(\round_in[0][1507] ) );
  AND U8391 ( .A(round_reg[1508]), .B(init), .Z(\round_in[0][1508] ) );
  AND U8392 ( .A(round_reg[1509]), .B(init), .Z(\round_in[0][1509] ) );
  NAND U8393 ( .A(init), .B(round_reg[150]), .Z(n2970) );
  NAND U8394 ( .A(n2778), .B(in[150]), .Z(n2969) );
  NAND U8395 ( .A(n2970), .B(n2969), .Z(\round_in[0][150] ) );
  AND U8396 ( .A(round_reg[1510]), .B(init), .Z(\round_in[0][1510] ) );
  AND U8397 ( .A(round_reg[1511]), .B(init), .Z(\round_in[0][1511] ) );
  AND U8398 ( .A(round_reg[1512]), .B(init), .Z(\round_in[0][1512] ) );
  AND U8399 ( .A(round_reg[1513]), .B(init), .Z(\round_in[0][1513] ) );
  AND U8400 ( .A(round_reg[1514]), .B(init), .Z(\round_in[0][1514] ) );
  AND U8401 ( .A(round_reg[1515]), .B(init), .Z(\round_in[0][1515] ) );
  AND U8402 ( .A(round_reg[1516]), .B(init), .Z(\round_in[0][1516] ) );
  AND U8403 ( .A(round_reg[1517]), .B(init), .Z(\round_in[0][1517] ) );
  AND U8404 ( .A(round_reg[1518]), .B(init), .Z(\round_in[0][1518] ) );
  AND U8405 ( .A(round_reg[1519]), .B(init), .Z(\round_in[0][1519] ) );
  NAND U8406 ( .A(init), .B(round_reg[151]), .Z(n2972) );
  NAND U8407 ( .A(n2778), .B(in[151]), .Z(n2971) );
  NAND U8408 ( .A(n2972), .B(n2971), .Z(\round_in[0][151] ) );
  AND U8409 ( .A(round_reg[1520]), .B(init), .Z(\round_in[0][1520] ) );
  AND U8410 ( .A(round_reg[1521]), .B(init), .Z(\round_in[0][1521] ) );
  AND U8411 ( .A(round_reg[1522]), .B(init), .Z(\round_in[0][1522] ) );
  AND U8412 ( .A(round_reg[1523]), .B(init), .Z(\round_in[0][1523] ) );
  AND U8413 ( .A(round_reg[1524]), .B(init), .Z(\round_in[0][1524] ) );
  AND U8414 ( .A(round_reg[1525]), .B(init), .Z(\round_in[0][1525] ) );
  AND U8415 ( .A(round_reg[1526]), .B(init), .Z(\round_in[0][1526] ) );
  AND U8416 ( .A(round_reg[1527]), .B(init), .Z(\round_in[0][1527] ) );
  AND U8417 ( .A(round_reg[1528]), .B(init), .Z(\round_in[0][1528] ) );
  AND U8418 ( .A(round_reg[1529]), .B(init), .Z(\round_in[0][1529] ) );
  NAND U8419 ( .A(init), .B(round_reg[152]), .Z(n2974) );
  NAND U8420 ( .A(n2778), .B(in[152]), .Z(n2973) );
  NAND U8421 ( .A(n2974), .B(n2973), .Z(\round_in[0][152] ) );
  AND U8422 ( .A(round_reg[1530]), .B(init), .Z(\round_in[0][1530] ) );
  AND U8423 ( .A(round_reg[1531]), .B(init), .Z(\round_in[0][1531] ) );
  AND U8424 ( .A(round_reg[1532]), .B(init), .Z(\round_in[0][1532] ) );
  AND U8425 ( .A(round_reg[1533]), .B(init), .Z(\round_in[0][1533] ) );
  AND U8426 ( .A(round_reg[1534]), .B(init), .Z(\round_in[0][1534] ) );
  AND U8427 ( .A(round_reg[1535]), .B(init), .Z(\round_in[0][1535] ) );
  AND U8428 ( .A(round_reg[1536]), .B(init), .Z(\round_in[0][1536] ) );
  AND U8429 ( .A(round_reg[1537]), .B(init), .Z(\round_in[0][1537] ) );
  AND U8430 ( .A(round_reg[1538]), .B(init), .Z(\round_in[0][1538] ) );
  AND U8431 ( .A(round_reg[1539]), .B(init), .Z(\round_in[0][1539] ) );
  NAND U8432 ( .A(init), .B(round_reg[153]), .Z(n2976) );
  NAND U8433 ( .A(n2778), .B(in[153]), .Z(n2975) );
  NAND U8434 ( .A(n2976), .B(n2975), .Z(\round_in[0][153] ) );
  AND U8435 ( .A(round_reg[1540]), .B(init), .Z(\round_in[0][1540] ) );
  AND U8436 ( .A(round_reg[1541]), .B(init), .Z(\round_in[0][1541] ) );
  AND U8437 ( .A(round_reg[1542]), .B(init), .Z(\round_in[0][1542] ) );
  AND U8438 ( .A(round_reg[1543]), .B(init), .Z(\round_in[0][1543] ) );
  AND U8439 ( .A(round_reg[1544]), .B(init), .Z(\round_in[0][1544] ) );
  AND U8440 ( .A(round_reg[1545]), .B(init), .Z(\round_in[0][1545] ) );
  AND U8441 ( .A(round_reg[1546]), .B(init), .Z(\round_in[0][1546] ) );
  AND U8442 ( .A(round_reg[1547]), .B(init), .Z(\round_in[0][1547] ) );
  AND U8443 ( .A(round_reg[1548]), .B(init), .Z(\round_in[0][1548] ) );
  AND U8444 ( .A(round_reg[1549]), .B(init), .Z(\round_in[0][1549] ) );
  NAND U8445 ( .A(init), .B(round_reg[154]), .Z(n2978) );
  NAND U8446 ( .A(n2778), .B(in[154]), .Z(n2977) );
  NAND U8447 ( .A(n2978), .B(n2977), .Z(\round_in[0][154] ) );
  AND U8448 ( .A(round_reg[1550]), .B(init), .Z(\round_in[0][1550] ) );
  AND U8449 ( .A(round_reg[1551]), .B(init), .Z(\round_in[0][1551] ) );
  AND U8450 ( .A(round_reg[1552]), .B(init), .Z(\round_in[0][1552] ) );
  AND U8451 ( .A(round_reg[1553]), .B(init), .Z(\round_in[0][1553] ) );
  AND U8452 ( .A(round_reg[1554]), .B(init), .Z(\round_in[0][1554] ) );
  AND U8453 ( .A(round_reg[1555]), .B(init), .Z(\round_in[0][1555] ) );
  AND U8454 ( .A(round_reg[1556]), .B(init), .Z(\round_in[0][1556] ) );
  AND U8455 ( .A(round_reg[1557]), .B(init), .Z(\round_in[0][1557] ) );
  AND U8456 ( .A(round_reg[1558]), .B(init), .Z(\round_in[0][1558] ) );
  AND U8457 ( .A(round_reg[1559]), .B(init), .Z(\round_in[0][1559] ) );
  NAND U8458 ( .A(init), .B(round_reg[155]), .Z(n2980) );
  NAND U8459 ( .A(n2779), .B(in[155]), .Z(n2979) );
  NAND U8460 ( .A(n2980), .B(n2979), .Z(\round_in[0][155] ) );
  AND U8461 ( .A(round_reg[1560]), .B(init), .Z(\round_in[0][1560] ) );
  AND U8462 ( .A(round_reg[1561]), .B(init), .Z(\round_in[0][1561] ) );
  AND U8463 ( .A(round_reg[1562]), .B(init), .Z(\round_in[0][1562] ) );
  AND U8464 ( .A(round_reg[1563]), .B(init), .Z(\round_in[0][1563] ) );
  AND U8465 ( .A(round_reg[1564]), .B(init), .Z(\round_in[0][1564] ) );
  AND U8466 ( .A(round_reg[1565]), .B(init), .Z(\round_in[0][1565] ) );
  AND U8467 ( .A(round_reg[1566]), .B(init), .Z(\round_in[0][1566] ) );
  AND U8468 ( .A(round_reg[1567]), .B(init), .Z(\round_in[0][1567] ) );
  AND U8469 ( .A(round_reg[1568]), .B(init), .Z(\round_in[0][1568] ) );
  AND U8470 ( .A(round_reg[1569]), .B(init), .Z(\round_in[0][1569] ) );
  NAND U8471 ( .A(init), .B(round_reg[156]), .Z(n2982) );
  NAND U8472 ( .A(n2779), .B(in[156]), .Z(n2981) );
  NAND U8473 ( .A(n2982), .B(n2981), .Z(\round_in[0][156] ) );
  AND U8474 ( .A(round_reg[1570]), .B(init), .Z(\round_in[0][1570] ) );
  AND U8475 ( .A(round_reg[1571]), .B(init), .Z(\round_in[0][1571] ) );
  AND U8476 ( .A(round_reg[1572]), .B(init), .Z(\round_in[0][1572] ) );
  AND U8477 ( .A(round_reg[1573]), .B(init), .Z(\round_in[0][1573] ) );
  AND U8478 ( .A(round_reg[1574]), .B(init), .Z(\round_in[0][1574] ) );
  AND U8479 ( .A(round_reg[1575]), .B(init), .Z(\round_in[0][1575] ) );
  AND U8480 ( .A(round_reg[1576]), .B(init), .Z(\round_in[0][1576] ) );
  AND U8481 ( .A(round_reg[1577]), .B(init), .Z(\round_in[0][1577] ) );
  AND U8482 ( .A(round_reg[1578]), .B(init), .Z(\round_in[0][1578] ) );
  AND U8483 ( .A(round_reg[1579]), .B(init), .Z(\round_in[0][1579] ) );
  NAND U8484 ( .A(init), .B(round_reg[157]), .Z(n2984) );
  NAND U8485 ( .A(n2779), .B(in[157]), .Z(n2983) );
  NAND U8486 ( .A(n2984), .B(n2983), .Z(\round_in[0][157] ) );
  AND U8487 ( .A(round_reg[1580]), .B(init), .Z(\round_in[0][1580] ) );
  AND U8488 ( .A(round_reg[1581]), .B(init), .Z(\round_in[0][1581] ) );
  AND U8489 ( .A(round_reg[1582]), .B(init), .Z(\round_in[0][1582] ) );
  AND U8490 ( .A(round_reg[1583]), .B(init), .Z(\round_in[0][1583] ) );
  AND U8491 ( .A(round_reg[1584]), .B(init), .Z(\round_in[0][1584] ) );
  AND U8492 ( .A(round_reg[1585]), .B(init), .Z(\round_in[0][1585] ) );
  AND U8493 ( .A(round_reg[1586]), .B(init), .Z(\round_in[0][1586] ) );
  AND U8494 ( .A(round_reg[1587]), .B(init), .Z(\round_in[0][1587] ) );
  AND U8495 ( .A(round_reg[1588]), .B(init), .Z(\round_in[0][1588] ) );
  AND U8496 ( .A(round_reg[1589]), .B(init), .Z(\round_in[0][1589] ) );
  NAND U8497 ( .A(init), .B(round_reg[158]), .Z(n2986) );
  NAND U8498 ( .A(n2779), .B(in[158]), .Z(n2985) );
  NAND U8499 ( .A(n2986), .B(n2985), .Z(\round_in[0][158] ) );
  AND U8500 ( .A(round_reg[1590]), .B(init), .Z(\round_in[0][1590] ) );
  AND U8501 ( .A(round_reg[1591]), .B(init), .Z(\round_in[0][1591] ) );
  AND U8502 ( .A(round_reg[1592]), .B(init), .Z(\round_in[0][1592] ) );
  AND U8503 ( .A(round_reg[1593]), .B(init), .Z(\round_in[0][1593] ) );
  AND U8504 ( .A(round_reg[1594]), .B(init), .Z(\round_in[0][1594] ) );
  AND U8505 ( .A(round_reg[1595]), .B(init), .Z(\round_in[0][1595] ) );
  AND U8506 ( .A(round_reg[1596]), .B(init), .Z(\round_in[0][1596] ) );
  AND U8507 ( .A(round_reg[1597]), .B(init), .Z(\round_in[0][1597] ) );
  AND U8508 ( .A(round_reg[1598]), .B(init), .Z(\round_in[0][1598] ) );
  AND U8509 ( .A(round_reg[1599]), .B(init), .Z(\round_in[0][1599] ) );
  NAND U8510 ( .A(init), .B(round_reg[159]), .Z(n2988) );
  NAND U8511 ( .A(n2779), .B(in[159]), .Z(n2987) );
  NAND U8512 ( .A(n2988), .B(n2987), .Z(\round_in[0][159] ) );
  NAND U8513 ( .A(init), .B(round_reg[15]), .Z(n2990) );
  NAND U8514 ( .A(n2779), .B(in[15]), .Z(n2989) );
  NAND U8515 ( .A(n2990), .B(n2989), .Z(\round_in[0][15] ) );
  NAND U8516 ( .A(init), .B(round_reg[160]), .Z(n2992) );
  NAND U8517 ( .A(n2779), .B(in[160]), .Z(n2991) );
  NAND U8518 ( .A(n2992), .B(n2991), .Z(\round_in[0][160] ) );
  NAND U8519 ( .A(init), .B(round_reg[161]), .Z(n2994) );
  NAND U8520 ( .A(n2780), .B(in[161]), .Z(n2993) );
  NAND U8521 ( .A(n2994), .B(n2993), .Z(\round_in[0][161] ) );
  NAND U8522 ( .A(init), .B(round_reg[162]), .Z(n2996) );
  NAND U8523 ( .A(n2780), .B(in[162]), .Z(n2995) );
  NAND U8524 ( .A(n2996), .B(n2995), .Z(\round_in[0][162] ) );
  NAND U8525 ( .A(init), .B(round_reg[163]), .Z(n2998) );
  NAND U8526 ( .A(n2780), .B(in[163]), .Z(n2997) );
  NAND U8527 ( .A(n2998), .B(n2997), .Z(\round_in[0][163] ) );
  NAND U8528 ( .A(init), .B(round_reg[164]), .Z(n3000) );
  NAND U8529 ( .A(n2780), .B(in[164]), .Z(n2999) );
  NAND U8530 ( .A(n3000), .B(n2999), .Z(\round_in[0][164] ) );
  NAND U8531 ( .A(init), .B(round_reg[165]), .Z(n3002) );
  NAND U8532 ( .A(n2780), .B(in[165]), .Z(n3001) );
  NAND U8533 ( .A(n3002), .B(n3001), .Z(\round_in[0][165] ) );
  NAND U8534 ( .A(init), .B(round_reg[166]), .Z(n3004) );
  NAND U8535 ( .A(n2780), .B(in[166]), .Z(n3003) );
  NAND U8536 ( .A(n3004), .B(n3003), .Z(\round_in[0][166] ) );
  NAND U8537 ( .A(init), .B(round_reg[167]), .Z(n3006) );
  NAND U8538 ( .A(n2780), .B(in[167]), .Z(n3005) );
  NAND U8539 ( .A(n3006), .B(n3005), .Z(\round_in[0][167] ) );
  NAND U8540 ( .A(init), .B(round_reg[168]), .Z(n3008) );
  NAND U8541 ( .A(n2781), .B(in[168]), .Z(n3007) );
  NAND U8542 ( .A(n3008), .B(n3007), .Z(\round_in[0][168] ) );
  NAND U8543 ( .A(init), .B(round_reg[169]), .Z(n3010) );
  NAND U8544 ( .A(n2781), .B(in[169]), .Z(n3009) );
  NAND U8545 ( .A(n3010), .B(n3009), .Z(\round_in[0][169] ) );
  NAND U8546 ( .A(init), .B(round_reg[16]), .Z(n3012) );
  NAND U8547 ( .A(n2781), .B(in[16]), .Z(n3011) );
  NAND U8548 ( .A(n3012), .B(n3011), .Z(\round_in[0][16] ) );
  NAND U8549 ( .A(init), .B(round_reg[170]), .Z(n3014) );
  NAND U8550 ( .A(n2781), .B(in[170]), .Z(n3013) );
  NAND U8551 ( .A(n3014), .B(n3013), .Z(\round_in[0][170] ) );
  NAND U8552 ( .A(init), .B(round_reg[171]), .Z(n3016) );
  NAND U8553 ( .A(n2781), .B(in[171]), .Z(n3015) );
  NAND U8554 ( .A(n3016), .B(n3015), .Z(\round_in[0][171] ) );
  NAND U8555 ( .A(init), .B(round_reg[172]), .Z(n3018) );
  NAND U8556 ( .A(n2781), .B(in[172]), .Z(n3017) );
  NAND U8557 ( .A(n3018), .B(n3017), .Z(\round_in[0][172] ) );
  NAND U8558 ( .A(init), .B(round_reg[173]), .Z(n3020) );
  NAND U8559 ( .A(n2781), .B(in[173]), .Z(n3019) );
  NAND U8560 ( .A(n3020), .B(n3019), .Z(\round_in[0][173] ) );
  NAND U8561 ( .A(init), .B(round_reg[174]), .Z(n3022) );
  NAND U8562 ( .A(n2782), .B(in[174]), .Z(n3021) );
  NAND U8563 ( .A(n3022), .B(n3021), .Z(\round_in[0][174] ) );
  NAND U8564 ( .A(init), .B(round_reg[175]), .Z(n3024) );
  NAND U8565 ( .A(n2782), .B(in[175]), .Z(n3023) );
  NAND U8566 ( .A(n3024), .B(n3023), .Z(\round_in[0][175] ) );
  NAND U8567 ( .A(init), .B(round_reg[176]), .Z(n3026) );
  NAND U8568 ( .A(n2782), .B(in[176]), .Z(n3025) );
  NAND U8569 ( .A(n3026), .B(n3025), .Z(\round_in[0][176] ) );
  NAND U8570 ( .A(init), .B(round_reg[177]), .Z(n3028) );
  NAND U8571 ( .A(n2782), .B(in[177]), .Z(n3027) );
  NAND U8572 ( .A(n3028), .B(n3027), .Z(\round_in[0][177] ) );
  NAND U8573 ( .A(init), .B(round_reg[178]), .Z(n3030) );
  NAND U8574 ( .A(n2782), .B(in[178]), .Z(n3029) );
  NAND U8575 ( .A(n3030), .B(n3029), .Z(\round_in[0][178] ) );
  NAND U8576 ( .A(init), .B(round_reg[179]), .Z(n3032) );
  NAND U8577 ( .A(n2782), .B(in[179]), .Z(n3031) );
  NAND U8578 ( .A(n3032), .B(n3031), .Z(\round_in[0][179] ) );
  NAND U8579 ( .A(init), .B(round_reg[17]), .Z(n3034) );
  NAND U8580 ( .A(n2782), .B(in[17]), .Z(n3033) );
  NAND U8581 ( .A(n3034), .B(n3033), .Z(\round_in[0][17] ) );
  NAND U8582 ( .A(init), .B(round_reg[180]), .Z(n3036) );
  NAND U8583 ( .A(n2783), .B(in[180]), .Z(n3035) );
  NAND U8584 ( .A(n3036), .B(n3035), .Z(\round_in[0][180] ) );
  NAND U8585 ( .A(init), .B(round_reg[181]), .Z(n3038) );
  NAND U8586 ( .A(n2783), .B(in[181]), .Z(n3037) );
  NAND U8587 ( .A(n3038), .B(n3037), .Z(\round_in[0][181] ) );
  NAND U8588 ( .A(init), .B(round_reg[182]), .Z(n3040) );
  NAND U8589 ( .A(n2783), .B(in[182]), .Z(n3039) );
  NAND U8590 ( .A(n3040), .B(n3039), .Z(\round_in[0][182] ) );
  NAND U8591 ( .A(init), .B(round_reg[183]), .Z(n3042) );
  NAND U8592 ( .A(n2783), .B(in[183]), .Z(n3041) );
  NAND U8593 ( .A(n3042), .B(n3041), .Z(\round_in[0][183] ) );
  NAND U8594 ( .A(init), .B(round_reg[184]), .Z(n3044) );
  NAND U8595 ( .A(n2783), .B(in[184]), .Z(n3043) );
  NAND U8596 ( .A(n3044), .B(n3043), .Z(\round_in[0][184] ) );
  NAND U8597 ( .A(init), .B(round_reg[185]), .Z(n3046) );
  NAND U8598 ( .A(n2783), .B(in[185]), .Z(n3045) );
  NAND U8599 ( .A(n3046), .B(n3045), .Z(\round_in[0][185] ) );
  NAND U8600 ( .A(init), .B(round_reg[186]), .Z(n3048) );
  NAND U8601 ( .A(n2783), .B(in[186]), .Z(n3047) );
  NAND U8602 ( .A(n3048), .B(n3047), .Z(\round_in[0][186] ) );
  NAND U8603 ( .A(init), .B(round_reg[187]), .Z(n3050) );
  NAND U8604 ( .A(n2784), .B(in[187]), .Z(n3049) );
  NAND U8605 ( .A(n3050), .B(n3049), .Z(\round_in[0][187] ) );
  NAND U8606 ( .A(init), .B(round_reg[188]), .Z(n3052) );
  NAND U8607 ( .A(n2784), .B(in[188]), .Z(n3051) );
  NAND U8608 ( .A(n3052), .B(n3051), .Z(\round_in[0][188] ) );
  NAND U8609 ( .A(init), .B(round_reg[189]), .Z(n3054) );
  NAND U8610 ( .A(n2784), .B(in[189]), .Z(n3053) );
  NAND U8611 ( .A(n3054), .B(n3053), .Z(\round_in[0][189] ) );
  NAND U8612 ( .A(init), .B(round_reg[18]), .Z(n3056) );
  NAND U8613 ( .A(n2784), .B(in[18]), .Z(n3055) );
  NAND U8614 ( .A(n3056), .B(n3055), .Z(\round_in[0][18] ) );
  NAND U8615 ( .A(init), .B(round_reg[190]), .Z(n3058) );
  NAND U8616 ( .A(n2784), .B(in[190]), .Z(n3057) );
  NAND U8617 ( .A(n3058), .B(n3057), .Z(\round_in[0][190] ) );
  NAND U8618 ( .A(init), .B(round_reg[191]), .Z(n3060) );
  NAND U8619 ( .A(n2784), .B(in[191]), .Z(n3059) );
  NAND U8620 ( .A(n3060), .B(n3059), .Z(\round_in[0][191] ) );
  NAND U8621 ( .A(init), .B(round_reg[192]), .Z(n3062) );
  NAND U8622 ( .A(n2784), .B(in[192]), .Z(n3061) );
  NAND U8623 ( .A(n3062), .B(n3061), .Z(\round_in[0][192] ) );
  NAND U8624 ( .A(init), .B(round_reg[193]), .Z(n3064) );
  NAND U8625 ( .A(n2785), .B(in[193]), .Z(n3063) );
  NAND U8626 ( .A(n3064), .B(n3063), .Z(\round_in[0][193] ) );
  NAND U8627 ( .A(init), .B(round_reg[194]), .Z(n3066) );
  NAND U8628 ( .A(n2785), .B(in[194]), .Z(n3065) );
  NAND U8629 ( .A(n3066), .B(n3065), .Z(\round_in[0][194] ) );
  NAND U8630 ( .A(init), .B(round_reg[195]), .Z(n3068) );
  NAND U8631 ( .A(n2785), .B(in[195]), .Z(n3067) );
  NAND U8632 ( .A(n3068), .B(n3067), .Z(\round_in[0][195] ) );
  NAND U8633 ( .A(init), .B(round_reg[196]), .Z(n3070) );
  NAND U8634 ( .A(n2785), .B(in[196]), .Z(n3069) );
  NAND U8635 ( .A(n3070), .B(n3069), .Z(\round_in[0][196] ) );
  NAND U8636 ( .A(init), .B(round_reg[197]), .Z(n3072) );
  NAND U8637 ( .A(n2785), .B(in[197]), .Z(n3071) );
  NAND U8638 ( .A(n3072), .B(n3071), .Z(\round_in[0][197] ) );
  NAND U8639 ( .A(init), .B(round_reg[198]), .Z(n3074) );
  NAND U8640 ( .A(n2785), .B(in[198]), .Z(n3073) );
  NAND U8641 ( .A(n3074), .B(n3073), .Z(\round_in[0][198] ) );
  NAND U8642 ( .A(init), .B(round_reg[199]), .Z(n3076) );
  NAND U8643 ( .A(n2785), .B(in[199]), .Z(n3075) );
  NAND U8644 ( .A(n3076), .B(n3075), .Z(\round_in[0][199] ) );
  NAND U8645 ( .A(init), .B(round_reg[19]), .Z(n3078) );
  NAND U8646 ( .A(n2786), .B(in[19]), .Z(n3077) );
  NAND U8647 ( .A(n3078), .B(n3077), .Z(\round_in[0][19] ) );
  NAND U8648 ( .A(init), .B(round_reg[1]), .Z(n3080) );
  NAND U8649 ( .A(n2786), .B(in[1]), .Z(n3079) );
  NAND U8650 ( .A(n3080), .B(n3079), .Z(\round_in[0][1] ) );
  NAND U8651 ( .A(init), .B(round_reg[200]), .Z(n3082) );
  NAND U8652 ( .A(n2786), .B(in[200]), .Z(n3081) );
  NAND U8653 ( .A(n3082), .B(n3081), .Z(\round_in[0][200] ) );
  NAND U8654 ( .A(init), .B(round_reg[201]), .Z(n3084) );
  NAND U8655 ( .A(n2786), .B(in[201]), .Z(n3083) );
  NAND U8656 ( .A(n3084), .B(n3083), .Z(\round_in[0][201] ) );
  NAND U8657 ( .A(init), .B(round_reg[202]), .Z(n3086) );
  NAND U8658 ( .A(n2786), .B(in[202]), .Z(n3085) );
  NAND U8659 ( .A(n3086), .B(n3085), .Z(\round_in[0][202] ) );
  NAND U8660 ( .A(init), .B(round_reg[203]), .Z(n3088) );
  NAND U8661 ( .A(n2786), .B(in[203]), .Z(n3087) );
  NAND U8662 ( .A(n3088), .B(n3087), .Z(\round_in[0][203] ) );
  NAND U8663 ( .A(init), .B(round_reg[204]), .Z(n3090) );
  NAND U8664 ( .A(n2786), .B(in[204]), .Z(n3089) );
  NAND U8665 ( .A(n3090), .B(n3089), .Z(\round_in[0][204] ) );
  NAND U8666 ( .A(init), .B(round_reg[205]), .Z(n3092) );
  NAND U8667 ( .A(n2787), .B(in[205]), .Z(n3091) );
  NAND U8668 ( .A(n3092), .B(n3091), .Z(\round_in[0][205] ) );
  NAND U8669 ( .A(init), .B(round_reg[206]), .Z(n3094) );
  NAND U8670 ( .A(n2787), .B(in[206]), .Z(n3093) );
  NAND U8671 ( .A(n3094), .B(n3093), .Z(\round_in[0][206] ) );
  NAND U8672 ( .A(init), .B(round_reg[207]), .Z(n3096) );
  NAND U8673 ( .A(n2787), .B(in[207]), .Z(n3095) );
  NAND U8674 ( .A(n3096), .B(n3095), .Z(\round_in[0][207] ) );
  NAND U8675 ( .A(init), .B(round_reg[208]), .Z(n3098) );
  NAND U8676 ( .A(n2787), .B(in[208]), .Z(n3097) );
  NAND U8677 ( .A(n3098), .B(n3097), .Z(\round_in[0][208] ) );
  NAND U8678 ( .A(init), .B(round_reg[209]), .Z(n3100) );
  NAND U8679 ( .A(n2787), .B(in[209]), .Z(n3099) );
  NAND U8680 ( .A(n3100), .B(n3099), .Z(\round_in[0][209] ) );
  NAND U8681 ( .A(init), .B(round_reg[20]), .Z(n3102) );
  NAND U8682 ( .A(n2787), .B(in[20]), .Z(n3101) );
  NAND U8683 ( .A(n3102), .B(n3101), .Z(\round_in[0][20] ) );
  NAND U8684 ( .A(init), .B(round_reg[210]), .Z(n3104) );
  NAND U8685 ( .A(n2787), .B(in[210]), .Z(n3103) );
  NAND U8686 ( .A(n3104), .B(n3103), .Z(\round_in[0][210] ) );
  NAND U8687 ( .A(init), .B(round_reg[211]), .Z(n3106) );
  NAND U8688 ( .A(n2788), .B(in[211]), .Z(n3105) );
  NAND U8689 ( .A(n3106), .B(n3105), .Z(\round_in[0][211] ) );
  NAND U8690 ( .A(init), .B(round_reg[212]), .Z(n3108) );
  NAND U8691 ( .A(n2788), .B(in[212]), .Z(n3107) );
  NAND U8692 ( .A(n3108), .B(n3107), .Z(\round_in[0][212] ) );
  NAND U8693 ( .A(init), .B(round_reg[213]), .Z(n3110) );
  NAND U8694 ( .A(n2788), .B(in[213]), .Z(n3109) );
  NAND U8695 ( .A(n3110), .B(n3109), .Z(\round_in[0][213] ) );
  NAND U8696 ( .A(init), .B(round_reg[214]), .Z(n3112) );
  NAND U8697 ( .A(n2788), .B(in[214]), .Z(n3111) );
  NAND U8698 ( .A(n3112), .B(n3111), .Z(\round_in[0][214] ) );
  NAND U8699 ( .A(init), .B(round_reg[215]), .Z(n3114) );
  NAND U8700 ( .A(n2788), .B(in[215]), .Z(n3113) );
  NAND U8701 ( .A(n3114), .B(n3113), .Z(\round_in[0][215] ) );
  NAND U8702 ( .A(init), .B(round_reg[216]), .Z(n3116) );
  NAND U8703 ( .A(n2788), .B(in[216]), .Z(n3115) );
  NAND U8704 ( .A(n3116), .B(n3115), .Z(\round_in[0][216] ) );
  NAND U8705 ( .A(init), .B(round_reg[217]), .Z(n3118) );
  NAND U8706 ( .A(n2788), .B(in[217]), .Z(n3117) );
  NAND U8707 ( .A(n3118), .B(n3117), .Z(\round_in[0][217] ) );
  NAND U8708 ( .A(init), .B(round_reg[218]), .Z(n3120) );
  NAND U8709 ( .A(n2789), .B(in[218]), .Z(n3119) );
  NAND U8710 ( .A(n3120), .B(n3119), .Z(\round_in[0][218] ) );
  NAND U8711 ( .A(init), .B(round_reg[219]), .Z(n3122) );
  NAND U8712 ( .A(n2789), .B(in[219]), .Z(n3121) );
  NAND U8713 ( .A(n3122), .B(n3121), .Z(\round_in[0][219] ) );
  NAND U8714 ( .A(init), .B(round_reg[21]), .Z(n3124) );
  NAND U8715 ( .A(n2789), .B(in[21]), .Z(n3123) );
  NAND U8716 ( .A(n3124), .B(n3123), .Z(\round_in[0][21] ) );
  NAND U8717 ( .A(init), .B(round_reg[220]), .Z(n3126) );
  NAND U8718 ( .A(n2789), .B(in[220]), .Z(n3125) );
  NAND U8719 ( .A(n3126), .B(n3125), .Z(\round_in[0][220] ) );
  NAND U8720 ( .A(init), .B(round_reg[221]), .Z(n3128) );
  NAND U8721 ( .A(n2789), .B(in[221]), .Z(n3127) );
  NAND U8722 ( .A(n3128), .B(n3127), .Z(\round_in[0][221] ) );
  NAND U8723 ( .A(init), .B(round_reg[222]), .Z(n3130) );
  NAND U8724 ( .A(n2789), .B(in[222]), .Z(n3129) );
  NAND U8725 ( .A(n3130), .B(n3129), .Z(\round_in[0][222] ) );
  NAND U8726 ( .A(init), .B(round_reg[223]), .Z(n3132) );
  NAND U8727 ( .A(n2789), .B(in[223]), .Z(n3131) );
  NAND U8728 ( .A(n3132), .B(n3131), .Z(\round_in[0][223] ) );
  NAND U8729 ( .A(init), .B(round_reg[224]), .Z(n3134) );
  NAND U8730 ( .A(n2790), .B(in[224]), .Z(n3133) );
  NAND U8731 ( .A(n3134), .B(n3133), .Z(\round_in[0][224] ) );
  NAND U8732 ( .A(init), .B(round_reg[225]), .Z(n3136) );
  NAND U8733 ( .A(n2790), .B(in[225]), .Z(n3135) );
  NAND U8734 ( .A(n3136), .B(n3135), .Z(\round_in[0][225] ) );
  NAND U8735 ( .A(init), .B(round_reg[226]), .Z(n3138) );
  NAND U8736 ( .A(n2790), .B(in[226]), .Z(n3137) );
  NAND U8737 ( .A(n3138), .B(n3137), .Z(\round_in[0][226] ) );
  NAND U8738 ( .A(init), .B(round_reg[227]), .Z(n3140) );
  NAND U8739 ( .A(n2790), .B(in[227]), .Z(n3139) );
  NAND U8740 ( .A(n3140), .B(n3139), .Z(\round_in[0][227] ) );
  NAND U8741 ( .A(init), .B(round_reg[228]), .Z(n3142) );
  NAND U8742 ( .A(n2790), .B(in[228]), .Z(n3141) );
  NAND U8743 ( .A(n3142), .B(n3141), .Z(\round_in[0][228] ) );
  NAND U8744 ( .A(init), .B(round_reg[229]), .Z(n3144) );
  NAND U8745 ( .A(n2790), .B(in[229]), .Z(n3143) );
  NAND U8746 ( .A(n3144), .B(n3143), .Z(\round_in[0][229] ) );
  NAND U8747 ( .A(init), .B(round_reg[22]), .Z(n3146) );
  NAND U8748 ( .A(n2790), .B(in[22]), .Z(n3145) );
  NAND U8749 ( .A(n3146), .B(n3145), .Z(\round_in[0][22] ) );
  NAND U8750 ( .A(init), .B(round_reg[230]), .Z(n3148) );
  NAND U8751 ( .A(n2791), .B(in[230]), .Z(n3147) );
  NAND U8752 ( .A(n3148), .B(n3147), .Z(\round_in[0][230] ) );
  NAND U8753 ( .A(init), .B(round_reg[231]), .Z(n3150) );
  NAND U8754 ( .A(n2791), .B(in[231]), .Z(n3149) );
  NAND U8755 ( .A(n3150), .B(n3149), .Z(\round_in[0][231] ) );
  NAND U8756 ( .A(init), .B(round_reg[232]), .Z(n3152) );
  NAND U8757 ( .A(n2791), .B(in[232]), .Z(n3151) );
  NAND U8758 ( .A(n3152), .B(n3151), .Z(\round_in[0][232] ) );
  NAND U8759 ( .A(init), .B(round_reg[233]), .Z(n3154) );
  NAND U8760 ( .A(n2791), .B(in[233]), .Z(n3153) );
  NAND U8761 ( .A(n3154), .B(n3153), .Z(\round_in[0][233] ) );
  NAND U8762 ( .A(init), .B(round_reg[234]), .Z(n3156) );
  NAND U8763 ( .A(n2791), .B(in[234]), .Z(n3155) );
  NAND U8764 ( .A(n3156), .B(n3155), .Z(\round_in[0][234] ) );
  NAND U8765 ( .A(init), .B(round_reg[235]), .Z(n3158) );
  NAND U8766 ( .A(n2791), .B(in[235]), .Z(n3157) );
  NAND U8767 ( .A(n3158), .B(n3157), .Z(\round_in[0][235] ) );
  NAND U8768 ( .A(init), .B(round_reg[236]), .Z(n3160) );
  NAND U8769 ( .A(n2791), .B(in[236]), .Z(n3159) );
  NAND U8770 ( .A(n3160), .B(n3159), .Z(\round_in[0][236] ) );
  NAND U8771 ( .A(init), .B(round_reg[237]), .Z(n3162) );
  NAND U8772 ( .A(n2792), .B(in[237]), .Z(n3161) );
  NAND U8773 ( .A(n3162), .B(n3161), .Z(\round_in[0][237] ) );
  NAND U8774 ( .A(init), .B(round_reg[238]), .Z(n3164) );
  NAND U8775 ( .A(n2792), .B(in[238]), .Z(n3163) );
  NAND U8776 ( .A(n3164), .B(n3163), .Z(\round_in[0][238] ) );
  NAND U8777 ( .A(init), .B(round_reg[239]), .Z(n3166) );
  NAND U8778 ( .A(n2792), .B(in[239]), .Z(n3165) );
  NAND U8779 ( .A(n3166), .B(n3165), .Z(\round_in[0][239] ) );
  NAND U8780 ( .A(init), .B(round_reg[23]), .Z(n3168) );
  NAND U8781 ( .A(n2792), .B(in[23]), .Z(n3167) );
  NAND U8782 ( .A(n3168), .B(n3167), .Z(\round_in[0][23] ) );
  NAND U8783 ( .A(init), .B(round_reg[240]), .Z(n3170) );
  NAND U8784 ( .A(n2792), .B(in[240]), .Z(n3169) );
  NAND U8785 ( .A(n3170), .B(n3169), .Z(\round_in[0][240] ) );
  NAND U8786 ( .A(init), .B(round_reg[241]), .Z(n3172) );
  NAND U8787 ( .A(n2792), .B(in[241]), .Z(n3171) );
  NAND U8788 ( .A(n3172), .B(n3171), .Z(\round_in[0][241] ) );
  NAND U8789 ( .A(init), .B(round_reg[242]), .Z(n3174) );
  NAND U8790 ( .A(n2792), .B(in[242]), .Z(n3173) );
  NAND U8791 ( .A(n3174), .B(n3173), .Z(\round_in[0][242] ) );
  NAND U8792 ( .A(init), .B(round_reg[243]), .Z(n3176) );
  NAND U8793 ( .A(n2793), .B(in[243]), .Z(n3175) );
  NAND U8794 ( .A(n3176), .B(n3175), .Z(\round_in[0][243] ) );
  NAND U8795 ( .A(init), .B(round_reg[244]), .Z(n3178) );
  NAND U8796 ( .A(n2793), .B(in[244]), .Z(n3177) );
  NAND U8797 ( .A(n3178), .B(n3177), .Z(\round_in[0][244] ) );
  NAND U8798 ( .A(init), .B(round_reg[245]), .Z(n3180) );
  NAND U8799 ( .A(n2793), .B(in[245]), .Z(n3179) );
  NAND U8800 ( .A(n3180), .B(n3179), .Z(\round_in[0][245] ) );
  NAND U8801 ( .A(init), .B(round_reg[246]), .Z(n3182) );
  NAND U8802 ( .A(n2793), .B(in[246]), .Z(n3181) );
  NAND U8803 ( .A(n3182), .B(n3181), .Z(\round_in[0][246] ) );
  NAND U8804 ( .A(init), .B(round_reg[247]), .Z(n3184) );
  NAND U8805 ( .A(n2793), .B(in[247]), .Z(n3183) );
  NAND U8806 ( .A(n3184), .B(n3183), .Z(\round_in[0][247] ) );
  NAND U8807 ( .A(init), .B(round_reg[248]), .Z(n3186) );
  NAND U8808 ( .A(n2793), .B(in[248]), .Z(n3185) );
  NAND U8809 ( .A(n3186), .B(n3185), .Z(\round_in[0][248] ) );
  NAND U8810 ( .A(init), .B(round_reg[249]), .Z(n3188) );
  NAND U8811 ( .A(n2793), .B(in[249]), .Z(n3187) );
  NAND U8812 ( .A(n3188), .B(n3187), .Z(\round_in[0][249] ) );
  NAND U8813 ( .A(init), .B(round_reg[24]), .Z(n3190) );
  NAND U8814 ( .A(n2794), .B(in[24]), .Z(n3189) );
  NAND U8815 ( .A(n3190), .B(n3189), .Z(\round_in[0][24] ) );
  NAND U8816 ( .A(init), .B(round_reg[250]), .Z(n3192) );
  NAND U8817 ( .A(n2794), .B(in[250]), .Z(n3191) );
  NAND U8818 ( .A(n3192), .B(n3191), .Z(\round_in[0][250] ) );
  NAND U8819 ( .A(init), .B(round_reg[251]), .Z(n3194) );
  NAND U8820 ( .A(n2794), .B(in[251]), .Z(n3193) );
  NAND U8821 ( .A(n3194), .B(n3193), .Z(\round_in[0][251] ) );
  NAND U8822 ( .A(init), .B(round_reg[252]), .Z(n3196) );
  NAND U8823 ( .A(n2794), .B(in[252]), .Z(n3195) );
  NAND U8824 ( .A(n3196), .B(n3195), .Z(\round_in[0][252] ) );
  NAND U8825 ( .A(init), .B(round_reg[253]), .Z(n3198) );
  NAND U8826 ( .A(n2794), .B(in[253]), .Z(n3197) );
  NAND U8827 ( .A(n3198), .B(n3197), .Z(\round_in[0][253] ) );
  NAND U8828 ( .A(init), .B(round_reg[254]), .Z(n3200) );
  NAND U8829 ( .A(n2794), .B(in[254]), .Z(n3199) );
  NAND U8830 ( .A(n3200), .B(n3199), .Z(\round_in[0][254] ) );
  NAND U8831 ( .A(init), .B(round_reg[255]), .Z(n3202) );
  NAND U8832 ( .A(n2794), .B(in[255]), .Z(n3201) );
  NAND U8833 ( .A(n3202), .B(n3201), .Z(\round_in[0][255] ) );
  NAND U8834 ( .A(init), .B(round_reg[256]), .Z(n3204) );
  NAND U8835 ( .A(n2795), .B(in[256]), .Z(n3203) );
  NAND U8836 ( .A(n3204), .B(n3203), .Z(\round_in[0][256] ) );
  NAND U8837 ( .A(init), .B(round_reg[257]), .Z(n3206) );
  NAND U8838 ( .A(n2795), .B(in[257]), .Z(n3205) );
  NAND U8839 ( .A(n3206), .B(n3205), .Z(\round_in[0][257] ) );
  NAND U8840 ( .A(init), .B(round_reg[258]), .Z(n3208) );
  NAND U8841 ( .A(n2795), .B(in[258]), .Z(n3207) );
  NAND U8842 ( .A(n3208), .B(n3207), .Z(\round_in[0][258] ) );
  NAND U8843 ( .A(init), .B(round_reg[259]), .Z(n3210) );
  NAND U8844 ( .A(n2795), .B(in[259]), .Z(n3209) );
  NAND U8845 ( .A(n3210), .B(n3209), .Z(\round_in[0][259] ) );
  NAND U8846 ( .A(init), .B(round_reg[25]), .Z(n3212) );
  NAND U8847 ( .A(n2795), .B(in[25]), .Z(n3211) );
  NAND U8848 ( .A(n3212), .B(n3211), .Z(\round_in[0][25] ) );
  NAND U8849 ( .A(init), .B(round_reg[260]), .Z(n3214) );
  NAND U8850 ( .A(n2795), .B(in[260]), .Z(n3213) );
  NAND U8851 ( .A(n3214), .B(n3213), .Z(\round_in[0][260] ) );
  NAND U8852 ( .A(init), .B(round_reg[261]), .Z(n3216) );
  NAND U8853 ( .A(n2795), .B(in[261]), .Z(n3215) );
  NAND U8854 ( .A(n3216), .B(n3215), .Z(\round_in[0][261] ) );
  NAND U8855 ( .A(init), .B(round_reg[262]), .Z(n3218) );
  NAND U8856 ( .A(n2796), .B(in[262]), .Z(n3217) );
  NAND U8857 ( .A(n3218), .B(n3217), .Z(\round_in[0][262] ) );
  NAND U8858 ( .A(init), .B(round_reg[263]), .Z(n3220) );
  NAND U8859 ( .A(n2796), .B(in[263]), .Z(n3219) );
  NAND U8860 ( .A(n3220), .B(n3219), .Z(\round_in[0][263] ) );
  NAND U8861 ( .A(init), .B(round_reg[264]), .Z(n3222) );
  NAND U8862 ( .A(n2796), .B(in[264]), .Z(n3221) );
  NAND U8863 ( .A(n3222), .B(n3221), .Z(\round_in[0][264] ) );
  NAND U8864 ( .A(init), .B(round_reg[265]), .Z(n3224) );
  NAND U8865 ( .A(n2796), .B(in[265]), .Z(n3223) );
  NAND U8866 ( .A(n3224), .B(n3223), .Z(\round_in[0][265] ) );
  NAND U8867 ( .A(init), .B(round_reg[266]), .Z(n3226) );
  NAND U8868 ( .A(n2796), .B(in[266]), .Z(n3225) );
  NAND U8869 ( .A(n3226), .B(n3225), .Z(\round_in[0][266] ) );
  NAND U8870 ( .A(init), .B(round_reg[267]), .Z(n3228) );
  NAND U8871 ( .A(n2796), .B(in[267]), .Z(n3227) );
  NAND U8872 ( .A(n3228), .B(n3227), .Z(\round_in[0][267] ) );
  NAND U8873 ( .A(init), .B(round_reg[268]), .Z(n3230) );
  NAND U8874 ( .A(n2796), .B(in[268]), .Z(n3229) );
  NAND U8875 ( .A(n3230), .B(n3229), .Z(\round_in[0][268] ) );
  NAND U8876 ( .A(init), .B(round_reg[269]), .Z(n3232) );
  NAND U8877 ( .A(n2797), .B(in[269]), .Z(n3231) );
  NAND U8878 ( .A(n3232), .B(n3231), .Z(\round_in[0][269] ) );
  NAND U8879 ( .A(init), .B(round_reg[26]), .Z(n3234) );
  NAND U8880 ( .A(n2797), .B(in[26]), .Z(n3233) );
  NAND U8881 ( .A(n3234), .B(n3233), .Z(\round_in[0][26] ) );
  NAND U8882 ( .A(init), .B(round_reg[270]), .Z(n3236) );
  NAND U8883 ( .A(n2797), .B(in[270]), .Z(n3235) );
  NAND U8884 ( .A(n3236), .B(n3235), .Z(\round_in[0][270] ) );
  NAND U8885 ( .A(init), .B(round_reg[271]), .Z(n3238) );
  NAND U8886 ( .A(n2797), .B(in[271]), .Z(n3237) );
  NAND U8887 ( .A(n3238), .B(n3237), .Z(\round_in[0][271] ) );
  NAND U8888 ( .A(init), .B(round_reg[272]), .Z(n3240) );
  NAND U8889 ( .A(n2797), .B(in[272]), .Z(n3239) );
  NAND U8890 ( .A(n3240), .B(n3239), .Z(\round_in[0][272] ) );
  NAND U8891 ( .A(init), .B(round_reg[273]), .Z(n3242) );
  NAND U8892 ( .A(n2797), .B(in[273]), .Z(n3241) );
  NAND U8893 ( .A(n3242), .B(n3241), .Z(\round_in[0][273] ) );
  NAND U8894 ( .A(init), .B(round_reg[274]), .Z(n3244) );
  NAND U8895 ( .A(n2797), .B(in[274]), .Z(n3243) );
  NAND U8896 ( .A(n3244), .B(n3243), .Z(\round_in[0][274] ) );
  NAND U8897 ( .A(init), .B(round_reg[275]), .Z(n3246) );
  NAND U8898 ( .A(n2798), .B(in[275]), .Z(n3245) );
  NAND U8899 ( .A(n3246), .B(n3245), .Z(\round_in[0][275] ) );
  NAND U8900 ( .A(init), .B(round_reg[276]), .Z(n3248) );
  NAND U8901 ( .A(n2798), .B(in[276]), .Z(n3247) );
  NAND U8902 ( .A(n3248), .B(n3247), .Z(\round_in[0][276] ) );
  NAND U8903 ( .A(init), .B(round_reg[277]), .Z(n3250) );
  NAND U8904 ( .A(n2798), .B(in[277]), .Z(n3249) );
  NAND U8905 ( .A(n3250), .B(n3249), .Z(\round_in[0][277] ) );
  NAND U8906 ( .A(init), .B(round_reg[278]), .Z(n3252) );
  NAND U8907 ( .A(n2798), .B(in[278]), .Z(n3251) );
  NAND U8908 ( .A(n3252), .B(n3251), .Z(\round_in[0][278] ) );
  NAND U8909 ( .A(init), .B(round_reg[279]), .Z(n3254) );
  NAND U8910 ( .A(n2798), .B(in[279]), .Z(n3253) );
  NAND U8911 ( .A(n3254), .B(n3253), .Z(\round_in[0][279] ) );
  NAND U8912 ( .A(init), .B(round_reg[27]), .Z(n3256) );
  NAND U8913 ( .A(n2798), .B(in[27]), .Z(n3255) );
  NAND U8914 ( .A(n3256), .B(n3255), .Z(\round_in[0][27] ) );
  NAND U8915 ( .A(init), .B(round_reg[280]), .Z(n3258) );
  NAND U8916 ( .A(n2798), .B(in[280]), .Z(n3257) );
  NAND U8917 ( .A(n3258), .B(n3257), .Z(\round_in[0][280] ) );
  NAND U8918 ( .A(init), .B(round_reg[281]), .Z(n3260) );
  NAND U8919 ( .A(n2799), .B(in[281]), .Z(n3259) );
  NAND U8920 ( .A(n3260), .B(n3259), .Z(\round_in[0][281] ) );
  NAND U8921 ( .A(init), .B(round_reg[282]), .Z(n3262) );
  NAND U8922 ( .A(n2799), .B(in[282]), .Z(n3261) );
  NAND U8923 ( .A(n3262), .B(n3261), .Z(\round_in[0][282] ) );
  NAND U8924 ( .A(init), .B(round_reg[283]), .Z(n3264) );
  NAND U8925 ( .A(n2799), .B(in[283]), .Z(n3263) );
  NAND U8926 ( .A(n3264), .B(n3263), .Z(\round_in[0][283] ) );
  NAND U8927 ( .A(init), .B(round_reg[284]), .Z(n3266) );
  NAND U8928 ( .A(n2799), .B(in[284]), .Z(n3265) );
  NAND U8929 ( .A(n3266), .B(n3265), .Z(\round_in[0][284] ) );
  NAND U8930 ( .A(init), .B(round_reg[285]), .Z(n3268) );
  NAND U8931 ( .A(n2799), .B(in[285]), .Z(n3267) );
  NAND U8932 ( .A(n3268), .B(n3267), .Z(\round_in[0][285] ) );
  NAND U8933 ( .A(init), .B(round_reg[286]), .Z(n3270) );
  NAND U8934 ( .A(n2799), .B(in[286]), .Z(n3269) );
  NAND U8935 ( .A(n3270), .B(n3269), .Z(\round_in[0][286] ) );
  NAND U8936 ( .A(init), .B(round_reg[287]), .Z(n3272) );
  NAND U8937 ( .A(n2799), .B(in[287]), .Z(n3271) );
  NAND U8938 ( .A(n3272), .B(n3271), .Z(\round_in[0][287] ) );
  NAND U8939 ( .A(init), .B(round_reg[288]), .Z(n3274) );
  NAND U8940 ( .A(n2800), .B(in[288]), .Z(n3273) );
  NAND U8941 ( .A(n3274), .B(n3273), .Z(\round_in[0][288] ) );
  NAND U8942 ( .A(init), .B(round_reg[289]), .Z(n3276) );
  NAND U8943 ( .A(n2800), .B(in[289]), .Z(n3275) );
  NAND U8944 ( .A(n3276), .B(n3275), .Z(\round_in[0][289] ) );
  NAND U8945 ( .A(init), .B(round_reg[28]), .Z(n3278) );
  NAND U8946 ( .A(n2800), .B(in[28]), .Z(n3277) );
  NAND U8947 ( .A(n3278), .B(n3277), .Z(\round_in[0][28] ) );
  NAND U8948 ( .A(init), .B(round_reg[290]), .Z(n3280) );
  NAND U8949 ( .A(n2800), .B(in[290]), .Z(n3279) );
  NAND U8950 ( .A(n3280), .B(n3279), .Z(\round_in[0][290] ) );
  NAND U8951 ( .A(init), .B(round_reg[291]), .Z(n3282) );
  NAND U8952 ( .A(n2800), .B(in[291]), .Z(n3281) );
  NAND U8953 ( .A(n3282), .B(n3281), .Z(\round_in[0][291] ) );
  NAND U8954 ( .A(init), .B(round_reg[292]), .Z(n3284) );
  NAND U8955 ( .A(n2800), .B(in[292]), .Z(n3283) );
  NAND U8956 ( .A(n3284), .B(n3283), .Z(\round_in[0][292] ) );
  NAND U8957 ( .A(init), .B(round_reg[293]), .Z(n3286) );
  NAND U8958 ( .A(n2800), .B(in[293]), .Z(n3285) );
  NAND U8959 ( .A(n3286), .B(n3285), .Z(\round_in[0][293] ) );
  NAND U8960 ( .A(init), .B(round_reg[294]), .Z(n3288) );
  NAND U8961 ( .A(n2801), .B(in[294]), .Z(n3287) );
  NAND U8962 ( .A(n3288), .B(n3287), .Z(\round_in[0][294] ) );
  NAND U8963 ( .A(init), .B(round_reg[295]), .Z(n3290) );
  NAND U8964 ( .A(n2801), .B(in[295]), .Z(n3289) );
  NAND U8965 ( .A(n3290), .B(n3289), .Z(\round_in[0][295] ) );
  NAND U8966 ( .A(init), .B(round_reg[296]), .Z(n3292) );
  NAND U8967 ( .A(n2801), .B(in[296]), .Z(n3291) );
  NAND U8968 ( .A(n3292), .B(n3291), .Z(\round_in[0][296] ) );
  NAND U8969 ( .A(init), .B(round_reg[297]), .Z(n3294) );
  NAND U8970 ( .A(n2801), .B(in[297]), .Z(n3293) );
  NAND U8971 ( .A(n3294), .B(n3293), .Z(\round_in[0][297] ) );
  NAND U8972 ( .A(init), .B(round_reg[298]), .Z(n3296) );
  NAND U8973 ( .A(n2801), .B(in[298]), .Z(n3295) );
  NAND U8974 ( .A(n3296), .B(n3295), .Z(\round_in[0][298] ) );
  NAND U8975 ( .A(init), .B(round_reg[299]), .Z(n3298) );
  NAND U8976 ( .A(n2801), .B(in[299]), .Z(n3297) );
  NAND U8977 ( .A(n3298), .B(n3297), .Z(\round_in[0][299] ) );
  NAND U8978 ( .A(init), .B(round_reg[29]), .Z(n3300) );
  NAND U8979 ( .A(n2801), .B(in[29]), .Z(n3299) );
  NAND U8980 ( .A(n3300), .B(n3299), .Z(\round_in[0][29] ) );
  NAND U8981 ( .A(init), .B(round_reg[2]), .Z(n3302) );
  NAND U8982 ( .A(n2802), .B(in[2]), .Z(n3301) );
  NAND U8983 ( .A(n3302), .B(n3301), .Z(\round_in[0][2] ) );
  NAND U8984 ( .A(init), .B(round_reg[300]), .Z(n3304) );
  NAND U8985 ( .A(n2802), .B(in[300]), .Z(n3303) );
  NAND U8986 ( .A(n3304), .B(n3303), .Z(\round_in[0][300] ) );
  NAND U8987 ( .A(init), .B(round_reg[301]), .Z(n3306) );
  NAND U8988 ( .A(n2802), .B(in[301]), .Z(n3305) );
  NAND U8989 ( .A(n3306), .B(n3305), .Z(\round_in[0][301] ) );
  NAND U8990 ( .A(init), .B(round_reg[302]), .Z(n3308) );
  NAND U8991 ( .A(n2802), .B(in[302]), .Z(n3307) );
  NAND U8992 ( .A(n3308), .B(n3307), .Z(\round_in[0][302] ) );
  NAND U8993 ( .A(init), .B(round_reg[303]), .Z(n3310) );
  NAND U8994 ( .A(n2802), .B(in[303]), .Z(n3309) );
  NAND U8995 ( .A(n3310), .B(n3309), .Z(\round_in[0][303] ) );
  NAND U8996 ( .A(init), .B(round_reg[304]), .Z(n3312) );
  NAND U8997 ( .A(n2802), .B(in[304]), .Z(n3311) );
  NAND U8998 ( .A(n3312), .B(n3311), .Z(\round_in[0][304] ) );
  NAND U8999 ( .A(init), .B(round_reg[305]), .Z(n3314) );
  NAND U9000 ( .A(n2802), .B(in[305]), .Z(n3313) );
  NAND U9001 ( .A(n3314), .B(n3313), .Z(\round_in[0][305] ) );
  NAND U9002 ( .A(init), .B(round_reg[306]), .Z(n3316) );
  NAND U9003 ( .A(n2803), .B(in[306]), .Z(n3315) );
  NAND U9004 ( .A(n3316), .B(n3315), .Z(\round_in[0][306] ) );
  NAND U9005 ( .A(init), .B(round_reg[307]), .Z(n3318) );
  NAND U9006 ( .A(n2803), .B(in[307]), .Z(n3317) );
  NAND U9007 ( .A(n3318), .B(n3317), .Z(\round_in[0][307] ) );
  NAND U9008 ( .A(init), .B(round_reg[308]), .Z(n3320) );
  NAND U9009 ( .A(n2803), .B(in[308]), .Z(n3319) );
  NAND U9010 ( .A(n3320), .B(n3319), .Z(\round_in[0][308] ) );
  NAND U9011 ( .A(init), .B(round_reg[309]), .Z(n3322) );
  NAND U9012 ( .A(n2803), .B(in[309]), .Z(n3321) );
  NAND U9013 ( .A(n3322), .B(n3321), .Z(\round_in[0][309] ) );
  NAND U9014 ( .A(init), .B(round_reg[30]), .Z(n3324) );
  NAND U9015 ( .A(n2803), .B(in[30]), .Z(n3323) );
  NAND U9016 ( .A(n3324), .B(n3323), .Z(\round_in[0][30] ) );
  NAND U9017 ( .A(init), .B(round_reg[310]), .Z(n3326) );
  NAND U9018 ( .A(n2803), .B(in[310]), .Z(n3325) );
  NAND U9019 ( .A(n3326), .B(n3325), .Z(\round_in[0][310] ) );
  NAND U9020 ( .A(init), .B(round_reg[311]), .Z(n3328) );
  NAND U9021 ( .A(n2803), .B(in[311]), .Z(n3327) );
  NAND U9022 ( .A(n3328), .B(n3327), .Z(\round_in[0][311] ) );
  NAND U9023 ( .A(init), .B(round_reg[312]), .Z(n3330) );
  NAND U9024 ( .A(n2804), .B(in[312]), .Z(n3329) );
  NAND U9025 ( .A(n3330), .B(n3329), .Z(\round_in[0][312] ) );
  NAND U9026 ( .A(init), .B(round_reg[313]), .Z(n3332) );
  NAND U9027 ( .A(n2804), .B(in[313]), .Z(n3331) );
  NAND U9028 ( .A(n3332), .B(n3331), .Z(\round_in[0][313] ) );
  NAND U9029 ( .A(init), .B(round_reg[314]), .Z(n3334) );
  NAND U9030 ( .A(n2804), .B(in[314]), .Z(n3333) );
  NAND U9031 ( .A(n3334), .B(n3333), .Z(\round_in[0][314] ) );
  NAND U9032 ( .A(init), .B(round_reg[315]), .Z(n3336) );
  NAND U9033 ( .A(n2804), .B(in[315]), .Z(n3335) );
  NAND U9034 ( .A(n3336), .B(n3335), .Z(\round_in[0][315] ) );
  NAND U9035 ( .A(init), .B(round_reg[316]), .Z(n3338) );
  NAND U9036 ( .A(n2804), .B(in[316]), .Z(n3337) );
  NAND U9037 ( .A(n3338), .B(n3337), .Z(\round_in[0][316] ) );
  NAND U9038 ( .A(init), .B(round_reg[317]), .Z(n3340) );
  NAND U9039 ( .A(n2804), .B(in[317]), .Z(n3339) );
  NAND U9040 ( .A(n3340), .B(n3339), .Z(\round_in[0][317] ) );
  NAND U9041 ( .A(init), .B(round_reg[318]), .Z(n3342) );
  NAND U9042 ( .A(n2804), .B(in[318]), .Z(n3341) );
  NAND U9043 ( .A(n3342), .B(n3341), .Z(\round_in[0][318] ) );
  NAND U9044 ( .A(init), .B(round_reg[319]), .Z(n3344) );
  NAND U9045 ( .A(n2805), .B(in[319]), .Z(n3343) );
  NAND U9046 ( .A(n3344), .B(n3343), .Z(\round_in[0][319] ) );
  NAND U9047 ( .A(init), .B(round_reg[31]), .Z(n3346) );
  NAND U9048 ( .A(n2805), .B(in[31]), .Z(n3345) );
  NAND U9049 ( .A(n3346), .B(n3345), .Z(\round_in[0][31] ) );
  NAND U9050 ( .A(init), .B(round_reg[320]), .Z(n3348) );
  NAND U9051 ( .A(n2805), .B(in[320]), .Z(n3347) );
  NAND U9052 ( .A(n3348), .B(n3347), .Z(\round_in[0][320] ) );
  NAND U9053 ( .A(init), .B(round_reg[321]), .Z(n3350) );
  NAND U9054 ( .A(n2805), .B(in[321]), .Z(n3349) );
  NAND U9055 ( .A(n3350), .B(n3349), .Z(\round_in[0][321] ) );
  NAND U9056 ( .A(init), .B(round_reg[322]), .Z(n3352) );
  NAND U9057 ( .A(n2805), .B(in[322]), .Z(n3351) );
  NAND U9058 ( .A(n3352), .B(n3351), .Z(\round_in[0][322] ) );
  NAND U9059 ( .A(init), .B(round_reg[323]), .Z(n3354) );
  NAND U9060 ( .A(n2805), .B(in[323]), .Z(n3353) );
  NAND U9061 ( .A(n3354), .B(n3353), .Z(\round_in[0][323] ) );
  NAND U9062 ( .A(init), .B(round_reg[324]), .Z(n3356) );
  NAND U9063 ( .A(n2805), .B(in[324]), .Z(n3355) );
  NAND U9064 ( .A(n3356), .B(n3355), .Z(\round_in[0][324] ) );
  NAND U9065 ( .A(init), .B(round_reg[325]), .Z(n3358) );
  NAND U9066 ( .A(n2806), .B(in[325]), .Z(n3357) );
  NAND U9067 ( .A(n3358), .B(n3357), .Z(\round_in[0][325] ) );
  NAND U9068 ( .A(init), .B(round_reg[326]), .Z(n3360) );
  NAND U9069 ( .A(n2806), .B(in[326]), .Z(n3359) );
  NAND U9070 ( .A(n3360), .B(n3359), .Z(\round_in[0][326] ) );
  NAND U9071 ( .A(init), .B(round_reg[327]), .Z(n3362) );
  NAND U9072 ( .A(n2806), .B(in[327]), .Z(n3361) );
  NAND U9073 ( .A(n3362), .B(n3361), .Z(\round_in[0][327] ) );
  NAND U9074 ( .A(init), .B(round_reg[328]), .Z(n3364) );
  NAND U9075 ( .A(n2806), .B(in[328]), .Z(n3363) );
  NAND U9076 ( .A(n3364), .B(n3363), .Z(\round_in[0][328] ) );
  NAND U9077 ( .A(init), .B(round_reg[329]), .Z(n3366) );
  NAND U9078 ( .A(n2806), .B(in[329]), .Z(n3365) );
  NAND U9079 ( .A(n3366), .B(n3365), .Z(\round_in[0][329] ) );
  NAND U9080 ( .A(init), .B(round_reg[32]), .Z(n3368) );
  NAND U9081 ( .A(n2806), .B(in[32]), .Z(n3367) );
  NAND U9082 ( .A(n3368), .B(n3367), .Z(\round_in[0][32] ) );
  NAND U9083 ( .A(init), .B(round_reg[330]), .Z(n3370) );
  NAND U9084 ( .A(n2806), .B(in[330]), .Z(n3369) );
  NAND U9085 ( .A(n3370), .B(n3369), .Z(\round_in[0][330] ) );
  NAND U9086 ( .A(init), .B(round_reg[331]), .Z(n3372) );
  NAND U9087 ( .A(n2807), .B(in[331]), .Z(n3371) );
  NAND U9088 ( .A(n3372), .B(n3371), .Z(\round_in[0][331] ) );
  NAND U9089 ( .A(init), .B(round_reg[332]), .Z(n3374) );
  NAND U9090 ( .A(n2807), .B(in[332]), .Z(n3373) );
  NAND U9091 ( .A(n3374), .B(n3373), .Z(\round_in[0][332] ) );
  NAND U9092 ( .A(init), .B(round_reg[333]), .Z(n3376) );
  NAND U9093 ( .A(n2807), .B(in[333]), .Z(n3375) );
  NAND U9094 ( .A(n3376), .B(n3375), .Z(\round_in[0][333] ) );
  NAND U9095 ( .A(init), .B(round_reg[334]), .Z(n3378) );
  NAND U9096 ( .A(n2807), .B(in[334]), .Z(n3377) );
  NAND U9097 ( .A(n3378), .B(n3377), .Z(\round_in[0][334] ) );
  NAND U9098 ( .A(init), .B(round_reg[335]), .Z(n3380) );
  NAND U9099 ( .A(n2807), .B(in[335]), .Z(n3379) );
  NAND U9100 ( .A(n3380), .B(n3379), .Z(\round_in[0][335] ) );
  NAND U9101 ( .A(init), .B(round_reg[336]), .Z(n3382) );
  NAND U9102 ( .A(n2807), .B(in[336]), .Z(n3381) );
  NAND U9103 ( .A(n3382), .B(n3381), .Z(\round_in[0][336] ) );
  NAND U9104 ( .A(init), .B(round_reg[337]), .Z(n3384) );
  NAND U9105 ( .A(n2807), .B(in[337]), .Z(n3383) );
  NAND U9106 ( .A(n3384), .B(n3383), .Z(\round_in[0][337] ) );
  NAND U9107 ( .A(init), .B(round_reg[338]), .Z(n3386) );
  NAND U9108 ( .A(n2808), .B(in[338]), .Z(n3385) );
  NAND U9109 ( .A(n3386), .B(n3385), .Z(\round_in[0][338] ) );
  NAND U9110 ( .A(init), .B(round_reg[339]), .Z(n3388) );
  NAND U9111 ( .A(n2808), .B(in[339]), .Z(n3387) );
  NAND U9112 ( .A(n3388), .B(n3387), .Z(\round_in[0][339] ) );
  NAND U9113 ( .A(init), .B(round_reg[33]), .Z(n3390) );
  NAND U9114 ( .A(n2808), .B(in[33]), .Z(n3389) );
  NAND U9115 ( .A(n3390), .B(n3389), .Z(\round_in[0][33] ) );
  NAND U9116 ( .A(init), .B(round_reg[340]), .Z(n3392) );
  NAND U9117 ( .A(n2808), .B(in[340]), .Z(n3391) );
  NAND U9118 ( .A(n3392), .B(n3391), .Z(\round_in[0][340] ) );
  NAND U9119 ( .A(init), .B(round_reg[341]), .Z(n3394) );
  NAND U9120 ( .A(n2808), .B(in[341]), .Z(n3393) );
  NAND U9121 ( .A(n3394), .B(n3393), .Z(\round_in[0][341] ) );
  NAND U9122 ( .A(init), .B(round_reg[342]), .Z(n3396) );
  NAND U9123 ( .A(n2808), .B(in[342]), .Z(n3395) );
  NAND U9124 ( .A(n3396), .B(n3395), .Z(\round_in[0][342] ) );
  NAND U9125 ( .A(init), .B(round_reg[343]), .Z(n3398) );
  NAND U9126 ( .A(n2808), .B(in[343]), .Z(n3397) );
  NAND U9127 ( .A(n3398), .B(n3397), .Z(\round_in[0][343] ) );
  NAND U9128 ( .A(init), .B(round_reg[344]), .Z(n3400) );
  NAND U9129 ( .A(n2809), .B(in[344]), .Z(n3399) );
  NAND U9130 ( .A(n3400), .B(n3399), .Z(\round_in[0][344] ) );
  NAND U9131 ( .A(init), .B(round_reg[345]), .Z(n3402) );
  NAND U9132 ( .A(n2809), .B(in[345]), .Z(n3401) );
  NAND U9133 ( .A(n3402), .B(n3401), .Z(\round_in[0][345] ) );
  NAND U9134 ( .A(init), .B(round_reg[346]), .Z(n3404) );
  NAND U9135 ( .A(n2809), .B(in[346]), .Z(n3403) );
  NAND U9136 ( .A(n3404), .B(n3403), .Z(\round_in[0][346] ) );
  NAND U9137 ( .A(init), .B(round_reg[347]), .Z(n3406) );
  NAND U9138 ( .A(n2809), .B(in[347]), .Z(n3405) );
  NAND U9139 ( .A(n3406), .B(n3405), .Z(\round_in[0][347] ) );
  NAND U9140 ( .A(init), .B(round_reg[348]), .Z(n3408) );
  NAND U9141 ( .A(n2809), .B(in[348]), .Z(n3407) );
  NAND U9142 ( .A(n3408), .B(n3407), .Z(\round_in[0][348] ) );
  NAND U9143 ( .A(init), .B(round_reg[349]), .Z(n3410) );
  NAND U9144 ( .A(n2809), .B(in[349]), .Z(n3409) );
  NAND U9145 ( .A(n3410), .B(n3409), .Z(\round_in[0][349] ) );
  NAND U9146 ( .A(init), .B(round_reg[34]), .Z(n3412) );
  NAND U9147 ( .A(n2809), .B(in[34]), .Z(n3411) );
  NAND U9148 ( .A(n3412), .B(n3411), .Z(\round_in[0][34] ) );
  NAND U9149 ( .A(init), .B(round_reg[350]), .Z(n3414) );
  NAND U9150 ( .A(n2810), .B(in[350]), .Z(n3413) );
  NAND U9151 ( .A(n3414), .B(n3413), .Z(\round_in[0][350] ) );
  NAND U9152 ( .A(init), .B(round_reg[351]), .Z(n3416) );
  NAND U9153 ( .A(n2810), .B(in[351]), .Z(n3415) );
  NAND U9154 ( .A(n3416), .B(n3415), .Z(\round_in[0][351] ) );
  NAND U9155 ( .A(init), .B(round_reg[352]), .Z(n3418) );
  NAND U9156 ( .A(n2810), .B(in[352]), .Z(n3417) );
  NAND U9157 ( .A(n3418), .B(n3417), .Z(\round_in[0][352] ) );
  NAND U9158 ( .A(init), .B(round_reg[353]), .Z(n3420) );
  NAND U9159 ( .A(n2810), .B(in[353]), .Z(n3419) );
  NAND U9160 ( .A(n3420), .B(n3419), .Z(\round_in[0][353] ) );
  NAND U9161 ( .A(init), .B(round_reg[354]), .Z(n3422) );
  NAND U9162 ( .A(n2810), .B(in[354]), .Z(n3421) );
  NAND U9163 ( .A(n3422), .B(n3421), .Z(\round_in[0][354] ) );
  NAND U9164 ( .A(init), .B(round_reg[355]), .Z(n3424) );
  NAND U9165 ( .A(n2810), .B(in[355]), .Z(n3423) );
  NAND U9166 ( .A(n3424), .B(n3423), .Z(\round_in[0][355] ) );
  NAND U9167 ( .A(init), .B(round_reg[356]), .Z(n3426) );
  NAND U9168 ( .A(n2810), .B(in[356]), .Z(n3425) );
  NAND U9169 ( .A(n3426), .B(n3425), .Z(\round_in[0][356] ) );
  NAND U9170 ( .A(init), .B(round_reg[357]), .Z(n3428) );
  NAND U9171 ( .A(n2811), .B(in[357]), .Z(n3427) );
  NAND U9172 ( .A(n3428), .B(n3427), .Z(\round_in[0][357] ) );
  NAND U9173 ( .A(init), .B(round_reg[358]), .Z(n3430) );
  NAND U9174 ( .A(n2811), .B(in[358]), .Z(n3429) );
  NAND U9175 ( .A(n3430), .B(n3429), .Z(\round_in[0][358] ) );
  NAND U9176 ( .A(init), .B(round_reg[359]), .Z(n3432) );
  NAND U9177 ( .A(n2811), .B(in[359]), .Z(n3431) );
  NAND U9178 ( .A(n3432), .B(n3431), .Z(\round_in[0][359] ) );
  NAND U9179 ( .A(init), .B(round_reg[35]), .Z(n3434) );
  NAND U9180 ( .A(n2811), .B(in[35]), .Z(n3433) );
  NAND U9181 ( .A(n3434), .B(n3433), .Z(\round_in[0][35] ) );
  NAND U9182 ( .A(init), .B(round_reg[360]), .Z(n3436) );
  NAND U9183 ( .A(n2811), .B(in[360]), .Z(n3435) );
  NAND U9184 ( .A(n3436), .B(n3435), .Z(\round_in[0][360] ) );
  NAND U9185 ( .A(init), .B(round_reg[361]), .Z(n3438) );
  NAND U9186 ( .A(n2811), .B(in[361]), .Z(n3437) );
  NAND U9187 ( .A(n3438), .B(n3437), .Z(\round_in[0][361] ) );
  NAND U9188 ( .A(init), .B(round_reg[362]), .Z(n3440) );
  NAND U9189 ( .A(n2811), .B(in[362]), .Z(n3439) );
  NAND U9190 ( .A(n3440), .B(n3439), .Z(\round_in[0][362] ) );
  NAND U9191 ( .A(init), .B(round_reg[363]), .Z(n3442) );
  NAND U9192 ( .A(n2812), .B(in[363]), .Z(n3441) );
  NAND U9193 ( .A(n3442), .B(n3441), .Z(\round_in[0][363] ) );
  NAND U9194 ( .A(init), .B(round_reg[364]), .Z(n3444) );
  NAND U9195 ( .A(n2812), .B(in[364]), .Z(n3443) );
  NAND U9196 ( .A(n3444), .B(n3443), .Z(\round_in[0][364] ) );
  NAND U9197 ( .A(init), .B(round_reg[365]), .Z(n3446) );
  NAND U9198 ( .A(n2812), .B(in[365]), .Z(n3445) );
  NAND U9199 ( .A(n3446), .B(n3445), .Z(\round_in[0][365] ) );
  NAND U9200 ( .A(init), .B(round_reg[366]), .Z(n3448) );
  NAND U9201 ( .A(n2812), .B(in[366]), .Z(n3447) );
  NAND U9202 ( .A(n3448), .B(n3447), .Z(\round_in[0][366] ) );
  NAND U9203 ( .A(init), .B(round_reg[367]), .Z(n3450) );
  NAND U9204 ( .A(n2812), .B(in[367]), .Z(n3449) );
  NAND U9205 ( .A(n3450), .B(n3449), .Z(\round_in[0][367] ) );
  NAND U9206 ( .A(init), .B(round_reg[368]), .Z(n3452) );
  NAND U9207 ( .A(n2812), .B(in[368]), .Z(n3451) );
  NAND U9208 ( .A(n3452), .B(n3451), .Z(\round_in[0][368] ) );
  NAND U9209 ( .A(init), .B(round_reg[369]), .Z(n3454) );
  NAND U9210 ( .A(n2812), .B(in[369]), .Z(n3453) );
  NAND U9211 ( .A(n3454), .B(n3453), .Z(\round_in[0][369] ) );
  NAND U9212 ( .A(init), .B(round_reg[36]), .Z(n3456) );
  NAND U9213 ( .A(n2813), .B(in[36]), .Z(n3455) );
  NAND U9214 ( .A(n3456), .B(n3455), .Z(\round_in[0][36] ) );
  NAND U9215 ( .A(init), .B(round_reg[370]), .Z(n3458) );
  NAND U9216 ( .A(n2813), .B(in[370]), .Z(n3457) );
  NAND U9217 ( .A(n3458), .B(n3457), .Z(\round_in[0][370] ) );
  NAND U9218 ( .A(init), .B(round_reg[371]), .Z(n3460) );
  NAND U9219 ( .A(n2813), .B(in[371]), .Z(n3459) );
  NAND U9220 ( .A(n3460), .B(n3459), .Z(\round_in[0][371] ) );
  NAND U9221 ( .A(init), .B(round_reg[372]), .Z(n3462) );
  NAND U9222 ( .A(n2813), .B(in[372]), .Z(n3461) );
  NAND U9223 ( .A(n3462), .B(n3461), .Z(\round_in[0][372] ) );
  NAND U9224 ( .A(init), .B(round_reg[373]), .Z(n3464) );
  NAND U9225 ( .A(n2813), .B(in[373]), .Z(n3463) );
  NAND U9226 ( .A(n3464), .B(n3463), .Z(\round_in[0][373] ) );
  NAND U9227 ( .A(init), .B(round_reg[374]), .Z(n3466) );
  NAND U9228 ( .A(n2813), .B(in[374]), .Z(n3465) );
  NAND U9229 ( .A(n3466), .B(n3465), .Z(\round_in[0][374] ) );
  NAND U9230 ( .A(init), .B(round_reg[375]), .Z(n3468) );
  NAND U9231 ( .A(n2813), .B(in[375]), .Z(n3467) );
  NAND U9232 ( .A(n3468), .B(n3467), .Z(\round_in[0][375] ) );
  NAND U9233 ( .A(init), .B(round_reg[376]), .Z(n3470) );
  NAND U9234 ( .A(n2814), .B(in[376]), .Z(n3469) );
  NAND U9235 ( .A(n3470), .B(n3469), .Z(\round_in[0][376] ) );
  NAND U9236 ( .A(init), .B(round_reg[377]), .Z(n3472) );
  NAND U9237 ( .A(n2814), .B(in[377]), .Z(n3471) );
  NAND U9238 ( .A(n3472), .B(n3471), .Z(\round_in[0][377] ) );
  NAND U9239 ( .A(init), .B(round_reg[378]), .Z(n3474) );
  NAND U9240 ( .A(n2814), .B(in[378]), .Z(n3473) );
  NAND U9241 ( .A(n3474), .B(n3473), .Z(\round_in[0][378] ) );
  NAND U9242 ( .A(init), .B(round_reg[379]), .Z(n3476) );
  NAND U9243 ( .A(n2814), .B(in[379]), .Z(n3475) );
  NAND U9244 ( .A(n3476), .B(n3475), .Z(\round_in[0][379] ) );
  NAND U9245 ( .A(init), .B(round_reg[37]), .Z(n3478) );
  NAND U9246 ( .A(n2814), .B(in[37]), .Z(n3477) );
  NAND U9247 ( .A(n3478), .B(n3477), .Z(\round_in[0][37] ) );
  NAND U9248 ( .A(init), .B(round_reg[380]), .Z(n3480) );
  NAND U9249 ( .A(n2814), .B(in[380]), .Z(n3479) );
  NAND U9250 ( .A(n3480), .B(n3479), .Z(\round_in[0][380] ) );
  NAND U9251 ( .A(init), .B(round_reg[381]), .Z(n3482) );
  NAND U9252 ( .A(n2814), .B(in[381]), .Z(n3481) );
  NAND U9253 ( .A(n3482), .B(n3481), .Z(\round_in[0][381] ) );
  NAND U9254 ( .A(init), .B(round_reg[382]), .Z(n3484) );
  NAND U9255 ( .A(n2815), .B(in[382]), .Z(n3483) );
  NAND U9256 ( .A(n3484), .B(n3483), .Z(\round_in[0][382] ) );
  NAND U9257 ( .A(init), .B(round_reg[383]), .Z(n3486) );
  NAND U9258 ( .A(n2815), .B(in[383]), .Z(n3485) );
  NAND U9259 ( .A(n3486), .B(n3485), .Z(\round_in[0][383] ) );
  NAND U9260 ( .A(init), .B(round_reg[384]), .Z(n3488) );
  NAND U9261 ( .A(n2815), .B(in[384]), .Z(n3487) );
  NAND U9262 ( .A(n3488), .B(n3487), .Z(\round_in[0][384] ) );
  NAND U9263 ( .A(init), .B(round_reg[385]), .Z(n3490) );
  NAND U9264 ( .A(n2815), .B(in[385]), .Z(n3489) );
  NAND U9265 ( .A(n3490), .B(n3489), .Z(\round_in[0][385] ) );
  NAND U9266 ( .A(init), .B(round_reg[386]), .Z(n3492) );
  NAND U9267 ( .A(n2815), .B(in[386]), .Z(n3491) );
  NAND U9268 ( .A(n3492), .B(n3491), .Z(\round_in[0][386] ) );
  NAND U9269 ( .A(init), .B(round_reg[387]), .Z(n3494) );
  NAND U9270 ( .A(n2815), .B(in[387]), .Z(n3493) );
  NAND U9271 ( .A(n3494), .B(n3493), .Z(\round_in[0][387] ) );
  NAND U9272 ( .A(init), .B(round_reg[388]), .Z(n3496) );
  NAND U9273 ( .A(n2815), .B(in[388]), .Z(n3495) );
  NAND U9274 ( .A(n3496), .B(n3495), .Z(\round_in[0][388] ) );
  NAND U9275 ( .A(init), .B(round_reg[389]), .Z(n3498) );
  NAND U9276 ( .A(n2816), .B(in[389]), .Z(n3497) );
  NAND U9277 ( .A(n3498), .B(n3497), .Z(\round_in[0][389] ) );
  NAND U9278 ( .A(init), .B(round_reg[38]), .Z(n3500) );
  NAND U9279 ( .A(n2816), .B(in[38]), .Z(n3499) );
  NAND U9280 ( .A(n3500), .B(n3499), .Z(\round_in[0][38] ) );
  NAND U9281 ( .A(init), .B(round_reg[390]), .Z(n3502) );
  NAND U9282 ( .A(n2816), .B(in[390]), .Z(n3501) );
  NAND U9283 ( .A(n3502), .B(n3501), .Z(\round_in[0][390] ) );
  NAND U9284 ( .A(init), .B(round_reg[391]), .Z(n3504) );
  NAND U9285 ( .A(n2816), .B(in[391]), .Z(n3503) );
  NAND U9286 ( .A(n3504), .B(n3503), .Z(\round_in[0][391] ) );
  NAND U9287 ( .A(init), .B(round_reg[392]), .Z(n3506) );
  NAND U9288 ( .A(n2816), .B(in[392]), .Z(n3505) );
  NAND U9289 ( .A(n3506), .B(n3505), .Z(\round_in[0][392] ) );
  NAND U9290 ( .A(init), .B(round_reg[393]), .Z(n3508) );
  NAND U9291 ( .A(n2816), .B(in[393]), .Z(n3507) );
  NAND U9292 ( .A(n3508), .B(n3507), .Z(\round_in[0][393] ) );
  NAND U9293 ( .A(init), .B(round_reg[394]), .Z(n3510) );
  NAND U9294 ( .A(n2816), .B(in[394]), .Z(n3509) );
  NAND U9295 ( .A(n3510), .B(n3509), .Z(\round_in[0][394] ) );
  NAND U9296 ( .A(init), .B(round_reg[395]), .Z(n3512) );
  NAND U9297 ( .A(n2817), .B(in[395]), .Z(n3511) );
  NAND U9298 ( .A(n3512), .B(n3511), .Z(\round_in[0][395] ) );
  NAND U9299 ( .A(init), .B(round_reg[396]), .Z(n3514) );
  NAND U9300 ( .A(n2817), .B(in[396]), .Z(n3513) );
  NAND U9301 ( .A(n3514), .B(n3513), .Z(\round_in[0][396] ) );
  NAND U9302 ( .A(init), .B(round_reg[397]), .Z(n3516) );
  NAND U9303 ( .A(n2817), .B(in[397]), .Z(n3515) );
  NAND U9304 ( .A(n3516), .B(n3515), .Z(\round_in[0][397] ) );
  NAND U9305 ( .A(init), .B(round_reg[398]), .Z(n3518) );
  NAND U9306 ( .A(n2817), .B(in[398]), .Z(n3517) );
  NAND U9307 ( .A(n3518), .B(n3517), .Z(\round_in[0][398] ) );
  NAND U9308 ( .A(init), .B(round_reg[399]), .Z(n3520) );
  NAND U9309 ( .A(n2817), .B(in[399]), .Z(n3519) );
  NAND U9310 ( .A(n3520), .B(n3519), .Z(\round_in[0][399] ) );
  NAND U9311 ( .A(init), .B(round_reg[39]), .Z(n3522) );
  NAND U9312 ( .A(n2817), .B(in[39]), .Z(n3521) );
  NAND U9313 ( .A(n3522), .B(n3521), .Z(\round_in[0][39] ) );
  NAND U9314 ( .A(init), .B(round_reg[3]), .Z(n3524) );
  NAND U9315 ( .A(n2817), .B(in[3]), .Z(n3523) );
  NAND U9316 ( .A(n3524), .B(n3523), .Z(\round_in[0][3] ) );
  NAND U9317 ( .A(init), .B(round_reg[400]), .Z(n3526) );
  NAND U9318 ( .A(n2818), .B(in[400]), .Z(n3525) );
  NAND U9319 ( .A(n3526), .B(n3525), .Z(\round_in[0][400] ) );
  NAND U9320 ( .A(init), .B(round_reg[401]), .Z(n3528) );
  NAND U9321 ( .A(n2818), .B(in[401]), .Z(n3527) );
  NAND U9322 ( .A(n3528), .B(n3527), .Z(\round_in[0][401] ) );
  NAND U9323 ( .A(init), .B(round_reg[402]), .Z(n3530) );
  NAND U9324 ( .A(n2818), .B(in[402]), .Z(n3529) );
  NAND U9325 ( .A(n3530), .B(n3529), .Z(\round_in[0][402] ) );
  NAND U9326 ( .A(init), .B(round_reg[403]), .Z(n3532) );
  NAND U9327 ( .A(n2818), .B(in[403]), .Z(n3531) );
  NAND U9328 ( .A(n3532), .B(n3531), .Z(\round_in[0][403] ) );
  NAND U9329 ( .A(init), .B(round_reg[404]), .Z(n3534) );
  NAND U9330 ( .A(n2818), .B(in[404]), .Z(n3533) );
  NAND U9331 ( .A(n3534), .B(n3533), .Z(\round_in[0][404] ) );
  NAND U9332 ( .A(init), .B(round_reg[405]), .Z(n3536) );
  NAND U9333 ( .A(n2818), .B(in[405]), .Z(n3535) );
  NAND U9334 ( .A(n3536), .B(n3535), .Z(\round_in[0][405] ) );
  NAND U9335 ( .A(init), .B(round_reg[406]), .Z(n3538) );
  NAND U9336 ( .A(n2818), .B(in[406]), .Z(n3537) );
  NAND U9337 ( .A(n3538), .B(n3537), .Z(\round_in[0][406] ) );
  NAND U9338 ( .A(init), .B(round_reg[407]), .Z(n3540) );
  NAND U9339 ( .A(n2819), .B(in[407]), .Z(n3539) );
  NAND U9340 ( .A(n3540), .B(n3539), .Z(\round_in[0][407] ) );
  NAND U9341 ( .A(init), .B(round_reg[408]), .Z(n3542) );
  NAND U9342 ( .A(n2819), .B(in[408]), .Z(n3541) );
  NAND U9343 ( .A(n3542), .B(n3541), .Z(\round_in[0][408] ) );
  NAND U9344 ( .A(init), .B(round_reg[409]), .Z(n3544) );
  NAND U9345 ( .A(n2819), .B(in[409]), .Z(n3543) );
  NAND U9346 ( .A(n3544), .B(n3543), .Z(\round_in[0][409] ) );
  NAND U9347 ( .A(init), .B(round_reg[40]), .Z(n3546) );
  NAND U9348 ( .A(n2819), .B(in[40]), .Z(n3545) );
  NAND U9349 ( .A(n3546), .B(n3545), .Z(\round_in[0][40] ) );
  NAND U9350 ( .A(init), .B(round_reg[410]), .Z(n3548) );
  NAND U9351 ( .A(n2819), .B(in[410]), .Z(n3547) );
  NAND U9352 ( .A(n3548), .B(n3547), .Z(\round_in[0][410] ) );
  NAND U9353 ( .A(init), .B(round_reg[411]), .Z(n3550) );
  NAND U9354 ( .A(n2819), .B(in[411]), .Z(n3549) );
  NAND U9355 ( .A(n3550), .B(n3549), .Z(\round_in[0][411] ) );
  NAND U9356 ( .A(init), .B(round_reg[412]), .Z(n3552) );
  NAND U9357 ( .A(n2819), .B(in[412]), .Z(n3551) );
  NAND U9358 ( .A(n3552), .B(n3551), .Z(\round_in[0][412] ) );
  NAND U9359 ( .A(init), .B(round_reg[413]), .Z(n3554) );
  NAND U9360 ( .A(n2820), .B(in[413]), .Z(n3553) );
  NAND U9361 ( .A(n3554), .B(n3553), .Z(\round_in[0][413] ) );
  NAND U9362 ( .A(init), .B(round_reg[414]), .Z(n3556) );
  NAND U9363 ( .A(n2820), .B(in[414]), .Z(n3555) );
  NAND U9364 ( .A(n3556), .B(n3555), .Z(\round_in[0][414] ) );
  NAND U9365 ( .A(init), .B(round_reg[415]), .Z(n3558) );
  NAND U9366 ( .A(n2820), .B(in[415]), .Z(n3557) );
  NAND U9367 ( .A(n3558), .B(n3557), .Z(\round_in[0][415] ) );
  NAND U9368 ( .A(init), .B(round_reg[416]), .Z(n3560) );
  NAND U9369 ( .A(n2820), .B(in[416]), .Z(n3559) );
  NAND U9370 ( .A(n3560), .B(n3559), .Z(\round_in[0][416] ) );
  NAND U9371 ( .A(init), .B(round_reg[417]), .Z(n3562) );
  NAND U9372 ( .A(n2820), .B(in[417]), .Z(n3561) );
  NAND U9373 ( .A(n3562), .B(n3561), .Z(\round_in[0][417] ) );
  NAND U9374 ( .A(init), .B(round_reg[418]), .Z(n3564) );
  NAND U9375 ( .A(n2820), .B(in[418]), .Z(n3563) );
  NAND U9376 ( .A(n3564), .B(n3563), .Z(\round_in[0][418] ) );
  NAND U9377 ( .A(init), .B(round_reg[419]), .Z(n3566) );
  NAND U9378 ( .A(n2820), .B(in[419]), .Z(n3565) );
  NAND U9379 ( .A(n3566), .B(n3565), .Z(\round_in[0][419] ) );
  NAND U9380 ( .A(init), .B(round_reg[41]), .Z(n3568) );
  NAND U9381 ( .A(n2821), .B(in[41]), .Z(n3567) );
  NAND U9382 ( .A(n3568), .B(n3567), .Z(\round_in[0][41] ) );
  NAND U9383 ( .A(init), .B(round_reg[420]), .Z(n3570) );
  NAND U9384 ( .A(n2821), .B(in[420]), .Z(n3569) );
  NAND U9385 ( .A(n3570), .B(n3569), .Z(\round_in[0][420] ) );
  NAND U9386 ( .A(init), .B(round_reg[421]), .Z(n3572) );
  NAND U9387 ( .A(n2821), .B(in[421]), .Z(n3571) );
  NAND U9388 ( .A(n3572), .B(n3571), .Z(\round_in[0][421] ) );
  NAND U9389 ( .A(init), .B(round_reg[422]), .Z(n3574) );
  NAND U9390 ( .A(n2821), .B(in[422]), .Z(n3573) );
  NAND U9391 ( .A(n3574), .B(n3573), .Z(\round_in[0][422] ) );
  NAND U9392 ( .A(init), .B(round_reg[423]), .Z(n3576) );
  NAND U9393 ( .A(n2821), .B(in[423]), .Z(n3575) );
  NAND U9394 ( .A(n3576), .B(n3575), .Z(\round_in[0][423] ) );
  NAND U9395 ( .A(init), .B(round_reg[424]), .Z(n3578) );
  NAND U9396 ( .A(n2821), .B(in[424]), .Z(n3577) );
  NAND U9397 ( .A(n3578), .B(n3577), .Z(\round_in[0][424] ) );
  NAND U9398 ( .A(init), .B(round_reg[425]), .Z(n3580) );
  NAND U9399 ( .A(n2821), .B(in[425]), .Z(n3579) );
  NAND U9400 ( .A(n3580), .B(n3579), .Z(\round_in[0][425] ) );
  NAND U9401 ( .A(init), .B(round_reg[426]), .Z(n3582) );
  NAND U9402 ( .A(n2822), .B(in[426]), .Z(n3581) );
  NAND U9403 ( .A(n3582), .B(n3581), .Z(\round_in[0][426] ) );
  NAND U9404 ( .A(init), .B(round_reg[427]), .Z(n3584) );
  NAND U9405 ( .A(n2822), .B(in[427]), .Z(n3583) );
  NAND U9406 ( .A(n3584), .B(n3583), .Z(\round_in[0][427] ) );
  NAND U9407 ( .A(init), .B(round_reg[428]), .Z(n3586) );
  NAND U9408 ( .A(n2822), .B(in[428]), .Z(n3585) );
  NAND U9409 ( .A(n3586), .B(n3585), .Z(\round_in[0][428] ) );
  NAND U9410 ( .A(init), .B(round_reg[429]), .Z(n3588) );
  NAND U9411 ( .A(n2822), .B(in[429]), .Z(n3587) );
  NAND U9412 ( .A(n3588), .B(n3587), .Z(\round_in[0][429] ) );
  NAND U9413 ( .A(init), .B(round_reg[42]), .Z(n3590) );
  NAND U9414 ( .A(n2822), .B(in[42]), .Z(n3589) );
  NAND U9415 ( .A(n3590), .B(n3589), .Z(\round_in[0][42] ) );
  NAND U9416 ( .A(init), .B(round_reg[430]), .Z(n3592) );
  NAND U9417 ( .A(n2822), .B(in[430]), .Z(n3591) );
  NAND U9418 ( .A(n3592), .B(n3591), .Z(\round_in[0][430] ) );
  NAND U9419 ( .A(init), .B(round_reg[431]), .Z(n3594) );
  NAND U9420 ( .A(n2822), .B(in[431]), .Z(n3593) );
  NAND U9421 ( .A(n3594), .B(n3593), .Z(\round_in[0][431] ) );
  NAND U9422 ( .A(init), .B(round_reg[432]), .Z(n3596) );
  NAND U9423 ( .A(n2823), .B(in[432]), .Z(n3595) );
  NAND U9424 ( .A(n3596), .B(n3595), .Z(\round_in[0][432] ) );
  NAND U9425 ( .A(init), .B(round_reg[433]), .Z(n3598) );
  NAND U9426 ( .A(n2823), .B(in[433]), .Z(n3597) );
  NAND U9427 ( .A(n3598), .B(n3597), .Z(\round_in[0][433] ) );
  NAND U9428 ( .A(init), .B(round_reg[434]), .Z(n3600) );
  NAND U9429 ( .A(n2823), .B(in[434]), .Z(n3599) );
  NAND U9430 ( .A(n3600), .B(n3599), .Z(\round_in[0][434] ) );
  NAND U9431 ( .A(init), .B(round_reg[435]), .Z(n3602) );
  NAND U9432 ( .A(n2823), .B(in[435]), .Z(n3601) );
  NAND U9433 ( .A(n3602), .B(n3601), .Z(\round_in[0][435] ) );
  NAND U9434 ( .A(init), .B(round_reg[436]), .Z(n3604) );
  NAND U9435 ( .A(n2823), .B(in[436]), .Z(n3603) );
  NAND U9436 ( .A(n3604), .B(n3603), .Z(\round_in[0][436] ) );
  NAND U9437 ( .A(init), .B(round_reg[437]), .Z(n3606) );
  NAND U9438 ( .A(n2823), .B(in[437]), .Z(n3605) );
  NAND U9439 ( .A(n3606), .B(n3605), .Z(\round_in[0][437] ) );
  NAND U9440 ( .A(init), .B(round_reg[438]), .Z(n3608) );
  NAND U9441 ( .A(n2823), .B(in[438]), .Z(n3607) );
  NAND U9442 ( .A(n3608), .B(n3607), .Z(\round_in[0][438] ) );
  NAND U9443 ( .A(init), .B(round_reg[439]), .Z(n3610) );
  NAND U9444 ( .A(n2824), .B(in[439]), .Z(n3609) );
  NAND U9445 ( .A(n3610), .B(n3609), .Z(\round_in[0][439] ) );
  NAND U9446 ( .A(init), .B(round_reg[43]), .Z(n3612) );
  NAND U9447 ( .A(n2824), .B(in[43]), .Z(n3611) );
  NAND U9448 ( .A(n3612), .B(n3611), .Z(\round_in[0][43] ) );
  NAND U9449 ( .A(init), .B(round_reg[440]), .Z(n3614) );
  NAND U9450 ( .A(n2824), .B(in[440]), .Z(n3613) );
  NAND U9451 ( .A(n3614), .B(n3613), .Z(\round_in[0][440] ) );
  NAND U9452 ( .A(init), .B(round_reg[441]), .Z(n3616) );
  NAND U9453 ( .A(n2824), .B(in[441]), .Z(n3615) );
  NAND U9454 ( .A(n3616), .B(n3615), .Z(\round_in[0][441] ) );
  NAND U9455 ( .A(init), .B(round_reg[442]), .Z(n3618) );
  NAND U9456 ( .A(n2824), .B(in[442]), .Z(n3617) );
  NAND U9457 ( .A(n3618), .B(n3617), .Z(\round_in[0][442] ) );
  NAND U9458 ( .A(init), .B(round_reg[443]), .Z(n3620) );
  NAND U9459 ( .A(n2824), .B(in[443]), .Z(n3619) );
  NAND U9460 ( .A(n3620), .B(n3619), .Z(\round_in[0][443] ) );
  NAND U9461 ( .A(init), .B(round_reg[444]), .Z(n3622) );
  NAND U9462 ( .A(n2824), .B(in[444]), .Z(n3621) );
  NAND U9463 ( .A(n3622), .B(n3621), .Z(\round_in[0][444] ) );
  NAND U9464 ( .A(init), .B(round_reg[445]), .Z(n3624) );
  NAND U9465 ( .A(n2825), .B(in[445]), .Z(n3623) );
  NAND U9466 ( .A(n3624), .B(n3623), .Z(\round_in[0][445] ) );
  NAND U9467 ( .A(init), .B(round_reg[446]), .Z(n3626) );
  NAND U9468 ( .A(n2825), .B(in[446]), .Z(n3625) );
  NAND U9469 ( .A(n3626), .B(n3625), .Z(\round_in[0][446] ) );
  NAND U9470 ( .A(init), .B(round_reg[447]), .Z(n3628) );
  NAND U9471 ( .A(n2825), .B(in[447]), .Z(n3627) );
  NAND U9472 ( .A(n3628), .B(n3627), .Z(\round_in[0][447] ) );
  NAND U9473 ( .A(init), .B(round_reg[448]), .Z(n3630) );
  NAND U9474 ( .A(n2825), .B(in[448]), .Z(n3629) );
  NAND U9475 ( .A(n3630), .B(n3629), .Z(\round_in[0][448] ) );
  NAND U9476 ( .A(init), .B(round_reg[449]), .Z(n3632) );
  NAND U9477 ( .A(n2825), .B(in[449]), .Z(n3631) );
  NAND U9478 ( .A(n3632), .B(n3631), .Z(\round_in[0][449] ) );
  NAND U9479 ( .A(init), .B(round_reg[44]), .Z(n3634) );
  NAND U9480 ( .A(n2825), .B(in[44]), .Z(n3633) );
  NAND U9481 ( .A(n3634), .B(n3633), .Z(\round_in[0][44] ) );
  NAND U9482 ( .A(init), .B(round_reg[450]), .Z(n3636) );
  NAND U9483 ( .A(n2825), .B(in[450]), .Z(n3635) );
  NAND U9484 ( .A(n3636), .B(n3635), .Z(\round_in[0][450] ) );
  NAND U9485 ( .A(init), .B(round_reg[451]), .Z(n3638) );
  NAND U9486 ( .A(n2826), .B(in[451]), .Z(n3637) );
  NAND U9487 ( .A(n3638), .B(n3637), .Z(\round_in[0][451] ) );
  NAND U9488 ( .A(init), .B(round_reg[452]), .Z(n3640) );
  NAND U9489 ( .A(n2826), .B(in[452]), .Z(n3639) );
  NAND U9490 ( .A(n3640), .B(n3639), .Z(\round_in[0][452] ) );
  NAND U9491 ( .A(init), .B(round_reg[453]), .Z(n3642) );
  NAND U9492 ( .A(n2826), .B(in[453]), .Z(n3641) );
  NAND U9493 ( .A(n3642), .B(n3641), .Z(\round_in[0][453] ) );
  NAND U9494 ( .A(init), .B(round_reg[454]), .Z(n3644) );
  NAND U9495 ( .A(n2826), .B(in[454]), .Z(n3643) );
  NAND U9496 ( .A(n3644), .B(n3643), .Z(\round_in[0][454] ) );
  NAND U9497 ( .A(init), .B(round_reg[455]), .Z(n3646) );
  NAND U9498 ( .A(n2826), .B(in[455]), .Z(n3645) );
  NAND U9499 ( .A(n3646), .B(n3645), .Z(\round_in[0][455] ) );
  NAND U9500 ( .A(init), .B(round_reg[456]), .Z(n3648) );
  NAND U9501 ( .A(n2826), .B(in[456]), .Z(n3647) );
  NAND U9502 ( .A(n3648), .B(n3647), .Z(\round_in[0][456] ) );
  NAND U9503 ( .A(init), .B(round_reg[457]), .Z(n3650) );
  NAND U9504 ( .A(n2826), .B(in[457]), .Z(n3649) );
  NAND U9505 ( .A(n3650), .B(n3649), .Z(\round_in[0][457] ) );
  NAND U9506 ( .A(init), .B(round_reg[458]), .Z(n3652) );
  NAND U9507 ( .A(n2827), .B(in[458]), .Z(n3651) );
  NAND U9508 ( .A(n3652), .B(n3651), .Z(\round_in[0][458] ) );
  NAND U9509 ( .A(init), .B(round_reg[459]), .Z(n3654) );
  NAND U9510 ( .A(n2827), .B(in[459]), .Z(n3653) );
  NAND U9511 ( .A(n3654), .B(n3653), .Z(\round_in[0][459] ) );
  NAND U9512 ( .A(init), .B(round_reg[45]), .Z(n3656) );
  NAND U9513 ( .A(n2827), .B(in[45]), .Z(n3655) );
  NAND U9514 ( .A(n3656), .B(n3655), .Z(\round_in[0][45] ) );
  NAND U9515 ( .A(init), .B(round_reg[460]), .Z(n3658) );
  NAND U9516 ( .A(n2827), .B(in[460]), .Z(n3657) );
  NAND U9517 ( .A(n3658), .B(n3657), .Z(\round_in[0][460] ) );
  NAND U9518 ( .A(init), .B(round_reg[461]), .Z(n3660) );
  NAND U9519 ( .A(n2827), .B(in[461]), .Z(n3659) );
  NAND U9520 ( .A(n3660), .B(n3659), .Z(\round_in[0][461] ) );
  NAND U9521 ( .A(init), .B(round_reg[462]), .Z(n3662) );
  NAND U9522 ( .A(n2827), .B(in[462]), .Z(n3661) );
  NAND U9523 ( .A(n3662), .B(n3661), .Z(\round_in[0][462] ) );
  NAND U9524 ( .A(init), .B(round_reg[463]), .Z(n3664) );
  NAND U9525 ( .A(n2827), .B(in[463]), .Z(n3663) );
  NAND U9526 ( .A(n3664), .B(n3663), .Z(\round_in[0][463] ) );
  NAND U9527 ( .A(init), .B(round_reg[464]), .Z(n3666) );
  NAND U9528 ( .A(n2828), .B(in[464]), .Z(n3665) );
  NAND U9529 ( .A(n3666), .B(n3665), .Z(\round_in[0][464] ) );
  NAND U9530 ( .A(init), .B(round_reg[465]), .Z(n3668) );
  NAND U9531 ( .A(n2828), .B(in[465]), .Z(n3667) );
  NAND U9532 ( .A(n3668), .B(n3667), .Z(\round_in[0][465] ) );
  NAND U9533 ( .A(init), .B(round_reg[466]), .Z(n3670) );
  NAND U9534 ( .A(n2828), .B(in[466]), .Z(n3669) );
  NAND U9535 ( .A(n3670), .B(n3669), .Z(\round_in[0][466] ) );
  NAND U9536 ( .A(init), .B(round_reg[467]), .Z(n3672) );
  NAND U9537 ( .A(n2828), .B(in[467]), .Z(n3671) );
  NAND U9538 ( .A(n3672), .B(n3671), .Z(\round_in[0][467] ) );
  NAND U9539 ( .A(init), .B(round_reg[468]), .Z(n3674) );
  NAND U9540 ( .A(n2828), .B(in[468]), .Z(n3673) );
  NAND U9541 ( .A(n3674), .B(n3673), .Z(\round_in[0][468] ) );
  NAND U9542 ( .A(init), .B(round_reg[469]), .Z(n3676) );
  NAND U9543 ( .A(n2828), .B(in[469]), .Z(n3675) );
  NAND U9544 ( .A(n3676), .B(n3675), .Z(\round_in[0][469] ) );
  NAND U9545 ( .A(init), .B(round_reg[46]), .Z(n3678) );
  NAND U9546 ( .A(n2828), .B(in[46]), .Z(n3677) );
  NAND U9547 ( .A(n3678), .B(n3677), .Z(\round_in[0][46] ) );
  NAND U9548 ( .A(init), .B(round_reg[470]), .Z(n3680) );
  NAND U9549 ( .A(n2829), .B(in[470]), .Z(n3679) );
  NAND U9550 ( .A(n3680), .B(n3679), .Z(\round_in[0][470] ) );
  NAND U9551 ( .A(init), .B(round_reg[471]), .Z(n3682) );
  NAND U9552 ( .A(n2829), .B(in[471]), .Z(n3681) );
  NAND U9553 ( .A(n3682), .B(n3681), .Z(\round_in[0][471] ) );
  NAND U9554 ( .A(init), .B(round_reg[472]), .Z(n3684) );
  NAND U9555 ( .A(n2829), .B(in[472]), .Z(n3683) );
  NAND U9556 ( .A(n3684), .B(n3683), .Z(\round_in[0][472] ) );
  NAND U9557 ( .A(init), .B(round_reg[473]), .Z(n3686) );
  NAND U9558 ( .A(n2829), .B(in[473]), .Z(n3685) );
  NAND U9559 ( .A(n3686), .B(n3685), .Z(\round_in[0][473] ) );
  NAND U9560 ( .A(init), .B(round_reg[474]), .Z(n3688) );
  NAND U9561 ( .A(n2829), .B(in[474]), .Z(n3687) );
  NAND U9562 ( .A(n3688), .B(n3687), .Z(\round_in[0][474] ) );
  NAND U9563 ( .A(init), .B(round_reg[475]), .Z(n3690) );
  NAND U9564 ( .A(n2829), .B(in[475]), .Z(n3689) );
  NAND U9565 ( .A(n3690), .B(n3689), .Z(\round_in[0][475] ) );
  NAND U9566 ( .A(init), .B(round_reg[476]), .Z(n3692) );
  NAND U9567 ( .A(n2829), .B(in[476]), .Z(n3691) );
  NAND U9568 ( .A(n3692), .B(n3691), .Z(\round_in[0][476] ) );
  NAND U9569 ( .A(init), .B(round_reg[477]), .Z(n3694) );
  NAND U9570 ( .A(n2830), .B(in[477]), .Z(n3693) );
  NAND U9571 ( .A(n3694), .B(n3693), .Z(\round_in[0][477] ) );
  NAND U9572 ( .A(init), .B(round_reg[478]), .Z(n3696) );
  NAND U9573 ( .A(n2830), .B(in[478]), .Z(n3695) );
  NAND U9574 ( .A(n3696), .B(n3695), .Z(\round_in[0][478] ) );
  NAND U9575 ( .A(init), .B(round_reg[479]), .Z(n3698) );
  NAND U9576 ( .A(n2830), .B(in[479]), .Z(n3697) );
  NAND U9577 ( .A(n3698), .B(n3697), .Z(\round_in[0][479] ) );
  NAND U9578 ( .A(init), .B(round_reg[47]), .Z(n3700) );
  NAND U9579 ( .A(n2830), .B(in[47]), .Z(n3699) );
  NAND U9580 ( .A(n3700), .B(n3699), .Z(\round_in[0][47] ) );
  NAND U9581 ( .A(init), .B(round_reg[480]), .Z(n3702) );
  NAND U9582 ( .A(n2830), .B(in[480]), .Z(n3701) );
  NAND U9583 ( .A(n3702), .B(n3701), .Z(\round_in[0][480] ) );
  NAND U9584 ( .A(init), .B(round_reg[481]), .Z(n3704) );
  NAND U9585 ( .A(n2830), .B(in[481]), .Z(n3703) );
  NAND U9586 ( .A(n3704), .B(n3703), .Z(\round_in[0][481] ) );
  NAND U9587 ( .A(init), .B(round_reg[482]), .Z(n3706) );
  NAND U9588 ( .A(n2830), .B(in[482]), .Z(n3705) );
  NAND U9589 ( .A(n3706), .B(n3705), .Z(\round_in[0][482] ) );
  NAND U9590 ( .A(init), .B(round_reg[483]), .Z(n3708) );
  NAND U9591 ( .A(n2831), .B(in[483]), .Z(n3707) );
  NAND U9592 ( .A(n3708), .B(n3707), .Z(\round_in[0][483] ) );
  NAND U9593 ( .A(init), .B(round_reg[484]), .Z(n3710) );
  NAND U9594 ( .A(n2831), .B(in[484]), .Z(n3709) );
  NAND U9595 ( .A(n3710), .B(n3709), .Z(\round_in[0][484] ) );
  NAND U9596 ( .A(init), .B(round_reg[485]), .Z(n3712) );
  NAND U9597 ( .A(n2831), .B(in[485]), .Z(n3711) );
  NAND U9598 ( .A(n3712), .B(n3711), .Z(\round_in[0][485] ) );
  NAND U9599 ( .A(init), .B(round_reg[486]), .Z(n3714) );
  NAND U9600 ( .A(n2831), .B(in[486]), .Z(n3713) );
  NAND U9601 ( .A(n3714), .B(n3713), .Z(\round_in[0][486] ) );
  NAND U9602 ( .A(init), .B(round_reg[487]), .Z(n3716) );
  NAND U9603 ( .A(n2831), .B(in[487]), .Z(n3715) );
  NAND U9604 ( .A(n3716), .B(n3715), .Z(\round_in[0][487] ) );
  NAND U9605 ( .A(init), .B(round_reg[488]), .Z(n3718) );
  NAND U9606 ( .A(n2831), .B(in[488]), .Z(n3717) );
  NAND U9607 ( .A(n3718), .B(n3717), .Z(\round_in[0][488] ) );
  NAND U9608 ( .A(init), .B(round_reg[489]), .Z(n3720) );
  NAND U9609 ( .A(n2831), .B(in[489]), .Z(n3719) );
  NAND U9610 ( .A(n3720), .B(n3719), .Z(\round_in[0][489] ) );
  NAND U9611 ( .A(init), .B(round_reg[48]), .Z(n3722) );
  NAND U9612 ( .A(n2832), .B(in[48]), .Z(n3721) );
  NAND U9613 ( .A(n3722), .B(n3721), .Z(\round_in[0][48] ) );
  NAND U9614 ( .A(init), .B(round_reg[490]), .Z(n3724) );
  NAND U9615 ( .A(n2832), .B(in[490]), .Z(n3723) );
  NAND U9616 ( .A(n3724), .B(n3723), .Z(\round_in[0][490] ) );
  NAND U9617 ( .A(init), .B(round_reg[491]), .Z(n3726) );
  NAND U9618 ( .A(n2832), .B(in[491]), .Z(n3725) );
  NAND U9619 ( .A(n3726), .B(n3725), .Z(\round_in[0][491] ) );
  NAND U9620 ( .A(init), .B(round_reg[492]), .Z(n3728) );
  NAND U9621 ( .A(n2832), .B(in[492]), .Z(n3727) );
  NAND U9622 ( .A(n3728), .B(n3727), .Z(\round_in[0][492] ) );
  NAND U9623 ( .A(init), .B(round_reg[493]), .Z(n3730) );
  NAND U9624 ( .A(n2832), .B(in[493]), .Z(n3729) );
  NAND U9625 ( .A(n3730), .B(n3729), .Z(\round_in[0][493] ) );
  NAND U9626 ( .A(init), .B(round_reg[494]), .Z(n3732) );
  NAND U9627 ( .A(n2832), .B(in[494]), .Z(n3731) );
  NAND U9628 ( .A(n3732), .B(n3731), .Z(\round_in[0][494] ) );
  NAND U9629 ( .A(init), .B(round_reg[495]), .Z(n3734) );
  NAND U9630 ( .A(n2832), .B(in[495]), .Z(n3733) );
  NAND U9631 ( .A(n3734), .B(n3733), .Z(\round_in[0][495] ) );
  NAND U9632 ( .A(init), .B(round_reg[496]), .Z(n3736) );
  NAND U9633 ( .A(n2833), .B(in[496]), .Z(n3735) );
  NAND U9634 ( .A(n3736), .B(n3735), .Z(\round_in[0][496] ) );
  NAND U9635 ( .A(init), .B(round_reg[497]), .Z(n3738) );
  NAND U9636 ( .A(n2833), .B(in[497]), .Z(n3737) );
  NAND U9637 ( .A(n3738), .B(n3737), .Z(\round_in[0][497] ) );
  NAND U9638 ( .A(init), .B(round_reg[498]), .Z(n3740) );
  NAND U9639 ( .A(n2833), .B(in[498]), .Z(n3739) );
  NAND U9640 ( .A(n3740), .B(n3739), .Z(\round_in[0][498] ) );
  NAND U9641 ( .A(init), .B(round_reg[499]), .Z(n3742) );
  NAND U9642 ( .A(n2833), .B(in[499]), .Z(n3741) );
  NAND U9643 ( .A(n3742), .B(n3741), .Z(\round_in[0][499] ) );
  NAND U9644 ( .A(init), .B(round_reg[49]), .Z(n3744) );
  NAND U9645 ( .A(n2833), .B(in[49]), .Z(n3743) );
  NAND U9646 ( .A(n3744), .B(n3743), .Z(\round_in[0][49] ) );
  NAND U9647 ( .A(init), .B(round_reg[4]), .Z(n3746) );
  NAND U9648 ( .A(n2833), .B(in[4]), .Z(n3745) );
  NAND U9649 ( .A(n3746), .B(n3745), .Z(\round_in[0][4] ) );
  NAND U9650 ( .A(init), .B(round_reg[500]), .Z(n3748) );
  NAND U9651 ( .A(n2833), .B(in[500]), .Z(n3747) );
  NAND U9652 ( .A(n3748), .B(n3747), .Z(\round_in[0][500] ) );
  NAND U9653 ( .A(init), .B(round_reg[501]), .Z(n3750) );
  NAND U9654 ( .A(n2834), .B(in[501]), .Z(n3749) );
  NAND U9655 ( .A(n3750), .B(n3749), .Z(\round_in[0][501] ) );
  NAND U9656 ( .A(init), .B(round_reg[502]), .Z(n3752) );
  NAND U9657 ( .A(n2834), .B(in[502]), .Z(n3751) );
  NAND U9658 ( .A(n3752), .B(n3751), .Z(\round_in[0][502] ) );
  NAND U9659 ( .A(init), .B(round_reg[503]), .Z(n3754) );
  NAND U9660 ( .A(n2834), .B(in[503]), .Z(n3753) );
  NAND U9661 ( .A(n3754), .B(n3753), .Z(\round_in[0][503] ) );
  NAND U9662 ( .A(init), .B(round_reg[504]), .Z(n3756) );
  NAND U9663 ( .A(n2834), .B(in[504]), .Z(n3755) );
  NAND U9664 ( .A(n3756), .B(n3755), .Z(\round_in[0][504] ) );
  NAND U9665 ( .A(init), .B(round_reg[505]), .Z(n3758) );
  NAND U9666 ( .A(n2834), .B(in[505]), .Z(n3757) );
  NAND U9667 ( .A(n3758), .B(n3757), .Z(\round_in[0][505] ) );
  NAND U9668 ( .A(init), .B(round_reg[506]), .Z(n3760) );
  NAND U9669 ( .A(n2834), .B(in[506]), .Z(n3759) );
  NAND U9670 ( .A(n3760), .B(n3759), .Z(\round_in[0][506] ) );
  NAND U9671 ( .A(init), .B(round_reg[507]), .Z(n3762) );
  NAND U9672 ( .A(n2834), .B(in[507]), .Z(n3761) );
  NAND U9673 ( .A(n3762), .B(n3761), .Z(\round_in[0][507] ) );
  NAND U9674 ( .A(init), .B(round_reg[508]), .Z(n3764) );
  NAND U9675 ( .A(n2835), .B(in[508]), .Z(n3763) );
  NAND U9676 ( .A(n3764), .B(n3763), .Z(\round_in[0][508] ) );
  NAND U9677 ( .A(init), .B(round_reg[509]), .Z(n3766) );
  NAND U9678 ( .A(n2835), .B(in[509]), .Z(n3765) );
  NAND U9679 ( .A(n3766), .B(n3765), .Z(\round_in[0][509] ) );
  NAND U9680 ( .A(init), .B(round_reg[50]), .Z(n3768) );
  NAND U9681 ( .A(n2835), .B(in[50]), .Z(n3767) );
  NAND U9682 ( .A(n3768), .B(n3767), .Z(\round_in[0][50] ) );
  NAND U9683 ( .A(init), .B(round_reg[510]), .Z(n3770) );
  NAND U9684 ( .A(n2835), .B(in[510]), .Z(n3769) );
  NAND U9685 ( .A(n3770), .B(n3769), .Z(\round_in[0][510] ) );
  NAND U9686 ( .A(init), .B(round_reg[511]), .Z(n3772) );
  NAND U9687 ( .A(n2835), .B(in[511]), .Z(n3771) );
  NAND U9688 ( .A(n3772), .B(n3771), .Z(\round_in[0][511] ) );
  NAND U9689 ( .A(init), .B(round_reg[512]), .Z(n3774) );
  NAND U9690 ( .A(n2835), .B(in[512]), .Z(n3773) );
  NAND U9691 ( .A(n3774), .B(n3773), .Z(\round_in[0][512] ) );
  NAND U9692 ( .A(init), .B(round_reg[513]), .Z(n3776) );
  NAND U9693 ( .A(n2835), .B(in[513]), .Z(n3775) );
  NAND U9694 ( .A(n3776), .B(n3775), .Z(\round_in[0][513] ) );
  NAND U9695 ( .A(init), .B(round_reg[514]), .Z(n3778) );
  NAND U9696 ( .A(n2836), .B(in[514]), .Z(n3777) );
  NAND U9697 ( .A(n3778), .B(n3777), .Z(\round_in[0][514] ) );
  NAND U9698 ( .A(init), .B(round_reg[515]), .Z(n3780) );
  NAND U9699 ( .A(n2836), .B(in[515]), .Z(n3779) );
  NAND U9700 ( .A(n3780), .B(n3779), .Z(\round_in[0][515] ) );
  NAND U9701 ( .A(init), .B(round_reg[516]), .Z(n3782) );
  NAND U9702 ( .A(n2836), .B(in[516]), .Z(n3781) );
  NAND U9703 ( .A(n3782), .B(n3781), .Z(\round_in[0][516] ) );
  NAND U9704 ( .A(init), .B(round_reg[517]), .Z(n3784) );
  NAND U9705 ( .A(n2836), .B(in[517]), .Z(n3783) );
  NAND U9706 ( .A(n3784), .B(n3783), .Z(\round_in[0][517] ) );
  NAND U9707 ( .A(init), .B(round_reg[518]), .Z(n3786) );
  NAND U9708 ( .A(n2836), .B(in[518]), .Z(n3785) );
  NAND U9709 ( .A(n3786), .B(n3785), .Z(\round_in[0][518] ) );
  NAND U9710 ( .A(init), .B(round_reg[519]), .Z(n3788) );
  NAND U9711 ( .A(n2836), .B(in[519]), .Z(n3787) );
  NAND U9712 ( .A(n3788), .B(n3787), .Z(\round_in[0][519] ) );
  NAND U9713 ( .A(init), .B(round_reg[51]), .Z(n3790) );
  NAND U9714 ( .A(n2836), .B(in[51]), .Z(n3789) );
  NAND U9715 ( .A(n3790), .B(n3789), .Z(\round_in[0][51] ) );
  NAND U9716 ( .A(init), .B(round_reg[520]), .Z(n3792) );
  NAND U9717 ( .A(n2837), .B(in[520]), .Z(n3791) );
  NAND U9718 ( .A(n3792), .B(n3791), .Z(\round_in[0][520] ) );
  NAND U9719 ( .A(init), .B(round_reg[521]), .Z(n3794) );
  NAND U9720 ( .A(n2837), .B(in[521]), .Z(n3793) );
  NAND U9721 ( .A(n3794), .B(n3793), .Z(\round_in[0][521] ) );
  NAND U9722 ( .A(init), .B(round_reg[522]), .Z(n3796) );
  NAND U9723 ( .A(n2837), .B(in[522]), .Z(n3795) );
  NAND U9724 ( .A(n3796), .B(n3795), .Z(\round_in[0][522] ) );
  NAND U9725 ( .A(init), .B(round_reg[523]), .Z(n3798) );
  NAND U9726 ( .A(n2837), .B(in[523]), .Z(n3797) );
  NAND U9727 ( .A(n3798), .B(n3797), .Z(\round_in[0][523] ) );
  NAND U9728 ( .A(init), .B(round_reg[524]), .Z(n3800) );
  NAND U9729 ( .A(n2837), .B(in[524]), .Z(n3799) );
  NAND U9730 ( .A(n3800), .B(n3799), .Z(\round_in[0][524] ) );
  NAND U9731 ( .A(init), .B(round_reg[525]), .Z(n3802) );
  NAND U9732 ( .A(n2837), .B(in[525]), .Z(n3801) );
  NAND U9733 ( .A(n3802), .B(n3801), .Z(\round_in[0][525] ) );
  NAND U9734 ( .A(init), .B(round_reg[526]), .Z(n3804) );
  NAND U9735 ( .A(n2837), .B(in[526]), .Z(n3803) );
  NAND U9736 ( .A(n3804), .B(n3803), .Z(\round_in[0][526] ) );
  NAND U9737 ( .A(init), .B(round_reg[527]), .Z(n3806) );
  NAND U9738 ( .A(n2838), .B(in[527]), .Z(n3805) );
  NAND U9739 ( .A(n3806), .B(n3805), .Z(\round_in[0][527] ) );
  NAND U9740 ( .A(init), .B(round_reg[528]), .Z(n3808) );
  NAND U9741 ( .A(n2838), .B(in[528]), .Z(n3807) );
  NAND U9742 ( .A(n3808), .B(n3807), .Z(\round_in[0][528] ) );
  NAND U9743 ( .A(init), .B(round_reg[529]), .Z(n3810) );
  NAND U9744 ( .A(n2838), .B(in[529]), .Z(n3809) );
  NAND U9745 ( .A(n3810), .B(n3809), .Z(\round_in[0][529] ) );
  NAND U9746 ( .A(init), .B(round_reg[52]), .Z(n3812) );
  NAND U9747 ( .A(n2838), .B(in[52]), .Z(n3811) );
  NAND U9748 ( .A(n3812), .B(n3811), .Z(\round_in[0][52] ) );
  NAND U9749 ( .A(init), .B(round_reg[530]), .Z(n3814) );
  NAND U9750 ( .A(n2838), .B(in[530]), .Z(n3813) );
  NAND U9751 ( .A(n3814), .B(n3813), .Z(\round_in[0][530] ) );
  NAND U9752 ( .A(init), .B(round_reg[531]), .Z(n3816) );
  NAND U9753 ( .A(n2838), .B(in[531]), .Z(n3815) );
  NAND U9754 ( .A(n3816), .B(n3815), .Z(\round_in[0][531] ) );
  NAND U9755 ( .A(init), .B(round_reg[532]), .Z(n3818) );
  NAND U9756 ( .A(n2838), .B(in[532]), .Z(n3817) );
  NAND U9757 ( .A(n3818), .B(n3817), .Z(\round_in[0][532] ) );
  NAND U9758 ( .A(init), .B(round_reg[533]), .Z(n3820) );
  NAND U9759 ( .A(n2839), .B(in[533]), .Z(n3819) );
  NAND U9760 ( .A(n3820), .B(n3819), .Z(\round_in[0][533] ) );
  NAND U9761 ( .A(init), .B(round_reg[534]), .Z(n3822) );
  NAND U9762 ( .A(n2839), .B(in[534]), .Z(n3821) );
  NAND U9763 ( .A(n3822), .B(n3821), .Z(\round_in[0][534] ) );
  NAND U9764 ( .A(init), .B(round_reg[535]), .Z(n3824) );
  NAND U9765 ( .A(n2839), .B(in[535]), .Z(n3823) );
  NAND U9766 ( .A(n3824), .B(n3823), .Z(\round_in[0][535] ) );
  NAND U9767 ( .A(init), .B(round_reg[536]), .Z(n3826) );
  NAND U9768 ( .A(n2839), .B(in[536]), .Z(n3825) );
  NAND U9769 ( .A(n3826), .B(n3825), .Z(\round_in[0][536] ) );
  NAND U9770 ( .A(init), .B(round_reg[537]), .Z(n3828) );
  NAND U9771 ( .A(n2839), .B(in[537]), .Z(n3827) );
  NAND U9772 ( .A(n3828), .B(n3827), .Z(\round_in[0][537] ) );
  NAND U9773 ( .A(init), .B(round_reg[538]), .Z(n3830) );
  NAND U9774 ( .A(n2839), .B(in[538]), .Z(n3829) );
  NAND U9775 ( .A(n3830), .B(n3829), .Z(\round_in[0][538] ) );
  NAND U9776 ( .A(init), .B(round_reg[539]), .Z(n3832) );
  NAND U9777 ( .A(n2839), .B(in[539]), .Z(n3831) );
  NAND U9778 ( .A(n3832), .B(n3831), .Z(\round_in[0][539] ) );
  NAND U9779 ( .A(init), .B(round_reg[53]), .Z(n3834) );
  NAND U9780 ( .A(n2840), .B(in[53]), .Z(n3833) );
  NAND U9781 ( .A(n3834), .B(n3833), .Z(\round_in[0][53] ) );
  NAND U9782 ( .A(init), .B(round_reg[540]), .Z(n3836) );
  NAND U9783 ( .A(n2840), .B(in[540]), .Z(n3835) );
  NAND U9784 ( .A(n3836), .B(n3835), .Z(\round_in[0][540] ) );
  NAND U9785 ( .A(init), .B(round_reg[541]), .Z(n3838) );
  NAND U9786 ( .A(n2840), .B(in[541]), .Z(n3837) );
  NAND U9787 ( .A(n3838), .B(n3837), .Z(\round_in[0][541] ) );
  NAND U9788 ( .A(init), .B(round_reg[542]), .Z(n3840) );
  NAND U9789 ( .A(n2840), .B(in[542]), .Z(n3839) );
  NAND U9790 ( .A(n3840), .B(n3839), .Z(\round_in[0][542] ) );
  NAND U9791 ( .A(init), .B(round_reg[543]), .Z(n3842) );
  NAND U9792 ( .A(n2840), .B(in[543]), .Z(n3841) );
  NAND U9793 ( .A(n3842), .B(n3841), .Z(\round_in[0][543] ) );
  NAND U9794 ( .A(init), .B(round_reg[544]), .Z(n3844) );
  NAND U9795 ( .A(n2840), .B(in[544]), .Z(n3843) );
  NAND U9796 ( .A(n3844), .B(n3843), .Z(\round_in[0][544] ) );
  NAND U9797 ( .A(init), .B(round_reg[545]), .Z(n3846) );
  NAND U9798 ( .A(n2840), .B(in[545]), .Z(n3845) );
  NAND U9799 ( .A(n3846), .B(n3845), .Z(\round_in[0][545] ) );
  NAND U9800 ( .A(init), .B(round_reg[546]), .Z(n3848) );
  NAND U9801 ( .A(n2841), .B(in[546]), .Z(n3847) );
  NAND U9802 ( .A(n3848), .B(n3847), .Z(\round_in[0][546] ) );
  NAND U9803 ( .A(init), .B(round_reg[547]), .Z(n3850) );
  NAND U9804 ( .A(n2841), .B(in[547]), .Z(n3849) );
  NAND U9805 ( .A(n3850), .B(n3849), .Z(\round_in[0][547] ) );
  NAND U9806 ( .A(init), .B(round_reg[548]), .Z(n3852) );
  NAND U9807 ( .A(n2841), .B(in[548]), .Z(n3851) );
  NAND U9808 ( .A(n3852), .B(n3851), .Z(\round_in[0][548] ) );
  NAND U9809 ( .A(init), .B(round_reg[549]), .Z(n3854) );
  NAND U9810 ( .A(n2841), .B(in[549]), .Z(n3853) );
  NAND U9811 ( .A(n3854), .B(n3853), .Z(\round_in[0][549] ) );
  NAND U9812 ( .A(init), .B(round_reg[54]), .Z(n3856) );
  NAND U9813 ( .A(n2841), .B(in[54]), .Z(n3855) );
  NAND U9814 ( .A(n3856), .B(n3855), .Z(\round_in[0][54] ) );
  NAND U9815 ( .A(init), .B(round_reg[550]), .Z(n3858) );
  NAND U9816 ( .A(n2841), .B(in[550]), .Z(n3857) );
  NAND U9817 ( .A(n3858), .B(n3857), .Z(\round_in[0][550] ) );
  NAND U9818 ( .A(init), .B(round_reg[551]), .Z(n3860) );
  NAND U9819 ( .A(n2841), .B(in[551]), .Z(n3859) );
  NAND U9820 ( .A(n3860), .B(n3859), .Z(\round_in[0][551] ) );
  NAND U9821 ( .A(init), .B(round_reg[552]), .Z(n3862) );
  NAND U9822 ( .A(n2842), .B(in[552]), .Z(n3861) );
  NAND U9823 ( .A(n3862), .B(n3861), .Z(\round_in[0][552] ) );
  NAND U9824 ( .A(init), .B(round_reg[553]), .Z(n3864) );
  NAND U9825 ( .A(n2842), .B(in[553]), .Z(n3863) );
  NAND U9826 ( .A(n3864), .B(n3863), .Z(\round_in[0][553] ) );
  NAND U9827 ( .A(init), .B(round_reg[554]), .Z(n3866) );
  NAND U9828 ( .A(n2842), .B(in[554]), .Z(n3865) );
  NAND U9829 ( .A(n3866), .B(n3865), .Z(\round_in[0][554] ) );
  NAND U9830 ( .A(init), .B(round_reg[555]), .Z(n3868) );
  NAND U9831 ( .A(n2842), .B(in[555]), .Z(n3867) );
  NAND U9832 ( .A(n3868), .B(n3867), .Z(\round_in[0][555] ) );
  NAND U9833 ( .A(init), .B(round_reg[556]), .Z(n3870) );
  NAND U9834 ( .A(n2842), .B(in[556]), .Z(n3869) );
  NAND U9835 ( .A(n3870), .B(n3869), .Z(\round_in[0][556] ) );
  NAND U9836 ( .A(init), .B(round_reg[557]), .Z(n3872) );
  NAND U9837 ( .A(n2842), .B(in[557]), .Z(n3871) );
  NAND U9838 ( .A(n3872), .B(n3871), .Z(\round_in[0][557] ) );
  NAND U9839 ( .A(init), .B(round_reg[558]), .Z(n3874) );
  NAND U9840 ( .A(n2842), .B(in[558]), .Z(n3873) );
  NAND U9841 ( .A(n3874), .B(n3873), .Z(\round_in[0][558] ) );
  NAND U9842 ( .A(init), .B(round_reg[559]), .Z(n3876) );
  NAND U9843 ( .A(n2843), .B(in[559]), .Z(n3875) );
  NAND U9844 ( .A(n3876), .B(n3875), .Z(\round_in[0][559] ) );
  NAND U9845 ( .A(init), .B(round_reg[55]), .Z(n3878) );
  NAND U9846 ( .A(n2843), .B(in[55]), .Z(n3877) );
  NAND U9847 ( .A(n3878), .B(n3877), .Z(\round_in[0][55] ) );
  NAND U9848 ( .A(init), .B(round_reg[560]), .Z(n3880) );
  NAND U9849 ( .A(n2843), .B(in[560]), .Z(n3879) );
  NAND U9850 ( .A(n3880), .B(n3879), .Z(\round_in[0][560] ) );
  NAND U9851 ( .A(init), .B(round_reg[561]), .Z(n3882) );
  NAND U9852 ( .A(n2843), .B(in[561]), .Z(n3881) );
  NAND U9853 ( .A(n3882), .B(n3881), .Z(\round_in[0][561] ) );
  NAND U9854 ( .A(init), .B(round_reg[562]), .Z(n3884) );
  NAND U9855 ( .A(n2843), .B(in[562]), .Z(n3883) );
  NAND U9856 ( .A(n3884), .B(n3883), .Z(\round_in[0][562] ) );
  NAND U9857 ( .A(init), .B(round_reg[563]), .Z(n3886) );
  NAND U9858 ( .A(n2843), .B(in[563]), .Z(n3885) );
  NAND U9859 ( .A(n3886), .B(n3885), .Z(\round_in[0][563] ) );
  NAND U9860 ( .A(init), .B(round_reg[564]), .Z(n3888) );
  NAND U9861 ( .A(n2843), .B(in[564]), .Z(n3887) );
  NAND U9862 ( .A(n3888), .B(n3887), .Z(\round_in[0][564] ) );
  NAND U9863 ( .A(init), .B(round_reg[565]), .Z(n3890) );
  NAND U9864 ( .A(n2844), .B(in[565]), .Z(n3889) );
  NAND U9865 ( .A(n3890), .B(n3889), .Z(\round_in[0][565] ) );
  NAND U9866 ( .A(init), .B(round_reg[566]), .Z(n3892) );
  NAND U9867 ( .A(n2844), .B(in[566]), .Z(n3891) );
  NAND U9868 ( .A(n3892), .B(n3891), .Z(\round_in[0][566] ) );
  NAND U9869 ( .A(init), .B(round_reg[567]), .Z(n3894) );
  NAND U9870 ( .A(n2844), .B(in[567]), .Z(n3893) );
  NAND U9871 ( .A(n3894), .B(n3893), .Z(\round_in[0][567] ) );
  NAND U9872 ( .A(init), .B(round_reg[568]), .Z(n3896) );
  NAND U9873 ( .A(n2844), .B(in[568]), .Z(n3895) );
  NAND U9874 ( .A(n3896), .B(n3895), .Z(\round_in[0][568] ) );
  NAND U9875 ( .A(init), .B(round_reg[569]), .Z(n3898) );
  NAND U9876 ( .A(n2844), .B(in[569]), .Z(n3897) );
  NAND U9877 ( .A(n3898), .B(n3897), .Z(\round_in[0][569] ) );
  NAND U9878 ( .A(init), .B(round_reg[56]), .Z(n3900) );
  NAND U9879 ( .A(n2844), .B(in[56]), .Z(n3899) );
  NAND U9880 ( .A(n3900), .B(n3899), .Z(\round_in[0][56] ) );
  NAND U9881 ( .A(init), .B(round_reg[570]), .Z(n3902) );
  NAND U9882 ( .A(n2844), .B(in[570]), .Z(n3901) );
  NAND U9883 ( .A(n3902), .B(n3901), .Z(\round_in[0][570] ) );
  NAND U9884 ( .A(init), .B(round_reg[571]), .Z(n3904) );
  NAND U9885 ( .A(n2845), .B(in[571]), .Z(n3903) );
  NAND U9886 ( .A(n3904), .B(n3903), .Z(\round_in[0][571] ) );
  NAND U9887 ( .A(init), .B(round_reg[572]), .Z(n3906) );
  NAND U9888 ( .A(n2845), .B(in[572]), .Z(n3905) );
  NAND U9889 ( .A(n3906), .B(n3905), .Z(\round_in[0][572] ) );
  NAND U9890 ( .A(init), .B(round_reg[573]), .Z(n3908) );
  NAND U9891 ( .A(n2845), .B(in[573]), .Z(n3907) );
  NAND U9892 ( .A(n3908), .B(n3907), .Z(\round_in[0][573] ) );
  NAND U9893 ( .A(init), .B(round_reg[574]), .Z(n3910) );
  NAND U9894 ( .A(n2845), .B(in[574]), .Z(n3909) );
  NAND U9895 ( .A(n3910), .B(n3909), .Z(\round_in[0][574] ) );
  NAND U9896 ( .A(init), .B(round_reg[575]), .Z(n3912) );
  NAND U9897 ( .A(n2845), .B(in[575]), .Z(n3911) );
  NAND U9898 ( .A(n3912), .B(n3911), .Z(\round_in[0][575] ) );
  AND U9899 ( .A(round_reg[576]), .B(init), .Z(\round_in[0][576] ) );
  AND U9900 ( .A(round_reg[577]), .B(init), .Z(\round_in[0][577] ) );
  AND U9901 ( .A(round_reg[578]), .B(init), .Z(\round_in[0][578] ) );
  AND U9902 ( .A(round_reg[579]), .B(init), .Z(\round_in[0][579] ) );
  NAND U9903 ( .A(init), .B(round_reg[57]), .Z(n3914) );
  NAND U9904 ( .A(n2845), .B(in[57]), .Z(n3913) );
  NAND U9905 ( .A(n3914), .B(n3913), .Z(\round_in[0][57] ) );
  AND U9906 ( .A(round_reg[580]), .B(init), .Z(\round_in[0][580] ) );
  AND U9907 ( .A(round_reg[581]), .B(init), .Z(\round_in[0][581] ) );
  AND U9908 ( .A(round_reg[582]), .B(init), .Z(\round_in[0][582] ) );
  AND U9909 ( .A(round_reg[583]), .B(init), .Z(\round_in[0][583] ) );
  AND U9910 ( .A(round_reg[584]), .B(init), .Z(\round_in[0][584] ) );
  AND U9911 ( .A(round_reg[585]), .B(init), .Z(\round_in[0][585] ) );
  AND U9912 ( .A(round_reg[586]), .B(init), .Z(\round_in[0][586] ) );
  AND U9913 ( .A(round_reg[587]), .B(init), .Z(\round_in[0][587] ) );
  AND U9914 ( .A(round_reg[588]), .B(init), .Z(\round_in[0][588] ) );
  AND U9915 ( .A(round_reg[589]), .B(init), .Z(\round_in[0][589] ) );
  NAND U9916 ( .A(init), .B(round_reg[58]), .Z(n3916) );
  NAND U9917 ( .A(n2845), .B(in[58]), .Z(n3915) );
  NAND U9918 ( .A(n3916), .B(n3915), .Z(\round_in[0][58] ) );
  AND U9919 ( .A(round_reg[590]), .B(init), .Z(\round_in[0][590] ) );
  AND U9920 ( .A(round_reg[591]), .B(init), .Z(\round_in[0][591] ) );
  AND U9921 ( .A(round_reg[592]), .B(init), .Z(\round_in[0][592] ) );
  AND U9922 ( .A(round_reg[593]), .B(init), .Z(\round_in[0][593] ) );
  AND U9923 ( .A(round_reg[594]), .B(init), .Z(\round_in[0][594] ) );
  AND U9924 ( .A(round_reg[595]), .B(init), .Z(\round_in[0][595] ) );
  AND U9925 ( .A(round_reg[596]), .B(init), .Z(\round_in[0][596] ) );
  AND U9926 ( .A(round_reg[597]), .B(init), .Z(\round_in[0][597] ) );
  AND U9927 ( .A(round_reg[598]), .B(init), .Z(\round_in[0][598] ) );
  AND U9928 ( .A(round_reg[599]), .B(init), .Z(\round_in[0][599] ) );
  NAND U9929 ( .A(init), .B(round_reg[59]), .Z(n3918) );
  NAND U9930 ( .A(n2846), .B(in[59]), .Z(n3917) );
  NAND U9931 ( .A(n3918), .B(n3917), .Z(\round_in[0][59] ) );
  NAND U9932 ( .A(init), .B(round_reg[5]), .Z(n3920) );
  NAND U9933 ( .A(n2846), .B(in[5]), .Z(n3919) );
  NAND U9934 ( .A(n3920), .B(n3919), .Z(\round_in[0][5] ) );
  AND U9935 ( .A(round_reg[600]), .B(init), .Z(\round_in[0][600] ) );
  AND U9936 ( .A(round_reg[601]), .B(init), .Z(\round_in[0][601] ) );
  AND U9937 ( .A(round_reg[602]), .B(init), .Z(\round_in[0][602] ) );
  AND U9938 ( .A(round_reg[603]), .B(init), .Z(\round_in[0][603] ) );
  AND U9939 ( .A(round_reg[604]), .B(init), .Z(\round_in[0][604] ) );
  AND U9940 ( .A(round_reg[605]), .B(init), .Z(\round_in[0][605] ) );
  AND U9941 ( .A(round_reg[606]), .B(init), .Z(\round_in[0][606] ) );
  AND U9942 ( .A(round_reg[607]), .B(init), .Z(\round_in[0][607] ) );
  AND U9943 ( .A(round_reg[608]), .B(init), .Z(\round_in[0][608] ) );
  AND U9944 ( .A(round_reg[609]), .B(init), .Z(\round_in[0][609] ) );
  NAND U9945 ( .A(init), .B(round_reg[60]), .Z(n3922) );
  NAND U9946 ( .A(n2846), .B(in[60]), .Z(n3921) );
  NAND U9947 ( .A(n3922), .B(n3921), .Z(\round_in[0][60] ) );
  AND U9948 ( .A(round_reg[610]), .B(init), .Z(\round_in[0][610] ) );
  AND U9949 ( .A(round_reg[611]), .B(init), .Z(\round_in[0][611] ) );
  AND U9950 ( .A(round_reg[612]), .B(init), .Z(\round_in[0][612] ) );
  AND U9951 ( .A(round_reg[613]), .B(init), .Z(\round_in[0][613] ) );
  AND U9952 ( .A(round_reg[614]), .B(init), .Z(\round_in[0][614] ) );
  AND U9953 ( .A(round_reg[615]), .B(init), .Z(\round_in[0][615] ) );
  AND U9954 ( .A(round_reg[616]), .B(init), .Z(\round_in[0][616] ) );
  AND U9955 ( .A(round_reg[617]), .B(init), .Z(\round_in[0][617] ) );
  AND U9956 ( .A(round_reg[618]), .B(init), .Z(\round_in[0][618] ) );
  AND U9957 ( .A(round_reg[619]), .B(init), .Z(\round_in[0][619] ) );
  NAND U9958 ( .A(init), .B(round_reg[61]), .Z(n3924) );
  NAND U9959 ( .A(n2846), .B(in[61]), .Z(n3923) );
  NAND U9960 ( .A(n3924), .B(n3923), .Z(\round_in[0][61] ) );
  AND U9961 ( .A(round_reg[620]), .B(init), .Z(\round_in[0][620] ) );
  AND U9962 ( .A(round_reg[621]), .B(init), .Z(\round_in[0][621] ) );
  AND U9963 ( .A(round_reg[622]), .B(init), .Z(\round_in[0][622] ) );
  AND U9964 ( .A(round_reg[623]), .B(init), .Z(\round_in[0][623] ) );
  AND U9965 ( .A(round_reg[624]), .B(init), .Z(\round_in[0][624] ) );
  AND U9966 ( .A(round_reg[625]), .B(init), .Z(\round_in[0][625] ) );
  AND U9967 ( .A(round_reg[626]), .B(init), .Z(\round_in[0][626] ) );
  AND U9968 ( .A(round_reg[627]), .B(init), .Z(\round_in[0][627] ) );
  AND U9969 ( .A(round_reg[628]), .B(init), .Z(\round_in[0][628] ) );
  AND U9970 ( .A(round_reg[629]), .B(init), .Z(\round_in[0][629] ) );
  NAND U9971 ( .A(init), .B(round_reg[62]), .Z(n3926) );
  NAND U9972 ( .A(n2846), .B(in[62]), .Z(n3925) );
  NAND U9973 ( .A(n3926), .B(n3925), .Z(\round_in[0][62] ) );
  AND U9974 ( .A(round_reg[630]), .B(init), .Z(\round_in[0][630] ) );
  AND U9975 ( .A(round_reg[631]), .B(init), .Z(\round_in[0][631] ) );
  AND U9976 ( .A(round_reg[632]), .B(init), .Z(\round_in[0][632] ) );
  AND U9977 ( .A(round_reg[633]), .B(init), .Z(\round_in[0][633] ) );
  AND U9978 ( .A(round_reg[634]), .B(init), .Z(\round_in[0][634] ) );
  AND U9979 ( .A(round_reg[635]), .B(init), .Z(\round_in[0][635] ) );
  AND U9980 ( .A(round_reg[636]), .B(init), .Z(\round_in[0][636] ) );
  AND U9981 ( .A(round_reg[637]), .B(init), .Z(\round_in[0][637] ) );
  AND U9982 ( .A(round_reg[638]), .B(init), .Z(\round_in[0][638] ) );
  AND U9983 ( .A(round_reg[639]), .B(init), .Z(\round_in[0][639] ) );
  NAND U9984 ( .A(init), .B(round_reg[63]), .Z(n3928) );
  NAND U9985 ( .A(n2846), .B(in[63]), .Z(n3927) );
  NAND U9986 ( .A(n3928), .B(n3927), .Z(\round_in[0][63] ) );
  AND U9987 ( .A(round_reg[640]), .B(init), .Z(\round_in[0][640] ) );
  AND U9988 ( .A(round_reg[641]), .B(init), .Z(\round_in[0][641] ) );
  AND U9989 ( .A(round_reg[642]), .B(init), .Z(\round_in[0][642] ) );
  AND U9990 ( .A(round_reg[643]), .B(init), .Z(\round_in[0][643] ) );
  AND U9991 ( .A(round_reg[644]), .B(init), .Z(\round_in[0][644] ) );
  AND U9992 ( .A(round_reg[645]), .B(init), .Z(\round_in[0][645] ) );
  AND U9993 ( .A(round_reg[646]), .B(init), .Z(\round_in[0][646] ) );
  AND U9994 ( .A(round_reg[647]), .B(init), .Z(\round_in[0][647] ) );
  AND U9995 ( .A(round_reg[648]), .B(init), .Z(\round_in[0][648] ) );
  AND U9996 ( .A(round_reg[649]), .B(init), .Z(\round_in[0][649] ) );
  NAND U9997 ( .A(init), .B(round_reg[64]), .Z(n3930) );
  NAND U9998 ( .A(n2846), .B(in[64]), .Z(n3929) );
  NAND U9999 ( .A(n3930), .B(n3929), .Z(\round_in[0][64] ) );
  AND U10000 ( .A(round_reg[650]), .B(init), .Z(\round_in[0][650] ) );
  AND U10001 ( .A(round_reg[651]), .B(init), .Z(\round_in[0][651] ) );
  AND U10002 ( .A(round_reg[652]), .B(init), .Z(\round_in[0][652] ) );
  AND U10003 ( .A(round_reg[653]), .B(init), .Z(\round_in[0][653] ) );
  AND U10004 ( .A(round_reg[654]), .B(init), .Z(\round_in[0][654] ) );
  AND U10005 ( .A(round_reg[655]), .B(init), .Z(\round_in[0][655] ) );
  AND U10006 ( .A(round_reg[656]), .B(init), .Z(\round_in[0][656] ) );
  AND U10007 ( .A(round_reg[657]), .B(init), .Z(\round_in[0][657] ) );
  AND U10008 ( .A(round_reg[658]), .B(init), .Z(\round_in[0][658] ) );
  AND U10009 ( .A(round_reg[659]), .B(init), .Z(\round_in[0][659] ) );
  NAND U10010 ( .A(init), .B(round_reg[65]), .Z(n3932) );
  NAND U10011 ( .A(n2847), .B(in[65]), .Z(n3931) );
  NAND U10012 ( .A(n3932), .B(n3931), .Z(\round_in[0][65] ) );
  AND U10013 ( .A(round_reg[660]), .B(init), .Z(\round_in[0][660] ) );
  AND U10014 ( .A(round_reg[661]), .B(init), .Z(\round_in[0][661] ) );
  AND U10015 ( .A(round_reg[662]), .B(init), .Z(\round_in[0][662] ) );
  AND U10016 ( .A(round_reg[663]), .B(init), .Z(\round_in[0][663] ) );
  AND U10017 ( .A(round_reg[664]), .B(init), .Z(\round_in[0][664] ) );
  AND U10018 ( .A(round_reg[665]), .B(init), .Z(\round_in[0][665] ) );
  AND U10019 ( .A(round_reg[666]), .B(init), .Z(\round_in[0][666] ) );
  AND U10020 ( .A(round_reg[667]), .B(init), .Z(\round_in[0][667] ) );
  AND U10021 ( .A(round_reg[668]), .B(init), .Z(\round_in[0][668] ) );
  AND U10022 ( .A(round_reg[669]), .B(init), .Z(\round_in[0][669] ) );
  NAND U10023 ( .A(init), .B(round_reg[66]), .Z(n3934) );
  NAND U10024 ( .A(n2847), .B(in[66]), .Z(n3933) );
  NAND U10025 ( .A(n3934), .B(n3933), .Z(\round_in[0][66] ) );
  AND U10026 ( .A(round_reg[670]), .B(init), .Z(\round_in[0][670] ) );
  AND U10027 ( .A(round_reg[671]), .B(init), .Z(\round_in[0][671] ) );
  AND U10028 ( .A(round_reg[672]), .B(init), .Z(\round_in[0][672] ) );
  AND U10029 ( .A(round_reg[673]), .B(init), .Z(\round_in[0][673] ) );
  AND U10030 ( .A(round_reg[674]), .B(init), .Z(\round_in[0][674] ) );
  AND U10031 ( .A(round_reg[675]), .B(init), .Z(\round_in[0][675] ) );
  AND U10032 ( .A(round_reg[676]), .B(init), .Z(\round_in[0][676] ) );
  AND U10033 ( .A(round_reg[677]), .B(init), .Z(\round_in[0][677] ) );
  AND U10034 ( .A(round_reg[678]), .B(init), .Z(\round_in[0][678] ) );
  AND U10035 ( .A(round_reg[679]), .B(init), .Z(\round_in[0][679] ) );
  NAND U10036 ( .A(init), .B(round_reg[67]), .Z(n3936) );
  NAND U10037 ( .A(n2847), .B(in[67]), .Z(n3935) );
  NAND U10038 ( .A(n3936), .B(n3935), .Z(\round_in[0][67] ) );
  AND U10039 ( .A(round_reg[680]), .B(init), .Z(\round_in[0][680] ) );
  AND U10040 ( .A(round_reg[681]), .B(init), .Z(\round_in[0][681] ) );
  AND U10041 ( .A(round_reg[682]), .B(init), .Z(\round_in[0][682] ) );
  AND U10042 ( .A(round_reg[683]), .B(init), .Z(\round_in[0][683] ) );
  AND U10043 ( .A(round_reg[684]), .B(init), .Z(\round_in[0][684] ) );
  AND U10044 ( .A(round_reg[685]), .B(init), .Z(\round_in[0][685] ) );
  AND U10045 ( .A(round_reg[686]), .B(init), .Z(\round_in[0][686] ) );
  AND U10046 ( .A(round_reg[687]), .B(init), .Z(\round_in[0][687] ) );
  AND U10047 ( .A(round_reg[688]), .B(init), .Z(\round_in[0][688] ) );
  AND U10048 ( .A(round_reg[689]), .B(init), .Z(\round_in[0][689] ) );
  NAND U10049 ( .A(init), .B(round_reg[68]), .Z(n3938) );
  NAND U10050 ( .A(n2847), .B(in[68]), .Z(n3937) );
  NAND U10051 ( .A(n3938), .B(n3937), .Z(\round_in[0][68] ) );
  AND U10052 ( .A(round_reg[690]), .B(init), .Z(\round_in[0][690] ) );
  AND U10053 ( .A(round_reg[691]), .B(init), .Z(\round_in[0][691] ) );
  AND U10054 ( .A(round_reg[692]), .B(init), .Z(\round_in[0][692] ) );
  AND U10055 ( .A(round_reg[693]), .B(init), .Z(\round_in[0][693] ) );
  AND U10056 ( .A(round_reg[694]), .B(init), .Z(\round_in[0][694] ) );
  AND U10057 ( .A(round_reg[695]), .B(init), .Z(\round_in[0][695] ) );
  AND U10058 ( .A(round_reg[696]), .B(init), .Z(\round_in[0][696] ) );
  AND U10059 ( .A(round_reg[697]), .B(init), .Z(\round_in[0][697] ) );
  AND U10060 ( .A(round_reg[698]), .B(init), .Z(\round_in[0][698] ) );
  AND U10061 ( .A(round_reg[699]), .B(init), .Z(\round_in[0][699] ) );
  NAND U10062 ( .A(init), .B(round_reg[69]), .Z(n3940) );
  NAND U10063 ( .A(n2847), .B(in[69]), .Z(n3939) );
  NAND U10064 ( .A(n3940), .B(n3939), .Z(\round_in[0][69] ) );
  NAND U10065 ( .A(init), .B(round_reg[6]), .Z(n3942) );
  NAND U10066 ( .A(n2847), .B(in[6]), .Z(n3941) );
  NAND U10067 ( .A(n3942), .B(n3941), .Z(\round_in[0][6] ) );
  AND U10068 ( .A(round_reg[700]), .B(init), .Z(\round_in[0][700] ) );
  AND U10069 ( .A(round_reg[701]), .B(init), .Z(\round_in[0][701] ) );
  AND U10070 ( .A(round_reg[702]), .B(init), .Z(\round_in[0][702] ) );
  AND U10071 ( .A(round_reg[703]), .B(init), .Z(\round_in[0][703] ) );
  AND U10072 ( .A(round_reg[704]), .B(init), .Z(\round_in[0][704] ) );
  AND U10073 ( .A(round_reg[705]), .B(init), .Z(\round_in[0][705] ) );
  AND U10074 ( .A(round_reg[706]), .B(init), .Z(\round_in[0][706] ) );
  AND U10075 ( .A(round_reg[707]), .B(init), .Z(\round_in[0][707] ) );
  AND U10076 ( .A(round_reg[708]), .B(init), .Z(\round_in[0][708] ) );
  AND U10077 ( .A(round_reg[709]), .B(init), .Z(\round_in[0][709] ) );
  NAND U10078 ( .A(init), .B(round_reg[70]), .Z(n3944) );
  NAND U10079 ( .A(n2847), .B(in[70]), .Z(n3943) );
  NAND U10080 ( .A(n3944), .B(n3943), .Z(\round_in[0][70] ) );
  AND U10081 ( .A(round_reg[710]), .B(init), .Z(\round_in[0][710] ) );
  AND U10082 ( .A(round_reg[711]), .B(init), .Z(\round_in[0][711] ) );
  AND U10083 ( .A(round_reg[712]), .B(init), .Z(\round_in[0][712] ) );
  AND U10084 ( .A(round_reg[713]), .B(init), .Z(\round_in[0][713] ) );
  AND U10085 ( .A(round_reg[714]), .B(init), .Z(\round_in[0][714] ) );
  AND U10086 ( .A(round_reg[715]), .B(init), .Z(\round_in[0][715] ) );
  AND U10087 ( .A(round_reg[716]), .B(init), .Z(\round_in[0][716] ) );
  AND U10088 ( .A(round_reg[717]), .B(init), .Z(\round_in[0][717] ) );
  AND U10089 ( .A(round_reg[718]), .B(init), .Z(\round_in[0][718] ) );
  AND U10090 ( .A(round_reg[719]), .B(init), .Z(\round_in[0][719] ) );
  NAND U10091 ( .A(init), .B(round_reg[71]), .Z(n3946) );
  NAND U10092 ( .A(n2848), .B(in[71]), .Z(n3945) );
  NAND U10093 ( .A(n3946), .B(n3945), .Z(\round_in[0][71] ) );
  AND U10094 ( .A(round_reg[720]), .B(init), .Z(\round_in[0][720] ) );
  AND U10095 ( .A(round_reg[721]), .B(init), .Z(\round_in[0][721] ) );
  AND U10096 ( .A(round_reg[722]), .B(init), .Z(\round_in[0][722] ) );
  AND U10097 ( .A(round_reg[723]), .B(init), .Z(\round_in[0][723] ) );
  AND U10098 ( .A(round_reg[724]), .B(init), .Z(\round_in[0][724] ) );
  AND U10099 ( .A(round_reg[725]), .B(init), .Z(\round_in[0][725] ) );
  AND U10100 ( .A(round_reg[726]), .B(init), .Z(\round_in[0][726] ) );
  AND U10101 ( .A(round_reg[727]), .B(init), .Z(\round_in[0][727] ) );
  AND U10102 ( .A(round_reg[728]), .B(init), .Z(\round_in[0][728] ) );
  AND U10103 ( .A(round_reg[729]), .B(init), .Z(\round_in[0][729] ) );
  NAND U10104 ( .A(init), .B(round_reg[72]), .Z(n3948) );
  NAND U10105 ( .A(n2848), .B(in[72]), .Z(n3947) );
  NAND U10106 ( .A(n3948), .B(n3947), .Z(\round_in[0][72] ) );
  AND U10107 ( .A(round_reg[730]), .B(init), .Z(\round_in[0][730] ) );
  AND U10108 ( .A(round_reg[731]), .B(init), .Z(\round_in[0][731] ) );
  AND U10109 ( .A(round_reg[732]), .B(init), .Z(\round_in[0][732] ) );
  AND U10110 ( .A(round_reg[733]), .B(init), .Z(\round_in[0][733] ) );
  AND U10111 ( .A(round_reg[734]), .B(init), .Z(\round_in[0][734] ) );
  AND U10112 ( .A(round_reg[735]), .B(init), .Z(\round_in[0][735] ) );
  AND U10113 ( .A(round_reg[736]), .B(init), .Z(\round_in[0][736] ) );
  AND U10114 ( .A(round_reg[737]), .B(init), .Z(\round_in[0][737] ) );
  AND U10115 ( .A(round_reg[738]), .B(init), .Z(\round_in[0][738] ) );
  AND U10116 ( .A(round_reg[739]), .B(init), .Z(\round_in[0][739] ) );
  NAND U10117 ( .A(init), .B(round_reg[73]), .Z(n3950) );
  NAND U10118 ( .A(n2848), .B(in[73]), .Z(n3949) );
  NAND U10119 ( .A(n3950), .B(n3949), .Z(\round_in[0][73] ) );
  AND U10120 ( .A(round_reg[740]), .B(init), .Z(\round_in[0][740] ) );
  AND U10121 ( .A(round_reg[741]), .B(init), .Z(\round_in[0][741] ) );
  AND U10122 ( .A(round_reg[742]), .B(init), .Z(\round_in[0][742] ) );
  AND U10123 ( .A(round_reg[743]), .B(init), .Z(\round_in[0][743] ) );
  AND U10124 ( .A(round_reg[744]), .B(init), .Z(\round_in[0][744] ) );
  AND U10125 ( .A(round_reg[745]), .B(init), .Z(\round_in[0][745] ) );
  AND U10126 ( .A(round_reg[746]), .B(init), .Z(\round_in[0][746] ) );
  AND U10127 ( .A(round_reg[747]), .B(init), .Z(\round_in[0][747] ) );
  AND U10128 ( .A(round_reg[748]), .B(init), .Z(\round_in[0][748] ) );
  AND U10129 ( .A(round_reg[749]), .B(init), .Z(\round_in[0][749] ) );
  NAND U10130 ( .A(init), .B(round_reg[74]), .Z(n3952) );
  NAND U10131 ( .A(n2848), .B(in[74]), .Z(n3951) );
  NAND U10132 ( .A(n3952), .B(n3951), .Z(\round_in[0][74] ) );
  AND U10133 ( .A(round_reg[750]), .B(init), .Z(\round_in[0][750] ) );
  AND U10134 ( .A(round_reg[751]), .B(init), .Z(\round_in[0][751] ) );
  AND U10135 ( .A(round_reg[752]), .B(init), .Z(\round_in[0][752] ) );
  AND U10136 ( .A(round_reg[753]), .B(init), .Z(\round_in[0][753] ) );
  AND U10137 ( .A(round_reg[754]), .B(init), .Z(\round_in[0][754] ) );
  AND U10138 ( .A(round_reg[755]), .B(init), .Z(\round_in[0][755] ) );
  AND U10139 ( .A(round_reg[756]), .B(init), .Z(\round_in[0][756] ) );
  AND U10140 ( .A(round_reg[757]), .B(init), .Z(\round_in[0][757] ) );
  AND U10141 ( .A(round_reg[758]), .B(init), .Z(\round_in[0][758] ) );
  AND U10142 ( .A(round_reg[759]), .B(init), .Z(\round_in[0][759] ) );
  NAND U10143 ( .A(init), .B(round_reg[75]), .Z(n3954) );
  NAND U10144 ( .A(n2848), .B(in[75]), .Z(n3953) );
  NAND U10145 ( .A(n3954), .B(n3953), .Z(\round_in[0][75] ) );
  AND U10146 ( .A(round_reg[760]), .B(init), .Z(\round_in[0][760] ) );
  AND U10147 ( .A(round_reg[761]), .B(init), .Z(\round_in[0][761] ) );
  AND U10148 ( .A(round_reg[762]), .B(init), .Z(\round_in[0][762] ) );
  AND U10149 ( .A(round_reg[763]), .B(init), .Z(\round_in[0][763] ) );
  AND U10150 ( .A(round_reg[764]), .B(init), .Z(\round_in[0][764] ) );
  AND U10151 ( .A(round_reg[765]), .B(init), .Z(\round_in[0][765] ) );
  AND U10152 ( .A(round_reg[766]), .B(init), .Z(\round_in[0][766] ) );
  AND U10153 ( .A(round_reg[767]), .B(init), .Z(\round_in[0][767] ) );
  AND U10154 ( .A(round_reg[768]), .B(init), .Z(\round_in[0][768] ) );
  AND U10155 ( .A(round_reg[769]), .B(init), .Z(\round_in[0][769] ) );
  NAND U10156 ( .A(init), .B(round_reg[76]), .Z(n3956) );
  NAND U10157 ( .A(n2848), .B(in[76]), .Z(n3955) );
  NAND U10158 ( .A(n3956), .B(n3955), .Z(\round_in[0][76] ) );
  AND U10159 ( .A(round_reg[770]), .B(init), .Z(\round_in[0][770] ) );
  AND U10160 ( .A(round_reg[771]), .B(init), .Z(\round_in[0][771] ) );
  AND U10161 ( .A(round_reg[772]), .B(init), .Z(\round_in[0][772] ) );
  AND U10162 ( .A(round_reg[773]), .B(init), .Z(\round_in[0][773] ) );
  AND U10163 ( .A(round_reg[774]), .B(init), .Z(\round_in[0][774] ) );
  AND U10164 ( .A(round_reg[775]), .B(init), .Z(\round_in[0][775] ) );
  AND U10165 ( .A(round_reg[776]), .B(init), .Z(\round_in[0][776] ) );
  AND U10166 ( .A(round_reg[777]), .B(init), .Z(\round_in[0][777] ) );
  AND U10167 ( .A(round_reg[778]), .B(init), .Z(\round_in[0][778] ) );
  AND U10168 ( .A(round_reg[779]), .B(init), .Z(\round_in[0][779] ) );
  NAND U10169 ( .A(init), .B(round_reg[77]), .Z(n3958) );
  NAND U10170 ( .A(n2848), .B(in[77]), .Z(n3957) );
  NAND U10171 ( .A(n3958), .B(n3957), .Z(\round_in[0][77] ) );
  AND U10172 ( .A(round_reg[780]), .B(init), .Z(\round_in[0][780] ) );
  AND U10173 ( .A(round_reg[781]), .B(init), .Z(\round_in[0][781] ) );
  AND U10174 ( .A(round_reg[782]), .B(init), .Z(\round_in[0][782] ) );
  AND U10175 ( .A(round_reg[783]), .B(init), .Z(\round_in[0][783] ) );
  AND U10176 ( .A(round_reg[784]), .B(init), .Z(\round_in[0][784] ) );
  AND U10177 ( .A(round_reg[785]), .B(init), .Z(\round_in[0][785] ) );
  AND U10178 ( .A(round_reg[786]), .B(init), .Z(\round_in[0][786] ) );
  AND U10179 ( .A(round_reg[787]), .B(init), .Z(\round_in[0][787] ) );
  AND U10180 ( .A(round_reg[788]), .B(init), .Z(\round_in[0][788] ) );
  AND U10181 ( .A(round_reg[789]), .B(init), .Z(\round_in[0][789] ) );
  NAND U10182 ( .A(init), .B(round_reg[78]), .Z(n3960) );
  NAND U10183 ( .A(n2849), .B(in[78]), .Z(n3959) );
  NAND U10184 ( .A(n3960), .B(n3959), .Z(\round_in[0][78] ) );
  AND U10185 ( .A(round_reg[790]), .B(init), .Z(\round_in[0][790] ) );
  AND U10186 ( .A(round_reg[791]), .B(init), .Z(\round_in[0][791] ) );
  AND U10187 ( .A(round_reg[792]), .B(init), .Z(\round_in[0][792] ) );
  AND U10188 ( .A(round_reg[793]), .B(init), .Z(\round_in[0][793] ) );
  AND U10189 ( .A(round_reg[794]), .B(init), .Z(\round_in[0][794] ) );
  AND U10190 ( .A(round_reg[795]), .B(init), .Z(\round_in[0][795] ) );
  AND U10191 ( .A(round_reg[796]), .B(init), .Z(\round_in[0][796] ) );
  AND U10192 ( .A(round_reg[797]), .B(init), .Z(\round_in[0][797] ) );
  AND U10193 ( .A(round_reg[798]), .B(init), .Z(\round_in[0][798] ) );
  AND U10194 ( .A(round_reg[799]), .B(init), .Z(\round_in[0][799] ) );
  NAND U10195 ( .A(init), .B(round_reg[79]), .Z(n3962) );
  NAND U10196 ( .A(n2849), .B(in[79]), .Z(n3961) );
  NAND U10197 ( .A(n3962), .B(n3961), .Z(\round_in[0][79] ) );
  NAND U10198 ( .A(init), .B(round_reg[7]), .Z(n3964) );
  NAND U10199 ( .A(n2849), .B(in[7]), .Z(n3963) );
  NAND U10200 ( .A(n3964), .B(n3963), .Z(\round_in[0][7] ) );
  AND U10201 ( .A(round_reg[800]), .B(init), .Z(\round_in[0][800] ) );
  AND U10202 ( .A(round_reg[801]), .B(init), .Z(\round_in[0][801] ) );
  AND U10203 ( .A(round_reg[802]), .B(init), .Z(\round_in[0][802] ) );
  AND U10204 ( .A(round_reg[803]), .B(init), .Z(\round_in[0][803] ) );
  AND U10205 ( .A(round_reg[804]), .B(init), .Z(\round_in[0][804] ) );
  AND U10206 ( .A(round_reg[805]), .B(init), .Z(\round_in[0][805] ) );
  AND U10207 ( .A(round_reg[806]), .B(init), .Z(\round_in[0][806] ) );
  AND U10208 ( .A(round_reg[807]), .B(init), .Z(\round_in[0][807] ) );
  AND U10209 ( .A(round_reg[808]), .B(init), .Z(\round_in[0][808] ) );
  AND U10210 ( .A(round_reg[809]), .B(init), .Z(\round_in[0][809] ) );
  NAND U10211 ( .A(init), .B(round_reg[80]), .Z(n3966) );
  NAND U10212 ( .A(n2849), .B(in[80]), .Z(n3965) );
  NAND U10213 ( .A(n3966), .B(n3965), .Z(\round_in[0][80] ) );
  AND U10214 ( .A(round_reg[810]), .B(init), .Z(\round_in[0][810] ) );
  AND U10215 ( .A(round_reg[811]), .B(init), .Z(\round_in[0][811] ) );
  AND U10216 ( .A(round_reg[812]), .B(init), .Z(\round_in[0][812] ) );
  AND U10217 ( .A(round_reg[813]), .B(init), .Z(\round_in[0][813] ) );
  AND U10218 ( .A(round_reg[814]), .B(init), .Z(\round_in[0][814] ) );
  AND U10219 ( .A(round_reg[815]), .B(init), .Z(\round_in[0][815] ) );
  AND U10220 ( .A(round_reg[816]), .B(init), .Z(\round_in[0][816] ) );
  AND U10221 ( .A(round_reg[817]), .B(init), .Z(\round_in[0][817] ) );
  AND U10222 ( .A(round_reg[818]), .B(init), .Z(\round_in[0][818] ) );
  AND U10223 ( .A(round_reg[819]), .B(init), .Z(\round_in[0][819] ) );
  NAND U10224 ( .A(init), .B(round_reg[81]), .Z(n3968) );
  NAND U10225 ( .A(n2849), .B(in[81]), .Z(n3967) );
  NAND U10226 ( .A(n3968), .B(n3967), .Z(\round_in[0][81] ) );
  AND U10227 ( .A(round_reg[820]), .B(init), .Z(\round_in[0][820] ) );
  AND U10228 ( .A(round_reg[821]), .B(init), .Z(\round_in[0][821] ) );
  AND U10229 ( .A(round_reg[822]), .B(init), .Z(\round_in[0][822] ) );
  AND U10230 ( .A(round_reg[823]), .B(init), .Z(\round_in[0][823] ) );
  AND U10231 ( .A(round_reg[824]), .B(init), .Z(\round_in[0][824] ) );
  AND U10232 ( .A(round_reg[825]), .B(init), .Z(\round_in[0][825] ) );
  AND U10233 ( .A(round_reg[826]), .B(init), .Z(\round_in[0][826] ) );
  AND U10234 ( .A(round_reg[827]), .B(init), .Z(\round_in[0][827] ) );
  AND U10235 ( .A(round_reg[828]), .B(init), .Z(\round_in[0][828] ) );
  AND U10236 ( .A(round_reg[829]), .B(init), .Z(\round_in[0][829] ) );
  NAND U10237 ( .A(init), .B(round_reg[82]), .Z(n3970) );
  NAND U10238 ( .A(n2849), .B(in[82]), .Z(n3969) );
  NAND U10239 ( .A(n3970), .B(n3969), .Z(\round_in[0][82] ) );
  AND U10240 ( .A(round_reg[830]), .B(init), .Z(\round_in[0][830] ) );
  AND U10241 ( .A(round_reg[831]), .B(init), .Z(\round_in[0][831] ) );
  AND U10242 ( .A(round_reg[832]), .B(init), .Z(\round_in[0][832] ) );
  AND U10243 ( .A(round_reg[833]), .B(init), .Z(\round_in[0][833] ) );
  AND U10244 ( .A(round_reg[834]), .B(init), .Z(\round_in[0][834] ) );
  AND U10245 ( .A(round_reg[835]), .B(init), .Z(\round_in[0][835] ) );
  AND U10246 ( .A(round_reg[836]), .B(init), .Z(\round_in[0][836] ) );
  AND U10247 ( .A(round_reg[837]), .B(init), .Z(\round_in[0][837] ) );
  AND U10248 ( .A(round_reg[838]), .B(init), .Z(\round_in[0][838] ) );
  AND U10249 ( .A(round_reg[839]), .B(init), .Z(\round_in[0][839] ) );
  NAND U10250 ( .A(init), .B(round_reg[83]), .Z(n3972) );
  NAND U10251 ( .A(n2849), .B(in[83]), .Z(n3971) );
  NAND U10252 ( .A(n3972), .B(n3971), .Z(\round_in[0][83] ) );
  AND U10253 ( .A(round_reg[840]), .B(init), .Z(\round_in[0][840] ) );
  AND U10254 ( .A(round_reg[841]), .B(init), .Z(\round_in[0][841] ) );
  AND U10255 ( .A(round_reg[842]), .B(init), .Z(\round_in[0][842] ) );
  AND U10256 ( .A(round_reg[843]), .B(init), .Z(\round_in[0][843] ) );
  AND U10257 ( .A(round_reg[844]), .B(init), .Z(\round_in[0][844] ) );
  AND U10258 ( .A(round_reg[845]), .B(init), .Z(\round_in[0][845] ) );
  AND U10259 ( .A(round_reg[846]), .B(init), .Z(\round_in[0][846] ) );
  AND U10260 ( .A(round_reg[847]), .B(init), .Z(\round_in[0][847] ) );
  AND U10261 ( .A(round_reg[848]), .B(init), .Z(\round_in[0][848] ) );
  AND U10262 ( .A(round_reg[849]), .B(init), .Z(\round_in[0][849] ) );
  NAND U10263 ( .A(init), .B(round_reg[84]), .Z(n3974) );
  NAND U10264 ( .A(n2850), .B(in[84]), .Z(n3973) );
  NAND U10265 ( .A(n3974), .B(n3973), .Z(\round_in[0][84] ) );
  AND U10266 ( .A(round_reg[850]), .B(init), .Z(\round_in[0][850] ) );
  AND U10267 ( .A(round_reg[851]), .B(init), .Z(\round_in[0][851] ) );
  AND U10268 ( .A(round_reg[852]), .B(init), .Z(\round_in[0][852] ) );
  AND U10269 ( .A(round_reg[853]), .B(init), .Z(\round_in[0][853] ) );
  AND U10270 ( .A(round_reg[854]), .B(init), .Z(\round_in[0][854] ) );
  AND U10271 ( .A(round_reg[855]), .B(init), .Z(\round_in[0][855] ) );
  AND U10272 ( .A(round_reg[856]), .B(init), .Z(\round_in[0][856] ) );
  AND U10273 ( .A(round_reg[857]), .B(init), .Z(\round_in[0][857] ) );
  AND U10274 ( .A(round_reg[858]), .B(init), .Z(\round_in[0][858] ) );
  AND U10275 ( .A(round_reg[859]), .B(init), .Z(\round_in[0][859] ) );
  NAND U10276 ( .A(init), .B(round_reg[85]), .Z(n3976) );
  NAND U10277 ( .A(n2850), .B(in[85]), .Z(n3975) );
  NAND U10278 ( .A(n3976), .B(n3975), .Z(\round_in[0][85] ) );
  AND U10279 ( .A(round_reg[860]), .B(init), .Z(\round_in[0][860] ) );
  AND U10280 ( .A(round_reg[861]), .B(init), .Z(\round_in[0][861] ) );
  AND U10281 ( .A(round_reg[862]), .B(init), .Z(\round_in[0][862] ) );
  AND U10282 ( .A(round_reg[863]), .B(init), .Z(\round_in[0][863] ) );
  AND U10283 ( .A(round_reg[864]), .B(init), .Z(\round_in[0][864] ) );
  AND U10284 ( .A(round_reg[865]), .B(init), .Z(\round_in[0][865] ) );
  AND U10285 ( .A(round_reg[866]), .B(init), .Z(\round_in[0][866] ) );
  AND U10286 ( .A(round_reg[867]), .B(init), .Z(\round_in[0][867] ) );
  AND U10287 ( .A(round_reg[868]), .B(init), .Z(\round_in[0][868] ) );
  AND U10288 ( .A(round_reg[869]), .B(init), .Z(\round_in[0][869] ) );
  NAND U10289 ( .A(init), .B(round_reg[86]), .Z(n3978) );
  NAND U10290 ( .A(n2850), .B(in[86]), .Z(n3977) );
  NAND U10291 ( .A(n3978), .B(n3977), .Z(\round_in[0][86] ) );
  AND U10292 ( .A(round_reg[870]), .B(init), .Z(\round_in[0][870] ) );
  AND U10293 ( .A(round_reg[871]), .B(init), .Z(\round_in[0][871] ) );
  AND U10294 ( .A(round_reg[872]), .B(init), .Z(\round_in[0][872] ) );
  AND U10295 ( .A(round_reg[873]), .B(init), .Z(\round_in[0][873] ) );
  AND U10296 ( .A(round_reg[874]), .B(init), .Z(\round_in[0][874] ) );
  AND U10297 ( .A(round_reg[875]), .B(init), .Z(\round_in[0][875] ) );
  AND U10298 ( .A(round_reg[876]), .B(init), .Z(\round_in[0][876] ) );
  AND U10299 ( .A(round_reg[877]), .B(init), .Z(\round_in[0][877] ) );
  AND U10300 ( .A(round_reg[878]), .B(init), .Z(\round_in[0][878] ) );
  AND U10301 ( .A(round_reg[879]), .B(init), .Z(\round_in[0][879] ) );
  NAND U10302 ( .A(init), .B(round_reg[87]), .Z(n3980) );
  NAND U10303 ( .A(n2850), .B(in[87]), .Z(n3979) );
  NAND U10304 ( .A(n3980), .B(n3979), .Z(\round_in[0][87] ) );
  AND U10305 ( .A(round_reg[880]), .B(init), .Z(\round_in[0][880] ) );
  AND U10306 ( .A(round_reg[881]), .B(init), .Z(\round_in[0][881] ) );
  AND U10307 ( .A(round_reg[882]), .B(init), .Z(\round_in[0][882] ) );
  AND U10308 ( .A(round_reg[883]), .B(init), .Z(\round_in[0][883] ) );
  AND U10309 ( .A(round_reg[884]), .B(init), .Z(\round_in[0][884] ) );
  AND U10310 ( .A(round_reg[885]), .B(init), .Z(\round_in[0][885] ) );
  AND U10311 ( .A(round_reg[886]), .B(init), .Z(\round_in[0][886] ) );
  AND U10312 ( .A(round_reg[887]), .B(init), .Z(\round_in[0][887] ) );
  AND U10313 ( .A(round_reg[888]), .B(init), .Z(\round_in[0][888] ) );
  AND U10314 ( .A(round_reg[889]), .B(init), .Z(\round_in[0][889] ) );
  NAND U10315 ( .A(init), .B(round_reg[88]), .Z(n3982) );
  NAND U10316 ( .A(n2850), .B(in[88]), .Z(n3981) );
  NAND U10317 ( .A(n3982), .B(n3981), .Z(\round_in[0][88] ) );
  AND U10318 ( .A(round_reg[890]), .B(init), .Z(\round_in[0][890] ) );
  AND U10319 ( .A(round_reg[891]), .B(init), .Z(\round_in[0][891] ) );
  AND U10320 ( .A(round_reg[892]), .B(init), .Z(\round_in[0][892] ) );
  AND U10321 ( .A(round_reg[893]), .B(init), .Z(\round_in[0][893] ) );
  AND U10322 ( .A(round_reg[894]), .B(init), .Z(\round_in[0][894] ) );
  AND U10323 ( .A(round_reg[895]), .B(init), .Z(\round_in[0][895] ) );
  AND U10324 ( .A(round_reg[896]), .B(init), .Z(\round_in[0][896] ) );
  AND U10325 ( .A(round_reg[897]), .B(init), .Z(\round_in[0][897] ) );
  AND U10326 ( .A(round_reg[898]), .B(init), .Z(\round_in[0][898] ) );
  AND U10327 ( .A(round_reg[899]), .B(init), .Z(\round_in[0][899] ) );
  NAND U10328 ( .A(init), .B(round_reg[89]), .Z(n3984) );
  NAND U10329 ( .A(n2850), .B(in[89]), .Z(n3983) );
  NAND U10330 ( .A(n3984), .B(n3983), .Z(\round_in[0][89] ) );
  NAND U10331 ( .A(init), .B(round_reg[8]), .Z(n3986) );
  NAND U10332 ( .A(n2850), .B(in[8]), .Z(n3985) );
  NAND U10333 ( .A(n3986), .B(n3985), .Z(\round_in[0][8] ) );
  AND U10334 ( .A(round_reg[900]), .B(init), .Z(\round_in[0][900] ) );
  AND U10335 ( .A(round_reg[901]), .B(init), .Z(\round_in[0][901] ) );
  AND U10336 ( .A(round_reg[902]), .B(init), .Z(\round_in[0][902] ) );
  AND U10337 ( .A(round_reg[903]), .B(init), .Z(\round_in[0][903] ) );
  AND U10338 ( .A(round_reg[904]), .B(init), .Z(\round_in[0][904] ) );
  AND U10339 ( .A(round_reg[905]), .B(init), .Z(\round_in[0][905] ) );
  AND U10340 ( .A(round_reg[906]), .B(init), .Z(\round_in[0][906] ) );
  AND U10341 ( .A(round_reg[907]), .B(init), .Z(\round_in[0][907] ) );
  AND U10342 ( .A(round_reg[908]), .B(init), .Z(\round_in[0][908] ) );
  AND U10343 ( .A(round_reg[909]), .B(init), .Z(\round_in[0][909] ) );
  NAND U10344 ( .A(init), .B(round_reg[90]), .Z(n3988) );
  NAND U10345 ( .A(n2851), .B(in[90]), .Z(n3987) );
  NAND U10346 ( .A(n3988), .B(n3987), .Z(\round_in[0][90] ) );
  AND U10347 ( .A(round_reg[910]), .B(init), .Z(\round_in[0][910] ) );
  AND U10348 ( .A(round_reg[911]), .B(init), .Z(\round_in[0][911] ) );
  AND U10349 ( .A(round_reg[912]), .B(init), .Z(\round_in[0][912] ) );
  AND U10350 ( .A(round_reg[913]), .B(init), .Z(\round_in[0][913] ) );
  AND U10351 ( .A(round_reg[914]), .B(init), .Z(\round_in[0][914] ) );
  AND U10352 ( .A(round_reg[915]), .B(init), .Z(\round_in[0][915] ) );
  AND U10353 ( .A(round_reg[916]), .B(init), .Z(\round_in[0][916] ) );
  AND U10354 ( .A(round_reg[917]), .B(init), .Z(\round_in[0][917] ) );
  AND U10355 ( .A(round_reg[918]), .B(init), .Z(\round_in[0][918] ) );
  AND U10356 ( .A(round_reg[919]), .B(init), .Z(\round_in[0][919] ) );
  NAND U10357 ( .A(init), .B(round_reg[91]), .Z(n3990) );
  NAND U10358 ( .A(n2851), .B(in[91]), .Z(n3989) );
  NAND U10359 ( .A(n3990), .B(n3989), .Z(\round_in[0][91] ) );
  AND U10360 ( .A(round_reg[920]), .B(init), .Z(\round_in[0][920] ) );
  AND U10361 ( .A(round_reg[921]), .B(init), .Z(\round_in[0][921] ) );
  AND U10362 ( .A(round_reg[922]), .B(init), .Z(\round_in[0][922] ) );
  AND U10363 ( .A(round_reg[923]), .B(init), .Z(\round_in[0][923] ) );
  AND U10364 ( .A(round_reg[924]), .B(init), .Z(\round_in[0][924] ) );
  AND U10365 ( .A(round_reg[925]), .B(init), .Z(\round_in[0][925] ) );
  AND U10366 ( .A(round_reg[926]), .B(init), .Z(\round_in[0][926] ) );
  AND U10367 ( .A(round_reg[927]), .B(init), .Z(\round_in[0][927] ) );
  AND U10368 ( .A(round_reg[928]), .B(init), .Z(\round_in[0][928] ) );
  AND U10369 ( .A(round_reg[929]), .B(init), .Z(\round_in[0][929] ) );
  NAND U10370 ( .A(init), .B(round_reg[92]), .Z(n3992) );
  NAND U10371 ( .A(n2851), .B(in[92]), .Z(n3991) );
  NAND U10372 ( .A(n3992), .B(n3991), .Z(\round_in[0][92] ) );
  AND U10373 ( .A(round_reg[930]), .B(init), .Z(\round_in[0][930] ) );
  AND U10374 ( .A(round_reg[931]), .B(init), .Z(\round_in[0][931] ) );
  AND U10375 ( .A(round_reg[932]), .B(init), .Z(\round_in[0][932] ) );
  AND U10376 ( .A(round_reg[933]), .B(init), .Z(\round_in[0][933] ) );
  AND U10377 ( .A(round_reg[934]), .B(init), .Z(\round_in[0][934] ) );
  AND U10378 ( .A(round_reg[935]), .B(init), .Z(\round_in[0][935] ) );
  AND U10379 ( .A(round_reg[936]), .B(init), .Z(\round_in[0][936] ) );
  AND U10380 ( .A(round_reg[937]), .B(init), .Z(\round_in[0][937] ) );
  AND U10381 ( .A(round_reg[938]), .B(init), .Z(\round_in[0][938] ) );
  AND U10382 ( .A(round_reg[939]), .B(init), .Z(\round_in[0][939] ) );
  NAND U10383 ( .A(init), .B(round_reg[93]), .Z(n3994) );
  NAND U10384 ( .A(n2851), .B(in[93]), .Z(n3993) );
  NAND U10385 ( .A(n3994), .B(n3993), .Z(\round_in[0][93] ) );
  AND U10386 ( .A(round_reg[940]), .B(init), .Z(\round_in[0][940] ) );
  AND U10387 ( .A(round_reg[941]), .B(init), .Z(\round_in[0][941] ) );
  AND U10388 ( .A(round_reg[942]), .B(init), .Z(\round_in[0][942] ) );
  AND U10389 ( .A(round_reg[943]), .B(init), .Z(\round_in[0][943] ) );
  AND U10390 ( .A(round_reg[944]), .B(init), .Z(\round_in[0][944] ) );
  AND U10391 ( .A(round_reg[945]), .B(init), .Z(\round_in[0][945] ) );
  AND U10392 ( .A(round_reg[946]), .B(init), .Z(\round_in[0][946] ) );
  AND U10393 ( .A(round_reg[947]), .B(init), .Z(\round_in[0][947] ) );
  AND U10394 ( .A(round_reg[948]), .B(init), .Z(\round_in[0][948] ) );
  AND U10395 ( .A(round_reg[949]), .B(init), .Z(\round_in[0][949] ) );
  NAND U10396 ( .A(init), .B(round_reg[94]), .Z(n3996) );
  NAND U10397 ( .A(n2851), .B(in[94]), .Z(n3995) );
  NAND U10398 ( .A(n3996), .B(n3995), .Z(\round_in[0][94] ) );
  AND U10399 ( .A(round_reg[950]), .B(init), .Z(\round_in[0][950] ) );
  AND U10400 ( .A(round_reg[951]), .B(init), .Z(\round_in[0][951] ) );
  AND U10401 ( .A(round_reg[952]), .B(init), .Z(\round_in[0][952] ) );
  AND U10402 ( .A(round_reg[953]), .B(init), .Z(\round_in[0][953] ) );
  AND U10403 ( .A(round_reg[954]), .B(init), .Z(\round_in[0][954] ) );
  AND U10404 ( .A(round_reg[955]), .B(init), .Z(\round_in[0][955] ) );
  AND U10405 ( .A(round_reg[956]), .B(init), .Z(\round_in[0][956] ) );
  AND U10406 ( .A(round_reg[957]), .B(init), .Z(\round_in[0][957] ) );
  AND U10407 ( .A(round_reg[958]), .B(init), .Z(\round_in[0][958] ) );
  AND U10408 ( .A(round_reg[959]), .B(init), .Z(\round_in[0][959] ) );
  NAND U10409 ( .A(init), .B(round_reg[95]), .Z(n3998) );
  NAND U10410 ( .A(n2851), .B(in[95]), .Z(n3997) );
  NAND U10411 ( .A(n3998), .B(n3997), .Z(\round_in[0][95] ) );
  AND U10412 ( .A(round_reg[960]), .B(init), .Z(\round_in[0][960] ) );
  AND U10413 ( .A(round_reg[961]), .B(init), .Z(\round_in[0][961] ) );
  AND U10414 ( .A(round_reg[962]), .B(init), .Z(\round_in[0][962] ) );
  AND U10415 ( .A(round_reg[963]), .B(init), .Z(\round_in[0][963] ) );
  AND U10416 ( .A(round_reg[964]), .B(init), .Z(\round_in[0][964] ) );
  AND U10417 ( .A(round_reg[965]), .B(init), .Z(\round_in[0][965] ) );
  AND U10418 ( .A(round_reg[966]), .B(init), .Z(\round_in[0][966] ) );
  AND U10419 ( .A(round_reg[967]), .B(init), .Z(\round_in[0][967] ) );
  AND U10420 ( .A(round_reg[968]), .B(init), .Z(\round_in[0][968] ) );
  AND U10421 ( .A(round_reg[969]), .B(init), .Z(\round_in[0][969] ) );
  NAND U10422 ( .A(init), .B(round_reg[96]), .Z(n4000) );
  NAND U10423 ( .A(n2851), .B(in[96]), .Z(n3999) );
  NAND U10424 ( .A(n4000), .B(n3999), .Z(\round_in[0][96] ) );
  AND U10425 ( .A(round_reg[970]), .B(init), .Z(\round_in[0][970] ) );
  AND U10426 ( .A(round_reg[971]), .B(init), .Z(\round_in[0][971] ) );
  AND U10427 ( .A(round_reg[972]), .B(init), .Z(\round_in[0][972] ) );
  AND U10428 ( .A(round_reg[973]), .B(init), .Z(\round_in[0][973] ) );
  AND U10429 ( .A(round_reg[974]), .B(init), .Z(\round_in[0][974] ) );
  AND U10430 ( .A(round_reg[975]), .B(init), .Z(\round_in[0][975] ) );
  AND U10431 ( .A(round_reg[976]), .B(init), .Z(\round_in[0][976] ) );
  AND U10432 ( .A(round_reg[977]), .B(init), .Z(\round_in[0][977] ) );
  AND U10433 ( .A(round_reg[978]), .B(init), .Z(\round_in[0][978] ) );
  AND U10434 ( .A(round_reg[979]), .B(init), .Z(\round_in[0][979] ) );
  NAND U10435 ( .A(init), .B(round_reg[97]), .Z(n4002) );
  NAND U10436 ( .A(n2852), .B(in[97]), .Z(n4001) );
  NAND U10437 ( .A(n4002), .B(n4001), .Z(\round_in[0][97] ) );
  AND U10438 ( .A(round_reg[980]), .B(init), .Z(\round_in[0][980] ) );
  AND U10439 ( .A(round_reg[981]), .B(init), .Z(\round_in[0][981] ) );
  AND U10440 ( .A(round_reg[982]), .B(init), .Z(\round_in[0][982] ) );
  AND U10441 ( .A(round_reg[983]), .B(init), .Z(\round_in[0][983] ) );
  AND U10442 ( .A(round_reg[984]), .B(init), .Z(\round_in[0][984] ) );
  AND U10443 ( .A(round_reg[985]), .B(init), .Z(\round_in[0][985] ) );
  AND U10444 ( .A(round_reg[986]), .B(init), .Z(\round_in[0][986] ) );
  AND U10445 ( .A(round_reg[987]), .B(init), .Z(\round_in[0][987] ) );
  AND U10446 ( .A(round_reg[988]), .B(init), .Z(\round_in[0][988] ) );
  AND U10447 ( .A(round_reg[989]), .B(init), .Z(\round_in[0][989] ) );
  NAND U10448 ( .A(init), .B(round_reg[98]), .Z(n4004) );
  NAND U10449 ( .A(n2852), .B(in[98]), .Z(n4003) );
  NAND U10450 ( .A(n4004), .B(n4003), .Z(\round_in[0][98] ) );
  AND U10451 ( .A(round_reg[990]), .B(init), .Z(\round_in[0][990] ) );
  AND U10452 ( .A(round_reg[991]), .B(init), .Z(\round_in[0][991] ) );
  AND U10453 ( .A(round_reg[992]), .B(init), .Z(\round_in[0][992] ) );
  AND U10454 ( .A(round_reg[993]), .B(init), .Z(\round_in[0][993] ) );
  AND U10455 ( .A(round_reg[994]), .B(init), .Z(\round_in[0][994] ) );
  AND U10456 ( .A(round_reg[995]), .B(init), .Z(\round_in[0][995] ) );
  AND U10457 ( .A(round_reg[996]), .B(init), .Z(\round_in[0][996] ) );
  AND U10458 ( .A(round_reg[997]), .B(init), .Z(\round_in[0][997] ) );
  AND U10459 ( .A(round_reg[998]), .B(init), .Z(\round_in[0][998] ) );
  AND U10460 ( .A(round_reg[999]), .B(init), .Z(\round_in[0][999] ) );
  NAND U10461 ( .A(init), .B(round_reg[99]), .Z(n4006) );
  NAND U10462 ( .A(n2852), .B(in[99]), .Z(n4005) );
  NAND U10463 ( .A(n4006), .B(n4005), .Z(\round_in[0][99] ) );
  NAND U10464 ( .A(init), .B(round_reg[9]), .Z(n4008) );
  NAND U10465 ( .A(n2852), .B(in[9]), .Z(n4007) );
  NAND U10466 ( .A(n4008), .B(n4007), .Z(\round_in[0][9] ) );
  OR U10467 ( .A(\RCONST[1].rconst_/N15 ), .B(rc_i[1]), .Z(n1610) );
endmodule

