
module hamming_N160_CC1 ( clk, rst, x, y, o );
  input [159:0] x;
  input [159:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;

  NAND U161 ( .A(n483), .B(n482), .Z(n1) );
  NAND U162 ( .A(n480), .B(n481), .Z(n2) );
  NAND U163 ( .A(n1), .B(n2), .Z(n750) );
  NAND U164 ( .A(n514), .B(n513), .Z(n3) );
  NAND U165 ( .A(n511), .B(n512), .Z(n4) );
  AND U166 ( .A(n3), .B(n4), .Z(n753) );
  XOR U167 ( .A(n768), .B(n769), .Z(n5) );
  XNOR U168 ( .A(n770), .B(n5), .Z(n740) );
  NAND U169 ( .A(n805), .B(n806), .Z(n6) );
  XOR U170 ( .A(n805), .B(n806), .Z(n7) );
  NANDN U171 ( .A(n804), .B(n7), .Z(n8) );
  NAND U172 ( .A(n6), .B(n8), .Z(n904) );
  NAND U173 ( .A(n502), .B(n503), .Z(n9) );
  XOR U174 ( .A(n502), .B(n503), .Z(n10) );
  NANDN U175 ( .A(n501), .B(n10), .Z(n11) );
  NAND U176 ( .A(n9), .B(n11), .Z(n827) );
  NAND U177 ( .A(n817), .B(n818), .Z(n12) );
  XOR U178 ( .A(n817), .B(n818), .Z(n13) );
  NANDN U179 ( .A(n816), .B(n13), .Z(n14) );
  NAND U180 ( .A(n12), .B(n14), .Z(n924) );
  NAND U181 ( .A(n547), .B(n548), .Z(n15) );
  XOR U182 ( .A(n547), .B(n548), .Z(n16) );
  NANDN U183 ( .A(n546), .B(n16), .Z(n17) );
  NAND U184 ( .A(n15), .B(n17), .Z(n830) );
  XOR U185 ( .A(n689), .B(n688), .Z(n18) );
  NANDN U186 ( .A(n690), .B(n18), .Z(n19) );
  NAND U187 ( .A(n689), .B(n688), .Z(n20) );
  AND U188 ( .A(n19), .B(n20), .Z(n863) );
  NAND U189 ( .A(n926), .B(n925), .Z(n21) );
  XOR U190 ( .A(n926), .B(n925), .Z(n22) );
  NANDN U191 ( .A(n927), .B(n22), .Z(n23) );
  NAND U192 ( .A(n21), .B(n23), .Z(n943) );
  NAND U193 ( .A(n870), .B(n871), .Z(n24) );
  XOR U194 ( .A(n870), .B(n871), .Z(n25) );
  NANDN U195 ( .A(n869), .B(n25), .Z(n26) );
  NAND U196 ( .A(n24), .B(n26), .Z(n974) );
  XNOR U197 ( .A(n557), .B(n556), .Z(n558) );
  XNOR U198 ( .A(n569), .B(n568), .Z(n570) );
  NAND U199 ( .A(n313), .B(n312), .Z(n27) );
  NAND U200 ( .A(n310), .B(n311), .Z(n28) );
  NAND U201 ( .A(n27), .B(n28), .Z(n809) );
  NAND U202 ( .A(n811), .B(n812), .Z(n29) );
  XOR U203 ( .A(n811), .B(n812), .Z(n30) );
  NANDN U204 ( .A(n810), .B(n30), .Z(n31) );
  NAND U205 ( .A(n29), .B(n31), .Z(n905) );
  NAND U206 ( .A(n752), .B(n753), .Z(n32) );
  XOR U207 ( .A(n752), .B(n753), .Z(n33) );
  NANDN U208 ( .A(n751), .B(n33), .Z(n34) );
  NAND U209 ( .A(n32), .B(n34), .Z(n899) );
  NAND U210 ( .A(n724), .B(n725), .Z(n35) );
  XOR U211 ( .A(n724), .B(n725), .Z(n36) );
  NANDN U212 ( .A(n723), .B(n36), .Z(n37) );
  NAND U213 ( .A(n35), .B(n37), .Z(n901) );
  NAND U214 ( .A(n540), .B(n541), .Z(n38) );
  XOR U215 ( .A(n540), .B(n541), .Z(n39) );
  NANDN U216 ( .A(n539), .B(n39), .Z(n40) );
  NAND U217 ( .A(n38), .B(n40), .Z(n741) );
  NAND U218 ( .A(n473), .B(n475), .Z(n41) );
  XOR U219 ( .A(n473), .B(n475), .Z(n42) );
  NAND U220 ( .A(n42), .B(n474), .Z(n43) );
  NAND U221 ( .A(n41), .B(n43), .Z(n841) );
  XOR U222 ( .A(n379), .B(n380), .Z(n44) );
  NANDN U223 ( .A(n381), .B(n44), .Z(n45) );
  NAND U224 ( .A(n379), .B(n380), .Z(n46) );
  AND U225 ( .A(n45), .B(n46), .Z(n793) );
  XOR U226 ( .A(n739), .B(n738), .Z(n47) );
  NAND U227 ( .A(n47), .B(n737), .Z(n48) );
  NAND U228 ( .A(n739), .B(n738), .Z(n49) );
  AND U229 ( .A(n48), .B(n49), .Z(n918) );
  XOR U230 ( .A(n705), .B(n703), .Z(n50) );
  NANDN U231 ( .A(n704), .B(n50), .Z(n51) );
  NAND U232 ( .A(n705), .B(n703), .Z(n52) );
  AND U233 ( .A(n51), .B(n52), .Z(n886) );
  XOR U234 ( .A(n721), .B(n719), .Z(n53) );
  NANDN U235 ( .A(n720), .B(n53), .Z(n54) );
  NAND U236 ( .A(n721), .B(n719), .Z(n55) );
  AND U237 ( .A(n54), .B(n55), .Z(n884) );
  NAND U238 ( .A(n601), .B(n603), .Z(n56) );
  XOR U239 ( .A(n601), .B(n603), .Z(n57) );
  NAND U240 ( .A(n57), .B(n602), .Z(n58) );
  NAND U241 ( .A(n56), .B(n58), .Z(n845) );
  NAND U242 ( .A(n357), .B(n358), .Z(n59) );
  XOR U243 ( .A(n357), .B(n358), .Z(n60) );
  NANDN U244 ( .A(n356), .B(n60), .Z(n61) );
  NAND U245 ( .A(n59), .B(n61), .Z(n686) );
  NAND U246 ( .A(n890), .B(n891), .Z(n62) );
  XOR U247 ( .A(n890), .B(n891), .Z(n63) );
  NANDN U248 ( .A(n889), .B(n63), .Z(n64) );
  NAND U249 ( .A(n62), .B(n64), .Z(n940) );
  NAND U250 ( .A(n552), .B(n553), .Z(n65) );
  NANDN U251 ( .A(n555), .B(n554), .Z(n66) );
  AND U252 ( .A(n65), .B(n66), .Z(n785) );
  NAND U253 ( .A(n929), .B(n930), .Z(n67) );
  XOR U254 ( .A(n929), .B(n930), .Z(n68) );
  NANDN U255 ( .A(n928), .B(n68), .Z(n69) );
  NAND U256 ( .A(n67), .B(n69), .Z(n971) );
  NAND U257 ( .A(n973), .B(n975), .Z(n70) );
  XOR U258 ( .A(n973), .B(n975), .Z(n71) );
  NAND U259 ( .A(n71), .B(n974), .Z(n72) );
  NAND U260 ( .A(n70), .B(n72), .Z(n986) );
  NAND U261 ( .A(n658), .B(n657), .Z(n73) );
  NAND U262 ( .A(n655), .B(n656), .Z(n74) );
  NAND U263 ( .A(n73), .B(n74), .Z(n812) );
  XNOR U264 ( .A(n528), .B(n527), .Z(n529) );
  XNOR U265 ( .A(n534), .B(n533), .Z(n535) );
  NAND U266 ( .A(n757), .B(n758), .Z(n75) );
  XOR U267 ( .A(n757), .B(n758), .Z(n76) );
  NANDN U268 ( .A(n756), .B(n76), .Z(n77) );
  NAND U269 ( .A(n75), .B(n77), .Z(n908) );
  NAND U270 ( .A(n808), .B(n809), .Z(n78) );
  XOR U271 ( .A(n808), .B(n809), .Z(n79) );
  NANDN U272 ( .A(n807), .B(n79), .Z(n80) );
  NAND U273 ( .A(n78), .B(n80), .Z(n906) );
  XOR U274 ( .A(n729), .B(n730), .Z(n81) );
  NANDN U275 ( .A(n731), .B(n81), .Z(n82) );
  NAND U276 ( .A(n729), .B(n730), .Z(n83) );
  AND U277 ( .A(n82), .B(n83), .Z(n902) );
  NAND U278 ( .A(n593), .B(n595), .Z(n84) );
  XOR U279 ( .A(n593), .B(n595), .Z(n85) );
  NAND U280 ( .A(n85), .B(n594), .Z(n86) );
  NAND U281 ( .A(n84), .B(n86), .Z(n836) );
  NAND U282 ( .A(n677), .B(n678), .Z(n87) );
  XOR U283 ( .A(n677), .B(n678), .Z(n88) );
  NANDN U284 ( .A(n676), .B(n88), .Z(n89) );
  NAND U285 ( .A(n87), .B(n89), .Z(n798) );
  NAND U286 ( .A(n476), .B(n478), .Z(n90) );
  XOR U287 ( .A(n476), .B(n478), .Z(n91) );
  NAND U288 ( .A(n91), .B(n477), .Z(n92) );
  NAND U289 ( .A(n90), .B(n92), .Z(n840) );
  XOR U290 ( .A(n442), .B(n443), .Z(n93) );
  NANDN U291 ( .A(n444), .B(n93), .Z(n94) );
  NAND U292 ( .A(n442), .B(n443), .Z(n95) );
  AND U293 ( .A(n94), .B(n95), .Z(n735) );
  NAND U294 ( .A(n717), .B(n718), .Z(n96) );
  XOR U295 ( .A(n717), .B(n718), .Z(n97) );
  NANDN U296 ( .A(n716), .B(n97), .Z(n98) );
  NAND U297 ( .A(n96), .B(n98), .Z(n885) );
  NAND U298 ( .A(n760), .B(n761), .Z(n99) );
  XOR U299 ( .A(n760), .B(n761), .Z(n100) );
  NANDN U300 ( .A(n759), .B(n100), .Z(n101) );
  NAND U301 ( .A(n99), .B(n101), .Z(n880) );
  NAND U302 ( .A(n827), .B(n828), .Z(n102) );
  XOR U303 ( .A(n827), .B(n828), .Z(n103) );
  NANDN U304 ( .A(n826), .B(n103), .Z(n104) );
  NAND U305 ( .A(n102), .B(n104), .Z(n923) );
  NAND U306 ( .A(n605), .B(n606), .Z(n105) );
  XOR U307 ( .A(n605), .B(n606), .Z(n106) );
  NANDN U308 ( .A(n604), .B(n106), .Z(n107) );
  NAND U309 ( .A(n105), .B(n107), .Z(n843) );
  XOR U310 ( .A(n719), .B(n720), .Z(n108) );
  XNOR U311 ( .A(n721), .B(n108), .Z(n821) );
  XOR U312 ( .A(n543), .B(n544), .Z(n109) );
  NANDN U313 ( .A(n545), .B(n109), .Z(n110) );
  NAND U314 ( .A(n543), .B(n544), .Z(n111) );
  AND U315 ( .A(n110), .B(n111), .Z(n831) );
  XOR U316 ( .A(n741), .B(n742), .Z(n112) );
  XNOR U317 ( .A(n743), .B(n112), .Z(n682) );
  XOR U318 ( .A(n687), .B(n685), .Z(n113) );
  NANDN U319 ( .A(n686), .B(n113), .Z(n114) );
  NAND U320 ( .A(n687), .B(n685), .Z(n115) );
  AND U321 ( .A(n114), .B(n115), .Z(n865) );
  NAND U322 ( .A(n886), .B(n888), .Z(n116) );
  XOR U323 ( .A(n886), .B(n888), .Z(n117) );
  NAND U324 ( .A(n117), .B(n887), .Z(n118) );
  NAND U325 ( .A(n116), .B(n118), .Z(n963) );
  NAND U326 ( .A(n867), .B(n868), .Z(n119) );
  XOR U327 ( .A(n867), .B(n868), .Z(n120) );
  NANDN U328 ( .A(n866), .B(n120), .Z(n121) );
  NAND U329 ( .A(n119), .B(n121), .Z(n975) );
  NAND U330 ( .A(n971), .B(n970), .Z(n122) );
  XOR U331 ( .A(n971), .B(n970), .Z(n123) );
  NANDN U332 ( .A(n972), .B(n123), .Z(n124) );
  NAND U333 ( .A(n122), .B(n124), .Z(n987) );
  XNOR U334 ( .A(n407), .B(n406), .Z(n408) );
  XNOR U335 ( .A(n395), .B(n394), .Z(n396) );
  XNOR U336 ( .A(n660), .B(n659), .Z(n661) );
  XNOR U337 ( .A(n401), .B(n400), .Z(n402) );
  NAND U338 ( .A(n498), .B(n500), .Z(n125) );
  XOR U339 ( .A(n498), .B(n500), .Z(n126) );
  NAND U340 ( .A(n126), .B(n499), .Z(n127) );
  NAND U341 ( .A(n125), .B(n127), .Z(n828) );
  XOR U342 ( .A(n726), .B(n727), .Z(n128) );
  NANDN U343 ( .A(n728), .B(n128), .Z(n129) );
  NAND U344 ( .A(n726), .B(n727), .Z(n130) );
  AND U345 ( .A(n129), .B(n130), .Z(n903) );
  NAND U346 ( .A(n749), .B(n750), .Z(n131) );
  XOR U347 ( .A(n749), .B(n750), .Z(n132) );
  NANDN U348 ( .A(n748), .B(n132), .Z(n133) );
  NAND U349 ( .A(n131), .B(n133), .Z(n910) );
  XNOR U350 ( .A(n666), .B(n665), .Z(n667) );
  XNOR U351 ( .A(n291), .B(n290), .Z(n292) );
  XNOR U352 ( .A(n303), .B(n302), .Z(n304) );
  XNOR U353 ( .A(n297), .B(n296), .Z(n298) );
  XNOR U354 ( .A(n383), .B(n382), .Z(n384) );
  XOR U355 ( .A(n713), .B(n714), .Z(n134) );
  XNOR U356 ( .A(n715), .B(n134), .Z(n838) );
  NAND U357 ( .A(n652), .B(n654), .Z(n135) );
  XOR U358 ( .A(n652), .B(n654), .Z(n136) );
  NAND U359 ( .A(n136), .B(n653), .Z(n137) );
  NAND U360 ( .A(n135), .B(n137), .Z(n776) );
  XNOR U361 ( .A(n752), .B(n751), .Z(n138) );
  XNOR U362 ( .A(n753), .B(n138), .Z(n743) );
  XOR U363 ( .A(n703), .B(n704), .Z(n139) );
  XNOR U364 ( .A(n705), .B(n139), .Z(n817) );
  NAND U365 ( .A(n735), .B(n736), .Z(n140) );
  XOR U366 ( .A(n735), .B(n736), .Z(n141) );
  NANDN U367 ( .A(n734), .B(n141), .Z(n142) );
  NAND U368 ( .A(n140), .B(n142), .Z(n917) );
  NAND U369 ( .A(n710), .B(n711), .Z(n143) );
  XOR U370 ( .A(n710), .B(n711), .Z(n144) );
  NANDN U371 ( .A(n709), .B(n144), .Z(n145) );
  NAND U372 ( .A(n143), .B(n145), .Z(n887) );
  XOR U373 ( .A(n770), .B(n768), .Z(n146) );
  NANDN U374 ( .A(n769), .B(n146), .Z(n147) );
  NAND U375 ( .A(n770), .B(n768), .Z(n148) );
  AND U376 ( .A(n147), .B(n148), .Z(n881) );
  NAND U377 ( .A(n920), .B(n921), .Z(n149) );
  XOR U378 ( .A(n920), .B(n921), .Z(n150) );
  NANDN U379 ( .A(n919), .B(n150), .Z(n151) );
  NAND U380 ( .A(n149), .B(n151), .Z(n949) );
  NAND U381 ( .A(n840), .B(n841), .Z(n152) );
  XOR U382 ( .A(n840), .B(n841), .Z(n153) );
  NANDN U383 ( .A(n839), .B(n153), .Z(n154) );
  NAND U384 ( .A(n152), .B(n154), .Z(n926) );
  NAND U385 ( .A(n645), .B(n647), .Z(n155) );
  XOR U386 ( .A(n645), .B(n647), .Z(n156) );
  NAND U387 ( .A(n156), .B(n646), .Z(n157) );
  NAND U388 ( .A(n155), .B(n157), .Z(n819) );
  NAND U389 ( .A(n415), .B(n416), .Z(n158) );
  XOR U390 ( .A(n415), .B(n416), .Z(n159) );
  NANDN U391 ( .A(n414), .B(n159), .Z(n160) );
  NAND U392 ( .A(n158), .B(n160), .Z(n790) );
  NAND U393 ( .A(n883), .B(n885), .Z(n161) );
  XOR U394 ( .A(n883), .B(n885), .Z(n162) );
  NAND U395 ( .A(n162), .B(n884), .Z(n163) );
  NAND U396 ( .A(n161), .B(n163), .Z(n964) );
  NAND U397 ( .A(n864), .B(n865), .Z(n164) );
  XOR U398 ( .A(n864), .B(n865), .Z(n165) );
  NANDN U399 ( .A(n863), .B(n165), .Z(n166) );
  NAND U400 ( .A(n164), .B(n166), .Z(n973) );
  XOR U401 ( .A(n694), .B(n692), .Z(n167) );
  NANDN U402 ( .A(n693), .B(n167), .Z(n168) );
  NAND U403 ( .A(n694), .B(n692), .Z(n169) );
  AND U404 ( .A(n168), .B(n169), .Z(n876) );
  NAND U405 ( .A(n932), .B(n933), .Z(n170) );
  XOR U406 ( .A(n932), .B(n933), .Z(n171) );
  NANDN U407 ( .A(n934), .B(n171), .Z(n172) );
  NAND U408 ( .A(n170), .B(n172), .Z(n977) );
  XNOR U409 ( .A(n997), .B(n998), .Z(n988) );
  XNOR U410 ( .A(n485), .B(n484), .Z(n486) );
  XNOR U411 ( .A(n516), .B(n515), .Z(n517) );
  XNOR U412 ( .A(n330), .B(n329), .Z(n331) );
  XNOR U413 ( .A(n342), .B(n341), .Z(n343) );
  XNOR U414 ( .A(n336), .B(n335), .Z(n337) );
  XNOR U415 ( .A(n373), .B(n372), .Z(n374) );
  XNOR U416 ( .A(n284), .B(n283), .Z(n285) );
  XNOR U417 ( .A(n276), .B(n275), .Z(n277) );
  XNOR U418 ( .A(n621), .B(n620), .Z(n622) );
  XNOR U419 ( .A(n270), .B(n269), .Z(n271) );
  XNOR U420 ( .A(n522), .B(n521), .Z(n523) );
  XNOR U421 ( .A(n389), .B(n388), .Z(n390) );
  NAND U422 ( .A(n674), .B(n675), .Z(n173) );
  XOR U423 ( .A(n674), .B(n675), .Z(n174) );
  NANDN U424 ( .A(n673), .B(n174), .Z(n175) );
  NAND U425 ( .A(n173), .B(n175), .Z(n799) );
  NAND U426 ( .A(n649), .B(n651), .Z(n176) );
  XOR U427 ( .A(n649), .B(n651), .Z(n177) );
  NAND U428 ( .A(n177), .B(n650), .Z(n178) );
  NAND U429 ( .A(n176), .B(n178), .Z(n774) );
  NAND U430 ( .A(n707), .B(n708), .Z(n179) );
  XOR U431 ( .A(n707), .B(n708), .Z(n180) );
  NANDN U432 ( .A(n706), .B(n180), .Z(n181) );
  NAND U433 ( .A(n179), .B(n181), .Z(n888) );
  XOR U434 ( .A(n715), .B(n713), .Z(n182) );
  NANDN U435 ( .A(n714), .B(n182), .Z(n183) );
  NAND U436 ( .A(n715), .B(n713), .Z(n184) );
  AND U437 ( .A(n183), .B(n184), .Z(n883) );
  NAND U438 ( .A(n904), .B(n906), .Z(n185) );
  XOR U439 ( .A(n904), .B(n906), .Z(n186) );
  NAND U440 ( .A(n186), .B(n905), .Z(n187) );
  NAND U441 ( .A(n185), .B(n187), .Z(n914) );
  NAND U442 ( .A(n901), .B(n903), .Z(n188) );
  XOR U443 ( .A(n901), .B(n903), .Z(n189) );
  NAND U444 ( .A(n189), .B(n902), .Z(n190) );
  NAND U445 ( .A(n188), .B(n190), .Z(n955) );
  NAND U446 ( .A(n917), .B(n918), .Z(n191) );
  XOR U447 ( .A(n917), .B(n918), .Z(n192) );
  NANDN U448 ( .A(n916), .B(n192), .Z(n193) );
  NAND U449 ( .A(n191), .B(n193), .Z(n950) );
  NAND U450 ( .A(n837), .B(n838), .Z(n194) );
  XOR U451 ( .A(n837), .B(n838), .Z(n195) );
  NANDN U452 ( .A(n836), .B(n195), .Z(n196) );
  NAND U453 ( .A(n194), .B(n196), .Z(n927) );
  XNOR U454 ( .A(n909), .B(n910), .Z(n891) );
  NAND U455 ( .A(n598), .B(n600), .Z(n197) );
  XOR U456 ( .A(n598), .B(n600), .Z(n198) );
  NAND U457 ( .A(n198), .B(n599), .Z(n199) );
  NAND U458 ( .A(n197), .B(n199), .Z(n842) );
  NAND U459 ( .A(n789), .B(n790), .Z(n200) );
  XOR U460 ( .A(n789), .B(n790), .Z(n201) );
  NANDN U461 ( .A(n788), .B(n201), .Z(n202) );
  NAND U462 ( .A(n200), .B(n202), .Z(n868) );
  NANDN U463 ( .A(n681), .B(n684), .Z(n203) );
  OR U464 ( .A(n684), .B(n683), .Z(n204) );
  NANDN U465 ( .A(n682), .B(n204), .Z(n205) );
  NAND U466 ( .A(n203), .B(n205), .Z(n864) );
  NAND U467 ( .A(n880), .B(n882), .Z(n206) );
  XOR U468 ( .A(n880), .B(n882), .Z(n207) );
  NAND U469 ( .A(n207), .B(n881), .Z(n208) );
  NAND U470 ( .A(n206), .B(n208), .Z(n966) );
  XOR U471 ( .A(n924), .B(n922), .Z(n209) );
  NANDN U472 ( .A(n923), .B(n209), .Z(n210) );
  NAND U473 ( .A(n924), .B(n922), .Z(n211) );
  AND U474 ( .A(n210), .B(n211), .Z(n944) );
  XNOR U475 ( .A(n539), .B(n540), .Z(n212) );
  XNOR U476 ( .A(n541), .B(n212), .Z(n543) );
  NAND U477 ( .A(n550), .B(n551), .Z(n213) );
  XOR U478 ( .A(n550), .B(n551), .Z(n214) );
  NANDN U479 ( .A(n549), .B(n214), .Z(n215) );
  NAND U480 ( .A(n213), .B(n215), .Z(n783) );
  XOR U481 ( .A(n247), .B(n248), .Z(n216) );
  NANDN U482 ( .A(n249), .B(n216), .Z(n217) );
  NAND U483 ( .A(n247), .B(n248), .Z(n218) );
  AND U484 ( .A(n217), .B(n218), .Z(n696) );
  NAND U485 ( .A(n978), .B(n979), .Z(n219) );
  XOR U486 ( .A(n978), .B(n979), .Z(n220) );
  NANDN U487 ( .A(n977), .B(n220), .Z(n221) );
  NAND U488 ( .A(n219), .B(n221), .Z(n990) );
  NAND U489 ( .A(n986), .B(n988), .Z(n222) );
  XOR U490 ( .A(n986), .B(n988), .Z(n223) );
  NAND U491 ( .A(n223), .B(n987), .Z(n224) );
  NAND U492 ( .A(n222), .B(n224), .Z(n1017) );
  XOR U493 ( .A(x[157]), .B(y[157]), .Z(n282) );
  XOR U494 ( .A(x[155]), .B(y[155]), .Z(n281) );
  XOR U495 ( .A(n282), .B(n281), .Z(n658) );
  XOR U496 ( .A(x[147]), .B(y[147]), .Z(n656) );
  XOR U497 ( .A(x[151]), .B(y[151]), .Z(n655) );
  XOR U498 ( .A(n656), .B(n655), .Z(n657) );
  XOR U499 ( .A(n658), .B(n657), .Z(n652) );
  XOR U500 ( .A(x[111]), .B(y[111]), .Z(n363) );
  XOR U501 ( .A(x[113]), .B(y[113]), .Z(n361) );
  XOR U502 ( .A(x[115]), .B(y[115]), .Z(n360) );
  XOR U503 ( .A(n361), .B(n360), .Z(n362) );
  XOR U504 ( .A(n363), .B(n362), .Z(n654) );
  XOR U505 ( .A(x[105]), .B(y[105]), .Z(n420) );
  XOR U506 ( .A(x[109]), .B(y[109]), .Z(n418) );
  XOR U507 ( .A(x[107]), .B(y[107]), .Z(n417) );
  XOR U508 ( .A(n418), .B(n417), .Z(n419) );
  XOR U509 ( .A(n420), .B(n419), .Z(n653) );
  XNOR U510 ( .A(n654), .B(n653), .Z(n225) );
  XOR U511 ( .A(n652), .B(n225), .Z(n438) );
  XOR U512 ( .A(x[135]), .B(y[135]), .Z(n565) );
  XOR U513 ( .A(x[139]), .B(y[139]), .Z(n562) );
  XNOR U514 ( .A(x[137]), .B(y[137]), .Z(n563) );
  XNOR U515 ( .A(n562), .B(n563), .Z(n564) );
  XOR U516 ( .A(n565), .B(n564), .Z(n437) );
  XOR U517 ( .A(x[129]), .B(y[129]), .Z(n508) );
  XOR U518 ( .A(x[133]), .B(y[133]), .Z(n505) );
  XNOR U519 ( .A(x[131]), .B(y[131]), .Z(n506) );
  XNOR U520 ( .A(n505), .B(n506), .Z(n507) );
  XNOR U521 ( .A(n508), .B(n507), .Z(n436) );
  XOR U522 ( .A(n437), .B(n436), .Z(n439) );
  XOR U523 ( .A(n438), .B(n439), .Z(n551) );
  XOR U524 ( .A(x[51]), .B(y[51]), .Z(n425) );
  XOR U525 ( .A(x[55]), .B(y[55]), .Z(n423) );
  XNOR U526 ( .A(x[53]), .B(y[53]), .Z(n424) );
  XOR U527 ( .A(n423), .B(n424), .Z(n426) );
  XNOR U528 ( .A(n425), .B(n426), .Z(n678) );
  XOR U529 ( .A(x[45]), .B(y[45]), .Z(n431) );
  XOR U530 ( .A(x[49]), .B(y[49]), .Z(n429) );
  XNOR U531 ( .A(x[47]), .B(y[47]), .Z(n430) );
  XOR U532 ( .A(n429), .B(n430), .Z(n432) );
  XNOR U533 ( .A(n431), .B(n432), .Z(n677) );
  XOR U534 ( .A(x[39]), .B(y[39]), .Z(n368) );
  XOR U535 ( .A(x[43]), .B(y[43]), .Z(n366) );
  XNOR U536 ( .A(x[41]), .B(y[41]), .Z(n367) );
  XOR U537 ( .A(n366), .B(n367), .Z(n369) );
  XOR U538 ( .A(n368), .B(n369), .Z(n676) );
  XOR U539 ( .A(n677), .B(n676), .Z(n226) );
  XNOR U540 ( .A(n678), .B(n226), .Z(n550) );
  XOR U541 ( .A(x[81]), .B(y[81]), .Z(n385) );
  XOR U542 ( .A(x[85]), .B(y[85]), .Z(n382) );
  XNOR U543 ( .A(x[83]), .B(y[83]), .Z(n383) );
  XOR U544 ( .A(n385), .B(n384), .Z(n601) );
  XOR U545 ( .A(x[87]), .B(y[87]), .Z(n524) );
  XOR U546 ( .A(x[91]), .B(y[91]), .Z(n521) );
  XNOR U547 ( .A(x[89]), .B(y[89]), .Z(n522) );
  XOR U548 ( .A(n524), .B(n523), .Z(n603) );
  XOR U549 ( .A(x[75]), .B(y[75]), .Z(n391) );
  XOR U550 ( .A(x[79]), .B(y[79]), .Z(n388) );
  XNOR U551 ( .A(x[77]), .B(y[77]), .Z(n389) );
  XOR U552 ( .A(n391), .B(n390), .Z(n602) );
  XNOR U553 ( .A(n603), .B(n602), .Z(n227) );
  XOR U554 ( .A(n601), .B(n227), .Z(n549) );
  XOR U555 ( .A(n550), .B(n549), .Z(n228) );
  XOR U556 ( .A(n551), .B(n228), .Z(n448) );
  XOR U557 ( .A(x[92]), .B(y[92]), .Z(n258) );
  XOR U558 ( .A(x[154]), .B(y[154]), .Z(n256) );
  XNOR U559 ( .A(x[90]), .B(y[90]), .Z(n257) );
  XOR U560 ( .A(n256), .B(n257), .Z(n259) );
  XOR U561 ( .A(n258), .B(n259), .Z(n443) );
  XOR U562 ( .A(x[88]), .B(y[88]), .Z(n252) );
  XOR U563 ( .A(x[156]), .B(y[156]), .Z(n250) );
  XNOR U564 ( .A(x[86]), .B(y[86]), .Z(n251) );
  XOR U565 ( .A(n250), .B(n251), .Z(n253) );
  XNOR U566 ( .A(n252), .B(n253), .Z(n444) );
  XOR U567 ( .A(x[96]), .B(y[96]), .Z(n264) );
  XOR U568 ( .A(x[152]), .B(y[152]), .Z(n262) );
  XNOR U569 ( .A(x[94]), .B(y[94]), .Z(n263) );
  XOR U570 ( .A(n262), .B(n263), .Z(n265) );
  XOR U571 ( .A(n264), .B(n265), .Z(n442) );
  XOR U572 ( .A(n444), .B(n442), .Z(n229) );
  XOR U573 ( .A(n443), .B(n229), .Z(n415) );
  XOR U574 ( .A(x[104]), .B(y[104]), .Z(n634) );
  XOR U575 ( .A(x[148]), .B(y[148]), .Z(n632) );
  XNOR U576 ( .A(x[102]), .B(y[102]), .Z(n633) );
  XOR U577 ( .A(n632), .B(n633), .Z(n635) );
  XOR U578 ( .A(n634), .B(n635), .Z(n380) );
  XOR U579 ( .A(x[100]), .B(y[100]), .Z(n628) );
  XOR U580 ( .A(x[150]), .B(y[150]), .Z(n626) );
  XNOR U581 ( .A(x[98]), .B(y[98]), .Z(n627) );
  XOR U582 ( .A(n626), .B(n627), .Z(n629) );
  XNOR U583 ( .A(n628), .B(n629), .Z(n381) );
  XOR U584 ( .A(x[108]), .B(y[108]), .Z(n640) );
  XOR U585 ( .A(x[146]), .B(y[146]), .Z(n638) );
  XNOR U586 ( .A(x[106]), .B(y[106]), .Z(n639) );
  XOR U587 ( .A(n638), .B(n639), .Z(n641) );
  XOR U588 ( .A(n640), .B(n641), .Z(n379) );
  XOR U589 ( .A(n381), .B(n379), .Z(n230) );
  XOR U590 ( .A(n380), .B(n230), .Z(n416) );
  XOR U591 ( .A(x[80]), .B(y[80]), .Z(n338) );
  XOR U592 ( .A(x[78]), .B(y[78]), .Z(n335) );
  XNOR U593 ( .A(x[76]), .B(y[76]), .Z(n336) );
  XOR U594 ( .A(n338), .B(n337), .Z(n476) );
  XOR U595 ( .A(x[74]), .B(y[74]), .Z(n332) );
  XOR U596 ( .A(x[72]), .B(y[72]), .Z(n329) );
  XNOR U597 ( .A(x[70]), .B(y[70]), .Z(n330) );
  XOR U598 ( .A(n332), .B(n331), .Z(n478) );
  XOR U599 ( .A(x[84]), .B(y[84]), .Z(n344) );
  XOR U600 ( .A(x[158]), .B(y[158]), .Z(n341) );
  XNOR U601 ( .A(x[82]), .B(y[82]), .Z(n342) );
  XOR U602 ( .A(n344), .B(n343), .Z(n477) );
  XNOR U603 ( .A(n478), .B(n477), .Z(n231) );
  XOR U604 ( .A(n476), .B(n231), .Z(n414) );
  XOR U605 ( .A(n416), .B(n414), .Z(n232) );
  XOR U606 ( .A(n415), .B(n232), .Z(n248) );
  XOR U607 ( .A(x[99]), .B(y[99]), .Z(n403) );
  XOR U608 ( .A(x[103]), .B(y[103]), .Z(n400) );
  XNOR U609 ( .A(x[101]), .B(y[101]), .Z(n401) );
  XOR U610 ( .A(n403), .B(n402), .Z(n600) );
  XOR U611 ( .A(x[93]), .B(y[93]), .Z(n536) );
  XOR U612 ( .A(x[97]), .B(y[97]), .Z(n533) );
  XNOR U613 ( .A(x[95]), .B(y[95]), .Z(n534) );
  XOR U614 ( .A(n536), .B(n535), .Z(n599) );
  XOR U615 ( .A(x[149]), .B(y[149]), .Z(n662) );
  XOR U616 ( .A(x[159]), .B(y[159]), .Z(n659) );
  XNOR U617 ( .A(x[153]), .B(y[153]), .Z(n660) );
  XOR U618 ( .A(n662), .B(n661), .Z(n598) );
  XNOR U619 ( .A(n599), .B(n598), .Z(n233) );
  XOR U620 ( .A(n600), .B(n233), .Z(n548) );
  XOR U621 ( .A(x[117]), .B(y[117]), .Z(n463) );
  XOR U622 ( .A(x[121]), .B(y[121]), .Z(n460) );
  XNOR U623 ( .A(x[119]), .B(y[119]), .Z(n461) );
  XNOR U624 ( .A(n460), .B(n461), .Z(n462) );
  XOR U625 ( .A(n463), .B(n462), .Z(n348) );
  XOR U626 ( .A(x[123]), .B(y[123]), .Z(n487) );
  XOR U627 ( .A(x[127]), .B(y[127]), .Z(n484) );
  XNOR U628 ( .A(x[125]), .B(y[125]), .Z(n485) );
  XOR U629 ( .A(n487), .B(n486), .Z(n352) );
  XOR U630 ( .A(x[141]), .B(y[141]), .Z(n588) );
  XOR U631 ( .A(x[145]), .B(y[145]), .Z(n586) );
  XNOR U632 ( .A(x[143]), .B(y[143]), .Z(n587) );
  XOR U633 ( .A(n586), .B(n587), .Z(n589) );
  XOR U634 ( .A(n588), .B(n589), .Z(n347) );
  XOR U635 ( .A(n352), .B(n347), .Z(n234) );
  XOR U636 ( .A(n348), .B(n234), .Z(n547) );
  XOR U637 ( .A(x[63]), .B(y[63]), .Z(n397) );
  XOR U638 ( .A(x[67]), .B(y[67]), .Z(n394) );
  XNOR U639 ( .A(x[65]), .B(y[65]), .Z(n395) );
  XOR U640 ( .A(n397), .B(n396), .Z(n674) );
  XOR U641 ( .A(x[69]), .B(y[69]), .Z(n530) );
  XOR U642 ( .A(x[73]), .B(y[73]), .Z(n527) );
  XNOR U643 ( .A(x[71]), .B(y[71]), .Z(n528) );
  XOR U644 ( .A(n530), .B(n529), .Z(n675) );
  XOR U645 ( .A(x[57]), .B(y[57]), .Z(n409) );
  XOR U646 ( .A(x[61]), .B(y[61]), .Z(n406) );
  XNOR U647 ( .A(x[59]), .B(y[59]), .Z(n407) );
  XNOR U648 ( .A(n409), .B(n408), .Z(n673) );
  XOR U649 ( .A(n675), .B(n673), .Z(n235) );
  XNOR U650 ( .A(n674), .B(n235), .Z(n546) );
  XOR U651 ( .A(n547), .B(n546), .Z(n236) );
  XOR U652 ( .A(n548), .B(n236), .Z(n249) );
  XOR U653 ( .A(x[2]), .B(y[2]), .Z(n518) );
  XOR U654 ( .A(x[1]), .B(y[1]), .Z(n515) );
  XNOR U655 ( .A(x[0]), .B(y[0]), .Z(n516) );
  XOR U656 ( .A(n518), .B(n517), .Z(n595) );
  XOR U657 ( .A(x[14]), .B(y[14]), .Z(n571) );
  XOR U658 ( .A(x[12]), .B(y[12]), .Z(n568) );
  XNOR U659 ( .A(x[10]), .B(y[10]), .Z(n569) );
  XOR U660 ( .A(n571), .B(n570), .Z(n594) );
  XOR U661 ( .A(x[8]), .B(y[8]), .Z(n559) );
  XOR U662 ( .A(x[6]), .B(y[6]), .Z(n556) );
  XNOR U663 ( .A(x[4]), .B(y[4]), .Z(n557) );
  XOR U664 ( .A(n559), .B(n558), .Z(n593) );
  XNOR U665 ( .A(n594), .B(n593), .Z(n237) );
  XNOR U666 ( .A(n595), .B(n237), .Z(n358) );
  XOR U667 ( .A(x[33]), .B(y[33]), .Z(n375) );
  XOR U668 ( .A(x[37]), .B(y[37]), .Z(n372) );
  XNOR U669 ( .A(x[35]), .B(y[35]), .Z(n373) );
  XOR U670 ( .A(n375), .B(n374), .Z(n606) );
  XOR U671 ( .A(x[21]), .B(y[21]), .Z(n468) );
  XOR U672 ( .A(x[25]), .B(y[25]), .Z(n466) );
  XNOR U673 ( .A(x[23]), .B(y[23]), .Z(n467) );
  XOR U674 ( .A(n466), .B(n467), .Z(n469) );
  XNOR U675 ( .A(n468), .B(n469), .Z(n605) );
  XOR U676 ( .A(x[27]), .B(y[27]), .Z(n456) );
  XOR U677 ( .A(x[31]), .B(y[31]), .Z(n454) );
  XNOR U678 ( .A(x[29]), .B(y[29]), .Z(n455) );
  XOR U679 ( .A(n454), .B(n455), .Z(n457) );
  XOR U680 ( .A(n456), .B(n457), .Z(n604) );
  XOR U681 ( .A(n605), .B(n604), .Z(n238) );
  XNOR U682 ( .A(n606), .B(n238), .Z(n357) );
  XOR U683 ( .A(x[9]), .B(y[9]), .Z(n493) );
  XOR U684 ( .A(x[13]), .B(y[13]), .Z(n491) );
  XOR U685 ( .A(x[11]), .B(y[11]), .Z(n490) );
  XOR U686 ( .A(n491), .B(n490), .Z(n492) );
  XOR U687 ( .A(n493), .B(n492), .Z(n649) );
  XOR U688 ( .A(x[15]), .B(y[15]), .Z(n483) );
  XOR U689 ( .A(x[19]), .B(y[19]), .Z(n481) );
  XOR U690 ( .A(x[17]), .B(y[17]), .Z(n480) );
  XOR U691 ( .A(n481), .B(n480), .Z(n482) );
  XOR U692 ( .A(n483), .B(n482), .Z(n651) );
  XOR U693 ( .A(x[3]), .B(y[3]), .Z(n514) );
  XOR U694 ( .A(x[7]), .B(y[7]), .Z(n512) );
  XOR U695 ( .A(x[5]), .B(y[5]), .Z(n511) );
  XOR U696 ( .A(n512), .B(n511), .Z(n513) );
  XOR U697 ( .A(n514), .B(n513), .Z(n650) );
  XNOR U698 ( .A(n651), .B(n650), .Z(n239) );
  XOR U699 ( .A(n649), .B(n239), .Z(n356) );
  XOR U700 ( .A(n357), .B(n356), .Z(n240) );
  XOR U701 ( .A(n358), .B(n240), .Z(n247) );
  XOR U702 ( .A(n249), .B(n247), .Z(n241) );
  XOR U703 ( .A(n248), .B(n241), .Z(n449) );
  XNOR U704 ( .A(n448), .B(n449), .Z(n451) );
  XOR U705 ( .A(x[44]), .B(y[44]), .Z(n317) );
  XOR U706 ( .A(x[42]), .B(y[42]), .Z(n315) );
  XOR U707 ( .A(x[40]), .B(y[40]), .Z(n314) );
  XOR U708 ( .A(n315), .B(n314), .Z(n316) );
  XOR U709 ( .A(n317), .B(n316), .Z(n498) );
  XOR U710 ( .A(x[38]), .B(y[38]), .Z(n313) );
  XOR U711 ( .A(x[36]), .B(y[36]), .Z(n311) );
  XOR U712 ( .A(x[34]), .B(y[34]), .Z(n310) );
  XOR U713 ( .A(n311), .B(n310), .Z(n312) );
  XOR U714 ( .A(n313), .B(n312), .Z(n500) );
  XOR U715 ( .A(x[50]), .B(y[50]), .Z(n324) );
  XOR U716 ( .A(x[48]), .B(y[48]), .Z(n322) );
  XOR U717 ( .A(x[46]), .B(y[46]), .Z(n321) );
  XOR U718 ( .A(n322), .B(n321), .Z(n323) );
  XOR U719 ( .A(n324), .B(n323), .Z(n499) );
  XNOR U720 ( .A(n500), .B(n499), .Z(n242) );
  XOR U721 ( .A(n498), .B(n242), .Z(n544) );
  XOR U722 ( .A(x[62]), .B(y[62]), .Z(n299) );
  XOR U723 ( .A(x[60]), .B(y[60]), .Z(n296) );
  XNOR U724 ( .A(x[58]), .B(y[58]), .Z(n297) );
  XOR U725 ( .A(n299), .B(n298), .Z(n473) );
  XOR U726 ( .A(x[56]), .B(y[56]), .Z(n293) );
  XOR U727 ( .A(x[54]), .B(y[54]), .Z(n290) );
  XNOR U728 ( .A(x[52]), .B(y[52]), .Z(n291) );
  XOR U729 ( .A(n293), .B(n292), .Z(n475) );
  XOR U730 ( .A(x[68]), .B(y[68]), .Z(n305) );
  XOR U731 ( .A(x[66]), .B(y[66]), .Z(n302) );
  XNOR U732 ( .A(x[64]), .B(y[64]), .Z(n303) );
  XOR U733 ( .A(n305), .B(n304), .Z(n474) );
  XNOR U734 ( .A(n475), .B(n474), .Z(n243) );
  XNOR U735 ( .A(n473), .B(n243), .Z(n545) );
  XOR U736 ( .A(x[26]), .B(y[26]), .Z(n576) );
  XOR U737 ( .A(x[24]), .B(y[24]), .Z(n574) );
  XNOR U738 ( .A(x[22]), .B(y[22]), .Z(n575) );
  XOR U739 ( .A(n574), .B(n575), .Z(n577) );
  XNOR U740 ( .A(n576), .B(n577), .Z(n541) );
  XOR U741 ( .A(x[32]), .B(y[32]), .Z(n668) );
  XOR U742 ( .A(x[30]), .B(y[30]), .Z(n665) );
  XNOR U743 ( .A(x[28]), .B(y[28]), .Z(n666) );
  XOR U744 ( .A(n668), .B(n667), .Z(n540) );
  XOR U745 ( .A(x[20]), .B(y[20]), .Z(n582) );
  XOR U746 ( .A(x[18]), .B(y[18]), .Z(n580) );
  XNOR U747 ( .A(x[16]), .B(y[16]), .Z(n581) );
  XOR U748 ( .A(n580), .B(n581), .Z(n583) );
  XOR U749 ( .A(n582), .B(n583), .Z(n539) );
  XOR U750 ( .A(n545), .B(n543), .Z(n244) );
  XOR U751 ( .A(n544), .B(n244), .Z(n555) );
  XOR U752 ( .A(x[124]), .B(y[124]), .Z(n272) );
  XOR U753 ( .A(x[138]), .B(y[138]), .Z(n269) );
  XNOR U754 ( .A(x[122]), .B(y[122]), .Z(n270) );
  XOR U755 ( .A(n272), .B(n271), .Z(n645) );
  XOR U756 ( .A(x[120]), .B(y[120]), .Z(n623) );
  XOR U757 ( .A(x[140]), .B(y[140]), .Z(n620) );
  XNOR U758 ( .A(x[118]), .B(y[118]), .Z(n621) );
  XOR U759 ( .A(n623), .B(n622), .Z(n647) );
  XOR U760 ( .A(x[132]), .B(y[132]), .Z(n278) );
  XOR U761 ( .A(x[136]), .B(y[136]), .Z(n275) );
  XNOR U762 ( .A(x[134]), .B(y[134]), .Z(n276) );
  XOR U763 ( .A(n278), .B(n277), .Z(n646) );
  XNOR U764 ( .A(n647), .B(n646), .Z(n245) );
  XOR U765 ( .A(n645), .B(n245), .Z(n552) );
  XOR U766 ( .A(x[116]), .B(y[116]), .Z(n616) );
  XOR U767 ( .A(x[142]), .B(y[142]), .Z(n614) );
  XNOR U768 ( .A(x[114]), .B(y[114]), .Z(n615) );
  XOR U769 ( .A(n614), .B(n615), .Z(n617) );
  XOR U770 ( .A(n616), .B(n617), .Z(n501) );
  XOR U771 ( .A(x[112]), .B(y[112]), .Z(n610) );
  XOR U772 ( .A(x[144]), .B(y[144]), .Z(n608) );
  XNOR U773 ( .A(x[110]), .B(y[110]), .Z(n609) );
  XOR U774 ( .A(n608), .B(n609), .Z(n611) );
  XNOR U775 ( .A(n610), .B(n611), .Z(n503) );
  XOR U776 ( .A(x[128]), .B(y[128]), .Z(n286) );
  XOR U777 ( .A(x[130]), .B(y[130]), .Z(n283) );
  XNOR U778 ( .A(x[126]), .B(y[126]), .Z(n284) );
  XOR U779 ( .A(n286), .B(n285), .Z(n502) );
  XNOR U780 ( .A(n503), .B(n502), .Z(n246) );
  XNOR U781 ( .A(n501), .B(n246), .Z(n553) );
  XOR U782 ( .A(n552), .B(n553), .Z(n554) );
  XNOR U783 ( .A(n555), .B(n554), .Z(n450) );
  XNOR U784 ( .A(n451), .B(n450), .Z(o[0]) );
  NANDN U785 ( .A(n251), .B(n250), .Z(n255) );
  NANDN U786 ( .A(n253), .B(n252), .Z(n254) );
  NAND U787 ( .A(n255), .B(n254), .Z(n711) );
  NANDN U788 ( .A(n257), .B(n256), .Z(n261) );
  NANDN U789 ( .A(n259), .B(n258), .Z(n260) );
  NAND U790 ( .A(n261), .B(n260), .Z(n710) );
  NANDN U791 ( .A(n263), .B(n262), .Z(n267) );
  NANDN U792 ( .A(n265), .B(n264), .Z(n266) );
  AND U793 ( .A(n267), .B(n266), .Z(n709) );
  XOR U794 ( .A(n710), .B(n709), .Z(n268) );
  XOR U795 ( .A(n711), .B(n268), .Z(n739) );
  NANDN U796 ( .A(n270), .B(n269), .Z(n274) );
  NAND U797 ( .A(n272), .B(n271), .Z(n273) );
  AND U798 ( .A(n274), .B(n273), .Z(n756) );
  NANDN U799 ( .A(n276), .B(n275), .Z(n280) );
  NAND U800 ( .A(n278), .B(n277), .Z(n279) );
  AND U801 ( .A(n280), .B(n279), .Z(n754) );
  AND U802 ( .A(n282), .B(n281), .Z(n755) );
  XNOR U803 ( .A(n754), .B(n755), .Z(n758) );
  NANDN U804 ( .A(n284), .B(n283), .Z(n288) );
  NAND U805 ( .A(n286), .B(n285), .Z(n287) );
  NAND U806 ( .A(n288), .B(n287), .Z(n757) );
  XOR U807 ( .A(n758), .B(n757), .Z(n289) );
  XOR U808 ( .A(n756), .B(n289), .Z(n737) );
  NANDN U809 ( .A(n291), .B(n290), .Z(n295) );
  NAND U810 ( .A(n293), .B(n292), .Z(n294) );
  NAND U811 ( .A(n295), .B(n294), .Z(n708) );
  NANDN U812 ( .A(n297), .B(n296), .Z(n301) );
  NAND U813 ( .A(n299), .B(n298), .Z(n300) );
  NAND U814 ( .A(n301), .B(n300), .Z(n707) );
  NANDN U815 ( .A(n303), .B(n302), .Z(n307) );
  NAND U816 ( .A(n305), .B(n304), .Z(n306) );
  AND U817 ( .A(n307), .B(n306), .Z(n706) );
  XOR U818 ( .A(n707), .B(n706), .Z(n308) );
  XOR U819 ( .A(n708), .B(n308), .Z(n738) );
  XOR U820 ( .A(n737), .B(n738), .Z(n309) );
  XOR U821 ( .A(n739), .B(n309), .Z(n685) );
  NAND U822 ( .A(n315), .B(n314), .Z(n320) );
  IV U823 ( .A(n316), .Z(n318) );
  NANDN U824 ( .A(n318), .B(n317), .Z(n319) );
  NAND U825 ( .A(n320), .B(n319), .Z(n808) );
  NAND U826 ( .A(n322), .B(n321), .Z(n327) );
  IV U827 ( .A(n323), .Z(n325) );
  NANDN U828 ( .A(n325), .B(n324), .Z(n326) );
  AND U829 ( .A(n327), .B(n326), .Z(n807) );
  XOR U830 ( .A(n808), .B(n807), .Z(n328) );
  XOR U831 ( .A(n809), .B(n328), .Z(n818) );
  NANDN U832 ( .A(n330), .B(n329), .Z(n334) );
  NAND U833 ( .A(n332), .B(n331), .Z(n333) );
  AND U834 ( .A(n334), .B(n333), .Z(n705) );
  NANDN U835 ( .A(n336), .B(n335), .Z(n340) );
  NAND U836 ( .A(n338), .B(n337), .Z(n339) );
  NAND U837 ( .A(n340), .B(n339), .Z(n704) );
  NANDN U838 ( .A(n342), .B(n341), .Z(n346) );
  NAND U839 ( .A(n344), .B(n343), .Z(n345) );
  AND U840 ( .A(n346), .B(n345), .Z(n703) );
  IV U841 ( .A(n347), .Z(n350) );
  IV U842 ( .A(n348), .Z(n349) );
  NANDN U843 ( .A(n350), .B(n349), .Z(n354) );
  ANDN U844 ( .B(n350), .A(n349), .Z(n351) );
  OR U845 ( .A(n352), .B(n351), .Z(n353) );
  AND U846 ( .A(n354), .B(n353), .Z(n816) );
  XNOR U847 ( .A(n817), .B(n816), .Z(n355) );
  XOR U848 ( .A(n818), .B(n355), .Z(n687) );
  XNOR U849 ( .A(n687), .B(n686), .Z(n359) );
  XOR U850 ( .A(n685), .B(n359), .Z(n699) );
  NAND U851 ( .A(n361), .B(n360), .Z(n365) );
  NAND U852 ( .A(n363), .B(n362), .Z(n364) );
  NAND U853 ( .A(n365), .B(n364), .Z(n727) );
  NANDN U854 ( .A(n367), .B(n366), .Z(n371) );
  NANDN U855 ( .A(n369), .B(n368), .Z(n370) );
  AND U856 ( .A(n371), .B(n370), .Z(n728) );
  NANDN U857 ( .A(n373), .B(n372), .Z(n377) );
  NAND U858 ( .A(n375), .B(n374), .Z(n376) );
  NAND U859 ( .A(n377), .B(n376), .Z(n726) );
  XOR U860 ( .A(n728), .B(n726), .Z(n378) );
  XOR U861 ( .A(n727), .B(n378), .Z(n794) );
  NANDN U862 ( .A(n383), .B(n382), .Z(n387) );
  NAND U863 ( .A(n385), .B(n384), .Z(n386) );
  AND U864 ( .A(n387), .B(n386), .Z(n762) );
  NANDN U865 ( .A(n389), .B(n388), .Z(n393) );
  NAND U866 ( .A(n391), .B(n390), .Z(n392) );
  NAND U867 ( .A(n393), .B(n392), .Z(n763) );
  XNOR U868 ( .A(n762), .B(n763), .Z(n765) );
  NANDN U869 ( .A(n395), .B(n394), .Z(n399) );
  NAND U870 ( .A(n397), .B(n396), .Z(n398) );
  NAND U871 ( .A(n399), .B(n398), .Z(n718) );
  NANDN U872 ( .A(n401), .B(n400), .Z(n405) );
  NAND U873 ( .A(n403), .B(n402), .Z(n404) );
  NAND U874 ( .A(n405), .B(n404), .Z(n717) );
  NANDN U875 ( .A(n407), .B(n406), .Z(n411) );
  NAND U876 ( .A(n409), .B(n408), .Z(n410) );
  AND U877 ( .A(n411), .B(n410), .Z(n716) );
  XOR U878 ( .A(n717), .B(n716), .Z(n412) );
  XOR U879 ( .A(n718), .B(n412), .Z(n764) );
  XOR U880 ( .A(n765), .B(n764), .Z(n792) );
  IV U881 ( .A(n792), .Z(n791) );
  XOR U882 ( .A(n793), .B(n791), .Z(n413) );
  XOR U883 ( .A(n794), .B(n413), .Z(n788) );
  NAND U884 ( .A(n418), .B(n417), .Z(n422) );
  NAND U885 ( .A(n420), .B(n419), .Z(n421) );
  NAND U886 ( .A(n422), .B(n421), .Z(n730) );
  NANDN U887 ( .A(n424), .B(n423), .Z(n428) );
  NANDN U888 ( .A(n426), .B(n425), .Z(n427) );
  AND U889 ( .A(n428), .B(n427), .Z(n731) );
  NANDN U890 ( .A(n430), .B(n429), .Z(n434) );
  NANDN U891 ( .A(n432), .B(n431), .Z(n433) );
  NAND U892 ( .A(n434), .B(n433), .Z(n729) );
  XOR U893 ( .A(n731), .B(n729), .Z(n435) );
  XOR U894 ( .A(n730), .B(n435), .Z(n734) );
  NANDN U895 ( .A(n437), .B(n436), .Z(n441) );
  NANDN U896 ( .A(n439), .B(n438), .Z(n440) );
  AND U897 ( .A(n441), .B(n440), .Z(n736) );
  XNOR U898 ( .A(n736), .B(n735), .Z(n445) );
  XOR U899 ( .A(n734), .B(n445), .Z(n789) );
  XNOR U900 ( .A(n790), .B(n789), .Z(n446) );
  XOR U901 ( .A(n788), .B(n446), .Z(n697) );
  IV U902 ( .A(n697), .Z(n695) );
  XOR U903 ( .A(n699), .B(n695), .Z(n447) );
  XNOR U904 ( .A(n696), .B(n447), .Z(n851) );
  NANDN U905 ( .A(n449), .B(n448), .Z(n453) );
  NAND U906 ( .A(n451), .B(n450), .Z(n452) );
  AND U907 ( .A(n453), .B(n452), .Z(n852) );
  XNOR U908 ( .A(n851), .B(n852), .Z(n854) );
  NANDN U909 ( .A(n455), .B(n454), .Z(n459) );
  NANDN U910 ( .A(n457), .B(n456), .Z(n458) );
  NAND U911 ( .A(n459), .B(n458), .Z(n761) );
  NANDN U912 ( .A(n461), .B(n460), .Z(n465) );
  NAND U913 ( .A(n463), .B(n462), .Z(n464) );
  NAND U914 ( .A(n465), .B(n464), .Z(n760) );
  NANDN U915 ( .A(n467), .B(n466), .Z(n471) );
  NANDN U916 ( .A(n469), .B(n468), .Z(n470) );
  AND U917 ( .A(n471), .B(n470), .Z(n759) );
  XOR U918 ( .A(n760), .B(n759), .Z(n472) );
  XOR U919 ( .A(n761), .B(n472), .Z(n839) );
  XNOR U920 ( .A(n841), .B(n840), .Z(n479) );
  XOR U921 ( .A(n839), .B(n479), .Z(n684) );
  NANDN U922 ( .A(n485), .B(n484), .Z(n489) );
  NAND U923 ( .A(n487), .B(n486), .Z(n488) );
  NAND U924 ( .A(n489), .B(n488), .Z(n749) );
  NAND U925 ( .A(n491), .B(n490), .Z(n496) );
  IV U926 ( .A(n492), .Z(n494) );
  NANDN U927 ( .A(n494), .B(n493), .Z(n495) );
  AND U928 ( .A(n496), .B(n495), .Z(n748) );
  XOR U929 ( .A(n749), .B(n748), .Z(n497) );
  XOR U930 ( .A(n750), .B(n497), .Z(n826) );
  XNOR U931 ( .A(n828), .B(n827), .Z(n504) );
  XOR U932 ( .A(n826), .B(n504), .Z(n683) );
  IV U933 ( .A(n683), .Z(n681) );
  NANDN U934 ( .A(n506), .B(n505), .Z(n510) );
  NAND U935 ( .A(n508), .B(n507), .Z(n509) );
  NAND U936 ( .A(n510), .B(n509), .Z(n751) );
  NANDN U937 ( .A(n516), .B(n515), .Z(n520) );
  NAND U938 ( .A(n518), .B(n517), .Z(n519) );
  AND U939 ( .A(n520), .B(n519), .Z(n752) );
  NANDN U940 ( .A(n522), .B(n521), .Z(n526) );
  NAND U941 ( .A(n524), .B(n523), .Z(n525) );
  AND U942 ( .A(n526), .B(n525), .Z(n770) );
  NANDN U943 ( .A(n528), .B(n527), .Z(n532) );
  NAND U944 ( .A(n530), .B(n529), .Z(n531) );
  NAND U945 ( .A(n532), .B(n531), .Z(n769) );
  NANDN U946 ( .A(n534), .B(n533), .Z(n538) );
  NAND U947 ( .A(n536), .B(n535), .Z(n537) );
  AND U948 ( .A(n538), .B(n537), .Z(n768) );
  IV U949 ( .A(n740), .Z(n742) );
  XOR U950 ( .A(n681), .B(n682), .Z(n542) );
  XOR U951 ( .A(n684), .B(n542), .Z(n833) );
  XNOR U952 ( .A(n831), .B(n830), .Z(n832) );
  XOR U953 ( .A(n833), .B(n832), .Z(n692) );
  NANDN U954 ( .A(n557), .B(n556), .Z(n561) );
  NAND U955 ( .A(n559), .B(n558), .Z(n560) );
  AND U956 ( .A(n561), .B(n560), .Z(n715) );
  NANDN U957 ( .A(n563), .B(n562), .Z(n567) );
  NAND U958 ( .A(n565), .B(n564), .Z(n566) );
  NAND U959 ( .A(n567), .B(n566), .Z(n714) );
  NANDN U960 ( .A(n569), .B(n568), .Z(n573) );
  NAND U961 ( .A(n571), .B(n570), .Z(n572) );
  AND U962 ( .A(n573), .B(n572), .Z(n713) );
  NANDN U963 ( .A(n575), .B(n574), .Z(n579) );
  NANDN U964 ( .A(n577), .B(n576), .Z(n578) );
  NAND U965 ( .A(n579), .B(n578), .Z(n723) );
  NANDN U966 ( .A(n581), .B(n580), .Z(n585) );
  NANDN U967 ( .A(n583), .B(n582), .Z(n584) );
  AND U968 ( .A(n585), .B(n584), .Z(n725) );
  NANDN U969 ( .A(n587), .B(n586), .Z(n591) );
  NANDN U970 ( .A(n589), .B(n588), .Z(n590) );
  AND U971 ( .A(n591), .B(n590), .Z(n724) );
  XNOR U972 ( .A(n725), .B(n724), .Z(n592) );
  XOR U973 ( .A(n723), .B(n592), .Z(n837) );
  XNOR U974 ( .A(n837), .B(n836), .Z(n596) );
  XOR U975 ( .A(n838), .B(n596), .Z(n782) );
  IV U976 ( .A(n782), .Z(n781) );
  XOR U977 ( .A(n785), .B(n781), .Z(n597) );
  XOR U978 ( .A(n783), .B(n597), .Z(n694) );
  XOR U979 ( .A(n845), .B(n843), .Z(n607) );
  XOR U980 ( .A(n842), .B(n607), .Z(n689) );
  NANDN U981 ( .A(n609), .B(n608), .Z(n613) );
  NANDN U982 ( .A(n611), .B(n610), .Z(n612) );
  AND U983 ( .A(n613), .B(n612), .Z(n721) );
  NANDN U984 ( .A(n615), .B(n614), .Z(n619) );
  NANDN U985 ( .A(n617), .B(n616), .Z(n618) );
  NAND U986 ( .A(n619), .B(n618), .Z(n720) );
  NANDN U987 ( .A(n621), .B(n620), .Z(n625) );
  NAND U988 ( .A(n623), .B(n622), .Z(n624) );
  AND U989 ( .A(n625), .B(n624), .Z(n719) );
  NANDN U990 ( .A(n627), .B(n626), .Z(n631) );
  NANDN U991 ( .A(n629), .B(n628), .Z(n630) );
  NAND U992 ( .A(n631), .B(n630), .Z(n806) );
  NANDN U993 ( .A(n633), .B(n632), .Z(n637) );
  NANDN U994 ( .A(n635), .B(n634), .Z(n636) );
  NAND U995 ( .A(n637), .B(n636), .Z(n805) );
  NANDN U996 ( .A(n639), .B(n638), .Z(n643) );
  NANDN U997 ( .A(n641), .B(n640), .Z(n642) );
  AND U998 ( .A(n643), .B(n642), .Z(n804) );
  XOR U999 ( .A(n805), .B(n804), .Z(n644) );
  XOR U1000 ( .A(n806), .B(n644), .Z(n820) );
  XNOR U1001 ( .A(n820), .B(n819), .Z(n648) );
  XOR U1002 ( .A(n821), .B(n648), .Z(n690) );
  NANDN U1003 ( .A(n660), .B(n659), .Z(n664) );
  NAND U1004 ( .A(n662), .B(n661), .Z(n663) );
  NAND U1005 ( .A(n664), .B(n663), .Z(n811) );
  NANDN U1006 ( .A(n666), .B(n665), .Z(n670) );
  NAND U1007 ( .A(n668), .B(n667), .Z(n669) );
  AND U1008 ( .A(n670), .B(n669), .Z(n810) );
  XOR U1009 ( .A(n811), .B(n810), .Z(n671) );
  XOR U1010 ( .A(n812), .B(n671), .Z(n773) );
  IV U1011 ( .A(n773), .Z(n772) );
  XOR U1012 ( .A(n776), .B(n772), .Z(n672) );
  XOR U1013 ( .A(n774), .B(n672), .Z(n801) );
  XOR U1014 ( .A(n799), .B(n798), .Z(n800) );
  XOR U1015 ( .A(n801), .B(n800), .Z(n688) );
  XOR U1016 ( .A(n690), .B(n688), .Z(n679) );
  XOR U1017 ( .A(n689), .B(n679), .Z(n693) );
  XNOR U1018 ( .A(n694), .B(n693), .Z(n680) );
  XNOR U1019 ( .A(n692), .B(n680), .Z(n853) );
  XNOR U1020 ( .A(n854), .B(n853), .Z(o[1]) );
  XOR U1021 ( .A(n865), .B(n863), .Z(n691) );
  XOR U1022 ( .A(n864), .B(n691), .Z(n875) );
  IV U1023 ( .A(n875), .Z(n873) );
  NANDN U1024 ( .A(n695), .B(n696), .Z(n701) );
  NOR U1025 ( .A(n697), .B(n696), .Z(n698) );
  OR U1026 ( .A(n699), .B(n698), .Z(n700) );
  AND U1027 ( .A(n701), .B(n700), .Z(n874) );
  XNOR U1028 ( .A(n876), .B(n874), .Z(n702) );
  XOR U1029 ( .A(n873), .B(n702), .Z(n860) );
  XNOR U1030 ( .A(n888), .B(n887), .Z(n712) );
  XOR U1031 ( .A(n886), .B(n712), .Z(n892) );
  XNOR U1032 ( .A(n885), .B(n884), .Z(n722) );
  XNOR U1033 ( .A(n883), .B(n722), .Z(n895) );
  XOR U1034 ( .A(n903), .B(n902), .Z(n732) );
  XNOR U1035 ( .A(n901), .B(n732), .Z(n893) );
  XOR U1036 ( .A(n895), .B(n893), .Z(n733) );
  XOR U1037 ( .A(n892), .B(n733), .Z(n869) );
  NANDN U1038 ( .A(n740), .B(n741), .Z(n746) );
  NOR U1039 ( .A(n742), .B(n741), .Z(n744) );
  NANDN U1040 ( .A(n744), .B(n743), .Z(n745) );
  AND U1041 ( .A(n746), .B(n745), .Z(n916) );
  XOR U1042 ( .A(n918), .B(n916), .Z(n747) );
  XNOR U1043 ( .A(n917), .B(n747), .Z(n871) );
  ANDN U1044 ( .B(n755), .A(n754), .Z(n900) );
  XOR U1045 ( .A(n899), .B(n900), .Z(n907) );
  XOR U1046 ( .A(n907), .B(n908), .Z(n909) );
  NANDN U1047 ( .A(n763), .B(n762), .Z(n767) );
  NAND U1048 ( .A(n765), .B(n764), .Z(n766) );
  AND U1049 ( .A(n767), .B(n766), .Z(n882) );
  XNOR U1050 ( .A(n882), .B(n881), .Z(n771) );
  XOR U1051 ( .A(n880), .B(n771), .Z(n889) );
  OR U1052 ( .A(n774), .B(n772), .Z(n778) );
  ANDN U1053 ( .B(n774), .A(n773), .Z(n775) );
  OR U1054 ( .A(n776), .B(n775), .Z(n777) );
  AND U1055 ( .A(n778), .B(n777), .Z(n890) );
  XOR U1056 ( .A(n889), .B(n890), .Z(n779) );
  XNOR U1057 ( .A(n891), .B(n779), .Z(n870) );
  XOR U1058 ( .A(n871), .B(n870), .Z(n780) );
  XOR U1059 ( .A(n869), .B(n780), .Z(n933) );
  OR U1060 ( .A(n783), .B(n781), .Z(n787) );
  ANDN U1061 ( .B(n783), .A(n782), .Z(n784) );
  OR U1062 ( .A(n785), .B(n784), .Z(n786) );
  AND U1063 ( .A(n787), .B(n786), .Z(n867) );
  OR U1064 ( .A(n793), .B(n791), .Z(n797) );
  ANDN U1065 ( .B(n793), .A(n792), .Z(n795) );
  NANDN U1066 ( .A(n795), .B(n794), .Z(n796) );
  AND U1067 ( .A(n797), .B(n796), .Z(n920) );
  OR U1068 ( .A(n799), .B(n798), .Z(n803) );
  NANDN U1069 ( .A(n801), .B(n800), .Z(n802) );
  AND U1070 ( .A(n803), .B(n802), .Z(n921) );
  XNOR U1071 ( .A(n906), .B(n905), .Z(n813) );
  XOR U1072 ( .A(n904), .B(n813), .Z(n919) );
  XOR U1073 ( .A(n921), .B(n919), .Z(n814) );
  XOR U1074 ( .A(n920), .B(n814), .Z(n866) );
  XOR U1075 ( .A(n868), .B(n866), .Z(n815) );
  XNOR U1076 ( .A(n867), .B(n815), .Z(n934) );
  NANDN U1077 ( .A(n820), .B(n819), .Z(n825) );
  ANDN U1078 ( .B(n820), .A(n819), .Z(n823) );
  IV U1079 ( .A(n821), .Z(n822) );
  NANDN U1080 ( .A(n823), .B(n822), .Z(n824) );
  AND U1081 ( .A(n825), .B(n824), .Z(n922) );
  XNOR U1082 ( .A(n922), .B(n923), .Z(n829) );
  XOR U1083 ( .A(n924), .B(n829), .Z(n928) );
  NANDN U1084 ( .A(n831), .B(n830), .Z(n835) );
  NANDN U1085 ( .A(n833), .B(n832), .Z(n834) );
  AND U1086 ( .A(n835), .B(n834), .Z(n930) );
  OR U1087 ( .A(n843), .B(n842), .Z(n847) );
  AND U1088 ( .A(n843), .B(n842), .Z(n844) );
  OR U1089 ( .A(n845), .B(n844), .Z(n846) );
  AND U1090 ( .A(n847), .B(n846), .Z(n925) );
  XOR U1091 ( .A(n926), .B(n925), .Z(n848) );
  XNOR U1092 ( .A(n927), .B(n848), .Z(n929) );
  XOR U1093 ( .A(n930), .B(n929), .Z(n849) );
  XOR U1094 ( .A(n928), .B(n849), .Z(n932) );
  XOR U1095 ( .A(n934), .B(n932), .Z(n850) );
  XOR U1096 ( .A(n933), .B(n850), .Z(n858) );
  NANDN U1097 ( .A(n852), .B(n851), .Z(n856) );
  NAND U1098 ( .A(n854), .B(n853), .Z(n855) );
  NAND U1099 ( .A(n856), .B(n855), .Z(n857) );
  XNOR U1100 ( .A(n858), .B(n857), .Z(n859) );
  XNOR U1101 ( .A(n860), .B(n859), .Z(o[2]) );
  NANDN U1102 ( .A(n858), .B(n857), .Z(n862) );
  NAND U1103 ( .A(n860), .B(n859), .Z(n861) );
  AND U1104 ( .A(n862), .B(n861), .Z(n981) );
  XOR U1105 ( .A(n975), .B(n974), .Z(n872) );
  XNOR U1106 ( .A(n973), .B(n872), .Z(n980) );
  XNOR U1107 ( .A(n981), .B(n980), .Z(n983) );
  NANDN U1108 ( .A(n873), .B(n874), .Z(n879) );
  NOR U1109 ( .A(n875), .B(n874), .Z(n877) );
  NANDN U1110 ( .A(n877), .B(n876), .Z(n878) );
  AND U1111 ( .A(n879), .B(n878), .Z(n979) );
  XOR U1112 ( .A(n964), .B(n963), .Z(n965) );
  XOR U1113 ( .A(n966), .B(n965), .Z(n936) );
  IV U1114 ( .A(n936), .Z(n937) );
  NANDN U1115 ( .A(n893), .B(n892), .Z(n897) );
  ANDN U1116 ( .B(n893), .A(n892), .Z(n894) );
  OR U1117 ( .A(n895), .B(n894), .Z(n896) );
  AND U1118 ( .A(n897), .B(n896), .Z(n938) );
  XNOR U1119 ( .A(n940), .B(n938), .Z(n898) );
  XOR U1120 ( .A(n937), .B(n898), .Z(n970) );
  ANDN U1121 ( .B(n900), .A(n899), .Z(n956) );
  XNOR U1122 ( .A(n956), .B(n955), .Z(n958) );
  NANDN U1123 ( .A(n908), .B(n907), .Z(n912) );
  OR U1124 ( .A(n910), .B(n909), .Z(n911) );
  AND U1125 ( .A(n912), .B(n911), .Z(n913) );
  NAND U1126 ( .A(n914), .B(n913), .Z(n1006) );
  IV U1127 ( .A(n1006), .Z(n957) );
  OR U1128 ( .A(n914), .B(n913), .Z(n960) );
  NANDN U1129 ( .A(n957), .B(n960), .Z(n915) );
  XOR U1130 ( .A(n958), .B(n915), .Z(n951) );
  XOR U1131 ( .A(n950), .B(n949), .Z(n952) );
  XOR U1132 ( .A(n951), .B(n952), .Z(n946) );
  XOR U1133 ( .A(n944), .B(n943), .Z(n945) );
  XOR U1134 ( .A(n946), .B(n945), .Z(n972) );
  XNOR U1135 ( .A(n972), .B(n971), .Z(n931) );
  XOR U1136 ( .A(n970), .B(n931), .Z(n978) );
  XNOR U1137 ( .A(n978), .B(n977), .Z(n935) );
  XNOR U1138 ( .A(n979), .B(n935), .Z(n982) );
  XNOR U1139 ( .A(n983), .B(n982), .Z(o[3]) );
  OR U1140 ( .A(n938), .B(n936), .Z(n942) );
  ANDN U1141 ( .B(n938), .A(n937), .Z(n939) );
  OR U1142 ( .A(n940), .B(n939), .Z(n941) );
  AND U1143 ( .A(n942), .B(n941), .Z(n998) );
  OR U1144 ( .A(n944), .B(n943), .Z(n948) );
  NAND U1145 ( .A(n946), .B(n945), .Z(n947) );
  NAND U1146 ( .A(n948), .B(n947), .Z(n996) );
  OR U1147 ( .A(n950), .B(n949), .Z(n954) );
  NAND U1148 ( .A(n952), .B(n951), .Z(n953) );
  AND U1149 ( .A(n954), .B(n953), .Z(n1004) );
  ANDN U1150 ( .B(n956), .A(n955), .Z(n1007) );
  XOR U1151 ( .A(n1006), .B(n1007), .Z(n962) );
  ANDN U1152 ( .B(n958), .A(n957), .Z(n959) );
  NAND U1153 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1154 ( .A(n962), .B(n961), .Z(n1002) );
  OR U1155 ( .A(n964), .B(n963), .Z(n968) );
  NANDN U1156 ( .A(n966), .B(n965), .Z(n967) );
  AND U1157 ( .A(n968), .B(n967), .Z(n1001) );
  XNOR U1158 ( .A(n1002), .B(n1001), .Z(n969) );
  XOR U1159 ( .A(n1004), .B(n969), .Z(n995) );
  XNOR U1160 ( .A(n996), .B(n995), .Z(n997) );
  XNOR U1161 ( .A(n987), .B(n986), .Z(n976) );
  XOR U1162 ( .A(n988), .B(n976), .Z(n992) );
  NANDN U1163 ( .A(n981), .B(n980), .Z(n985) );
  NAND U1164 ( .A(n983), .B(n982), .Z(n984) );
  NAND U1165 ( .A(n985), .B(n984), .Z(n989) );
  XNOR U1166 ( .A(n990), .B(n989), .Z(n991) );
  XNOR U1167 ( .A(n992), .B(n991), .Z(o[4]) );
  NANDN U1168 ( .A(n990), .B(n989), .Z(n994) );
  NAND U1169 ( .A(n992), .B(n991), .Z(n993) );
  NAND U1170 ( .A(n994), .B(n993), .Z(n1016) );
  XNOR U1171 ( .A(n1017), .B(n1016), .Z(n1019) );
  NAND U1172 ( .A(n996), .B(n995), .Z(n1000) );
  OR U1173 ( .A(n998), .B(n997), .Z(n999) );
  NAND U1174 ( .A(n1000), .B(n999), .Z(n1012) );
  NAND U1175 ( .A(n1001), .B(n1002), .Z(n1005) );
  OR U1176 ( .A(n1002), .B(n1001), .Z(n1003) );
  AND U1177 ( .A(n1004), .B(n1003), .Z(n1009) );
  ANDN U1178 ( .B(n1005), .A(n1009), .Z(n1008) );
  ANDN U1179 ( .B(n1007), .A(n1006), .Z(n1010) );
  ANDN U1180 ( .B(n1008), .A(n1010), .Z(n1013) );
  NAND U1181 ( .A(n1010), .B(n1009), .Z(n1015) );
  NANDN U1182 ( .A(n1013), .B(n1015), .Z(n1011) );
  XNOR U1183 ( .A(n1012), .B(n1011), .Z(n1018) );
  XNOR U1184 ( .A(n1019), .B(n1018), .Z(o[5]) );
  OR U1185 ( .A(n1013), .B(n1012), .Z(n1014) );
  AND U1186 ( .A(n1015), .B(n1014), .Z(n1022) );
  NANDN U1187 ( .A(n1017), .B(n1016), .Z(n1021) );
  NAND U1188 ( .A(n1019), .B(n1018), .Z(n1020) );
  AND U1189 ( .A(n1021), .B(n1020), .Z(n1023) );
  XNOR U1190 ( .A(n1022), .B(n1023), .Z(o[6]) );
  ANDN U1191 ( .B(n1023), .A(n1022), .Z(o[7]) );
endmodule

