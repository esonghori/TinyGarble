
module stackMachine_N16 ( clk, rst, x, opcode, o );
  input [15:0] x;
  input [2:0] opcode;
  output [15:0] o;
  input clk, rst;
  wire   \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \stack[0][15] , \stack[0][14] , \stack[0][13] , \stack[0][12] ,
         \stack[0][11] , \stack[0][10] , \stack[0][9] , \stack[0][8] ,
         \stack[0][7] , \stack[0][6] , \stack[0][5] , \stack[0][4] ,
         \stack[0][3] , \stack[0][2] , \stack[0][1] , \stack[0][0] , n1013,
         n1020, n1027, n1036, n1045, n1054, n1063, n1072, n1081, n1090, n1099,
         n1108, n1117, n1126, n1135, n1144, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084;

  DFF \stack_reg[0][0]  ( .D(n1267), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][0] ) );
  DFF \stack_reg[1][0]  ( .D(n1251), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][0] ) );
  DFF \stack_reg[0][15]  ( .D(n1252), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][15] ) );
  DFF \stack_reg[1][15]  ( .D(n1236), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][15] ) );
  DFF \stack_reg[0][1]  ( .D(n1266), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][1] ) );
  DFF \stack_reg[1][1]  ( .D(n1250), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][1] ) );
  DFF \stack_reg[2][1]  ( .D(n1234), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][1] ) );
  DFF \stack_reg[3][1]  ( .D(n1218), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][1] ) );
  DFF \stack_reg[4][1]  ( .D(n1202), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][1] ) );
  DFF \stack_reg[5][1]  ( .D(n1186), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][1] ) );
  DFF \stack_reg[6][1]  ( .D(n1170), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][1] ) );
  DFF \stack_reg[7][1]  ( .D(n1144), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][1] ) );
  DFF \stack_reg[0][2]  ( .D(n1265), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][2] ) );
  DFF \stack_reg[1][2]  ( .D(n1249), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][2] ) );
  DFF \stack_reg[2][2]  ( .D(n1233), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][2] ) );
  DFF \stack_reg[3][2]  ( .D(n1217), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][2] ) );
  DFF \stack_reg[4][2]  ( .D(n1201), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][2] ) );
  DFF \stack_reg[5][2]  ( .D(n1185), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][2] ) );
  DFF \stack_reg[6][2]  ( .D(n1169), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][2] ) );
  DFF \stack_reg[7][2]  ( .D(n1135), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][2] ) );
  DFF \stack_reg[0][3]  ( .D(n1264), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][3] ) );
  DFF \stack_reg[1][3]  ( .D(n1248), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][3] ) );
  DFF \stack_reg[2][3]  ( .D(n1232), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][3] ) );
  DFF \stack_reg[3][3]  ( .D(n1216), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][3] ) );
  DFF \stack_reg[4][3]  ( .D(n1200), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][3] ) );
  DFF \stack_reg[5][3]  ( .D(n1184), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][3] ) );
  DFF \stack_reg[6][3]  ( .D(n1168), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][3] ) );
  DFF \stack_reg[7][3]  ( .D(n1126), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][3] ) );
  DFF \stack_reg[0][4]  ( .D(n1263), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][4] ) );
  DFF \stack_reg[1][4]  ( .D(n1247), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][4] ) );
  DFF \stack_reg[2][4]  ( .D(n1231), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][4] ) );
  DFF \stack_reg[3][4]  ( .D(n1215), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][4] ) );
  DFF \stack_reg[4][4]  ( .D(n1199), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][4] ) );
  DFF \stack_reg[5][4]  ( .D(n1183), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][4] ) );
  DFF \stack_reg[6][4]  ( .D(n1167), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][4] ) );
  DFF \stack_reg[7][4]  ( .D(n1117), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][4] ) );
  DFF \stack_reg[0][5]  ( .D(n1262), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][5] ) );
  DFF \stack_reg[1][5]  ( .D(n1246), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][5] ) );
  DFF \stack_reg[2][5]  ( .D(n1230), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][5] ) );
  DFF \stack_reg[3][5]  ( .D(n1214), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][5] ) );
  DFF \stack_reg[4][5]  ( .D(n1198), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][5] ) );
  DFF \stack_reg[5][5]  ( .D(n1182), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][5] ) );
  DFF \stack_reg[6][5]  ( .D(n1166), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][5] ) );
  DFF \stack_reg[7][5]  ( .D(n1108), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][5] ) );
  DFF \stack_reg[0][6]  ( .D(n1261), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][6] ) );
  DFF \stack_reg[1][6]  ( .D(n1245), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][6] ) );
  DFF \stack_reg[2][6]  ( .D(n1229), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][6] ) );
  DFF \stack_reg[3][6]  ( .D(n1213), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][6] ) );
  DFF \stack_reg[4][6]  ( .D(n1197), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][6] ) );
  DFF \stack_reg[5][6]  ( .D(n1181), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][6] ) );
  DFF \stack_reg[6][6]  ( .D(n1165), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][6] ) );
  DFF \stack_reg[7][6]  ( .D(n1099), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][6] ) );
  DFF \stack_reg[0][7]  ( .D(n1260), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][7] ) );
  DFF \stack_reg[1][7]  ( .D(n1244), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][7] ) );
  DFF \stack_reg[2][7]  ( .D(n1228), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][7] ) );
  DFF \stack_reg[3][7]  ( .D(n1212), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][7] ) );
  DFF \stack_reg[4][7]  ( .D(n1196), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][7] ) );
  DFF \stack_reg[5][7]  ( .D(n1180), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][7] ) );
  DFF \stack_reg[6][7]  ( .D(n1164), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][7] ) );
  DFF \stack_reg[7][7]  ( .D(n1090), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][7] ) );
  DFF \stack_reg[0][8]  ( .D(n1259), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][8] ) );
  DFF \stack_reg[1][8]  ( .D(n1243), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][8] ) );
  DFF \stack_reg[2][8]  ( .D(n1227), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][8] ) );
  DFF \stack_reg[3][8]  ( .D(n1211), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][8] ) );
  DFF \stack_reg[4][8]  ( .D(n1195), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][8] ) );
  DFF \stack_reg[5][8]  ( .D(n1179), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][8] ) );
  DFF \stack_reg[6][8]  ( .D(n1163), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][8] ) );
  DFF \stack_reg[7][8]  ( .D(n1081), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][8] ) );
  DFF \stack_reg[0][9]  ( .D(n1258), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][9] ) );
  DFF \stack_reg[1][9]  ( .D(n1242), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][9] ) );
  DFF \stack_reg[2][9]  ( .D(n1226), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][9] ) );
  DFF \stack_reg[3][9]  ( .D(n1210), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][9] ) );
  DFF \stack_reg[4][9]  ( .D(n1194), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][9] ) );
  DFF \stack_reg[5][9]  ( .D(n1178), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][9] ) );
  DFF \stack_reg[6][9]  ( .D(n1162), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][9] ) );
  DFF \stack_reg[7][9]  ( .D(n1072), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][9] ) );
  DFF \stack_reg[0][10]  ( .D(n1257), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][10] ) );
  DFF \stack_reg[1][10]  ( .D(n1241), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][10] ) );
  DFF \stack_reg[2][10]  ( .D(n1225), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][10] ) );
  DFF \stack_reg[3][10]  ( .D(n1209), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][10] ) );
  DFF \stack_reg[4][10]  ( .D(n1193), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][10] ) );
  DFF \stack_reg[5][10]  ( .D(n1177), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][10] ) );
  DFF \stack_reg[6][10]  ( .D(n1161), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][10] ) );
  DFF \stack_reg[7][10]  ( .D(n1063), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][10] ) );
  DFF \stack_reg[0][11]  ( .D(n1256), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][11] ) );
  DFF \stack_reg[1][11]  ( .D(n1240), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][11] ) );
  DFF \stack_reg[2][11]  ( .D(n1224), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][11] ) );
  DFF \stack_reg[3][11]  ( .D(n1208), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][11] ) );
  DFF \stack_reg[4][11]  ( .D(n1192), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][11] ) );
  DFF \stack_reg[5][11]  ( .D(n1176), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][11] ) );
  DFF \stack_reg[6][11]  ( .D(n1160), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][11] ) );
  DFF \stack_reg[7][11]  ( .D(n1054), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][11] ) );
  DFF \stack_reg[0][12]  ( .D(n1255), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][12] ) );
  DFF \stack_reg[1][12]  ( .D(n1239), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][12] ) );
  DFF \stack_reg[2][12]  ( .D(n1223), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][12] ) );
  DFF \stack_reg[3][12]  ( .D(n1207), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][12] ) );
  DFF \stack_reg[4][12]  ( .D(n1191), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][12] ) );
  DFF \stack_reg[5][12]  ( .D(n1175), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][12] ) );
  DFF \stack_reg[6][12]  ( .D(n1159), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][12] ) );
  DFF \stack_reg[7][12]  ( .D(n1045), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][12] ) );
  DFF \stack_reg[0][13]  ( .D(n1254), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][13] ) );
  DFF \stack_reg[1][13]  ( .D(n1238), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][13] ) );
  DFF \stack_reg[2][13]  ( .D(n1222), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][13] ) );
  DFF \stack_reg[3][13]  ( .D(n1206), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][13] ) );
  DFF \stack_reg[4][13]  ( .D(n1190), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][13] ) );
  DFF \stack_reg[5][13]  ( .D(n1174), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][13] ) );
  DFF \stack_reg[6][13]  ( .D(n1158), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][13] ) );
  DFF \stack_reg[7][13]  ( .D(n1036), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][13] ) );
  DFF \stack_reg[0][14]  ( .D(n1253), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[0][14] ) );
  DFF \stack_reg[1][14]  ( .D(n1237), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[1][14] ) );
  DFF \stack_reg[2][14]  ( .D(n1221), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][14] ) );
  DFF \stack_reg[3][14]  ( .D(n1205), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][14] ) );
  DFF \stack_reg[4][14]  ( .D(n1189), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][14] ) );
  DFF \stack_reg[5][14]  ( .D(n1173), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][14] ) );
  DFF \stack_reg[6][14]  ( .D(n1157), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][14] ) );
  DFF \stack_reg[7][14]  ( .D(n1027), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][14] ) );
  DFF \stack_reg[2][15]  ( .D(n1220), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][15] ) );
  DFF \stack_reg[3][15]  ( .D(n1204), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][15] ) );
  DFF \stack_reg[4][15]  ( .D(n1188), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][15] ) );
  DFF \stack_reg[5][15]  ( .D(n1172), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][15] ) );
  DFF \stack_reg[6][15]  ( .D(n1156), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][15] ) );
  DFF \stack_reg[7][15]  ( .D(n1020), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][15] ) );
  DFF \stack_reg[2][0]  ( .D(n1235), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[2][0] ) );
  DFF \stack_reg[3][0]  ( .D(n1219), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[3][0] ) );
  DFF \stack_reg[4][0]  ( .D(n1203), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[4][0] ) );
  DFF \stack_reg[5][0]  ( .D(n1187), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[5][0] ) );
  DFF \stack_reg[6][0]  ( .D(n1171), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[6][0] ) );
  DFF \stack_reg[7][0]  ( .D(n1013), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        \stack[7][0] ) );
  OR U1280 ( .A(\stack[0][13] ), .B(\stack[1][13] ), .Z(n1641) );
  OR U1281 ( .A(\stack[0][12] ), .B(\stack[1][12] ), .Z(n1618) );
  OR U1282 ( .A(n1704), .B(n1703), .Z(n1706) );
  NANDN U1283 ( .A(\stack[0][2] ), .B(n1380), .Z(n1379) );
  OR U1284 ( .A(n2221), .B(n2223), .Z(n2271) );
  OR U1285 ( .A(n2096), .B(n2098), .Z(n2161) );
  OR U1286 ( .A(n1716), .B(n1715), .Z(n1718) );
  OR U1287 ( .A(n1941), .B(n1943), .Z(n2021) );
  NANDN U1288 ( .A(n1551), .B(n1553), .Z(n2438) );
  XNOR U1289 ( .A(\stack[1][15] ), .B(\stack[0][15] ), .Z(n1687) );
  NANDN U1290 ( .A(\stack[0][1] ), .B(n1357), .Z(n1356) );
  OR U1291 ( .A(n1740), .B(n1739), .Z(n1742) );
  OR U1292 ( .A(n1754), .B(n1753), .Z(n1756) );
  OR U1293 ( .A(n1774), .B(n1773), .Z(n1776) );
  OR U1294 ( .A(n1800), .B(n1799), .Z(n1802) );
  NANDN U1295 ( .A(n1814), .B(n1813), .Z(n1816) );
  NANDN U1296 ( .A(n1539), .B(n1541), .Z(n1836) );
  NANDN U1297 ( .A(n1339), .B(n1341), .Z(n2473) );
  OR U1298 ( .A(\stack[0][15] ), .B(\stack[1][15] ), .Z(n2398) );
  NANDN U1299 ( .A(n1268), .B(n1269), .Z(o[9]) );
  NANDN U1300 ( .A(n1270), .B(n1271), .Z(n1269) );
  NANDN U1301 ( .A(n1272), .B(n1273), .Z(o[8]) );
  NANDN U1302 ( .A(n1274), .B(n1271), .Z(n1273) );
  NANDN U1303 ( .A(n1275), .B(n1276), .Z(o[7]) );
  NANDN U1304 ( .A(n1277), .B(n1271), .Z(n1276) );
  NANDN U1305 ( .A(n1278), .B(n1279), .Z(o[6]) );
  NANDN U1306 ( .A(n1280), .B(n1271), .Z(n1279) );
  NANDN U1307 ( .A(n1281), .B(n1282), .Z(o[5]) );
  NANDN U1308 ( .A(n1283), .B(n1271), .Z(n1282) );
  NANDN U1309 ( .A(n1284), .B(n1285), .Z(o[4]) );
  NANDN U1310 ( .A(n1286), .B(n1271), .Z(n1285) );
  NANDN U1311 ( .A(n1287), .B(n1288), .Z(o[3]) );
  NANDN U1312 ( .A(n1289), .B(n1271), .Z(n1288) );
  NANDN U1313 ( .A(n1290), .B(n1291), .Z(o[2]) );
  NANDN U1314 ( .A(n1292), .B(n1271), .Z(n1291) );
  NANDN U1315 ( .A(n1293), .B(n1294), .Z(o[1]) );
  NANDN U1316 ( .A(n1295), .B(n1271), .Z(n1294) );
  NANDN U1317 ( .A(n1296), .B(n1297), .Z(o[15]) );
  NANDN U1318 ( .A(n1298), .B(n1271), .Z(n1297) );
  NANDN U1319 ( .A(n1299), .B(n1300), .Z(o[14]) );
  NANDN U1320 ( .A(n1301), .B(n1271), .Z(n1300) );
  NANDN U1321 ( .A(n1302), .B(n1303), .Z(o[13]) );
  NANDN U1322 ( .A(n1304), .B(n1271), .Z(n1303) );
  NANDN U1323 ( .A(n1305), .B(n1306), .Z(o[12]) );
  NANDN U1324 ( .A(n1307), .B(n1271), .Z(n1306) );
  NANDN U1325 ( .A(n1308), .B(n1309), .Z(o[11]) );
  NANDN U1326 ( .A(n1310), .B(n1271), .Z(n1309) );
  NANDN U1327 ( .A(n1311), .B(n1312), .Z(o[10]) );
  NANDN U1328 ( .A(n1313), .B(n1271), .Z(n1312) );
  NANDN U1329 ( .A(n1314), .B(n1315), .Z(o[0]) );
  NANDN U1330 ( .A(n1316), .B(n1271), .Z(n1315) );
  NAND U1331 ( .A(n1317), .B(n1318), .Z(n1267) );
  NANDN U1332 ( .A(n1319), .B(\stack[0][0] ), .Z(n1318) );
  ANDN U1333 ( .B(n1320), .A(n1314), .Z(n1317) );
  ANDN U1334 ( .B(x[0]), .A(n1271), .Z(n1314) );
  NANDN U1335 ( .A(n1316), .B(n1321), .Z(n1320) );
  AND U1336 ( .A(n1322), .B(n1323), .Z(n1316) );
  AND U1337 ( .A(n1324), .B(n1325), .Z(n1323) );
  NAND U1338 ( .A(n1326), .B(n1327), .Z(n1325) );
  AND U1339 ( .A(\stack[0][0] ), .B(\stack[1][0] ), .Z(n1326) );
  AND U1340 ( .A(n1328), .B(n1329), .Z(n1324) );
  NAND U1341 ( .A(\stack[1][0] ), .B(n1330), .Z(n1329) );
  ANDN U1342 ( .B(\stack[0][0] ), .A(n1331), .Z(n1330) );
  NAND U1343 ( .A(n1332), .B(n1333), .Z(n1328) );
  NAND U1344 ( .A(n1334), .B(n1335), .Z(n1332) );
  AND U1345 ( .A(n1336), .B(n1337), .Z(n1322) );
  NAND U1346 ( .A(\stack[0][0] ), .B(n1338), .Z(n1337) );
  XOR U1347 ( .A(n1339), .B(n1340), .Z(n1336) );
  XNOR U1348 ( .A(n1341), .B(n1342), .Z(n1340) );
  NAND U1349 ( .A(n1343), .B(n1344), .Z(n1266) );
  NANDN U1350 ( .A(n1319), .B(\stack[0][1] ), .Z(n1344) );
  ANDN U1351 ( .B(n1345), .A(n1293), .Z(n1343) );
  ANDN U1352 ( .B(x[1]), .A(n1271), .Z(n1293) );
  NANDN U1353 ( .A(n1295), .B(n1321), .Z(n1345) );
  AND U1354 ( .A(n1346), .B(n1347), .Z(n1295) );
  AND U1355 ( .A(n1348), .B(n1349), .Z(n1347) );
  NAND U1356 ( .A(n1350), .B(n1327), .Z(n1349) );
  XOR U1357 ( .A(n1351), .B(n1352), .Z(n1350) );
  AND U1358 ( .A(n1353), .B(n1354), .Z(n1348) );
  NAND U1359 ( .A(\stack[1][1] ), .B(n1355), .Z(n1354) );
  ANDN U1360 ( .B(\stack[0][1] ), .A(n1331), .Z(n1355) );
  NAND U1361 ( .A(n1356), .B(n1333), .Z(n1353) );
  AND U1362 ( .A(n1358), .B(n1359), .Z(n1346) );
  NAND U1363 ( .A(\stack[0][1] ), .B(n1338), .Z(n1359) );
  XNOR U1364 ( .A(n1360), .B(n1361), .Z(n1358) );
  XNOR U1365 ( .A(n1362), .B(n1363), .Z(n1361) );
  NAND U1366 ( .A(n1364), .B(n1365), .Z(n1265) );
  NANDN U1367 ( .A(n1319), .B(\stack[0][2] ), .Z(n1365) );
  ANDN U1368 ( .B(n1366), .A(n1290), .Z(n1364) );
  ANDN U1369 ( .B(x[2]), .A(n1271), .Z(n1290) );
  NANDN U1370 ( .A(n1292), .B(n1321), .Z(n1366) );
  AND U1371 ( .A(n1367), .B(n1368), .Z(n1292) );
  AND U1372 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1373 ( .A(n1371), .B(n1327), .Z(n1370) );
  XNOR U1374 ( .A(n1372), .B(n1373), .Z(n1371) );
  XNOR U1375 ( .A(n1374), .B(n1375), .Z(n1373) );
  AND U1376 ( .A(n1376), .B(n1377), .Z(n1369) );
  NAND U1377 ( .A(\stack[1][2] ), .B(n1378), .Z(n1377) );
  ANDN U1378 ( .B(\stack[0][2] ), .A(n1331), .Z(n1378) );
  NAND U1379 ( .A(n1379), .B(n1333), .Z(n1376) );
  AND U1380 ( .A(n1381), .B(n1382), .Z(n1367) );
  NAND U1381 ( .A(\stack[0][2] ), .B(n1338), .Z(n1382) );
  XNOR U1382 ( .A(n1383), .B(n1384), .Z(n1381) );
  XNOR U1383 ( .A(n1385), .B(n1386), .Z(n1384) );
  NAND U1384 ( .A(n1387), .B(n1388), .Z(n1264) );
  NANDN U1385 ( .A(n1319), .B(\stack[0][3] ), .Z(n1388) );
  ANDN U1386 ( .B(n1389), .A(n1287), .Z(n1387) );
  ANDN U1387 ( .B(x[3]), .A(n1271), .Z(n1287) );
  NANDN U1388 ( .A(n1289), .B(n1321), .Z(n1389) );
  AND U1389 ( .A(n1390), .B(n1391), .Z(n1289) );
  AND U1390 ( .A(n1392), .B(n1393), .Z(n1391) );
  NAND U1391 ( .A(n1394), .B(n1327), .Z(n1393) );
  XNOR U1392 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U1393 ( .A(n1397), .B(n1398), .Z(n1396) );
  AND U1394 ( .A(n1399), .B(n1400), .Z(n1392) );
  NAND U1395 ( .A(\stack[1][3] ), .B(n1401), .Z(n1400) );
  ANDN U1396 ( .B(\stack[0][3] ), .A(n1331), .Z(n1401) );
  NAND U1397 ( .A(n1402), .B(n1333), .Z(n1399) );
  NAND U1398 ( .A(n1403), .B(n1404), .Z(n1402) );
  AND U1399 ( .A(n1405), .B(n1406), .Z(n1390) );
  NAND U1400 ( .A(\stack[0][3] ), .B(n1338), .Z(n1406) );
  XNOR U1401 ( .A(n1407), .B(n1408), .Z(n1405) );
  XNOR U1402 ( .A(n1409), .B(n1410), .Z(n1408) );
  NAND U1403 ( .A(n1411), .B(n1412), .Z(n1263) );
  NANDN U1404 ( .A(n1319), .B(\stack[0][4] ), .Z(n1412) );
  ANDN U1405 ( .B(n1413), .A(n1284), .Z(n1411) );
  ANDN U1406 ( .B(x[4]), .A(n1271), .Z(n1284) );
  NANDN U1407 ( .A(n1286), .B(n1321), .Z(n1413) );
  AND U1408 ( .A(n1414), .B(n1415), .Z(n1286) );
  AND U1409 ( .A(n1416), .B(n1417), .Z(n1415) );
  NAND U1410 ( .A(n1418), .B(n1327), .Z(n1417) );
  XOR U1411 ( .A(n1419), .B(n1420), .Z(n1418) );
  XNOR U1412 ( .A(n1421), .B(n1422), .Z(n1420) );
  AND U1413 ( .A(n1423), .B(n1424), .Z(n1416) );
  NAND U1414 ( .A(\stack[1][4] ), .B(n1425), .Z(n1424) );
  ANDN U1415 ( .B(\stack[0][4] ), .A(n1331), .Z(n1425) );
  NAND U1416 ( .A(n1426), .B(n1333), .Z(n1423) );
  NAND U1417 ( .A(n1427), .B(n1428), .Z(n1426) );
  AND U1418 ( .A(n1429), .B(n1430), .Z(n1414) );
  NAND U1419 ( .A(\stack[0][4] ), .B(n1338), .Z(n1430) );
  XNOR U1420 ( .A(n1431), .B(n1432), .Z(n1429) );
  XNOR U1421 ( .A(n1433), .B(n1434), .Z(n1432) );
  NAND U1422 ( .A(n1435), .B(n1436), .Z(n1262) );
  NANDN U1423 ( .A(n1319), .B(\stack[0][5] ), .Z(n1436) );
  ANDN U1424 ( .B(n1437), .A(n1281), .Z(n1435) );
  ANDN U1425 ( .B(x[5]), .A(n1271), .Z(n1281) );
  NANDN U1426 ( .A(n1283), .B(n1321), .Z(n1437) );
  AND U1427 ( .A(n1438), .B(n1439), .Z(n1283) );
  AND U1428 ( .A(n1440), .B(n1441), .Z(n1439) );
  NAND U1429 ( .A(n1442), .B(n1327), .Z(n1441) );
  XNOR U1430 ( .A(n1443), .B(n1444), .Z(n1442) );
  XOR U1431 ( .A(n1445), .B(n1446), .Z(n1444) );
  AND U1432 ( .A(n1447), .B(n1448), .Z(n1440) );
  NAND U1433 ( .A(\stack[0][5] ), .B(n1449), .Z(n1448) );
  ANDN U1434 ( .B(\stack[1][5] ), .A(n1331), .Z(n1449) );
  NAND U1435 ( .A(n1450), .B(n1333), .Z(n1447) );
  NAND U1436 ( .A(n1451), .B(n1452), .Z(n1450) );
  AND U1437 ( .A(n1453), .B(n1454), .Z(n1438) );
  NAND U1438 ( .A(\stack[0][5] ), .B(n1338), .Z(n1454) );
  XNOR U1439 ( .A(n1455), .B(n1456), .Z(n1453) );
  XNOR U1440 ( .A(n1457), .B(n1458), .Z(n1456) );
  NAND U1441 ( .A(n1459), .B(n1460), .Z(n1261) );
  NANDN U1442 ( .A(n1319), .B(\stack[0][6] ), .Z(n1460) );
  ANDN U1443 ( .B(n1461), .A(n1278), .Z(n1459) );
  ANDN U1444 ( .B(x[6]), .A(n1271), .Z(n1278) );
  NANDN U1445 ( .A(n1280), .B(n1321), .Z(n1461) );
  AND U1446 ( .A(n1462), .B(n1463), .Z(n1280) );
  AND U1447 ( .A(n1464), .B(n1465), .Z(n1463) );
  NAND U1448 ( .A(n1466), .B(n1327), .Z(n1465) );
  XOR U1449 ( .A(n1467), .B(n1468), .Z(n1466) );
  XNOR U1450 ( .A(n1469), .B(n1470), .Z(n1468) );
  AND U1451 ( .A(n1471), .B(n1472), .Z(n1464) );
  NAND U1452 ( .A(\stack[0][6] ), .B(n1473), .Z(n1472) );
  ANDN U1453 ( .B(\stack[1][6] ), .A(n1331), .Z(n1473) );
  NAND U1454 ( .A(n1474), .B(n1333), .Z(n1471) );
  NAND U1455 ( .A(n1475), .B(n1476), .Z(n1474) );
  AND U1456 ( .A(n1477), .B(n1478), .Z(n1462) );
  NAND U1457 ( .A(\stack[0][6] ), .B(n1338), .Z(n1478) );
  XNOR U1458 ( .A(n1479), .B(n1480), .Z(n1477) );
  XNOR U1459 ( .A(n1481), .B(n1482), .Z(n1480) );
  NAND U1460 ( .A(n1483), .B(n1484), .Z(n1260) );
  NANDN U1461 ( .A(n1319), .B(\stack[0][7] ), .Z(n1484) );
  ANDN U1462 ( .B(n1485), .A(n1275), .Z(n1483) );
  ANDN U1463 ( .B(x[7]), .A(n1271), .Z(n1275) );
  NANDN U1464 ( .A(n1277), .B(n1321), .Z(n1485) );
  AND U1465 ( .A(n1486), .B(n1487), .Z(n1277) );
  AND U1466 ( .A(n1488), .B(n1489), .Z(n1487) );
  NAND U1467 ( .A(n1490), .B(n1327), .Z(n1489) );
  XNOR U1468 ( .A(n1491), .B(n1492), .Z(n1490) );
  XOR U1469 ( .A(n1493), .B(n1494), .Z(n1492) );
  AND U1470 ( .A(n1495), .B(n1496), .Z(n1488) );
  NAND U1471 ( .A(\stack[0][7] ), .B(n1497), .Z(n1496) );
  ANDN U1472 ( .B(\stack[1][7] ), .A(n1331), .Z(n1497) );
  NAND U1473 ( .A(n1498), .B(n1333), .Z(n1495) );
  NAND U1474 ( .A(n1499), .B(n1500), .Z(n1498) );
  AND U1475 ( .A(n1501), .B(n1502), .Z(n1486) );
  NAND U1476 ( .A(\stack[0][7] ), .B(n1338), .Z(n1502) );
  XNOR U1477 ( .A(n1503), .B(n1504), .Z(n1501) );
  XNOR U1478 ( .A(n1505), .B(n1506), .Z(n1504) );
  NAND U1479 ( .A(n1507), .B(n1508), .Z(n1259) );
  NANDN U1480 ( .A(n1319), .B(\stack[0][8] ), .Z(n1508) );
  ANDN U1481 ( .B(n1509), .A(n1272), .Z(n1507) );
  ANDN U1482 ( .B(x[8]), .A(n1271), .Z(n1272) );
  NANDN U1483 ( .A(n1274), .B(n1321), .Z(n1509) );
  AND U1484 ( .A(n1510), .B(n1511), .Z(n1274) );
  AND U1485 ( .A(n1512), .B(n1513), .Z(n1511) );
  NAND U1486 ( .A(n1514), .B(n1327), .Z(n1513) );
  XOR U1487 ( .A(n1515), .B(n1516), .Z(n1514) );
  XNOR U1488 ( .A(n1517), .B(n1518), .Z(n1516) );
  AND U1489 ( .A(n1519), .B(n1520), .Z(n1512) );
  NAND U1490 ( .A(\stack[0][8] ), .B(n1521), .Z(n1520) );
  ANDN U1491 ( .B(\stack[1][8] ), .A(n1331), .Z(n1521) );
  NAND U1492 ( .A(n1522), .B(n1333), .Z(n1519) );
  NAND U1493 ( .A(n1523), .B(n1524), .Z(n1522) );
  AND U1494 ( .A(n1525), .B(n1526), .Z(n1510) );
  NAND U1495 ( .A(\stack[0][8] ), .B(n1338), .Z(n1526) );
  XNOR U1496 ( .A(n1527), .B(n1528), .Z(n1525) );
  XNOR U1497 ( .A(n1529), .B(n1530), .Z(n1528) );
  NAND U1498 ( .A(n1531), .B(n1532), .Z(n1258) );
  NANDN U1499 ( .A(n1319), .B(\stack[0][9] ), .Z(n1532) );
  ANDN U1500 ( .B(n1533), .A(n1268), .Z(n1531) );
  ANDN U1501 ( .B(x[9]), .A(n1271), .Z(n1268) );
  NANDN U1502 ( .A(n1270), .B(n1321), .Z(n1533) );
  AND U1503 ( .A(n1534), .B(n1535), .Z(n1270) );
  AND U1504 ( .A(n1536), .B(n1537), .Z(n1535) );
  NAND U1505 ( .A(n1538), .B(n1327), .Z(n1537) );
  XOR U1506 ( .A(n1539), .B(n1540), .Z(n1538) );
  XNOR U1507 ( .A(n1541), .B(n1542), .Z(n1540) );
  AND U1508 ( .A(n1543), .B(n1544), .Z(n1536) );
  NAND U1509 ( .A(\stack[1][9] ), .B(n1545), .Z(n1544) );
  ANDN U1510 ( .B(\stack[0][9] ), .A(n1331), .Z(n1545) );
  NAND U1511 ( .A(n1546), .B(n1333), .Z(n1543) );
  NAND U1512 ( .A(n1547), .B(n1548), .Z(n1546) );
  AND U1513 ( .A(n1549), .B(n1550), .Z(n1534) );
  NAND U1514 ( .A(\stack[0][9] ), .B(n1338), .Z(n1550) );
  XOR U1515 ( .A(n1551), .B(n1552), .Z(n1549) );
  XNOR U1516 ( .A(n1553), .B(n1554), .Z(n1552) );
  NAND U1517 ( .A(n1555), .B(n1556), .Z(n1257) );
  NANDN U1518 ( .A(n1319), .B(\stack[0][10] ), .Z(n1556) );
  ANDN U1519 ( .B(n1557), .A(n1311), .Z(n1555) );
  ANDN U1520 ( .B(x[10]), .A(n1271), .Z(n1311) );
  NANDN U1521 ( .A(n1313), .B(n1321), .Z(n1557) );
  AND U1522 ( .A(n1558), .B(n1559), .Z(n1313) );
  AND U1523 ( .A(n1560), .B(n1561), .Z(n1559) );
  NAND U1524 ( .A(n1562), .B(n1327), .Z(n1561) );
  XOR U1525 ( .A(n1563), .B(n1564), .Z(n1562) );
  XNOR U1526 ( .A(n1565), .B(n1566), .Z(n1564) );
  AND U1527 ( .A(n1567), .B(n1568), .Z(n1560) );
  NAND U1528 ( .A(\stack[0][10] ), .B(n1569), .Z(n1568) );
  ANDN U1529 ( .B(\stack[1][10] ), .A(n1331), .Z(n1569) );
  NAND U1530 ( .A(n1570), .B(n1333), .Z(n1567) );
  NAND U1531 ( .A(n1571), .B(n1572), .Z(n1570) );
  AND U1532 ( .A(n1573), .B(n1574), .Z(n1558) );
  NAND U1533 ( .A(\stack[0][10] ), .B(n1338), .Z(n1574) );
  XNOR U1534 ( .A(n1575), .B(n1576), .Z(n1573) );
  XNOR U1535 ( .A(n1577), .B(n1578), .Z(n1576) );
  NAND U1536 ( .A(n1579), .B(n1580), .Z(n1256) );
  NANDN U1537 ( .A(n1319), .B(\stack[0][11] ), .Z(n1580) );
  ANDN U1538 ( .B(n1581), .A(n1308), .Z(n1579) );
  ANDN U1539 ( .B(x[11]), .A(n1271), .Z(n1308) );
  NANDN U1540 ( .A(n1310), .B(n1321), .Z(n1581) );
  AND U1541 ( .A(n1582), .B(n1583), .Z(n1310) );
  AND U1542 ( .A(n1584), .B(n1585), .Z(n1583) );
  NAND U1543 ( .A(n1586), .B(n1327), .Z(n1585) );
  XNOR U1544 ( .A(n1587), .B(n1588), .Z(n1586) );
  XOR U1545 ( .A(n1589), .B(n1590), .Z(n1588) );
  AND U1546 ( .A(n1591), .B(n1592), .Z(n1584) );
  NAND U1547 ( .A(\stack[0][11] ), .B(n1593), .Z(n1592) );
  ANDN U1548 ( .B(\stack[1][11] ), .A(n1331), .Z(n1593) );
  NAND U1549 ( .A(n1594), .B(n1333), .Z(n1591) );
  NAND U1550 ( .A(n1595), .B(n1596), .Z(n1594) );
  AND U1551 ( .A(n1597), .B(n1598), .Z(n1582) );
  NAND U1552 ( .A(\stack[0][11] ), .B(n1338), .Z(n1598) );
  XNOR U1553 ( .A(n1599), .B(n1600), .Z(n1597) );
  XNOR U1554 ( .A(n1601), .B(n1602), .Z(n1600) );
  NAND U1555 ( .A(n1603), .B(n1604), .Z(n1255) );
  NANDN U1556 ( .A(n1319), .B(\stack[0][12] ), .Z(n1604) );
  ANDN U1557 ( .B(n1605), .A(n1305), .Z(n1603) );
  ANDN U1558 ( .B(x[12]), .A(n1271), .Z(n1305) );
  NANDN U1559 ( .A(n1307), .B(n1321), .Z(n1605) );
  AND U1560 ( .A(n1606), .B(n1607), .Z(n1307) );
  AND U1561 ( .A(n1608), .B(n1609), .Z(n1607) );
  NAND U1562 ( .A(n1610), .B(n1327), .Z(n1609) );
  XOR U1563 ( .A(n1611), .B(n1612), .Z(n1610) );
  XNOR U1564 ( .A(n1613), .B(n1614), .Z(n1612) );
  AND U1565 ( .A(n1615), .B(n1616), .Z(n1608) );
  NAND U1566 ( .A(\stack[1][12] ), .B(n1617), .Z(n1616) );
  ANDN U1567 ( .B(\stack[0][12] ), .A(n1331), .Z(n1617) );
  NAND U1568 ( .A(n1618), .B(n1333), .Z(n1615) );
  AND U1569 ( .A(n1620), .B(n1621), .Z(n1606) );
  NAND U1570 ( .A(\stack[0][12] ), .B(n1338), .Z(n1621) );
  XNOR U1571 ( .A(n1622), .B(n1623), .Z(n1620) );
  XNOR U1572 ( .A(n1624), .B(n1625), .Z(n1623) );
  NAND U1573 ( .A(n1626), .B(n1627), .Z(n1254) );
  NANDN U1574 ( .A(n1319), .B(\stack[0][13] ), .Z(n1627) );
  ANDN U1575 ( .B(n1628), .A(n1302), .Z(n1626) );
  ANDN U1576 ( .B(x[13]), .A(n1271), .Z(n1302) );
  NANDN U1577 ( .A(n1304), .B(n1321), .Z(n1628) );
  AND U1578 ( .A(n1629), .B(n1630), .Z(n1304) );
  AND U1579 ( .A(n1631), .B(n1632), .Z(n1630) );
  NAND U1580 ( .A(n1633), .B(n1327), .Z(n1632) );
  XOR U1581 ( .A(n1634), .B(n1635), .Z(n1633) );
  XNOR U1582 ( .A(n1636), .B(n1637), .Z(n1635) );
  AND U1583 ( .A(n1638), .B(n1639), .Z(n1631) );
  NAND U1584 ( .A(\stack[0][13] ), .B(n1640), .Z(n1639) );
  ANDN U1585 ( .B(\stack[1][13] ), .A(n1331), .Z(n1640) );
  NAND U1586 ( .A(n1641), .B(n1333), .Z(n1638) );
  AND U1587 ( .A(n1643), .B(n1644), .Z(n1629) );
  NAND U1588 ( .A(\stack[0][13] ), .B(n1338), .Z(n1644) );
  XNOR U1589 ( .A(n1645), .B(n1646), .Z(n1643) );
  XNOR U1590 ( .A(n1647), .B(n1648), .Z(n1646) );
  NAND U1591 ( .A(n1649), .B(n1650), .Z(n1253) );
  NANDN U1592 ( .A(n1319), .B(\stack[0][14] ), .Z(n1650) );
  ANDN U1593 ( .B(n1651), .A(n1299), .Z(n1649) );
  ANDN U1594 ( .B(x[14]), .A(n1271), .Z(n1299) );
  NANDN U1595 ( .A(n1301), .B(n1321), .Z(n1651) );
  AND U1596 ( .A(n1652), .B(n1653), .Z(n1301) );
  AND U1597 ( .A(n1654), .B(n1655), .Z(n1653) );
  NAND U1598 ( .A(n1656), .B(n1327), .Z(n1655) );
  XOR U1599 ( .A(n1657), .B(n1658), .Z(n1656) );
  XNOR U1600 ( .A(n1659), .B(n1660), .Z(n1658) );
  AND U1601 ( .A(n1661), .B(n1662), .Z(n1654) );
  NAND U1602 ( .A(\stack[0][14] ), .B(n1663), .Z(n1662) );
  ANDN U1603 ( .B(\stack[1][14] ), .A(n1331), .Z(n1663) );
  NAND U1604 ( .A(n1664), .B(n1333), .Z(n1661) );
  NAND U1605 ( .A(n1665), .B(n1666), .Z(n1664) );
  IV U1606 ( .A(\stack[1][14] ), .Z(n1666) );
  AND U1607 ( .A(n1667), .B(n1668), .Z(n1652) );
  NAND U1608 ( .A(\stack[0][14] ), .B(n1338), .Z(n1668) );
  XOR U1609 ( .A(n1669), .B(n1670), .Z(n1667) );
  XOR U1610 ( .A(n1671), .B(n1672), .Z(n1670) );
  NAND U1611 ( .A(n1673), .B(n1674), .Z(n1252) );
  NANDN U1612 ( .A(n1319), .B(\stack[0][15] ), .Z(n1674) );
  NANDN U1613 ( .A(n1675), .B(n1676), .Z(n1319) );
  ANDN U1614 ( .B(n1271), .A(n1677), .Z(n1676) );
  ANDN U1615 ( .B(n1678), .A(n1296), .Z(n1673) );
  ANDN U1616 ( .B(x[15]), .A(n1271), .Z(n1296) );
  NANDN U1617 ( .A(n1298), .B(n1321), .Z(n1678) );
  OR U1618 ( .A(n1677), .B(n1675), .Z(n1321) );
  AND U1619 ( .A(n1679), .B(n1680), .Z(n1298) );
  AND U1620 ( .A(n1681), .B(n1682), .Z(n1680) );
  NAND U1621 ( .A(n1683), .B(n1327), .Z(n1682) );
  AND U1622 ( .A(n1684), .B(n1685), .Z(n1683) );
  NANDN U1623 ( .A(n1686), .B(n1687), .Z(n1685) );
  NAND U1624 ( .A(n1688), .B(n1686), .Z(n1684) );
  XOR U1625 ( .A(n1689), .B(n1690), .Z(n1686) );
  XOR U1626 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U1627 ( .A(n1693), .B(n1694), .Z(n1692) );
  XOR U1628 ( .A(n1695), .B(n1696), .Z(n1694) );
  XOR U1629 ( .A(n1697), .B(n1698), .Z(n1696) );
  XOR U1630 ( .A(n1699), .B(n1700), .Z(n1698) );
  NAND U1631 ( .A(n1701), .B(n1702), .Z(n1700) );
  NAND U1632 ( .A(n1703), .B(n1704), .Z(n1702) );
  NANDN U1633 ( .A(n1705), .B(n1706), .Z(n1701) );
  AND U1634 ( .A(\stack[1][1] ), .B(\stack[0][14] ), .Z(n1699) );
  XOR U1635 ( .A(n1707), .B(n1708), .Z(n1697) );
  XOR U1636 ( .A(n1709), .B(n1710), .Z(n1708) );
  XOR U1637 ( .A(n1711), .B(n1712), .Z(n1710) );
  AND U1638 ( .A(n1713), .B(n1714), .Z(n1712) );
  NAND U1639 ( .A(n1715), .B(n1716), .Z(n1714) );
  NANDN U1640 ( .A(n1717), .B(n1718), .Z(n1713) );
  AND U1641 ( .A(\stack[1][3] ), .B(\stack[0][12] ), .Z(n1711) );
  XOR U1642 ( .A(n1719), .B(n1720), .Z(n1709) );
  XOR U1643 ( .A(n1721), .B(n1722), .Z(n1720) );
  XOR U1644 ( .A(n1723), .B(n1724), .Z(n1722) );
  XOR U1645 ( .A(n1725), .B(n1726), .Z(n1724) );
  XOR U1646 ( .A(n1727), .B(n1728), .Z(n1726) );
  AND U1647 ( .A(\stack[0][2] ), .B(\stack[1][13] ), .Z(n1728) );
  ANDN U1648 ( .B(n1729), .A(n1730), .Z(n1727) );
  AND U1649 ( .A(\stack[0][0] ), .B(\stack[1][14] ), .Z(n1729) );
  XOR U1650 ( .A(n1731), .B(n1732), .Z(n1725) );
  AND U1651 ( .A(n1334), .B(\stack[1][15] ), .Z(n1732) );
  IV U1652 ( .A(\stack[0][0] ), .Z(n1334) );
  AND U1653 ( .A(\stack[0][1] ), .B(\stack[1][14] ), .Z(n1731) );
  XOR U1654 ( .A(n1733), .B(n1734), .Z(n1723) );
  XOR U1655 ( .A(n1735), .B(n1736), .Z(n1734) );
  AND U1656 ( .A(n1737), .B(n1738), .Z(n1736) );
  NAND U1657 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1658 ( .A(n1741), .B(n1742), .Z(n1737) );
  AND U1659 ( .A(\stack[0][4] ), .B(\stack[1][11] ), .Z(n1735) );
  XOR U1660 ( .A(n1743), .B(n1744), .Z(n1733) );
  AND U1661 ( .A(n1745), .B(n1746), .Z(n1744) );
  NAND U1662 ( .A(n1747), .B(n1748), .Z(n1746) );
  NANDN U1663 ( .A(n1749), .B(n1750), .Z(n1745) );
  OR U1664 ( .A(n1747), .B(n1748), .Z(n1750) );
  AND U1665 ( .A(\stack[0][3] ), .B(\stack[1][12] ), .Z(n1743) );
  AND U1666 ( .A(n1751), .B(n1752), .Z(n1721) );
  NAND U1667 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1668 ( .A(n1755), .B(n1756), .Z(n1751) );
  XOR U1669 ( .A(n1757), .B(n1758), .Z(n1719) );
  XOR U1670 ( .A(n1759), .B(n1760), .Z(n1758) );
  AND U1671 ( .A(n1761), .B(n1762), .Z(n1760) );
  NANDN U1672 ( .A(n1763), .B(n1764), .Z(n1762) );
  NANDN U1673 ( .A(n1765), .B(n1766), .Z(n1761) );
  NANDN U1674 ( .A(n1764), .B(n1763), .Z(n1766) );
  AND U1675 ( .A(\stack[1][8] ), .B(\stack[0][7] ), .Z(n1759) );
  AND U1676 ( .A(\stack[1][7] ), .B(\stack[0][8] ), .Z(n1757) );
  XOR U1677 ( .A(n1767), .B(n1768), .Z(n1707) );
  XOR U1678 ( .A(n1769), .B(n1770), .Z(n1768) );
  AND U1679 ( .A(n1771), .B(n1772), .Z(n1770) );
  NAND U1680 ( .A(n1773), .B(n1774), .Z(n1772) );
  NANDN U1681 ( .A(n1775), .B(n1776), .Z(n1771) );
  AND U1682 ( .A(\stack[1][9] ), .B(\stack[0][6] ), .Z(n1769) );
  XOR U1683 ( .A(n1777), .B(n1778), .Z(n1767) );
  AND U1684 ( .A(n1779), .B(n1780), .Z(n1778) );
  NANDN U1685 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1686 ( .A(n1783), .B(n1784), .Z(n1779) );
  NANDN U1687 ( .A(n1782), .B(n1781), .Z(n1784) );
  AND U1688 ( .A(\stack[0][5] ), .B(\stack[1][10] ), .Z(n1777) );
  XOR U1689 ( .A(n1785), .B(n1786), .Z(n1695) );
  AND U1690 ( .A(n1787), .B(n1788), .Z(n1786) );
  NANDN U1691 ( .A(n1789), .B(n1790), .Z(n1788) );
  NANDN U1692 ( .A(n1791), .B(n1792), .Z(n1787) );
  NANDN U1693 ( .A(n1790), .B(n1789), .Z(n1792) );
  AND U1694 ( .A(\stack[1][4] ), .B(\stack[0][11] ), .Z(n1785) );
  XOR U1695 ( .A(n1793), .B(n1794), .Z(n1693) );
  XOR U1696 ( .A(n1795), .B(n1796), .Z(n1794) );
  AND U1697 ( .A(n1797), .B(n1798), .Z(n1796) );
  NAND U1698 ( .A(n1799), .B(n1800), .Z(n1798) );
  NANDN U1699 ( .A(n1801), .B(n1802), .Z(n1797) );
  AND U1700 ( .A(\stack[1][5] ), .B(\stack[0][10] ), .Z(n1795) );
  XOR U1701 ( .A(n1803), .B(n1804), .Z(n1793) );
  AND U1702 ( .A(n1805), .B(n1806), .Z(n1804) );
  NANDN U1703 ( .A(n1807), .B(n1808), .Z(n1806) );
  NANDN U1704 ( .A(n1809), .B(n1810), .Z(n1805) );
  NANDN U1705 ( .A(n1808), .B(n1807), .Z(n1810) );
  AND U1706 ( .A(\stack[0][9] ), .B(\stack[1][6] ), .Z(n1803) );
  AND U1707 ( .A(n1811), .B(n1812), .Z(n1691) );
  NANDN U1708 ( .A(n1813), .B(n1814), .Z(n1812) );
  NANDN U1709 ( .A(n1815), .B(n1816), .Z(n1811) );
  XOR U1710 ( .A(n1817), .B(n1818), .Z(n1689) );
  AND U1711 ( .A(\stack[1][2] ), .B(\stack[0][13] ), .Z(n1818) );
  AND U1712 ( .A(n1819), .B(n1820), .Z(n1817) );
  NAND U1713 ( .A(n1821), .B(n1660), .Z(n1820) );
  NAND U1714 ( .A(n1822), .B(n1823), .Z(n1660) );
  NANDN U1715 ( .A(n1637), .B(n1824), .Z(n1823) );
  OR U1716 ( .A(n1636), .B(n1634), .Z(n1824) );
  AND U1717 ( .A(n1825), .B(n1826), .Z(n1637) );
  OR U1718 ( .A(n1611), .B(n1613), .Z(n1826) );
  NANDN U1719 ( .A(n1614), .B(n1827), .Z(n1825) );
  NAND U1720 ( .A(n1611), .B(n1613), .Z(n1827) );
  AND U1721 ( .A(n1828), .B(n1829), .Z(n1613) );
  OR U1722 ( .A(n1587), .B(n1589), .Z(n1829) );
  NANDN U1723 ( .A(n1590), .B(n1830), .Z(n1828) );
  NAND U1724 ( .A(n1587), .B(n1589), .Z(n1830) );
  AND U1725 ( .A(n1831), .B(n1832), .Z(n1589) );
  OR U1726 ( .A(n1563), .B(n1565), .Z(n1832) );
  NANDN U1727 ( .A(n1566), .B(n1833), .Z(n1831) );
  NAND U1728 ( .A(n1563), .B(n1565), .Z(n1833) );
  AND U1729 ( .A(n1834), .B(n1835), .Z(n1565) );
  NANDN U1730 ( .A(n1541), .B(n1539), .Z(n1835) );
  NAND U1731 ( .A(n1836), .B(n1542), .Z(n1834) );
  ANDN U1732 ( .B(\stack[0][9] ), .A(n1335), .Z(n1542) );
  AND U1733 ( .A(n1837), .B(n1838), .Z(n1541) );
  OR U1734 ( .A(n1515), .B(n1517), .Z(n1838) );
  NANDN U1735 ( .A(n1518), .B(n1839), .Z(n1837) );
  NAND U1736 ( .A(n1515), .B(n1517), .Z(n1839) );
  AND U1737 ( .A(n1840), .B(n1841), .Z(n1517) );
  OR U1738 ( .A(n1491), .B(n1493), .Z(n1841) );
  NANDN U1739 ( .A(n1494), .B(n1842), .Z(n1840) );
  NAND U1740 ( .A(n1491), .B(n1493), .Z(n1842) );
  AND U1741 ( .A(n1843), .B(n1844), .Z(n1493) );
  OR U1742 ( .A(n1467), .B(n1469), .Z(n1844) );
  NANDN U1743 ( .A(n1470), .B(n1845), .Z(n1843) );
  NAND U1744 ( .A(n1467), .B(n1469), .Z(n1845) );
  AND U1745 ( .A(n1846), .B(n1847), .Z(n1469) );
  OR U1746 ( .A(n1443), .B(n1445), .Z(n1847) );
  NANDN U1747 ( .A(n1446), .B(n1848), .Z(n1846) );
  NAND U1748 ( .A(n1443), .B(n1445), .Z(n1848) );
  AND U1749 ( .A(n1849), .B(n1850), .Z(n1445) );
  OR U1750 ( .A(n1419), .B(n1421), .Z(n1850) );
  NANDN U1751 ( .A(n1422), .B(n1851), .Z(n1849) );
  NAND U1752 ( .A(n1419), .B(n1421), .Z(n1851) );
  AND U1753 ( .A(n1852), .B(n1853), .Z(n1421) );
  NANDN U1754 ( .A(n1395), .B(n1397), .Z(n1853) );
  NANDN U1755 ( .A(n1398), .B(n1854), .Z(n1852) );
  NANDN U1756 ( .A(n1397), .B(n1395), .Z(n1854) );
  XNOR U1757 ( .A(n1855), .B(n1856), .Z(n1395) );
  XNOR U1758 ( .A(n1857), .B(n1858), .Z(n1856) );
  AND U1759 ( .A(\stack[1][0] ), .B(\stack[0][3] ), .Z(n1397) );
  AND U1760 ( .A(n1859), .B(n1860), .Z(n1398) );
  NANDN U1761 ( .A(n1372), .B(n1374), .Z(n1860) );
  NANDN U1762 ( .A(n1375), .B(n1861), .Z(n1859) );
  NANDN U1763 ( .A(n1374), .B(n1372), .Z(n1861) );
  XNOR U1764 ( .A(n1862), .B(n1863), .Z(n1372) );
  NAND U1765 ( .A(\stack[0][0] ), .B(\stack[1][2] ), .Z(n1863) );
  NOR U1766 ( .A(n1351), .B(n1352), .Z(n1374) );
  NAND U1767 ( .A(\stack[1][0] ), .B(\stack[0][1] ), .Z(n1352) );
  NAND U1768 ( .A(\stack[1][1] ), .B(\stack[0][0] ), .Z(n1351) );
  NAND U1769 ( .A(\stack[1][0] ), .B(\stack[0][2] ), .Z(n1375) );
  XOR U1770 ( .A(n1864), .B(n1865), .Z(n1419) );
  XNOR U1771 ( .A(n1866), .B(n1867), .Z(n1865) );
  NAND U1772 ( .A(\stack[1][0] ), .B(\stack[0][4] ), .Z(n1422) );
  XOR U1773 ( .A(n1868), .B(n1869), .Z(n1443) );
  XOR U1774 ( .A(n1870), .B(n1871), .Z(n1869) );
  NAND U1775 ( .A(\stack[0][5] ), .B(\stack[1][0] ), .Z(n1446) );
  XOR U1776 ( .A(n1872), .B(n1873), .Z(n1467) );
  XNOR U1777 ( .A(n1874), .B(n1875), .Z(n1873) );
  NAND U1778 ( .A(\stack[1][0] ), .B(\stack[0][6] ), .Z(n1470) );
  XOR U1779 ( .A(n1876), .B(n1877), .Z(n1491) );
  XOR U1780 ( .A(n1878), .B(n1879), .Z(n1877) );
  NAND U1781 ( .A(\stack[0][7] ), .B(\stack[1][0] ), .Z(n1494) );
  XOR U1782 ( .A(n1880), .B(n1881), .Z(n1515) );
  XNOR U1783 ( .A(n1882), .B(n1883), .Z(n1881) );
  NAND U1784 ( .A(\stack[1][0] ), .B(\stack[0][8] ), .Z(n1518) );
  XOR U1785 ( .A(n1884), .B(n1885), .Z(n1539) );
  XNOR U1786 ( .A(n1886), .B(n1887), .Z(n1885) );
  XOR U1787 ( .A(n1888), .B(n1889), .Z(n1563) );
  XNOR U1788 ( .A(n1890), .B(n1891), .Z(n1889) );
  NAND U1789 ( .A(\stack[0][10] ), .B(\stack[1][0] ), .Z(n1566) );
  XOR U1790 ( .A(n1892), .B(n1893), .Z(n1587) );
  XOR U1791 ( .A(n1894), .B(n1895), .Z(n1893) );
  NAND U1792 ( .A(\stack[1][0] ), .B(\stack[0][11] ), .Z(n1590) );
  XOR U1793 ( .A(n1896), .B(n1897), .Z(n1611) );
  XNOR U1794 ( .A(n1898), .B(n1899), .Z(n1897) );
  NAND U1795 ( .A(\stack[0][12] ), .B(\stack[1][0] ), .Z(n1614) );
  NAND U1796 ( .A(n1634), .B(n1636), .Z(n1822) );
  ANDN U1797 ( .B(\stack[1][0] ), .A(n1642), .Z(n1636) );
  XNOR U1798 ( .A(n1900), .B(n1901), .Z(n1634) );
  XOR U1799 ( .A(n1902), .B(n1903), .Z(n1901) );
  NANDN U1800 ( .A(n1659), .B(n1657), .Z(n1821) );
  AND U1801 ( .A(n1904), .B(n1905), .Z(n1819) );
  NAND U1802 ( .A(\stack[0][15] ), .B(n1335), .Z(n1905) );
  IV U1803 ( .A(\stack[1][0] ), .Z(n1335) );
  NANDN U1804 ( .A(n1657), .B(n1659), .Z(n1904) );
  ANDN U1805 ( .B(\stack[1][0] ), .A(n1665), .Z(n1659) );
  IV U1806 ( .A(\stack[0][14] ), .Z(n1665) );
  XNOR U1807 ( .A(n1704), .B(n1906), .Z(n1657) );
  XNOR U1808 ( .A(n1703), .B(n1705), .Z(n1906) );
  AND U1809 ( .A(n1907), .B(n1908), .Z(n1705) );
  NANDN U1810 ( .A(n1900), .B(n1909), .Z(n1908) );
  NANDN U1811 ( .A(n1903), .B(n1910), .Z(n1907) );
  NAND U1812 ( .A(n1902), .B(n1900), .Z(n1910) );
  XOR U1813 ( .A(n1911), .B(n1912), .Z(n1900) );
  XNOR U1814 ( .A(n1913), .B(n1914), .Z(n1912) );
  IV U1815 ( .A(n1909), .Z(n1902) );
  NOR U1816 ( .A(n1619), .B(n1357), .Z(n1909) );
  AND U1817 ( .A(n1915), .B(n1916), .Z(n1903) );
  NANDN U1818 ( .A(n1896), .B(n1898), .Z(n1916) );
  NANDN U1819 ( .A(n1899), .B(n1917), .Z(n1915) );
  NANDN U1820 ( .A(n1898), .B(n1896), .Z(n1917) );
  XOR U1821 ( .A(n1918), .B(n1919), .Z(n1896) );
  XOR U1822 ( .A(n1920), .B(n1921), .Z(n1919) );
  AND U1823 ( .A(\stack[0][11] ), .B(\stack[1][1] ), .Z(n1898) );
  AND U1824 ( .A(n1922), .B(n1923), .Z(n1899) );
  NANDN U1825 ( .A(n1892), .B(n1924), .Z(n1923) );
  NANDN U1826 ( .A(n1895), .B(n1925), .Z(n1922) );
  NAND U1827 ( .A(n1894), .B(n1892), .Z(n1925) );
  XOR U1828 ( .A(n1926), .B(n1927), .Z(n1892) );
  XNOR U1829 ( .A(n1928), .B(n1929), .Z(n1927) );
  IV U1830 ( .A(n1924), .Z(n1894) );
  NOR U1831 ( .A(n1571), .B(n1357), .Z(n1924) );
  AND U1832 ( .A(n1930), .B(n1931), .Z(n1895) );
  NANDN U1833 ( .A(n1888), .B(n1890), .Z(n1931) );
  NANDN U1834 ( .A(n1891), .B(n1932), .Z(n1930) );
  NANDN U1835 ( .A(n1890), .B(n1888), .Z(n1932) );
  XOR U1836 ( .A(n1933), .B(n1934), .Z(n1888) );
  XOR U1837 ( .A(n1935), .B(n1936), .Z(n1934) );
  AND U1838 ( .A(\stack[1][1] ), .B(\stack[0][9] ), .Z(n1890) );
  AND U1839 ( .A(n1937), .B(n1938), .Z(n1891) );
  NAND U1840 ( .A(n1884), .B(n1886), .Z(n1938) );
  IV U1841 ( .A(n1939), .Z(n1884) );
  NANDN U1842 ( .A(n1887), .B(n1940), .Z(n1937) );
  NANDN U1843 ( .A(n1886), .B(n1939), .Z(n1940) );
  XNOR U1844 ( .A(n1941), .B(n1942), .Z(n1939) );
  XNOR U1845 ( .A(n1943), .B(n1944), .Z(n1942) );
  ANDN U1846 ( .B(\stack[0][8] ), .A(n1357), .Z(n1886) );
  AND U1847 ( .A(n1945), .B(n1946), .Z(n1887) );
  NANDN U1848 ( .A(n1880), .B(n1882), .Z(n1946) );
  NANDN U1849 ( .A(n1883), .B(n1947), .Z(n1945) );
  NANDN U1850 ( .A(n1882), .B(n1880), .Z(n1947) );
  XOR U1851 ( .A(n1948), .B(n1949), .Z(n1880) );
  XOR U1852 ( .A(n1950), .B(n1951), .Z(n1949) );
  AND U1853 ( .A(\stack[1][1] ), .B(\stack[0][7] ), .Z(n1882) );
  AND U1854 ( .A(n1952), .B(n1953), .Z(n1883) );
  NANDN U1855 ( .A(n1876), .B(n1954), .Z(n1953) );
  NANDN U1856 ( .A(n1879), .B(n1955), .Z(n1952) );
  NAND U1857 ( .A(n1878), .B(n1876), .Z(n1955) );
  XOR U1858 ( .A(n1956), .B(n1957), .Z(n1876) );
  XNOR U1859 ( .A(n1958), .B(n1959), .Z(n1957) );
  IV U1860 ( .A(n1954), .Z(n1878) );
  NOR U1861 ( .A(n1357), .B(n1475), .Z(n1954) );
  AND U1862 ( .A(n1960), .B(n1961), .Z(n1879) );
  NANDN U1863 ( .A(n1872), .B(n1874), .Z(n1961) );
  NANDN U1864 ( .A(n1875), .B(n1962), .Z(n1960) );
  NANDN U1865 ( .A(n1874), .B(n1872), .Z(n1962) );
  XOR U1866 ( .A(n1963), .B(n1964), .Z(n1872) );
  XOR U1867 ( .A(n1965), .B(n1966), .Z(n1964) );
  AND U1868 ( .A(\stack[1][1] ), .B(\stack[0][5] ), .Z(n1874) );
  AND U1869 ( .A(n1967), .B(n1968), .Z(n1875) );
  NANDN U1870 ( .A(n1868), .B(n1969), .Z(n1968) );
  NANDN U1871 ( .A(n1871), .B(n1970), .Z(n1967) );
  NAND U1872 ( .A(n1870), .B(n1868), .Z(n1970) );
  XOR U1873 ( .A(n1971), .B(n1972), .Z(n1868) );
  XNOR U1874 ( .A(n1973), .B(n1974), .Z(n1972) );
  IV U1875 ( .A(n1969), .Z(n1870) );
  NOR U1876 ( .A(n1357), .B(n1427), .Z(n1969) );
  AND U1877 ( .A(n1975), .B(n1976), .Z(n1871) );
  NANDN U1878 ( .A(n1864), .B(n1866), .Z(n1976) );
  NANDN U1879 ( .A(n1867), .B(n1977), .Z(n1975) );
  NANDN U1880 ( .A(n1866), .B(n1864), .Z(n1977) );
  XNOR U1881 ( .A(n1978), .B(n1979), .Z(n1864) );
  XNOR U1882 ( .A(n1980), .B(n1981), .Z(n1979) );
  AND U1883 ( .A(\stack[1][1] ), .B(\stack[0][3] ), .Z(n1866) );
  AND U1884 ( .A(n1982), .B(n1983), .Z(n1867) );
  NANDN U1885 ( .A(n1855), .B(n1857), .Z(n1983) );
  NAND U1886 ( .A(n1984), .B(n1858), .Z(n1982) );
  ANDN U1887 ( .B(n1985), .A(n1862), .Z(n1858) );
  NAND U1888 ( .A(\stack[1][1] ), .B(\stack[0][1] ), .Z(n1862) );
  AND U1889 ( .A(\stack[0][0] ), .B(\stack[1][2] ), .Z(n1985) );
  NANDN U1890 ( .A(n1857), .B(n1855), .Z(n1984) );
  XNOR U1891 ( .A(n1986), .B(n1987), .Z(n1855) );
  NAND U1892 ( .A(\stack[0][0] ), .B(\stack[1][3] ), .Z(n1987) );
  AND U1893 ( .A(\stack[1][1] ), .B(\stack[0][2] ), .Z(n1857) );
  NOR U1894 ( .A(n1642), .B(n1357), .Z(n1703) );
  IV U1895 ( .A(\stack[1][1] ), .Z(n1357) );
  IV U1896 ( .A(\stack[0][13] ), .Z(n1642) );
  XNOR U1897 ( .A(n1813), .B(n1988), .Z(n1704) );
  XNOR U1898 ( .A(n1814), .B(n1815), .Z(n1988) );
  AND U1899 ( .A(n1989), .B(n1990), .Z(n1815) );
  NANDN U1900 ( .A(n1911), .B(n1913), .Z(n1990) );
  NANDN U1901 ( .A(n1914), .B(n1991), .Z(n1989) );
  NANDN U1902 ( .A(n1913), .B(n1911), .Z(n1991) );
  XOR U1903 ( .A(n1992), .B(n1993), .Z(n1911) );
  XOR U1904 ( .A(n1994), .B(n1995), .Z(n1993) );
  AND U1905 ( .A(\stack[0][11] ), .B(\stack[1][2] ), .Z(n1913) );
  AND U1906 ( .A(n1996), .B(n1997), .Z(n1914) );
  NANDN U1907 ( .A(n1918), .B(n1998), .Z(n1997) );
  NANDN U1908 ( .A(n1921), .B(n1999), .Z(n1996) );
  NAND U1909 ( .A(n1920), .B(n1918), .Z(n1999) );
  XOR U1910 ( .A(n2000), .B(n2001), .Z(n1918) );
  XNOR U1911 ( .A(n2002), .B(n2003), .Z(n2001) );
  IV U1912 ( .A(n1998), .Z(n1920) );
  NOR U1913 ( .A(n1571), .B(n1380), .Z(n1998) );
  AND U1914 ( .A(n2004), .B(n2005), .Z(n1921) );
  NANDN U1915 ( .A(n1926), .B(n1928), .Z(n2005) );
  NANDN U1916 ( .A(n1929), .B(n2006), .Z(n2004) );
  NANDN U1917 ( .A(n1928), .B(n1926), .Z(n2006) );
  XOR U1918 ( .A(n2007), .B(n2008), .Z(n1926) );
  XOR U1919 ( .A(n2009), .B(n2010), .Z(n2008) );
  AND U1920 ( .A(\stack[1][2] ), .B(\stack[0][9] ), .Z(n1928) );
  AND U1921 ( .A(n2011), .B(n2012), .Z(n1929) );
  NANDN U1922 ( .A(n1933), .B(n2013), .Z(n2012) );
  NANDN U1923 ( .A(n1936), .B(n2014), .Z(n2011) );
  NAND U1924 ( .A(n1935), .B(n1933), .Z(n2014) );
  XOR U1925 ( .A(n2015), .B(n2016), .Z(n1933) );
  XNOR U1926 ( .A(n2017), .B(n2018), .Z(n2016) );
  IV U1927 ( .A(n2013), .Z(n1935) );
  NOR U1928 ( .A(n1523), .B(n1380), .Z(n2013) );
  AND U1929 ( .A(n2019), .B(n2020), .Z(n1936) );
  NAND U1930 ( .A(n1943), .B(n1941), .Z(n2020) );
  NANDN U1931 ( .A(n1944), .B(n2021), .Z(n2019) );
  NOR U1932 ( .A(n1380), .B(n1499), .Z(n1943) );
  XNOR U1933 ( .A(n2022), .B(n2023), .Z(n1941) );
  XNOR U1934 ( .A(n2024), .B(n2025), .Z(n2023) );
  AND U1935 ( .A(n2026), .B(n2027), .Z(n1944) );
  NANDN U1936 ( .A(n1948), .B(n2028), .Z(n2027) );
  NANDN U1937 ( .A(n1951), .B(n2029), .Z(n2026) );
  NAND U1938 ( .A(n1950), .B(n1948), .Z(n2029) );
  XOR U1939 ( .A(n2030), .B(n2031), .Z(n1948) );
  XNOR U1940 ( .A(n2032), .B(n2033), .Z(n2031) );
  IV U1941 ( .A(n2028), .Z(n1950) );
  NOR U1942 ( .A(n1380), .B(n1475), .Z(n2028) );
  AND U1943 ( .A(n2034), .B(n2035), .Z(n1951) );
  NANDN U1944 ( .A(n1956), .B(n1958), .Z(n2035) );
  NANDN U1945 ( .A(n1959), .B(n2036), .Z(n2034) );
  NANDN U1946 ( .A(n1958), .B(n1956), .Z(n2036) );
  XOR U1947 ( .A(n2037), .B(n2038), .Z(n1956) );
  XOR U1948 ( .A(n2039), .B(n2040), .Z(n2038) );
  AND U1949 ( .A(\stack[1][2] ), .B(\stack[0][5] ), .Z(n1958) );
  AND U1950 ( .A(n2041), .B(n2042), .Z(n1959) );
  NANDN U1951 ( .A(n1963), .B(n2043), .Z(n2042) );
  NANDN U1952 ( .A(n1966), .B(n2044), .Z(n2041) );
  NAND U1953 ( .A(n1965), .B(n1963), .Z(n2044) );
  XOR U1954 ( .A(n2045), .B(n2046), .Z(n1963) );
  XNOR U1955 ( .A(n2047), .B(n2048), .Z(n2046) );
  IV U1956 ( .A(n2043), .Z(n1965) );
  NOR U1957 ( .A(n1380), .B(n1427), .Z(n2043) );
  AND U1958 ( .A(n2049), .B(n2050), .Z(n1966) );
  NANDN U1959 ( .A(n1971), .B(n1973), .Z(n2050) );
  NANDN U1960 ( .A(n1974), .B(n2051), .Z(n2049) );
  NANDN U1961 ( .A(n1973), .B(n1971), .Z(n2051) );
  XNOR U1962 ( .A(n2052), .B(n2053), .Z(n1971) );
  XNOR U1963 ( .A(n2054), .B(n2055), .Z(n2053) );
  AND U1964 ( .A(\stack[1][2] ), .B(\stack[0][3] ), .Z(n1973) );
  AND U1965 ( .A(n2056), .B(n2057), .Z(n1974) );
  NANDN U1966 ( .A(n1978), .B(n1980), .Z(n2057) );
  NAND U1967 ( .A(n2058), .B(n1981), .Z(n2056) );
  ANDN U1968 ( .B(n2059), .A(n1986), .Z(n1981) );
  NAND U1969 ( .A(\stack[1][2] ), .B(\stack[0][1] ), .Z(n1986) );
  AND U1970 ( .A(\stack[0][0] ), .B(\stack[1][3] ), .Z(n2059) );
  NANDN U1971 ( .A(n1980), .B(n1978), .Z(n2058) );
  XNOR U1972 ( .A(n2060), .B(n2061), .Z(n1978) );
  NAND U1973 ( .A(\stack[0][0] ), .B(\stack[1][4] ), .Z(n2061) );
  AND U1974 ( .A(\stack[1][2] ), .B(\stack[0][2] ), .Z(n1980) );
  NOR U1975 ( .A(n1619), .B(n1380), .Z(n1814) );
  IV U1976 ( .A(\stack[1][2] ), .Z(n1380) );
  IV U1977 ( .A(\stack[0][12] ), .Z(n1619) );
  XNOR U1978 ( .A(n1716), .B(n2062), .Z(n1813) );
  XNOR U1979 ( .A(n1715), .B(n1717), .Z(n2062) );
  AND U1980 ( .A(n2063), .B(n2064), .Z(n1717) );
  NANDN U1981 ( .A(n1992), .B(n2065), .Z(n2064) );
  NANDN U1982 ( .A(n1995), .B(n2066), .Z(n2063) );
  NAND U1983 ( .A(n1994), .B(n1992), .Z(n2066) );
  XOR U1984 ( .A(n2067), .B(n2068), .Z(n1992) );
  XNOR U1985 ( .A(n2069), .B(n2070), .Z(n2068) );
  IV U1986 ( .A(n2065), .Z(n1994) );
  NOR U1987 ( .A(n1571), .B(n1404), .Z(n2065) );
  AND U1988 ( .A(n2071), .B(n2072), .Z(n1995) );
  NANDN U1989 ( .A(n2000), .B(n2002), .Z(n2072) );
  NANDN U1990 ( .A(n2003), .B(n2073), .Z(n2071) );
  NANDN U1991 ( .A(n2002), .B(n2000), .Z(n2073) );
  XOR U1992 ( .A(n2074), .B(n2075), .Z(n2000) );
  XOR U1993 ( .A(n2076), .B(n2077), .Z(n2075) );
  AND U1994 ( .A(\stack[1][3] ), .B(\stack[0][9] ), .Z(n2002) );
  AND U1995 ( .A(n2078), .B(n2079), .Z(n2003) );
  NANDN U1996 ( .A(n2007), .B(n2080), .Z(n2079) );
  NANDN U1997 ( .A(n2010), .B(n2081), .Z(n2078) );
  NAND U1998 ( .A(n2009), .B(n2007), .Z(n2081) );
  XOR U1999 ( .A(n2082), .B(n2083), .Z(n2007) );
  XNOR U2000 ( .A(n2084), .B(n2085), .Z(n2083) );
  IV U2001 ( .A(n2080), .Z(n2009) );
  NOR U2002 ( .A(n1523), .B(n1404), .Z(n2080) );
  AND U2003 ( .A(n2086), .B(n2087), .Z(n2010) );
  NANDN U2004 ( .A(n2015), .B(n2017), .Z(n2087) );
  NANDN U2005 ( .A(n2018), .B(n2088), .Z(n2086) );
  NANDN U2006 ( .A(n2017), .B(n2015), .Z(n2088) );
  XOR U2007 ( .A(n2089), .B(n2090), .Z(n2015) );
  XOR U2008 ( .A(n2091), .B(n2092), .Z(n2090) );
  AND U2009 ( .A(\stack[0][7] ), .B(\stack[1][3] ), .Z(n2017) );
  AND U2010 ( .A(n2093), .B(n2094), .Z(n2018) );
  NANDN U2011 ( .A(n2022), .B(n2024), .Z(n2094) );
  NANDN U2012 ( .A(n2025), .B(n2095), .Z(n2093) );
  NANDN U2013 ( .A(n2024), .B(n2022), .Z(n2095) );
  XNOR U2014 ( .A(n2096), .B(n2097), .Z(n2022) );
  XNOR U2015 ( .A(n2098), .B(n2099), .Z(n2097) );
  ANDN U2016 ( .B(\stack[0][6] ), .A(n1404), .Z(n2024) );
  AND U2017 ( .A(n2100), .B(n2101), .Z(n2025) );
  NANDN U2018 ( .A(n2030), .B(n2032), .Z(n2101) );
  NANDN U2019 ( .A(n2033), .B(n2102), .Z(n2100) );
  NANDN U2020 ( .A(n2032), .B(n2030), .Z(n2102) );
  XOR U2021 ( .A(n2103), .B(n2104), .Z(n2030) );
  XOR U2022 ( .A(n2105), .B(n2106), .Z(n2104) );
  AND U2023 ( .A(\stack[1][3] ), .B(\stack[0][5] ), .Z(n2032) );
  AND U2024 ( .A(n2107), .B(n2108), .Z(n2033) );
  NANDN U2025 ( .A(n2037), .B(n2109), .Z(n2108) );
  NANDN U2026 ( .A(n2040), .B(n2110), .Z(n2107) );
  NAND U2027 ( .A(n2039), .B(n2037), .Z(n2110) );
  XOR U2028 ( .A(n2111), .B(n2112), .Z(n2037) );
  XNOR U2029 ( .A(n2113), .B(n2114), .Z(n2112) );
  IV U2030 ( .A(n2109), .Z(n2039) );
  NOR U2031 ( .A(n1404), .B(n1427), .Z(n2109) );
  AND U2032 ( .A(n2115), .B(n2116), .Z(n2040) );
  NANDN U2033 ( .A(n2045), .B(n2047), .Z(n2116) );
  NANDN U2034 ( .A(n2048), .B(n2117), .Z(n2115) );
  NANDN U2035 ( .A(n2047), .B(n2045), .Z(n2117) );
  XNOR U2036 ( .A(n2118), .B(n2119), .Z(n2045) );
  XNOR U2037 ( .A(n2120), .B(n2121), .Z(n2119) );
  AND U2038 ( .A(\stack[1][3] ), .B(\stack[0][3] ), .Z(n2047) );
  AND U2039 ( .A(n2122), .B(n2123), .Z(n2048) );
  NANDN U2040 ( .A(n2052), .B(n2054), .Z(n2123) );
  NAND U2041 ( .A(n2124), .B(n2055), .Z(n2122) );
  ANDN U2042 ( .B(n2125), .A(n2060), .Z(n2055) );
  NAND U2043 ( .A(\stack[1][3] ), .B(\stack[0][1] ), .Z(n2060) );
  AND U2044 ( .A(\stack[0][0] ), .B(\stack[1][4] ), .Z(n2125) );
  NANDN U2045 ( .A(n2054), .B(n2052), .Z(n2124) );
  XNOR U2046 ( .A(n2126), .B(n2127), .Z(n2052) );
  NAND U2047 ( .A(\stack[0][0] ), .B(\stack[1][5] ), .Z(n2127) );
  AND U2048 ( .A(\stack[1][3] ), .B(\stack[0][2] ), .Z(n2054) );
  NOR U2049 ( .A(n1595), .B(n1404), .Z(n1715) );
  IV U2050 ( .A(\stack[1][3] ), .Z(n1404) );
  IV U2051 ( .A(\stack[0][11] ), .Z(n1595) );
  XNOR U2052 ( .A(n1789), .B(n2128), .Z(n1716) );
  XNOR U2053 ( .A(n1790), .B(n1791), .Z(n2128) );
  AND U2054 ( .A(n2129), .B(n2130), .Z(n1791) );
  NANDN U2055 ( .A(n2067), .B(n2069), .Z(n2130) );
  NANDN U2056 ( .A(n2070), .B(n2131), .Z(n2129) );
  NANDN U2057 ( .A(n2069), .B(n2067), .Z(n2131) );
  XOR U2058 ( .A(n2132), .B(n2133), .Z(n2067) );
  XOR U2059 ( .A(n2134), .B(n2135), .Z(n2133) );
  AND U2060 ( .A(\stack[1][4] ), .B(\stack[0][9] ), .Z(n2069) );
  AND U2061 ( .A(n2136), .B(n2137), .Z(n2070) );
  NANDN U2062 ( .A(n2074), .B(n2138), .Z(n2137) );
  NANDN U2063 ( .A(n2077), .B(n2139), .Z(n2136) );
  NAND U2064 ( .A(n2076), .B(n2074), .Z(n2139) );
  XOR U2065 ( .A(n2140), .B(n2141), .Z(n2074) );
  XNOR U2066 ( .A(n2142), .B(n2143), .Z(n2141) );
  IV U2067 ( .A(n2138), .Z(n2076) );
  NOR U2068 ( .A(n1523), .B(n1428), .Z(n2138) );
  AND U2069 ( .A(n2144), .B(n2145), .Z(n2077) );
  NANDN U2070 ( .A(n2082), .B(n2084), .Z(n2145) );
  NANDN U2071 ( .A(n2085), .B(n2146), .Z(n2144) );
  NANDN U2072 ( .A(n2084), .B(n2082), .Z(n2146) );
  XOR U2073 ( .A(n2147), .B(n2148), .Z(n2082) );
  XOR U2074 ( .A(n2149), .B(n2150), .Z(n2148) );
  AND U2075 ( .A(\stack[0][7] ), .B(\stack[1][4] ), .Z(n2084) );
  AND U2076 ( .A(n2151), .B(n2152), .Z(n2085) );
  NANDN U2077 ( .A(n2089), .B(n2153), .Z(n2152) );
  NANDN U2078 ( .A(n2092), .B(n2154), .Z(n2151) );
  NAND U2079 ( .A(n2091), .B(n2089), .Z(n2154) );
  XOR U2080 ( .A(n2155), .B(n2156), .Z(n2089) );
  XNOR U2081 ( .A(n2157), .B(n2158), .Z(n2156) );
  IV U2082 ( .A(n2153), .Z(n2091) );
  NOR U2083 ( .A(n1475), .B(n1428), .Z(n2153) );
  AND U2084 ( .A(n2159), .B(n2160), .Z(n2092) );
  NAND U2085 ( .A(n2098), .B(n2096), .Z(n2160) );
  NANDN U2086 ( .A(n2099), .B(n2161), .Z(n2159) );
  NOR U2087 ( .A(n1428), .B(n1451), .Z(n2098) );
  XNOR U2088 ( .A(n2162), .B(n2163), .Z(n2096) );
  XNOR U2089 ( .A(n2164), .B(n2165), .Z(n2163) );
  AND U2090 ( .A(n2166), .B(n2167), .Z(n2099) );
  NANDN U2091 ( .A(n2103), .B(n2168), .Z(n2167) );
  NANDN U2092 ( .A(n2106), .B(n2169), .Z(n2166) );
  NAND U2093 ( .A(n2105), .B(n2103), .Z(n2169) );
  XOR U2094 ( .A(n2170), .B(n2171), .Z(n2103) );
  XNOR U2095 ( .A(n2172), .B(n2173), .Z(n2171) );
  IV U2096 ( .A(n2168), .Z(n2105) );
  NOR U2097 ( .A(n1428), .B(n1427), .Z(n2168) );
  IV U2098 ( .A(\stack[1][4] ), .Z(n1428) );
  AND U2099 ( .A(n2174), .B(n2175), .Z(n2106) );
  NANDN U2100 ( .A(n2111), .B(n2113), .Z(n2175) );
  NANDN U2101 ( .A(n2114), .B(n2176), .Z(n2174) );
  NANDN U2102 ( .A(n2113), .B(n2111), .Z(n2176) );
  XNOR U2103 ( .A(n2177), .B(n2178), .Z(n2111) );
  XNOR U2104 ( .A(n2179), .B(n2180), .Z(n2178) );
  AND U2105 ( .A(\stack[1][4] ), .B(\stack[0][3] ), .Z(n2113) );
  AND U2106 ( .A(n2181), .B(n2182), .Z(n2114) );
  NANDN U2107 ( .A(n2118), .B(n2120), .Z(n2182) );
  NAND U2108 ( .A(n2183), .B(n2121), .Z(n2181) );
  ANDN U2109 ( .B(n2184), .A(n2126), .Z(n2121) );
  NAND U2110 ( .A(\stack[1][4] ), .B(\stack[0][1] ), .Z(n2126) );
  AND U2111 ( .A(\stack[0][0] ), .B(\stack[1][5] ), .Z(n2184) );
  NANDN U2112 ( .A(n2120), .B(n2118), .Z(n2183) );
  XNOR U2113 ( .A(n2185), .B(n2186), .Z(n2118) );
  NAND U2114 ( .A(\stack[0][0] ), .B(\stack[1][6] ), .Z(n2186) );
  AND U2115 ( .A(\stack[1][4] ), .B(\stack[0][2] ), .Z(n2120) );
  ANDN U2116 ( .B(\stack[1][4] ), .A(n1571), .Z(n1790) );
  IV U2117 ( .A(\stack[0][10] ), .Z(n1571) );
  XNOR U2118 ( .A(n1800), .B(n2187), .Z(n1789) );
  XNOR U2119 ( .A(n1799), .B(n1801), .Z(n2187) );
  AND U2120 ( .A(n2188), .B(n2189), .Z(n1801) );
  NANDN U2121 ( .A(n2132), .B(n2190), .Z(n2189) );
  NANDN U2122 ( .A(n2135), .B(n2191), .Z(n2188) );
  NAND U2123 ( .A(n2134), .B(n2132), .Z(n2191) );
  XOR U2124 ( .A(n2192), .B(n2193), .Z(n2132) );
  XNOR U2125 ( .A(n2194), .B(n2195), .Z(n2193) );
  IV U2126 ( .A(n2190), .Z(n2134) );
  NOR U2127 ( .A(n1523), .B(n1452), .Z(n2190) );
  AND U2128 ( .A(n2196), .B(n2197), .Z(n2135) );
  NANDN U2129 ( .A(n2140), .B(n2142), .Z(n2197) );
  NANDN U2130 ( .A(n2143), .B(n2198), .Z(n2196) );
  NANDN U2131 ( .A(n2142), .B(n2140), .Z(n2198) );
  XOR U2132 ( .A(n2199), .B(n2200), .Z(n2140) );
  XOR U2133 ( .A(n2201), .B(n2202), .Z(n2200) );
  AND U2134 ( .A(\stack[0][7] ), .B(\stack[1][5] ), .Z(n2142) );
  AND U2135 ( .A(n2203), .B(n2204), .Z(n2143) );
  NANDN U2136 ( .A(n2147), .B(n2205), .Z(n2204) );
  NANDN U2137 ( .A(n2150), .B(n2206), .Z(n2203) );
  NAND U2138 ( .A(n2149), .B(n2147), .Z(n2206) );
  XOR U2139 ( .A(n2207), .B(n2208), .Z(n2147) );
  XNOR U2140 ( .A(n2209), .B(n2210), .Z(n2208) );
  IV U2141 ( .A(n2205), .Z(n2149) );
  NOR U2142 ( .A(n1475), .B(n1452), .Z(n2205) );
  AND U2143 ( .A(n2211), .B(n2212), .Z(n2150) );
  NANDN U2144 ( .A(n2155), .B(n2157), .Z(n2212) );
  NANDN U2145 ( .A(n2158), .B(n2213), .Z(n2211) );
  NANDN U2146 ( .A(n2157), .B(n2155), .Z(n2213) );
  XOR U2147 ( .A(n2214), .B(n2215), .Z(n2155) );
  XOR U2148 ( .A(n2216), .B(n2217), .Z(n2215) );
  AND U2149 ( .A(\stack[0][5] ), .B(\stack[1][5] ), .Z(n2157) );
  AND U2150 ( .A(n2218), .B(n2219), .Z(n2158) );
  NANDN U2151 ( .A(n2162), .B(n2164), .Z(n2219) );
  NANDN U2152 ( .A(n2165), .B(n2220), .Z(n2218) );
  NANDN U2153 ( .A(n2164), .B(n2162), .Z(n2220) );
  XNOR U2154 ( .A(n2221), .B(n2222), .Z(n2162) );
  XNOR U2155 ( .A(n2223), .B(n2224), .Z(n2222) );
  ANDN U2156 ( .B(\stack[0][4] ), .A(n1452), .Z(n2164) );
  AND U2157 ( .A(n2225), .B(n2226), .Z(n2165) );
  NANDN U2158 ( .A(n2170), .B(n2172), .Z(n2226) );
  NANDN U2159 ( .A(n2173), .B(n2227), .Z(n2225) );
  NANDN U2160 ( .A(n2172), .B(n2170), .Z(n2227) );
  XNOR U2161 ( .A(n2228), .B(n2229), .Z(n2170) );
  XNOR U2162 ( .A(n2230), .B(n2231), .Z(n2229) );
  AND U2163 ( .A(\stack[1][5] ), .B(\stack[0][3] ), .Z(n2172) );
  AND U2164 ( .A(n2232), .B(n2233), .Z(n2173) );
  NANDN U2165 ( .A(n2177), .B(n2179), .Z(n2233) );
  NAND U2166 ( .A(n2234), .B(n2180), .Z(n2232) );
  ANDN U2167 ( .B(n2235), .A(n2185), .Z(n2180) );
  NAND U2168 ( .A(\stack[1][5] ), .B(\stack[0][1] ), .Z(n2185) );
  AND U2169 ( .A(\stack[0][0] ), .B(\stack[1][6] ), .Z(n2235) );
  NANDN U2170 ( .A(n2179), .B(n2177), .Z(n2234) );
  XNOR U2171 ( .A(n2236), .B(n2237), .Z(n2177) );
  NAND U2172 ( .A(\stack[0][0] ), .B(\stack[1][7] ), .Z(n2237) );
  AND U2173 ( .A(\stack[1][5] ), .B(\stack[0][2] ), .Z(n2179) );
  NOR U2174 ( .A(n1452), .B(n1547), .Z(n1799) );
  IV U2175 ( .A(\stack[0][9] ), .Z(n1547) );
  IV U2176 ( .A(\stack[1][5] ), .Z(n1452) );
  XNOR U2177 ( .A(n1807), .B(n2238), .Z(n1800) );
  XNOR U2178 ( .A(n1808), .B(n1809), .Z(n2238) );
  AND U2179 ( .A(n2239), .B(n2240), .Z(n1809) );
  NANDN U2180 ( .A(n2192), .B(n2194), .Z(n2240) );
  NANDN U2181 ( .A(n2195), .B(n2241), .Z(n2239) );
  NANDN U2182 ( .A(n2194), .B(n2192), .Z(n2241) );
  XOR U2183 ( .A(n2242), .B(n2243), .Z(n2192) );
  XOR U2184 ( .A(n2244), .B(n2245), .Z(n2243) );
  AND U2185 ( .A(\stack[0][7] ), .B(\stack[1][6] ), .Z(n2194) );
  AND U2186 ( .A(n2246), .B(n2247), .Z(n2195) );
  NANDN U2187 ( .A(n2199), .B(n2248), .Z(n2247) );
  NANDN U2188 ( .A(n2202), .B(n2249), .Z(n2246) );
  NAND U2189 ( .A(n2201), .B(n2199), .Z(n2249) );
  XOR U2190 ( .A(n2250), .B(n2251), .Z(n2199) );
  XNOR U2191 ( .A(n2252), .B(n2253), .Z(n2251) );
  IV U2192 ( .A(n2248), .Z(n2201) );
  NOR U2193 ( .A(n1475), .B(n1476), .Z(n2248) );
  AND U2194 ( .A(n2254), .B(n2255), .Z(n2202) );
  NANDN U2195 ( .A(n2207), .B(n2209), .Z(n2255) );
  NANDN U2196 ( .A(n2210), .B(n2256), .Z(n2254) );
  NANDN U2197 ( .A(n2209), .B(n2207), .Z(n2256) );
  XOR U2198 ( .A(n2257), .B(n2258), .Z(n2207) );
  XOR U2199 ( .A(n2259), .B(n2260), .Z(n2258) );
  AND U2200 ( .A(\stack[0][5] ), .B(\stack[1][6] ), .Z(n2209) );
  AND U2201 ( .A(n2261), .B(n2262), .Z(n2210) );
  NANDN U2202 ( .A(n2214), .B(n2263), .Z(n2262) );
  NANDN U2203 ( .A(n2217), .B(n2264), .Z(n2261) );
  NAND U2204 ( .A(n2216), .B(n2214), .Z(n2264) );
  XOR U2205 ( .A(n2265), .B(n2266), .Z(n2214) );
  XNOR U2206 ( .A(n2267), .B(n2268), .Z(n2266) );
  IV U2207 ( .A(n2263), .Z(n2216) );
  NOR U2208 ( .A(n1427), .B(n1476), .Z(n2263) );
  AND U2209 ( .A(n2269), .B(n2270), .Z(n2217) );
  NAND U2210 ( .A(n2223), .B(n2221), .Z(n2270) );
  NANDN U2211 ( .A(n2224), .B(n2271), .Z(n2269) );
  NOR U2212 ( .A(n1476), .B(n1403), .Z(n2223) );
  IV U2213 ( .A(\stack[1][6] ), .Z(n1476) );
  XNOR U2214 ( .A(n2272), .B(n2273), .Z(n2221) );
  XOR U2215 ( .A(n2274), .B(n2275), .Z(n2273) );
  AND U2216 ( .A(n2276), .B(n2277), .Z(n2224) );
  NANDN U2217 ( .A(n2228), .B(n2230), .Z(n2277) );
  NAND U2218 ( .A(n2278), .B(n2231), .Z(n2276) );
  ANDN U2219 ( .B(n2279), .A(n2236), .Z(n2231) );
  NAND U2220 ( .A(\stack[1][6] ), .B(\stack[0][1] ), .Z(n2236) );
  AND U2221 ( .A(\stack[0][0] ), .B(\stack[1][7] ), .Z(n2279) );
  NANDN U2222 ( .A(n2230), .B(n2228), .Z(n2278) );
  XNOR U2223 ( .A(n2280), .B(n2281), .Z(n2228) );
  NAND U2224 ( .A(\stack[1][8] ), .B(\stack[0][0] ), .Z(n2281) );
  AND U2225 ( .A(\stack[1][6] ), .B(\stack[0][2] ), .Z(n2230) );
  ANDN U2226 ( .B(\stack[1][6] ), .A(n1523), .Z(n1808) );
  IV U2227 ( .A(\stack[0][8] ), .Z(n1523) );
  XNOR U2228 ( .A(n1754), .B(n2282), .Z(n1807) );
  XNOR U2229 ( .A(n1753), .B(n1755), .Z(n2282) );
  AND U2230 ( .A(n2283), .B(n2284), .Z(n1755) );
  NANDN U2231 ( .A(n2242), .B(n2285), .Z(n2284) );
  NANDN U2232 ( .A(n2245), .B(n2286), .Z(n2283) );
  NAND U2233 ( .A(n2244), .B(n2242), .Z(n2286) );
  XOR U2234 ( .A(n2287), .B(n2288), .Z(n2242) );
  XNOR U2235 ( .A(n2289), .B(n2290), .Z(n2288) );
  IV U2236 ( .A(n2285), .Z(n2244) );
  NOR U2237 ( .A(n1475), .B(n1500), .Z(n2285) );
  AND U2238 ( .A(n2291), .B(n2292), .Z(n2245) );
  NANDN U2239 ( .A(n2250), .B(n2252), .Z(n2292) );
  NANDN U2240 ( .A(n2253), .B(n2293), .Z(n2291) );
  NANDN U2241 ( .A(n2252), .B(n2250), .Z(n2293) );
  XOR U2242 ( .A(n2294), .B(n2295), .Z(n2250) );
  XOR U2243 ( .A(n2296), .B(n2297), .Z(n2295) );
  AND U2244 ( .A(\stack[0][5] ), .B(\stack[1][7] ), .Z(n2252) );
  AND U2245 ( .A(n2298), .B(n2299), .Z(n2253) );
  NANDN U2246 ( .A(n2257), .B(n2300), .Z(n2299) );
  NANDN U2247 ( .A(n2260), .B(n2301), .Z(n2298) );
  NAND U2248 ( .A(n2259), .B(n2257), .Z(n2301) );
  XOR U2249 ( .A(n2302), .B(n2303), .Z(n2257) );
  XNOR U2250 ( .A(n2304), .B(n2305), .Z(n2303) );
  IV U2251 ( .A(n2300), .Z(n2259) );
  NOR U2252 ( .A(n1427), .B(n1500), .Z(n2300) );
  AND U2253 ( .A(n2306), .B(n2307), .Z(n2260) );
  NANDN U2254 ( .A(n2265), .B(n2267), .Z(n2307) );
  NANDN U2255 ( .A(n2268), .B(n2308), .Z(n2306) );
  NANDN U2256 ( .A(n2267), .B(n2265), .Z(n2308) );
  XNOR U2257 ( .A(n2309), .B(n2310), .Z(n2265) );
  XOR U2258 ( .A(n2311), .B(n2312), .Z(n2310) );
  AND U2259 ( .A(\stack[0][3] ), .B(\stack[1][7] ), .Z(n2267) );
  AND U2260 ( .A(n2313), .B(n2314), .Z(n2268) );
  NAND U2261 ( .A(n2272), .B(n2275), .Z(n2314) );
  NANDN U2262 ( .A(n2274), .B(n2315), .Z(n2313) );
  OR U2263 ( .A(n2272), .B(n2275), .Z(n2315) );
  AND U2264 ( .A(\stack[0][2] ), .B(\stack[1][7] ), .Z(n2275) );
  XOR U2265 ( .A(n2316), .B(n2317), .Z(n2272) );
  NAND U2266 ( .A(\stack[1][9] ), .B(\stack[0][0] ), .Z(n2317) );
  NANDN U2267 ( .A(n2280), .B(n2318), .Z(n2274) );
  AND U2268 ( .A(\stack[1][8] ), .B(\stack[0][0] ), .Z(n2318) );
  NAND U2269 ( .A(\stack[1][7] ), .B(\stack[0][1] ), .Z(n2280) );
  NOR U2270 ( .A(n1499), .B(n1500), .Z(n1753) );
  IV U2271 ( .A(\stack[1][7] ), .Z(n1500) );
  IV U2272 ( .A(\stack[0][7] ), .Z(n1499) );
  XNOR U2273 ( .A(n1763), .B(n2319), .Z(n1754) );
  XNOR U2274 ( .A(n1764), .B(n1765), .Z(n2319) );
  AND U2275 ( .A(n2320), .B(n2321), .Z(n1765) );
  NANDN U2276 ( .A(n2287), .B(n2289), .Z(n2321) );
  NANDN U2277 ( .A(n2290), .B(n2322), .Z(n2320) );
  NANDN U2278 ( .A(n2289), .B(n2287), .Z(n2322) );
  XOR U2279 ( .A(n2323), .B(n2324), .Z(n2287) );
  XOR U2280 ( .A(n2325), .B(n2326), .Z(n2324) );
  AND U2281 ( .A(\stack[0][5] ), .B(\stack[1][8] ), .Z(n2289) );
  AND U2282 ( .A(n2327), .B(n2328), .Z(n2290) );
  NANDN U2283 ( .A(n2294), .B(n2329), .Z(n2328) );
  NANDN U2284 ( .A(n2297), .B(n2330), .Z(n2327) );
  NAND U2285 ( .A(n2296), .B(n2294), .Z(n2330) );
  XOR U2286 ( .A(n2331), .B(n2332), .Z(n2294) );
  XNOR U2287 ( .A(n2333), .B(n2334), .Z(n2332) );
  IV U2288 ( .A(n2329), .Z(n2296) );
  NOR U2289 ( .A(n1427), .B(n1524), .Z(n2329) );
  IV U2290 ( .A(\stack[1][8] ), .Z(n1524) );
  AND U2291 ( .A(n2335), .B(n2336), .Z(n2297) );
  NANDN U2292 ( .A(n2302), .B(n2304), .Z(n2336) );
  NANDN U2293 ( .A(n2305), .B(n2337), .Z(n2335) );
  NANDN U2294 ( .A(n2304), .B(n2302), .Z(n2337) );
  XNOR U2295 ( .A(n2338), .B(n2339), .Z(n2302) );
  XNOR U2296 ( .A(n2340), .B(n2341), .Z(n2339) );
  AND U2297 ( .A(\stack[0][3] ), .B(\stack[1][8] ), .Z(n2304) );
  AND U2298 ( .A(n2342), .B(n2343), .Z(n2305) );
  NANDN U2299 ( .A(n2309), .B(n2311), .Z(n2343) );
  NANDN U2300 ( .A(n2312), .B(n2344), .Z(n2342) );
  NANDN U2301 ( .A(n2311), .B(n2309), .Z(n2344) );
  XNOR U2302 ( .A(n2345), .B(n2346), .Z(n2309) );
  NAND U2303 ( .A(\stack[0][0] ), .B(\stack[1][10] ), .Z(n2346) );
  AND U2304 ( .A(\stack[0][2] ), .B(\stack[1][8] ), .Z(n2311) );
  NANDN U2305 ( .A(n2316), .B(n2347), .Z(n2312) );
  AND U2306 ( .A(\stack[1][9] ), .B(\stack[0][0] ), .Z(n2347) );
  NAND U2307 ( .A(\stack[1][8] ), .B(\stack[0][1] ), .Z(n2316) );
  ANDN U2308 ( .B(\stack[1][8] ), .A(n1475), .Z(n1764) );
  IV U2309 ( .A(\stack[0][6] ), .Z(n1475) );
  XNOR U2310 ( .A(n1774), .B(n2348), .Z(n1763) );
  XNOR U2311 ( .A(n1773), .B(n1775), .Z(n2348) );
  AND U2312 ( .A(n2349), .B(n2350), .Z(n1775) );
  NANDN U2313 ( .A(n2323), .B(n2351), .Z(n2350) );
  NANDN U2314 ( .A(n2326), .B(n2352), .Z(n2349) );
  NAND U2315 ( .A(n2325), .B(n2323), .Z(n2352) );
  XOR U2316 ( .A(n2353), .B(n2354), .Z(n2323) );
  XNOR U2317 ( .A(n2355), .B(n2356), .Z(n2354) );
  IV U2318 ( .A(n2351), .Z(n2325) );
  NOR U2319 ( .A(n1427), .B(n1548), .Z(n2351) );
  IV U2320 ( .A(\stack[0][4] ), .Z(n1427) );
  AND U2321 ( .A(n2357), .B(n2358), .Z(n2326) );
  NANDN U2322 ( .A(n2331), .B(n2333), .Z(n2358) );
  NANDN U2323 ( .A(n2334), .B(n2359), .Z(n2357) );
  NANDN U2324 ( .A(n2333), .B(n2331), .Z(n2359) );
  XNOR U2325 ( .A(n2360), .B(n2361), .Z(n2331) );
  XNOR U2326 ( .A(n2362), .B(n2363), .Z(n2361) );
  AND U2327 ( .A(\stack[0][3] ), .B(\stack[1][9] ), .Z(n2333) );
  AND U2328 ( .A(n2364), .B(n2365), .Z(n2334) );
  NANDN U2329 ( .A(n2338), .B(n2340), .Z(n2365) );
  NAND U2330 ( .A(n2366), .B(n2341), .Z(n2364) );
  ANDN U2331 ( .B(n2367), .A(n2345), .Z(n2341) );
  NAND U2332 ( .A(\stack[0][1] ), .B(\stack[1][9] ), .Z(n2345) );
  AND U2333 ( .A(\stack[0][0] ), .B(\stack[1][10] ), .Z(n2367) );
  NANDN U2334 ( .A(n2340), .B(n2338), .Z(n2366) );
  XNOR U2335 ( .A(n2368), .B(n2369), .Z(n2338) );
  NAND U2336 ( .A(\stack[0][0] ), .B(\stack[1][11] ), .Z(n2369) );
  AND U2337 ( .A(\stack[0][2] ), .B(\stack[1][9] ), .Z(n2340) );
  NOR U2338 ( .A(n1451), .B(n1548), .Z(n1773) );
  IV U2339 ( .A(\stack[1][9] ), .Z(n1548) );
  IV U2340 ( .A(\stack[0][5] ), .Z(n1451) );
  XNOR U2341 ( .A(n1781), .B(n2370), .Z(n1774) );
  XNOR U2342 ( .A(n1782), .B(n1783), .Z(n2370) );
  AND U2343 ( .A(n2371), .B(n2372), .Z(n1783) );
  NANDN U2344 ( .A(n2353), .B(n2355), .Z(n2372) );
  NANDN U2345 ( .A(n2356), .B(n2373), .Z(n2371) );
  NANDN U2346 ( .A(n2355), .B(n2353), .Z(n2373) );
  XNOR U2347 ( .A(n2374), .B(n2375), .Z(n2353) );
  XNOR U2348 ( .A(n2376), .B(n2377), .Z(n2375) );
  AND U2349 ( .A(\stack[1][10] ), .B(\stack[0][3] ), .Z(n2355) );
  AND U2350 ( .A(n2378), .B(n2379), .Z(n2356) );
  NANDN U2351 ( .A(n2360), .B(n2362), .Z(n2379) );
  NAND U2352 ( .A(n2380), .B(n2363), .Z(n2378) );
  ANDN U2353 ( .B(n2381), .A(n2368), .Z(n2363) );
  NAND U2354 ( .A(\stack[1][10] ), .B(\stack[0][1] ), .Z(n2368) );
  AND U2355 ( .A(\stack[0][0] ), .B(\stack[1][11] ), .Z(n2381) );
  NANDN U2356 ( .A(n2362), .B(n2360), .Z(n2380) );
  XNOR U2357 ( .A(n2382), .B(n2383), .Z(n2360) );
  NAND U2358 ( .A(\stack[0][0] ), .B(\stack[1][12] ), .Z(n2383) );
  AND U2359 ( .A(\stack[1][10] ), .B(\stack[0][2] ), .Z(n2362) );
  ANDN U2360 ( .B(\stack[0][4] ), .A(n1572), .Z(n1782) );
  IV U2361 ( .A(\stack[1][10] ), .Z(n1572) );
  XNOR U2362 ( .A(n1740), .B(n2384), .Z(n1781) );
  XNOR U2363 ( .A(n1739), .B(n1741), .Z(n2384) );
  AND U2364 ( .A(n2385), .B(n2386), .Z(n1741) );
  NANDN U2365 ( .A(n2374), .B(n2376), .Z(n2386) );
  NAND U2366 ( .A(n2387), .B(n2377), .Z(n2385) );
  ANDN U2367 ( .B(n2388), .A(n2382), .Z(n2377) );
  NAND U2368 ( .A(\stack[1][11] ), .B(\stack[0][1] ), .Z(n2382) );
  AND U2369 ( .A(\stack[0][0] ), .B(\stack[1][12] ), .Z(n2388) );
  NANDN U2370 ( .A(n2376), .B(n2374), .Z(n2387) );
  XNOR U2371 ( .A(n2389), .B(n2390), .Z(n2374) );
  NAND U2372 ( .A(\stack[0][0] ), .B(\stack[1][13] ), .Z(n2390) );
  AND U2373 ( .A(\stack[1][11] ), .B(\stack[0][2] ), .Z(n2376) );
  NOR U2374 ( .A(n1596), .B(n1403), .Z(n1739) );
  IV U2375 ( .A(\stack[0][3] ), .Z(n1403) );
  IV U2376 ( .A(\stack[1][11] ), .Z(n1596) );
  XNOR U2377 ( .A(n1747), .B(n2391), .Z(n1740) );
  XOR U2378 ( .A(n1749), .B(n1748), .Z(n2391) );
  AND U2379 ( .A(\stack[1][12] ), .B(\stack[0][2] ), .Z(n1748) );
  NANDN U2380 ( .A(n2389), .B(n2392), .Z(n1749) );
  AND U2381 ( .A(\stack[0][0] ), .B(\stack[1][13] ), .Z(n2392) );
  NAND U2382 ( .A(\stack[1][12] ), .B(\stack[0][1] ), .Z(n2389) );
  XOR U2383 ( .A(n1730), .B(n2393), .Z(n1747) );
  NAND U2384 ( .A(\stack[0][0] ), .B(\stack[1][14] ), .Z(n2393) );
  NAND U2385 ( .A(\stack[1][13] ), .B(\stack[0][1] ), .Z(n1730) );
  XOR U2386 ( .A(\stack[1][15] ), .B(\stack[0][15] ), .Z(n1688) );
  AND U2387 ( .A(n2394), .B(n2395), .Z(n1681) );
  NAND U2388 ( .A(\stack[1][15] ), .B(n2396), .Z(n2395) );
  ANDN U2389 ( .B(\stack[0][15] ), .A(n1331), .Z(n2396) );
  NAND U2390 ( .A(n2397), .B(opcode[2]), .Z(n1331) );
  NAND U2391 ( .A(n2398), .B(n1333), .Z(n2394) );
  ANDN U2392 ( .B(opcode[0]), .A(n2399), .Z(n1333) );
  AND U2393 ( .A(n2400), .B(n2401), .Z(n1679) );
  NAND U2394 ( .A(\stack[0][15] ), .B(n1338), .Z(n2401) );
  ANDN U2395 ( .B(n2402), .A(opcode[0]), .Z(n1338) );
  XOR U2396 ( .A(n2403), .B(n2404), .Z(n2400) );
  XOR U2397 ( .A(n2405), .B(n2406), .Z(n2404) );
  NAND U2398 ( .A(n2407), .B(n2408), .Z(n2406) );
  NANDN U2399 ( .A(n1672), .B(n2409), .Z(n2408) );
  OR U2400 ( .A(n1671), .B(n1669), .Z(n2409) );
  AND U2401 ( .A(n2410), .B(n2411), .Z(n1672) );
  NAND U2402 ( .A(\stack[0][14] ), .B(n2412), .Z(n2411) );
  NAND U2403 ( .A(\stack[0][14] ), .B(n2413), .Z(n2410) );
  NAND U2404 ( .A(n1671), .B(n1669), .Z(n2407) );
  XOR U2405 ( .A(n2414), .B(n2415), .Z(n1669) );
  NAND U2406 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND U2407 ( .A(\stack[1][14] ), .B(n2413), .Z(n2417) );
  AND U2408 ( .A(n2418), .B(n2419), .Z(n2416) );
  NAND U2409 ( .A(\stack[0][14] ), .B(n1677), .Z(n2419) );
  NAND U2410 ( .A(\stack[1][14] ), .B(n2412), .Z(n2418) );
  NAND U2411 ( .A(n2420), .B(n2421), .Z(n1671) );
  NANDN U2412 ( .A(n1647), .B(n2422), .Z(n2421) );
  NANDN U2413 ( .A(n1648), .B(n2423), .Z(n2420) );
  NAND U2414 ( .A(n1645), .B(n1647), .Z(n2423) );
  AND U2415 ( .A(n2424), .B(n2425), .Z(n1647) );
  NANDN U2416 ( .A(n1624), .B(n2426), .Z(n2425) );
  NANDN U2417 ( .A(n1625), .B(n2427), .Z(n2424) );
  NAND U2418 ( .A(n1622), .B(n1624), .Z(n2427) );
  AND U2419 ( .A(n2428), .B(n2429), .Z(n1624) );
  NANDN U2420 ( .A(n1601), .B(n2430), .Z(n2429) );
  NANDN U2421 ( .A(n1602), .B(n2431), .Z(n2428) );
  NAND U2422 ( .A(n1599), .B(n1601), .Z(n2431) );
  AND U2423 ( .A(n2432), .B(n2433), .Z(n1601) );
  NANDN U2424 ( .A(n1577), .B(n2434), .Z(n2433) );
  NANDN U2425 ( .A(n1578), .B(n2435), .Z(n2432) );
  NAND U2426 ( .A(n1575), .B(n1577), .Z(n2435) );
  AND U2427 ( .A(n2436), .B(n2437), .Z(n1577) );
  NANDN U2428 ( .A(n1553), .B(n1551), .Z(n2437) );
  NANDN U2429 ( .A(n1554), .B(n2438), .Z(n2436) );
  AND U2430 ( .A(n2439), .B(n2440), .Z(n1553) );
  NANDN U2431 ( .A(n1529), .B(n2441), .Z(n2440) );
  NANDN U2432 ( .A(n1530), .B(n2442), .Z(n2439) );
  NAND U2433 ( .A(n1527), .B(n1529), .Z(n2442) );
  AND U2434 ( .A(n2443), .B(n2444), .Z(n1529) );
  NANDN U2435 ( .A(n1505), .B(n2445), .Z(n2444) );
  NANDN U2436 ( .A(n1506), .B(n2446), .Z(n2443) );
  NAND U2437 ( .A(n1503), .B(n1505), .Z(n2446) );
  AND U2438 ( .A(n2447), .B(n2448), .Z(n1505) );
  NANDN U2439 ( .A(n1481), .B(n2449), .Z(n2448) );
  NANDN U2440 ( .A(n1482), .B(n2450), .Z(n2447) );
  NAND U2441 ( .A(n1479), .B(n1481), .Z(n2450) );
  AND U2442 ( .A(n2451), .B(n2452), .Z(n1481) );
  NANDN U2443 ( .A(n1457), .B(n2453), .Z(n2452) );
  NANDN U2444 ( .A(n1458), .B(n2454), .Z(n2451) );
  NAND U2445 ( .A(n1455), .B(n1457), .Z(n2454) );
  AND U2446 ( .A(n2455), .B(n2456), .Z(n1457) );
  NANDN U2447 ( .A(n1433), .B(n2457), .Z(n2456) );
  NANDN U2448 ( .A(n1434), .B(n2458), .Z(n2455) );
  NAND U2449 ( .A(n1431), .B(n1433), .Z(n2458) );
  AND U2450 ( .A(n2459), .B(n2460), .Z(n1433) );
  NANDN U2451 ( .A(n1409), .B(n2461), .Z(n2460) );
  NANDN U2452 ( .A(n1410), .B(n2462), .Z(n2459) );
  NAND U2453 ( .A(n1407), .B(n1409), .Z(n2462) );
  AND U2454 ( .A(n2463), .B(n2464), .Z(n1409) );
  NANDN U2455 ( .A(n1385), .B(n2465), .Z(n2464) );
  NANDN U2456 ( .A(n1386), .B(n2466), .Z(n2463) );
  NAND U2457 ( .A(n1383), .B(n1385), .Z(n2466) );
  AND U2458 ( .A(n2467), .B(n2468), .Z(n1385) );
  NANDN U2459 ( .A(n1362), .B(n2469), .Z(n2468) );
  NANDN U2460 ( .A(n1363), .B(n2470), .Z(n2467) );
  NAND U2461 ( .A(n1360), .B(n1362), .Z(n2470) );
  AND U2462 ( .A(n2471), .B(n2472), .Z(n1362) );
  NAND U2463 ( .A(n2414), .B(n1339), .Z(n2472) );
  NANDN U2464 ( .A(n1342), .B(n2473), .Z(n2471) );
  XOR U2465 ( .A(n2414), .B(n2474), .Z(n1339) );
  NAND U2466 ( .A(n2475), .B(n2476), .Z(n2474) );
  NAND U2467 ( .A(\stack[1][0] ), .B(n2413), .Z(n2476) );
  AND U2468 ( .A(n2477), .B(n2478), .Z(n2475) );
  NAND U2469 ( .A(\stack[0][0] ), .B(n1677), .Z(n2478) );
  NAND U2470 ( .A(\stack[1][0] ), .B(n2412), .Z(n2477) );
  AND U2471 ( .A(n2479), .B(n2480), .Z(n1342) );
  NAND U2472 ( .A(\stack[0][0] ), .B(n2412), .Z(n2480) );
  NAND U2473 ( .A(\stack[0][0] ), .B(n2413), .Z(n2479) );
  IV U2474 ( .A(n2469), .Z(n1360) );
  XOR U2475 ( .A(n2414), .B(n2481), .Z(n2469) );
  NAND U2476 ( .A(n2482), .B(n2483), .Z(n2481) );
  NAND U2477 ( .A(\stack[1][1] ), .B(n2413), .Z(n2483) );
  AND U2478 ( .A(n2484), .B(n2485), .Z(n2482) );
  NAND U2479 ( .A(\stack[0][1] ), .B(n1677), .Z(n2485) );
  NAND U2480 ( .A(\stack[1][1] ), .B(n2412), .Z(n2484) );
  AND U2481 ( .A(n2486), .B(n2487), .Z(n1363) );
  NAND U2482 ( .A(\stack[0][1] ), .B(n2412), .Z(n2487) );
  NAND U2483 ( .A(\stack[0][1] ), .B(n2413), .Z(n2486) );
  IV U2484 ( .A(n2465), .Z(n1383) );
  XOR U2485 ( .A(n2414), .B(n2488), .Z(n2465) );
  NAND U2486 ( .A(n2489), .B(n2490), .Z(n2488) );
  NAND U2487 ( .A(\stack[1][2] ), .B(n2413), .Z(n2490) );
  AND U2488 ( .A(n2491), .B(n2492), .Z(n2489) );
  NAND U2489 ( .A(\stack[0][2] ), .B(n1677), .Z(n2492) );
  NAND U2490 ( .A(\stack[1][2] ), .B(n2412), .Z(n2491) );
  AND U2491 ( .A(n2493), .B(n2494), .Z(n1386) );
  NAND U2492 ( .A(\stack[0][2] ), .B(n2412), .Z(n2494) );
  NAND U2493 ( .A(\stack[0][2] ), .B(n2413), .Z(n2493) );
  IV U2494 ( .A(n2461), .Z(n1407) );
  XOR U2495 ( .A(n2414), .B(n2495), .Z(n2461) );
  NAND U2496 ( .A(n2496), .B(n2497), .Z(n2495) );
  NAND U2497 ( .A(\stack[1][3] ), .B(n2413), .Z(n2497) );
  AND U2498 ( .A(n2498), .B(n2499), .Z(n2496) );
  NAND U2499 ( .A(\stack[0][3] ), .B(n1677), .Z(n2499) );
  NAND U2500 ( .A(\stack[1][3] ), .B(n2412), .Z(n2498) );
  AND U2501 ( .A(n2500), .B(n2501), .Z(n1410) );
  NAND U2502 ( .A(\stack[0][3] ), .B(n2412), .Z(n2501) );
  NAND U2503 ( .A(\stack[0][3] ), .B(n2413), .Z(n2500) );
  IV U2504 ( .A(n2457), .Z(n1431) );
  XOR U2505 ( .A(n2414), .B(n2502), .Z(n2457) );
  NAND U2506 ( .A(n2503), .B(n2504), .Z(n2502) );
  NAND U2507 ( .A(\stack[1][4] ), .B(n2413), .Z(n2504) );
  AND U2508 ( .A(n2505), .B(n2506), .Z(n2503) );
  NAND U2509 ( .A(\stack[0][4] ), .B(n1677), .Z(n2506) );
  NAND U2510 ( .A(\stack[1][4] ), .B(n2412), .Z(n2505) );
  AND U2511 ( .A(n2507), .B(n2508), .Z(n1434) );
  NAND U2512 ( .A(\stack[0][4] ), .B(n2412), .Z(n2508) );
  NAND U2513 ( .A(\stack[0][4] ), .B(n2413), .Z(n2507) );
  IV U2514 ( .A(n2453), .Z(n1455) );
  XOR U2515 ( .A(n2414), .B(n2509), .Z(n2453) );
  NAND U2516 ( .A(n2510), .B(n2511), .Z(n2509) );
  NAND U2517 ( .A(\stack[1][5] ), .B(n2413), .Z(n2511) );
  AND U2518 ( .A(n2512), .B(n2513), .Z(n2510) );
  NAND U2519 ( .A(\stack[0][5] ), .B(n1677), .Z(n2513) );
  NAND U2520 ( .A(\stack[1][5] ), .B(n2412), .Z(n2512) );
  AND U2521 ( .A(n2514), .B(n2515), .Z(n1458) );
  NAND U2522 ( .A(\stack[0][5] ), .B(n2412), .Z(n2515) );
  NAND U2523 ( .A(\stack[0][5] ), .B(n2413), .Z(n2514) );
  IV U2524 ( .A(n2449), .Z(n1479) );
  XOR U2525 ( .A(n2414), .B(n2516), .Z(n2449) );
  NAND U2526 ( .A(n2517), .B(n2518), .Z(n2516) );
  NAND U2527 ( .A(\stack[1][6] ), .B(n2413), .Z(n2518) );
  AND U2528 ( .A(n2519), .B(n2520), .Z(n2517) );
  NAND U2529 ( .A(\stack[0][6] ), .B(n1677), .Z(n2520) );
  NAND U2530 ( .A(\stack[1][6] ), .B(n2412), .Z(n2519) );
  AND U2531 ( .A(n2521), .B(n2522), .Z(n1482) );
  NAND U2532 ( .A(\stack[0][6] ), .B(n2412), .Z(n2522) );
  NAND U2533 ( .A(\stack[0][6] ), .B(n2413), .Z(n2521) );
  IV U2534 ( .A(n2445), .Z(n1503) );
  XOR U2535 ( .A(n2414), .B(n2523), .Z(n2445) );
  NAND U2536 ( .A(n2524), .B(n2525), .Z(n2523) );
  NAND U2537 ( .A(\stack[1][7] ), .B(n2413), .Z(n2525) );
  AND U2538 ( .A(n2526), .B(n2527), .Z(n2524) );
  NAND U2539 ( .A(\stack[0][7] ), .B(n1677), .Z(n2527) );
  NAND U2540 ( .A(\stack[1][7] ), .B(n2412), .Z(n2526) );
  AND U2541 ( .A(n2528), .B(n2529), .Z(n1506) );
  NAND U2542 ( .A(\stack[0][7] ), .B(n2412), .Z(n2529) );
  NAND U2543 ( .A(\stack[0][7] ), .B(n2413), .Z(n2528) );
  IV U2544 ( .A(n2441), .Z(n1527) );
  XOR U2545 ( .A(n2414), .B(n2530), .Z(n2441) );
  NAND U2546 ( .A(n2531), .B(n2532), .Z(n2530) );
  NAND U2547 ( .A(\stack[1][8] ), .B(n2413), .Z(n2532) );
  AND U2548 ( .A(n2533), .B(n2534), .Z(n2531) );
  NAND U2549 ( .A(\stack[0][8] ), .B(n1677), .Z(n2534) );
  NAND U2550 ( .A(\stack[1][8] ), .B(n2412), .Z(n2533) );
  AND U2551 ( .A(n2535), .B(n2536), .Z(n1530) );
  NAND U2552 ( .A(\stack[0][8] ), .B(n2412), .Z(n2536) );
  NAND U2553 ( .A(\stack[0][8] ), .B(n2413), .Z(n2535) );
  XOR U2554 ( .A(n2537), .B(n1341), .Z(n1551) );
  AND U2555 ( .A(n2538), .B(n2539), .Z(n2537) );
  NAND U2556 ( .A(\stack[1][9] ), .B(n2413), .Z(n2539) );
  AND U2557 ( .A(n2540), .B(n2541), .Z(n2538) );
  NAND U2558 ( .A(\stack[0][9] ), .B(n1677), .Z(n2541) );
  NAND U2559 ( .A(\stack[1][9] ), .B(n2412), .Z(n2540) );
  AND U2560 ( .A(n2542), .B(n2543), .Z(n1554) );
  NAND U2561 ( .A(\stack[0][9] ), .B(n2412), .Z(n2543) );
  NAND U2562 ( .A(\stack[0][9] ), .B(n2413), .Z(n2542) );
  IV U2563 ( .A(n2434), .Z(n1575) );
  XOR U2564 ( .A(n2414), .B(n2544), .Z(n2434) );
  NAND U2565 ( .A(n2545), .B(n2546), .Z(n2544) );
  NAND U2566 ( .A(\stack[1][10] ), .B(n2413), .Z(n2546) );
  AND U2567 ( .A(n2547), .B(n2548), .Z(n2545) );
  NAND U2568 ( .A(\stack[0][10] ), .B(n1677), .Z(n2548) );
  NAND U2569 ( .A(\stack[1][10] ), .B(n2412), .Z(n2547) );
  AND U2570 ( .A(n2549), .B(n2550), .Z(n1578) );
  NAND U2571 ( .A(\stack[0][10] ), .B(n2412), .Z(n2550) );
  NAND U2572 ( .A(\stack[0][10] ), .B(n2413), .Z(n2549) );
  IV U2573 ( .A(n2430), .Z(n1599) );
  XOR U2574 ( .A(n2414), .B(n2551), .Z(n2430) );
  NAND U2575 ( .A(n2552), .B(n2553), .Z(n2551) );
  NAND U2576 ( .A(\stack[1][11] ), .B(n2413), .Z(n2553) );
  AND U2577 ( .A(n2554), .B(n2555), .Z(n2552) );
  NAND U2578 ( .A(\stack[0][11] ), .B(n1677), .Z(n2555) );
  NAND U2579 ( .A(\stack[1][11] ), .B(n2412), .Z(n2554) );
  AND U2580 ( .A(n2556), .B(n2557), .Z(n1602) );
  NAND U2581 ( .A(\stack[0][11] ), .B(n2412), .Z(n2557) );
  NAND U2582 ( .A(\stack[0][11] ), .B(n2413), .Z(n2556) );
  IV U2583 ( .A(n2426), .Z(n1622) );
  XOR U2584 ( .A(n2414), .B(n2558), .Z(n2426) );
  NAND U2585 ( .A(n2559), .B(n2560), .Z(n2558) );
  NAND U2586 ( .A(\stack[1][12] ), .B(n2413), .Z(n2560) );
  AND U2587 ( .A(n2561), .B(n2562), .Z(n2559) );
  NAND U2588 ( .A(\stack[0][12] ), .B(n1677), .Z(n2562) );
  NAND U2589 ( .A(\stack[1][12] ), .B(n2412), .Z(n2561) );
  AND U2590 ( .A(n2563), .B(n2564), .Z(n1625) );
  NAND U2591 ( .A(\stack[0][12] ), .B(n2412), .Z(n2564) );
  NAND U2592 ( .A(\stack[0][12] ), .B(n2413), .Z(n2563) );
  IV U2593 ( .A(n2422), .Z(n1645) );
  XOR U2594 ( .A(n2414), .B(n2565), .Z(n2422) );
  NAND U2595 ( .A(n2566), .B(n2567), .Z(n2565) );
  NAND U2596 ( .A(\stack[1][13] ), .B(n2413), .Z(n2567) );
  AND U2597 ( .A(n2568), .B(n2569), .Z(n2566) );
  NAND U2598 ( .A(\stack[0][13] ), .B(n1677), .Z(n2569) );
  NAND U2599 ( .A(\stack[1][13] ), .B(n2412), .Z(n2568) );
  IV U2600 ( .A(n1341), .Z(n2414) );
  AND U2601 ( .A(n2570), .B(n2571), .Z(n1648) );
  NAND U2602 ( .A(\stack[0][13] ), .B(n2412), .Z(n2571) );
  NAND U2603 ( .A(\stack[0][13] ), .B(n2413), .Z(n2570) );
  AND U2604 ( .A(n2572), .B(n2573), .Z(n2405) );
  NAND U2605 ( .A(\stack[0][15] ), .B(n2412), .Z(n2573) );
  NAND U2606 ( .A(\stack[0][15] ), .B(n2413), .Z(n2572) );
  XOR U2607 ( .A(n1341), .B(n2574), .Z(n2403) );
  AND U2608 ( .A(n2575), .B(n2576), .Z(n2574) );
  NAND U2609 ( .A(\stack[1][15] ), .B(n2413), .Z(n2576) );
  AND U2610 ( .A(n2577), .B(n2578), .Z(n2575) );
  NAND U2611 ( .A(\stack[0][15] ), .B(n1677), .Z(n2578) );
  NAND U2612 ( .A(\stack[1][15] ), .B(n2412), .Z(n2577) );
  NOR U2613 ( .A(n1677), .B(n2413), .Z(n1341) );
  ANDN U2614 ( .B(n2579), .A(n2397), .Z(n1677) );
  AND U2615 ( .A(n2402), .B(opcode[2]), .Z(n2579) );
  NAND U2616 ( .A(n2580), .B(n2581), .Z(n1251) );
  NAND U2617 ( .A(\stack[1][0] ), .B(n2582), .Z(n2581) );
  NAND U2618 ( .A(n2583), .B(n2584), .Z(n2580) );
  NAND U2619 ( .A(n2585), .B(n2586), .Z(n2584) );
  NAND U2620 ( .A(n1271), .B(\stack[2][0] ), .Z(n2586) );
  NAND U2621 ( .A(\stack[0][0] ), .B(n2587), .Z(n2585) );
  NAND U2622 ( .A(n2588), .B(n2589), .Z(n1250) );
  NAND U2623 ( .A(\stack[1][1] ), .B(n2582), .Z(n2589) );
  NAND U2624 ( .A(n2583), .B(n2590), .Z(n2588) );
  NAND U2625 ( .A(n2591), .B(n2592), .Z(n2590) );
  NAND U2626 ( .A(n1271), .B(\stack[2][1] ), .Z(n2592) );
  NAND U2627 ( .A(\stack[0][1] ), .B(n2587), .Z(n2591) );
  NAND U2628 ( .A(n2593), .B(n2594), .Z(n1249) );
  NAND U2629 ( .A(\stack[1][2] ), .B(n2582), .Z(n2594) );
  NAND U2630 ( .A(n2583), .B(n2595), .Z(n2593) );
  NAND U2631 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND U2632 ( .A(n1271), .B(\stack[2][2] ), .Z(n2597) );
  NAND U2633 ( .A(\stack[0][2] ), .B(n2587), .Z(n2596) );
  NAND U2634 ( .A(n2598), .B(n2599), .Z(n1248) );
  NAND U2635 ( .A(\stack[1][3] ), .B(n2582), .Z(n2599) );
  NAND U2636 ( .A(n2583), .B(n2600), .Z(n2598) );
  NAND U2637 ( .A(n2601), .B(n2602), .Z(n2600) );
  NAND U2638 ( .A(n1271), .B(\stack[2][3] ), .Z(n2602) );
  NAND U2639 ( .A(\stack[0][3] ), .B(n2587), .Z(n2601) );
  NAND U2640 ( .A(n2603), .B(n2604), .Z(n1247) );
  NAND U2641 ( .A(\stack[1][4] ), .B(n2582), .Z(n2604) );
  NAND U2642 ( .A(n2583), .B(n2605), .Z(n2603) );
  NAND U2643 ( .A(n2606), .B(n2607), .Z(n2605) );
  NAND U2644 ( .A(n1271), .B(\stack[2][4] ), .Z(n2607) );
  NAND U2645 ( .A(\stack[0][4] ), .B(n2587), .Z(n2606) );
  NAND U2646 ( .A(n2608), .B(n2609), .Z(n1246) );
  NAND U2647 ( .A(\stack[1][5] ), .B(n2582), .Z(n2609) );
  NAND U2648 ( .A(n2583), .B(n2610), .Z(n2608) );
  NAND U2649 ( .A(n2611), .B(n2612), .Z(n2610) );
  NAND U2650 ( .A(n1271), .B(\stack[2][5] ), .Z(n2612) );
  NAND U2651 ( .A(\stack[0][5] ), .B(n2587), .Z(n2611) );
  NAND U2652 ( .A(n2613), .B(n2614), .Z(n1245) );
  NAND U2653 ( .A(\stack[1][6] ), .B(n2582), .Z(n2614) );
  NAND U2654 ( .A(n2583), .B(n2615), .Z(n2613) );
  NAND U2655 ( .A(n2616), .B(n2617), .Z(n2615) );
  NAND U2656 ( .A(n1271), .B(\stack[2][6] ), .Z(n2617) );
  NAND U2657 ( .A(\stack[0][6] ), .B(n2587), .Z(n2616) );
  NAND U2658 ( .A(n2618), .B(n2619), .Z(n1244) );
  NAND U2659 ( .A(\stack[1][7] ), .B(n2582), .Z(n2619) );
  NAND U2660 ( .A(n2583), .B(n2620), .Z(n2618) );
  NAND U2661 ( .A(n2621), .B(n2622), .Z(n2620) );
  NAND U2662 ( .A(n1271), .B(\stack[2][7] ), .Z(n2622) );
  NAND U2663 ( .A(\stack[0][7] ), .B(n2587), .Z(n2621) );
  NAND U2664 ( .A(n2623), .B(n2624), .Z(n1243) );
  NAND U2665 ( .A(\stack[1][8] ), .B(n2582), .Z(n2624) );
  NAND U2666 ( .A(n2583), .B(n2625), .Z(n2623) );
  NAND U2667 ( .A(n2626), .B(n2627), .Z(n2625) );
  NAND U2668 ( .A(n1271), .B(\stack[2][8] ), .Z(n2627) );
  NAND U2669 ( .A(\stack[0][8] ), .B(n2587), .Z(n2626) );
  NAND U2670 ( .A(n2628), .B(n2629), .Z(n1242) );
  NAND U2671 ( .A(\stack[1][9] ), .B(n2582), .Z(n2629) );
  NAND U2672 ( .A(n2583), .B(n2630), .Z(n2628) );
  NAND U2673 ( .A(n2631), .B(n2632), .Z(n2630) );
  NAND U2674 ( .A(n1271), .B(\stack[2][9] ), .Z(n2632) );
  NAND U2675 ( .A(\stack[0][9] ), .B(n2587), .Z(n2631) );
  NAND U2676 ( .A(n2633), .B(n2634), .Z(n1241) );
  NAND U2677 ( .A(\stack[1][10] ), .B(n2582), .Z(n2634) );
  NAND U2678 ( .A(n2583), .B(n2635), .Z(n2633) );
  NAND U2679 ( .A(n2636), .B(n2637), .Z(n2635) );
  NAND U2680 ( .A(n1271), .B(\stack[2][10] ), .Z(n2637) );
  NAND U2681 ( .A(n2587), .B(\stack[0][10] ), .Z(n2636) );
  NAND U2682 ( .A(n2638), .B(n2639), .Z(n1240) );
  NAND U2683 ( .A(\stack[1][11] ), .B(n2582), .Z(n2639) );
  NAND U2684 ( .A(n2583), .B(n2640), .Z(n2638) );
  NAND U2685 ( .A(n2641), .B(n2642), .Z(n2640) );
  NAND U2686 ( .A(n1271), .B(\stack[2][11] ), .Z(n2642) );
  NAND U2687 ( .A(n2587), .B(\stack[0][11] ), .Z(n2641) );
  NAND U2688 ( .A(n2643), .B(n2644), .Z(n1239) );
  NAND U2689 ( .A(\stack[1][12] ), .B(n2582), .Z(n2644) );
  NAND U2690 ( .A(n2583), .B(n2645), .Z(n2643) );
  NAND U2691 ( .A(n2646), .B(n2647), .Z(n2645) );
  NAND U2692 ( .A(n1271), .B(\stack[2][12] ), .Z(n2647) );
  NAND U2693 ( .A(n2587), .B(\stack[0][12] ), .Z(n2646) );
  NAND U2694 ( .A(n2648), .B(n2649), .Z(n1238) );
  NAND U2695 ( .A(\stack[1][13] ), .B(n2582), .Z(n2649) );
  NAND U2696 ( .A(n2583), .B(n2650), .Z(n2648) );
  NAND U2697 ( .A(n2651), .B(n2652), .Z(n2650) );
  NAND U2698 ( .A(n1271), .B(\stack[2][13] ), .Z(n2652) );
  NAND U2699 ( .A(n2587), .B(\stack[0][13] ), .Z(n2651) );
  NAND U2700 ( .A(n2653), .B(n2654), .Z(n1237) );
  NAND U2701 ( .A(\stack[1][14] ), .B(n2582), .Z(n2654) );
  NAND U2702 ( .A(n2583), .B(n2655), .Z(n2653) );
  NAND U2703 ( .A(n2656), .B(n2657), .Z(n2655) );
  NAND U2704 ( .A(n1271), .B(\stack[2][14] ), .Z(n2657) );
  NAND U2705 ( .A(n2587), .B(\stack[0][14] ), .Z(n2656) );
  NAND U2706 ( .A(n2658), .B(n2659), .Z(n1236) );
  NAND U2707 ( .A(\stack[1][15] ), .B(n2582), .Z(n2659) );
  NAND U2708 ( .A(n2583), .B(n2660), .Z(n2658) );
  NAND U2709 ( .A(n2661), .B(n2662), .Z(n2660) );
  NAND U2710 ( .A(n1271), .B(\stack[2][15] ), .Z(n2662) );
  NAND U2711 ( .A(n2587), .B(\stack[0][15] ), .Z(n2661) );
  NAND U2712 ( .A(n2663), .B(n2664), .Z(n1235) );
  NAND U2713 ( .A(n2582), .B(\stack[2][0] ), .Z(n2664) );
  NAND U2714 ( .A(n2583), .B(n2665), .Z(n2663) );
  NAND U2715 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2716 ( .A(n1271), .B(\stack[3][0] ), .Z(n2667) );
  NAND U2717 ( .A(\stack[1][0] ), .B(n2587), .Z(n2666) );
  NAND U2718 ( .A(n2668), .B(n2669), .Z(n1234) );
  NAND U2719 ( .A(n2582), .B(\stack[2][1] ), .Z(n2669) );
  NAND U2720 ( .A(n2583), .B(n2670), .Z(n2668) );
  NAND U2721 ( .A(n2671), .B(n2672), .Z(n2670) );
  NAND U2722 ( .A(n1271), .B(\stack[3][1] ), .Z(n2672) );
  NAND U2723 ( .A(\stack[1][1] ), .B(n2587), .Z(n2671) );
  NAND U2724 ( .A(n2673), .B(n2674), .Z(n1233) );
  NAND U2725 ( .A(n2582), .B(\stack[2][2] ), .Z(n2674) );
  NAND U2726 ( .A(n2583), .B(n2675), .Z(n2673) );
  NAND U2727 ( .A(n2676), .B(n2677), .Z(n2675) );
  NAND U2728 ( .A(n1271), .B(\stack[3][2] ), .Z(n2677) );
  NAND U2729 ( .A(\stack[1][2] ), .B(n2587), .Z(n2676) );
  NAND U2730 ( .A(n2678), .B(n2679), .Z(n1232) );
  NAND U2731 ( .A(n2582), .B(\stack[2][3] ), .Z(n2679) );
  NAND U2732 ( .A(n2583), .B(n2680), .Z(n2678) );
  NAND U2733 ( .A(n2681), .B(n2682), .Z(n2680) );
  NAND U2734 ( .A(n1271), .B(\stack[3][3] ), .Z(n2682) );
  NAND U2735 ( .A(\stack[1][3] ), .B(n2587), .Z(n2681) );
  NAND U2736 ( .A(n2683), .B(n2684), .Z(n1231) );
  NAND U2737 ( .A(n2582), .B(\stack[2][4] ), .Z(n2684) );
  NAND U2738 ( .A(n2583), .B(n2685), .Z(n2683) );
  NAND U2739 ( .A(n2686), .B(n2687), .Z(n2685) );
  NAND U2740 ( .A(n1271), .B(\stack[3][4] ), .Z(n2687) );
  NAND U2741 ( .A(\stack[1][4] ), .B(n2587), .Z(n2686) );
  NAND U2742 ( .A(n2688), .B(n2689), .Z(n1230) );
  NAND U2743 ( .A(n2582), .B(\stack[2][5] ), .Z(n2689) );
  NAND U2744 ( .A(n2583), .B(n2690), .Z(n2688) );
  NAND U2745 ( .A(n2691), .B(n2692), .Z(n2690) );
  NAND U2746 ( .A(n1271), .B(\stack[3][5] ), .Z(n2692) );
  NAND U2747 ( .A(\stack[1][5] ), .B(n2587), .Z(n2691) );
  NAND U2748 ( .A(n2693), .B(n2694), .Z(n1229) );
  NAND U2749 ( .A(n2582), .B(\stack[2][6] ), .Z(n2694) );
  NAND U2750 ( .A(n2583), .B(n2695), .Z(n2693) );
  NAND U2751 ( .A(n2696), .B(n2697), .Z(n2695) );
  NAND U2752 ( .A(n1271), .B(\stack[3][6] ), .Z(n2697) );
  NAND U2753 ( .A(\stack[1][6] ), .B(n2587), .Z(n2696) );
  NAND U2754 ( .A(n2698), .B(n2699), .Z(n1228) );
  NAND U2755 ( .A(n2582), .B(\stack[2][7] ), .Z(n2699) );
  NAND U2756 ( .A(n2583), .B(n2700), .Z(n2698) );
  NAND U2757 ( .A(n2701), .B(n2702), .Z(n2700) );
  NAND U2758 ( .A(n1271), .B(\stack[3][7] ), .Z(n2702) );
  NAND U2759 ( .A(\stack[1][7] ), .B(n2587), .Z(n2701) );
  NAND U2760 ( .A(n2703), .B(n2704), .Z(n1227) );
  NAND U2761 ( .A(n2582), .B(\stack[2][8] ), .Z(n2704) );
  NAND U2762 ( .A(n2583), .B(n2705), .Z(n2703) );
  NAND U2763 ( .A(n2706), .B(n2707), .Z(n2705) );
  NAND U2764 ( .A(n1271), .B(\stack[3][8] ), .Z(n2707) );
  NAND U2765 ( .A(\stack[1][8] ), .B(n2587), .Z(n2706) );
  NAND U2766 ( .A(n2708), .B(n2709), .Z(n1226) );
  NAND U2767 ( .A(n2582), .B(\stack[2][9] ), .Z(n2709) );
  NAND U2768 ( .A(n2583), .B(n2710), .Z(n2708) );
  NAND U2769 ( .A(n2711), .B(n2712), .Z(n2710) );
  NAND U2770 ( .A(n1271), .B(\stack[3][9] ), .Z(n2712) );
  NAND U2771 ( .A(\stack[1][9] ), .B(n2587), .Z(n2711) );
  NAND U2772 ( .A(n2713), .B(n2714), .Z(n1225) );
  NAND U2773 ( .A(n2582), .B(\stack[2][10] ), .Z(n2714) );
  NAND U2774 ( .A(n2583), .B(n2715), .Z(n2713) );
  NAND U2775 ( .A(n2716), .B(n2717), .Z(n2715) );
  NAND U2776 ( .A(n1271), .B(\stack[3][10] ), .Z(n2717) );
  NAND U2777 ( .A(n2587), .B(\stack[1][10] ), .Z(n2716) );
  NAND U2778 ( .A(n2718), .B(n2719), .Z(n1224) );
  NAND U2779 ( .A(n2582), .B(\stack[2][11] ), .Z(n2719) );
  NAND U2780 ( .A(n2583), .B(n2720), .Z(n2718) );
  NAND U2781 ( .A(n2721), .B(n2722), .Z(n2720) );
  NAND U2782 ( .A(n1271), .B(\stack[3][11] ), .Z(n2722) );
  NAND U2783 ( .A(n2587), .B(\stack[1][11] ), .Z(n2721) );
  NAND U2784 ( .A(n2723), .B(n2724), .Z(n1223) );
  NAND U2785 ( .A(n2582), .B(\stack[2][12] ), .Z(n2724) );
  NAND U2786 ( .A(n2583), .B(n2725), .Z(n2723) );
  NAND U2787 ( .A(n2726), .B(n2727), .Z(n2725) );
  NAND U2788 ( .A(n1271), .B(\stack[3][12] ), .Z(n2727) );
  NAND U2789 ( .A(n2587), .B(\stack[1][12] ), .Z(n2726) );
  NAND U2790 ( .A(n2728), .B(n2729), .Z(n1222) );
  NAND U2791 ( .A(n2582), .B(\stack[2][13] ), .Z(n2729) );
  NAND U2792 ( .A(n2583), .B(n2730), .Z(n2728) );
  NAND U2793 ( .A(n2731), .B(n2732), .Z(n2730) );
  NAND U2794 ( .A(n1271), .B(\stack[3][13] ), .Z(n2732) );
  NAND U2795 ( .A(n2587), .B(\stack[1][13] ), .Z(n2731) );
  NAND U2796 ( .A(n2733), .B(n2734), .Z(n1221) );
  NAND U2797 ( .A(n2582), .B(\stack[2][14] ), .Z(n2734) );
  NAND U2798 ( .A(n2583), .B(n2735), .Z(n2733) );
  NAND U2799 ( .A(n2736), .B(n2737), .Z(n2735) );
  NAND U2800 ( .A(n1271), .B(\stack[3][14] ), .Z(n2737) );
  NAND U2801 ( .A(n2587), .B(\stack[1][14] ), .Z(n2736) );
  NAND U2802 ( .A(n2738), .B(n2739), .Z(n1220) );
  NAND U2803 ( .A(n2582), .B(\stack[2][15] ), .Z(n2739) );
  NAND U2804 ( .A(n2583), .B(n2740), .Z(n2738) );
  NAND U2805 ( .A(n2741), .B(n2742), .Z(n2740) );
  NAND U2806 ( .A(n1271), .B(\stack[3][15] ), .Z(n2742) );
  NAND U2807 ( .A(n2587), .B(\stack[1][15] ), .Z(n2741) );
  NAND U2808 ( .A(n2743), .B(n2744), .Z(n1219) );
  NAND U2809 ( .A(n2582), .B(\stack[3][0] ), .Z(n2744) );
  NAND U2810 ( .A(n2583), .B(n2745), .Z(n2743) );
  NAND U2811 ( .A(n2746), .B(n2747), .Z(n2745) );
  NAND U2812 ( .A(n1271), .B(\stack[4][0] ), .Z(n2747) );
  NAND U2813 ( .A(n2587), .B(\stack[2][0] ), .Z(n2746) );
  NAND U2814 ( .A(n2748), .B(n2749), .Z(n1218) );
  NAND U2815 ( .A(n2582), .B(\stack[3][1] ), .Z(n2749) );
  NAND U2816 ( .A(n2583), .B(n2750), .Z(n2748) );
  NAND U2817 ( .A(n2751), .B(n2752), .Z(n2750) );
  NAND U2818 ( .A(n1271), .B(\stack[4][1] ), .Z(n2752) );
  NAND U2819 ( .A(n2587), .B(\stack[2][1] ), .Z(n2751) );
  NAND U2820 ( .A(n2753), .B(n2754), .Z(n1217) );
  NAND U2821 ( .A(n2582), .B(\stack[3][2] ), .Z(n2754) );
  NAND U2822 ( .A(n2583), .B(n2755), .Z(n2753) );
  NAND U2823 ( .A(n2756), .B(n2757), .Z(n2755) );
  NAND U2824 ( .A(n1271), .B(\stack[4][2] ), .Z(n2757) );
  NAND U2825 ( .A(n2587), .B(\stack[2][2] ), .Z(n2756) );
  NAND U2826 ( .A(n2758), .B(n2759), .Z(n1216) );
  NAND U2827 ( .A(n2582), .B(\stack[3][3] ), .Z(n2759) );
  NAND U2828 ( .A(n2583), .B(n2760), .Z(n2758) );
  NAND U2829 ( .A(n2761), .B(n2762), .Z(n2760) );
  NAND U2830 ( .A(n1271), .B(\stack[4][3] ), .Z(n2762) );
  NAND U2831 ( .A(n2587), .B(\stack[2][3] ), .Z(n2761) );
  NAND U2832 ( .A(n2763), .B(n2764), .Z(n1215) );
  NAND U2833 ( .A(n2582), .B(\stack[3][4] ), .Z(n2764) );
  NAND U2834 ( .A(n2583), .B(n2765), .Z(n2763) );
  NAND U2835 ( .A(n2766), .B(n2767), .Z(n2765) );
  NAND U2836 ( .A(n1271), .B(\stack[4][4] ), .Z(n2767) );
  NAND U2837 ( .A(n2587), .B(\stack[2][4] ), .Z(n2766) );
  NAND U2838 ( .A(n2768), .B(n2769), .Z(n1214) );
  NAND U2839 ( .A(n2582), .B(\stack[3][5] ), .Z(n2769) );
  NAND U2840 ( .A(n2583), .B(n2770), .Z(n2768) );
  NAND U2841 ( .A(n2771), .B(n2772), .Z(n2770) );
  NAND U2842 ( .A(n1271), .B(\stack[4][5] ), .Z(n2772) );
  NAND U2843 ( .A(n2587), .B(\stack[2][5] ), .Z(n2771) );
  NAND U2844 ( .A(n2773), .B(n2774), .Z(n1213) );
  NAND U2845 ( .A(n2582), .B(\stack[3][6] ), .Z(n2774) );
  NAND U2846 ( .A(n2583), .B(n2775), .Z(n2773) );
  NAND U2847 ( .A(n2776), .B(n2777), .Z(n2775) );
  NAND U2848 ( .A(n1271), .B(\stack[4][6] ), .Z(n2777) );
  NAND U2849 ( .A(n2587), .B(\stack[2][6] ), .Z(n2776) );
  NAND U2850 ( .A(n2778), .B(n2779), .Z(n1212) );
  NAND U2851 ( .A(n2582), .B(\stack[3][7] ), .Z(n2779) );
  NAND U2852 ( .A(n2583), .B(n2780), .Z(n2778) );
  NAND U2853 ( .A(n2781), .B(n2782), .Z(n2780) );
  NAND U2854 ( .A(n1271), .B(\stack[4][7] ), .Z(n2782) );
  NAND U2855 ( .A(n2587), .B(\stack[2][7] ), .Z(n2781) );
  NAND U2856 ( .A(n2783), .B(n2784), .Z(n1211) );
  NAND U2857 ( .A(n2582), .B(\stack[3][8] ), .Z(n2784) );
  NAND U2858 ( .A(n2583), .B(n2785), .Z(n2783) );
  NAND U2859 ( .A(n2786), .B(n2787), .Z(n2785) );
  NAND U2860 ( .A(n1271), .B(\stack[4][8] ), .Z(n2787) );
  NAND U2861 ( .A(n2587), .B(\stack[2][8] ), .Z(n2786) );
  NAND U2862 ( .A(n2788), .B(n2789), .Z(n1210) );
  NAND U2863 ( .A(n2582), .B(\stack[3][9] ), .Z(n2789) );
  NAND U2864 ( .A(n2583), .B(n2790), .Z(n2788) );
  NAND U2865 ( .A(n2791), .B(n2792), .Z(n2790) );
  NAND U2866 ( .A(n1271), .B(\stack[4][9] ), .Z(n2792) );
  NAND U2867 ( .A(n2587), .B(\stack[2][9] ), .Z(n2791) );
  NAND U2868 ( .A(n2793), .B(n2794), .Z(n1209) );
  NAND U2869 ( .A(n2582), .B(\stack[3][10] ), .Z(n2794) );
  NAND U2870 ( .A(n2583), .B(n2795), .Z(n2793) );
  NAND U2871 ( .A(n2796), .B(n2797), .Z(n2795) );
  NAND U2872 ( .A(n1271), .B(\stack[4][10] ), .Z(n2797) );
  NAND U2873 ( .A(n2587), .B(\stack[2][10] ), .Z(n2796) );
  NAND U2874 ( .A(n2798), .B(n2799), .Z(n1208) );
  NAND U2875 ( .A(n2582), .B(\stack[3][11] ), .Z(n2799) );
  NAND U2876 ( .A(n2583), .B(n2800), .Z(n2798) );
  NAND U2877 ( .A(n2801), .B(n2802), .Z(n2800) );
  NAND U2878 ( .A(n1271), .B(\stack[4][11] ), .Z(n2802) );
  NAND U2879 ( .A(n2587), .B(\stack[2][11] ), .Z(n2801) );
  NAND U2880 ( .A(n2803), .B(n2804), .Z(n1207) );
  NAND U2881 ( .A(n2582), .B(\stack[3][12] ), .Z(n2804) );
  NAND U2882 ( .A(n2583), .B(n2805), .Z(n2803) );
  NAND U2883 ( .A(n2806), .B(n2807), .Z(n2805) );
  NAND U2884 ( .A(n1271), .B(\stack[4][12] ), .Z(n2807) );
  NAND U2885 ( .A(n2587), .B(\stack[2][12] ), .Z(n2806) );
  NAND U2886 ( .A(n2808), .B(n2809), .Z(n1206) );
  NAND U2887 ( .A(n2582), .B(\stack[3][13] ), .Z(n2809) );
  NAND U2888 ( .A(n2583), .B(n2810), .Z(n2808) );
  NAND U2889 ( .A(n2811), .B(n2812), .Z(n2810) );
  NAND U2890 ( .A(n1271), .B(\stack[4][13] ), .Z(n2812) );
  NAND U2891 ( .A(n2587), .B(\stack[2][13] ), .Z(n2811) );
  NAND U2892 ( .A(n2813), .B(n2814), .Z(n1205) );
  NAND U2893 ( .A(n2582), .B(\stack[3][14] ), .Z(n2814) );
  NAND U2894 ( .A(n2583), .B(n2815), .Z(n2813) );
  NAND U2895 ( .A(n2816), .B(n2817), .Z(n2815) );
  NAND U2896 ( .A(n1271), .B(\stack[4][14] ), .Z(n2817) );
  NAND U2897 ( .A(n2587), .B(\stack[2][14] ), .Z(n2816) );
  NAND U2898 ( .A(n2818), .B(n2819), .Z(n1204) );
  NAND U2899 ( .A(n2582), .B(\stack[3][15] ), .Z(n2819) );
  NAND U2900 ( .A(n2583), .B(n2820), .Z(n2818) );
  NAND U2901 ( .A(n2821), .B(n2822), .Z(n2820) );
  NAND U2902 ( .A(n1271), .B(\stack[4][15] ), .Z(n2822) );
  NAND U2903 ( .A(n2587), .B(\stack[2][15] ), .Z(n2821) );
  NAND U2904 ( .A(n2823), .B(n2824), .Z(n1203) );
  NAND U2905 ( .A(n2582), .B(\stack[4][0] ), .Z(n2824) );
  NAND U2906 ( .A(n2583), .B(n2825), .Z(n2823) );
  NAND U2907 ( .A(n2826), .B(n2827), .Z(n2825) );
  NAND U2908 ( .A(n1271), .B(\stack[5][0] ), .Z(n2827) );
  NAND U2909 ( .A(n2587), .B(\stack[3][0] ), .Z(n2826) );
  NAND U2910 ( .A(n2828), .B(n2829), .Z(n1202) );
  NAND U2911 ( .A(n2582), .B(\stack[4][1] ), .Z(n2829) );
  NAND U2912 ( .A(n2583), .B(n2830), .Z(n2828) );
  NAND U2913 ( .A(n2831), .B(n2832), .Z(n2830) );
  NAND U2914 ( .A(n1271), .B(\stack[5][1] ), .Z(n2832) );
  NAND U2915 ( .A(n2587), .B(\stack[3][1] ), .Z(n2831) );
  NAND U2916 ( .A(n2833), .B(n2834), .Z(n1201) );
  NAND U2917 ( .A(n2582), .B(\stack[4][2] ), .Z(n2834) );
  NAND U2918 ( .A(n2583), .B(n2835), .Z(n2833) );
  NAND U2919 ( .A(n2836), .B(n2837), .Z(n2835) );
  NAND U2920 ( .A(n1271), .B(\stack[5][2] ), .Z(n2837) );
  NAND U2921 ( .A(n2587), .B(\stack[3][2] ), .Z(n2836) );
  NAND U2922 ( .A(n2838), .B(n2839), .Z(n1200) );
  NAND U2923 ( .A(n2582), .B(\stack[4][3] ), .Z(n2839) );
  NAND U2924 ( .A(n2583), .B(n2840), .Z(n2838) );
  NAND U2925 ( .A(n2841), .B(n2842), .Z(n2840) );
  NAND U2926 ( .A(n1271), .B(\stack[5][3] ), .Z(n2842) );
  NAND U2927 ( .A(n2587), .B(\stack[3][3] ), .Z(n2841) );
  NAND U2928 ( .A(n2843), .B(n2844), .Z(n1199) );
  NAND U2929 ( .A(n2582), .B(\stack[4][4] ), .Z(n2844) );
  NAND U2930 ( .A(n2583), .B(n2845), .Z(n2843) );
  NAND U2931 ( .A(n2846), .B(n2847), .Z(n2845) );
  NAND U2932 ( .A(n1271), .B(\stack[5][4] ), .Z(n2847) );
  NAND U2933 ( .A(n2587), .B(\stack[3][4] ), .Z(n2846) );
  NAND U2934 ( .A(n2848), .B(n2849), .Z(n1198) );
  NAND U2935 ( .A(n2582), .B(\stack[4][5] ), .Z(n2849) );
  NAND U2936 ( .A(n2583), .B(n2850), .Z(n2848) );
  NAND U2937 ( .A(n2851), .B(n2852), .Z(n2850) );
  NAND U2938 ( .A(n1271), .B(\stack[5][5] ), .Z(n2852) );
  NAND U2939 ( .A(n2587), .B(\stack[3][5] ), .Z(n2851) );
  NAND U2940 ( .A(n2853), .B(n2854), .Z(n1197) );
  NAND U2941 ( .A(n2582), .B(\stack[4][6] ), .Z(n2854) );
  NAND U2942 ( .A(n2583), .B(n2855), .Z(n2853) );
  NAND U2943 ( .A(n2856), .B(n2857), .Z(n2855) );
  NAND U2944 ( .A(n1271), .B(\stack[5][6] ), .Z(n2857) );
  NAND U2945 ( .A(n2587), .B(\stack[3][6] ), .Z(n2856) );
  NAND U2946 ( .A(n2858), .B(n2859), .Z(n1196) );
  NAND U2947 ( .A(n2582), .B(\stack[4][7] ), .Z(n2859) );
  NAND U2948 ( .A(n2583), .B(n2860), .Z(n2858) );
  NAND U2949 ( .A(n2861), .B(n2862), .Z(n2860) );
  NAND U2950 ( .A(n1271), .B(\stack[5][7] ), .Z(n2862) );
  NAND U2951 ( .A(n2587), .B(\stack[3][7] ), .Z(n2861) );
  NAND U2952 ( .A(n2863), .B(n2864), .Z(n1195) );
  NAND U2953 ( .A(n2582), .B(\stack[4][8] ), .Z(n2864) );
  NAND U2954 ( .A(n2583), .B(n2865), .Z(n2863) );
  NAND U2955 ( .A(n2866), .B(n2867), .Z(n2865) );
  NAND U2956 ( .A(n1271), .B(\stack[5][8] ), .Z(n2867) );
  NAND U2957 ( .A(n2587), .B(\stack[3][8] ), .Z(n2866) );
  NAND U2958 ( .A(n2868), .B(n2869), .Z(n1194) );
  NAND U2959 ( .A(n2582), .B(\stack[4][9] ), .Z(n2869) );
  NAND U2960 ( .A(n2583), .B(n2870), .Z(n2868) );
  NAND U2961 ( .A(n2871), .B(n2872), .Z(n2870) );
  NAND U2962 ( .A(n1271), .B(\stack[5][9] ), .Z(n2872) );
  NAND U2963 ( .A(n2587), .B(\stack[3][9] ), .Z(n2871) );
  NAND U2964 ( .A(n2873), .B(n2874), .Z(n1193) );
  NAND U2965 ( .A(n2582), .B(\stack[4][10] ), .Z(n2874) );
  NAND U2966 ( .A(n2583), .B(n2875), .Z(n2873) );
  NAND U2967 ( .A(n2876), .B(n2877), .Z(n2875) );
  NAND U2968 ( .A(n1271), .B(\stack[5][10] ), .Z(n2877) );
  NAND U2969 ( .A(n2587), .B(\stack[3][10] ), .Z(n2876) );
  NAND U2970 ( .A(n2878), .B(n2879), .Z(n1192) );
  NAND U2971 ( .A(n2582), .B(\stack[4][11] ), .Z(n2879) );
  NAND U2972 ( .A(n2583), .B(n2880), .Z(n2878) );
  NAND U2973 ( .A(n2881), .B(n2882), .Z(n2880) );
  NAND U2974 ( .A(n1271), .B(\stack[5][11] ), .Z(n2882) );
  NAND U2975 ( .A(n2587), .B(\stack[3][11] ), .Z(n2881) );
  NAND U2976 ( .A(n2883), .B(n2884), .Z(n1191) );
  NAND U2977 ( .A(n2582), .B(\stack[4][12] ), .Z(n2884) );
  NAND U2978 ( .A(n2583), .B(n2885), .Z(n2883) );
  NAND U2979 ( .A(n2886), .B(n2887), .Z(n2885) );
  NAND U2980 ( .A(n1271), .B(\stack[5][12] ), .Z(n2887) );
  NAND U2981 ( .A(n2587), .B(\stack[3][12] ), .Z(n2886) );
  NAND U2982 ( .A(n2888), .B(n2889), .Z(n1190) );
  NAND U2983 ( .A(n2582), .B(\stack[4][13] ), .Z(n2889) );
  NAND U2984 ( .A(n2583), .B(n2890), .Z(n2888) );
  NAND U2985 ( .A(n2891), .B(n2892), .Z(n2890) );
  NAND U2986 ( .A(n1271), .B(\stack[5][13] ), .Z(n2892) );
  NAND U2987 ( .A(n2587), .B(\stack[3][13] ), .Z(n2891) );
  NAND U2988 ( .A(n2893), .B(n2894), .Z(n1189) );
  NAND U2989 ( .A(n2582), .B(\stack[4][14] ), .Z(n2894) );
  NAND U2990 ( .A(n2583), .B(n2895), .Z(n2893) );
  NAND U2991 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U2992 ( .A(n1271), .B(\stack[5][14] ), .Z(n2897) );
  NAND U2993 ( .A(n2587), .B(\stack[3][14] ), .Z(n2896) );
  NAND U2994 ( .A(n2898), .B(n2899), .Z(n1188) );
  NAND U2995 ( .A(n2582), .B(\stack[4][15] ), .Z(n2899) );
  NAND U2996 ( .A(n2583), .B(n2900), .Z(n2898) );
  NAND U2997 ( .A(n2901), .B(n2902), .Z(n2900) );
  NAND U2998 ( .A(n1271), .B(\stack[5][15] ), .Z(n2902) );
  NAND U2999 ( .A(n2587), .B(\stack[3][15] ), .Z(n2901) );
  NAND U3000 ( .A(n2903), .B(n2904), .Z(n1187) );
  NAND U3001 ( .A(n2582), .B(\stack[5][0] ), .Z(n2904) );
  NAND U3002 ( .A(n2583), .B(n2905), .Z(n2903) );
  NAND U3003 ( .A(n2906), .B(n2907), .Z(n2905) );
  NAND U3004 ( .A(n1271), .B(\stack[6][0] ), .Z(n2907) );
  NAND U3005 ( .A(n2587), .B(\stack[4][0] ), .Z(n2906) );
  NAND U3006 ( .A(n2908), .B(n2909), .Z(n1186) );
  NAND U3007 ( .A(n2582), .B(\stack[5][1] ), .Z(n2909) );
  NAND U3008 ( .A(n2583), .B(n2910), .Z(n2908) );
  NAND U3009 ( .A(n2911), .B(n2912), .Z(n2910) );
  NAND U3010 ( .A(n1271), .B(\stack[6][1] ), .Z(n2912) );
  NAND U3011 ( .A(n2587), .B(\stack[4][1] ), .Z(n2911) );
  NAND U3012 ( .A(n2913), .B(n2914), .Z(n1185) );
  NAND U3013 ( .A(n2582), .B(\stack[5][2] ), .Z(n2914) );
  NAND U3014 ( .A(n2583), .B(n2915), .Z(n2913) );
  NAND U3015 ( .A(n2916), .B(n2917), .Z(n2915) );
  NAND U3016 ( .A(n1271), .B(\stack[6][2] ), .Z(n2917) );
  NAND U3017 ( .A(n2587), .B(\stack[4][2] ), .Z(n2916) );
  NAND U3018 ( .A(n2918), .B(n2919), .Z(n1184) );
  NAND U3019 ( .A(n2582), .B(\stack[5][3] ), .Z(n2919) );
  NAND U3020 ( .A(n2583), .B(n2920), .Z(n2918) );
  NAND U3021 ( .A(n2921), .B(n2922), .Z(n2920) );
  NAND U3022 ( .A(n1271), .B(\stack[6][3] ), .Z(n2922) );
  NAND U3023 ( .A(n2587), .B(\stack[4][3] ), .Z(n2921) );
  NAND U3024 ( .A(n2923), .B(n2924), .Z(n1183) );
  NAND U3025 ( .A(n2582), .B(\stack[5][4] ), .Z(n2924) );
  NAND U3026 ( .A(n2583), .B(n2925), .Z(n2923) );
  NAND U3027 ( .A(n2926), .B(n2927), .Z(n2925) );
  NAND U3028 ( .A(n1271), .B(\stack[6][4] ), .Z(n2927) );
  NAND U3029 ( .A(n2587), .B(\stack[4][4] ), .Z(n2926) );
  NAND U3030 ( .A(n2928), .B(n2929), .Z(n1182) );
  NAND U3031 ( .A(n2582), .B(\stack[5][5] ), .Z(n2929) );
  NAND U3032 ( .A(n2583), .B(n2930), .Z(n2928) );
  NAND U3033 ( .A(n2931), .B(n2932), .Z(n2930) );
  NAND U3034 ( .A(n1271), .B(\stack[6][5] ), .Z(n2932) );
  NAND U3035 ( .A(n2587), .B(\stack[4][5] ), .Z(n2931) );
  NAND U3036 ( .A(n2933), .B(n2934), .Z(n1181) );
  NAND U3037 ( .A(n2582), .B(\stack[5][6] ), .Z(n2934) );
  NAND U3038 ( .A(n2583), .B(n2935), .Z(n2933) );
  NAND U3039 ( .A(n2936), .B(n2937), .Z(n2935) );
  NAND U3040 ( .A(n1271), .B(\stack[6][6] ), .Z(n2937) );
  NAND U3041 ( .A(n2587), .B(\stack[4][6] ), .Z(n2936) );
  NAND U3042 ( .A(n2938), .B(n2939), .Z(n1180) );
  NAND U3043 ( .A(n2582), .B(\stack[5][7] ), .Z(n2939) );
  NAND U3044 ( .A(n2583), .B(n2940), .Z(n2938) );
  NAND U3045 ( .A(n2941), .B(n2942), .Z(n2940) );
  NAND U3046 ( .A(n1271), .B(\stack[6][7] ), .Z(n2942) );
  NAND U3047 ( .A(n2587), .B(\stack[4][7] ), .Z(n2941) );
  NAND U3048 ( .A(n2943), .B(n2944), .Z(n1179) );
  NAND U3049 ( .A(n2582), .B(\stack[5][8] ), .Z(n2944) );
  NAND U3050 ( .A(n2583), .B(n2945), .Z(n2943) );
  NAND U3051 ( .A(n2946), .B(n2947), .Z(n2945) );
  NAND U3052 ( .A(n1271), .B(\stack[6][8] ), .Z(n2947) );
  NAND U3053 ( .A(n2587), .B(\stack[4][8] ), .Z(n2946) );
  NAND U3054 ( .A(n2948), .B(n2949), .Z(n1178) );
  NAND U3055 ( .A(n2582), .B(\stack[5][9] ), .Z(n2949) );
  NAND U3056 ( .A(n2583), .B(n2950), .Z(n2948) );
  NAND U3057 ( .A(n2951), .B(n2952), .Z(n2950) );
  NAND U3058 ( .A(n1271), .B(\stack[6][9] ), .Z(n2952) );
  NAND U3059 ( .A(n2587), .B(\stack[4][9] ), .Z(n2951) );
  NAND U3060 ( .A(n2953), .B(n2954), .Z(n1177) );
  NAND U3061 ( .A(n2582), .B(\stack[5][10] ), .Z(n2954) );
  NAND U3062 ( .A(n2583), .B(n2955), .Z(n2953) );
  NAND U3063 ( .A(n2956), .B(n2957), .Z(n2955) );
  NAND U3064 ( .A(n1271), .B(\stack[6][10] ), .Z(n2957) );
  NAND U3065 ( .A(n2587), .B(\stack[4][10] ), .Z(n2956) );
  NAND U3066 ( .A(n2958), .B(n2959), .Z(n1176) );
  NAND U3067 ( .A(n2582), .B(\stack[5][11] ), .Z(n2959) );
  NAND U3068 ( .A(n2583), .B(n2960), .Z(n2958) );
  NAND U3069 ( .A(n2961), .B(n2962), .Z(n2960) );
  NAND U3070 ( .A(n1271), .B(\stack[6][11] ), .Z(n2962) );
  NAND U3071 ( .A(n2587), .B(\stack[4][11] ), .Z(n2961) );
  NAND U3072 ( .A(n2963), .B(n2964), .Z(n1175) );
  NAND U3073 ( .A(n2582), .B(\stack[5][12] ), .Z(n2964) );
  NAND U3074 ( .A(n2583), .B(n2965), .Z(n2963) );
  NAND U3075 ( .A(n2966), .B(n2967), .Z(n2965) );
  NAND U3076 ( .A(n1271), .B(\stack[6][12] ), .Z(n2967) );
  NAND U3077 ( .A(n2587), .B(\stack[4][12] ), .Z(n2966) );
  NAND U3078 ( .A(n2968), .B(n2969), .Z(n1174) );
  NAND U3079 ( .A(n2582), .B(\stack[5][13] ), .Z(n2969) );
  NAND U3080 ( .A(n2583), .B(n2970), .Z(n2968) );
  NAND U3081 ( .A(n2971), .B(n2972), .Z(n2970) );
  NAND U3082 ( .A(n1271), .B(\stack[6][13] ), .Z(n2972) );
  NAND U3083 ( .A(n2587), .B(\stack[4][13] ), .Z(n2971) );
  NAND U3084 ( .A(n2973), .B(n2974), .Z(n1173) );
  NAND U3085 ( .A(n2582), .B(\stack[5][14] ), .Z(n2974) );
  NAND U3086 ( .A(n2583), .B(n2975), .Z(n2973) );
  NAND U3087 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U3088 ( .A(n1271), .B(\stack[6][14] ), .Z(n2977) );
  NAND U3089 ( .A(n2587), .B(\stack[4][14] ), .Z(n2976) );
  NAND U3090 ( .A(n2978), .B(n2979), .Z(n1172) );
  NAND U3091 ( .A(n2582), .B(\stack[5][15] ), .Z(n2979) );
  NAND U3092 ( .A(n2583), .B(n2980), .Z(n2978) );
  NAND U3093 ( .A(n2981), .B(n2982), .Z(n2980) );
  NAND U3094 ( .A(n1271), .B(\stack[6][15] ), .Z(n2982) );
  NAND U3095 ( .A(n2587), .B(\stack[4][15] ), .Z(n2981) );
  NAND U3096 ( .A(n2983), .B(n2984), .Z(n1171) );
  NAND U3097 ( .A(n2582), .B(\stack[6][0] ), .Z(n2984) );
  NAND U3098 ( .A(n2583), .B(n2985), .Z(n2983) );
  NANDN U3099 ( .A(n2986), .B(n2987), .Z(n2985) );
  NAND U3100 ( .A(n2587), .B(\stack[5][0] ), .Z(n2987) );
  NAND U3101 ( .A(n2988), .B(n2989), .Z(n1170) );
  NAND U3102 ( .A(n2582), .B(\stack[6][1] ), .Z(n2989) );
  NAND U3103 ( .A(n2583), .B(n2990), .Z(n2988) );
  NANDN U3104 ( .A(n2991), .B(n2992), .Z(n2990) );
  NAND U3105 ( .A(n2587), .B(\stack[5][1] ), .Z(n2992) );
  NAND U3106 ( .A(n2993), .B(n2994), .Z(n1169) );
  NAND U3107 ( .A(n2582), .B(\stack[6][2] ), .Z(n2994) );
  NAND U3108 ( .A(n2583), .B(n2995), .Z(n2993) );
  NANDN U3109 ( .A(n2996), .B(n2997), .Z(n2995) );
  NAND U3110 ( .A(n2587), .B(\stack[5][2] ), .Z(n2997) );
  NAND U3111 ( .A(n2998), .B(n2999), .Z(n1168) );
  NAND U3112 ( .A(n2582), .B(\stack[6][3] ), .Z(n2999) );
  NAND U3113 ( .A(n2583), .B(n3000), .Z(n2998) );
  NANDN U3114 ( .A(n3001), .B(n3002), .Z(n3000) );
  NAND U3115 ( .A(n2587), .B(\stack[5][3] ), .Z(n3002) );
  NAND U3116 ( .A(n3003), .B(n3004), .Z(n1167) );
  NAND U3117 ( .A(n2582), .B(\stack[6][4] ), .Z(n3004) );
  NAND U3118 ( .A(n2583), .B(n3005), .Z(n3003) );
  NANDN U3119 ( .A(n3006), .B(n3007), .Z(n3005) );
  NAND U3120 ( .A(n2587), .B(\stack[5][4] ), .Z(n3007) );
  NAND U3121 ( .A(n3008), .B(n3009), .Z(n1166) );
  NAND U3122 ( .A(n2582), .B(\stack[6][5] ), .Z(n3009) );
  NAND U3123 ( .A(n2583), .B(n3010), .Z(n3008) );
  NANDN U3124 ( .A(n3011), .B(n3012), .Z(n3010) );
  NAND U3125 ( .A(n2587), .B(\stack[5][5] ), .Z(n3012) );
  NAND U3126 ( .A(n3013), .B(n3014), .Z(n1165) );
  NAND U3127 ( .A(n2582), .B(\stack[6][6] ), .Z(n3014) );
  NAND U3128 ( .A(n2583), .B(n3015), .Z(n3013) );
  NANDN U3129 ( .A(n3016), .B(n3017), .Z(n3015) );
  NAND U3130 ( .A(n2587), .B(\stack[5][6] ), .Z(n3017) );
  NAND U3131 ( .A(n3018), .B(n3019), .Z(n1164) );
  NAND U3132 ( .A(n2582), .B(\stack[6][7] ), .Z(n3019) );
  NAND U3133 ( .A(n2583), .B(n3020), .Z(n3018) );
  NANDN U3134 ( .A(n3021), .B(n3022), .Z(n3020) );
  NAND U3135 ( .A(n2587), .B(\stack[5][7] ), .Z(n3022) );
  NAND U3136 ( .A(n3023), .B(n3024), .Z(n1163) );
  NAND U3137 ( .A(n2582), .B(\stack[6][8] ), .Z(n3024) );
  NAND U3138 ( .A(n2583), .B(n3025), .Z(n3023) );
  NANDN U3139 ( .A(n3026), .B(n3027), .Z(n3025) );
  NAND U3140 ( .A(n2587), .B(\stack[5][8] ), .Z(n3027) );
  NAND U3141 ( .A(n3028), .B(n3029), .Z(n1162) );
  NAND U3142 ( .A(n2582), .B(\stack[6][9] ), .Z(n3029) );
  NAND U3143 ( .A(n2583), .B(n3030), .Z(n3028) );
  NANDN U3144 ( .A(n3031), .B(n3032), .Z(n3030) );
  NAND U3145 ( .A(n2587), .B(\stack[5][9] ), .Z(n3032) );
  NAND U3146 ( .A(n3033), .B(n3034), .Z(n1161) );
  NAND U3147 ( .A(n2582), .B(\stack[6][10] ), .Z(n3034) );
  NAND U3148 ( .A(n2583), .B(n3035), .Z(n3033) );
  NANDN U3149 ( .A(n3036), .B(n3037), .Z(n3035) );
  NAND U3150 ( .A(n2587), .B(\stack[5][10] ), .Z(n3037) );
  NAND U3151 ( .A(n3038), .B(n3039), .Z(n1160) );
  NAND U3152 ( .A(n2582), .B(\stack[6][11] ), .Z(n3039) );
  NAND U3153 ( .A(n2583), .B(n3040), .Z(n3038) );
  NANDN U3154 ( .A(n3041), .B(n3042), .Z(n3040) );
  NAND U3155 ( .A(n2587), .B(\stack[5][11] ), .Z(n3042) );
  NAND U3156 ( .A(n3043), .B(n3044), .Z(n1159) );
  NAND U3157 ( .A(n2582), .B(\stack[6][12] ), .Z(n3044) );
  NAND U3158 ( .A(n2583), .B(n3045), .Z(n3043) );
  NANDN U3159 ( .A(n3046), .B(n3047), .Z(n3045) );
  NAND U3160 ( .A(n2587), .B(\stack[5][12] ), .Z(n3047) );
  NAND U3161 ( .A(n3048), .B(n3049), .Z(n1158) );
  NAND U3162 ( .A(n2582), .B(\stack[6][13] ), .Z(n3049) );
  NAND U3163 ( .A(n2583), .B(n3050), .Z(n3048) );
  NANDN U3164 ( .A(n3051), .B(n3052), .Z(n3050) );
  NAND U3165 ( .A(n2587), .B(\stack[5][13] ), .Z(n3052) );
  NAND U3166 ( .A(n3053), .B(n3054), .Z(n1157) );
  NAND U3167 ( .A(n2582), .B(\stack[6][14] ), .Z(n3054) );
  NAND U3168 ( .A(n2583), .B(n3055), .Z(n3053) );
  NANDN U3169 ( .A(n3056), .B(n3057), .Z(n3055) );
  NAND U3170 ( .A(n2587), .B(\stack[5][14] ), .Z(n3057) );
  NAND U3171 ( .A(n3058), .B(n3059), .Z(n1156) );
  NAND U3172 ( .A(n2582), .B(\stack[6][15] ), .Z(n3059) );
  NAND U3173 ( .A(n2583), .B(n3060), .Z(n3058) );
  NANDN U3174 ( .A(n3061), .B(n3062), .Z(n3060) );
  NAND U3175 ( .A(n2587), .B(\stack[5][15] ), .Z(n3062) );
  IV U3176 ( .A(n2582), .Z(n2583) );
  ANDN U3177 ( .B(n1271), .A(n1675), .Z(n2582) );
  NAND U3178 ( .A(n3063), .B(n3064), .Z(n1675) );
  NOR U3179 ( .A(n1327), .B(n2413), .Z(n3064) );
  NOR U3180 ( .A(opcode[0]), .B(n3065), .Z(n2413) );
  ANDN U3181 ( .B(opcode[0]), .A(n3065), .Z(n1327) );
  NAND U3182 ( .A(n3066), .B(opcode[1]), .Z(n3065) );
  ANDN U3183 ( .B(n2399), .A(n2412), .Z(n3063) );
  ANDN U3184 ( .B(n3067), .A(n2397), .Z(n2412) );
  AND U3185 ( .A(n2402), .B(n3066), .Z(n3067) );
  NAND U3186 ( .A(opcode[2]), .B(opcode[1]), .Z(n2399) );
  IV U3187 ( .A(n2587), .Z(n1271) );
  NANDN U3188 ( .A(n2991), .B(n3068), .Z(n1144) );
  NAND U3189 ( .A(n2587), .B(\stack[6][1] ), .Z(n3068) );
  ANDN U3190 ( .B(\stack[7][1] ), .A(n2587), .Z(n2991) );
  NANDN U3191 ( .A(n2996), .B(n3069), .Z(n1135) );
  NAND U3192 ( .A(n2587), .B(\stack[6][2] ), .Z(n3069) );
  ANDN U3193 ( .B(\stack[7][2] ), .A(n2587), .Z(n2996) );
  NANDN U3194 ( .A(n3001), .B(n3070), .Z(n1126) );
  NAND U3195 ( .A(n2587), .B(\stack[6][3] ), .Z(n3070) );
  ANDN U3196 ( .B(\stack[7][3] ), .A(n2587), .Z(n3001) );
  NANDN U3197 ( .A(n3006), .B(n3071), .Z(n1117) );
  NAND U3198 ( .A(n2587), .B(\stack[6][4] ), .Z(n3071) );
  ANDN U3199 ( .B(\stack[7][4] ), .A(n2587), .Z(n3006) );
  NANDN U3200 ( .A(n3011), .B(n3072), .Z(n1108) );
  NAND U3201 ( .A(n2587), .B(\stack[6][5] ), .Z(n3072) );
  ANDN U3202 ( .B(\stack[7][5] ), .A(n2587), .Z(n3011) );
  NANDN U3203 ( .A(n3016), .B(n3073), .Z(n1099) );
  NAND U3204 ( .A(n2587), .B(\stack[6][6] ), .Z(n3073) );
  ANDN U3205 ( .B(\stack[7][6] ), .A(n2587), .Z(n3016) );
  NANDN U3206 ( .A(n3021), .B(n3074), .Z(n1090) );
  NAND U3207 ( .A(n2587), .B(\stack[6][7] ), .Z(n3074) );
  ANDN U3208 ( .B(\stack[7][7] ), .A(n2587), .Z(n3021) );
  NANDN U3209 ( .A(n3026), .B(n3075), .Z(n1081) );
  NAND U3210 ( .A(n2587), .B(\stack[6][8] ), .Z(n3075) );
  ANDN U3211 ( .B(\stack[7][8] ), .A(n2587), .Z(n3026) );
  NANDN U3212 ( .A(n3031), .B(n3076), .Z(n1072) );
  NAND U3213 ( .A(n2587), .B(\stack[6][9] ), .Z(n3076) );
  ANDN U3214 ( .B(\stack[7][9] ), .A(n2587), .Z(n3031) );
  NANDN U3215 ( .A(n3036), .B(n3077), .Z(n1063) );
  NAND U3216 ( .A(n2587), .B(\stack[6][10] ), .Z(n3077) );
  ANDN U3217 ( .B(\stack[7][10] ), .A(n2587), .Z(n3036) );
  NANDN U3218 ( .A(n3041), .B(n3078), .Z(n1054) );
  NAND U3219 ( .A(n2587), .B(\stack[6][11] ), .Z(n3078) );
  ANDN U3220 ( .B(\stack[7][11] ), .A(n2587), .Z(n3041) );
  NANDN U3221 ( .A(n3046), .B(n3079), .Z(n1045) );
  NAND U3222 ( .A(n2587), .B(\stack[6][12] ), .Z(n3079) );
  ANDN U3223 ( .B(\stack[7][12] ), .A(n2587), .Z(n3046) );
  NANDN U3224 ( .A(n3051), .B(n3080), .Z(n1036) );
  NAND U3225 ( .A(n2587), .B(\stack[6][13] ), .Z(n3080) );
  ANDN U3226 ( .B(\stack[7][13] ), .A(n2587), .Z(n3051) );
  NANDN U3227 ( .A(n3056), .B(n3081), .Z(n1027) );
  NAND U3228 ( .A(n2587), .B(\stack[6][14] ), .Z(n3081) );
  ANDN U3229 ( .B(\stack[7][14] ), .A(n2587), .Z(n3056) );
  NANDN U3230 ( .A(n3061), .B(n3082), .Z(n1020) );
  NAND U3231 ( .A(n2587), .B(\stack[6][15] ), .Z(n3082) );
  ANDN U3232 ( .B(\stack[7][15] ), .A(n2587), .Z(n3061) );
  NANDN U3233 ( .A(n2986), .B(n3083), .Z(n1013) );
  NAND U3234 ( .A(n2587), .B(\stack[6][0] ), .Z(n3083) );
  ANDN U3235 ( .B(\stack[7][0] ), .A(n2587), .Z(n2986) );
  ANDN U3236 ( .B(n3084), .A(n3066), .Z(n2587) );
  IV U3237 ( .A(opcode[2]), .Z(n3066) );
  AND U3238 ( .A(n2397), .B(n2402), .Z(n3084) );
  IV U3239 ( .A(opcode[1]), .Z(n2402) );
  IV U3240 ( .A(opcode[0]), .Z(n2397) );
endmodule

