
module sha3_seq_CC24 ( clk, rst, in, out );
  input [575:0] in;
  output [1599:0] out;
  input clk, rst;
  wire   init, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237;
  wire   [23:0] rc_i;
  wire   [1599:0] round_reg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .I(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(n1050), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[0])
         );
  DFF \rc_i_reg[1]  ( .D(rc_i[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[1])
         );
  DFF \rc_i_reg[2]  ( .D(rc_i[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[2])
         );
  DFF \rc_i_reg[3]  ( .D(rc_i[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[3])
         );
  DFF \rc_i_reg[4]  ( .D(rc_i[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[4])
         );
  DFF \rc_i_reg[5]  ( .D(rc_i[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[5])
         );
  DFF \rc_i_reg[6]  ( .D(rc_i[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[6])
         );
  DFF \rc_i_reg[7]  ( .D(rc_i[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[7])
         );
  DFF \rc_i_reg[8]  ( .D(rc_i[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[8])
         );
  DFF \rc_i_reg[9]  ( .D(rc_i[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[9])
         );
  DFF \rc_i_reg[10]  ( .D(rc_i[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[10]) );
  DFF \rc_i_reg[11]  ( .D(rc_i[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[11]) );
  DFF \rc_i_reg[12]  ( .D(rc_i[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[12]) );
  DFF \rc_i_reg[13]  ( .D(rc_i[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[13]) );
  DFF \rc_i_reg[14]  ( .D(rc_i[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[14]) );
  DFF \rc_i_reg[15]  ( .D(rc_i[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[15]) );
  DFF \rc_i_reg[16]  ( .D(rc_i[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[16]) );
  DFF \rc_i_reg[17]  ( .D(rc_i[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[17]) );
  DFF \rc_i_reg[18]  ( .D(rc_i[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[18]) );
  DFF \rc_i_reg[19]  ( .D(rc_i[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[19]) );
  DFF \rc_i_reg[20]  ( .D(rc_i[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[20]) );
  DFF \rc_i_reg[21]  ( .D(rc_i[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[21]) );
  DFF \rc_i_reg[22]  ( .D(rc_i[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[22]) );
  DFF \rc_i_reg[23]  ( .D(rc_i[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[23]) );
  DFF \round_reg_reg[0]  ( .D(out[0]), .CLK(clk), .RST(rst), .I(in[0]), .Q(
        round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(out[1]), .CLK(clk), .RST(rst), .I(in[1]), .Q(
        round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(out[2]), .CLK(clk), .RST(rst), .I(in[2]), .Q(
        round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(out[3]), .CLK(clk), .RST(rst), .I(in[3]), .Q(
        round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(out[4]), .CLK(clk), .RST(rst), .I(in[4]), .Q(
        round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(out[5]), .CLK(clk), .RST(rst), .I(in[5]), .Q(
        round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(out[6]), .CLK(clk), .RST(rst), .I(in[6]), .Q(
        round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(out[7]), .CLK(clk), .RST(rst), .I(in[7]), .Q(
        round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(out[8]), .CLK(clk), .RST(rst), .I(in[8]), .Q(
        round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(out[9]), .CLK(clk), .RST(rst), .I(in[9]), .Q(
        round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(out[10]), .CLK(clk), .RST(rst), .I(in[10]), .Q(
        round_reg[10]) );
  DFF \round_reg_reg[11]  ( .D(out[11]), .CLK(clk), .RST(rst), .I(in[11]), .Q(
        round_reg[11]) );
  DFF \round_reg_reg[12]  ( .D(out[12]), .CLK(clk), .RST(rst), .I(in[12]), .Q(
        round_reg[12]) );
  DFF \round_reg_reg[13]  ( .D(out[13]), .CLK(clk), .RST(rst), .I(in[13]), .Q(
        round_reg[13]) );
  DFF \round_reg_reg[14]  ( .D(out[14]), .CLK(clk), .RST(rst), .I(in[14]), .Q(
        round_reg[14]) );
  DFF \round_reg_reg[15]  ( .D(out[15]), .CLK(clk), .RST(rst), .I(in[15]), .Q(
        round_reg[15]) );
  DFF \round_reg_reg[16]  ( .D(out[16]), .CLK(clk), .RST(rst), .I(in[16]), .Q(
        round_reg[16]) );
  DFF \round_reg_reg[17]  ( .D(out[17]), .CLK(clk), .RST(rst), .I(in[17]), .Q(
        round_reg[17]) );
  DFF \round_reg_reg[18]  ( .D(out[18]), .CLK(clk), .RST(rst), .I(in[18]), .Q(
        round_reg[18]) );
  DFF \round_reg_reg[19]  ( .D(out[19]), .CLK(clk), .RST(rst), .I(in[19]), .Q(
        round_reg[19]) );
  DFF \round_reg_reg[20]  ( .D(out[20]), .CLK(clk), .RST(rst), .I(in[20]), .Q(
        round_reg[20]) );
  DFF \round_reg_reg[21]  ( .D(out[21]), .CLK(clk), .RST(rst), .I(in[21]), .Q(
        round_reg[21]) );
  DFF \round_reg_reg[22]  ( .D(out[22]), .CLK(clk), .RST(rst), .I(in[22]), .Q(
        round_reg[22]) );
  DFF \round_reg_reg[23]  ( .D(out[23]), .CLK(clk), .RST(rst), .I(in[23]), .Q(
        round_reg[23]) );
  DFF \round_reg_reg[24]  ( .D(out[24]), .CLK(clk), .RST(rst), .I(in[24]), .Q(
        round_reg[24]) );
  DFF \round_reg_reg[25]  ( .D(out[25]), .CLK(clk), .RST(rst), .I(in[25]), .Q(
        round_reg[25]) );
  DFF \round_reg_reg[26]  ( .D(out[26]), .CLK(clk), .RST(rst), .I(in[26]), .Q(
        round_reg[26]) );
  DFF \round_reg_reg[27]  ( .D(out[27]), .CLK(clk), .RST(rst), .I(in[27]), .Q(
        round_reg[27]) );
  DFF \round_reg_reg[28]  ( .D(out[28]), .CLK(clk), .RST(rst), .I(in[28]), .Q(
        round_reg[28]) );
  DFF \round_reg_reg[29]  ( .D(out[29]), .CLK(clk), .RST(rst), .I(in[29]), .Q(
        round_reg[29]) );
  DFF \round_reg_reg[30]  ( .D(out[30]), .CLK(clk), .RST(rst), .I(in[30]), .Q(
        round_reg[30]) );
  DFF \round_reg_reg[31]  ( .D(out[31]), .CLK(clk), .RST(rst), .I(in[31]), .Q(
        round_reg[31]) );
  DFF \round_reg_reg[32]  ( .D(out[32]), .CLK(clk), .RST(rst), .I(in[32]), .Q(
        round_reg[32]) );
  DFF \round_reg_reg[33]  ( .D(out[33]), .CLK(clk), .RST(rst), .I(in[33]), .Q(
        round_reg[33]) );
  DFF \round_reg_reg[34]  ( .D(out[34]), .CLK(clk), .RST(rst), .I(in[34]), .Q(
        round_reg[34]) );
  DFF \round_reg_reg[35]  ( .D(out[35]), .CLK(clk), .RST(rst), .I(in[35]), .Q(
        round_reg[35]) );
  DFF \round_reg_reg[36]  ( .D(out[36]), .CLK(clk), .RST(rst), .I(in[36]), .Q(
        round_reg[36]) );
  DFF \round_reg_reg[37]  ( .D(out[37]), .CLK(clk), .RST(rst), .I(in[37]), .Q(
        round_reg[37]) );
  DFF \round_reg_reg[38]  ( .D(out[38]), .CLK(clk), .RST(rst), .I(in[38]), .Q(
        round_reg[38]) );
  DFF \round_reg_reg[39]  ( .D(out[39]), .CLK(clk), .RST(rst), .I(in[39]), .Q(
        round_reg[39]) );
  DFF \round_reg_reg[40]  ( .D(out[40]), .CLK(clk), .RST(rst), .I(in[40]), .Q(
        round_reg[40]) );
  DFF \round_reg_reg[41]  ( .D(out[41]), .CLK(clk), .RST(rst), .I(in[41]), .Q(
        round_reg[41]) );
  DFF \round_reg_reg[42]  ( .D(out[42]), .CLK(clk), .RST(rst), .I(in[42]), .Q(
        round_reg[42]) );
  DFF \round_reg_reg[43]  ( .D(out[43]), .CLK(clk), .RST(rst), .I(in[43]), .Q(
        round_reg[43]) );
  DFF \round_reg_reg[44]  ( .D(out[44]), .CLK(clk), .RST(rst), .I(in[44]), .Q(
        round_reg[44]) );
  DFF \round_reg_reg[45]  ( .D(out[45]), .CLK(clk), .RST(rst), .I(in[45]), .Q(
        round_reg[45]) );
  DFF \round_reg_reg[46]  ( .D(out[46]), .CLK(clk), .RST(rst), .I(in[46]), .Q(
        round_reg[46]) );
  DFF \round_reg_reg[47]  ( .D(out[47]), .CLK(clk), .RST(rst), .I(in[47]), .Q(
        round_reg[47]) );
  DFF \round_reg_reg[48]  ( .D(out[48]), .CLK(clk), .RST(rst), .I(in[48]), .Q(
        round_reg[48]) );
  DFF \round_reg_reg[49]  ( .D(out[49]), .CLK(clk), .RST(rst), .I(in[49]), .Q(
        round_reg[49]) );
  DFF \round_reg_reg[50]  ( .D(out[50]), .CLK(clk), .RST(rst), .I(in[50]), .Q(
        round_reg[50]) );
  DFF \round_reg_reg[51]  ( .D(out[51]), .CLK(clk), .RST(rst), .I(in[51]), .Q(
        round_reg[51]) );
  DFF \round_reg_reg[52]  ( .D(out[52]), .CLK(clk), .RST(rst), .I(in[52]), .Q(
        round_reg[52]) );
  DFF \round_reg_reg[53]  ( .D(out[53]), .CLK(clk), .RST(rst), .I(in[53]), .Q(
        round_reg[53]) );
  DFF \round_reg_reg[54]  ( .D(out[54]), .CLK(clk), .RST(rst), .I(in[54]), .Q(
        round_reg[54]) );
  DFF \round_reg_reg[55]  ( .D(out[55]), .CLK(clk), .RST(rst), .I(in[55]), .Q(
        round_reg[55]) );
  DFF \round_reg_reg[56]  ( .D(out[56]), .CLK(clk), .RST(rst), .I(in[56]), .Q(
        round_reg[56]) );
  DFF \round_reg_reg[57]  ( .D(out[57]), .CLK(clk), .RST(rst), .I(in[57]), .Q(
        round_reg[57]) );
  DFF \round_reg_reg[58]  ( .D(out[58]), .CLK(clk), .RST(rst), .I(in[58]), .Q(
        round_reg[58]) );
  DFF \round_reg_reg[59]  ( .D(out[59]), .CLK(clk), .RST(rst), .I(in[59]), .Q(
        round_reg[59]) );
  DFF \round_reg_reg[60]  ( .D(out[60]), .CLK(clk), .RST(rst), .I(in[60]), .Q(
        round_reg[60]) );
  DFF \round_reg_reg[61]  ( .D(out[61]), .CLK(clk), .RST(rst), .I(in[61]), .Q(
        round_reg[61]) );
  DFF \round_reg_reg[62]  ( .D(out[62]), .CLK(clk), .RST(rst), .I(in[62]), .Q(
        round_reg[62]) );
  DFF \round_reg_reg[63]  ( .D(out[63]), .CLK(clk), .RST(rst), .I(in[63]), .Q(
        round_reg[63]) );
  DFF \round_reg_reg[64]  ( .D(out[64]), .CLK(clk), .RST(rst), .I(in[64]), .Q(
        round_reg[64]) );
  DFF \round_reg_reg[65]  ( .D(out[65]), .CLK(clk), .RST(rst), .I(in[65]), .Q(
        round_reg[65]) );
  DFF \round_reg_reg[66]  ( .D(out[66]), .CLK(clk), .RST(rst), .I(in[66]), .Q(
        round_reg[66]) );
  DFF \round_reg_reg[67]  ( .D(out[67]), .CLK(clk), .RST(rst), .I(in[67]), .Q(
        round_reg[67]) );
  DFF \round_reg_reg[68]  ( .D(out[68]), .CLK(clk), .RST(rst), .I(in[68]), .Q(
        round_reg[68]) );
  DFF \round_reg_reg[69]  ( .D(out[69]), .CLK(clk), .RST(rst), .I(in[69]), .Q(
        round_reg[69]) );
  DFF \round_reg_reg[70]  ( .D(out[70]), .CLK(clk), .RST(rst), .I(in[70]), .Q(
        round_reg[70]) );
  DFF \round_reg_reg[71]  ( .D(out[71]), .CLK(clk), .RST(rst), .I(in[71]), .Q(
        round_reg[71]) );
  DFF \round_reg_reg[72]  ( .D(out[72]), .CLK(clk), .RST(rst), .I(in[72]), .Q(
        round_reg[72]) );
  DFF \round_reg_reg[73]  ( .D(out[73]), .CLK(clk), .RST(rst), .I(in[73]), .Q(
        round_reg[73]) );
  DFF \round_reg_reg[74]  ( .D(out[74]), .CLK(clk), .RST(rst), .I(in[74]), .Q(
        round_reg[74]) );
  DFF \round_reg_reg[75]  ( .D(out[75]), .CLK(clk), .RST(rst), .I(in[75]), .Q(
        round_reg[75]) );
  DFF \round_reg_reg[76]  ( .D(out[76]), .CLK(clk), .RST(rst), .I(in[76]), .Q(
        round_reg[76]) );
  DFF \round_reg_reg[77]  ( .D(out[77]), .CLK(clk), .RST(rst), .I(in[77]), .Q(
        round_reg[77]) );
  DFF \round_reg_reg[78]  ( .D(out[78]), .CLK(clk), .RST(rst), .I(in[78]), .Q(
        round_reg[78]) );
  DFF \round_reg_reg[79]  ( .D(out[79]), .CLK(clk), .RST(rst), .I(in[79]), .Q(
        round_reg[79]) );
  DFF \round_reg_reg[80]  ( .D(out[80]), .CLK(clk), .RST(rst), .I(in[80]), .Q(
        round_reg[80]) );
  DFF \round_reg_reg[81]  ( .D(out[81]), .CLK(clk), .RST(rst), .I(in[81]), .Q(
        round_reg[81]) );
  DFF \round_reg_reg[82]  ( .D(out[82]), .CLK(clk), .RST(rst), .I(in[82]), .Q(
        round_reg[82]) );
  DFF \round_reg_reg[83]  ( .D(out[83]), .CLK(clk), .RST(rst), .I(in[83]), .Q(
        round_reg[83]) );
  DFF \round_reg_reg[84]  ( .D(out[84]), .CLK(clk), .RST(rst), .I(in[84]), .Q(
        round_reg[84]) );
  DFF \round_reg_reg[85]  ( .D(out[85]), .CLK(clk), .RST(rst), .I(in[85]), .Q(
        round_reg[85]) );
  DFF \round_reg_reg[86]  ( .D(out[86]), .CLK(clk), .RST(rst), .I(in[86]), .Q(
        round_reg[86]) );
  DFF \round_reg_reg[87]  ( .D(out[87]), .CLK(clk), .RST(rst), .I(in[87]), .Q(
        round_reg[87]) );
  DFF \round_reg_reg[88]  ( .D(out[88]), .CLK(clk), .RST(rst), .I(in[88]), .Q(
        round_reg[88]) );
  DFF \round_reg_reg[89]  ( .D(out[89]), .CLK(clk), .RST(rst), .I(in[89]), .Q(
        round_reg[89]) );
  DFF \round_reg_reg[90]  ( .D(out[90]), .CLK(clk), .RST(rst), .I(in[90]), .Q(
        round_reg[90]) );
  DFF \round_reg_reg[91]  ( .D(out[91]), .CLK(clk), .RST(rst), .I(in[91]), .Q(
        round_reg[91]) );
  DFF \round_reg_reg[92]  ( .D(out[92]), .CLK(clk), .RST(rst), .I(in[92]), .Q(
        round_reg[92]) );
  DFF \round_reg_reg[93]  ( .D(out[93]), .CLK(clk), .RST(rst), .I(in[93]), .Q(
        round_reg[93]) );
  DFF \round_reg_reg[94]  ( .D(out[94]), .CLK(clk), .RST(rst), .I(in[94]), .Q(
        round_reg[94]) );
  DFF \round_reg_reg[95]  ( .D(out[95]), .CLK(clk), .RST(rst), .I(in[95]), .Q(
        round_reg[95]) );
  DFF \round_reg_reg[96]  ( .D(out[96]), .CLK(clk), .RST(rst), .I(in[96]), .Q(
        round_reg[96]) );
  DFF \round_reg_reg[97]  ( .D(out[97]), .CLK(clk), .RST(rst), .I(in[97]), .Q(
        round_reg[97]) );
  DFF \round_reg_reg[98]  ( .D(out[98]), .CLK(clk), .RST(rst), .I(in[98]), .Q(
        round_reg[98]) );
  DFF \round_reg_reg[99]  ( .D(out[99]), .CLK(clk), .RST(rst), .I(in[99]), .Q(
        round_reg[99]) );
  DFF \round_reg_reg[100]  ( .D(out[100]), .CLK(clk), .RST(rst), .I(in[100]), 
        .Q(round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(out[101]), .CLK(clk), .RST(rst), .I(in[101]), 
        .Q(round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(out[102]), .CLK(clk), .RST(rst), .I(in[102]), 
        .Q(round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(out[103]), .CLK(clk), .RST(rst), .I(in[103]), 
        .Q(round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(out[104]), .CLK(clk), .RST(rst), .I(in[104]), 
        .Q(round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(out[105]), .CLK(clk), .RST(rst), .I(in[105]), 
        .Q(round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(out[106]), .CLK(clk), .RST(rst), .I(in[106]), 
        .Q(round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(out[107]), .CLK(clk), .RST(rst), .I(in[107]), 
        .Q(round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(out[108]), .CLK(clk), .RST(rst), .I(in[108]), 
        .Q(round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(out[109]), .CLK(clk), .RST(rst), .I(in[109]), 
        .Q(round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(out[110]), .CLK(clk), .RST(rst), .I(in[110]), 
        .Q(round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(out[111]), .CLK(clk), .RST(rst), .I(in[111]), 
        .Q(round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(out[112]), .CLK(clk), .RST(rst), .I(in[112]), 
        .Q(round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(out[113]), .CLK(clk), .RST(rst), .I(in[113]), 
        .Q(round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(out[114]), .CLK(clk), .RST(rst), .I(in[114]), 
        .Q(round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(out[115]), .CLK(clk), .RST(rst), .I(in[115]), 
        .Q(round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(out[116]), .CLK(clk), .RST(rst), .I(in[116]), 
        .Q(round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(out[117]), .CLK(clk), .RST(rst), .I(in[117]), 
        .Q(round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(out[118]), .CLK(clk), .RST(rst), .I(in[118]), 
        .Q(round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(out[119]), .CLK(clk), .RST(rst), .I(in[119]), 
        .Q(round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(out[120]), .CLK(clk), .RST(rst), .I(in[120]), 
        .Q(round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(out[121]), .CLK(clk), .RST(rst), .I(in[121]), 
        .Q(round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(out[122]), .CLK(clk), .RST(rst), .I(in[122]), 
        .Q(round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(out[123]), .CLK(clk), .RST(rst), .I(in[123]), 
        .Q(round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(out[124]), .CLK(clk), .RST(rst), .I(in[124]), 
        .Q(round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(out[125]), .CLK(clk), .RST(rst), .I(in[125]), 
        .Q(round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(out[126]), .CLK(clk), .RST(rst), .I(in[126]), 
        .Q(round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(out[127]), .CLK(clk), .RST(rst), .I(in[127]), 
        .Q(round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(out[128]), .CLK(clk), .RST(rst), .I(in[128]), 
        .Q(round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(out[129]), .CLK(clk), .RST(rst), .I(in[129]), 
        .Q(round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(out[130]), .CLK(clk), .RST(rst), .I(in[130]), 
        .Q(round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(out[131]), .CLK(clk), .RST(rst), .I(in[131]), 
        .Q(round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(out[132]), .CLK(clk), .RST(rst), .I(in[132]), 
        .Q(round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(out[133]), .CLK(clk), .RST(rst), .I(in[133]), 
        .Q(round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(out[134]), .CLK(clk), .RST(rst), .I(in[134]), 
        .Q(round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(out[135]), .CLK(clk), .RST(rst), .I(in[135]), 
        .Q(round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(out[136]), .CLK(clk), .RST(rst), .I(in[136]), 
        .Q(round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(out[137]), .CLK(clk), .RST(rst), .I(in[137]), 
        .Q(round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(out[138]), .CLK(clk), .RST(rst), .I(in[138]), 
        .Q(round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(out[139]), .CLK(clk), .RST(rst), .I(in[139]), 
        .Q(round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(out[140]), .CLK(clk), .RST(rst), .I(in[140]), 
        .Q(round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(out[141]), .CLK(clk), .RST(rst), .I(in[141]), 
        .Q(round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(out[142]), .CLK(clk), .RST(rst), .I(in[142]), 
        .Q(round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(out[143]), .CLK(clk), .RST(rst), .I(in[143]), 
        .Q(round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(out[144]), .CLK(clk), .RST(rst), .I(in[144]), 
        .Q(round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(out[145]), .CLK(clk), .RST(rst), .I(in[145]), 
        .Q(round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(out[146]), .CLK(clk), .RST(rst), .I(in[146]), 
        .Q(round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(out[147]), .CLK(clk), .RST(rst), .I(in[147]), 
        .Q(round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(out[148]), .CLK(clk), .RST(rst), .I(in[148]), 
        .Q(round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(out[149]), .CLK(clk), .RST(rst), .I(in[149]), 
        .Q(round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(out[150]), .CLK(clk), .RST(rst), .I(in[150]), 
        .Q(round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(out[151]), .CLK(clk), .RST(rst), .I(in[151]), 
        .Q(round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(out[152]), .CLK(clk), .RST(rst), .I(in[152]), 
        .Q(round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(out[153]), .CLK(clk), .RST(rst), .I(in[153]), 
        .Q(round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(out[154]), .CLK(clk), .RST(rst), .I(in[154]), 
        .Q(round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(out[155]), .CLK(clk), .RST(rst), .I(in[155]), 
        .Q(round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(out[156]), .CLK(clk), .RST(rst), .I(in[156]), 
        .Q(round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(out[157]), .CLK(clk), .RST(rst), .I(in[157]), 
        .Q(round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(out[158]), .CLK(clk), .RST(rst), .I(in[158]), 
        .Q(round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(out[159]), .CLK(clk), .RST(rst), .I(in[159]), 
        .Q(round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(out[160]), .CLK(clk), .RST(rst), .I(in[160]), 
        .Q(round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(out[161]), .CLK(clk), .RST(rst), .I(in[161]), 
        .Q(round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(out[162]), .CLK(clk), .RST(rst), .I(in[162]), 
        .Q(round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(out[163]), .CLK(clk), .RST(rst), .I(in[163]), 
        .Q(round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(out[164]), .CLK(clk), .RST(rst), .I(in[164]), 
        .Q(round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(out[165]), .CLK(clk), .RST(rst), .I(in[165]), 
        .Q(round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(out[166]), .CLK(clk), .RST(rst), .I(in[166]), 
        .Q(round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(out[167]), .CLK(clk), .RST(rst), .I(in[167]), 
        .Q(round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(out[168]), .CLK(clk), .RST(rst), .I(in[168]), 
        .Q(round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(out[169]), .CLK(clk), .RST(rst), .I(in[169]), 
        .Q(round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(out[170]), .CLK(clk), .RST(rst), .I(in[170]), 
        .Q(round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(out[171]), .CLK(clk), .RST(rst), .I(in[171]), 
        .Q(round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(out[172]), .CLK(clk), .RST(rst), .I(in[172]), 
        .Q(round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(out[173]), .CLK(clk), .RST(rst), .I(in[173]), 
        .Q(round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(out[174]), .CLK(clk), .RST(rst), .I(in[174]), 
        .Q(round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(out[175]), .CLK(clk), .RST(rst), .I(in[175]), 
        .Q(round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(out[176]), .CLK(clk), .RST(rst), .I(in[176]), 
        .Q(round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(out[177]), .CLK(clk), .RST(rst), .I(in[177]), 
        .Q(round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(out[178]), .CLK(clk), .RST(rst), .I(in[178]), 
        .Q(round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(out[179]), .CLK(clk), .RST(rst), .I(in[179]), 
        .Q(round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(out[180]), .CLK(clk), .RST(rst), .I(in[180]), 
        .Q(round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(out[181]), .CLK(clk), .RST(rst), .I(in[181]), 
        .Q(round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(out[182]), .CLK(clk), .RST(rst), .I(in[182]), 
        .Q(round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(out[183]), .CLK(clk), .RST(rst), .I(in[183]), 
        .Q(round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(out[184]), .CLK(clk), .RST(rst), .I(in[184]), 
        .Q(round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(out[185]), .CLK(clk), .RST(rst), .I(in[185]), 
        .Q(round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(out[186]), .CLK(clk), .RST(rst), .I(in[186]), 
        .Q(round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(out[187]), .CLK(clk), .RST(rst), .I(in[187]), 
        .Q(round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(out[188]), .CLK(clk), .RST(rst), .I(in[188]), 
        .Q(round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(out[189]), .CLK(clk), .RST(rst), .I(in[189]), 
        .Q(round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(out[190]), .CLK(clk), .RST(rst), .I(in[190]), 
        .Q(round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(out[191]), .CLK(clk), .RST(rst), .I(in[191]), 
        .Q(round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(out[192]), .CLK(clk), .RST(rst), .I(in[192]), 
        .Q(round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(out[193]), .CLK(clk), .RST(rst), .I(in[193]), 
        .Q(round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(out[194]), .CLK(clk), .RST(rst), .I(in[194]), 
        .Q(round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(out[195]), .CLK(clk), .RST(rst), .I(in[195]), 
        .Q(round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(out[196]), .CLK(clk), .RST(rst), .I(in[196]), 
        .Q(round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(out[197]), .CLK(clk), .RST(rst), .I(in[197]), 
        .Q(round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(out[198]), .CLK(clk), .RST(rst), .I(in[198]), 
        .Q(round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(out[199]), .CLK(clk), .RST(rst), .I(in[199]), 
        .Q(round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(out[200]), .CLK(clk), .RST(rst), .I(in[200]), 
        .Q(round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(out[201]), .CLK(clk), .RST(rst), .I(in[201]), 
        .Q(round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(out[202]), .CLK(clk), .RST(rst), .I(in[202]), 
        .Q(round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(out[203]), .CLK(clk), .RST(rst), .I(in[203]), 
        .Q(round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(out[204]), .CLK(clk), .RST(rst), .I(in[204]), 
        .Q(round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(out[205]), .CLK(clk), .RST(rst), .I(in[205]), 
        .Q(round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(out[206]), .CLK(clk), .RST(rst), .I(in[206]), 
        .Q(round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(out[207]), .CLK(clk), .RST(rst), .I(in[207]), 
        .Q(round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(out[208]), .CLK(clk), .RST(rst), .I(in[208]), 
        .Q(round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(out[209]), .CLK(clk), .RST(rst), .I(in[209]), 
        .Q(round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(out[210]), .CLK(clk), .RST(rst), .I(in[210]), 
        .Q(round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(out[211]), .CLK(clk), .RST(rst), .I(in[211]), 
        .Q(round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(out[212]), .CLK(clk), .RST(rst), .I(in[212]), 
        .Q(round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(out[213]), .CLK(clk), .RST(rst), .I(in[213]), 
        .Q(round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(out[214]), .CLK(clk), .RST(rst), .I(in[214]), 
        .Q(round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(out[215]), .CLK(clk), .RST(rst), .I(in[215]), 
        .Q(round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(out[216]), .CLK(clk), .RST(rst), .I(in[216]), 
        .Q(round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(out[217]), .CLK(clk), .RST(rst), .I(in[217]), 
        .Q(round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(out[218]), .CLK(clk), .RST(rst), .I(in[218]), 
        .Q(round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(out[219]), .CLK(clk), .RST(rst), .I(in[219]), 
        .Q(round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(out[220]), .CLK(clk), .RST(rst), .I(in[220]), 
        .Q(round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(out[221]), .CLK(clk), .RST(rst), .I(in[221]), 
        .Q(round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(out[222]), .CLK(clk), .RST(rst), .I(in[222]), 
        .Q(round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(out[223]), .CLK(clk), .RST(rst), .I(in[223]), 
        .Q(round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(out[224]), .CLK(clk), .RST(rst), .I(in[224]), 
        .Q(round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(out[225]), .CLK(clk), .RST(rst), .I(in[225]), 
        .Q(round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(out[226]), .CLK(clk), .RST(rst), .I(in[226]), 
        .Q(round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(out[227]), .CLK(clk), .RST(rst), .I(in[227]), 
        .Q(round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(out[228]), .CLK(clk), .RST(rst), .I(in[228]), 
        .Q(round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(out[229]), .CLK(clk), .RST(rst), .I(in[229]), 
        .Q(round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(out[230]), .CLK(clk), .RST(rst), .I(in[230]), 
        .Q(round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(out[231]), .CLK(clk), .RST(rst), .I(in[231]), 
        .Q(round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(out[232]), .CLK(clk), .RST(rst), .I(in[232]), 
        .Q(round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(out[233]), .CLK(clk), .RST(rst), .I(in[233]), 
        .Q(round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(out[234]), .CLK(clk), .RST(rst), .I(in[234]), 
        .Q(round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(out[235]), .CLK(clk), .RST(rst), .I(in[235]), 
        .Q(round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(out[236]), .CLK(clk), .RST(rst), .I(in[236]), 
        .Q(round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(out[237]), .CLK(clk), .RST(rst), .I(in[237]), 
        .Q(round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(out[238]), .CLK(clk), .RST(rst), .I(in[238]), 
        .Q(round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(out[239]), .CLK(clk), .RST(rst), .I(in[239]), 
        .Q(round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(out[240]), .CLK(clk), .RST(rst), .I(in[240]), 
        .Q(round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(out[241]), .CLK(clk), .RST(rst), .I(in[241]), 
        .Q(round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(out[242]), .CLK(clk), .RST(rst), .I(in[242]), 
        .Q(round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(out[243]), .CLK(clk), .RST(rst), .I(in[243]), 
        .Q(round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(out[244]), .CLK(clk), .RST(rst), .I(in[244]), 
        .Q(round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(out[245]), .CLK(clk), .RST(rst), .I(in[245]), 
        .Q(round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(out[246]), .CLK(clk), .RST(rst), .I(in[246]), 
        .Q(round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(out[247]), .CLK(clk), .RST(rst), .I(in[247]), 
        .Q(round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(out[248]), .CLK(clk), .RST(rst), .I(in[248]), 
        .Q(round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(out[249]), .CLK(clk), .RST(rst), .I(in[249]), 
        .Q(round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(out[250]), .CLK(clk), .RST(rst), .I(in[250]), 
        .Q(round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(out[251]), .CLK(clk), .RST(rst), .I(in[251]), 
        .Q(round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(out[252]), .CLK(clk), .RST(rst), .I(in[252]), 
        .Q(round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(out[253]), .CLK(clk), .RST(rst), .I(in[253]), 
        .Q(round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(out[254]), .CLK(clk), .RST(rst), .I(in[254]), 
        .Q(round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(out[255]), .CLK(clk), .RST(rst), .I(in[255]), 
        .Q(round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(out[256]), .CLK(clk), .RST(rst), .I(in[256]), 
        .Q(round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(out[257]), .CLK(clk), .RST(rst), .I(in[257]), 
        .Q(round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(out[258]), .CLK(clk), .RST(rst), .I(in[258]), 
        .Q(round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(out[259]), .CLK(clk), .RST(rst), .I(in[259]), 
        .Q(round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(out[260]), .CLK(clk), .RST(rst), .I(in[260]), 
        .Q(round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(out[261]), .CLK(clk), .RST(rst), .I(in[261]), 
        .Q(round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(out[262]), .CLK(clk), .RST(rst), .I(in[262]), 
        .Q(round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(out[263]), .CLK(clk), .RST(rst), .I(in[263]), 
        .Q(round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(out[264]), .CLK(clk), .RST(rst), .I(in[264]), 
        .Q(round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(out[265]), .CLK(clk), .RST(rst), .I(in[265]), 
        .Q(round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(out[266]), .CLK(clk), .RST(rst), .I(in[266]), 
        .Q(round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(out[267]), .CLK(clk), .RST(rst), .I(in[267]), 
        .Q(round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(out[268]), .CLK(clk), .RST(rst), .I(in[268]), 
        .Q(round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(out[269]), .CLK(clk), .RST(rst), .I(in[269]), 
        .Q(round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(out[270]), .CLK(clk), .RST(rst), .I(in[270]), 
        .Q(round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(out[271]), .CLK(clk), .RST(rst), .I(in[271]), 
        .Q(round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(out[272]), .CLK(clk), .RST(rst), .I(in[272]), 
        .Q(round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(out[273]), .CLK(clk), .RST(rst), .I(in[273]), 
        .Q(round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(out[274]), .CLK(clk), .RST(rst), .I(in[274]), 
        .Q(round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(out[275]), .CLK(clk), .RST(rst), .I(in[275]), 
        .Q(round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(out[276]), .CLK(clk), .RST(rst), .I(in[276]), 
        .Q(round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(out[277]), .CLK(clk), .RST(rst), .I(in[277]), 
        .Q(round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(out[278]), .CLK(clk), .RST(rst), .I(in[278]), 
        .Q(round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(out[279]), .CLK(clk), .RST(rst), .I(in[279]), 
        .Q(round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(out[280]), .CLK(clk), .RST(rst), .I(in[280]), 
        .Q(round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(out[281]), .CLK(clk), .RST(rst), .I(in[281]), 
        .Q(round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(out[282]), .CLK(clk), .RST(rst), .I(in[282]), 
        .Q(round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(out[283]), .CLK(clk), .RST(rst), .I(in[283]), 
        .Q(round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(out[284]), .CLK(clk), .RST(rst), .I(in[284]), 
        .Q(round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(out[285]), .CLK(clk), .RST(rst), .I(in[285]), 
        .Q(round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(out[286]), .CLK(clk), .RST(rst), .I(in[286]), 
        .Q(round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(out[287]), .CLK(clk), .RST(rst), .I(in[287]), 
        .Q(round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(out[288]), .CLK(clk), .RST(rst), .I(in[288]), 
        .Q(round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(out[289]), .CLK(clk), .RST(rst), .I(in[289]), 
        .Q(round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(out[290]), .CLK(clk), .RST(rst), .I(in[290]), 
        .Q(round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(out[291]), .CLK(clk), .RST(rst), .I(in[291]), 
        .Q(round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(out[292]), .CLK(clk), .RST(rst), .I(in[292]), 
        .Q(round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(out[293]), .CLK(clk), .RST(rst), .I(in[293]), 
        .Q(round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(out[294]), .CLK(clk), .RST(rst), .I(in[294]), 
        .Q(round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(out[295]), .CLK(clk), .RST(rst), .I(in[295]), 
        .Q(round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(out[296]), .CLK(clk), .RST(rst), .I(in[296]), 
        .Q(round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(out[297]), .CLK(clk), .RST(rst), .I(in[297]), 
        .Q(round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(out[298]), .CLK(clk), .RST(rst), .I(in[298]), 
        .Q(round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(out[299]), .CLK(clk), .RST(rst), .I(in[299]), 
        .Q(round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(out[300]), .CLK(clk), .RST(rst), .I(in[300]), 
        .Q(round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(out[301]), .CLK(clk), .RST(rst), .I(in[301]), 
        .Q(round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(out[302]), .CLK(clk), .RST(rst), .I(in[302]), 
        .Q(round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(out[303]), .CLK(clk), .RST(rst), .I(in[303]), 
        .Q(round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(out[304]), .CLK(clk), .RST(rst), .I(in[304]), 
        .Q(round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(out[305]), .CLK(clk), .RST(rst), .I(in[305]), 
        .Q(round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(out[306]), .CLK(clk), .RST(rst), .I(in[306]), 
        .Q(round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(out[307]), .CLK(clk), .RST(rst), .I(in[307]), 
        .Q(round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(out[308]), .CLK(clk), .RST(rst), .I(in[308]), 
        .Q(round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(out[309]), .CLK(clk), .RST(rst), .I(in[309]), 
        .Q(round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(out[310]), .CLK(clk), .RST(rst), .I(in[310]), 
        .Q(round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(out[311]), .CLK(clk), .RST(rst), .I(in[311]), 
        .Q(round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(out[312]), .CLK(clk), .RST(rst), .I(in[312]), 
        .Q(round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(out[313]), .CLK(clk), .RST(rst), .I(in[313]), 
        .Q(round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(out[314]), .CLK(clk), .RST(rst), .I(in[314]), 
        .Q(round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(out[315]), .CLK(clk), .RST(rst), .I(in[315]), 
        .Q(round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(out[316]), .CLK(clk), .RST(rst), .I(in[316]), 
        .Q(round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(out[317]), .CLK(clk), .RST(rst), .I(in[317]), 
        .Q(round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(out[318]), .CLK(clk), .RST(rst), .I(in[318]), 
        .Q(round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(out[319]), .CLK(clk), .RST(rst), .I(in[319]), 
        .Q(round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(out[320]), .CLK(clk), .RST(rst), .I(in[320]), 
        .Q(round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(out[321]), .CLK(clk), .RST(rst), .I(in[321]), 
        .Q(round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(out[322]), .CLK(clk), .RST(rst), .I(in[322]), 
        .Q(round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(out[323]), .CLK(clk), .RST(rst), .I(in[323]), 
        .Q(round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(out[324]), .CLK(clk), .RST(rst), .I(in[324]), 
        .Q(round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(out[325]), .CLK(clk), .RST(rst), .I(in[325]), 
        .Q(round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(out[326]), .CLK(clk), .RST(rst), .I(in[326]), 
        .Q(round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(out[327]), .CLK(clk), .RST(rst), .I(in[327]), 
        .Q(round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(out[328]), .CLK(clk), .RST(rst), .I(in[328]), 
        .Q(round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(out[329]), .CLK(clk), .RST(rst), .I(in[329]), 
        .Q(round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(out[330]), .CLK(clk), .RST(rst), .I(in[330]), 
        .Q(round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(out[331]), .CLK(clk), .RST(rst), .I(in[331]), 
        .Q(round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(out[332]), .CLK(clk), .RST(rst), .I(in[332]), 
        .Q(round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(out[333]), .CLK(clk), .RST(rst), .I(in[333]), 
        .Q(round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(out[334]), .CLK(clk), .RST(rst), .I(in[334]), 
        .Q(round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(out[335]), .CLK(clk), .RST(rst), .I(in[335]), 
        .Q(round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(out[336]), .CLK(clk), .RST(rst), .I(in[336]), 
        .Q(round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(out[337]), .CLK(clk), .RST(rst), .I(in[337]), 
        .Q(round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(out[338]), .CLK(clk), .RST(rst), .I(in[338]), 
        .Q(round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(out[339]), .CLK(clk), .RST(rst), .I(in[339]), 
        .Q(round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(out[340]), .CLK(clk), .RST(rst), .I(in[340]), 
        .Q(round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(out[341]), .CLK(clk), .RST(rst), .I(in[341]), 
        .Q(round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(out[342]), .CLK(clk), .RST(rst), .I(in[342]), 
        .Q(round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(out[343]), .CLK(clk), .RST(rst), .I(in[343]), 
        .Q(round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(out[344]), .CLK(clk), .RST(rst), .I(in[344]), 
        .Q(round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(out[345]), .CLK(clk), .RST(rst), .I(in[345]), 
        .Q(round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(out[346]), .CLK(clk), .RST(rst), .I(in[346]), 
        .Q(round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(out[347]), .CLK(clk), .RST(rst), .I(in[347]), 
        .Q(round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(out[348]), .CLK(clk), .RST(rst), .I(in[348]), 
        .Q(round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(out[349]), .CLK(clk), .RST(rst), .I(in[349]), 
        .Q(round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(out[350]), .CLK(clk), .RST(rst), .I(in[350]), 
        .Q(round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(out[351]), .CLK(clk), .RST(rst), .I(in[351]), 
        .Q(round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(out[352]), .CLK(clk), .RST(rst), .I(in[352]), 
        .Q(round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(out[353]), .CLK(clk), .RST(rst), .I(in[353]), 
        .Q(round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(out[354]), .CLK(clk), .RST(rst), .I(in[354]), 
        .Q(round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(out[355]), .CLK(clk), .RST(rst), .I(in[355]), 
        .Q(round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(out[356]), .CLK(clk), .RST(rst), .I(in[356]), 
        .Q(round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(out[357]), .CLK(clk), .RST(rst), .I(in[357]), 
        .Q(round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(out[358]), .CLK(clk), .RST(rst), .I(in[358]), 
        .Q(round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(out[359]), .CLK(clk), .RST(rst), .I(in[359]), 
        .Q(round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(out[360]), .CLK(clk), .RST(rst), .I(in[360]), 
        .Q(round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(out[361]), .CLK(clk), .RST(rst), .I(in[361]), 
        .Q(round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(out[362]), .CLK(clk), .RST(rst), .I(in[362]), 
        .Q(round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(out[363]), .CLK(clk), .RST(rst), .I(in[363]), 
        .Q(round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(out[364]), .CLK(clk), .RST(rst), .I(in[364]), 
        .Q(round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(out[365]), .CLK(clk), .RST(rst), .I(in[365]), 
        .Q(round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(out[366]), .CLK(clk), .RST(rst), .I(in[366]), 
        .Q(round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(out[367]), .CLK(clk), .RST(rst), .I(in[367]), 
        .Q(round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(out[368]), .CLK(clk), .RST(rst), .I(in[368]), 
        .Q(round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(out[369]), .CLK(clk), .RST(rst), .I(in[369]), 
        .Q(round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(out[370]), .CLK(clk), .RST(rst), .I(in[370]), 
        .Q(round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(out[371]), .CLK(clk), .RST(rst), .I(in[371]), 
        .Q(round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(out[372]), .CLK(clk), .RST(rst), .I(in[372]), 
        .Q(round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(out[373]), .CLK(clk), .RST(rst), .I(in[373]), 
        .Q(round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(out[374]), .CLK(clk), .RST(rst), .I(in[374]), 
        .Q(round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(out[375]), .CLK(clk), .RST(rst), .I(in[375]), 
        .Q(round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(out[376]), .CLK(clk), .RST(rst), .I(in[376]), 
        .Q(round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(out[377]), .CLK(clk), .RST(rst), .I(in[377]), 
        .Q(round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(out[378]), .CLK(clk), .RST(rst), .I(in[378]), 
        .Q(round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(out[379]), .CLK(clk), .RST(rst), .I(in[379]), 
        .Q(round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(out[380]), .CLK(clk), .RST(rst), .I(in[380]), 
        .Q(round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(out[381]), .CLK(clk), .RST(rst), .I(in[381]), 
        .Q(round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(out[382]), .CLK(clk), .RST(rst), .I(in[382]), 
        .Q(round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(out[383]), .CLK(clk), .RST(rst), .I(in[383]), 
        .Q(round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(out[384]), .CLK(clk), .RST(rst), .I(in[384]), 
        .Q(round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(out[385]), .CLK(clk), .RST(rst), .I(in[385]), 
        .Q(round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(out[386]), .CLK(clk), .RST(rst), .I(in[386]), 
        .Q(round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(out[387]), .CLK(clk), .RST(rst), .I(in[387]), 
        .Q(round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(out[388]), .CLK(clk), .RST(rst), .I(in[388]), 
        .Q(round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(out[389]), .CLK(clk), .RST(rst), .I(in[389]), 
        .Q(round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(out[390]), .CLK(clk), .RST(rst), .I(in[390]), 
        .Q(round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(out[391]), .CLK(clk), .RST(rst), .I(in[391]), 
        .Q(round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(out[392]), .CLK(clk), .RST(rst), .I(in[392]), 
        .Q(round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(out[393]), .CLK(clk), .RST(rst), .I(in[393]), 
        .Q(round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(out[394]), .CLK(clk), .RST(rst), .I(in[394]), 
        .Q(round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(out[395]), .CLK(clk), .RST(rst), .I(in[395]), 
        .Q(round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(out[396]), .CLK(clk), .RST(rst), .I(in[396]), 
        .Q(round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(out[397]), .CLK(clk), .RST(rst), .I(in[397]), 
        .Q(round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(out[398]), .CLK(clk), .RST(rst), .I(in[398]), 
        .Q(round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(out[399]), .CLK(clk), .RST(rst), .I(in[399]), 
        .Q(round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(out[400]), .CLK(clk), .RST(rst), .I(in[400]), 
        .Q(round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(out[401]), .CLK(clk), .RST(rst), .I(in[401]), 
        .Q(round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(out[402]), .CLK(clk), .RST(rst), .I(in[402]), 
        .Q(round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(out[403]), .CLK(clk), .RST(rst), .I(in[403]), 
        .Q(round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(out[404]), .CLK(clk), .RST(rst), .I(in[404]), 
        .Q(round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(out[405]), .CLK(clk), .RST(rst), .I(in[405]), 
        .Q(round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(out[406]), .CLK(clk), .RST(rst), .I(in[406]), 
        .Q(round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(out[407]), .CLK(clk), .RST(rst), .I(in[407]), 
        .Q(round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(out[408]), .CLK(clk), .RST(rst), .I(in[408]), 
        .Q(round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(out[409]), .CLK(clk), .RST(rst), .I(in[409]), 
        .Q(round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(out[410]), .CLK(clk), .RST(rst), .I(in[410]), 
        .Q(round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(out[411]), .CLK(clk), .RST(rst), .I(in[411]), 
        .Q(round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(out[412]), .CLK(clk), .RST(rst), .I(in[412]), 
        .Q(round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(out[413]), .CLK(clk), .RST(rst), .I(in[413]), 
        .Q(round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(out[414]), .CLK(clk), .RST(rst), .I(in[414]), 
        .Q(round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(out[415]), .CLK(clk), .RST(rst), .I(in[415]), 
        .Q(round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(out[416]), .CLK(clk), .RST(rst), .I(in[416]), 
        .Q(round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(out[417]), .CLK(clk), .RST(rst), .I(in[417]), 
        .Q(round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(out[418]), .CLK(clk), .RST(rst), .I(in[418]), 
        .Q(round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(out[419]), .CLK(clk), .RST(rst), .I(in[419]), 
        .Q(round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(out[420]), .CLK(clk), .RST(rst), .I(in[420]), 
        .Q(round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(out[421]), .CLK(clk), .RST(rst), .I(in[421]), 
        .Q(round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(out[422]), .CLK(clk), .RST(rst), .I(in[422]), 
        .Q(round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(out[423]), .CLK(clk), .RST(rst), .I(in[423]), 
        .Q(round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(out[424]), .CLK(clk), .RST(rst), .I(in[424]), 
        .Q(round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(out[425]), .CLK(clk), .RST(rst), .I(in[425]), 
        .Q(round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(out[426]), .CLK(clk), .RST(rst), .I(in[426]), 
        .Q(round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(out[427]), .CLK(clk), .RST(rst), .I(in[427]), 
        .Q(round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(out[428]), .CLK(clk), .RST(rst), .I(in[428]), 
        .Q(round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(out[429]), .CLK(clk), .RST(rst), .I(in[429]), 
        .Q(round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(out[430]), .CLK(clk), .RST(rst), .I(in[430]), 
        .Q(round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(out[431]), .CLK(clk), .RST(rst), .I(in[431]), 
        .Q(round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(out[432]), .CLK(clk), .RST(rst), .I(in[432]), 
        .Q(round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(out[433]), .CLK(clk), .RST(rst), .I(in[433]), 
        .Q(round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(out[434]), .CLK(clk), .RST(rst), .I(in[434]), 
        .Q(round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(out[435]), .CLK(clk), .RST(rst), .I(in[435]), 
        .Q(round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(out[436]), .CLK(clk), .RST(rst), .I(in[436]), 
        .Q(round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(out[437]), .CLK(clk), .RST(rst), .I(in[437]), 
        .Q(round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(out[438]), .CLK(clk), .RST(rst), .I(in[438]), 
        .Q(round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(out[439]), .CLK(clk), .RST(rst), .I(in[439]), 
        .Q(round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(out[440]), .CLK(clk), .RST(rst), .I(in[440]), 
        .Q(round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(out[441]), .CLK(clk), .RST(rst), .I(in[441]), 
        .Q(round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(out[442]), .CLK(clk), .RST(rst), .I(in[442]), 
        .Q(round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(out[443]), .CLK(clk), .RST(rst), .I(in[443]), 
        .Q(round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(out[444]), .CLK(clk), .RST(rst), .I(in[444]), 
        .Q(round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(out[445]), .CLK(clk), .RST(rst), .I(in[445]), 
        .Q(round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(out[446]), .CLK(clk), .RST(rst), .I(in[446]), 
        .Q(round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(out[447]), .CLK(clk), .RST(rst), .I(in[447]), 
        .Q(round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(out[448]), .CLK(clk), .RST(rst), .I(in[448]), 
        .Q(round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(out[449]), .CLK(clk), .RST(rst), .I(in[449]), 
        .Q(round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(out[450]), .CLK(clk), .RST(rst), .I(in[450]), 
        .Q(round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(out[451]), .CLK(clk), .RST(rst), .I(in[451]), 
        .Q(round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(out[452]), .CLK(clk), .RST(rst), .I(in[452]), 
        .Q(round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(out[453]), .CLK(clk), .RST(rst), .I(in[453]), 
        .Q(round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(out[454]), .CLK(clk), .RST(rst), .I(in[454]), 
        .Q(round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(out[455]), .CLK(clk), .RST(rst), .I(in[455]), 
        .Q(round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(out[456]), .CLK(clk), .RST(rst), .I(in[456]), 
        .Q(round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(out[457]), .CLK(clk), .RST(rst), .I(in[457]), 
        .Q(round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(out[458]), .CLK(clk), .RST(rst), .I(in[458]), 
        .Q(round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(out[459]), .CLK(clk), .RST(rst), .I(in[459]), 
        .Q(round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(out[460]), .CLK(clk), .RST(rst), .I(in[460]), 
        .Q(round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(out[461]), .CLK(clk), .RST(rst), .I(in[461]), 
        .Q(round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(out[462]), .CLK(clk), .RST(rst), .I(in[462]), 
        .Q(round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(out[463]), .CLK(clk), .RST(rst), .I(in[463]), 
        .Q(round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(out[464]), .CLK(clk), .RST(rst), .I(in[464]), 
        .Q(round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(out[465]), .CLK(clk), .RST(rst), .I(in[465]), 
        .Q(round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(out[466]), .CLK(clk), .RST(rst), .I(in[466]), 
        .Q(round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(out[467]), .CLK(clk), .RST(rst), .I(in[467]), 
        .Q(round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(out[468]), .CLK(clk), .RST(rst), .I(in[468]), 
        .Q(round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(out[469]), .CLK(clk), .RST(rst), .I(in[469]), 
        .Q(round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(out[470]), .CLK(clk), .RST(rst), .I(in[470]), 
        .Q(round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(out[471]), .CLK(clk), .RST(rst), .I(in[471]), 
        .Q(round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(out[472]), .CLK(clk), .RST(rst), .I(in[472]), 
        .Q(round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(out[473]), .CLK(clk), .RST(rst), .I(in[473]), 
        .Q(round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(out[474]), .CLK(clk), .RST(rst), .I(in[474]), 
        .Q(round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(out[475]), .CLK(clk), .RST(rst), .I(in[475]), 
        .Q(round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(out[476]), .CLK(clk), .RST(rst), .I(in[476]), 
        .Q(round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(out[477]), .CLK(clk), .RST(rst), .I(in[477]), 
        .Q(round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(out[478]), .CLK(clk), .RST(rst), .I(in[478]), 
        .Q(round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(out[479]), .CLK(clk), .RST(rst), .I(in[479]), 
        .Q(round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(out[480]), .CLK(clk), .RST(rst), .I(in[480]), 
        .Q(round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(out[481]), .CLK(clk), .RST(rst), .I(in[481]), 
        .Q(round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(out[482]), .CLK(clk), .RST(rst), .I(in[482]), 
        .Q(round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(out[483]), .CLK(clk), .RST(rst), .I(in[483]), 
        .Q(round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(out[484]), .CLK(clk), .RST(rst), .I(in[484]), 
        .Q(round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(out[485]), .CLK(clk), .RST(rst), .I(in[485]), 
        .Q(round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(out[486]), .CLK(clk), .RST(rst), .I(in[486]), 
        .Q(round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(out[487]), .CLK(clk), .RST(rst), .I(in[487]), 
        .Q(round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(out[488]), .CLK(clk), .RST(rst), .I(in[488]), 
        .Q(round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(out[489]), .CLK(clk), .RST(rst), .I(in[489]), 
        .Q(round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(out[490]), .CLK(clk), .RST(rst), .I(in[490]), 
        .Q(round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(out[491]), .CLK(clk), .RST(rst), .I(in[491]), 
        .Q(round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(out[492]), .CLK(clk), .RST(rst), .I(in[492]), 
        .Q(round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(out[493]), .CLK(clk), .RST(rst), .I(in[493]), 
        .Q(round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(out[494]), .CLK(clk), .RST(rst), .I(in[494]), 
        .Q(round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(out[495]), .CLK(clk), .RST(rst), .I(in[495]), 
        .Q(round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(out[496]), .CLK(clk), .RST(rst), .I(in[496]), 
        .Q(round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(out[497]), .CLK(clk), .RST(rst), .I(in[497]), 
        .Q(round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(out[498]), .CLK(clk), .RST(rst), .I(in[498]), 
        .Q(round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(out[499]), .CLK(clk), .RST(rst), .I(in[499]), 
        .Q(round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(out[500]), .CLK(clk), .RST(rst), .I(in[500]), 
        .Q(round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(out[501]), .CLK(clk), .RST(rst), .I(in[501]), 
        .Q(round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(out[502]), .CLK(clk), .RST(rst), .I(in[502]), 
        .Q(round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(out[503]), .CLK(clk), .RST(rst), .I(in[503]), 
        .Q(round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(out[504]), .CLK(clk), .RST(rst), .I(in[504]), 
        .Q(round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(out[505]), .CLK(clk), .RST(rst), .I(in[505]), 
        .Q(round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(out[506]), .CLK(clk), .RST(rst), .I(in[506]), 
        .Q(round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(out[507]), .CLK(clk), .RST(rst), .I(in[507]), 
        .Q(round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(out[508]), .CLK(clk), .RST(rst), .I(in[508]), 
        .Q(round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(out[509]), .CLK(clk), .RST(rst), .I(in[509]), 
        .Q(round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(out[510]), .CLK(clk), .RST(rst), .I(in[510]), 
        .Q(round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(out[511]), .CLK(clk), .RST(rst), .I(in[511]), 
        .Q(round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(out[512]), .CLK(clk), .RST(rst), .I(in[512]), 
        .Q(round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(out[513]), .CLK(clk), .RST(rst), .I(in[513]), 
        .Q(round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(out[514]), .CLK(clk), .RST(rst), .I(in[514]), 
        .Q(round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(out[515]), .CLK(clk), .RST(rst), .I(in[515]), 
        .Q(round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(out[516]), .CLK(clk), .RST(rst), .I(in[516]), 
        .Q(round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(out[517]), .CLK(clk), .RST(rst), .I(in[517]), 
        .Q(round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(out[518]), .CLK(clk), .RST(rst), .I(in[518]), 
        .Q(round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(out[519]), .CLK(clk), .RST(rst), .I(in[519]), 
        .Q(round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(out[520]), .CLK(clk), .RST(rst), .I(in[520]), 
        .Q(round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(out[521]), .CLK(clk), .RST(rst), .I(in[521]), 
        .Q(round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(out[522]), .CLK(clk), .RST(rst), .I(in[522]), 
        .Q(round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(out[523]), .CLK(clk), .RST(rst), .I(in[523]), 
        .Q(round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(out[524]), .CLK(clk), .RST(rst), .I(in[524]), 
        .Q(round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(out[525]), .CLK(clk), .RST(rst), .I(in[525]), 
        .Q(round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(out[526]), .CLK(clk), .RST(rst), .I(in[526]), 
        .Q(round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(out[527]), .CLK(clk), .RST(rst), .I(in[527]), 
        .Q(round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(out[528]), .CLK(clk), .RST(rst), .I(in[528]), 
        .Q(round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(out[529]), .CLK(clk), .RST(rst), .I(in[529]), 
        .Q(round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(out[530]), .CLK(clk), .RST(rst), .I(in[530]), 
        .Q(round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(out[531]), .CLK(clk), .RST(rst), .I(in[531]), 
        .Q(round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(out[532]), .CLK(clk), .RST(rst), .I(in[532]), 
        .Q(round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(out[533]), .CLK(clk), .RST(rst), .I(in[533]), 
        .Q(round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(out[534]), .CLK(clk), .RST(rst), .I(in[534]), 
        .Q(round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(out[535]), .CLK(clk), .RST(rst), .I(in[535]), 
        .Q(round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(out[536]), .CLK(clk), .RST(rst), .I(in[536]), 
        .Q(round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(out[537]), .CLK(clk), .RST(rst), .I(in[537]), 
        .Q(round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(out[538]), .CLK(clk), .RST(rst), .I(in[538]), 
        .Q(round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(out[539]), .CLK(clk), .RST(rst), .I(in[539]), 
        .Q(round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(out[540]), .CLK(clk), .RST(rst), .I(in[540]), 
        .Q(round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(out[541]), .CLK(clk), .RST(rst), .I(in[541]), 
        .Q(round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(out[542]), .CLK(clk), .RST(rst), .I(in[542]), 
        .Q(round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(out[543]), .CLK(clk), .RST(rst), .I(in[543]), 
        .Q(round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(out[544]), .CLK(clk), .RST(rst), .I(in[544]), 
        .Q(round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(out[545]), .CLK(clk), .RST(rst), .I(in[545]), 
        .Q(round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(out[546]), .CLK(clk), .RST(rst), .I(in[546]), 
        .Q(round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(out[547]), .CLK(clk), .RST(rst), .I(in[547]), 
        .Q(round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(out[548]), .CLK(clk), .RST(rst), .I(in[548]), 
        .Q(round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(out[549]), .CLK(clk), .RST(rst), .I(in[549]), 
        .Q(round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(out[550]), .CLK(clk), .RST(rst), .I(in[550]), 
        .Q(round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(out[551]), .CLK(clk), .RST(rst), .I(in[551]), 
        .Q(round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(out[552]), .CLK(clk), .RST(rst), .I(in[552]), 
        .Q(round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(out[553]), .CLK(clk), .RST(rst), .I(in[553]), 
        .Q(round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(out[554]), .CLK(clk), .RST(rst), .I(in[554]), 
        .Q(round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(out[555]), .CLK(clk), .RST(rst), .I(in[555]), 
        .Q(round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(out[556]), .CLK(clk), .RST(rst), .I(in[556]), 
        .Q(round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(out[557]), .CLK(clk), .RST(rst), .I(in[557]), 
        .Q(round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(out[558]), .CLK(clk), .RST(rst), .I(in[558]), 
        .Q(round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(out[559]), .CLK(clk), .RST(rst), .I(in[559]), 
        .Q(round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(out[560]), .CLK(clk), .RST(rst), .I(in[560]), 
        .Q(round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(out[561]), .CLK(clk), .RST(rst), .I(in[561]), 
        .Q(round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(out[562]), .CLK(clk), .RST(rst), .I(in[562]), 
        .Q(round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(out[563]), .CLK(clk), .RST(rst), .I(in[563]), 
        .Q(round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(out[564]), .CLK(clk), .RST(rst), .I(in[564]), 
        .Q(round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(out[565]), .CLK(clk), .RST(rst), .I(in[565]), 
        .Q(round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(out[566]), .CLK(clk), .RST(rst), .I(in[566]), 
        .Q(round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(out[567]), .CLK(clk), .RST(rst), .I(in[567]), 
        .Q(round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(out[568]), .CLK(clk), .RST(rst), .I(in[568]), 
        .Q(round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(out[569]), .CLK(clk), .RST(rst), .I(in[569]), 
        .Q(round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(out[570]), .CLK(clk), .RST(rst), .I(in[570]), 
        .Q(round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(out[571]), .CLK(clk), .RST(rst), .I(in[571]), 
        .Q(round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(out[572]), .CLK(clk), .RST(rst), .I(in[572]), 
        .Q(round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(out[573]), .CLK(clk), .RST(rst), .I(in[573]), 
        .Q(round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(out[574]), .CLK(clk), .RST(rst), .I(in[574]), 
        .Q(round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(out[575]), .CLK(clk), .RST(rst), .I(in[575]), 
        .Q(round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(out[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(out[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(out[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(out[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(out[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(out[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(out[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(out[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(out[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(out[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(out[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(out[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(out[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(out[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(out[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(out[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(out[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(out[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(out[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(out[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(out[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(out[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(out[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(out[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(out[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(out[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(out[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(out[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(out[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(out[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(out[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(out[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(out[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(out[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(out[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(out[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(out[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(out[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(out[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(out[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(out[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(out[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(out[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(out[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(out[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(out[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(out[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(out[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(out[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(out[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(out[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(out[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(out[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(out[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(out[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(out[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(out[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(out[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(out[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(out[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(out[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(out[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(out[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(out[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(out[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(out[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(out[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(out[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(out[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(out[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(out[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(out[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(out[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(out[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(out[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(out[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(out[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(out[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(out[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(out[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(out[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(out[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(out[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(out[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(out[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(out[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(out[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(out[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(out[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(out[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(out[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(out[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(out[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(out[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(out[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(out[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(out[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(out[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(out[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(out[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(out[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(out[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(out[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(out[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(out[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(out[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(out[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(out[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(out[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(out[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(out[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(out[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(out[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(out[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(out[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(out[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(out[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(out[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(out[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(out[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(out[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(out[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(out[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(out[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(out[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(out[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(out[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(out[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(out[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(out[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(out[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(out[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(out[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(out[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(out[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(out[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(out[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(out[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(out[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(out[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(out[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(out[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(out[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(out[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(out[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(out[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(out[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(out[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(out[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(out[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(out[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(out[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(out[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(out[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(out[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(out[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(out[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(out[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(out[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(out[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(out[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(out[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(out[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(out[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(out[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(out[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(out[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(out[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(out[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(out[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(out[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(out[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(out[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(out[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(out[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(out[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(out[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(out[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(out[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(out[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(out[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(out[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(out[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(out[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(out[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(out[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(out[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(out[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(out[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(out[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(out[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(out[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(out[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(out[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(out[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(out[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(out[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(out[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(out[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(out[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(out[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(out[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(out[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(out[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(out[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(out[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(out[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(out[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(out[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(out[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(out[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(out[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(out[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(out[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(out[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(out[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(out[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(out[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(out[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(out[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(out[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(out[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(out[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(out[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(out[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(out[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(out[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(out[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(out[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(out[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(out[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(out[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(out[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(out[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(out[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(out[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(out[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(out[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(out[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(out[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(out[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(out[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(out[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(out[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(out[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(out[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(out[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(out[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(out[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(out[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(out[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(out[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(out[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(out[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(out[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(out[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(out[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(out[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(out[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(out[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(out[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(out[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(out[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(out[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(out[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(out[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(out[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(out[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(out[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(out[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(out[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(out[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(out[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(out[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(out[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(out[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(out[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(out[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(out[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(out[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(out[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(out[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(out[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(out[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(out[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(out[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(out[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(out[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(out[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(out[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(out[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(out[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(out[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(out[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(out[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(out[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(out[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(out[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(out[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(out[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(out[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(out[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(out[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(out[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(out[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(out[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(out[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(out[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(out[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(out[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(out[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(out[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(out[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(out[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(out[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(out[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(out[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(out[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(out[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(out[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(out[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(out[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(out[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(out[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(out[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(out[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(out[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(out[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(out[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(out[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(out[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(out[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(out[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(out[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(out[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(out[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(out[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(out[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(out[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(out[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(out[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(out[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(out[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(out[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(out[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(out[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(out[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(out[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(out[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(out[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(out[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(out[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(out[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(out[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(out[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(out[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(out[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(out[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(out[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(out[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(out[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(out[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(out[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(out[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(out[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(out[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(out[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(out[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(out[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(out[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(out[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(out[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(out[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(out[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(out[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(out[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(out[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(out[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(out[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(out[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(out[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(out[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(out[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(out[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(out[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(out[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(out[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(out[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(out[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(out[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(out[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(out[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(out[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(out[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(out[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(out[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(out[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(out[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(out[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(out[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(out[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(out[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(out[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(out[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(out[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(out[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(out[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(out[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(out[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(out[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(out[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(out[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(out[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(out[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(out[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(out[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(out[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(out[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(out[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(out[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(out[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(out[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(out[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(out[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(out[1000]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(out[1001]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(out[1002]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(out[1003]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(out[1004]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(out[1005]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(out[1006]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(out[1007]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(out[1008]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(out[1009]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(out[1010]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(out[1011]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(out[1012]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(out[1013]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(out[1014]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(out[1015]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(out[1016]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(out[1017]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(out[1018]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(out[1019]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(out[1020]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(out[1021]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(out[1022]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(out[1023]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(out[1024]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(out[1025]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(out[1026]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(out[1027]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(out[1028]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(out[1029]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(out[1030]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(out[1031]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(out[1032]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(out[1033]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(out[1034]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(out[1035]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(out[1036]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(out[1037]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(out[1038]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(out[1039]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(out[1040]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(out[1041]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(out[1042]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(out[1043]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(out[1044]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(out[1045]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(out[1046]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(out[1047]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(out[1048]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(out[1049]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(out[1050]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(out[1051]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(out[1052]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(out[1053]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(out[1054]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(out[1055]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(out[1056]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(out[1057]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(out[1058]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(out[1059]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(out[1060]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(out[1061]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(out[1062]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(out[1063]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(out[1064]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(out[1065]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(out[1066]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(out[1067]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(out[1068]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(out[1069]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(out[1070]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(out[1071]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(out[1072]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(out[1073]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(out[1074]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(out[1075]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(out[1076]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(out[1077]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(out[1078]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(out[1079]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(out[1080]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(out[1081]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(out[1082]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(out[1083]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(out[1084]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(out[1085]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(out[1086]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(out[1087]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(out[1088]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(out[1089]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(out[1090]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(out[1091]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(out[1092]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(out[1093]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(out[1094]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(out[1095]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(out[1096]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(out[1097]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(out[1098]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(out[1099]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(out[1100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(out[1101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(out[1102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(out[1103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(out[1104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(out[1105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(out[1106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(out[1107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(out[1108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(out[1109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(out[1110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(out[1111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(out[1112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(out[1113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(out[1114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(out[1115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(out[1116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(out[1117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(out[1118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(out[1119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(out[1120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(out[1121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(out[1122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(out[1123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(out[1124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(out[1125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(out[1126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(out[1127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(out[1128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(out[1129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(out[1130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(out[1131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(out[1132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(out[1133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(out[1134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(out[1135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(out[1136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(out[1137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(out[1138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(out[1139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(out[1140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(out[1141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(out[1142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(out[1143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(out[1144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(out[1145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(out[1146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(out[1147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(out[1148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(out[1149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(out[1150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(out[1151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(out[1152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(out[1153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(out[1154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(out[1155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(out[1156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(out[1157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(out[1158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(out[1159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(out[1160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(out[1161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(out[1162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(out[1163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(out[1164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(out[1165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(out[1166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(out[1167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(out[1168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(out[1169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(out[1170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(out[1171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(out[1172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(out[1173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(out[1174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(out[1175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(out[1176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(out[1177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(out[1178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(out[1179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(out[1180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(out[1181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(out[1182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(out[1183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(out[1184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(out[1185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(out[1186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(out[1187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(out[1188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(out[1189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(out[1190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(out[1191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(out[1192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(out[1193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(out[1194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(out[1195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(out[1196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(out[1197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(out[1198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(out[1199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(out[1200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(out[1201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(out[1202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(out[1203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(out[1204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(out[1205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(out[1206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(out[1207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(out[1208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(out[1209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(out[1210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(out[1211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(out[1212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(out[1213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(out[1214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(out[1215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(out[1216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(out[1217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(out[1218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(out[1219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(out[1220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(out[1221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(out[1222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(out[1223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(out[1224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(out[1225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(out[1226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(out[1227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(out[1228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(out[1229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(out[1230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(out[1231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(out[1232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(out[1233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(out[1234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(out[1235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(out[1236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(out[1237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(out[1238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(out[1239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(out[1240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(out[1241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(out[1242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(out[1243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(out[1244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(out[1245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(out[1246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(out[1247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(out[1248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(out[1249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(out[1250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(out[1251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(out[1252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(out[1253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(out[1254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(out[1255]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(out[1256]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(out[1257]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(out[1258]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(out[1259]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(out[1260]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(out[1261]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(out[1262]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(out[1263]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(out[1264]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(out[1265]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(out[1266]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(out[1267]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(out[1268]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(out[1269]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(out[1270]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(out[1271]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(out[1272]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(out[1273]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(out[1274]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(out[1275]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(out[1276]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(out[1277]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(out[1278]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(out[1279]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(out[1280]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(out[1281]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(out[1282]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(out[1283]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(out[1284]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(out[1285]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(out[1286]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(out[1287]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(out[1288]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(out[1289]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(out[1290]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(out[1291]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(out[1292]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(out[1293]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(out[1294]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(out[1295]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(out[1296]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(out[1297]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(out[1298]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(out[1299]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(out[1300]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(out[1301]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(out[1302]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(out[1303]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(out[1304]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(out[1305]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(out[1306]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(out[1307]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(out[1308]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(out[1309]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(out[1310]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(out[1311]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(out[1312]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(out[1313]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(out[1314]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(out[1315]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(out[1316]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(out[1317]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(out[1318]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(out[1319]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(out[1320]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(out[1321]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(out[1322]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(out[1323]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(out[1324]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(out[1325]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(out[1326]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(out[1327]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(out[1328]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(out[1329]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(out[1330]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(out[1331]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(out[1332]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(out[1333]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(out[1334]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(out[1335]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(out[1336]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(out[1337]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(out[1338]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(out[1339]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(out[1340]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(out[1341]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(out[1342]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(out[1343]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(out[1344]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(out[1345]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(out[1346]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(out[1347]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(out[1348]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(out[1349]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(out[1350]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(out[1351]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(out[1352]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(out[1353]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(out[1354]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(out[1355]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(out[1356]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(out[1357]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(out[1358]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(out[1359]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(out[1360]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(out[1361]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(out[1362]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(out[1363]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(out[1364]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(out[1365]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(out[1366]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(out[1367]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(out[1368]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(out[1369]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(out[1370]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(out[1371]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(out[1372]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(out[1373]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(out[1374]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(out[1375]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(out[1376]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(out[1377]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(out[1378]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(out[1379]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(out[1380]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(out[1381]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(out[1382]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(out[1383]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(out[1384]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(out[1385]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(out[1386]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(out[1387]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(out[1388]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(out[1389]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(out[1390]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(out[1391]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(out[1392]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(out[1393]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(out[1394]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(out[1395]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(out[1396]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(out[1397]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(out[1398]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(out[1399]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(out[1400]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(out[1401]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(out[1402]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(out[1403]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(out[1404]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(out[1405]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(out[1406]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(out[1407]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(out[1408]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(out[1409]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(out[1410]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(out[1411]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(out[1412]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(out[1413]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(out[1414]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(out[1415]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(out[1416]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(out[1417]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(out[1418]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(out[1419]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(out[1420]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(out[1421]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(out[1422]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(out[1423]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(out[1424]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(out[1425]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(out[1426]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(out[1427]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(out[1428]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(out[1429]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(out[1430]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(out[1431]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(out[1432]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(out[1433]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(out[1434]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(out[1435]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(out[1436]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(out[1437]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(out[1438]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(out[1439]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(out[1440]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(out[1441]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(out[1442]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(out[1443]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(out[1444]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(out[1445]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(out[1446]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(out[1447]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(out[1448]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(out[1449]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(out[1450]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(out[1451]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(out[1452]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(out[1453]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(out[1454]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(out[1455]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(out[1456]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(out[1457]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(out[1458]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(out[1459]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(out[1460]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(out[1461]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(out[1462]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(out[1463]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(out[1464]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(out[1465]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(out[1466]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(out[1467]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(out[1468]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(out[1469]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(out[1470]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(out[1471]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(out[1472]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(out[1473]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(out[1474]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(out[1475]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(out[1476]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(out[1477]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(out[1478]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(out[1479]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(out[1480]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(out[1481]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(out[1482]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(out[1483]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(out[1484]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(out[1485]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(out[1486]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(out[1487]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(out[1488]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(out[1489]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(out[1490]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(out[1491]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(out[1492]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(out[1493]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(out[1494]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(out[1495]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(out[1496]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(out[1497]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(out[1498]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(out[1499]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(out[1500]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(out[1501]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(out[1502]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(out[1503]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(out[1504]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(out[1505]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(out[1506]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(out[1507]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(out[1508]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(out[1509]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(out[1510]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(out[1511]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(out[1512]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(out[1513]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(out[1514]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(out[1515]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(out[1516]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(out[1517]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(out[1518]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(out[1519]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(out[1520]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(out[1521]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(out[1522]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(out[1523]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(out[1524]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(out[1525]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(out[1526]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(out[1527]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(out[1528]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(out[1529]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(out[1530]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(out[1531]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(out[1532]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(out[1533]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(out[1534]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(out[1535]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(out[1536]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(out[1537]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(out[1538]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(out[1539]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(out[1540]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(out[1541]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(out[1542]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(out[1543]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(out[1544]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(out[1545]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(out[1546]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(out[1547]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(out[1548]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(out[1549]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(out[1550]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(out[1551]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(out[1552]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(out[1553]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(out[1554]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(out[1555]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(out[1556]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(out[1557]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(out[1558]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(out[1559]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(out[1560]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(out[1561]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(out[1562]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(out[1563]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(out[1564]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(out[1565]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(out[1566]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(out[1567]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(out[1568]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(out[1569]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(out[1570]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(out[1571]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(out[1572]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(out[1573]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(out[1574]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(out[1575]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(out[1576]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(out[1577]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(out[1578]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(out[1579]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(out[1580]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(out[1581]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(out[1582]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(out[1583]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(out[1584]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(out[1585]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(out[1586]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(out[1587]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(out[1588]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(out[1589]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(out[1590]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(out[1591]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(out[1592]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(out[1593]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(out[1594]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(out[1595]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(out[1596]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(out[1597]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(out[1598]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(out[1599]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(round_reg[1599]) );
  XNOR U1053 ( .A(n4998), .B(n5049), .Z(n4243) );
  ANDN U1054 ( .B(n3786), .A(n3787), .Z(n3784) );
  ANDN U1055 ( .B(n3790), .A(n3791), .Z(n3788) );
  ANDN U1056 ( .B(n4123), .A(n3981), .Z(n4122) );
  ANDN U1057 ( .B(n4136), .A(n3990), .Z(n4135) );
  ANDN U1058 ( .B(n3626), .A(n4081), .Z(n4217) );
  ANDN U1059 ( .B(n3680), .A(n4109), .Z(n4237) );
  ANDN U1060 ( .B(n1556), .A(n1290), .Z(n1555) );
  ANDN U1061 ( .B(n1583), .A(n1338), .Z(n1582) );
  ANDN U1062 ( .B(n1585), .A(n1342), .Z(n1584) );
  ANDN U1063 ( .B(n1587), .A(n1346), .Z(n1586) );
  ANDN U1064 ( .B(n4121), .A(n3978), .Z(n4120) );
  ANDN U1065 ( .B(n1520), .A(n1238), .Z(n1519) );
  ANDN U1066 ( .B(n1522), .A(n1242), .Z(n1521) );
  ANDN U1067 ( .B(n1524), .A(n1246), .Z(n1523) );
  ANDN U1068 ( .B(n1558), .A(n1294), .Z(n1557) );
  ANDN U1069 ( .B(n1581), .A(n1334), .Z(n1580) );
  ANDN U1070 ( .B(n1593), .A(n1350), .Z(n1592) );
  ANDN U1071 ( .B(n1710), .A(n1518), .Z(n1709) );
  ANDN U1072 ( .B(n1757), .A(n1556), .Z(n1755) );
  ANDN U1073 ( .B(n1794), .A(n1583), .Z(n1792) );
  ANDN U1074 ( .B(n1797), .A(n1585), .Z(n1795) );
  ANDN U1075 ( .B(n1800), .A(n1587), .Z(n1798) );
  XNOR U1076 ( .A(n4795), .B(n4794), .Z(n4401) );
  XOR U1077 ( .A(n4922), .B(n5398), .Z(n1930) );
  XOR U1078 ( .A(n4939), .B(n5495), .Z(n1722) );
  ANDN U1079 ( .B(n3782), .A(n3783), .Z(n3780) );
  ANDN U1080 ( .B(n3794), .A(n3795), .Z(n3792) );
  ANDN U1081 ( .B(n3798), .A(n3799), .Z(n3796) );
  ANDN U1082 ( .B(n3993), .A(n3727), .Z(n3992) );
  ANDN U1083 ( .B(n3675), .A(n4107), .Z(n4236) );
  ANDN U1084 ( .B(n4436), .A(n4437), .Z(n4434) );
  ANDN U1085 ( .B(n1579), .A(n1330), .Z(n1578) );
  ANDN U1086 ( .B(n1706), .A(n1510), .Z(n1705) );
  ANDN U1087 ( .B(n1713), .A(n1520), .Z(n1711) );
  ANDN U1088 ( .B(n1791), .A(n1581), .Z(n1789) );
  ANDN U1089 ( .B(n1803), .A(n1593), .Z(n1801) );
  ANDN U1090 ( .B(n1934), .A(n1710), .Z(n1932) );
  NOR U1091 ( .A(n1757), .B(n1288), .Z(n1972) );
  NOR U1092 ( .A(n1760), .B(n1292), .Z(n1974) );
  ANDN U1093 ( .B(n2829), .A(n2638), .Z(n2828) );
  ANDN U1094 ( .B(n2994), .A(n2835), .Z(n2992) );
  ANDN U1095 ( .B(n2996), .A(n2837), .Z(n2995) );
  ANDN U1096 ( .B(n2998), .A(n2840), .Z(n2997) );
  XNOR U1097 ( .A(n4787), .B(n4786), .Z(n4397) );
  XNOR U1098 ( .A(n4791), .B(n4790), .Z(n4399) );
  XOR U1099 ( .A(n4906), .B(n5339), .Z(n1914) );
  XOR U1100 ( .A(n5527), .B(n5526), .Z(n2243) );
  XOR U1101 ( .A(n5542), .B(n5541), .Z(n2247) );
  XOR U1102 ( .A(n5557), .B(n5556), .Z(n2251) );
  XOR U1103 ( .A(n5572), .B(n5571), .Z(n2255) );
  XOR U1104 ( .A(n5587), .B(n5586), .Z(n2263) );
  XOR U1105 ( .A(n4928), .B(n5411), .Z(n1933) );
  XOR U1106 ( .A(n4932), .B(n5424), .Z(n1712) );
  XOR U1107 ( .A(n4936), .B(n5437), .Z(n1715) );
  XOR U1108 ( .A(n4942), .B(n5654), .Z(n1725) );
  XOR U1109 ( .A(n4970), .B(n5601), .Z(n1756) );
  ANDN U1110 ( .B(n3648), .A(n3649), .Z(n3646) );
  ANDN U1111 ( .B(n3697), .A(n3698), .Z(n3695) );
  ANDN U1112 ( .B(n4432), .A(n4433), .Z(n4430) );
  ANDN U1113 ( .B(n4440), .A(n4441), .Z(n4438) );
  ANDN U1114 ( .B(n4470), .A(n4471), .Z(n4468) );
  ANDN U1115 ( .B(n4474), .A(n4475), .Z(n4472) );
  ANDN U1116 ( .B(n1560), .A(n1298), .Z(n1559) );
  ANDN U1117 ( .B(n1562), .A(n1302), .Z(n1561) );
  ANDN U1118 ( .B(n1568), .A(n1306), .Z(n1567) );
  ANDN U1119 ( .B(n1570), .A(n1310), .Z(n1569) );
  ANDN U1120 ( .B(n1702), .A(n1494), .Z(n1701) );
  ANDN U1121 ( .B(n1704), .A(n1506), .Z(n1703) );
  ANDN U1122 ( .B(n1708), .A(n1514), .Z(n1707) );
  ANDN U1123 ( .B(n1723), .A(n1524), .Z(n1721) );
  ANDN U1124 ( .B(n1784), .A(n1579), .Z(n1782) );
  ANDN U1125 ( .B(n1909), .A(n1694), .Z(n1907) );
  NOR U1126 ( .A(n1791), .B(n1332), .Z(n2003) );
  NOR U1127 ( .A(n1797), .B(n1340), .Z(n2007) );
  NOR U1128 ( .A(n1800), .B(n1344), .Z(n2009) );
  NOR U1129 ( .A(n1803), .B(n1348), .Z(n2011) );
  ANDN U1130 ( .B(n2804), .A(n2594), .Z(n2803) );
  ANDN U1131 ( .B(n2991), .A(n2829), .Z(n2989) );
  ANDN U1132 ( .B(n3001), .A(n2843), .Z(n2999) );
  NOR U1133 ( .A(n2994), .B(n2640), .Z(n3125) );
  NOR U1134 ( .A(n2996), .B(n2644), .Z(n3126) );
  NOR U1135 ( .A(n2998), .B(n2648), .Z(n3131) );
  XNOR U1136 ( .A(n4783), .B(n4782), .Z(n4395) );
  XOR U1137 ( .A(n4910), .B(n5361), .Z(n1917) );
  XOR U1138 ( .A(n4914), .B(n5372), .Z(n1920) );
  XOR U1139 ( .A(n4918), .B(n5385), .Z(n1923) );
  ANDN U1140 ( .B(n3599), .A(n3600), .Z(n3588) );
  ANDN U1141 ( .B(n3778), .A(n3779), .Z(n3776) );
  ANDN U1142 ( .B(n3802), .A(n3803), .Z(n3800) );
  ANDN U1143 ( .B(n3819), .A(n3820), .Z(n3806) );
  ANDN U1144 ( .B(n3823), .A(n3824), .Z(n3821) );
  ANDN U1145 ( .B(n3828), .A(n3829), .Z(n3826) );
  ANDN U1146 ( .B(n3832), .A(n3833), .Z(n3830) );
  ANDN U1147 ( .B(n3836), .A(n3837), .Z(n3834) );
  ANDN U1148 ( .B(n3840), .A(n3841), .Z(n3838) );
  ANDN U1149 ( .B(n3844), .A(n3845), .Z(n3842) );
  ANDN U1150 ( .B(n3848), .A(n3849), .Z(n3846) );
  ANDN U1151 ( .B(n3868), .A(n3869), .Z(n3866) );
  ANDN U1152 ( .B(n3872), .A(n3873), .Z(n3870) );
  ANDN U1153 ( .B(n3876), .A(n3877), .Z(n3874) );
  ANDN U1154 ( .B(n3894), .A(n3895), .Z(n3881) );
  ANDN U1155 ( .B(n3898), .A(n3899), .Z(n3896) );
  ANDN U1156 ( .B(n3923), .A(n3924), .Z(n3915) );
  ANDN U1157 ( .B(n3622), .A(n4079), .Z(n4216) );
  ANDN U1158 ( .B(n4424), .A(n4425), .Z(n4422) );
  ANDN U1159 ( .B(n4428), .A(n4429), .Z(n4426) );
  ANDN U1160 ( .B(n4478), .A(n4479), .Z(n4476) );
  ANDN U1161 ( .B(n4486), .A(n4487), .Z(n4484) );
  ANDN U1162 ( .B(n4492), .A(n4493), .Z(n4490) );
  ANDN U1163 ( .B(n4496), .A(n4497), .Z(n4494) );
  ANDN U1164 ( .B(n1526), .A(n1250), .Z(n1525) );
  ANDN U1165 ( .B(n1572), .A(n1314), .Z(n1571) );
  ANDN U1166 ( .B(n1574), .A(n1318), .Z(n1573) );
  ANDN U1167 ( .B(n1700), .A(n1490), .Z(n1699) );
  ANDN U1168 ( .B(n1716), .A(n1522), .Z(n1714) );
  ANDN U1169 ( .B(n1760), .A(n1558), .Z(n1758) );
  ANDN U1170 ( .B(n1244), .A(n1723), .Z(n1939) );
  NOR U1171 ( .A(n1794), .B(n1336), .Z(n2005) );
  ANDN U1172 ( .B(n2676), .A(n2395), .Z(n2675) );
  ANDN U1173 ( .B(n2678), .A(n2399), .Z(n2677) );
  ANDN U1174 ( .B(n2680), .A(n2403), .Z(n2679) );
  ANDN U1175 ( .B(n2682), .A(n2407), .Z(n2681) );
  ANDN U1176 ( .B(n2684), .A(n2411), .Z(n2683) );
  ANDN U1177 ( .B(n2692), .A(n2419), .Z(n2691) );
  ANDN U1178 ( .B(n2694), .A(n2423), .Z(n2693) );
  ANDN U1179 ( .B(n2788), .A(n2555), .Z(n2787) );
  ANDN U1180 ( .B(n2790), .A(n2559), .Z(n2789) );
  ANDN U1181 ( .B(n2792), .A(n2563), .Z(n2791) );
  ANDN U1182 ( .B(n2794), .A(n2574), .Z(n2793) );
  ANDN U1183 ( .B(n2798), .A(n2582), .Z(n2797) );
  ANDN U1184 ( .B(n2800), .A(n2586), .Z(n2799) );
  ANDN U1185 ( .B(n2802), .A(n2590), .Z(n2801) );
  ANDN U1186 ( .B(n2819), .A(n2618), .Z(n2818) );
  ANDN U1187 ( .B(n2821), .A(n2622), .Z(n2820) );
  ANDN U1188 ( .B(n2835), .A(n2642), .Z(n2834) );
  ANDN U1189 ( .B(n2847), .A(n2666), .Z(n2846) );
  ANDN U1190 ( .B(n2849), .A(n2670), .Z(n2848) );
  ANDN U1191 ( .B(n2851), .A(n2674), .Z(n2850) );
  NOR U1192 ( .A(n2930), .B(n2529), .Z(n3071) );
  NOR U1193 ( .A(n2936), .B(n2533), .Z(n3072) );
  NOR U1194 ( .A(n2938), .B(n2537), .Z(n3073) );
  NOR U1195 ( .A(n2966), .B(n2592), .Z(n3099) );
  NOR U1196 ( .A(n2991), .B(n2636), .Z(n3124) );
  NOR U1197 ( .A(n3001), .B(n2652), .Z(n3132) );
  ANDN U1198 ( .B(n3401), .A(n2122), .Z(n3400) );
  ANDN U1199 ( .B(n3403), .A(n2565), .Z(n3402) );
  ANDN U1200 ( .B(n3405), .A(n2881), .Z(n3404) );
  ANDN U1201 ( .B(n3417), .A(n3418), .Z(n3415) );
  NOR U1202 ( .A(n3395), .B(n2046), .Z(n3516) );
  XNOR U1203 ( .A(n5260), .B(n4935), .Z(n2206) );
  XOR U1204 ( .A(n4751), .B(n4750), .Z(n2086) );
  XOR U1205 ( .A(n4973), .B(n5616), .Z(n1759) );
  XOR U1206 ( .A(n4976), .B(n5631), .Z(n1762) );
  XOR U1207 ( .A(n4979), .B(n5657), .Z(n1765) );
  XOR U1208 ( .A(n4982), .B(n5672), .Z(n1768) );
  XOR U1209 ( .A(n4985), .B(n5687), .Z(n1771) );
  XOR U1210 ( .A(n4988), .B(n5702), .Z(n1774) );
  XOR U1211 ( .A(n4992), .B(n5717), .Z(n1777) );
  ANDN U1212 ( .B(n3693), .A(n3694), .Z(n3691) );
  ANDN U1213 ( .B(n3765), .A(n3766), .Z(n3763) );
  ANDN U1214 ( .B(n3769), .A(n3770), .Z(n3767) );
  ANDN U1215 ( .B(n3774), .A(n3775), .Z(n3772) );
  ANDN U1216 ( .B(n3864), .A(n3865), .Z(n3852) );
  ANDN U1217 ( .B(n3911), .A(n3912), .Z(n3902) );
  ANDN U1218 ( .B(n4416), .A(n4417), .Z(n4414) );
  ANDN U1219 ( .B(n4420), .A(n4421), .Z(n4418) );
  ANDN U1220 ( .B(n4482), .A(n4483), .Z(n4480) );
  ANDN U1221 ( .B(n4500), .A(n4501), .Z(n4498) );
  ANDN U1222 ( .B(n4504), .A(n4505), .Z(n4502) );
  NOR U1223 ( .A(n1784), .B(n1328), .Z(n2001) );
  ANDN U1224 ( .B(n2686), .A(n2415), .Z(n2685) );
  ANDN U1225 ( .B(n2739), .A(n2487), .Z(n2738) );
  ANDN U1226 ( .B(n2741), .A(n2491), .Z(n2740) );
  ANDN U1227 ( .B(n2743), .A(n2495), .Z(n2742) );
  ANDN U1228 ( .B(n2745), .A(n2499), .Z(n2744) );
  ANDN U1229 ( .B(n2747), .A(n2503), .Z(n2746) );
  ANDN U1230 ( .B(n2780), .A(n2547), .Z(n2779) );
  ANDN U1231 ( .B(n2786), .A(n2551), .Z(n2785) );
  ANDN U1232 ( .B(n2796), .A(n2578), .Z(n2795) );
  ANDN U1233 ( .B(n2813), .A(n2602), .Z(n2812) );
  ANDN U1234 ( .B(n2815), .A(n2606), .Z(n2814) );
  ANDN U1235 ( .B(n2817), .A(n2610), .Z(n2816) );
  ANDN U1236 ( .B(n2823), .A(n2626), .Z(n2822) );
  ANDN U1237 ( .B(n2825), .A(n2630), .Z(n2824) );
  ANDN U1238 ( .B(n2827), .A(n2634), .Z(n2826) );
  ANDN U1239 ( .B(n2843), .A(n2654), .Z(n2842) );
  ANDN U1240 ( .B(n2845), .A(n2662), .Z(n2844) );
  NOR U1241 ( .A(n2922), .B(n2509), .Z(n3063) );
  NOR U1242 ( .A(n2924), .B(n2513), .Z(n3068) );
  NOR U1243 ( .A(n2926), .B(n2517), .Z(n3069) );
  NOR U1244 ( .A(n2928), .B(n2525), .Z(n3070) );
  ANDN U1245 ( .B(n3320), .A(n3321), .Z(n3318) );
  ANDN U1246 ( .B(n3324), .A(n3325), .Z(n3322) );
  ANDN U1247 ( .B(n3408), .A(n3105), .Z(n3407) );
  ANDN U1248 ( .B(n3413), .A(n3414), .Z(n3411) );
  NOR U1249 ( .A(n3311), .B(n1232), .Z(n3483) );
  NOR U1250 ( .A(n3313), .B(n1276), .Z(n3484) );
  NOR U1251 ( .A(n3315), .B(n1320), .Z(n3485) );
  NOR U1252 ( .A(n3317), .B(n1364), .Z(n3486) );
  NOR U1253 ( .A(n3358), .B(n1718), .Z(n3497) );
  NOR U1254 ( .A(n3362), .B(n1752), .Z(n3499) );
  NOR U1255 ( .A(n3398), .B(n2068), .Z(n3519) );
  NOR U1256 ( .A(n3401), .B(n2090), .Z(n3520) );
  NOR U1257 ( .A(n3403), .B(n2125), .Z(n3521) );
  NOR U1258 ( .A(n3405), .B(n2169), .Z(n3522) );
  NOR U1259 ( .A(n3433), .B(n2656), .Z(n3541) );
  NOR U1260 ( .A(n3435), .B(n2688), .Z(n3542) );
  NOR U1261 ( .A(n3437), .B(n2720), .Z(n3543) );
  NOR U1262 ( .A(n3439), .B(n2749), .Z(n3544) );
  NOR U1263 ( .A(n3441), .B(n2782), .Z(n3545) );
  NOR U1264 ( .A(n3443), .B(n2806), .Z(n3546) );
  ANDN U1265 ( .B(n1893), .A(n1894), .Z(n1891) );
  ANDN U1266 ( .B(n1927), .A(n1928), .Z(n1925) );
  ANDN U1267 ( .B(n1958), .A(n1959), .Z(n1956) );
  ANDN U1268 ( .B(n1990), .A(n1991), .Z(n1988) );
  ANDN U1269 ( .B(n2346), .A(n2347), .Z(n2344) );
  ANDN U1270 ( .B(n3084), .A(n3085), .Z(n3082) );
  ANDN U1271 ( .B(n3109), .A(n3110), .Z(n3107) );
  ANDN U1272 ( .B(n3129), .A(n3130), .Z(n3127) );
  ANDN U1273 ( .B(n3143), .A(n3144), .Z(n3141) );
  ANDN U1274 ( .B(n3157), .A(n3158), .Z(n3155) );
  XOR U1275 ( .A(n1051), .B(n1052), .Z(out[9]) );
  ANDN U1276 ( .B(n1053), .A(n1054), .Z(n1051) );
  XOR U1277 ( .A(n1055), .B(n1056), .Z(out[99]) );
  ANDN U1278 ( .B(n1057), .A(n1058), .Z(n1055) );
  XOR U1279 ( .A(n1059), .B(n1060), .Z(out[999]) );
  ANDN U1280 ( .B(n1061), .A(n1062), .Z(n1059) );
  XOR U1281 ( .A(n1063), .B(n1064), .Z(out[998]) );
  AND U1282 ( .A(n1065), .B(n1066), .Z(n1063) );
  XOR U1283 ( .A(n1067), .B(n1068), .Z(out[997]) );
  ANDN U1284 ( .B(n1069), .A(n1070), .Z(n1067) );
  XOR U1285 ( .A(n1071), .B(n1072), .Z(out[996]) );
  ANDN U1286 ( .B(n1073), .A(n1074), .Z(n1071) );
  XOR U1287 ( .A(n1075), .B(n1076), .Z(out[995]) );
  ANDN U1288 ( .B(n1077), .A(n1078), .Z(n1075) );
  XOR U1289 ( .A(n1079), .B(n1080), .Z(out[994]) );
  ANDN U1290 ( .B(n1081), .A(n1082), .Z(n1079) );
  XOR U1291 ( .A(n1083), .B(n1084), .Z(out[993]) );
  ANDN U1292 ( .B(n1085), .A(n1086), .Z(n1083) );
  XOR U1293 ( .A(n1087), .B(n1088), .Z(out[992]) );
  ANDN U1294 ( .B(n1089), .A(n1090), .Z(n1087) );
  XOR U1295 ( .A(n1091), .B(n1092), .Z(out[991]) );
  ANDN U1296 ( .B(n1093), .A(n1094), .Z(n1091) );
  XOR U1297 ( .A(n1095), .B(n1096), .Z(out[990]) );
  ANDN U1298 ( .B(n1097), .A(n1098), .Z(n1095) );
  XOR U1299 ( .A(n1099), .B(n1100), .Z(out[98]) );
  ANDN U1300 ( .B(n1101), .A(n1102), .Z(n1099) );
  XNOR U1301 ( .A(n1103), .B(n1104), .Z(out[989]) );
  ANDN U1302 ( .B(n1105), .A(n1106), .Z(n1103) );
  XNOR U1303 ( .A(n1107), .B(n1108), .Z(out[988]) );
  ANDN U1304 ( .B(n1109), .A(n1110), .Z(n1107) );
  XOR U1305 ( .A(n1111), .B(n1112), .Z(out[987]) );
  ANDN U1306 ( .B(n1113), .A(n1114), .Z(n1111) );
  XOR U1307 ( .A(n1115), .B(n1116), .Z(out[986]) );
  ANDN U1308 ( .B(n1117), .A(n1118), .Z(n1115) );
  XOR U1309 ( .A(n1119), .B(n1120), .Z(out[985]) );
  ANDN U1310 ( .B(n1121), .A(n1122), .Z(n1119) );
  XOR U1311 ( .A(n1123), .B(n1124), .Z(out[984]) );
  ANDN U1312 ( .B(n1125), .A(n1126), .Z(n1123) );
  XOR U1313 ( .A(n1127), .B(n1128), .Z(out[983]) );
  ANDN U1314 ( .B(n1129), .A(n1130), .Z(n1127) );
  XOR U1315 ( .A(n1131), .B(n1132), .Z(out[982]) );
  ANDN U1316 ( .B(n1133), .A(n1134), .Z(n1131) );
  XOR U1317 ( .A(n1135), .B(n1136), .Z(out[981]) );
  ANDN U1318 ( .B(n1137), .A(n1138), .Z(n1135) );
  XOR U1319 ( .A(n1139), .B(n1140), .Z(out[980]) );
  ANDN U1320 ( .B(n1141), .A(n1142), .Z(n1139) );
  XOR U1321 ( .A(n1143), .B(n1144), .Z(out[97]) );
  AND U1322 ( .A(n1145), .B(n1146), .Z(n1143) );
  XOR U1323 ( .A(n1147), .B(n1148), .Z(out[979]) );
  NOR U1324 ( .A(n1149), .B(n1150), .Z(n1147) );
  XOR U1325 ( .A(n1151), .B(n1152), .Z(out[978]) );
  ANDN U1326 ( .B(n1153), .A(n1154), .Z(n1151) );
  XOR U1327 ( .A(n1155), .B(n1156), .Z(out[977]) );
  ANDN U1328 ( .B(n1157), .A(n1158), .Z(n1155) );
  XOR U1329 ( .A(n1159), .B(n1160), .Z(out[976]) );
  ANDN U1330 ( .B(n1161), .A(n1162), .Z(n1159) );
  XNOR U1331 ( .A(n1163), .B(n1164), .Z(out[975]) );
  ANDN U1332 ( .B(n1165), .A(n1166), .Z(n1163) );
  XOR U1333 ( .A(n1167), .B(n1168), .Z(out[974]) );
  ANDN U1334 ( .B(n1169), .A(n1170), .Z(n1167) );
  XOR U1335 ( .A(n1171), .B(n1172), .Z(out[973]) );
  ANDN U1336 ( .B(n1173), .A(n1174), .Z(n1171) );
  XOR U1337 ( .A(n1175), .B(n1176), .Z(out[972]) );
  NOR U1338 ( .A(n1177), .B(n1178), .Z(n1175) );
  XOR U1339 ( .A(n1179), .B(n1180), .Z(out[971]) );
  NOR U1340 ( .A(n1181), .B(n1182), .Z(n1179) );
  XOR U1341 ( .A(n1183), .B(n1184), .Z(out[970]) );
  NOR U1342 ( .A(n1185), .B(n1186), .Z(n1183) );
  XNOR U1343 ( .A(n1187), .B(n1188), .Z(out[96]) );
  AND U1344 ( .A(n1189), .B(n1190), .Z(n1187) );
  XOR U1345 ( .A(n1191), .B(n1192), .Z(out[969]) );
  NOR U1346 ( .A(n1193), .B(n1194), .Z(n1191) );
  XNOR U1347 ( .A(n1195), .B(n1196), .Z(out[968]) );
  ANDN U1348 ( .B(n1197), .A(n1198), .Z(n1195) );
  XNOR U1349 ( .A(n1199), .B(n1200), .Z(out[967]) );
  ANDN U1350 ( .B(n1201), .A(n1202), .Z(n1199) );
  XNOR U1351 ( .A(n1203), .B(n1204), .Z(out[966]) );
  ANDN U1352 ( .B(n1205), .A(n1206), .Z(n1203) );
  XNOR U1353 ( .A(n1207), .B(n1208), .Z(out[965]) );
  AND U1354 ( .A(n1209), .B(n1210), .Z(n1207) );
  XNOR U1355 ( .A(n1211), .B(n1212), .Z(out[964]) );
  AND U1356 ( .A(n1213), .B(n1214), .Z(n1211) );
  XNOR U1357 ( .A(n1215), .B(n1216), .Z(out[963]) );
  AND U1358 ( .A(n1217), .B(n1218), .Z(n1215) );
  XNOR U1359 ( .A(n1219), .B(n1220), .Z(out[962]) );
  AND U1360 ( .A(n1221), .B(n1222), .Z(n1219) );
  XNOR U1361 ( .A(n1223), .B(n1224), .Z(out[961]) );
  AND U1362 ( .A(n1225), .B(n1226), .Z(n1223) );
  XNOR U1363 ( .A(n1227), .B(n1228), .Z(out[960]) );
  AND U1364 ( .A(n1229), .B(n1230), .Z(n1227) );
  XNOR U1365 ( .A(n1231), .B(n1232), .Z(out[95]) );
  AND U1366 ( .A(n1233), .B(n1234), .Z(n1231) );
  XOR U1367 ( .A(n1235), .B(n1236), .Z(out[959]) );
  AND U1368 ( .A(n1237), .B(n1238), .Z(n1235) );
  XOR U1369 ( .A(n1239), .B(n1240), .Z(out[958]) );
  AND U1370 ( .A(n1241), .B(n1242), .Z(n1239) );
  XOR U1371 ( .A(n1243), .B(n1244), .Z(out[957]) );
  AND U1372 ( .A(n1245), .B(n1246), .Z(n1243) );
  XOR U1373 ( .A(n1247), .B(n1248), .Z(out[956]) );
  AND U1374 ( .A(n1249), .B(n1250), .Z(n1247) );
  XOR U1375 ( .A(n1251), .B(n1252), .Z(out[955]) );
  AND U1376 ( .A(n1253), .B(n1254), .Z(n1251) );
  XNOR U1377 ( .A(n1255), .B(n1256), .Z(out[954]) );
  AND U1378 ( .A(n1257), .B(n1258), .Z(n1255) );
  XNOR U1379 ( .A(n1259), .B(n1260), .Z(out[953]) );
  AND U1380 ( .A(n1261), .B(n1262), .Z(n1259) );
  XNOR U1381 ( .A(n1263), .B(n1264), .Z(out[952]) );
  AND U1382 ( .A(n1265), .B(n1266), .Z(n1263) );
  XNOR U1383 ( .A(n1267), .B(n1268), .Z(out[951]) );
  AND U1384 ( .A(n1269), .B(n1270), .Z(n1267) );
  XNOR U1385 ( .A(n1271), .B(n1272), .Z(out[950]) );
  AND U1386 ( .A(n1273), .B(n1274), .Z(n1271) );
  XNOR U1387 ( .A(n1275), .B(n1276), .Z(out[94]) );
  AND U1388 ( .A(n1277), .B(n1278), .Z(n1275) );
  XNOR U1389 ( .A(n1279), .B(n1280), .Z(out[949]) );
  AND U1390 ( .A(n1281), .B(n1282), .Z(n1279) );
  XNOR U1391 ( .A(n1283), .B(n1284), .Z(out[948]) );
  AND U1392 ( .A(n1285), .B(n1286), .Z(n1283) );
  XNOR U1393 ( .A(n1287), .B(n1288), .Z(out[947]) );
  AND U1394 ( .A(n1289), .B(n1290), .Z(n1287) );
  XNOR U1395 ( .A(n1291), .B(n1292), .Z(out[946]) );
  AND U1396 ( .A(n1293), .B(n1294), .Z(n1291) );
  XNOR U1397 ( .A(n1295), .B(n1296), .Z(out[945]) );
  AND U1398 ( .A(n1297), .B(n1298), .Z(n1295) );
  XNOR U1399 ( .A(n1299), .B(n1300), .Z(out[944]) );
  AND U1400 ( .A(n1301), .B(n1302), .Z(n1299) );
  XNOR U1401 ( .A(n1303), .B(n1304), .Z(out[943]) );
  AND U1402 ( .A(n1305), .B(n1306), .Z(n1303) );
  XNOR U1403 ( .A(n1307), .B(n1308), .Z(out[942]) );
  AND U1404 ( .A(n1309), .B(n1310), .Z(n1307) );
  XNOR U1405 ( .A(n1311), .B(n1312), .Z(out[941]) );
  AND U1406 ( .A(n1313), .B(n1314), .Z(n1311) );
  XNOR U1407 ( .A(n1315), .B(n1316), .Z(out[940]) );
  AND U1408 ( .A(n1317), .B(n1318), .Z(n1315) );
  XNOR U1409 ( .A(n1319), .B(n1320), .Z(out[93]) );
  AND U1410 ( .A(n1321), .B(n1322), .Z(n1319) );
  XNOR U1411 ( .A(n1323), .B(n1324), .Z(out[939]) );
  AND U1412 ( .A(n1325), .B(n1326), .Z(n1323) );
  XNOR U1413 ( .A(n1327), .B(n1328), .Z(out[938]) );
  AND U1414 ( .A(n1329), .B(n1330), .Z(n1327) );
  XNOR U1415 ( .A(n1331), .B(n1332), .Z(out[937]) );
  AND U1416 ( .A(n1333), .B(n1334), .Z(n1331) );
  XNOR U1417 ( .A(n1335), .B(n1336), .Z(out[936]) );
  AND U1418 ( .A(n1337), .B(n1338), .Z(n1335) );
  XNOR U1419 ( .A(n1339), .B(n1340), .Z(out[935]) );
  AND U1420 ( .A(n1341), .B(n1342), .Z(n1339) );
  XNOR U1421 ( .A(n1343), .B(n1344), .Z(out[934]) );
  AND U1422 ( .A(n1345), .B(n1346), .Z(n1343) );
  XNOR U1423 ( .A(n1347), .B(n1348), .Z(out[933]) );
  AND U1424 ( .A(n1349), .B(n1350), .Z(n1347) );
  XNOR U1425 ( .A(n1351), .B(n1352), .Z(out[932]) );
  AND U1426 ( .A(n1353), .B(n1354), .Z(n1351) );
  XNOR U1427 ( .A(n1355), .B(n1356), .Z(out[931]) );
  AND U1428 ( .A(n1357), .B(n1358), .Z(n1355) );
  XNOR U1429 ( .A(n1359), .B(n1360), .Z(out[930]) );
  AND U1430 ( .A(n1361), .B(n1362), .Z(n1359) );
  XNOR U1431 ( .A(n1363), .B(n1364), .Z(out[92]) );
  AND U1432 ( .A(n1365), .B(n1366), .Z(n1363) );
  XNOR U1433 ( .A(n1367), .B(n1368), .Z(out[929]) );
  AND U1434 ( .A(n1369), .B(n1370), .Z(n1367) );
  XNOR U1435 ( .A(n1371), .B(n1372), .Z(out[928]) );
  AND U1436 ( .A(n1373), .B(n1374), .Z(n1371) );
  XNOR U1437 ( .A(n1375), .B(n1376), .Z(out[927]) );
  AND U1438 ( .A(n1377), .B(n1378), .Z(n1375) );
  XNOR U1439 ( .A(n1379), .B(n1380), .Z(out[926]) );
  AND U1440 ( .A(n1381), .B(n1382), .Z(n1379) );
  XNOR U1441 ( .A(n1383), .B(n1384), .Z(out[925]) );
  AND U1442 ( .A(n1385), .B(n1386), .Z(n1383) );
  XNOR U1443 ( .A(n1387), .B(n1388), .Z(out[924]) );
  AND U1444 ( .A(n1389), .B(n1390), .Z(n1387) );
  XNOR U1445 ( .A(n1391), .B(n1392), .Z(out[923]) );
  AND U1446 ( .A(n1393), .B(n1394), .Z(n1391) );
  XNOR U1447 ( .A(n1395), .B(n1396), .Z(out[922]) );
  AND U1448 ( .A(n1397), .B(n1398), .Z(n1395) );
  XNOR U1449 ( .A(n1399), .B(n1400), .Z(out[921]) );
  AND U1450 ( .A(n1401), .B(n1402), .Z(n1399) );
  XNOR U1451 ( .A(n1403), .B(n1404), .Z(out[920]) );
  AND U1452 ( .A(n1405), .B(n1406), .Z(n1403) );
  XNOR U1453 ( .A(n1407), .B(n1408), .Z(out[91]) );
  AND U1454 ( .A(n1409), .B(n1410), .Z(n1407) );
  XNOR U1455 ( .A(n1411), .B(n1412), .Z(out[919]) );
  AND U1456 ( .A(n1413), .B(n1414), .Z(n1411) );
  XNOR U1457 ( .A(n1415), .B(n1416), .Z(out[918]) );
  AND U1458 ( .A(n1417), .B(n1418), .Z(n1415) );
  XNOR U1459 ( .A(n1419), .B(n1420), .Z(out[917]) );
  AND U1460 ( .A(n1421), .B(n1422), .Z(n1419) );
  XNOR U1461 ( .A(n1423), .B(n1424), .Z(out[916]) );
  AND U1462 ( .A(n1425), .B(n1426), .Z(n1423) );
  XNOR U1463 ( .A(n1427), .B(n1428), .Z(out[915]) );
  AND U1464 ( .A(n1429), .B(n1430), .Z(n1427) );
  XNOR U1465 ( .A(n1431), .B(n1432), .Z(out[914]) );
  AND U1466 ( .A(n1433), .B(n1434), .Z(n1431) );
  XNOR U1467 ( .A(n1435), .B(n1436), .Z(out[913]) );
  AND U1468 ( .A(n1437), .B(n1438), .Z(n1435) );
  XNOR U1469 ( .A(n1439), .B(n1440), .Z(out[912]) );
  AND U1470 ( .A(n1441), .B(n1442), .Z(n1439) );
  XNOR U1471 ( .A(n1443), .B(n1444), .Z(out[911]) );
  AND U1472 ( .A(n1445), .B(n1446), .Z(n1443) );
  XNOR U1473 ( .A(n1447), .B(n1448), .Z(out[910]) );
  AND U1474 ( .A(n1449), .B(n1450), .Z(n1447) );
  XNOR U1475 ( .A(n1451), .B(n1452), .Z(out[90]) );
  AND U1476 ( .A(n1453), .B(n1454), .Z(n1451) );
  XNOR U1477 ( .A(n1455), .B(n1456), .Z(out[909]) );
  AND U1478 ( .A(n1457), .B(n1458), .Z(n1455) );
  XNOR U1479 ( .A(n1459), .B(n1460), .Z(out[908]) );
  AND U1480 ( .A(n1461), .B(n1462), .Z(n1459) );
  XNOR U1481 ( .A(n1463), .B(n1464), .Z(out[907]) );
  AND U1482 ( .A(n1465), .B(n1466), .Z(n1463) );
  XNOR U1483 ( .A(n1467), .B(n1468), .Z(out[906]) );
  AND U1484 ( .A(n1469), .B(n1470), .Z(n1467) );
  XNOR U1485 ( .A(n1471), .B(n1472), .Z(out[905]) );
  AND U1486 ( .A(n1473), .B(n1474), .Z(n1471) );
  XNOR U1487 ( .A(n1475), .B(n1476), .Z(out[904]) );
  AND U1488 ( .A(n1477), .B(n1478), .Z(n1475) );
  XNOR U1489 ( .A(n1479), .B(n1480), .Z(out[903]) );
  AND U1490 ( .A(n1481), .B(n1482), .Z(n1479) );
  XNOR U1491 ( .A(n1483), .B(n1484), .Z(out[902]) );
  AND U1492 ( .A(n1485), .B(n1486), .Z(n1483) );
  XNOR U1493 ( .A(n1487), .B(n1488), .Z(out[901]) );
  AND U1494 ( .A(n1489), .B(n1490), .Z(n1487) );
  XNOR U1495 ( .A(n1491), .B(n1492), .Z(out[900]) );
  AND U1496 ( .A(n1493), .B(n1494), .Z(n1491) );
  XNOR U1497 ( .A(n1495), .B(n1496), .Z(out[8]) );
  NOR U1498 ( .A(n1497), .B(n1498), .Z(n1495) );
  XNOR U1499 ( .A(n1499), .B(n1500), .Z(out[89]) );
  AND U1500 ( .A(n1501), .B(n1502), .Z(n1499) );
  XNOR U1501 ( .A(n1503), .B(n1504), .Z(out[899]) );
  AND U1502 ( .A(n1505), .B(n1506), .Z(n1503) );
  XNOR U1503 ( .A(n1507), .B(n1508), .Z(out[898]) );
  AND U1504 ( .A(n1509), .B(n1510), .Z(n1507) );
  XNOR U1505 ( .A(n1511), .B(n1512), .Z(out[897]) );
  AND U1506 ( .A(n1513), .B(n1514), .Z(n1511) );
  XNOR U1507 ( .A(n1515), .B(n1516), .Z(out[896]) );
  AND U1508 ( .A(n1517), .B(n1518), .Z(n1515) );
  XNOR U1509 ( .A(n1519), .B(n1237), .Z(out[895]) );
  XNOR U1510 ( .A(n1521), .B(n1241), .Z(out[894]) );
  XNOR U1511 ( .A(n1523), .B(n1245), .Z(out[893]) );
  XNOR U1512 ( .A(n1525), .B(n1249), .Z(out[892]) );
  XNOR U1513 ( .A(n1527), .B(n1253), .Z(out[891]) );
  AND U1514 ( .A(n1528), .B(n1529), .Z(n1527) );
  XNOR U1515 ( .A(n1530), .B(n1257), .Z(out[890]) );
  AND U1516 ( .A(n1531), .B(n1532), .Z(n1530) );
  XNOR U1517 ( .A(n1533), .B(n1534), .Z(out[88]) );
  AND U1518 ( .A(n1535), .B(n1536), .Z(n1533) );
  XNOR U1519 ( .A(n1537), .B(n1261), .Z(out[889]) );
  AND U1520 ( .A(n1538), .B(n1539), .Z(n1537) );
  XNOR U1521 ( .A(n1540), .B(n1265), .Z(out[888]) );
  AND U1522 ( .A(n1541), .B(n1542), .Z(n1540) );
  XNOR U1523 ( .A(n1543), .B(n1269), .Z(out[887]) );
  AND U1524 ( .A(n1544), .B(n1545), .Z(n1543) );
  XNOR U1525 ( .A(n1546), .B(n1273), .Z(out[886]) );
  AND U1526 ( .A(n1547), .B(n1548), .Z(n1546) );
  XNOR U1527 ( .A(n1549), .B(n1281), .Z(out[885]) );
  AND U1528 ( .A(n1550), .B(n1551), .Z(n1549) );
  XNOR U1529 ( .A(n1552), .B(n1285), .Z(out[884]) );
  AND U1530 ( .A(n1553), .B(n1554), .Z(n1552) );
  XNOR U1531 ( .A(n1555), .B(n1289), .Z(out[883]) );
  XNOR U1532 ( .A(n1557), .B(n1293), .Z(out[882]) );
  XNOR U1533 ( .A(n1559), .B(n1297), .Z(out[881]) );
  XNOR U1534 ( .A(n1561), .B(n1301), .Z(out[880]) );
  XNOR U1535 ( .A(n1563), .B(n1564), .Z(out[87]) );
  AND U1536 ( .A(n1565), .B(n1566), .Z(n1563) );
  XNOR U1537 ( .A(n1567), .B(n1305), .Z(out[879]) );
  XNOR U1538 ( .A(n1569), .B(n1309), .Z(out[878]) );
  XNOR U1539 ( .A(n1571), .B(n1313), .Z(out[877]) );
  XNOR U1540 ( .A(n1573), .B(n1317), .Z(out[876]) );
  XNOR U1541 ( .A(n1575), .B(n1325), .Z(out[875]) );
  AND U1542 ( .A(n1576), .B(n1577), .Z(n1575) );
  XNOR U1543 ( .A(n1578), .B(n1329), .Z(out[874]) );
  XNOR U1544 ( .A(n1580), .B(n1333), .Z(out[873]) );
  XNOR U1545 ( .A(n1582), .B(n1337), .Z(out[872]) );
  XNOR U1546 ( .A(n1584), .B(n1341), .Z(out[871]) );
  XNOR U1547 ( .A(n1586), .B(n1345), .Z(out[870]) );
  XNOR U1548 ( .A(n1588), .B(n1589), .Z(out[86]) );
  AND U1549 ( .A(n1590), .B(n1591), .Z(n1588) );
  XNOR U1550 ( .A(n1592), .B(n1349), .Z(out[869]) );
  XNOR U1551 ( .A(n1594), .B(n1353), .Z(out[868]) );
  AND U1552 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1553 ( .A(n1597), .B(n1357), .Z(out[867]) );
  AND U1554 ( .A(n1598), .B(n1599), .Z(n1597) );
  XNOR U1555 ( .A(n1600), .B(n1361), .Z(out[866]) );
  AND U1556 ( .A(n1601), .B(n1602), .Z(n1600) );
  XNOR U1557 ( .A(n1603), .B(n1369), .Z(out[865]) );
  AND U1558 ( .A(n1604), .B(n1605), .Z(n1603) );
  XNOR U1559 ( .A(n1606), .B(n1373), .Z(out[864]) );
  AND U1560 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1561 ( .A(n1609), .B(n1377), .Z(out[863]) );
  AND U1562 ( .A(n1610), .B(n1611), .Z(n1609) );
  XNOR U1563 ( .A(n1612), .B(n1381), .Z(out[862]) );
  AND U1564 ( .A(n1613), .B(n1614), .Z(n1612) );
  XNOR U1565 ( .A(n1615), .B(n1385), .Z(out[861]) );
  AND U1566 ( .A(n1616), .B(n1617), .Z(n1615) );
  XNOR U1567 ( .A(n1618), .B(n1389), .Z(out[860]) );
  AND U1568 ( .A(n1619), .B(n1620), .Z(n1618) );
  XNOR U1569 ( .A(n1621), .B(n1622), .Z(out[85]) );
  AND U1570 ( .A(n1623), .B(n1624), .Z(n1621) );
  XNOR U1571 ( .A(n1625), .B(n1393), .Z(out[859]) );
  AND U1572 ( .A(n1626), .B(n1627), .Z(n1625) );
  XNOR U1573 ( .A(n1628), .B(n1397), .Z(out[858]) );
  AND U1574 ( .A(n1629), .B(n1630), .Z(n1628) );
  XNOR U1575 ( .A(n1631), .B(n1401), .Z(out[857]) );
  AND U1576 ( .A(n1632), .B(n1633), .Z(n1631) );
  XNOR U1577 ( .A(n1634), .B(n1405), .Z(out[856]) );
  AND U1578 ( .A(n1635), .B(n1636), .Z(n1634) );
  XNOR U1579 ( .A(n1637), .B(n1413), .Z(out[855]) );
  AND U1580 ( .A(n1638), .B(n1639), .Z(n1637) );
  XNOR U1581 ( .A(n1640), .B(n1417), .Z(out[854]) );
  AND U1582 ( .A(n1641), .B(n1642), .Z(n1640) );
  XNOR U1583 ( .A(n1643), .B(n1421), .Z(out[853]) );
  AND U1584 ( .A(n1644), .B(n1645), .Z(n1643) );
  XNOR U1585 ( .A(n1646), .B(n1425), .Z(out[852]) );
  AND U1586 ( .A(n1647), .B(n1648), .Z(n1646) );
  XNOR U1587 ( .A(n1649), .B(n1429), .Z(out[851]) );
  AND U1588 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1589 ( .A(n1652), .B(n1433), .Z(out[850]) );
  AND U1590 ( .A(n1653), .B(n1654), .Z(n1652) );
  XNOR U1591 ( .A(n1655), .B(n1656), .Z(out[84]) );
  AND U1592 ( .A(n1657), .B(n1658), .Z(n1655) );
  XNOR U1593 ( .A(n1659), .B(n1437), .Z(out[849]) );
  AND U1594 ( .A(n1660), .B(n1661), .Z(n1659) );
  XNOR U1595 ( .A(n1662), .B(n1441), .Z(out[848]) );
  AND U1596 ( .A(n1663), .B(n1664), .Z(n1662) );
  XNOR U1597 ( .A(n1665), .B(n1445), .Z(out[847]) );
  AND U1598 ( .A(n1666), .B(n1667), .Z(n1665) );
  XNOR U1599 ( .A(n1668), .B(n1449), .Z(out[846]) );
  AND U1600 ( .A(n1669), .B(n1670), .Z(n1668) );
  XNOR U1601 ( .A(n1671), .B(n1457), .Z(out[845]) );
  AND U1602 ( .A(n1672), .B(n1673), .Z(n1671) );
  XNOR U1603 ( .A(n1674), .B(n1461), .Z(out[844]) );
  AND U1604 ( .A(n1675), .B(n1676), .Z(n1674) );
  XNOR U1605 ( .A(n1677), .B(n1465), .Z(out[843]) );
  AND U1606 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U1607 ( .A(n1680), .B(n1469), .Z(out[842]) );
  AND U1608 ( .A(n1681), .B(n1682), .Z(n1680) );
  XNOR U1609 ( .A(n1683), .B(n1473), .Z(out[841]) );
  AND U1610 ( .A(n1684), .B(n1685), .Z(n1683) );
  XNOR U1611 ( .A(n1686), .B(n1477), .Z(out[840]) );
  AND U1612 ( .A(n1687), .B(n1688), .Z(n1686) );
  XNOR U1613 ( .A(n1689), .B(n1690), .Z(out[83]) );
  AND U1614 ( .A(n1691), .B(n1692), .Z(n1689) );
  XNOR U1615 ( .A(n1693), .B(n1481), .Z(out[839]) );
  AND U1616 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U1617 ( .A(n1696), .B(n1485), .Z(out[838]) );
  AND U1618 ( .A(n1697), .B(n1698), .Z(n1696) );
  XNOR U1619 ( .A(n1699), .B(n1489), .Z(out[837]) );
  XNOR U1620 ( .A(n1701), .B(n1493), .Z(out[836]) );
  XNOR U1621 ( .A(n1703), .B(n1505), .Z(out[835]) );
  XNOR U1622 ( .A(n1705), .B(n1509), .Z(out[834]) );
  XNOR U1623 ( .A(n1707), .B(n1513), .Z(out[833]) );
  XNOR U1624 ( .A(n1709), .B(n1517), .Z(out[832]) );
  XOR U1625 ( .A(n1711), .B(n1238), .Z(out[831]) );
  XNOR U1626 ( .A(round_reg[742]), .B(n1712), .Z(n1238) );
  XOR U1627 ( .A(n1714), .B(n1242), .Z(out[830]) );
  XNOR U1628 ( .A(round_reg[741]), .B(n1715), .Z(n1242) );
  XNOR U1629 ( .A(n1717), .B(n1718), .Z(out[82]) );
  AND U1630 ( .A(n1719), .B(n1720), .Z(n1717) );
  XOR U1631 ( .A(n1721), .B(n1246), .Z(out[829]) );
  XNOR U1632 ( .A(round_reg[740]), .B(n1722), .Z(n1246) );
  XOR U1633 ( .A(n1724), .B(n1250), .Z(out[828]) );
  XNOR U1634 ( .A(round_reg[739]), .B(n1725), .Z(n1250) );
  NOR U1635 ( .A(n1726), .B(n1526), .Z(n1724) );
  XOR U1636 ( .A(n1727), .B(n1254), .Z(out[827]) );
  IV U1637 ( .A(n1529), .Z(n1254) );
  XNOR U1638 ( .A(round_reg[738]), .B(n1728), .Z(n1529) );
  NOR U1639 ( .A(n1729), .B(n1528), .Z(n1727) );
  XOR U1640 ( .A(n1730), .B(n1258), .Z(out[826]) );
  IV U1641 ( .A(n1532), .Z(n1258) );
  XNOR U1642 ( .A(round_reg[737]), .B(n1731), .Z(n1532) );
  NOR U1643 ( .A(n1732), .B(n1531), .Z(n1730) );
  XOR U1644 ( .A(n1733), .B(n1262), .Z(out[825]) );
  IV U1645 ( .A(n1539), .Z(n1262) );
  XNOR U1646 ( .A(round_reg[736]), .B(n1734), .Z(n1539) );
  NOR U1647 ( .A(n1735), .B(n1538), .Z(n1733) );
  XOR U1648 ( .A(n1736), .B(n1266), .Z(out[824]) );
  IV U1649 ( .A(n1542), .Z(n1266) );
  XNOR U1650 ( .A(round_reg[735]), .B(n1737), .Z(n1542) );
  NOR U1651 ( .A(n1738), .B(n1541), .Z(n1736) );
  XOR U1652 ( .A(n1739), .B(n1270), .Z(out[823]) );
  IV U1653 ( .A(n1545), .Z(n1270) );
  XNOR U1654 ( .A(round_reg[734]), .B(n1740), .Z(n1545) );
  NOR U1655 ( .A(n1741), .B(n1544), .Z(n1739) );
  XOR U1656 ( .A(n1742), .B(n1274), .Z(out[822]) );
  IV U1657 ( .A(n1548), .Z(n1274) );
  XNOR U1658 ( .A(round_reg[733]), .B(n1743), .Z(n1548) );
  NOR U1659 ( .A(n1744), .B(n1547), .Z(n1742) );
  XOR U1660 ( .A(n1745), .B(n1282), .Z(out[821]) );
  IV U1661 ( .A(n1551), .Z(n1282) );
  XNOR U1662 ( .A(round_reg[732]), .B(n1746), .Z(n1551) );
  NOR U1663 ( .A(n1747), .B(n1550), .Z(n1745) );
  XOR U1664 ( .A(n1748), .B(n1286), .Z(out[820]) );
  IV U1665 ( .A(n1554), .Z(n1286) );
  XNOR U1666 ( .A(round_reg[731]), .B(n1749), .Z(n1554) );
  NOR U1667 ( .A(n1750), .B(n1553), .Z(n1748) );
  XNOR U1668 ( .A(n1751), .B(n1752), .Z(out[81]) );
  AND U1669 ( .A(n1753), .B(n1754), .Z(n1751) );
  XOR U1670 ( .A(n1755), .B(n1290), .Z(out[819]) );
  XNOR U1671 ( .A(round_reg[730]), .B(n1756), .Z(n1290) );
  XOR U1672 ( .A(n1758), .B(n1294), .Z(out[818]) );
  XNOR U1673 ( .A(round_reg[729]), .B(n1759), .Z(n1294) );
  XOR U1674 ( .A(n1761), .B(n1298), .Z(out[817]) );
  XNOR U1675 ( .A(round_reg[728]), .B(n1762), .Z(n1298) );
  NOR U1676 ( .A(n1763), .B(n1560), .Z(n1761) );
  XOR U1677 ( .A(n1764), .B(n1302), .Z(out[816]) );
  XNOR U1678 ( .A(round_reg[727]), .B(n1765), .Z(n1302) );
  NOR U1679 ( .A(n1766), .B(n1562), .Z(n1764) );
  XOR U1680 ( .A(n1767), .B(n1306), .Z(out[815]) );
  XNOR U1681 ( .A(round_reg[726]), .B(n1768), .Z(n1306) );
  NOR U1682 ( .A(n1769), .B(n1568), .Z(n1767) );
  XOR U1683 ( .A(n1770), .B(n1310), .Z(out[814]) );
  XNOR U1684 ( .A(round_reg[725]), .B(n1771), .Z(n1310) );
  NOR U1685 ( .A(n1772), .B(n1570), .Z(n1770) );
  XOR U1686 ( .A(n1773), .B(n1314), .Z(out[813]) );
  XNOR U1687 ( .A(round_reg[724]), .B(n1774), .Z(n1314) );
  NOR U1688 ( .A(n1775), .B(n1572), .Z(n1773) );
  XOR U1689 ( .A(n1776), .B(n1318), .Z(out[812]) );
  XNOR U1690 ( .A(round_reg[723]), .B(n1777), .Z(n1318) );
  NOR U1691 ( .A(n1778), .B(n1574), .Z(n1776) );
  XOR U1692 ( .A(n1779), .B(n1326), .Z(out[811]) );
  IV U1693 ( .A(n1577), .Z(n1326) );
  XNOR U1694 ( .A(round_reg[722]), .B(n1780), .Z(n1577) );
  NOR U1695 ( .A(n1781), .B(n1576), .Z(n1779) );
  XOR U1696 ( .A(n1782), .B(n1330), .Z(out[810]) );
  XOR U1697 ( .A(round_reg[721]), .B(n1783), .Z(n1330) );
  XNOR U1698 ( .A(n1785), .B(n1786), .Z(out[80]) );
  AND U1699 ( .A(n1787), .B(n1788), .Z(n1785) );
  XOR U1700 ( .A(n1789), .B(n1334), .Z(out[809]) );
  XOR U1701 ( .A(round_reg[720]), .B(n1790), .Z(n1334) );
  XOR U1702 ( .A(n1792), .B(n1338), .Z(out[808]) );
  XOR U1703 ( .A(round_reg[719]), .B(n1793), .Z(n1338) );
  XOR U1704 ( .A(n1795), .B(n1342), .Z(out[807]) );
  XOR U1705 ( .A(round_reg[718]), .B(n1796), .Z(n1342) );
  XOR U1706 ( .A(n1798), .B(n1346), .Z(out[806]) );
  XOR U1707 ( .A(round_reg[717]), .B(n1799), .Z(n1346) );
  XOR U1708 ( .A(n1801), .B(n1350), .Z(out[805]) );
  XOR U1709 ( .A(round_reg[716]), .B(n1802), .Z(n1350) );
  XOR U1710 ( .A(n1804), .B(n1354), .Z(out[804]) );
  IV U1711 ( .A(n1596), .Z(n1354) );
  XNOR U1712 ( .A(round_reg[715]), .B(n1805), .Z(n1596) );
  NOR U1713 ( .A(n1806), .B(n1595), .Z(n1804) );
  XOR U1714 ( .A(n1807), .B(n1358), .Z(out[803]) );
  IV U1715 ( .A(n1599), .Z(n1358) );
  XNOR U1716 ( .A(round_reg[714]), .B(n1808), .Z(n1599) );
  ANDN U1717 ( .B(n1809), .A(n1598), .Z(n1807) );
  XOR U1718 ( .A(n1810), .B(n1362), .Z(out[802]) );
  IV U1719 ( .A(n1602), .Z(n1362) );
  XNOR U1720 ( .A(round_reg[713]), .B(n1811), .Z(n1602) );
  NOR U1721 ( .A(n1812), .B(n1601), .Z(n1810) );
  XOR U1722 ( .A(n1813), .B(n1370), .Z(out[801]) );
  IV U1723 ( .A(n1605), .Z(n1370) );
  XNOR U1724 ( .A(round_reg[712]), .B(n1814), .Z(n1605) );
  NOR U1725 ( .A(n1815), .B(n1604), .Z(n1813) );
  XOR U1726 ( .A(n1816), .B(n1374), .Z(out[800]) );
  IV U1727 ( .A(n1608), .Z(n1374) );
  XNOR U1728 ( .A(round_reg[711]), .B(n1817), .Z(n1608) );
  NOR U1729 ( .A(n1818), .B(n1607), .Z(n1816) );
  XNOR U1730 ( .A(n1819), .B(n1820), .Z(out[7]) );
  NOR U1731 ( .A(n1821), .B(n1822), .Z(n1819) );
  XNOR U1732 ( .A(n1823), .B(n1824), .Z(out[79]) );
  AND U1733 ( .A(n1825), .B(n1826), .Z(n1823) );
  XOR U1734 ( .A(n1827), .B(n1378), .Z(out[799]) );
  IV U1735 ( .A(n1611), .Z(n1378) );
  XNOR U1736 ( .A(round_reg[710]), .B(n1828), .Z(n1611) );
  NOR U1737 ( .A(n1829), .B(n1610), .Z(n1827) );
  XOR U1738 ( .A(n1830), .B(n1382), .Z(out[798]) );
  IV U1739 ( .A(n1614), .Z(n1382) );
  XNOR U1740 ( .A(round_reg[709]), .B(n1831), .Z(n1614) );
  NOR U1741 ( .A(n1832), .B(n1613), .Z(n1830) );
  XOR U1742 ( .A(n1833), .B(n1386), .Z(out[797]) );
  IV U1743 ( .A(n1617), .Z(n1386) );
  XNOR U1744 ( .A(round_reg[708]), .B(n1834), .Z(n1617) );
  NOR U1745 ( .A(n1835), .B(n1616), .Z(n1833) );
  XOR U1746 ( .A(n1836), .B(n1390), .Z(out[796]) );
  IV U1747 ( .A(n1620), .Z(n1390) );
  XNOR U1748 ( .A(round_reg[707]), .B(n1837), .Z(n1620) );
  ANDN U1749 ( .B(n1838), .A(n1619), .Z(n1836) );
  XOR U1750 ( .A(n1839), .B(n1394), .Z(out[795]) );
  IV U1751 ( .A(n1627), .Z(n1394) );
  XNOR U1752 ( .A(round_reg[706]), .B(n1840), .Z(n1627) );
  ANDN U1753 ( .B(n1841), .A(n1626), .Z(n1839) );
  XOR U1754 ( .A(n1842), .B(n1398), .Z(out[794]) );
  IV U1755 ( .A(n1630), .Z(n1398) );
  XNOR U1756 ( .A(round_reg[705]), .B(n1843), .Z(n1630) );
  ANDN U1757 ( .B(n1844), .A(n1629), .Z(n1842) );
  XOR U1758 ( .A(n1845), .B(n1402), .Z(out[793]) );
  IV U1759 ( .A(n1633), .Z(n1402) );
  XNOR U1760 ( .A(round_reg[704]), .B(n1846), .Z(n1633) );
  ANDN U1761 ( .B(n1847), .A(n1632), .Z(n1845) );
  XOR U1762 ( .A(n1848), .B(n1406), .Z(out[792]) );
  IV U1763 ( .A(n1636), .Z(n1406) );
  XNOR U1764 ( .A(round_reg[767]), .B(n1849), .Z(n1636) );
  ANDN U1765 ( .B(n1850), .A(n1635), .Z(n1848) );
  XOR U1766 ( .A(n1851), .B(n1414), .Z(out[791]) );
  IV U1767 ( .A(n1639), .Z(n1414) );
  XNOR U1768 ( .A(round_reg[766]), .B(n1852), .Z(n1639) );
  ANDN U1769 ( .B(n1853), .A(n1638), .Z(n1851) );
  XOR U1770 ( .A(n1854), .B(n1418), .Z(out[790]) );
  IV U1771 ( .A(n1642), .Z(n1418) );
  XNOR U1772 ( .A(round_reg[765]), .B(n1855), .Z(n1642) );
  ANDN U1773 ( .B(n1856), .A(n1641), .Z(n1854) );
  XNOR U1774 ( .A(n1857), .B(n1858), .Z(out[78]) );
  AND U1775 ( .A(n1859), .B(n1860), .Z(n1857) );
  XOR U1776 ( .A(n1861), .B(n1422), .Z(out[789]) );
  IV U1777 ( .A(n1645), .Z(n1422) );
  XNOR U1778 ( .A(round_reg[764]), .B(n1862), .Z(n1645) );
  ANDN U1779 ( .B(n1863), .A(n1644), .Z(n1861) );
  XOR U1780 ( .A(n1864), .B(n1426), .Z(out[788]) );
  IV U1781 ( .A(n1648), .Z(n1426) );
  XNOR U1782 ( .A(round_reg[763]), .B(n1865), .Z(n1648) );
  ANDN U1783 ( .B(n1866), .A(n1647), .Z(n1864) );
  XOR U1784 ( .A(n1867), .B(n1430), .Z(out[787]) );
  IV U1785 ( .A(n1651), .Z(n1430) );
  XNOR U1786 ( .A(round_reg[762]), .B(n1868), .Z(n1651) );
  ANDN U1787 ( .B(n1869), .A(n1650), .Z(n1867) );
  XOR U1788 ( .A(n1870), .B(n1434), .Z(out[786]) );
  IV U1789 ( .A(n1654), .Z(n1434) );
  XNOR U1790 ( .A(round_reg[761]), .B(n1871), .Z(n1654) );
  ANDN U1791 ( .B(n1872), .A(n1653), .Z(n1870) );
  XOR U1792 ( .A(n1873), .B(n1438), .Z(out[785]) );
  IV U1793 ( .A(n1661), .Z(n1438) );
  XNOR U1794 ( .A(round_reg[760]), .B(n1874), .Z(n1661) );
  ANDN U1795 ( .B(n1875), .A(n1660), .Z(n1873) );
  XOR U1796 ( .A(n1876), .B(n1442), .Z(out[784]) );
  IV U1797 ( .A(n1664), .Z(n1442) );
  XNOR U1798 ( .A(round_reg[759]), .B(n1877), .Z(n1664) );
  ANDN U1799 ( .B(n1878), .A(n1663), .Z(n1876) );
  XOR U1800 ( .A(n1879), .B(n1446), .Z(out[783]) );
  IV U1801 ( .A(n1667), .Z(n1446) );
  XNOR U1802 ( .A(round_reg[758]), .B(n1880), .Z(n1667) );
  ANDN U1803 ( .B(n1881), .A(n1666), .Z(n1879) );
  XOR U1804 ( .A(n1882), .B(n1450), .Z(out[782]) );
  IV U1805 ( .A(n1670), .Z(n1450) );
  XNOR U1806 ( .A(round_reg[757]), .B(n1883), .Z(n1670) );
  ANDN U1807 ( .B(n1884), .A(n1669), .Z(n1882) );
  XOR U1808 ( .A(n1885), .B(n1458), .Z(out[781]) );
  IV U1809 ( .A(n1673), .Z(n1458) );
  XNOR U1810 ( .A(round_reg[756]), .B(n1886), .Z(n1673) );
  ANDN U1811 ( .B(n1887), .A(n1672), .Z(n1885) );
  XOR U1812 ( .A(n1888), .B(n1462), .Z(out[780]) );
  IV U1813 ( .A(n1676), .Z(n1462) );
  XNOR U1814 ( .A(round_reg[755]), .B(n1889), .Z(n1676) );
  ANDN U1815 ( .B(n1890), .A(n1675), .Z(n1888) );
  XNOR U1816 ( .A(n1891), .B(n1892), .Z(out[77]) );
  XOR U1817 ( .A(n1895), .B(n1466), .Z(out[779]) );
  IV U1818 ( .A(n1679), .Z(n1466) );
  XNOR U1819 ( .A(round_reg[754]), .B(n1896), .Z(n1679) );
  ANDN U1820 ( .B(n1897), .A(n1678), .Z(n1895) );
  XOR U1821 ( .A(n1898), .B(n1470), .Z(out[778]) );
  IV U1822 ( .A(n1682), .Z(n1470) );
  XNOR U1823 ( .A(round_reg[753]), .B(n1899), .Z(n1682) );
  ANDN U1824 ( .B(n1900), .A(n1681), .Z(n1898) );
  XOR U1825 ( .A(n1901), .B(n1474), .Z(out[777]) );
  IV U1826 ( .A(n1685), .Z(n1474) );
  XNOR U1827 ( .A(round_reg[752]), .B(n1902), .Z(n1685) );
  ANDN U1828 ( .B(n1903), .A(n1684), .Z(n1901) );
  XOR U1829 ( .A(n1904), .B(n1478), .Z(out[776]) );
  IV U1830 ( .A(n1688), .Z(n1478) );
  XNOR U1831 ( .A(round_reg[751]), .B(n1905), .Z(n1688) );
  ANDN U1832 ( .B(n1906), .A(n1687), .Z(n1904) );
  XOR U1833 ( .A(n1907), .B(n1482), .Z(out[775]) );
  IV U1834 ( .A(n1695), .Z(n1482) );
  XNOR U1835 ( .A(round_reg[750]), .B(n1908), .Z(n1695) );
  XOR U1836 ( .A(n1910), .B(n1486), .Z(out[774]) );
  IV U1837 ( .A(n1698), .Z(n1486) );
  XNOR U1838 ( .A(round_reg[749]), .B(n1911), .Z(n1698) );
  ANDN U1839 ( .B(n1912), .A(n1697), .Z(n1910) );
  XOR U1840 ( .A(n1913), .B(n1490), .Z(out[773]) );
  XNOR U1841 ( .A(round_reg[748]), .B(n1914), .Z(n1490) );
  ANDN U1842 ( .B(n1915), .A(n1700), .Z(n1913) );
  XOR U1843 ( .A(n1916), .B(n1494), .Z(out[772]) );
  XNOR U1844 ( .A(round_reg[747]), .B(n1917), .Z(n1494) );
  ANDN U1845 ( .B(n1918), .A(n1702), .Z(n1916) );
  XOR U1846 ( .A(n1919), .B(n1506), .Z(out[771]) );
  XNOR U1847 ( .A(round_reg[746]), .B(n1920), .Z(n1506) );
  ANDN U1848 ( .B(n1921), .A(n1704), .Z(n1919) );
  XOR U1849 ( .A(n1922), .B(n1510), .Z(out[770]) );
  XNOR U1850 ( .A(round_reg[745]), .B(n1923), .Z(n1510) );
  ANDN U1851 ( .B(n1924), .A(n1706), .Z(n1922) );
  XNOR U1852 ( .A(n1925), .B(n1926), .Z(out[76]) );
  XOR U1853 ( .A(n1929), .B(n1514), .Z(out[769]) );
  XNOR U1854 ( .A(round_reg[744]), .B(n1930), .Z(n1514) );
  ANDN U1855 ( .B(n1931), .A(n1708), .Z(n1929) );
  XOR U1856 ( .A(n1932), .B(n1518), .Z(out[768]) );
  XNOR U1857 ( .A(round_reg[743]), .B(n1933), .Z(n1518) );
  XOR U1858 ( .A(n1935), .B(n1520), .Z(out[767]) );
  XOR U1859 ( .A(round_reg[375]), .B(n1936), .Z(n1520) );
  ANDN U1860 ( .B(n1236), .A(n1713), .Z(n1935) );
  XOR U1861 ( .A(n1937), .B(n1522), .Z(out[766]) );
  XOR U1862 ( .A(round_reg[374]), .B(n1938), .Z(n1522) );
  ANDN U1863 ( .B(n1240), .A(n1716), .Z(n1937) );
  XOR U1864 ( .A(n1939), .B(n1524), .Z(out[765]) );
  XOR U1865 ( .A(round_reg[373]), .B(n1940), .Z(n1524) );
  XOR U1866 ( .A(n1941), .B(n1526), .Z(out[764]) );
  XOR U1867 ( .A(round_reg[372]), .B(n1942), .Z(n1526) );
  AND U1868 ( .A(n1248), .B(n1726), .Z(n1941) );
  IV U1869 ( .A(n1943), .Z(n1726) );
  XOR U1870 ( .A(n1944), .B(n1528), .Z(out[763]) );
  XOR U1871 ( .A(round_reg[371]), .B(n1945), .Z(n1528) );
  AND U1872 ( .A(n1252), .B(n1729), .Z(n1944) );
  IV U1873 ( .A(n1946), .Z(n1729) );
  XOR U1874 ( .A(n1947), .B(n1531), .Z(out[762]) );
  XOR U1875 ( .A(round_reg[370]), .B(n1948), .Z(n1531) );
  ANDN U1876 ( .B(n1732), .A(n1256), .Z(n1947) );
  IV U1877 ( .A(n1949), .Z(n1732) );
  XOR U1878 ( .A(n1950), .B(n1538), .Z(out[761]) );
  XOR U1879 ( .A(round_reg[369]), .B(n1951), .Z(n1538) );
  ANDN U1880 ( .B(n1735), .A(n1260), .Z(n1950) );
  IV U1881 ( .A(n1952), .Z(n1735) );
  XOR U1882 ( .A(n1953), .B(n1541), .Z(out[760]) );
  XOR U1883 ( .A(round_reg[368]), .B(n1954), .Z(n1541) );
  ANDN U1884 ( .B(n1738), .A(n1264), .Z(n1953) );
  IV U1885 ( .A(n1955), .Z(n1738) );
  XNOR U1886 ( .A(n1956), .B(n1957), .Z(out[75]) );
  XOR U1887 ( .A(n1960), .B(n1544), .Z(out[759]) );
  XOR U1888 ( .A(round_reg[367]), .B(n1961), .Z(n1544) );
  ANDN U1889 ( .B(n1741), .A(n1268), .Z(n1960) );
  IV U1890 ( .A(n1962), .Z(n1741) );
  XOR U1891 ( .A(n1963), .B(n1547), .Z(out[758]) );
  XOR U1892 ( .A(round_reg[366]), .B(n1964), .Z(n1547) );
  ANDN U1893 ( .B(n1744), .A(n1272), .Z(n1963) );
  IV U1894 ( .A(n1965), .Z(n1744) );
  XOR U1895 ( .A(n1966), .B(n1550), .Z(out[757]) );
  XOR U1896 ( .A(round_reg[365]), .B(n1967), .Z(n1550) );
  ANDN U1897 ( .B(n1747), .A(n1280), .Z(n1966) );
  IV U1898 ( .A(n1968), .Z(n1747) );
  XOR U1899 ( .A(n1969), .B(n1553), .Z(out[756]) );
  XOR U1900 ( .A(round_reg[364]), .B(n1970), .Z(n1553) );
  ANDN U1901 ( .B(n1750), .A(n1284), .Z(n1969) );
  IV U1902 ( .A(n1971), .Z(n1750) );
  XOR U1903 ( .A(n1972), .B(n1556), .Z(out[755]) );
  XOR U1904 ( .A(round_reg[363]), .B(n1973), .Z(n1556) );
  XOR U1905 ( .A(n1974), .B(n1558), .Z(out[754]) );
  XOR U1906 ( .A(round_reg[362]), .B(n1975), .Z(n1558) );
  XOR U1907 ( .A(n1976), .B(n1560), .Z(out[753]) );
  XOR U1908 ( .A(round_reg[361]), .B(n1977), .Z(n1560) );
  ANDN U1909 ( .B(n1763), .A(n1296), .Z(n1976) );
  IV U1910 ( .A(n1978), .Z(n1763) );
  XOR U1911 ( .A(n1979), .B(n1562), .Z(out[752]) );
  XOR U1912 ( .A(round_reg[360]), .B(n1980), .Z(n1562) );
  ANDN U1913 ( .B(n1766), .A(n1300), .Z(n1979) );
  IV U1914 ( .A(n1981), .Z(n1766) );
  XOR U1915 ( .A(n1982), .B(n1568), .Z(out[751]) );
  XOR U1916 ( .A(round_reg[359]), .B(n1983), .Z(n1568) );
  ANDN U1917 ( .B(n1769), .A(n1304), .Z(n1982) );
  IV U1918 ( .A(n1984), .Z(n1769) );
  XOR U1919 ( .A(n1985), .B(n1570), .Z(out[750]) );
  XOR U1920 ( .A(round_reg[358]), .B(n1986), .Z(n1570) );
  ANDN U1921 ( .B(n1772), .A(n1308), .Z(n1985) );
  IV U1922 ( .A(n1987), .Z(n1772) );
  XNOR U1923 ( .A(n1988), .B(n1989), .Z(out[74]) );
  XOR U1924 ( .A(n1992), .B(n1572), .Z(out[749]) );
  XOR U1925 ( .A(round_reg[357]), .B(n1993), .Z(n1572) );
  ANDN U1926 ( .B(n1775), .A(n1312), .Z(n1992) );
  IV U1927 ( .A(n1994), .Z(n1775) );
  XOR U1928 ( .A(n1995), .B(n1574), .Z(out[748]) );
  XOR U1929 ( .A(round_reg[356]), .B(n1996), .Z(n1574) );
  ANDN U1930 ( .B(n1778), .A(n1316), .Z(n1995) );
  IV U1931 ( .A(n1997), .Z(n1778) );
  XOR U1932 ( .A(n1998), .B(n1576), .Z(out[747]) );
  XOR U1933 ( .A(round_reg[355]), .B(n1999), .Z(n1576) );
  ANDN U1934 ( .B(n1781), .A(n1324), .Z(n1998) );
  IV U1935 ( .A(n2000), .Z(n1781) );
  XOR U1936 ( .A(n2001), .B(n1579), .Z(out[746]) );
  XOR U1937 ( .A(round_reg[354]), .B(n2002), .Z(n1579) );
  XOR U1938 ( .A(n2003), .B(n1581), .Z(out[745]) );
  XOR U1939 ( .A(round_reg[353]), .B(n2004), .Z(n1581) );
  XOR U1940 ( .A(n2005), .B(n1583), .Z(out[744]) );
  XOR U1941 ( .A(round_reg[352]), .B(n2006), .Z(n1583) );
  XOR U1942 ( .A(n2007), .B(n1585), .Z(out[743]) );
  XOR U1943 ( .A(round_reg[351]), .B(n2008), .Z(n1585) );
  XOR U1944 ( .A(n2009), .B(n1587), .Z(out[742]) );
  XOR U1945 ( .A(round_reg[350]), .B(n2010), .Z(n1587) );
  XOR U1946 ( .A(n2011), .B(n1593), .Z(out[741]) );
  XOR U1947 ( .A(round_reg[349]), .B(n2012), .Z(n1593) );
  XOR U1948 ( .A(n2013), .B(n1595), .Z(out[740]) );
  XOR U1949 ( .A(round_reg[348]), .B(n2014), .Z(n1595) );
  ANDN U1950 ( .B(n1806), .A(n1352), .Z(n2013) );
  IV U1951 ( .A(n2015), .Z(n1806) );
  XNOR U1952 ( .A(n2016), .B(n2017), .Z(out[73]) );
  AND U1953 ( .A(n1054), .B(n2018), .Z(n2016) );
  XOR U1954 ( .A(n2019), .B(n1598), .Z(out[739]) );
  XOR U1955 ( .A(round_reg[347]), .B(n2020), .Z(n1598) );
  NOR U1956 ( .A(n1809), .B(n1356), .Z(n2019) );
  XOR U1957 ( .A(n2021), .B(n1601), .Z(out[738]) );
  XOR U1958 ( .A(round_reg[346]), .B(n2022), .Z(n1601) );
  ANDN U1959 ( .B(n1812), .A(n1360), .Z(n2021) );
  IV U1960 ( .A(n2023), .Z(n1812) );
  XOR U1961 ( .A(n2024), .B(n1604), .Z(out[737]) );
  XOR U1962 ( .A(round_reg[345]), .B(n2025), .Z(n1604) );
  ANDN U1963 ( .B(n1815), .A(n1368), .Z(n2024) );
  IV U1964 ( .A(n2026), .Z(n1815) );
  XOR U1965 ( .A(n2027), .B(n1607), .Z(out[736]) );
  XOR U1966 ( .A(round_reg[344]), .B(n2028), .Z(n1607) );
  ANDN U1967 ( .B(n1818), .A(n1372), .Z(n2027) );
  IV U1968 ( .A(n2029), .Z(n1818) );
  XOR U1969 ( .A(n2030), .B(n1610), .Z(out[735]) );
  XOR U1970 ( .A(round_reg[343]), .B(n2031), .Z(n1610) );
  ANDN U1971 ( .B(n1829), .A(n1376), .Z(n2030) );
  IV U1972 ( .A(n2032), .Z(n1829) );
  XOR U1973 ( .A(n2033), .B(n1613), .Z(out[734]) );
  XOR U1974 ( .A(round_reg[342]), .B(n2034), .Z(n1613) );
  ANDN U1975 ( .B(n1832), .A(n1380), .Z(n2033) );
  IV U1976 ( .A(n2035), .Z(n1832) );
  XOR U1977 ( .A(n2036), .B(n1616), .Z(out[733]) );
  XOR U1978 ( .A(round_reg[341]), .B(n2037), .Z(n1616) );
  ANDN U1979 ( .B(n1835), .A(n1384), .Z(n2036) );
  IV U1980 ( .A(n2038), .Z(n1835) );
  XOR U1981 ( .A(n2039), .B(n1619), .Z(out[732]) );
  XOR U1982 ( .A(round_reg[340]), .B(n2040), .Z(n1619) );
  NOR U1983 ( .A(n1838), .B(n1388), .Z(n2039) );
  XOR U1984 ( .A(n2041), .B(n1626), .Z(out[731]) );
  XOR U1985 ( .A(round_reg[339]), .B(n2042), .Z(n1626) );
  NOR U1986 ( .A(n1841), .B(n1392), .Z(n2041) );
  XOR U1987 ( .A(n2043), .B(n1629), .Z(out[730]) );
  XOR U1988 ( .A(round_reg[338]), .B(n2044), .Z(n1629) );
  NOR U1989 ( .A(n1844), .B(n1396), .Z(n2043) );
  XNOR U1990 ( .A(n2045), .B(n2046), .Z(out[72]) );
  AND U1991 ( .A(n1498), .B(n1496), .Z(n2045) );
  XOR U1992 ( .A(n2047), .B(n1632), .Z(out[729]) );
  XOR U1993 ( .A(round_reg[337]), .B(n2048), .Z(n1632) );
  NOR U1994 ( .A(n1847), .B(n1400), .Z(n2047) );
  XOR U1995 ( .A(n2049), .B(n1635), .Z(out[728]) );
  XOR U1996 ( .A(round_reg[336]), .B(n2050), .Z(n1635) );
  NOR U1997 ( .A(n1850), .B(n1404), .Z(n2049) );
  XOR U1998 ( .A(n2051), .B(n1638), .Z(out[727]) );
  XOR U1999 ( .A(round_reg[335]), .B(n2052), .Z(n1638) );
  NOR U2000 ( .A(n1853), .B(n1412), .Z(n2051) );
  XOR U2001 ( .A(n2053), .B(n1641), .Z(out[726]) );
  XOR U2002 ( .A(round_reg[334]), .B(n2054), .Z(n1641) );
  NOR U2003 ( .A(n1856), .B(n1416), .Z(n2053) );
  XOR U2004 ( .A(n2055), .B(n1644), .Z(out[725]) );
  XOR U2005 ( .A(round_reg[333]), .B(n2056), .Z(n1644) );
  NOR U2006 ( .A(n1863), .B(n1420), .Z(n2055) );
  XOR U2007 ( .A(n2057), .B(n1647), .Z(out[724]) );
  XOR U2008 ( .A(round_reg[332]), .B(n2058), .Z(n1647) );
  NOR U2009 ( .A(n1866), .B(n1424), .Z(n2057) );
  XOR U2010 ( .A(n2059), .B(n1650), .Z(out[723]) );
  XOR U2011 ( .A(round_reg[331]), .B(n2060), .Z(n1650) );
  NOR U2012 ( .A(n1869), .B(n1428), .Z(n2059) );
  XOR U2013 ( .A(n2061), .B(n1653), .Z(out[722]) );
  XOR U2014 ( .A(round_reg[330]), .B(n2062), .Z(n1653) );
  NOR U2015 ( .A(n1872), .B(n1432), .Z(n2061) );
  XOR U2016 ( .A(n2063), .B(n1660), .Z(out[721]) );
  XOR U2017 ( .A(round_reg[329]), .B(n2064), .Z(n1660) );
  NOR U2018 ( .A(n1875), .B(n1436), .Z(n2063) );
  XOR U2019 ( .A(n2065), .B(n1663), .Z(out[720]) );
  XOR U2020 ( .A(round_reg[328]), .B(n2066), .Z(n1663) );
  NOR U2021 ( .A(n1878), .B(n1440), .Z(n2065) );
  XNOR U2022 ( .A(n2067), .B(n2068), .Z(out[71]) );
  AND U2023 ( .A(n1822), .B(n1820), .Z(n2067) );
  XOR U2024 ( .A(n2069), .B(n1666), .Z(out[719]) );
  XOR U2025 ( .A(round_reg[327]), .B(n2070), .Z(n1666) );
  NOR U2026 ( .A(n1881), .B(n1444), .Z(n2069) );
  XOR U2027 ( .A(n2071), .B(n1669), .Z(out[718]) );
  XOR U2028 ( .A(round_reg[326]), .B(n2072), .Z(n1669) );
  NOR U2029 ( .A(n1884), .B(n1448), .Z(n2071) );
  XOR U2030 ( .A(n2073), .B(n1672), .Z(out[717]) );
  XOR U2031 ( .A(round_reg[325]), .B(n2074), .Z(n1672) );
  NOR U2032 ( .A(n1887), .B(n1456), .Z(n2073) );
  XOR U2033 ( .A(n2075), .B(n1675), .Z(out[716]) );
  XOR U2034 ( .A(round_reg[324]), .B(n2076), .Z(n1675) );
  NOR U2035 ( .A(n1890), .B(n1460), .Z(n2075) );
  XOR U2036 ( .A(n2077), .B(n1678), .Z(out[715]) );
  XOR U2037 ( .A(round_reg[323]), .B(n2078), .Z(n1678) );
  NOR U2038 ( .A(n1897), .B(n1464), .Z(n2077) );
  XOR U2039 ( .A(n2079), .B(n1681), .Z(out[714]) );
  XOR U2040 ( .A(round_reg[322]), .B(n2080), .Z(n1681) );
  NOR U2041 ( .A(n1900), .B(n1468), .Z(n2079) );
  XOR U2042 ( .A(n2081), .B(n1684), .Z(out[713]) );
  XOR U2043 ( .A(round_reg[321]), .B(n2082), .Z(n1684) );
  NOR U2044 ( .A(n1903), .B(n1472), .Z(n2081) );
  XOR U2045 ( .A(n2083), .B(n1687), .Z(out[712]) );
  XOR U2046 ( .A(round_reg[320]), .B(n2084), .Z(n1687) );
  NOR U2047 ( .A(n1906), .B(n1476), .Z(n2083) );
  XOR U2048 ( .A(n2085), .B(n1694), .Z(out[711]) );
  XNOR U2049 ( .A(round_reg[383]), .B(n2086), .Z(n1694) );
  NOR U2050 ( .A(n1909), .B(n1480), .Z(n2085) );
  XOR U2051 ( .A(n2087), .B(n1697), .Z(out[710]) );
  XOR U2052 ( .A(round_reg[382]), .B(n2088), .Z(n1697) );
  NOR U2053 ( .A(n1912), .B(n1484), .Z(n2087) );
  XNOR U2054 ( .A(n2089), .B(n2090), .Z(out[70]) );
  AND U2055 ( .A(n2091), .B(n2092), .Z(n2089) );
  XOR U2056 ( .A(n2093), .B(n1700), .Z(out[709]) );
  XOR U2057 ( .A(round_reg[381]), .B(n2094), .Z(n1700) );
  NOR U2058 ( .A(n1915), .B(n1488), .Z(n2093) );
  XOR U2059 ( .A(n2095), .B(n1702), .Z(out[708]) );
  XOR U2060 ( .A(round_reg[380]), .B(n2096), .Z(n1702) );
  NOR U2061 ( .A(n1918), .B(n1492), .Z(n2095) );
  XOR U2062 ( .A(n2097), .B(n1704), .Z(out[707]) );
  XOR U2063 ( .A(round_reg[379]), .B(n2098), .Z(n1704) );
  NOR U2064 ( .A(n1921), .B(n1504), .Z(n2097) );
  XOR U2065 ( .A(n2099), .B(n1706), .Z(out[706]) );
  XOR U2066 ( .A(round_reg[378]), .B(n2100), .Z(n1706) );
  NOR U2067 ( .A(n1924), .B(n1508), .Z(n2099) );
  XOR U2068 ( .A(n2101), .B(n1708), .Z(out[705]) );
  XOR U2069 ( .A(round_reg[377]), .B(n2102), .Z(n1708) );
  NOR U2070 ( .A(n1931), .B(n1512), .Z(n2101) );
  XOR U2071 ( .A(n2103), .B(n1710), .Z(out[704]) );
  XOR U2072 ( .A(round_reg[376]), .B(n2104), .Z(n1710) );
  NOR U2073 ( .A(n1934), .B(n1516), .Z(n2103) );
  XOR U2074 ( .A(n2105), .B(n1713), .Z(out[703]) );
  XOR U2075 ( .A(round_reg[301]), .B(n2106), .Z(n1713) );
  NOR U2076 ( .A(n1237), .B(n1236), .Z(n2105) );
  XNOR U2077 ( .A(round_reg[1534]), .B(n2107), .Z(n1236) );
  XNOR U2078 ( .A(round_reg[1145]), .B(n2108), .Z(n1237) );
  XOR U2079 ( .A(n2109), .B(n1716), .Z(out[702]) );
  XOR U2080 ( .A(round_reg[300]), .B(n2110), .Z(n1716) );
  NOR U2081 ( .A(n1241), .B(n1240), .Z(n2109) );
  XNOR U2082 ( .A(round_reg[1533]), .B(n2111), .Z(n1240) );
  XNOR U2083 ( .A(round_reg[1144]), .B(n2112), .Z(n1241) );
  XOR U2084 ( .A(n2113), .B(n1723), .Z(out[701]) );
  XOR U2085 ( .A(round_reg[299]), .B(n2114), .Z(n1723) );
  NOR U2086 ( .A(n1245), .B(n1244), .Z(n2113) );
  XOR U2087 ( .A(round_reg[1532]), .B(n2115), .Z(n1244) );
  XNOR U2088 ( .A(round_reg[1143]), .B(n2116), .Z(n1245) );
  XOR U2089 ( .A(n2117), .B(n1943), .Z(out[700]) );
  XOR U2090 ( .A(round_reg[298]), .B(n2118), .Z(n1943) );
  NOR U2091 ( .A(n1249), .B(n1248), .Z(n2117) );
  XOR U2092 ( .A(round_reg[1531]), .B(n2119), .Z(n1248) );
  XNOR U2093 ( .A(round_reg[1142]), .B(n2120), .Z(n1249) );
  XNOR U2094 ( .A(n2121), .B(n2091), .Z(out[6]) );
  AND U2095 ( .A(n2122), .B(n2123), .Z(n2121) );
  XNOR U2096 ( .A(n2124), .B(n2125), .Z(out[69]) );
  AND U2097 ( .A(n2126), .B(n2127), .Z(n2124) );
  XOR U2098 ( .A(n2128), .B(n1946), .Z(out[699]) );
  XOR U2099 ( .A(round_reg[297]), .B(n2129), .Z(n1946) );
  NOR U2100 ( .A(n1253), .B(n1252), .Z(n2128) );
  XNOR U2101 ( .A(round_reg[1530]), .B(n2130), .Z(n1252) );
  XNOR U2102 ( .A(round_reg[1141]), .B(n2131), .Z(n1253) );
  XOR U2103 ( .A(n2132), .B(n1949), .Z(out[698]) );
  XOR U2104 ( .A(round_reg[296]), .B(n2133), .Z(n1949) );
  ANDN U2105 ( .B(n1256), .A(n1257), .Z(n2132) );
  XNOR U2106 ( .A(round_reg[1140]), .B(n2134), .Z(n1257) );
  XNOR U2107 ( .A(round_reg[1529]), .B(n2135), .Z(n1256) );
  XOR U2108 ( .A(n2136), .B(n1952), .Z(out[697]) );
  XOR U2109 ( .A(round_reg[295]), .B(n2137), .Z(n1952) );
  ANDN U2110 ( .B(n1260), .A(n1261), .Z(n2136) );
  XNOR U2111 ( .A(round_reg[1139]), .B(n2138), .Z(n1261) );
  XNOR U2112 ( .A(round_reg[1528]), .B(n2139), .Z(n1260) );
  XOR U2113 ( .A(n2140), .B(n1955), .Z(out[696]) );
  XOR U2114 ( .A(round_reg[294]), .B(n2141), .Z(n1955) );
  ANDN U2115 ( .B(n1264), .A(n1265), .Z(n2140) );
  XNOR U2116 ( .A(round_reg[1138]), .B(n2142), .Z(n1265) );
  XNOR U2117 ( .A(round_reg[1527]), .B(n2143), .Z(n1264) );
  XOR U2118 ( .A(n2144), .B(n1962), .Z(out[695]) );
  XOR U2119 ( .A(round_reg[293]), .B(n2145), .Z(n1962) );
  ANDN U2120 ( .B(n1268), .A(n1269), .Z(n2144) );
  XNOR U2121 ( .A(round_reg[1137]), .B(n2146), .Z(n1269) );
  XNOR U2122 ( .A(round_reg[1526]), .B(n2147), .Z(n1268) );
  XOR U2123 ( .A(n2148), .B(n1965), .Z(out[694]) );
  XOR U2124 ( .A(round_reg[292]), .B(n2149), .Z(n1965) );
  ANDN U2125 ( .B(n1272), .A(n1273), .Z(n2148) );
  XNOR U2126 ( .A(round_reg[1136]), .B(n2150), .Z(n1273) );
  XNOR U2127 ( .A(round_reg[1525]), .B(n2151), .Z(n1272) );
  XOR U2128 ( .A(n2152), .B(n1968), .Z(out[693]) );
  XOR U2129 ( .A(round_reg[291]), .B(n2153), .Z(n1968) );
  ANDN U2130 ( .B(n1280), .A(n1281), .Z(n2152) );
  XNOR U2131 ( .A(round_reg[1135]), .B(n2154), .Z(n1281) );
  XNOR U2132 ( .A(round_reg[1524]), .B(n2155), .Z(n1280) );
  XOR U2133 ( .A(n2156), .B(n1971), .Z(out[692]) );
  XOR U2134 ( .A(round_reg[290]), .B(n2157), .Z(n1971) );
  ANDN U2135 ( .B(n1284), .A(n1285), .Z(n2156) );
  XNOR U2136 ( .A(round_reg[1134]), .B(n2158), .Z(n1285) );
  XNOR U2137 ( .A(round_reg[1523]), .B(n2159), .Z(n1284) );
  XOR U2138 ( .A(n2160), .B(n1757), .Z(out[691]) );
  XOR U2139 ( .A(round_reg[289]), .B(n2161), .Z(n1757) );
  ANDN U2140 ( .B(n1288), .A(n1289), .Z(n2160) );
  XNOR U2141 ( .A(round_reg[1133]), .B(n2162), .Z(n1289) );
  XNOR U2142 ( .A(round_reg[1522]), .B(n2163), .Z(n1288) );
  XOR U2143 ( .A(n2164), .B(n1760), .Z(out[690]) );
  XOR U2144 ( .A(round_reg[288]), .B(n2165), .Z(n1760) );
  ANDN U2145 ( .B(n1292), .A(n1293), .Z(n2164) );
  XNOR U2146 ( .A(round_reg[1132]), .B(n2166), .Z(n1293) );
  XNOR U2147 ( .A(round_reg[1521]), .B(n2167), .Z(n1292) );
  XNOR U2148 ( .A(n2168), .B(n2169), .Z(out[68]) );
  AND U2149 ( .A(n2170), .B(n2171), .Z(n2168) );
  XOR U2150 ( .A(n2172), .B(n1978), .Z(out[689]) );
  XOR U2151 ( .A(round_reg[287]), .B(n2173), .Z(n1978) );
  ANDN U2152 ( .B(n1296), .A(n1297), .Z(n2172) );
  XNOR U2153 ( .A(round_reg[1131]), .B(n2174), .Z(n1297) );
  XNOR U2154 ( .A(round_reg[1520]), .B(n2175), .Z(n1296) );
  XOR U2155 ( .A(n2176), .B(n1981), .Z(out[688]) );
  XOR U2156 ( .A(round_reg[286]), .B(n2177), .Z(n1981) );
  ANDN U2157 ( .B(n1300), .A(n1301), .Z(n2176) );
  XNOR U2158 ( .A(round_reg[1130]), .B(n2178), .Z(n1301) );
  XNOR U2159 ( .A(round_reg[1519]), .B(n2179), .Z(n1300) );
  XOR U2160 ( .A(n2180), .B(n1984), .Z(out[687]) );
  XOR U2161 ( .A(round_reg[285]), .B(n2181), .Z(n1984) );
  ANDN U2162 ( .B(n1304), .A(n1305), .Z(n2180) );
  XNOR U2163 ( .A(round_reg[1129]), .B(n2182), .Z(n1305) );
  XNOR U2164 ( .A(round_reg[1518]), .B(n2183), .Z(n1304) );
  XOR U2165 ( .A(n2184), .B(n1987), .Z(out[686]) );
  XOR U2166 ( .A(round_reg[284]), .B(n2185), .Z(n1987) );
  ANDN U2167 ( .B(n1308), .A(n1309), .Z(n2184) );
  XNOR U2168 ( .A(round_reg[1128]), .B(n2186), .Z(n1309) );
  XNOR U2169 ( .A(round_reg[1517]), .B(n2187), .Z(n1308) );
  XOR U2170 ( .A(n2188), .B(n1994), .Z(out[685]) );
  XOR U2171 ( .A(round_reg[283]), .B(n2189), .Z(n1994) );
  ANDN U2172 ( .B(n1312), .A(n1313), .Z(n2188) );
  XNOR U2173 ( .A(round_reg[1127]), .B(n2190), .Z(n1313) );
  XNOR U2174 ( .A(round_reg[1516]), .B(n2191), .Z(n1312) );
  XOR U2175 ( .A(n2192), .B(n1997), .Z(out[684]) );
  XOR U2176 ( .A(round_reg[282]), .B(n2193), .Z(n1997) );
  ANDN U2177 ( .B(n1316), .A(n1317), .Z(n2192) );
  XNOR U2178 ( .A(round_reg[1126]), .B(n2194), .Z(n1317) );
  XNOR U2179 ( .A(round_reg[1515]), .B(n2195), .Z(n1316) );
  XOR U2180 ( .A(n2196), .B(n2000), .Z(out[683]) );
  XOR U2181 ( .A(round_reg[281]), .B(n2197), .Z(n2000) );
  ANDN U2182 ( .B(n1324), .A(n1325), .Z(n2196) );
  XNOR U2183 ( .A(round_reg[1125]), .B(n2198), .Z(n1325) );
  XNOR U2184 ( .A(round_reg[1514]), .B(n2199), .Z(n1324) );
  XOR U2185 ( .A(n2200), .B(n1784), .Z(out[682]) );
  XOR U2186 ( .A(round_reg[280]), .B(n2201), .Z(n1784) );
  ANDN U2187 ( .B(n1328), .A(n1329), .Z(n2200) );
  XNOR U2188 ( .A(round_reg[1124]), .B(n2202), .Z(n1329) );
  XNOR U2189 ( .A(round_reg[1513]), .B(n2203), .Z(n1328) );
  XOR U2190 ( .A(n2204), .B(n1791), .Z(out[681]) );
  XOR U2191 ( .A(round_reg[279]), .B(n2205), .Z(n1791) );
  ANDN U2192 ( .B(n1332), .A(n1333), .Z(n2204) );
  XNOR U2193 ( .A(round_reg[1123]), .B(n2206), .Z(n1333) );
  XNOR U2194 ( .A(round_reg[1512]), .B(n2207), .Z(n1332) );
  XOR U2195 ( .A(n2208), .B(n1794), .Z(out[680]) );
  XOR U2196 ( .A(round_reg[278]), .B(n2209), .Z(n1794) );
  ANDN U2197 ( .B(n1336), .A(n1337), .Z(n2208) );
  XNOR U2198 ( .A(round_reg[1122]), .B(n2210), .Z(n1337) );
  XNOR U2199 ( .A(round_reg[1511]), .B(n2211), .Z(n1336) );
  XNOR U2200 ( .A(n2212), .B(n2213), .Z(out[67]) );
  AND U2201 ( .A(n2214), .B(n2215), .Z(n2212) );
  XOR U2202 ( .A(n2216), .B(n1797), .Z(out[679]) );
  XOR U2203 ( .A(round_reg[277]), .B(n2217), .Z(n1797) );
  ANDN U2204 ( .B(n1340), .A(n1341), .Z(n2216) );
  XNOR U2205 ( .A(round_reg[1121]), .B(n2218), .Z(n1341) );
  XNOR U2206 ( .A(round_reg[1510]), .B(n2219), .Z(n1340) );
  XOR U2207 ( .A(n2220), .B(n1800), .Z(out[678]) );
  XOR U2208 ( .A(round_reg[276]), .B(n2221), .Z(n1800) );
  ANDN U2209 ( .B(n1344), .A(n1345), .Z(n2220) );
  XNOR U2210 ( .A(round_reg[1120]), .B(n2222), .Z(n1345) );
  XNOR U2211 ( .A(round_reg[1509]), .B(n2223), .Z(n1344) );
  XOR U2212 ( .A(n2224), .B(n1803), .Z(out[677]) );
  XOR U2213 ( .A(round_reg[275]), .B(n2225), .Z(n1803) );
  ANDN U2214 ( .B(n1348), .A(n1349), .Z(n2224) );
  XNOR U2215 ( .A(round_reg[1119]), .B(n2226), .Z(n1349) );
  XNOR U2216 ( .A(round_reg[1508]), .B(n2227), .Z(n1348) );
  XOR U2217 ( .A(n2228), .B(n2015), .Z(out[676]) );
  XOR U2218 ( .A(round_reg[274]), .B(n2229), .Z(n2015) );
  ANDN U2219 ( .B(n1352), .A(n1353), .Z(n2228) );
  XNOR U2220 ( .A(round_reg[1118]), .B(n2230), .Z(n1353) );
  XNOR U2221 ( .A(round_reg[1507]), .B(n2231), .Z(n1352) );
  XOR U2222 ( .A(n2232), .B(n1809), .Z(out[675]) );
  XOR U2223 ( .A(round_reg[273]), .B(n2233), .Z(n1809) );
  ANDN U2224 ( .B(n1356), .A(n1357), .Z(n2232) );
  XNOR U2225 ( .A(round_reg[1117]), .B(n2234), .Z(n1357) );
  XNOR U2226 ( .A(round_reg[1506]), .B(n2235), .Z(n1356) );
  XOR U2227 ( .A(n2236), .B(n2023), .Z(out[674]) );
  XOR U2228 ( .A(round_reg[272]), .B(n2237), .Z(n2023) );
  ANDN U2229 ( .B(n1360), .A(n1361), .Z(n2236) );
  XNOR U2230 ( .A(round_reg[1116]), .B(n2238), .Z(n1361) );
  XNOR U2231 ( .A(round_reg[1505]), .B(n2239), .Z(n1360) );
  XOR U2232 ( .A(n2240), .B(n2026), .Z(out[673]) );
  XOR U2233 ( .A(round_reg[271]), .B(n2241), .Z(n2026) );
  ANDN U2234 ( .B(n1368), .A(n1369), .Z(n2240) );
  XNOR U2235 ( .A(round_reg[1115]), .B(n2242), .Z(n1369) );
  XOR U2236 ( .A(round_reg[1504]), .B(n2243), .Z(n1368) );
  XOR U2237 ( .A(n2244), .B(n2029), .Z(out[672]) );
  XOR U2238 ( .A(round_reg[270]), .B(n2245), .Z(n2029) );
  ANDN U2239 ( .B(n1372), .A(n1373), .Z(n2244) );
  XNOR U2240 ( .A(round_reg[1114]), .B(n2246), .Z(n1373) );
  XOR U2241 ( .A(round_reg[1503]), .B(n2247), .Z(n1372) );
  XOR U2242 ( .A(n2248), .B(n2032), .Z(out[671]) );
  XOR U2243 ( .A(round_reg[269]), .B(n2249), .Z(n2032) );
  ANDN U2244 ( .B(n1376), .A(n1377), .Z(n2248) );
  XNOR U2245 ( .A(round_reg[1113]), .B(n2250), .Z(n1377) );
  XOR U2246 ( .A(round_reg[1502]), .B(n2251), .Z(n1376) );
  XOR U2247 ( .A(n2252), .B(n2035), .Z(out[670]) );
  XOR U2248 ( .A(round_reg[268]), .B(n2253), .Z(n2035) );
  ANDN U2249 ( .B(n1380), .A(n1381), .Z(n2252) );
  XNOR U2250 ( .A(round_reg[1112]), .B(n2254), .Z(n1381) );
  XOR U2251 ( .A(round_reg[1501]), .B(n2255), .Z(n1380) );
  XNOR U2252 ( .A(n2256), .B(n2257), .Z(out[66]) );
  AND U2253 ( .A(n2258), .B(n2259), .Z(n2256) );
  XOR U2254 ( .A(n2260), .B(n2038), .Z(out[669]) );
  XOR U2255 ( .A(round_reg[267]), .B(n2261), .Z(n2038) );
  ANDN U2256 ( .B(n1384), .A(n1385), .Z(n2260) );
  XNOR U2257 ( .A(round_reg[1111]), .B(n2262), .Z(n1385) );
  XOR U2258 ( .A(round_reg[1500]), .B(n2263), .Z(n1384) );
  XOR U2259 ( .A(n2264), .B(n1838), .Z(out[668]) );
  XOR U2260 ( .A(round_reg[266]), .B(n2265), .Z(n1838) );
  ANDN U2261 ( .B(n1388), .A(n1389), .Z(n2264) );
  XNOR U2262 ( .A(round_reg[1110]), .B(n2266), .Z(n1389) );
  XNOR U2263 ( .A(round_reg[1499]), .B(n2267), .Z(n1388) );
  XOR U2264 ( .A(n2268), .B(n1841), .Z(out[667]) );
  XOR U2265 ( .A(round_reg[265]), .B(n2269), .Z(n1841) );
  ANDN U2266 ( .B(n1392), .A(n1393), .Z(n2268) );
  XNOR U2267 ( .A(round_reg[1109]), .B(n2270), .Z(n1393) );
  XNOR U2268 ( .A(round_reg[1498]), .B(n2271), .Z(n1392) );
  XOR U2269 ( .A(n2272), .B(n1844), .Z(out[666]) );
  XOR U2270 ( .A(round_reg[264]), .B(n2273), .Z(n1844) );
  ANDN U2271 ( .B(n1396), .A(n1397), .Z(n2272) );
  XNOR U2272 ( .A(round_reg[1108]), .B(n2274), .Z(n1397) );
  XNOR U2273 ( .A(round_reg[1497]), .B(n2275), .Z(n1396) );
  XOR U2274 ( .A(n2276), .B(n1847), .Z(out[665]) );
  XOR U2275 ( .A(round_reg[263]), .B(n2277), .Z(n1847) );
  ANDN U2276 ( .B(n1400), .A(n1401), .Z(n2276) );
  XNOR U2277 ( .A(round_reg[1107]), .B(n2278), .Z(n1401) );
  XNOR U2278 ( .A(round_reg[1496]), .B(n2279), .Z(n1400) );
  XOR U2279 ( .A(n2280), .B(n1850), .Z(out[664]) );
  XOR U2280 ( .A(round_reg[262]), .B(n2281), .Z(n1850) );
  ANDN U2281 ( .B(n1404), .A(n1405), .Z(n2280) );
  XNOR U2282 ( .A(round_reg[1106]), .B(n2282), .Z(n1405) );
  XNOR U2283 ( .A(round_reg[1495]), .B(n2283), .Z(n1404) );
  XOR U2284 ( .A(n2284), .B(n1853), .Z(out[663]) );
  XOR U2285 ( .A(round_reg[261]), .B(n2285), .Z(n1853) );
  ANDN U2286 ( .B(n1412), .A(n1413), .Z(n2284) );
  XNOR U2287 ( .A(round_reg[1105]), .B(n2286), .Z(n1413) );
  XNOR U2288 ( .A(round_reg[1494]), .B(n2287), .Z(n1412) );
  XOR U2289 ( .A(n2288), .B(n1856), .Z(out[662]) );
  XOR U2290 ( .A(round_reg[260]), .B(n2289), .Z(n1856) );
  ANDN U2291 ( .B(n1416), .A(n1417), .Z(n2288) );
  XNOR U2292 ( .A(round_reg[1104]), .B(n2290), .Z(n1417) );
  XNOR U2293 ( .A(round_reg[1493]), .B(n2291), .Z(n1416) );
  XOR U2294 ( .A(n2292), .B(n1863), .Z(out[661]) );
  XOR U2295 ( .A(round_reg[259]), .B(n2293), .Z(n1863) );
  ANDN U2296 ( .B(n1420), .A(n1421), .Z(n2292) );
  XNOR U2297 ( .A(round_reg[1103]), .B(n2294), .Z(n1421) );
  XNOR U2298 ( .A(round_reg[1492]), .B(n2295), .Z(n1420) );
  XOR U2299 ( .A(n2296), .B(n1866), .Z(out[660]) );
  XOR U2300 ( .A(round_reg[258]), .B(n2297), .Z(n1866) );
  ANDN U2301 ( .B(n1424), .A(n1425), .Z(n2296) );
  XNOR U2302 ( .A(round_reg[1102]), .B(n2298), .Z(n1425) );
  XNOR U2303 ( .A(round_reg[1491]), .B(n2299), .Z(n1424) );
  XNOR U2304 ( .A(n2300), .B(n2301), .Z(out[65]) );
  AND U2305 ( .A(n2302), .B(n2303), .Z(n2300) );
  XOR U2306 ( .A(n2304), .B(n1869), .Z(out[659]) );
  XOR U2307 ( .A(round_reg[257]), .B(n2305), .Z(n1869) );
  ANDN U2308 ( .B(n1428), .A(n1429), .Z(n2304) );
  XNOR U2309 ( .A(round_reg[1101]), .B(n2306), .Z(n1429) );
  XNOR U2310 ( .A(round_reg[1490]), .B(n2307), .Z(n1428) );
  XOR U2311 ( .A(n2308), .B(n1872), .Z(out[658]) );
  XOR U2312 ( .A(round_reg[256]), .B(n2309), .Z(n1872) );
  ANDN U2313 ( .B(n1432), .A(n1433), .Z(n2308) );
  XNOR U2314 ( .A(round_reg[1100]), .B(n2310), .Z(n1433) );
  XNOR U2315 ( .A(round_reg[1489]), .B(n2311), .Z(n1432) );
  XOR U2316 ( .A(n2312), .B(n1875), .Z(out[657]) );
  XOR U2317 ( .A(round_reg[319]), .B(n2313), .Z(n1875) );
  ANDN U2318 ( .B(n1436), .A(n1437), .Z(n2312) );
  XNOR U2319 ( .A(round_reg[1099]), .B(n2314), .Z(n1437) );
  XNOR U2320 ( .A(round_reg[1488]), .B(n2315), .Z(n1436) );
  XOR U2321 ( .A(n2316), .B(n1878), .Z(out[656]) );
  XOR U2322 ( .A(round_reg[318]), .B(n2317), .Z(n1878) );
  ANDN U2323 ( .B(n1440), .A(n1441), .Z(n2316) );
  XNOR U2324 ( .A(round_reg[1098]), .B(n2318), .Z(n1441) );
  XNOR U2325 ( .A(round_reg[1487]), .B(n2319), .Z(n1440) );
  XOR U2326 ( .A(n2320), .B(n1881), .Z(out[655]) );
  XOR U2327 ( .A(round_reg[317]), .B(n2321), .Z(n1881) );
  ANDN U2328 ( .B(n1444), .A(n1445), .Z(n2320) );
  XNOR U2329 ( .A(round_reg[1097]), .B(n2322), .Z(n1445) );
  XNOR U2330 ( .A(round_reg[1486]), .B(n2323), .Z(n1444) );
  XOR U2331 ( .A(n2324), .B(n1884), .Z(out[654]) );
  XOR U2332 ( .A(round_reg[316]), .B(n2325), .Z(n1884) );
  ANDN U2333 ( .B(n1448), .A(n1449), .Z(n2324) );
  XNOR U2334 ( .A(round_reg[1096]), .B(n2326), .Z(n1449) );
  XNOR U2335 ( .A(round_reg[1485]), .B(n2327), .Z(n1448) );
  XOR U2336 ( .A(n2328), .B(n1887), .Z(out[653]) );
  XOR U2337 ( .A(round_reg[315]), .B(n2329), .Z(n1887) );
  ANDN U2338 ( .B(n1456), .A(n1457), .Z(n2328) );
  XNOR U2339 ( .A(round_reg[1095]), .B(n2330), .Z(n1457) );
  XNOR U2340 ( .A(round_reg[1484]), .B(n2331), .Z(n1456) );
  XOR U2341 ( .A(n2332), .B(n1890), .Z(out[652]) );
  XOR U2342 ( .A(round_reg[314]), .B(n2333), .Z(n1890) );
  ANDN U2343 ( .B(n1460), .A(n1461), .Z(n2332) );
  XNOR U2344 ( .A(round_reg[1094]), .B(n2334), .Z(n1461) );
  XNOR U2345 ( .A(round_reg[1483]), .B(n2335), .Z(n1460) );
  XOR U2346 ( .A(n2336), .B(n1897), .Z(out[651]) );
  XOR U2347 ( .A(round_reg[313]), .B(n2337), .Z(n1897) );
  ANDN U2348 ( .B(n1464), .A(n1465), .Z(n2336) );
  XNOR U2349 ( .A(round_reg[1093]), .B(n2338), .Z(n1465) );
  XNOR U2350 ( .A(round_reg[1482]), .B(n2339), .Z(n1464) );
  XOR U2351 ( .A(n2340), .B(n1900), .Z(out[650]) );
  XOR U2352 ( .A(round_reg[312]), .B(n2341), .Z(n1900) );
  ANDN U2353 ( .B(n1468), .A(n1469), .Z(n2340) );
  XNOR U2354 ( .A(round_reg[1092]), .B(n2342), .Z(n1469) );
  XNOR U2355 ( .A(round_reg[1481]), .B(n2343), .Z(n1468) );
  XNOR U2356 ( .A(n2344), .B(n2345), .Z(out[64]) );
  XOR U2357 ( .A(n2348), .B(n1903), .Z(out[649]) );
  XOR U2358 ( .A(round_reg[311]), .B(n2349), .Z(n1903) );
  ANDN U2359 ( .B(n1472), .A(n1473), .Z(n2348) );
  XNOR U2360 ( .A(round_reg[1091]), .B(n2350), .Z(n1473) );
  XNOR U2361 ( .A(round_reg[1480]), .B(n2351), .Z(n1472) );
  XOR U2362 ( .A(n2352), .B(n1906), .Z(out[648]) );
  XOR U2363 ( .A(round_reg[310]), .B(n2353), .Z(n1906) );
  ANDN U2364 ( .B(n1476), .A(n1477), .Z(n2352) );
  XNOR U2365 ( .A(round_reg[1090]), .B(n2354), .Z(n1477) );
  XNOR U2366 ( .A(round_reg[1479]), .B(n2355), .Z(n1476) );
  XOR U2367 ( .A(n2356), .B(n1909), .Z(out[647]) );
  XOR U2368 ( .A(round_reg[309]), .B(n2357), .Z(n1909) );
  ANDN U2369 ( .B(n1480), .A(n1481), .Z(n2356) );
  XNOR U2370 ( .A(round_reg[1089]), .B(n2358), .Z(n1481) );
  XNOR U2371 ( .A(round_reg[1478]), .B(n2359), .Z(n1480) );
  XOR U2372 ( .A(n2360), .B(n1912), .Z(out[646]) );
  XOR U2373 ( .A(round_reg[308]), .B(n2361), .Z(n1912) );
  ANDN U2374 ( .B(n1484), .A(n1485), .Z(n2360) );
  XNOR U2375 ( .A(round_reg[1088]), .B(n2362), .Z(n1485) );
  XNOR U2376 ( .A(round_reg[1477]), .B(n2363), .Z(n1484) );
  XOR U2377 ( .A(n2364), .B(n1915), .Z(out[645]) );
  XOR U2378 ( .A(round_reg[307]), .B(n2365), .Z(n1915) );
  ANDN U2379 ( .B(n1488), .A(n1489), .Z(n2364) );
  XNOR U2380 ( .A(round_reg[1151]), .B(n2366), .Z(n1489) );
  XNOR U2381 ( .A(round_reg[1476]), .B(n2367), .Z(n1488) );
  XOR U2382 ( .A(n2368), .B(n1918), .Z(out[644]) );
  XOR U2383 ( .A(round_reg[306]), .B(n2369), .Z(n1918) );
  ANDN U2384 ( .B(n1492), .A(n1493), .Z(n2368) );
  XNOR U2385 ( .A(round_reg[1150]), .B(n2370), .Z(n1493) );
  XNOR U2386 ( .A(round_reg[1475]), .B(n2371), .Z(n1492) );
  XOR U2387 ( .A(n2372), .B(n1921), .Z(out[643]) );
  XOR U2388 ( .A(round_reg[305]), .B(n2373), .Z(n1921) );
  ANDN U2389 ( .B(n1504), .A(n1505), .Z(n2372) );
  XNOR U2390 ( .A(round_reg[1149]), .B(n2374), .Z(n1505) );
  XNOR U2391 ( .A(round_reg[1474]), .B(n2375), .Z(n1504) );
  XOR U2392 ( .A(n2376), .B(n1924), .Z(out[642]) );
  XOR U2393 ( .A(round_reg[304]), .B(n2377), .Z(n1924) );
  ANDN U2394 ( .B(n1508), .A(n1509), .Z(n2376) );
  XNOR U2395 ( .A(round_reg[1148]), .B(n2378), .Z(n1509) );
  XNOR U2396 ( .A(round_reg[1473]), .B(n2379), .Z(n1508) );
  XOR U2397 ( .A(n2380), .B(n1931), .Z(out[641]) );
  XOR U2398 ( .A(round_reg[303]), .B(n2381), .Z(n1931) );
  ANDN U2399 ( .B(n1512), .A(n1513), .Z(n2380) );
  XNOR U2400 ( .A(round_reg[1147]), .B(n2382), .Z(n1513) );
  XNOR U2401 ( .A(round_reg[1472]), .B(n2383), .Z(n1512) );
  XOR U2402 ( .A(n2384), .B(n1934), .Z(out[640]) );
  XOR U2403 ( .A(round_reg[302]), .B(n2385), .Z(n1934) );
  ANDN U2404 ( .B(n1516), .A(n1517), .Z(n2384) );
  XNOR U2405 ( .A(round_reg[1146]), .B(n2386), .Z(n1517) );
  XNOR U2406 ( .A(round_reg[1535]), .B(n2387), .Z(n1516) );
  XNOR U2407 ( .A(n2388), .B(n2389), .Z(out[63]) );
  AND U2408 ( .A(n2390), .B(n2391), .Z(n2388) );
  XNOR U2409 ( .A(n2392), .B(n2393), .Z(out[639]) );
  AND U2410 ( .A(n2394), .B(n2395), .Z(n2392) );
  XNOR U2411 ( .A(n2396), .B(n2397), .Z(out[638]) );
  AND U2412 ( .A(n2398), .B(n2399), .Z(n2396) );
  XNOR U2413 ( .A(n2400), .B(n2401), .Z(out[637]) );
  AND U2414 ( .A(n2402), .B(n2403), .Z(n2400) );
  XNOR U2415 ( .A(n2404), .B(n2405), .Z(out[636]) );
  AND U2416 ( .A(n2406), .B(n2407), .Z(n2404) );
  XNOR U2417 ( .A(n2408), .B(n2409), .Z(out[635]) );
  AND U2418 ( .A(n2410), .B(n2411), .Z(n2408) );
  XNOR U2419 ( .A(n2412), .B(n2413), .Z(out[634]) );
  AND U2420 ( .A(n2414), .B(n2415), .Z(n2412) );
  XNOR U2421 ( .A(n2416), .B(n2417), .Z(out[633]) );
  AND U2422 ( .A(n2418), .B(n2419), .Z(n2416) );
  XNOR U2423 ( .A(n2420), .B(n2421), .Z(out[632]) );
  AND U2424 ( .A(n2422), .B(n2423), .Z(n2420) );
  XNOR U2425 ( .A(n2424), .B(n2425), .Z(out[631]) );
  AND U2426 ( .A(n2426), .B(n2427), .Z(n2424) );
  XNOR U2427 ( .A(n2428), .B(n2429), .Z(out[630]) );
  AND U2428 ( .A(n2430), .B(n2431), .Z(n2428) );
  XNOR U2429 ( .A(n2432), .B(n2433), .Z(out[62]) );
  AND U2430 ( .A(n2434), .B(n2435), .Z(n2432) );
  XNOR U2431 ( .A(n2436), .B(n2437), .Z(out[629]) );
  AND U2432 ( .A(n2438), .B(n2439), .Z(n2436) );
  XNOR U2433 ( .A(n2440), .B(n2441), .Z(out[628]) );
  AND U2434 ( .A(n2442), .B(n2443), .Z(n2440) );
  XNOR U2435 ( .A(n2444), .B(n2445), .Z(out[627]) );
  AND U2436 ( .A(n2446), .B(n2447), .Z(n2444) );
  XNOR U2437 ( .A(n2448), .B(n2449), .Z(out[626]) );
  AND U2438 ( .A(n2450), .B(n2451), .Z(n2448) );
  XNOR U2439 ( .A(n2452), .B(n2453), .Z(out[625]) );
  AND U2440 ( .A(n2454), .B(n2455), .Z(n2452) );
  XNOR U2441 ( .A(n2456), .B(n2457), .Z(out[624]) );
  AND U2442 ( .A(n2458), .B(n2459), .Z(n2456) );
  XNOR U2443 ( .A(n2460), .B(n2461), .Z(out[623]) );
  AND U2444 ( .A(n2462), .B(n2463), .Z(n2460) );
  XNOR U2445 ( .A(n2464), .B(n2465), .Z(out[622]) );
  AND U2446 ( .A(n2466), .B(n2467), .Z(n2464) );
  XNOR U2447 ( .A(n2468), .B(n2469), .Z(out[621]) );
  AND U2448 ( .A(n2470), .B(n2471), .Z(n2468) );
  XNOR U2449 ( .A(n2472), .B(n2473), .Z(out[620]) );
  AND U2450 ( .A(n2474), .B(n2475), .Z(n2472) );
  XNOR U2451 ( .A(n2476), .B(n2477), .Z(out[61]) );
  AND U2452 ( .A(n2478), .B(n2479), .Z(n2476) );
  XNOR U2453 ( .A(n2480), .B(n2481), .Z(out[619]) );
  AND U2454 ( .A(n2482), .B(n2483), .Z(n2480) );
  XNOR U2455 ( .A(n2484), .B(n2485), .Z(out[618]) );
  AND U2456 ( .A(n2486), .B(n2487), .Z(n2484) );
  XNOR U2457 ( .A(n2488), .B(n2489), .Z(out[617]) );
  AND U2458 ( .A(n2490), .B(n2491), .Z(n2488) );
  XNOR U2459 ( .A(n2492), .B(n2493), .Z(out[616]) );
  AND U2460 ( .A(n2494), .B(n2495), .Z(n2492) );
  XNOR U2461 ( .A(n2496), .B(n2497), .Z(out[615]) );
  AND U2462 ( .A(n2498), .B(n2499), .Z(n2496) );
  XNOR U2463 ( .A(n2500), .B(n2501), .Z(out[614]) );
  AND U2464 ( .A(n2502), .B(n2503), .Z(n2500) );
  XNOR U2465 ( .A(n2504), .B(n2505), .Z(out[613]) );
  AND U2466 ( .A(n2506), .B(n2507), .Z(n2504) );
  XNOR U2467 ( .A(n2508), .B(n2509), .Z(out[612]) );
  AND U2468 ( .A(n2510), .B(n2511), .Z(n2508) );
  XNOR U2469 ( .A(n2512), .B(n2513), .Z(out[611]) );
  AND U2470 ( .A(n2514), .B(n2515), .Z(n2512) );
  XNOR U2471 ( .A(n2516), .B(n2517), .Z(out[610]) );
  AND U2472 ( .A(n2518), .B(n2519), .Z(n2516) );
  XNOR U2473 ( .A(n2520), .B(n2521), .Z(out[60]) );
  AND U2474 ( .A(n2522), .B(n2523), .Z(n2520) );
  XNOR U2475 ( .A(n2524), .B(n2525), .Z(out[609]) );
  AND U2476 ( .A(n2526), .B(n2527), .Z(n2524) );
  XNOR U2477 ( .A(n2528), .B(n2529), .Z(out[608]) );
  AND U2478 ( .A(n2530), .B(n2531), .Z(n2528) );
  XNOR U2479 ( .A(n2532), .B(n2533), .Z(out[607]) );
  AND U2480 ( .A(n2534), .B(n2535), .Z(n2532) );
  XNOR U2481 ( .A(n2536), .B(n2537), .Z(out[606]) );
  AND U2482 ( .A(n2538), .B(n2539), .Z(n2536) );
  XNOR U2483 ( .A(n2540), .B(n2541), .Z(out[605]) );
  AND U2484 ( .A(n2542), .B(n2543), .Z(n2540) );
  XNOR U2485 ( .A(n2544), .B(n2545), .Z(out[604]) );
  AND U2486 ( .A(n2546), .B(n2547), .Z(n2544) );
  XNOR U2487 ( .A(n2548), .B(n2549), .Z(out[603]) );
  AND U2488 ( .A(n2550), .B(n2551), .Z(n2548) );
  XNOR U2489 ( .A(n2552), .B(n2553), .Z(out[602]) );
  AND U2490 ( .A(n2554), .B(n2555), .Z(n2552) );
  XNOR U2491 ( .A(n2556), .B(n2557), .Z(out[601]) );
  AND U2492 ( .A(n2558), .B(n2559), .Z(n2556) );
  XNOR U2493 ( .A(n2560), .B(n2561), .Z(out[600]) );
  AND U2494 ( .A(n2562), .B(n2563), .Z(n2560) );
  XNOR U2495 ( .A(n2564), .B(n2126), .Z(out[5]) );
  AND U2496 ( .A(n2565), .B(n2566), .Z(n2564) );
  XNOR U2497 ( .A(n2567), .B(n2568), .Z(out[59]) );
  AND U2498 ( .A(n2569), .B(n2570), .Z(n2567) );
  XNOR U2499 ( .A(n2571), .B(n2572), .Z(out[599]) );
  AND U2500 ( .A(n2573), .B(n2574), .Z(n2571) );
  XNOR U2501 ( .A(n2575), .B(n2576), .Z(out[598]) );
  AND U2502 ( .A(n2577), .B(n2578), .Z(n2575) );
  XNOR U2503 ( .A(n2579), .B(n2580), .Z(out[597]) );
  AND U2504 ( .A(n2581), .B(n2582), .Z(n2579) );
  XNOR U2505 ( .A(n2583), .B(n2584), .Z(out[596]) );
  AND U2506 ( .A(n2585), .B(n2586), .Z(n2583) );
  XNOR U2507 ( .A(n2587), .B(n2588), .Z(out[595]) );
  AND U2508 ( .A(n2589), .B(n2590), .Z(n2587) );
  XNOR U2509 ( .A(n2591), .B(n2592), .Z(out[594]) );
  AND U2510 ( .A(n2593), .B(n2594), .Z(n2591) );
  XNOR U2511 ( .A(n2595), .B(n2596), .Z(out[593]) );
  AND U2512 ( .A(n2597), .B(n2598), .Z(n2595) );
  XNOR U2513 ( .A(n2599), .B(n2600), .Z(out[592]) );
  AND U2514 ( .A(n2601), .B(n2602), .Z(n2599) );
  XNOR U2515 ( .A(n2603), .B(n2604), .Z(out[591]) );
  AND U2516 ( .A(n2605), .B(n2606), .Z(n2603) );
  XNOR U2517 ( .A(n2607), .B(n2608), .Z(out[590]) );
  AND U2518 ( .A(n2609), .B(n2610), .Z(n2607) );
  XNOR U2519 ( .A(n2611), .B(n2612), .Z(out[58]) );
  AND U2520 ( .A(n2613), .B(n2614), .Z(n2611) );
  XNOR U2521 ( .A(n2615), .B(n2616), .Z(out[589]) );
  AND U2522 ( .A(n2617), .B(n2618), .Z(n2615) );
  XNOR U2523 ( .A(n2619), .B(n2620), .Z(out[588]) );
  AND U2524 ( .A(n2621), .B(n2622), .Z(n2619) );
  XNOR U2525 ( .A(n2623), .B(n2624), .Z(out[587]) );
  AND U2526 ( .A(n2625), .B(n2626), .Z(n2623) );
  XNOR U2527 ( .A(n2627), .B(n2628), .Z(out[586]) );
  AND U2528 ( .A(n2629), .B(n2630), .Z(n2627) );
  XNOR U2529 ( .A(n2631), .B(n2632), .Z(out[585]) );
  AND U2530 ( .A(n2633), .B(n2634), .Z(n2631) );
  XNOR U2531 ( .A(n2635), .B(n2636), .Z(out[584]) );
  AND U2532 ( .A(n2637), .B(n2638), .Z(n2635) );
  XNOR U2533 ( .A(n2639), .B(n2640), .Z(out[583]) );
  AND U2534 ( .A(n2641), .B(n2642), .Z(n2639) );
  XNOR U2535 ( .A(n2643), .B(n2644), .Z(out[582]) );
  AND U2536 ( .A(n2645), .B(n2646), .Z(n2643) );
  XNOR U2537 ( .A(n2647), .B(n2648), .Z(out[581]) );
  AND U2538 ( .A(n2649), .B(n2650), .Z(n2647) );
  XNOR U2539 ( .A(n2651), .B(n2652), .Z(out[580]) );
  AND U2540 ( .A(n2653), .B(n2654), .Z(n2651) );
  XNOR U2541 ( .A(n2655), .B(n2656), .Z(out[57]) );
  AND U2542 ( .A(n2657), .B(n2658), .Z(n2655) );
  XNOR U2543 ( .A(n2659), .B(n2660), .Z(out[579]) );
  AND U2544 ( .A(n2661), .B(n2662), .Z(n2659) );
  XNOR U2545 ( .A(n2663), .B(n2664), .Z(out[578]) );
  AND U2546 ( .A(n2665), .B(n2666), .Z(n2663) );
  XNOR U2547 ( .A(n2667), .B(n2668), .Z(out[577]) );
  AND U2548 ( .A(n2669), .B(n2670), .Z(n2667) );
  XNOR U2549 ( .A(n2671), .B(n2672), .Z(out[576]) );
  AND U2550 ( .A(n2673), .B(n2674), .Z(n2671) );
  XNOR U2551 ( .A(n2675), .B(n2394), .Z(out[575]) );
  XNOR U2552 ( .A(n2677), .B(n2398), .Z(out[574]) );
  XNOR U2553 ( .A(n2679), .B(n2402), .Z(out[573]) );
  XNOR U2554 ( .A(n2681), .B(n2406), .Z(out[572]) );
  XNOR U2555 ( .A(n2683), .B(n2410), .Z(out[571]) );
  XNOR U2556 ( .A(n2685), .B(n2414), .Z(out[570]) );
  XNOR U2557 ( .A(n2687), .B(n2688), .Z(out[56]) );
  AND U2558 ( .A(n2689), .B(n2690), .Z(n2687) );
  XNOR U2559 ( .A(n2691), .B(n2418), .Z(out[569]) );
  XNOR U2560 ( .A(n2693), .B(n2422), .Z(out[568]) );
  XNOR U2561 ( .A(n2695), .B(n2426), .Z(out[567]) );
  AND U2562 ( .A(n2696), .B(n2697), .Z(n2695) );
  XNOR U2563 ( .A(n2698), .B(n2430), .Z(out[566]) );
  AND U2564 ( .A(n2699), .B(n2700), .Z(n2698) );
  XNOR U2565 ( .A(n2701), .B(n2438), .Z(out[565]) );
  AND U2566 ( .A(n2702), .B(n2703), .Z(n2701) );
  XNOR U2567 ( .A(n2704), .B(n2442), .Z(out[564]) );
  AND U2568 ( .A(n2705), .B(n2706), .Z(n2704) );
  XNOR U2569 ( .A(n2707), .B(n2446), .Z(out[563]) );
  AND U2570 ( .A(n2708), .B(n2709), .Z(n2707) );
  XNOR U2571 ( .A(n2710), .B(n2450), .Z(out[562]) );
  AND U2572 ( .A(n2711), .B(n2712), .Z(n2710) );
  XNOR U2573 ( .A(n2713), .B(n2454), .Z(out[561]) );
  AND U2574 ( .A(n2714), .B(n2715), .Z(n2713) );
  XNOR U2575 ( .A(n2716), .B(n2458), .Z(out[560]) );
  AND U2576 ( .A(n2717), .B(n2718), .Z(n2716) );
  XNOR U2577 ( .A(n2719), .B(n2720), .Z(out[55]) );
  AND U2578 ( .A(n2721), .B(n2722), .Z(n2719) );
  XNOR U2579 ( .A(n2723), .B(n2462), .Z(out[559]) );
  AND U2580 ( .A(n2724), .B(n2725), .Z(n2723) );
  XNOR U2581 ( .A(n2726), .B(n2466), .Z(out[558]) );
  AND U2582 ( .A(n2727), .B(n2728), .Z(n2726) );
  XNOR U2583 ( .A(n2729), .B(n2470), .Z(out[557]) );
  AND U2584 ( .A(n2730), .B(n2731), .Z(n2729) );
  XNOR U2585 ( .A(n2732), .B(n2474), .Z(out[556]) );
  AND U2586 ( .A(n2733), .B(n2734), .Z(n2732) );
  XNOR U2587 ( .A(n2735), .B(n2482), .Z(out[555]) );
  AND U2588 ( .A(n2736), .B(n2737), .Z(n2735) );
  XNOR U2589 ( .A(n2738), .B(n2486), .Z(out[554]) );
  XNOR U2590 ( .A(n2740), .B(n2490), .Z(out[553]) );
  XNOR U2591 ( .A(n2742), .B(n2494), .Z(out[552]) );
  XNOR U2592 ( .A(n2744), .B(n2498), .Z(out[551]) );
  XNOR U2593 ( .A(n2746), .B(n2502), .Z(out[550]) );
  XNOR U2594 ( .A(n2748), .B(n2749), .Z(out[54]) );
  AND U2595 ( .A(n2750), .B(n2751), .Z(n2748) );
  XNOR U2596 ( .A(n2752), .B(n2506), .Z(out[549]) );
  AND U2597 ( .A(n2753), .B(n2754), .Z(n2752) );
  XNOR U2598 ( .A(n2755), .B(n2510), .Z(out[548]) );
  AND U2599 ( .A(n2756), .B(n2757), .Z(n2755) );
  XNOR U2600 ( .A(n2758), .B(n2514), .Z(out[547]) );
  AND U2601 ( .A(n2759), .B(n2760), .Z(n2758) );
  XNOR U2602 ( .A(n2761), .B(n2518), .Z(out[546]) );
  AND U2603 ( .A(n2762), .B(n2763), .Z(n2761) );
  XNOR U2604 ( .A(n2764), .B(n2526), .Z(out[545]) );
  AND U2605 ( .A(n2765), .B(n2766), .Z(n2764) );
  XNOR U2606 ( .A(n2767), .B(n2530), .Z(out[544]) );
  AND U2607 ( .A(n2768), .B(n2769), .Z(n2767) );
  XNOR U2608 ( .A(n2770), .B(n2534), .Z(out[543]) );
  AND U2609 ( .A(n2771), .B(n2772), .Z(n2770) );
  XNOR U2610 ( .A(n2773), .B(n2538), .Z(out[542]) );
  AND U2611 ( .A(n2774), .B(n2775), .Z(n2773) );
  XNOR U2612 ( .A(n2776), .B(n2542), .Z(out[541]) );
  AND U2613 ( .A(n2777), .B(n2778), .Z(n2776) );
  XNOR U2614 ( .A(n2779), .B(n2546), .Z(out[540]) );
  XNOR U2615 ( .A(n2781), .B(n2782), .Z(out[53]) );
  AND U2616 ( .A(n2783), .B(n2784), .Z(n2781) );
  XNOR U2617 ( .A(n2785), .B(n2550), .Z(out[539]) );
  XNOR U2618 ( .A(n2787), .B(n2554), .Z(out[538]) );
  XNOR U2619 ( .A(n2789), .B(n2558), .Z(out[537]) );
  XNOR U2620 ( .A(n2791), .B(n2562), .Z(out[536]) );
  XNOR U2621 ( .A(n2793), .B(n2573), .Z(out[535]) );
  XNOR U2622 ( .A(n2795), .B(n2577), .Z(out[534]) );
  XNOR U2623 ( .A(n2797), .B(n2581), .Z(out[533]) );
  XNOR U2624 ( .A(n2799), .B(n2585), .Z(out[532]) );
  XNOR U2625 ( .A(n2801), .B(n2589), .Z(out[531]) );
  XNOR U2626 ( .A(n2803), .B(n2593), .Z(out[530]) );
  XNOR U2627 ( .A(n2805), .B(n2806), .Z(out[52]) );
  AND U2628 ( .A(n2807), .B(n2808), .Z(n2805) );
  XNOR U2629 ( .A(n2809), .B(n2597), .Z(out[529]) );
  AND U2630 ( .A(n2810), .B(n2811), .Z(n2809) );
  XNOR U2631 ( .A(n2812), .B(n2601), .Z(out[528]) );
  XNOR U2632 ( .A(n2814), .B(n2605), .Z(out[527]) );
  XNOR U2633 ( .A(n2816), .B(n2609), .Z(out[526]) );
  XNOR U2634 ( .A(n2818), .B(n2617), .Z(out[525]) );
  XNOR U2635 ( .A(n2820), .B(n2621), .Z(out[524]) );
  XNOR U2636 ( .A(n2822), .B(n2625), .Z(out[523]) );
  XNOR U2637 ( .A(n2824), .B(n2629), .Z(out[522]) );
  XNOR U2638 ( .A(n2826), .B(n2633), .Z(out[521]) );
  XNOR U2639 ( .A(n2828), .B(n2637), .Z(out[520]) );
  XNOR U2640 ( .A(n2830), .B(n2831), .Z(out[51]) );
  AND U2641 ( .A(n2832), .B(n2833), .Z(n2830) );
  XNOR U2642 ( .A(n2834), .B(n2641), .Z(out[519]) );
  XNOR U2643 ( .A(n2836), .B(n2645), .Z(out[518]) );
  AND U2644 ( .A(n2837), .B(n2838), .Z(n2836) );
  XNOR U2645 ( .A(n2839), .B(n2649), .Z(out[517]) );
  AND U2646 ( .A(n2840), .B(n2841), .Z(n2839) );
  XNOR U2647 ( .A(n2842), .B(n2653), .Z(out[516]) );
  XNOR U2648 ( .A(n2844), .B(n2661), .Z(out[515]) );
  XNOR U2649 ( .A(n2846), .B(n2665), .Z(out[514]) );
  XNOR U2650 ( .A(n2848), .B(n2669), .Z(out[513]) );
  XNOR U2651 ( .A(n2850), .B(n2673), .Z(out[512]) );
  XOR U2652 ( .A(n2852), .B(n2395), .Z(out[511]) );
  XOR U2653 ( .A(round_reg[885]), .B(n2151), .Z(n2395) );
  ANDN U2654 ( .B(n2853), .A(n2676), .Z(n2852) );
  XOR U2655 ( .A(n2854), .B(n2399), .Z(out[510]) );
  XOR U2656 ( .A(round_reg[884]), .B(n2155), .Z(n2399) );
  ANDN U2657 ( .B(n2855), .A(n2678), .Z(n2854) );
  XNOR U2658 ( .A(n2856), .B(n2857), .Z(out[50]) );
  AND U2659 ( .A(n2858), .B(n2859), .Z(n2856) );
  XOR U2660 ( .A(n2860), .B(n2403), .Z(out[509]) );
  XOR U2661 ( .A(round_reg[883]), .B(n2159), .Z(n2403) );
  ANDN U2662 ( .B(n2861), .A(n2680), .Z(n2860) );
  XOR U2663 ( .A(n2862), .B(n2407), .Z(out[508]) );
  XOR U2664 ( .A(round_reg[882]), .B(n2163), .Z(n2407) );
  ANDN U2665 ( .B(n2863), .A(n2682), .Z(n2862) );
  XOR U2666 ( .A(n2864), .B(n2411), .Z(out[507]) );
  XOR U2667 ( .A(round_reg[881]), .B(n2167), .Z(n2411) );
  ANDN U2668 ( .B(n2865), .A(n2684), .Z(n2864) );
  XOR U2669 ( .A(n2866), .B(n2415), .Z(out[506]) );
  XOR U2670 ( .A(round_reg[880]), .B(n2175), .Z(n2415) );
  ANDN U2671 ( .B(n2867), .A(n2686), .Z(n2866) );
  XOR U2672 ( .A(n2868), .B(n2419), .Z(out[505]) );
  XOR U2673 ( .A(round_reg[879]), .B(n2179), .Z(n2419) );
  ANDN U2674 ( .B(n2869), .A(n2692), .Z(n2868) );
  XOR U2675 ( .A(n2870), .B(n2423), .Z(out[504]) );
  XOR U2676 ( .A(round_reg[878]), .B(n2183), .Z(n2423) );
  ANDN U2677 ( .B(n2871), .A(n2694), .Z(n2870) );
  XOR U2678 ( .A(n2872), .B(n2427), .Z(out[503]) );
  IV U2679 ( .A(n2697), .Z(n2427) );
  XNOR U2680 ( .A(round_reg[877]), .B(n2187), .Z(n2697) );
  ANDN U2681 ( .B(n2873), .A(n2696), .Z(n2872) );
  XOR U2682 ( .A(n2874), .B(n2431), .Z(out[502]) );
  IV U2683 ( .A(n2700), .Z(n2431) );
  XNOR U2684 ( .A(round_reg[876]), .B(n2191), .Z(n2700) );
  ANDN U2685 ( .B(n2875), .A(n2699), .Z(n2874) );
  XOR U2686 ( .A(n2876), .B(n2439), .Z(out[501]) );
  IV U2687 ( .A(n2703), .Z(n2439) );
  XNOR U2688 ( .A(round_reg[875]), .B(n2195), .Z(n2703) );
  ANDN U2689 ( .B(n2877), .A(n2702), .Z(n2876) );
  XOR U2690 ( .A(n2878), .B(n2443), .Z(out[500]) );
  IV U2691 ( .A(n2706), .Z(n2443) );
  XNOR U2692 ( .A(round_reg[874]), .B(n2199), .Z(n2706) );
  ANDN U2693 ( .B(n2879), .A(n2705), .Z(n2878) );
  XNOR U2694 ( .A(n2880), .B(n2170), .Z(out[4]) );
  AND U2695 ( .A(n2881), .B(n2882), .Z(n2880) );
  XNOR U2696 ( .A(n2883), .B(n2884), .Z(out[49]) );
  AND U2697 ( .A(n2885), .B(n2886), .Z(n2883) );
  XOR U2698 ( .A(n2887), .B(n2447), .Z(out[499]) );
  IV U2699 ( .A(n2709), .Z(n2447) );
  XNOR U2700 ( .A(round_reg[873]), .B(n2203), .Z(n2709) );
  ANDN U2701 ( .B(n2888), .A(n2708), .Z(n2887) );
  XOR U2702 ( .A(n2889), .B(n2451), .Z(out[498]) );
  IV U2703 ( .A(n2712), .Z(n2451) );
  XNOR U2704 ( .A(round_reg[872]), .B(n2207), .Z(n2712) );
  ANDN U2705 ( .B(n2890), .A(n2711), .Z(n2889) );
  XOR U2706 ( .A(n2891), .B(n2455), .Z(out[497]) );
  IV U2707 ( .A(n2715), .Z(n2455) );
  XNOR U2708 ( .A(round_reg[871]), .B(n2211), .Z(n2715) );
  ANDN U2709 ( .B(n2892), .A(n2714), .Z(n2891) );
  XOR U2710 ( .A(n2893), .B(n2459), .Z(out[496]) );
  IV U2711 ( .A(n2718), .Z(n2459) );
  XNOR U2712 ( .A(round_reg[870]), .B(n2219), .Z(n2718) );
  ANDN U2713 ( .B(n2894), .A(n2717), .Z(n2893) );
  XOR U2714 ( .A(n2895), .B(n2463), .Z(out[495]) );
  IV U2715 ( .A(n2725), .Z(n2463) );
  XNOR U2716 ( .A(round_reg[869]), .B(n2223), .Z(n2725) );
  ANDN U2717 ( .B(n2896), .A(n2724), .Z(n2895) );
  XOR U2718 ( .A(n2897), .B(n2467), .Z(out[494]) );
  IV U2719 ( .A(n2728), .Z(n2467) );
  XNOR U2720 ( .A(round_reg[868]), .B(n2227), .Z(n2728) );
  ANDN U2721 ( .B(n2898), .A(n2727), .Z(n2897) );
  XOR U2722 ( .A(n2899), .B(n2471), .Z(out[493]) );
  IV U2723 ( .A(n2731), .Z(n2471) );
  XNOR U2724 ( .A(round_reg[867]), .B(n2231), .Z(n2731) );
  ANDN U2725 ( .B(n2900), .A(n2730), .Z(n2899) );
  XOR U2726 ( .A(n2901), .B(n2475), .Z(out[492]) );
  IV U2727 ( .A(n2734), .Z(n2475) );
  XNOR U2728 ( .A(round_reg[866]), .B(n2235), .Z(n2734) );
  ANDN U2729 ( .B(n2902), .A(n2733), .Z(n2901) );
  XOR U2730 ( .A(n2903), .B(n2483), .Z(out[491]) );
  IV U2731 ( .A(n2737), .Z(n2483) );
  XNOR U2732 ( .A(round_reg[865]), .B(n2239), .Z(n2737) );
  ANDN U2733 ( .B(n2904), .A(n2736), .Z(n2903) );
  XOR U2734 ( .A(n2905), .B(n2487), .Z(out[490]) );
  XNOR U2735 ( .A(round_reg[864]), .B(n2243), .Z(n2487) );
  ANDN U2736 ( .B(n2906), .A(n2739), .Z(n2905) );
  XNOR U2737 ( .A(n2907), .B(n2908), .Z(out[48]) );
  AND U2738 ( .A(n2909), .B(n2910), .Z(n2907) );
  XOR U2739 ( .A(n2911), .B(n2491), .Z(out[489]) );
  XNOR U2740 ( .A(round_reg[863]), .B(n2247), .Z(n2491) );
  ANDN U2741 ( .B(n2912), .A(n2741), .Z(n2911) );
  XOR U2742 ( .A(n2913), .B(n2495), .Z(out[488]) );
  XNOR U2743 ( .A(round_reg[862]), .B(n2251), .Z(n2495) );
  ANDN U2744 ( .B(n2914), .A(n2743), .Z(n2913) );
  XOR U2745 ( .A(n2915), .B(n2499), .Z(out[487]) );
  XNOR U2746 ( .A(round_reg[861]), .B(n2255), .Z(n2499) );
  ANDN U2747 ( .B(n2916), .A(n2745), .Z(n2915) );
  XOR U2748 ( .A(n2917), .B(n2503), .Z(out[486]) );
  XNOR U2749 ( .A(round_reg[860]), .B(n2263), .Z(n2503) );
  ANDN U2750 ( .B(n2918), .A(n2747), .Z(n2917) );
  XOR U2751 ( .A(n2919), .B(n2507), .Z(out[485]) );
  IV U2752 ( .A(n2754), .Z(n2507) );
  XNOR U2753 ( .A(round_reg[859]), .B(n2267), .Z(n2754) );
  ANDN U2754 ( .B(n2920), .A(n2753), .Z(n2919) );
  XOR U2755 ( .A(n2921), .B(n2511), .Z(out[484]) );
  IV U2756 ( .A(n2757), .Z(n2511) );
  XNOR U2757 ( .A(round_reg[858]), .B(n2271), .Z(n2757) );
  ANDN U2758 ( .B(n2922), .A(n2756), .Z(n2921) );
  XOR U2759 ( .A(n2923), .B(n2515), .Z(out[483]) );
  IV U2760 ( .A(n2760), .Z(n2515) );
  XNOR U2761 ( .A(round_reg[857]), .B(n2275), .Z(n2760) );
  ANDN U2762 ( .B(n2924), .A(n2759), .Z(n2923) );
  XOR U2763 ( .A(n2925), .B(n2519), .Z(out[482]) );
  IV U2764 ( .A(n2763), .Z(n2519) );
  XNOR U2765 ( .A(round_reg[856]), .B(n2279), .Z(n2763) );
  ANDN U2766 ( .B(n2926), .A(n2762), .Z(n2925) );
  XOR U2767 ( .A(n2927), .B(n2527), .Z(out[481]) );
  IV U2768 ( .A(n2766), .Z(n2527) );
  XNOR U2769 ( .A(round_reg[855]), .B(n2283), .Z(n2766) );
  ANDN U2770 ( .B(n2928), .A(n2765), .Z(n2927) );
  XOR U2771 ( .A(n2929), .B(n2531), .Z(out[480]) );
  IV U2772 ( .A(n2769), .Z(n2531) );
  XNOR U2773 ( .A(round_reg[854]), .B(n2287), .Z(n2769) );
  ANDN U2774 ( .B(n2930), .A(n2768), .Z(n2929) );
  XNOR U2775 ( .A(n2931), .B(n2932), .Z(out[47]) );
  AND U2776 ( .A(n2933), .B(n2934), .Z(n2931) );
  XOR U2777 ( .A(n2935), .B(n2535), .Z(out[479]) );
  IV U2778 ( .A(n2772), .Z(n2535) );
  XNOR U2779 ( .A(round_reg[853]), .B(n2291), .Z(n2772) );
  ANDN U2780 ( .B(n2936), .A(n2771), .Z(n2935) );
  XOR U2781 ( .A(n2937), .B(n2539), .Z(out[478]) );
  IV U2782 ( .A(n2775), .Z(n2539) );
  XNOR U2783 ( .A(round_reg[852]), .B(n2295), .Z(n2775) );
  ANDN U2784 ( .B(n2938), .A(n2774), .Z(n2937) );
  XOR U2785 ( .A(n2939), .B(n2543), .Z(out[477]) );
  IV U2786 ( .A(n2778), .Z(n2543) );
  XNOR U2787 ( .A(round_reg[851]), .B(n2299), .Z(n2778) );
  NOR U2788 ( .A(n2940), .B(n2777), .Z(n2939) );
  XOR U2789 ( .A(n2941), .B(n2547), .Z(out[476]) );
  XOR U2790 ( .A(round_reg[850]), .B(n2307), .Z(n2547) );
  NOR U2791 ( .A(n2942), .B(n2780), .Z(n2941) );
  XOR U2792 ( .A(n2943), .B(n2551), .Z(out[475]) );
  XOR U2793 ( .A(round_reg[849]), .B(n2311), .Z(n2551) );
  NOR U2794 ( .A(n2944), .B(n2786), .Z(n2943) );
  XOR U2795 ( .A(n2945), .B(n2555), .Z(out[474]) );
  XOR U2796 ( .A(round_reg[848]), .B(n2315), .Z(n2555) );
  ANDN U2797 ( .B(n2946), .A(n2788), .Z(n2945) );
  XOR U2798 ( .A(n2947), .B(n2559), .Z(out[473]) );
  XOR U2799 ( .A(round_reg[847]), .B(n2319), .Z(n2559) );
  ANDN U2800 ( .B(n2948), .A(n2790), .Z(n2947) );
  XOR U2801 ( .A(n2949), .B(n2563), .Z(out[472]) );
  XOR U2802 ( .A(round_reg[846]), .B(n2323), .Z(n2563) );
  ANDN U2803 ( .B(n2950), .A(n2792), .Z(n2949) );
  XOR U2804 ( .A(n2951), .B(n2574), .Z(out[471]) );
  XOR U2805 ( .A(round_reg[845]), .B(n2327), .Z(n2574) );
  ANDN U2806 ( .B(n2952), .A(n2794), .Z(n2951) );
  XOR U2807 ( .A(n2953), .B(n2578), .Z(out[470]) );
  XOR U2808 ( .A(round_reg[844]), .B(n2331), .Z(n2578) );
  ANDN U2809 ( .B(n2954), .A(n2796), .Z(n2953) );
  XNOR U2810 ( .A(n2955), .B(n2956), .Z(out[46]) );
  AND U2811 ( .A(n2957), .B(n2958), .Z(n2955) );
  XOR U2812 ( .A(n2959), .B(n2582), .Z(out[469]) );
  XOR U2813 ( .A(round_reg[843]), .B(n2335), .Z(n2582) );
  ANDN U2814 ( .B(n2960), .A(n2798), .Z(n2959) );
  XOR U2815 ( .A(n2961), .B(n2586), .Z(out[468]) );
  XOR U2816 ( .A(round_reg[842]), .B(n2339), .Z(n2586) );
  ANDN U2817 ( .B(n2962), .A(n2800), .Z(n2961) );
  XOR U2818 ( .A(n2963), .B(n2590), .Z(out[467]) );
  XOR U2819 ( .A(round_reg[841]), .B(n2343), .Z(n2590) );
  ANDN U2820 ( .B(n2964), .A(n2802), .Z(n2963) );
  XOR U2821 ( .A(n2965), .B(n2594), .Z(out[466]) );
  XOR U2822 ( .A(round_reg[840]), .B(n2351), .Z(n2594) );
  ANDN U2823 ( .B(n2966), .A(n2804), .Z(n2965) );
  XOR U2824 ( .A(n2967), .B(n2598), .Z(out[465]) );
  IV U2825 ( .A(n2811), .Z(n2598) );
  XNOR U2826 ( .A(round_reg[839]), .B(n2355), .Z(n2811) );
  NOR U2827 ( .A(n2968), .B(n2810), .Z(n2967) );
  XOR U2828 ( .A(n2969), .B(n2602), .Z(out[464]) );
  XOR U2829 ( .A(round_reg[838]), .B(n2359), .Z(n2602) );
  NOR U2830 ( .A(n2970), .B(n2813), .Z(n2969) );
  XOR U2831 ( .A(n2971), .B(n2606), .Z(out[463]) );
  XOR U2832 ( .A(round_reg[837]), .B(n2363), .Z(n2606) );
  NOR U2833 ( .A(n2972), .B(n2815), .Z(n2971) );
  XOR U2834 ( .A(n2973), .B(n2610), .Z(out[462]) );
  XOR U2835 ( .A(round_reg[836]), .B(n2367), .Z(n2610) );
  NOR U2836 ( .A(n2974), .B(n2817), .Z(n2973) );
  XOR U2837 ( .A(n2975), .B(n2618), .Z(out[461]) );
  XOR U2838 ( .A(round_reg[835]), .B(n2371), .Z(n2618) );
  NOR U2839 ( .A(n2976), .B(n2819), .Z(n2975) );
  XOR U2840 ( .A(n2977), .B(n2622), .Z(out[460]) );
  XOR U2841 ( .A(round_reg[834]), .B(n2375), .Z(n2622) );
  NOR U2842 ( .A(n2978), .B(n2821), .Z(n2977) );
  XNOR U2843 ( .A(n2979), .B(n2980), .Z(out[45]) );
  AND U2844 ( .A(n2981), .B(n2982), .Z(n2979) );
  XOR U2845 ( .A(n2983), .B(n2626), .Z(out[459]) );
  XOR U2846 ( .A(round_reg[833]), .B(n2379), .Z(n2626) );
  NOR U2847 ( .A(n2984), .B(n2823), .Z(n2983) );
  XOR U2848 ( .A(n2985), .B(n2630), .Z(out[458]) );
  XOR U2849 ( .A(round_reg[832]), .B(n2383), .Z(n2630) );
  ANDN U2850 ( .B(n2986), .A(n2825), .Z(n2985) );
  XOR U2851 ( .A(n2987), .B(n2634), .Z(out[457]) );
  XOR U2852 ( .A(round_reg[895]), .B(n2387), .Z(n2634) );
  NOR U2853 ( .A(n2988), .B(n2827), .Z(n2987) );
  XOR U2854 ( .A(n2989), .B(n2638), .Z(out[456]) );
  XOR U2855 ( .A(round_reg[894]), .B(n2990), .Z(n2638) );
  XOR U2856 ( .A(n2992), .B(n2642), .Z(out[455]) );
  XOR U2857 ( .A(round_reg[893]), .B(n2993), .Z(n2642) );
  XOR U2858 ( .A(n2995), .B(n2646), .Z(out[454]) );
  IV U2859 ( .A(n2838), .Z(n2646) );
  XNOR U2860 ( .A(round_reg[892]), .B(n2115), .Z(n2838) );
  XOR U2861 ( .A(n2997), .B(n2650), .Z(out[453]) );
  IV U2862 ( .A(n2841), .Z(n2650) );
  XNOR U2863 ( .A(round_reg[891]), .B(n2119), .Z(n2841) );
  XOR U2864 ( .A(n2999), .B(n2654), .Z(out[452]) );
  XOR U2865 ( .A(round_reg[890]), .B(n3000), .Z(n2654) );
  XOR U2866 ( .A(n3002), .B(n2662), .Z(out[451]) );
  XOR U2867 ( .A(round_reg[889]), .B(n2135), .Z(n2662) );
  ANDN U2868 ( .B(n3003), .A(n2845), .Z(n3002) );
  XOR U2869 ( .A(n3004), .B(n2666), .Z(out[450]) );
  XOR U2870 ( .A(round_reg[888]), .B(n2139), .Z(n2666) );
  ANDN U2871 ( .B(n3005), .A(n2847), .Z(n3004) );
  XNOR U2872 ( .A(n3006), .B(n3007), .Z(out[44]) );
  AND U2873 ( .A(n3008), .B(n3009), .Z(n3006) );
  XOR U2874 ( .A(n3010), .B(n2670), .Z(out[449]) );
  XOR U2875 ( .A(round_reg[887]), .B(n2143), .Z(n2670) );
  ANDN U2876 ( .B(n3011), .A(n2849), .Z(n3010) );
  XOR U2877 ( .A(n3012), .B(n2674), .Z(out[448]) );
  XOR U2878 ( .A(round_reg[886]), .B(n2147), .Z(n2674) );
  ANDN U2879 ( .B(n3013), .A(n2851), .Z(n3012) );
  XOR U2880 ( .A(n3014), .B(n2676), .Z(out[447]) );
  XOR U2881 ( .A(round_reg[496]), .B(n2150), .Z(n2676) );
  NOR U2882 ( .A(n2853), .B(n2393), .Z(n3014) );
  XOR U2883 ( .A(n3015), .B(n2678), .Z(out[446]) );
  XOR U2884 ( .A(round_reg[495]), .B(n2154), .Z(n2678) );
  NOR U2885 ( .A(n2855), .B(n2397), .Z(n3015) );
  XOR U2886 ( .A(n3016), .B(n2680), .Z(out[445]) );
  XOR U2887 ( .A(round_reg[494]), .B(n2158), .Z(n2680) );
  NOR U2888 ( .A(n2861), .B(n2401), .Z(n3016) );
  XOR U2889 ( .A(n3017), .B(n2682), .Z(out[444]) );
  XOR U2890 ( .A(round_reg[493]), .B(n2162), .Z(n2682) );
  NOR U2891 ( .A(n2863), .B(n2405), .Z(n3017) );
  XOR U2892 ( .A(n3018), .B(n2684), .Z(out[443]) );
  XOR U2893 ( .A(round_reg[492]), .B(n2166), .Z(n2684) );
  NOR U2894 ( .A(n2865), .B(n2409), .Z(n3018) );
  XOR U2895 ( .A(n3019), .B(n2686), .Z(out[442]) );
  XOR U2896 ( .A(round_reg[491]), .B(n2174), .Z(n2686) );
  NOR U2897 ( .A(n2867), .B(n2413), .Z(n3019) );
  XOR U2898 ( .A(n3020), .B(n2692), .Z(out[441]) );
  XOR U2899 ( .A(round_reg[490]), .B(n2178), .Z(n2692) );
  NOR U2900 ( .A(n2869), .B(n2417), .Z(n3020) );
  XOR U2901 ( .A(n3021), .B(n2694), .Z(out[440]) );
  XOR U2902 ( .A(round_reg[489]), .B(n2182), .Z(n2694) );
  NOR U2903 ( .A(n2871), .B(n2421), .Z(n3021) );
  XNOR U2904 ( .A(n3022), .B(n3023), .Z(out[43]) );
  AND U2905 ( .A(n3024), .B(n3025), .Z(n3022) );
  XOR U2906 ( .A(n3026), .B(n2696), .Z(out[439]) );
  XOR U2907 ( .A(round_reg[488]), .B(n2186), .Z(n2696) );
  NOR U2908 ( .A(n2873), .B(n2425), .Z(n3026) );
  XOR U2909 ( .A(n3027), .B(n2699), .Z(out[438]) );
  XOR U2910 ( .A(round_reg[487]), .B(n2190), .Z(n2699) );
  NOR U2911 ( .A(n2875), .B(n2429), .Z(n3027) );
  XOR U2912 ( .A(n3028), .B(n2702), .Z(out[437]) );
  XOR U2913 ( .A(round_reg[486]), .B(n2194), .Z(n2702) );
  NOR U2914 ( .A(n2877), .B(n2437), .Z(n3028) );
  XOR U2915 ( .A(n3029), .B(n2705), .Z(out[436]) );
  XOR U2916 ( .A(round_reg[485]), .B(n2198), .Z(n2705) );
  NOR U2917 ( .A(n2441), .B(n2879), .Z(n3029) );
  XOR U2918 ( .A(n3030), .B(n2708), .Z(out[435]) );
  XOR U2919 ( .A(round_reg[484]), .B(n2202), .Z(n2708) );
  NOR U2920 ( .A(n2445), .B(n2888), .Z(n3030) );
  XOR U2921 ( .A(n3031), .B(n2711), .Z(out[434]) );
  XNOR U2922 ( .A(round_reg[483]), .B(n3032), .Z(n2711) );
  NOR U2923 ( .A(n2449), .B(n2890), .Z(n3031) );
  XOR U2924 ( .A(n3033), .B(n2714), .Z(out[433]) );
  XOR U2925 ( .A(round_reg[482]), .B(n2210), .Z(n2714) );
  ANDN U2926 ( .B(n3034), .A(n2453), .Z(n3033) );
  XOR U2927 ( .A(n3035), .B(n2717), .Z(out[432]) );
  XOR U2928 ( .A(round_reg[481]), .B(n2218), .Z(n2717) );
  ANDN U2929 ( .B(n3036), .A(n2457), .Z(n3035) );
  XOR U2930 ( .A(n3037), .B(n2724), .Z(out[431]) );
  XOR U2931 ( .A(round_reg[480]), .B(n2222), .Z(n2724) );
  ANDN U2932 ( .B(n3038), .A(n2461), .Z(n3037) );
  XOR U2933 ( .A(n3039), .B(n2727), .Z(out[430]) );
  XOR U2934 ( .A(round_reg[479]), .B(n2226), .Z(n2727) );
  ANDN U2935 ( .B(n3040), .A(n2465), .Z(n3039) );
  XNOR U2936 ( .A(n3041), .B(n3042), .Z(out[42]) );
  AND U2937 ( .A(n3043), .B(n3044), .Z(n3041) );
  XOR U2938 ( .A(n3045), .B(n2730), .Z(out[429]) );
  XOR U2939 ( .A(round_reg[478]), .B(n2230), .Z(n2730) );
  ANDN U2940 ( .B(n3046), .A(n2469), .Z(n3045) );
  XOR U2941 ( .A(n3047), .B(n2733), .Z(out[428]) );
  XOR U2942 ( .A(round_reg[477]), .B(n2234), .Z(n2733) );
  ANDN U2943 ( .B(n3048), .A(n2473), .Z(n3047) );
  XOR U2944 ( .A(n3049), .B(n2736), .Z(out[427]) );
  XOR U2945 ( .A(round_reg[476]), .B(n2238), .Z(n2736) );
  ANDN U2946 ( .B(n3050), .A(n2481), .Z(n3049) );
  XOR U2947 ( .A(n3051), .B(n2739), .Z(out[426]) );
  XOR U2948 ( .A(round_reg[475]), .B(n2242), .Z(n2739) );
  ANDN U2949 ( .B(n3052), .A(n2485), .Z(n3051) );
  XOR U2950 ( .A(n3053), .B(n2741), .Z(out[425]) );
  XOR U2951 ( .A(round_reg[474]), .B(n2246), .Z(n2741) );
  ANDN U2952 ( .B(n3054), .A(n2489), .Z(n3053) );
  XOR U2953 ( .A(n3055), .B(n2743), .Z(out[424]) );
  XOR U2954 ( .A(round_reg[473]), .B(n2250), .Z(n2743) );
  ANDN U2955 ( .B(n3056), .A(n2493), .Z(n3055) );
  XOR U2956 ( .A(n3057), .B(n2745), .Z(out[423]) );
  XOR U2957 ( .A(round_reg[472]), .B(n2254), .Z(n2745) );
  ANDN U2958 ( .B(n3058), .A(n2497), .Z(n3057) );
  XOR U2959 ( .A(n3059), .B(n2747), .Z(out[422]) );
  XOR U2960 ( .A(round_reg[471]), .B(n2262), .Z(n2747) );
  ANDN U2961 ( .B(n3060), .A(n2501), .Z(n3059) );
  XOR U2962 ( .A(n3061), .B(n2753), .Z(out[421]) );
  XOR U2963 ( .A(round_reg[470]), .B(n2266), .Z(n2753) );
  ANDN U2964 ( .B(n3062), .A(n2505), .Z(n3061) );
  XOR U2965 ( .A(n3063), .B(n2756), .Z(out[420]) );
  XOR U2966 ( .A(round_reg[469]), .B(n2270), .Z(n2756) );
  XNOR U2967 ( .A(n3064), .B(n3065), .Z(out[41]) );
  AND U2968 ( .A(n3066), .B(n3067), .Z(n3064) );
  XOR U2969 ( .A(n3068), .B(n2759), .Z(out[419]) );
  XOR U2970 ( .A(round_reg[468]), .B(n2274), .Z(n2759) );
  XOR U2971 ( .A(n3069), .B(n2762), .Z(out[418]) );
  XOR U2972 ( .A(round_reg[467]), .B(n2278), .Z(n2762) );
  XOR U2973 ( .A(n3070), .B(n2765), .Z(out[417]) );
  XOR U2974 ( .A(round_reg[466]), .B(n2282), .Z(n2765) );
  XOR U2975 ( .A(n3071), .B(n2768), .Z(out[416]) );
  XOR U2976 ( .A(round_reg[465]), .B(n2286), .Z(n2768) );
  XOR U2977 ( .A(n3072), .B(n2771), .Z(out[415]) );
  XOR U2978 ( .A(round_reg[464]), .B(n2290), .Z(n2771) );
  XOR U2979 ( .A(n3073), .B(n2774), .Z(out[414]) );
  XOR U2980 ( .A(round_reg[463]), .B(n2294), .Z(n2774) );
  XOR U2981 ( .A(n3074), .B(n2777), .Z(out[413]) );
  XOR U2982 ( .A(round_reg[462]), .B(n2298), .Z(n2777) );
  ANDN U2983 ( .B(n2940), .A(n2541), .Z(n3074) );
  IV U2984 ( .A(n3075), .Z(n2940) );
  XOR U2985 ( .A(n3076), .B(n2780), .Z(out[412]) );
  XOR U2986 ( .A(round_reg[461]), .B(n2306), .Z(n2780) );
  ANDN U2987 ( .B(n2942), .A(n2545), .Z(n3076) );
  IV U2988 ( .A(n3077), .Z(n2942) );
  XOR U2989 ( .A(n3078), .B(n2786), .Z(out[411]) );
  XOR U2990 ( .A(round_reg[460]), .B(n2310), .Z(n2786) );
  ANDN U2991 ( .B(n2944), .A(n2549), .Z(n3078) );
  IV U2992 ( .A(n3079), .Z(n2944) );
  XOR U2993 ( .A(n3080), .B(n2788), .Z(out[410]) );
  XOR U2994 ( .A(round_reg[459]), .B(n2314), .Z(n2788) );
  ANDN U2995 ( .B(n3081), .A(n2553), .Z(n3080) );
  XNOR U2996 ( .A(n3082), .B(n3083), .Z(out[40]) );
  XOR U2997 ( .A(n3086), .B(n2790), .Z(out[409]) );
  XOR U2998 ( .A(round_reg[458]), .B(n2318), .Z(n2790) );
  NOR U2999 ( .A(n2948), .B(n2557), .Z(n3086) );
  XOR U3000 ( .A(n3087), .B(n2792), .Z(out[408]) );
  XOR U3001 ( .A(round_reg[457]), .B(n2322), .Z(n2792) );
  ANDN U3002 ( .B(n3088), .A(n2561), .Z(n3087) );
  XOR U3003 ( .A(n3089), .B(n2794), .Z(out[407]) );
  XOR U3004 ( .A(round_reg[456]), .B(n2326), .Z(n2794) );
  ANDN U3005 ( .B(n3090), .A(n2572), .Z(n3089) );
  XOR U3006 ( .A(n3091), .B(n2796), .Z(out[406]) );
  XOR U3007 ( .A(round_reg[455]), .B(n2330), .Z(n2796) );
  ANDN U3008 ( .B(n3092), .A(n2576), .Z(n3091) );
  XOR U3009 ( .A(n3093), .B(n2798), .Z(out[405]) );
  XOR U3010 ( .A(round_reg[454]), .B(n2334), .Z(n2798) );
  ANDN U3011 ( .B(n3094), .A(n2580), .Z(n3093) );
  XOR U3012 ( .A(n3095), .B(n2800), .Z(out[404]) );
  XOR U3013 ( .A(round_reg[453]), .B(n2338), .Z(n2800) );
  ANDN U3014 ( .B(n3096), .A(n2584), .Z(n3095) );
  XOR U3015 ( .A(n3097), .B(n2802), .Z(out[403]) );
  XOR U3016 ( .A(round_reg[452]), .B(n2342), .Z(n2802) );
  ANDN U3017 ( .B(n3098), .A(n2588), .Z(n3097) );
  XOR U3018 ( .A(n3099), .B(n2804), .Z(out[402]) );
  XOR U3019 ( .A(round_reg[451]), .B(n2350), .Z(n2804) );
  XOR U3020 ( .A(n3100), .B(n2810), .Z(out[401]) );
  XOR U3021 ( .A(round_reg[450]), .B(n2354), .Z(n2810) );
  ANDN U3022 ( .B(n2968), .A(n2596), .Z(n3100) );
  IV U3023 ( .A(n3101), .Z(n2968) );
  XOR U3024 ( .A(n3102), .B(n2813), .Z(out[400]) );
  XOR U3025 ( .A(round_reg[449]), .B(n2358), .Z(n2813) );
  ANDN U3026 ( .B(n2970), .A(n2600), .Z(n3102) );
  IV U3027 ( .A(n3103), .Z(n2970) );
  XNOR U3028 ( .A(n3104), .B(n2214), .Z(out[3]) );
  AND U3029 ( .A(n3105), .B(n3106), .Z(n3104) );
  XNOR U3030 ( .A(n3107), .B(n3108), .Z(out[39]) );
  XOR U3031 ( .A(n3111), .B(n2815), .Z(out[399]) );
  XOR U3032 ( .A(round_reg[448]), .B(n2362), .Z(n2815) );
  ANDN U3033 ( .B(n2972), .A(n2604), .Z(n3111) );
  IV U3034 ( .A(n3112), .Z(n2972) );
  XOR U3035 ( .A(n3113), .B(n2817), .Z(out[398]) );
  XOR U3036 ( .A(round_reg[511]), .B(n2366), .Z(n2817) );
  ANDN U3037 ( .B(n2974), .A(n2608), .Z(n3113) );
  IV U3038 ( .A(n3114), .Z(n2974) );
  XOR U3039 ( .A(n3115), .B(n2819), .Z(out[397]) );
  XOR U3040 ( .A(round_reg[510]), .B(n2370), .Z(n2819) );
  ANDN U3041 ( .B(n2976), .A(n2616), .Z(n3115) );
  IV U3042 ( .A(n3116), .Z(n2976) );
  XOR U3043 ( .A(n3117), .B(n2821), .Z(out[396]) );
  XOR U3044 ( .A(round_reg[509]), .B(n2374), .Z(n2821) );
  ANDN U3045 ( .B(n2978), .A(n2620), .Z(n3117) );
  IV U3046 ( .A(n3118), .Z(n2978) );
  XOR U3047 ( .A(n3119), .B(n2823), .Z(out[395]) );
  XOR U3048 ( .A(round_reg[508]), .B(n2378), .Z(n2823) );
  ANDN U3049 ( .B(n2984), .A(n2624), .Z(n3119) );
  IV U3050 ( .A(n3120), .Z(n2984) );
  XOR U3051 ( .A(n3121), .B(n2825), .Z(out[394]) );
  XOR U3052 ( .A(round_reg[507]), .B(n2382), .Z(n2825) );
  NOR U3053 ( .A(n2986), .B(n2628), .Z(n3121) );
  XOR U3054 ( .A(n3122), .B(n2827), .Z(out[393]) );
  XOR U3055 ( .A(round_reg[506]), .B(n2386), .Z(n2827) );
  ANDN U3056 ( .B(n2988), .A(n2632), .Z(n3122) );
  IV U3057 ( .A(n3123), .Z(n2988) );
  XOR U3058 ( .A(n3124), .B(n2829), .Z(out[392]) );
  XOR U3059 ( .A(round_reg[505]), .B(n2108), .Z(n2829) );
  XOR U3060 ( .A(n3125), .B(n2835), .Z(out[391]) );
  XOR U3061 ( .A(round_reg[504]), .B(n2112), .Z(n2835) );
  XOR U3062 ( .A(n3126), .B(n2837), .Z(out[390]) );
  XOR U3063 ( .A(round_reg[503]), .B(n2116), .Z(n2837) );
  XNOR U3064 ( .A(n3127), .B(n3128), .Z(out[38]) );
  XOR U3065 ( .A(n3131), .B(n2840), .Z(out[389]) );
  XOR U3066 ( .A(round_reg[502]), .B(n2120), .Z(n2840) );
  XOR U3067 ( .A(n3132), .B(n2843), .Z(out[388]) );
  XOR U3068 ( .A(round_reg[501]), .B(n2131), .Z(n2843) );
  XOR U3069 ( .A(n3133), .B(n2845), .Z(out[387]) );
  XOR U3070 ( .A(round_reg[500]), .B(n2134), .Z(n2845) );
  NOR U3071 ( .A(n3003), .B(n2660), .Z(n3133) );
  XOR U3072 ( .A(n3134), .B(n2847), .Z(out[386]) );
  XOR U3073 ( .A(round_reg[499]), .B(n2138), .Z(n2847) );
  NOR U3074 ( .A(n3005), .B(n2664), .Z(n3134) );
  XOR U3075 ( .A(n3135), .B(n2849), .Z(out[385]) );
  XOR U3076 ( .A(round_reg[498]), .B(n2142), .Z(n2849) );
  NOR U3077 ( .A(n3011), .B(n2668), .Z(n3135) );
  XOR U3078 ( .A(n3136), .B(n2851), .Z(out[384]) );
  XOR U3079 ( .A(round_reg[497]), .B(n2146), .Z(n2851) );
  NOR U3080 ( .A(n3013), .B(n2672), .Z(n3136) );
  XOR U3081 ( .A(n3137), .B(n2853), .Z(out[383]) );
  XOR U3082 ( .A(round_reg[71]), .B(n1817), .Z(n2853) );
  ANDN U3083 ( .B(n2393), .A(n2394), .Z(n3137) );
  XNOR U3084 ( .A(round_reg[1243]), .B(n2189), .Z(n2394) );
  XNOR U3085 ( .A(round_reg[1316]), .B(n1996), .Z(n2393) );
  XOR U3086 ( .A(n3138), .B(n2855), .Z(out[382]) );
  XOR U3087 ( .A(round_reg[70]), .B(n1828), .Z(n2855) );
  ANDN U3088 ( .B(n2397), .A(n2398), .Z(n3138) );
  XNOR U3089 ( .A(round_reg[1242]), .B(n2193), .Z(n2398) );
  XNOR U3090 ( .A(round_reg[1315]), .B(n1999), .Z(n2397) );
  XOR U3091 ( .A(n3139), .B(n2861), .Z(out[381]) );
  XOR U3092 ( .A(round_reg[69]), .B(n1831), .Z(n2861) );
  ANDN U3093 ( .B(n2401), .A(n2402), .Z(n3139) );
  XNOR U3094 ( .A(round_reg[1241]), .B(n2197), .Z(n2402) );
  XNOR U3095 ( .A(round_reg[1314]), .B(n2002), .Z(n2401) );
  XOR U3096 ( .A(n3140), .B(n2863), .Z(out[380]) );
  XOR U3097 ( .A(round_reg[68]), .B(n1834), .Z(n2863) );
  ANDN U3098 ( .B(n2405), .A(n2406), .Z(n3140) );
  XNOR U3099 ( .A(round_reg[1240]), .B(n2201), .Z(n2406) );
  XNOR U3100 ( .A(round_reg[1313]), .B(n2004), .Z(n2405) );
  XNOR U3101 ( .A(n3141), .B(n3142), .Z(out[37]) );
  XOR U3102 ( .A(n3145), .B(n2865), .Z(out[379]) );
  XOR U3103 ( .A(round_reg[67]), .B(n1837), .Z(n2865) );
  ANDN U3104 ( .B(n2409), .A(n2410), .Z(n3145) );
  XNOR U3105 ( .A(round_reg[1239]), .B(n2205), .Z(n2410) );
  XNOR U3106 ( .A(round_reg[1312]), .B(n2006), .Z(n2409) );
  XOR U3107 ( .A(n3146), .B(n2867), .Z(out[378]) );
  XOR U3108 ( .A(round_reg[66]), .B(n1840), .Z(n2867) );
  ANDN U3109 ( .B(n2413), .A(n2414), .Z(n3146) );
  XNOR U3110 ( .A(round_reg[1238]), .B(n2209), .Z(n2414) );
  XNOR U3111 ( .A(round_reg[1311]), .B(n2008), .Z(n2413) );
  XOR U3112 ( .A(n3147), .B(n2869), .Z(out[377]) );
  XOR U3113 ( .A(round_reg[65]), .B(n1843), .Z(n2869) );
  ANDN U3114 ( .B(n2417), .A(n2418), .Z(n3147) );
  XNOR U3115 ( .A(round_reg[1237]), .B(n2217), .Z(n2418) );
  XNOR U3116 ( .A(round_reg[1310]), .B(n2010), .Z(n2417) );
  XOR U3117 ( .A(n3148), .B(n2871), .Z(out[376]) );
  XOR U3118 ( .A(round_reg[64]), .B(n1846), .Z(n2871) );
  ANDN U3119 ( .B(n2421), .A(n2422), .Z(n3148) );
  XNOR U3120 ( .A(round_reg[1236]), .B(n2221), .Z(n2422) );
  XNOR U3121 ( .A(round_reg[1309]), .B(n2012), .Z(n2421) );
  XOR U3122 ( .A(n3149), .B(n2873), .Z(out[375]) );
  XOR U3123 ( .A(round_reg[127]), .B(n1849), .Z(n2873) );
  ANDN U3124 ( .B(n2425), .A(n2426), .Z(n3149) );
  XNOR U3125 ( .A(round_reg[1235]), .B(n2225), .Z(n2426) );
  XNOR U3126 ( .A(round_reg[1308]), .B(n2014), .Z(n2425) );
  XOR U3127 ( .A(n3150), .B(n2875), .Z(out[374]) );
  XOR U3128 ( .A(round_reg[126]), .B(n1852), .Z(n2875) );
  ANDN U3129 ( .B(n2429), .A(n2430), .Z(n3150) );
  XNOR U3130 ( .A(round_reg[1234]), .B(n2229), .Z(n2430) );
  XNOR U3131 ( .A(round_reg[1307]), .B(n2020), .Z(n2429) );
  XOR U3132 ( .A(n3151), .B(n2877), .Z(out[373]) );
  XOR U3133 ( .A(round_reg[125]), .B(n1855), .Z(n2877) );
  ANDN U3134 ( .B(n2437), .A(n2438), .Z(n3151) );
  XNOR U3135 ( .A(round_reg[1233]), .B(n2233), .Z(n2438) );
  XNOR U3136 ( .A(round_reg[1306]), .B(n2022), .Z(n2437) );
  XOR U3137 ( .A(n3152), .B(n2879), .Z(out[372]) );
  XOR U3138 ( .A(round_reg[124]), .B(n1862), .Z(n2879) );
  ANDN U3139 ( .B(n2441), .A(n2442), .Z(n3152) );
  XNOR U3140 ( .A(round_reg[1232]), .B(n2237), .Z(n2442) );
  XNOR U3141 ( .A(round_reg[1305]), .B(n2025), .Z(n2441) );
  XOR U3142 ( .A(n3153), .B(n2888), .Z(out[371]) );
  XOR U3143 ( .A(round_reg[123]), .B(n1865), .Z(n2888) );
  ANDN U3144 ( .B(n2445), .A(n2446), .Z(n3153) );
  XNOR U3145 ( .A(round_reg[1231]), .B(n2241), .Z(n2446) );
  XNOR U3146 ( .A(round_reg[1304]), .B(n2028), .Z(n2445) );
  XOR U3147 ( .A(n3154), .B(n2890), .Z(out[370]) );
  XOR U3148 ( .A(round_reg[122]), .B(n1868), .Z(n2890) );
  ANDN U3149 ( .B(n2449), .A(n2450), .Z(n3154) );
  XNOR U3150 ( .A(round_reg[1230]), .B(n2245), .Z(n2450) );
  XNOR U3151 ( .A(round_reg[1303]), .B(n2031), .Z(n2449) );
  XNOR U3152 ( .A(n3155), .B(n3156), .Z(out[36]) );
  XOR U3153 ( .A(n3159), .B(n2892), .Z(out[369]) );
  IV U3154 ( .A(n3034), .Z(n2892) );
  XNOR U3155 ( .A(round_reg[121]), .B(n1871), .Z(n3034) );
  ANDN U3156 ( .B(n2453), .A(n2454), .Z(n3159) );
  XNOR U3157 ( .A(round_reg[1229]), .B(n2249), .Z(n2454) );
  XNOR U3158 ( .A(round_reg[1302]), .B(n2034), .Z(n2453) );
  XOR U3159 ( .A(n3160), .B(n2894), .Z(out[368]) );
  IV U3160 ( .A(n3036), .Z(n2894) );
  XNOR U3161 ( .A(round_reg[120]), .B(n1874), .Z(n3036) );
  ANDN U3162 ( .B(n2457), .A(n2458), .Z(n3160) );
  XNOR U3163 ( .A(round_reg[1228]), .B(n2253), .Z(n2458) );
  XNOR U3164 ( .A(round_reg[1301]), .B(n2037), .Z(n2457) );
  XOR U3165 ( .A(n3161), .B(n2896), .Z(out[367]) );
  IV U3166 ( .A(n3038), .Z(n2896) );
  XNOR U3167 ( .A(round_reg[119]), .B(n1877), .Z(n3038) );
  ANDN U3168 ( .B(n2461), .A(n2462), .Z(n3161) );
  XNOR U3169 ( .A(round_reg[1227]), .B(n2261), .Z(n2462) );
  XNOR U3170 ( .A(round_reg[1300]), .B(n2040), .Z(n2461) );
  XOR U3171 ( .A(n3162), .B(n2898), .Z(out[366]) );
  IV U3172 ( .A(n3040), .Z(n2898) );
  XNOR U3173 ( .A(round_reg[118]), .B(n1880), .Z(n3040) );
  ANDN U3174 ( .B(n2465), .A(n2466), .Z(n3162) );
  XNOR U3175 ( .A(round_reg[1226]), .B(n2265), .Z(n2466) );
  XNOR U3176 ( .A(round_reg[1299]), .B(n2042), .Z(n2465) );
  XOR U3177 ( .A(n3163), .B(n2900), .Z(out[365]) );
  IV U3178 ( .A(n3046), .Z(n2900) );
  XNOR U3179 ( .A(round_reg[117]), .B(n1883), .Z(n3046) );
  ANDN U3180 ( .B(n2469), .A(n2470), .Z(n3163) );
  XNOR U3181 ( .A(round_reg[1225]), .B(n2269), .Z(n2470) );
  XNOR U3182 ( .A(round_reg[1298]), .B(n2044), .Z(n2469) );
  XOR U3183 ( .A(n3164), .B(n2902), .Z(out[364]) );
  IV U3184 ( .A(n3048), .Z(n2902) );
  XNOR U3185 ( .A(round_reg[116]), .B(n1886), .Z(n3048) );
  ANDN U3186 ( .B(n2473), .A(n2474), .Z(n3164) );
  XNOR U3187 ( .A(round_reg[1224]), .B(n2273), .Z(n2474) );
  XNOR U3188 ( .A(round_reg[1297]), .B(n2048), .Z(n2473) );
  XOR U3189 ( .A(n3165), .B(n2904), .Z(out[363]) );
  IV U3190 ( .A(n3050), .Z(n2904) );
  XNOR U3191 ( .A(round_reg[115]), .B(n1889), .Z(n3050) );
  ANDN U3192 ( .B(n2481), .A(n2482), .Z(n3165) );
  XNOR U3193 ( .A(round_reg[1223]), .B(n2277), .Z(n2482) );
  XNOR U3194 ( .A(round_reg[1296]), .B(n2050), .Z(n2481) );
  XOR U3195 ( .A(n3166), .B(n2906), .Z(out[362]) );
  IV U3196 ( .A(n3052), .Z(n2906) );
  XNOR U3197 ( .A(round_reg[114]), .B(n1896), .Z(n3052) );
  ANDN U3198 ( .B(n2485), .A(n2486), .Z(n3166) );
  XNOR U3199 ( .A(round_reg[1222]), .B(n2281), .Z(n2486) );
  XNOR U3200 ( .A(round_reg[1295]), .B(n2052), .Z(n2485) );
  XOR U3201 ( .A(n3167), .B(n2912), .Z(out[361]) );
  IV U3202 ( .A(n3054), .Z(n2912) );
  XNOR U3203 ( .A(round_reg[113]), .B(n1899), .Z(n3054) );
  ANDN U3204 ( .B(n2489), .A(n2490), .Z(n3167) );
  XNOR U3205 ( .A(round_reg[1221]), .B(n2285), .Z(n2490) );
  XNOR U3206 ( .A(round_reg[1294]), .B(n2054), .Z(n2489) );
  XOR U3207 ( .A(n3168), .B(n2914), .Z(out[360]) );
  IV U3208 ( .A(n3056), .Z(n2914) );
  XNOR U3209 ( .A(round_reg[112]), .B(n1902), .Z(n3056) );
  ANDN U3210 ( .B(n2493), .A(n2494), .Z(n3168) );
  XNOR U3211 ( .A(round_reg[1220]), .B(n2289), .Z(n2494) );
  XNOR U3212 ( .A(round_reg[1293]), .B(n2056), .Z(n2493) );
  XOR U3213 ( .A(n3169), .B(n1058), .Z(out[35]) );
  ANDN U3214 ( .B(n3170), .A(n1057), .Z(n3169) );
  XOR U3215 ( .A(n3171), .B(n2916), .Z(out[359]) );
  IV U3216 ( .A(n3058), .Z(n2916) );
  XNOR U3217 ( .A(round_reg[111]), .B(n1905), .Z(n3058) );
  ANDN U3218 ( .B(n2497), .A(n2498), .Z(n3171) );
  XNOR U3219 ( .A(round_reg[1219]), .B(n2293), .Z(n2498) );
  XNOR U3220 ( .A(round_reg[1292]), .B(n2058), .Z(n2497) );
  XOR U3221 ( .A(n3172), .B(n2918), .Z(out[358]) );
  IV U3222 ( .A(n3060), .Z(n2918) );
  XNOR U3223 ( .A(round_reg[110]), .B(n1908), .Z(n3060) );
  ANDN U3224 ( .B(n2501), .A(n2502), .Z(n3172) );
  XNOR U3225 ( .A(round_reg[1218]), .B(n2297), .Z(n2502) );
  XNOR U3226 ( .A(round_reg[1291]), .B(n2060), .Z(n2501) );
  XOR U3227 ( .A(n3173), .B(n2920), .Z(out[357]) );
  IV U3228 ( .A(n3062), .Z(n2920) );
  XNOR U3229 ( .A(round_reg[109]), .B(n1911), .Z(n3062) );
  ANDN U3230 ( .B(n2505), .A(n2506), .Z(n3173) );
  XNOR U3231 ( .A(round_reg[1217]), .B(n2305), .Z(n2506) );
  XNOR U3232 ( .A(round_reg[1290]), .B(n2062), .Z(n2505) );
  XOR U3233 ( .A(n3174), .B(n2922), .Z(out[356]) );
  XNOR U3234 ( .A(round_reg[108]), .B(n1914), .Z(n2922) );
  ANDN U3235 ( .B(n2509), .A(n2510), .Z(n3174) );
  XNOR U3236 ( .A(round_reg[1216]), .B(n2309), .Z(n2510) );
  XNOR U3237 ( .A(round_reg[1289]), .B(n2064), .Z(n2509) );
  XOR U3238 ( .A(n3175), .B(n2924), .Z(out[355]) );
  XNOR U3239 ( .A(round_reg[107]), .B(n1917), .Z(n2924) );
  ANDN U3240 ( .B(n2513), .A(n2514), .Z(n3175) );
  XNOR U3241 ( .A(round_reg[1279]), .B(n2313), .Z(n2514) );
  XNOR U3242 ( .A(round_reg[1288]), .B(n2066), .Z(n2513) );
  XOR U3243 ( .A(n3176), .B(n2926), .Z(out[354]) );
  XNOR U3244 ( .A(round_reg[106]), .B(n1920), .Z(n2926) );
  ANDN U3245 ( .B(n2517), .A(n2518), .Z(n3176) );
  XNOR U3246 ( .A(round_reg[1278]), .B(n2317), .Z(n2518) );
  XNOR U3247 ( .A(round_reg[1287]), .B(n2070), .Z(n2517) );
  XOR U3248 ( .A(n3177), .B(n2928), .Z(out[353]) );
  XNOR U3249 ( .A(round_reg[105]), .B(n1923), .Z(n2928) );
  ANDN U3250 ( .B(n2525), .A(n2526), .Z(n3177) );
  XNOR U3251 ( .A(round_reg[1277]), .B(n2321), .Z(n2526) );
  XNOR U3252 ( .A(round_reg[1286]), .B(n2072), .Z(n2525) );
  XOR U3253 ( .A(n3178), .B(n2930), .Z(out[352]) );
  XNOR U3254 ( .A(round_reg[104]), .B(n1930), .Z(n2930) );
  ANDN U3255 ( .B(n2529), .A(n2530), .Z(n3178) );
  XNOR U3256 ( .A(round_reg[1276]), .B(n2325), .Z(n2530) );
  XNOR U3257 ( .A(round_reg[1285]), .B(n2074), .Z(n2529) );
  XOR U3258 ( .A(n3179), .B(n2936), .Z(out[351]) );
  XNOR U3259 ( .A(round_reg[103]), .B(n1933), .Z(n2936) );
  ANDN U3260 ( .B(n2533), .A(n2534), .Z(n3179) );
  XNOR U3261 ( .A(round_reg[1275]), .B(n2329), .Z(n2534) );
  XNOR U3262 ( .A(round_reg[1284]), .B(n2076), .Z(n2533) );
  XOR U3263 ( .A(n3180), .B(n2938), .Z(out[350]) );
  XNOR U3264 ( .A(round_reg[102]), .B(n1712), .Z(n2938) );
  ANDN U3265 ( .B(n2537), .A(n2538), .Z(n3180) );
  XNOR U3266 ( .A(round_reg[1274]), .B(n2333), .Z(n2538) );
  XNOR U3267 ( .A(round_reg[1283]), .B(n2078), .Z(n2537) );
  XOR U3268 ( .A(n3181), .B(n1102), .Z(out[34]) );
  ANDN U3269 ( .B(n3182), .A(n1101), .Z(n3181) );
  XOR U3270 ( .A(n3183), .B(n3075), .Z(out[349]) );
  XNOR U3271 ( .A(round_reg[101]), .B(n1715), .Z(n3075) );
  ANDN U3272 ( .B(n2541), .A(n2542), .Z(n3183) );
  XNOR U3273 ( .A(round_reg[1273]), .B(n2337), .Z(n2542) );
  XNOR U3274 ( .A(round_reg[1282]), .B(n2080), .Z(n2541) );
  XOR U3275 ( .A(n3184), .B(n3077), .Z(out[348]) );
  XNOR U3276 ( .A(round_reg[100]), .B(n1722), .Z(n3077) );
  ANDN U3277 ( .B(n2545), .A(n2546), .Z(n3184) );
  XNOR U3278 ( .A(round_reg[1272]), .B(n2341), .Z(n2546) );
  XNOR U3279 ( .A(round_reg[1281]), .B(n2082), .Z(n2545) );
  XOR U3280 ( .A(n3185), .B(n3079), .Z(out[347]) );
  XNOR U3281 ( .A(round_reg[99]), .B(n1725), .Z(n3079) );
  ANDN U3282 ( .B(n2549), .A(n2550), .Z(n3185) );
  XNOR U3283 ( .A(round_reg[1271]), .B(n2349), .Z(n2550) );
  XNOR U3284 ( .A(round_reg[1280]), .B(n2084), .Z(n2549) );
  XOR U3285 ( .A(n3186), .B(n2946), .Z(out[346]) );
  IV U3286 ( .A(n3081), .Z(n2946) );
  XNOR U3287 ( .A(round_reg[98]), .B(n1728), .Z(n3081) );
  ANDN U3288 ( .B(n2553), .A(n2554), .Z(n3186) );
  XNOR U3289 ( .A(round_reg[1270]), .B(n2353), .Z(n2554) );
  XOR U3290 ( .A(round_reg[1343]), .B(n2086), .Z(n2553) );
  XOR U3291 ( .A(n3187), .B(n2948), .Z(out[345]) );
  XOR U3292 ( .A(round_reg[97]), .B(n1731), .Z(n2948) );
  ANDN U3293 ( .B(n2557), .A(n2558), .Z(n3187) );
  XNOR U3294 ( .A(round_reg[1269]), .B(n2357), .Z(n2558) );
  XNOR U3295 ( .A(round_reg[1342]), .B(n2088), .Z(n2557) );
  XOR U3296 ( .A(n3188), .B(n2950), .Z(out[344]) );
  IV U3297 ( .A(n3088), .Z(n2950) );
  XNOR U3298 ( .A(round_reg[96]), .B(n1734), .Z(n3088) );
  ANDN U3299 ( .B(n2561), .A(n2562), .Z(n3188) );
  XNOR U3300 ( .A(round_reg[1268]), .B(n2361), .Z(n2562) );
  XNOR U3301 ( .A(round_reg[1341]), .B(n2094), .Z(n2561) );
  XOR U3302 ( .A(n3189), .B(n2952), .Z(out[343]) );
  IV U3303 ( .A(n3090), .Z(n2952) );
  XNOR U3304 ( .A(round_reg[95]), .B(n1737), .Z(n3090) );
  ANDN U3305 ( .B(n2572), .A(n2573), .Z(n3189) );
  XNOR U3306 ( .A(round_reg[1267]), .B(n2365), .Z(n2573) );
  XNOR U3307 ( .A(round_reg[1340]), .B(n2096), .Z(n2572) );
  XOR U3308 ( .A(n3190), .B(n2954), .Z(out[342]) );
  IV U3309 ( .A(n3092), .Z(n2954) );
  XNOR U3310 ( .A(round_reg[94]), .B(n1740), .Z(n3092) );
  ANDN U3311 ( .B(n2576), .A(n2577), .Z(n3190) );
  XNOR U3312 ( .A(round_reg[1266]), .B(n2369), .Z(n2577) );
  XNOR U3313 ( .A(round_reg[1339]), .B(n2098), .Z(n2576) );
  XOR U3314 ( .A(n3191), .B(n2960), .Z(out[341]) );
  IV U3315 ( .A(n3094), .Z(n2960) );
  XNOR U3316 ( .A(round_reg[93]), .B(n1743), .Z(n3094) );
  ANDN U3317 ( .B(n2580), .A(n2581), .Z(n3191) );
  XNOR U3318 ( .A(round_reg[1265]), .B(n2373), .Z(n2581) );
  XNOR U3319 ( .A(round_reg[1338]), .B(n2100), .Z(n2580) );
  XOR U3320 ( .A(n3192), .B(n2962), .Z(out[340]) );
  IV U3321 ( .A(n3096), .Z(n2962) );
  XNOR U3322 ( .A(round_reg[92]), .B(n1746), .Z(n3096) );
  ANDN U3323 ( .B(n2584), .A(n2585), .Z(n3192) );
  XNOR U3324 ( .A(round_reg[1264]), .B(n2377), .Z(n2585) );
  XNOR U3325 ( .A(round_reg[1337]), .B(n2102), .Z(n2584) );
  XNOR U3326 ( .A(n3193), .B(n1146), .Z(out[33]) );
  ANDN U3327 ( .B(n3194), .A(n1145), .Z(n3193) );
  XOR U3328 ( .A(n3195), .B(n2964), .Z(out[339]) );
  IV U3329 ( .A(n3098), .Z(n2964) );
  XNOR U3330 ( .A(round_reg[91]), .B(n1749), .Z(n3098) );
  ANDN U3331 ( .B(n2588), .A(n2589), .Z(n3195) );
  XNOR U3332 ( .A(round_reg[1263]), .B(n2381), .Z(n2589) );
  XNOR U3333 ( .A(round_reg[1336]), .B(n2104), .Z(n2588) );
  XOR U3334 ( .A(n3196), .B(n2966), .Z(out[338]) );
  XNOR U3335 ( .A(round_reg[90]), .B(n1756), .Z(n2966) );
  ANDN U3336 ( .B(n2592), .A(n2593), .Z(n3196) );
  XNOR U3337 ( .A(round_reg[1262]), .B(n2385), .Z(n2593) );
  XNOR U3338 ( .A(round_reg[1335]), .B(n1936), .Z(n2592) );
  XOR U3339 ( .A(n3197), .B(n3101), .Z(out[337]) );
  XNOR U3340 ( .A(round_reg[89]), .B(n1759), .Z(n3101) );
  ANDN U3341 ( .B(n2596), .A(n2597), .Z(n3197) );
  XNOR U3342 ( .A(round_reg[1261]), .B(n2106), .Z(n2597) );
  XNOR U3343 ( .A(round_reg[1334]), .B(n1938), .Z(n2596) );
  XOR U3344 ( .A(n3198), .B(n3103), .Z(out[336]) );
  XNOR U3345 ( .A(round_reg[88]), .B(n1762), .Z(n3103) );
  ANDN U3346 ( .B(n2600), .A(n2601), .Z(n3198) );
  XNOR U3347 ( .A(round_reg[1260]), .B(n2110), .Z(n2601) );
  XNOR U3348 ( .A(round_reg[1333]), .B(n1940), .Z(n2600) );
  XOR U3349 ( .A(n3199), .B(n3112), .Z(out[335]) );
  XNOR U3350 ( .A(round_reg[87]), .B(n1765), .Z(n3112) );
  ANDN U3351 ( .B(n2604), .A(n2605), .Z(n3199) );
  XNOR U3352 ( .A(round_reg[1259]), .B(n2114), .Z(n2605) );
  XNOR U3353 ( .A(round_reg[1332]), .B(n1942), .Z(n2604) );
  XOR U3354 ( .A(n3200), .B(n3114), .Z(out[334]) );
  XNOR U3355 ( .A(round_reg[86]), .B(n1768), .Z(n3114) );
  ANDN U3356 ( .B(n2608), .A(n2609), .Z(n3200) );
  XNOR U3357 ( .A(round_reg[1258]), .B(n2118), .Z(n2609) );
  XNOR U3358 ( .A(round_reg[1331]), .B(n1945), .Z(n2608) );
  XOR U3359 ( .A(n3201), .B(n3116), .Z(out[333]) );
  XNOR U3360 ( .A(round_reg[85]), .B(n1771), .Z(n3116) );
  ANDN U3361 ( .B(n2616), .A(n2617), .Z(n3201) );
  XNOR U3362 ( .A(round_reg[1257]), .B(n2129), .Z(n2617) );
  XNOR U3363 ( .A(round_reg[1330]), .B(n1948), .Z(n2616) );
  XOR U3364 ( .A(n3202), .B(n3118), .Z(out[332]) );
  XNOR U3365 ( .A(round_reg[84]), .B(n1774), .Z(n3118) );
  ANDN U3366 ( .B(n2620), .A(n2621), .Z(n3202) );
  XNOR U3367 ( .A(round_reg[1256]), .B(n2133), .Z(n2621) );
  XNOR U3368 ( .A(round_reg[1329]), .B(n1951), .Z(n2620) );
  XOR U3369 ( .A(n3203), .B(n3120), .Z(out[331]) );
  XNOR U3370 ( .A(round_reg[83]), .B(n1777), .Z(n3120) );
  ANDN U3371 ( .B(n2624), .A(n2625), .Z(n3203) );
  XNOR U3372 ( .A(round_reg[1255]), .B(n2137), .Z(n2625) );
  XNOR U3373 ( .A(round_reg[1328]), .B(n1954), .Z(n2624) );
  XOR U3374 ( .A(n3204), .B(n2986), .Z(out[330]) );
  XOR U3375 ( .A(round_reg[82]), .B(n1780), .Z(n2986) );
  ANDN U3376 ( .B(n2628), .A(n2629), .Z(n3204) );
  XNOR U3377 ( .A(round_reg[1254]), .B(n2141), .Z(n2629) );
  XNOR U3378 ( .A(round_reg[1327]), .B(n1961), .Z(n2628) );
  XNOR U3379 ( .A(n3205), .B(n1190), .Z(out[32]) );
  ANDN U3380 ( .B(n3206), .A(n1189), .Z(n3205) );
  XOR U3381 ( .A(n3207), .B(n3123), .Z(out[329]) );
  XOR U3382 ( .A(round_reg[81]), .B(n1783), .Z(n3123) );
  ANDN U3383 ( .B(n2632), .A(n2633), .Z(n3207) );
  XNOR U3384 ( .A(round_reg[1253]), .B(n2145), .Z(n2633) );
  XNOR U3385 ( .A(round_reg[1326]), .B(n1964), .Z(n2632) );
  XOR U3386 ( .A(n3208), .B(n2991), .Z(out[328]) );
  XOR U3387 ( .A(round_reg[80]), .B(n1790), .Z(n2991) );
  ANDN U3388 ( .B(n2636), .A(n2637), .Z(n3208) );
  XNOR U3389 ( .A(round_reg[1252]), .B(n2149), .Z(n2637) );
  XNOR U3390 ( .A(round_reg[1325]), .B(n1967), .Z(n2636) );
  XOR U3391 ( .A(n3209), .B(n2994), .Z(out[327]) );
  XOR U3392 ( .A(round_reg[79]), .B(n1793), .Z(n2994) );
  ANDN U3393 ( .B(n2640), .A(n2641), .Z(n3209) );
  XNOR U3394 ( .A(round_reg[1251]), .B(n2153), .Z(n2641) );
  XNOR U3395 ( .A(round_reg[1324]), .B(n1970), .Z(n2640) );
  XOR U3396 ( .A(n3210), .B(n2996), .Z(out[326]) );
  XOR U3397 ( .A(round_reg[78]), .B(n1796), .Z(n2996) );
  ANDN U3398 ( .B(n2644), .A(n2645), .Z(n3210) );
  XNOR U3399 ( .A(round_reg[1250]), .B(n2157), .Z(n2645) );
  XNOR U3400 ( .A(round_reg[1323]), .B(n1973), .Z(n2644) );
  XOR U3401 ( .A(n3211), .B(n2998), .Z(out[325]) );
  XOR U3402 ( .A(round_reg[77]), .B(n1799), .Z(n2998) );
  ANDN U3403 ( .B(n2648), .A(n2649), .Z(n3211) );
  XNOR U3404 ( .A(round_reg[1249]), .B(n2161), .Z(n2649) );
  XNOR U3405 ( .A(round_reg[1322]), .B(n1975), .Z(n2648) );
  XOR U3406 ( .A(n3212), .B(n3001), .Z(out[324]) );
  XOR U3407 ( .A(round_reg[76]), .B(n1802), .Z(n3001) );
  ANDN U3408 ( .B(n2652), .A(n2653), .Z(n3212) );
  XNOR U3409 ( .A(round_reg[1248]), .B(n2165), .Z(n2653) );
  XNOR U3410 ( .A(round_reg[1321]), .B(n1977), .Z(n2652) );
  XOR U3411 ( .A(n3213), .B(n3003), .Z(out[323]) );
  XOR U3412 ( .A(round_reg[75]), .B(n1805), .Z(n3003) );
  ANDN U3413 ( .B(n2660), .A(n2661), .Z(n3213) );
  XNOR U3414 ( .A(round_reg[1247]), .B(n2173), .Z(n2661) );
  XNOR U3415 ( .A(round_reg[1320]), .B(n1980), .Z(n2660) );
  XOR U3416 ( .A(n3214), .B(n3005), .Z(out[322]) );
  XOR U3417 ( .A(round_reg[74]), .B(n1808), .Z(n3005) );
  ANDN U3418 ( .B(n2664), .A(n2665), .Z(n3214) );
  XNOR U3419 ( .A(round_reg[1246]), .B(n2177), .Z(n2665) );
  XNOR U3420 ( .A(round_reg[1319]), .B(n1983), .Z(n2664) );
  XOR U3421 ( .A(n3215), .B(n3011), .Z(out[321]) );
  XOR U3422 ( .A(round_reg[73]), .B(n1811), .Z(n3011) );
  ANDN U3423 ( .B(n2668), .A(n2669), .Z(n3215) );
  XNOR U3424 ( .A(round_reg[1245]), .B(n2181), .Z(n2669) );
  XNOR U3425 ( .A(round_reg[1318]), .B(n1986), .Z(n2668) );
  XOR U3426 ( .A(n3216), .B(n3013), .Z(out[320]) );
  XOR U3427 ( .A(round_reg[72]), .B(n1814), .Z(n3013) );
  ANDN U3428 ( .B(n2672), .A(n2673), .Z(n3216) );
  XNOR U3429 ( .A(round_reg[1244]), .B(n2185), .Z(n2673) );
  XNOR U3430 ( .A(round_reg[1317]), .B(n1993), .Z(n2672) );
  XNOR U3431 ( .A(n3217), .B(n1234), .Z(out[31]) );
  ANDN U3432 ( .B(n3218), .A(n1233), .Z(n3217) );
  XNOR U3433 ( .A(n3219), .B(n2390), .Z(out[319]) );
  AND U3434 ( .A(n3220), .B(n3221), .Z(n3219) );
  XNOR U3435 ( .A(n3222), .B(n2434), .Z(out[318]) );
  AND U3436 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U3437 ( .A(n3225), .B(n2478), .Z(out[317]) );
  AND U3438 ( .A(n3226), .B(n3227), .Z(n3225) );
  XNOR U3439 ( .A(n3228), .B(n2522), .Z(out[316]) );
  AND U3440 ( .A(n3229), .B(n3230), .Z(n3228) );
  XNOR U3441 ( .A(n3231), .B(n2569), .Z(out[315]) );
  AND U3442 ( .A(n3232), .B(n3233), .Z(n3231) );
  XNOR U3443 ( .A(n3234), .B(n2613), .Z(out[314]) );
  AND U3444 ( .A(n3235), .B(n3236), .Z(n3234) );
  XNOR U3445 ( .A(n3237), .B(n2657), .Z(out[313]) );
  AND U3446 ( .A(n3238), .B(n3239), .Z(n3237) );
  XNOR U3447 ( .A(n3240), .B(n2689), .Z(out[312]) );
  AND U3448 ( .A(n3241), .B(n3242), .Z(n3240) );
  XNOR U3449 ( .A(n3243), .B(n2721), .Z(out[311]) );
  AND U3450 ( .A(n3244), .B(n3245), .Z(n3243) );
  XNOR U3451 ( .A(n3246), .B(n2750), .Z(out[310]) );
  AND U3452 ( .A(n3247), .B(n3248), .Z(n3246) );
  XNOR U3453 ( .A(n3249), .B(n1277), .Z(out[30]) );
  AND U3454 ( .A(n3250), .B(n3251), .Z(n3249) );
  XNOR U3455 ( .A(n3252), .B(n2783), .Z(out[309]) );
  AND U3456 ( .A(n3253), .B(n3254), .Z(n3252) );
  XNOR U3457 ( .A(n3255), .B(n2807), .Z(out[308]) );
  AND U3458 ( .A(n3256), .B(n3257), .Z(n3255) );
  XNOR U3459 ( .A(n3258), .B(n2832), .Z(out[307]) );
  AND U3460 ( .A(n3259), .B(n3260), .Z(n3258) );
  XNOR U3461 ( .A(n3261), .B(n2858), .Z(out[306]) );
  AND U3462 ( .A(n3262), .B(n3263), .Z(n3261) );
  XNOR U3463 ( .A(n3264), .B(n2885), .Z(out[305]) );
  AND U3464 ( .A(n3265), .B(n3266), .Z(n3264) );
  XNOR U3465 ( .A(n3267), .B(n2910), .Z(out[304]) );
  ANDN U3466 ( .B(n3268), .A(n2909), .Z(n3267) );
  XNOR U3467 ( .A(n3269), .B(n2934), .Z(out[303]) );
  ANDN U3468 ( .B(n3270), .A(n2933), .Z(n3269) );
  XNOR U3469 ( .A(n3271), .B(n2958), .Z(out[302]) );
  ANDN U3470 ( .B(n3272), .A(n2957), .Z(n3271) );
  XNOR U3471 ( .A(n3273), .B(n2982), .Z(out[301]) );
  ANDN U3472 ( .B(n3274), .A(n2981), .Z(n3273) );
  XNOR U3473 ( .A(n3275), .B(n3009), .Z(out[300]) );
  ANDN U3474 ( .B(n3276), .A(n3008), .Z(n3275) );
  XNOR U3475 ( .A(n3277), .B(n2258), .Z(out[2]) );
  AND U3476 ( .A(n3278), .B(n3279), .Z(n3277) );
  XNOR U3477 ( .A(n3280), .B(n1321), .Z(out[29]) );
  AND U3478 ( .A(n3281), .B(n3282), .Z(n3280) );
  XNOR U3479 ( .A(n3283), .B(n3025), .Z(out[299]) );
  ANDN U3480 ( .B(n3284), .A(n3024), .Z(n3283) );
  XNOR U3481 ( .A(n3285), .B(n3044), .Z(out[298]) );
  ANDN U3482 ( .B(n3286), .A(n3043), .Z(n3285) );
  XNOR U3483 ( .A(n3287), .B(n3067), .Z(out[297]) );
  ANDN U3484 ( .B(n3288), .A(n3066), .Z(n3287) );
  XOR U3485 ( .A(n3289), .B(n3085), .Z(out[296]) );
  ANDN U3486 ( .B(n3290), .A(n3084), .Z(n3289) );
  XOR U3487 ( .A(n3291), .B(n3110), .Z(out[295]) );
  ANDN U3488 ( .B(n3292), .A(n3109), .Z(n3291) );
  XOR U3489 ( .A(n3293), .B(n3130), .Z(out[294]) );
  ANDN U3490 ( .B(n3294), .A(n3129), .Z(n3293) );
  XOR U3491 ( .A(n3295), .B(n3144), .Z(out[293]) );
  ANDN U3492 ( .B(n3296), .A(n3143), .Z(n3295) );
  XOR U3493 ( .A(n3297), .B(n3158), .Z(out[292]) );
  ANDN U3494 ( .B(n3298), .A(n3157), .Z(n3297) );
  XOR U3495 ( .A(n3299), .B(n1057), .Z(out[291]) );
  XOR U3496 ( .A(round_reg[1445]), .B(n2198), .Z(n1057) );
  ANDN U3497 ( .B(n3300), .A(n3170), .Z(n3299) );
  XOR U3498 ( .A(n3301), .B(n1101), .Z(out[290]) );
  XOR U3499 ( .A(round_reg[1444]), .B(n2202), .Z(n1101) );
  ANDN U3500 ( .B(n3302), .A(n3182), .Z(n3301) );
  XNOR U3501 ( .A(n3303), .B(n1365), .Z(out[28]) );
  AND U3502 ( .A(n3304), .B(n3305), .Z(n3303) );
  XOR U3503 ( .A(n3306), .B(n1145), .Z(out[289]) );
  XNOR U3504 ( .A(round_reg[1443]), .B(n3032), .Z(n1145) );
  ANDN U3505 ( .B(n3307), .A(n3194), .Z(n3306) );
  XOR U3506 ( .A(n3308), .B(n1189), .Z(out[288]) );
  XOR U3507 ( .A(round_reg[1442]), .B(n2210), .Z(n1189) );
  ANDN U3508 ( .B(n3309), .A(n3206), .Z(n3308) );
  XOR U3509 ( .A(n3310), .B(n1233), .Z(out[287]) );
  XOR U3510 ( .A(round_reg[1441]), .B(n2218), .Z(n1233) );
  ANDN U3511 ( .B(n3311), .A(n3218), .Z(n3310) );
  XOR U3512 ( .A(n3312), .B(n1278), .Z(out[286]) );
  IV U3513 ( .A(n3251), .Z(n1278) );
  XNOR U3514 ( .A(round_reg[1440]), .B(n2222), .Z(n3251) );
  ANDN U3515 ( .B(n3313), .A(n3250), .Z(n3312) );
  XOR U3516 ( .A(n3314), .B(n1322), .Z(out[285]) );
  IV U3517 ( .A(n3282), .Z(n1322) );
  XNOR U3518 ( .A(round_reg[1439]), .B(n2226), .Z(n3282) );
  ANDN U3519 ( .B(n3315), .A(n3281), .Z(n3314) );
  XOR U3520 ( .A(n3316), .B(n1366), .Z(out[284]) );
  IV U3521 ( .A(n3305), .Z(n1366) );
  XNOR U3522 ( .A(round_reg[1438]), .B(n2230), .Z(n3305) );
  ANDN U3523 ( .B(n3317), .A(n3304), .Z(n3316) );
  XOR U3524 ( .A(n3318), .B(n1410), .Z(out[283]) );
  IV U3525 ( .A(n3319), .Z(n1410) );
  XOR U3526 ( .A(n3322), .B(n1454), .Z(out[282]) );
  IV U3527 ( .A(n3323), .Z(n1454) );
  XOR U3528 ( .A(n3326), .B(n1502), .Z(out[281]) );
  IV U3529 ( .A(n3327), .Z(n1502) );
  ANDN U3530 ( .B(n3328), .A(n3329), .Z(n3326) );
  XOR U3531 ( .A(n3330), .B(n1536), .Z(out[280]) );
  IV U3532 ( .A(n3331), .Z(n1536) );
  ANDN U3533 ( .B(n3332), .A(n3333), .Z(n3330) );
  XNOR U3534 ( .A(n3334), .B(n1409), .Z(out[27]) );
  AND U3535 ( .A(n3321), .B(n3319), .Z(n3334) );
  XNOR U3536 ( .A(round_reg[1437]), .B(n2234), .Z(n3319) );
  XOR U3537 ( .A(n3335), .B(n1566), .Z(out[279]) );
  IV U3538 ( .A(n3336), .Z(n1566) );
  ANDN U3539 ( .B(n3337), .A(n3338), .Z(n3335) );
  XOR U3540 ( .A(n3339), .B(n1591), .Z(out[278]) );
  IV U3541 ( .A(n3340), .Z(n1591) );
  ANDN U3542 ( .B(n3341), .A(n3342), .Z(n3339) );
  XOR U3543 ( .A(n3343), .B(n1624), .Z(out[277]) );
  IV U3544 ( .A(n3344), .Z(n1624) );
  ANDN U3545 ( .B(n3345), .A(n3346), .Z(n3343) );
  XOR U3546 ( .A(n3347), .B(n1658), .Z(out[276]) );
  IV U3547 ( .A(n3348), .Z(n1658) );
  AND U3548 ( .A(n3349), .B(n3350), .Z(n3347) );
  XOR U3549 ( .A(n3351), .B(n1692), .Z(out[275]) );
  IV U3550 ( .A(n3352), .Z(n1692) );
  AND U3551 ( .A(n3353), .B(n3354), .Z(n3351) );
  XOR U3552 ( .A(n3355), .B(n1720), .Z(out[274]) );
  IV U3553 ( .A(n3356), .Z(n1720) );
  AND U3554 ( .A(n3357), .B(n3358), .Z(n3355) );
  XOR U3555 ( .A(n3359), .B(n1754), .Z(out[273]) );
  IV U3556 ( .A(n3360), .Z(n1754) );
  AND U3557 ( .A(n3361), .B(n3362), .Z(n3359) );
  XOR U3558 ( .A(n3363), .B(n1788), .Z(out[272]) );
  IV U3559 ( .A(n3364), .Z(n1788) );
  AND U3560 ( .A(n3365), .B(n3366), .Z(n3363) );
  XOR U3561 ( .A(n3367), .B(n1826), .Z(out[271]) );
  IV U3562 ( .A(n3368), .Z(n1826) );
  AND U3563 ( .A(n3369), .B(n3370), .Z(n3367) );
  XOR U3564 ( .A(n3371), .B(n1860), .Z(out[270]) );
  IV U3565 ( .A(n3372), .Z(n1860) );
  AND U3566 ( .A(n3373), .B(n3374), .Z(n3371) );
  XNOR U3567 ( .A(n3375), .B(n1453), .Z(out[26]) );
  AND U3568 ( .A(n3325), .B(n3323), .Z(n3375) );
  XNOR U3569 ( .A(round_reg[1436]), .B(n2238), .Z(n3323) );
  XOR U3570 ( .A(n3376), .B(n1893), .Z(out[269]) );
  IV U3571 ( .A(n3377), .Z(n1893) );
  AND U3572 ( .A(n3378), .B(n3379), .Z(n3376) );
  XOR U3573 ( .A(n3380), .B(n1927), .Z(out[268]) );
  IV U3574 ( .A(n3381), .Z(n1927) );
  AND U3575 ( .A(n3382), .B(n3383), .Z(n3380) );
  XOR U3576 ( .A(n3384), .B(n1958), .Z(out[267]) );
  IV U3577 ( .A(n3385), .Z(n1958) );
  AND U3578 ( .A(n3386), .B(n3387), .Z(n3384) );
  XOR U3579 ( .A(n3388), .B(n1990), .Z(out[266]) );
  IV U3580 ( .A(n3389), .Z(n1990) );
  AND U3581 ( .A(n3390), .B(n3391), .Z(n3388) );
  XOR U3582 ( .A(n3392), .B(n1054), .Z(out[265]) );
  XOR U3583 ( .A(round_reg[1419]), .B(n2314), .Z(n1054) );
  NOR U3584 ( .A(n3393), .B(n1053), .Z(n3392) );
  XOR U3585 ( .A(n3394), .B(n1498), .Z(out[264]) );
  XOR U3586 ( .A(round_reg[1418]), .B(n2318), .Z(n1498) );
  AND U3587 ( .A(n3395), .B(n1497), .Z(n3394) );
  IV U3588 ( .A(n3396), .Z(n1497) );
  XOR U3589 ( .A(n3397), .B(n1822), .Z(out[263]) );
  XOR U3590 ( .A(round_reg[1417]), .B(n2322), .Z(n1822) );
  AND U3591 ( .A(n3398), .B(n1821), .Z(n3397) );
  IV U3592 ( .A(n3399), .Z(n1821) );
  XOR U3593 ( .A(n3400), .B(n2092), .Z(out[262]) );
  IV U3594 ( .A(n2123), .Z(n2092) );
  XNOR U3595 ( .A(round_reg[1416]), .B(n2326), .Z(n2123) );
  XOR U3596 ( .A(n3402), .B(n2127), .Z(out[261]) );
  IV U3597 ( .A(n2566), .Z(n2127) );
  XNOR U3598 ( .A(round_reg[1415]), .B(n2330), .Z(n2566) );
  XOR U3599 ( .A(n3404), .B(n2171), .Z(out[260]) );
  IV U3600 ( .A(n2882), .Z(n2171) );
  XNOR U3601 ( .A(round_reg[1414]), .B(n2334), .Z(n2882) );
  XNOR U3602 ( .A(n3406), .B(n1501), .Z(out[25]) );
  AND U3603 ( .A(n3329), .B(n3327), .Z(n3406) );
  XNOR U3604 ( .A(round_reg[1435]), .B(n2242), .Z(n3327) );
  XOR U3605 ( .A(n3407), .B(n2215), .Z(out[259]) );
  IV U3606 ( .A(n3106), .Z(n2215) );
  XNOR U3607 ( .A(round_reg[1413]), .B(n2338), .Z(n3106) );
  XOR U3608 ( .A(n3409), .B(n2259), .Z(out[258]) );
  IV U3609 ( .A(n3279), .Z(n2259) );
  XNOR U3610 ( .A(round_reg[1412]), .B(n2342), .Z(n3279) );
  ANDN U3611 ( .B(n3410), .A(n3278), .Z(n3409) );
  XOR U3612 ( .A(n3411), .B(n2303), .Z(out[257]) );
  IV U3613 ( .A(n3412), .Z(n2303) );
  XOR U3614 ( .A(n3415), .B(n2346), .Z(out[256]) );
  IV U3615 ( .A(n3416), .Z(n2346) );
  XOR U3616 ( .A(n3419), .B(n2391), .Z(out[255]) );
  IV U3617 ( .A(n3221), .Z(n2391) );
  XNOR U3618 ( .A(round_reg[1032]), .B(n1814), .Z(n3221) );
  NOR U3619 ( .A(n3420), .B(n3220), .Z(n3419) );
  XOR U3620 ( .A(n3421), .B(n2435), .Z(out[254]) );
  IV U3621 ( .A(n3224), .Z(n2435) );
  XNOR U3622 ( .A(round_reg[1031]), .B(n1817), .Z(n3224) );
  NOR U3623 ( .A(n3422), .B(n3223), .Z(n3421) );
  XOR U3624 ( .A(n3423), .B(n2479), .Z(out[253]) );
  IV U3625 ( .A(n3227), .Z(n2479) );
  XNOR U3626 ( .A(round_reg[1030]), .B(n1828), .Z(n3227) );
  NOR U3627 ( .A(n3424), .B(n3226), .Z(n3423) );
  XOR U3628 ( .A(n3425), .B(n2523), .Z(out[252]) );
  IV U3629 ( .A(n3230), .Z(n2523) );
  XNOR U3630 ( .A(round_reg[1029]), .B(n1831), .Z(n3230) );
  NOR U3631 ( .A(n3426), .B(n3229), .Z(n3425) );
  XOR U3632 ( .A(n3427), .B(n2570), .Z(out[251]) );
  IV U3633 ( .A(n3233), .Z(n2570) );
  XNOR U3634 ( .A(round_reg[1028]), .B(n1834), .Z(n3233) );
  NOR U3635 ( .A(n3428), .B(n3232), .Z(n3427) );
  XOR U3636 ( .A(n3429), .B(n2614), .Z(out[250]) );
  IV U3637 ( .A(n3236), .Z(n2614) );
  XNOR U3638 ( .A(round_reg[1027]), .B(n1837), .Z(n3236) );
  ANDN U3639 ( .B(n3430), .A(n3235), .Z(n3429) );
  XNOR U3640 ( .A(n3431), .B(n1535), .Z(out[24]) );
  AND U3641 ( .A(n3333), .B(n3331), .Z(n3431) );
  XNOR U3642 ( .A(round_reg[1434]), .B(n2246), .Z(n3331) );
  XOR U3643 ( .A(n3432), .B(n2658), .Z(out[249]) );
  IV U3644 ( .A(n3239), .Z(n2658) );
  XNOR U3645 ( .A(round_reg[1026]), .B(n1840), .Z(n3239) );
  ANDN U3646 ( .B(n3433), .A(n3238), .Z(n3432) );
  XOR U3647 ( .A(n3434), .B(n2690), .Z(out[248]) );
  IV U3648 ( .A(n3242), .Z(n2690) );
  XNOR U3649 ( .A(round_reg[1025]), .B(n1843), .Z(n3242) );
  ANDN U3650 ( .B(n3435), .A(n3241), .Z(n3434) );
  XOR U3651 ( .A(n3436), .B(n2722), .Z(out[247]) );
  IV U3652 ( .A(n3245), .Z(n2722) );
  XNOR U3653 ( .A(round_reg[1024]), .B(n1846), .Z(n3245) );
  ANDN U3654 ( .B(n3437), .A(n3244), .Z(n3436) );
  XOR U3655 ( .A(n3438), .B(n2751), .Z(out[246]) );
  IV U3656 ( .A(n3248), .Z(n2751) );
  XNOR U3657 ( .A(round_reg[1087]), .B(n1849), .Z(n3248) );
  ANDN U3658 ( .B(n3439), .A(n3247), .Z(n3438) );
  XOR U3659 ( .A(n3440), .B(n2784), .Z(out[245]) );
  IV U3660 ( .A(n3254), .Z(n2784) );
  XNOR U3661 ( .A(round_reg[1086]), .B(n1852), .Z(n3254) );
  ANDN U3662 ( .B(n3441), .A(n3253), .Z(n3440) );
  XOR U3663 ( .A(n3442), .B(n2808), .Z(out[244]) );
  IV U3664 ( .A(n3257), .Z(n2808) );
  XNOR U3665 ( .A(round_reg[1085]), .B(n1855), .Z(n3257) );
  ANDN U3666 ( .B(n3443), .A(n3256), .Z(n3442) );
  XOR U3667 ( .A(n3444), .B(n2833), .Z(out[243]) );
  IV U3668 ( .A(n3260), .Z(n2833) );
  XNOR U3669 ( .A(round_reg[1084]), .B(n1862), .Z(n3260) );
  ANDN U3670 ( .B(n3445), .A(n3259), .Z(n3444) );
  XOR U3671 ( .A(n3446), .B(n2859), .Z(out[242]) );
  IV U3672 ( .A(n3263), .Z(n2859) );
  XNOR U3673 ( .A(round_reg[1083]), .B(n1865), .Z(n3263) );
  ANDN U3674 ( .B(n3447), .A(n3262), .Z(n3446) );
  XOR U3675 ( .A(n3448), .B(n2886), .Z(out[241]) );
  IV U3676 ( .A(n3266), .Z(n2886) );
  XNOR U3677 ( .A(round_reg[1082]), .B(n1868), .Z(n3266) );
  ANDN U3678 ( .B(n3449), .A(n3265), .Z(n3448) );
  XOR U3679 ( .A(n3450), .B(n2909), .Z(out[240]) );
  XOR U3680 ( .A(round_reg[1081]), .B(n1871), .Z(n2909) );
  ANDN U3681 ( .B(n3451), .A(n3268), .Z(n3450) );
  XNOR U3682 ( .A(n3452), .B(n1565), .Z(out[23]) );
  AND U3683 ( .A(n3338), .B(n3336), .Z(n3452) );
  XNOR U3684 ( .A(round_reg[1433]), .B(n2250), .Z(n3336) );
  XOR U3685 ( .A(n3453), .B(n2933), .Z(out[239]) );
  XOR U3686 ( .A(round_reg[1080]), .B(n1874), .Z(n2933) );
  AND U3687 ( .A(n3454), .B(n3455), .Z(n3453) );
  XOR U3688 ( .A(n3456), .B(n2957), .Z(out[238]) );
  XOR U3689 ( .A(round_reg[1079]), .B(n1877), .Z(n2957) );
  ANDN U3690 ( .B(n3457), .A(n3272), .Z(n3456) );
  XOR U3691 ( .A(n3458), .B(n2981), .Z(out[237]) );
  XOR U3692 ( .A(round_reg[1078]), .B(n1880), .Z(n2981) );
  ANDN U3693 ( .B(n3459), .A(n3274), .Z(n3458) );
  XOR U3694 ( .A(n3460), .B(n3008), .Z(out[236]) );
  XOR U3695 ( .A(round_reg[1077]), .B(n1883), .Z(n3008) );
  ANDN U3696 ( .B(n3461), .A(n3276), .Z(n3460) );
  XOR U3697 ( .A(n3462), .B(n3024), .Z(out[235]) );
  XOR U3698 ( .A(round_reg[1076]), .B(n1886), .Z(n3024) );
  ANDN U3699 ( .B(n3463), .A(n3284), .Z(n3462) );
  XOR U3700 ( .A(n3464), .B(n3043), .Z(out[234]) );
  XOR U3701 ( .A(round_reg[1075]), .B(n1889), .Z(n3043) );
  ANDN U3702 ( .B(n3465), .A(n3286), .Z(n3464) );
  XOR U3703 ( .A(n3466), .B(n3066), .Z(out[233]) );
  XOR U3704 ( .A(round_reg[1074]), .B(n1896), .Z(n3066) );
  ANDN U3705 ( .B(n3467), .A(n3288), .Z(n3466) );
  XOR U3706 ( .A(n3468), .B(n3084), .Z(out[232]) );
  XOR U3707 ( .A(round_reg[1073]), .B(n1899), .Z(n3084) );
  ANDN U3708 ( .B(n3469), .A(n3290), .Z(n3468) );
  XOR U3709 ( .A(n3470), .B(n3109), .Z(out[231]) );
  XOR U3710 ( .A(round_reg[1072]), .B(n1902), .Z(n3109) );
  ANDN U3711 ( .B(n3471), .A(n3292), .Z(n3470) );
  XOR U3712 ( .A(n3472), .B(n3129), .Z(out[230]) );
  XOR U3713 ( .A(round_reg[1071]), .B(n1905), .Z(n3129) );
  ANDN U3714 ( .B(n3473), .A(n3294), .Z(n3472) );
  XNOR U3715 ( .A(n3474), .B(n1590), .Z(out[22]) );
  AND U3716 ( .A(n3342), .B(n3340), .Z(n3474) );
  XNOR U3717 ( .A(round_reg[1432]), .B(n2254), .Z(n3340) );
  XOR U3718 ( .A(n3475), .B(n3143), .Z(out[229]) );
  XOR U3719 ( .A(round_reg[1070]), .B(n1908), .Z(n3143) );
  ANDN U3720 ( .B(n3476), .A(n3296), .Z(n3475) );
  XOR U3721 ( .A(n3477), .B(n3157), .Z(out[228]) );
  XOR U3722 ( .A(round_reg[1069]), .B(n1911), .Z(n3157) );
  ANDN U3723 ( .B(n3478), .A(n3298), .Z(n3477) );
  XOR U3724 ( .A(n3479), .B(n3170), .Z(out[227]) );
  XNOR U3725 ( .A(round_reg[1068]), .B(n1914), .Z(n3170) );
  ANDN U3726 ( .B(n1056), .A(n3300), .Z(n3479) );
  XOR U3727 ( .A(n3480), .B(n3182), .Z(out[226]) );
  XNOR U3728 ( .A(round_reg[1067]), .B(n1917), .Z(n3182) );
  ANDN U3729 ( .B(n1100), .A(n3302), .Z(n3480) );
  XOR U3730 ( .A(n3481), .B(n3194), .Z(out[225]) );
  XNOR U3731 ( .A(round_reg[1066]), .B(n1920), .Z(n3194) );
  ANDN U3732 ( .B(n1144), .A(n3307), .Z(n3481) );
  XOR U3733 ( .A(n3482), .B(n3206), .Z(out[224]) );
  XNOR U3734 ( .A(round_reg[1065]), .B(n1923), .Z(n3206) );
  NOR U3735 ( .A(n1188), .B(n3309), .Z(n3482) );
  XOR U3736 ( .A(n3483), .B(n3218), .Z(out[223]) );
  XNOR U3737 ( .A(round_reg[1064]), .B(n1930), .Z(n3218) );
  XOR U3738 ( .A(n3484), .B(n3250), .Z(out[222]) );
  XNOR U3739 ( .A(round_reg[1063]), .B(n1933), .Z(n3250) );
  XOR U3740 ( .A(n3485), .B(n3281), .Z(out[221]) );
  XNOR U3741 ( .A(round_reg[1062]), .B(n1712), .Z(n3281) );
  XOR U3742 ( .A(n3486), .B(n3304), .Z(out[220]) );
  XNOR U3743 ( .A(round_reg[1061]), .B(n1715), .Z(n3304) );
  XNOR U3744 ( .A(n3487), .B(n1623), .Z(out[21]) );
  AND U3745 ( .A(n3346), .B(n3344), .Z(n3487) );
  XNOR U3746 ( .A(round_reg[1431]), .B(n2262), .Z(n3344) );
  XOR U3747 ( .A(n3488), .B(n3321), .Z(out[219]) );
  XNOR U3748 ( .A(round_reg[1060]), .B(n1722), .Z(n3321) );
  NOR U3749 ( .A(n3320), .B(n1408), .Z(n3488) );
  XOR U3750 ( .A(n3489), .B(n3325), .Z(out[218]) );
  XNOR U3751 ( .A(round_reg[1059]), .B(n1725), .Z(n3325) );
  NOR U3752 ( .A(n3324), .B(n1452), .Z(n3489) );
  XOR U3753 ( .A(n3490), .B(n3329), .Z(out[217]) );
  XOR U3754 ( .A(round_reg[1058]), .B(n1728), .Z(n3329) );
  NOR U3755 ( .A(n3328), .B(n1500), .Z(n3490) );
  XOR U3756 ( .A(n3491), .B(n3333), .Z(out[216]) );
  XOR U3757 ( .A(round_reg[1057]), .B(n1731), .Z(n3333) );
  NOR U3758 ( .A(n3332), .B(n1534), .Z(n3491) );
  XOR U3759 ( .A(n3492), .B(n3338), .Z(out[215]) );
  XOR U3760 ( .A(round_reg[1056]), .B(n1734), .Z(n3338) );
  NOR U3761 ( .A(n3337), .B(n1564), .Z(n3492) );
  XOR U3762 ( .A(n3493), .B(n3342), .Z(out[214]) );
  XOR U3763 ( .A(round_reg[1055]), .B(n1737), .Z(n3342) );
  NOR U3764 ( .A(n3341), .B(n1589), .Z(n3493) );
  XOR U3765 ( .A(n3494), .B(n3346), .Z(out[213]) );
  XOR U3766 ( .A(round_reg[1054]), .B(n1740), .Z(n3346) );
  NOR U3767 ( .A(n3345), .B(n1622), .Z(n3494) );
  XNOR U3768 ( .A(n3495), .B(n3350), .Z(out[212]) );
  NOR U3769 ( .A(n3349), .B(n1656), .Z(n3495) );
  XNOR U3770 ( .A(n3496), .B(n3354), .Z(out[211]) );
  NOR U3771 ( .A(n3353), .B(n1690), .Z(n3496) );
  XNOR U3772 ( .A(n3497), .B(n3357), .Z(out[210]) );
  XNOR U3773 ( .A(n3498), .B(n1657), .Z(out[20]) );
  ANDN U3774 ( .B(n3348), .A(n3350), .Z(n3498) );
  XNOR U3775 ( .A(round_reg[1053]), .B(n1743), .Z(n3350) );
  XNOR U3776 ( .A(round_reg[1430]), .B(n2266), .Z(n3348) );
  XNOR U3777 ( .A(n3499), .B(n3361), .Z(out[209]) );
  XNOR U3778 ( .A(n3500), .B(n3365), .Z(out[208]) );
  ANDN U3779 ( .B(n3501), .A(n1786), .Z(n3500) );
  XNOR U3780 ( .A(n3502), .B(n3369), .Z(out[207]) );
  ANDN U3781 ( .B(n3503), .A(n1824), .Z(n3502) );
  XNOR U3782 ( .A(n3504), .B(n3373), .Z(out[206]) );
  ANDN U3783 ( .B(n3505), .A(n1858), .Z(n3504) );
  XNOR U3784 ( .A(n3506), .B(n3378), .Z(out[205]) );
  ANDN U3785 ( .B(n3507), .A(n1892), .Z(n3506) );
  XNOR U3786 ( .A(n3508), .B(n3382), .Z(out[204]) );
  ANDN U3787 ( .B(n3509), .A(n1926), .Z(n3508) );
  XNOR U3788 ( .A(n3510), .B(n3386), .Z(out[203]) );
  ANDN U3789 ( .B(n3511), .A(n1957), .Z(n3510) );
  XNOR U3790 ( .A(n3512), .B(n3390), .Z(out[202]) );
  ANDN U3791 ( .B(n3513), .A(n1989), .Z(n3512) );
  XOR U3792 ( .A(n3514), .B(n1053), .Z(out[201]) );
  XOR U3793 ( .A(round_reg[1042]), .B(n1780), .Z(n1053) );
  ANDN U3794 ( .B(n3393), .A(n2017), .Z(n3514) );
  IV U3795 ( .A(n3515), .Z(n3393) );
  XOR U3796 ( .A(n3516), .B(n3396), .Z(out[200]) );
  XOR U3797 ( .A(round_reg[1041]), .B(n1783), .Z(n3396) );
  XNOR U3798 ( .A(n3517), .B(n2302), .Z(out[1]) );
  AND U3799 ( .A(n3414), .B(n3412), .Z(n3517) );
  XNOR U3800 ( .A(round_reg[1411]), .B(n2350), .Z(n3412) );
  XNOR U3801 ( .A(n3518), .B(n1691), .Z(out[19]) );
  ANDN U3802 ( .B(n3352), .A(n3354), .Z(n3518) );
  XNOR U3803 ( .A(round_reg[1052]), .B(n1746), .Z(n3354) );
  XNOR U3804 ( .A(round_reg[1429]), .B(n2270), .Z(n3352) );
  XOR U3805 ( .A(n3519), .B(n3399), .Z(out[199]) );
  XOR U3806 ( .A(round_reg[1040]), .B(n1790), .Z(n3399) );
  XOR U3807 ( .A(n3520), .B(n2122), .Z(out[198]) );
  XOR U3808 ( .A(round_reg[1039]), .B(n1793), .Z(n2122) );
  XOR U3809 ( .A(n3521), .B(n2565), .Z(out[197]) );
  XOR U3810 ( .A(round_reg[1038]), .B(n1796), .Z(n2565) );
  XOR U3811 ( .A(n3522), .B(n2881), .Z(out[196]) );
  XOR U3812 ( .A(round_reg[1037]), .B(n1799), .Z(n2881) );
  XOR U3813 ( .A(n3523), .B(n3105), .Z(out[195]) );
  XOR U3814 ( .A(round_reg[1036]), .B(n1802), .Z(n3105) );
  NOR U3815 ( .A(n3408), .B(n2213), .Z(n3523) );
  XOR U3816 ( .A(n3524), .B(n3278), .Z(out[194]) );
  XOR U3817 ( .A(round_reg[1035]), .B(n1805), .Z(n3278) );
  ANDN U3818 ( .B(n3525), .A(n2257), .Z(n3524) );
  XOR U3819 ( .A(n3526), .B(n3414), .Z(out[193]) );
  XOR U3820 ( .A(round_reg[1034]), .B(n1808), .Z(n3414) );
  NOR U3821 ( .A(n3413), .B(n2301), .Z(n3526) );
  XOR U3822 ( .A(n3527), .B(n3418), .Z(out[192]) );
  NOR U3823 ( .A(n3417), .B(n2345), .Z(n3527) );
  XOR U3824 ( .A(n3528), .B(n3220), .Z(out[191]) );
  XOR U3825 ( .A(round_reg[664]), .B(n2028), .Z(n3220) );
  ANDN U3826 ( .B(n3420), .A(n2389), .Z(n3528) );
  IV U3827 ( .A(n3529), .Z(n3420) );
  XOR U3828 ( .A(n3530), .B(n3223), .Z(out[190]) );
  XOR U3829 ( .A(round_reg[663]), .B(n2031), .Z(n3223) );
  ANDN U3830 ( .B(n3422), .A(n2433), .Z(n3530) );
  IV U3831 ( .A(n3531), .Z(n3422) );
  XNOR U3832 ( .A(n3532), .B(n1719), .Z(out[18]) );
  ANDN U3833 ( .B(n3356), .A(n3357), .Z(n3532) );
  XNOR U3834 ( .A(round_reg[1051]), .B(n1749), .Z(n3357) );
  XNOR U3835 ( .A(round_reg[1428]), .B(n2274), .Z(n3356) );
  XOR U3836 ( .A(n3533), .B(n3226), .Z(out[189]) );
  XOR U3837 ( .A(round_reg[662]), .B(n2034), .Z(n3226) );
  ANDN U3838 ( .B(n3424), .A(n2477), .Z(n3533) );
  IV U3839 ( .A(n3534), .Z(n3424) );
  XOR U3840 ( .A(n3535), .B(n3229), .Z(out[188]) );
  XOR U3841 ( .A(round_reg[661]), .B(n2037), .Z(n3229) );
  ANDN U3842 ( .B(n3426), .A(n2521), .Z(n3535) );
  IV U3843 ( .A(n3536), .Z(n3426) );
  XOR U3844 ( .A(n3537), .B(n3232), .Z(out[187]) );
  XOR U3845 ( .A(round_reg[660]), .B(n2040), .Z(n3232) );
  ANDN U3846 ( .B(n3428), .A(n2568), .Z(n3537) );
  IV U3847 ( .A(n3538), .Z(n3428) );
  XOR U3848 ( .A(n3539), .B(n3235), .Z(out[186]) );
  XOR U3849 ( .A(round_reg[659]), .B(n2042), .Z(n3235) );
  ANDN U3850 ( .B(n3540), .A(n2612), .Z(n3539) );
  XOR U3851 ( .A(n3541), .B(n3238), .Z(out[185]) );
  XOR U3852 ( .A(round_reg[658]), .B(n2044), .Z(n3238) );
  XOR U3853 ( .A(n3542), .B(n3241), .Z(out[184]) );
  XOR U3854 ( .A(round_reg[657]), .B(n2048), .Z(n3241) );
  XOR U3855 ( .A(n3543), .B(n3244), .Z(out[183]) );
  XOR U3856 ( .A(round_reg[656]), .B(n2050), .Z(n3244) );
  XOR U3857 ( .A(n3544), .B(n3247), .Z(out[182]) );
  XOR U3858 ( .A(round_reg[655]), .B(n2052), .Z(n3247) );
  XOR U3859 ( .A(n3545), .B(n3253), .Z(out[181]) );
  XOR U3860 ( .A(round_reg[654]), .B(n2054), .Z(n3253) );
  XOR U3861 ( .A(n3546), .B(n3256), .Z(out[180]) );
  XOR U3862 ( .A(round_reg[653]), .B(n2056), .Z(n3256) );
  XNOR U3863 ( .A(n3547), .B(n1753), .Z(out[17]) );
  ANDN U3864 ( .B(n3360), .A(n3361), .Z(n3547) );
  XOR U3865 ( .A(round_reg[1050]), .B(n1756), .Z(n3361) );
  XNOR U3866 ( .A(round_reg[1427]), .B(n2278), .Z(n3360) );
  XOR U3867 ( .A(n3548), .B(n3259), .Z(out[179]) );
  XOR U3868 ( .A(round_reg[652]), .B(n2058), .Z(n3259) );
  ANDN U3869 ( .B(n3549), .A(n2831), .Z(n3548) );
  XOR U3870 ( .A(n3550), .B(n3262), .Z(out[178]) );
  XOR U3871 ( .A(round_reg[651]), .B(n2060), .Z(n3262) );
  ANDN U3872 ( .B(n3551), .A(n2857), .Z(n3550) );
  XOR U3873 ( .A(n3552), .B(n3265), .Z(out[177]) );
  XOR U3874 ( .A(round_reg[650]), .B(n2062), .Z(n3265) );
  ANDN U3875 ( .B(n3553), .A(n2884), .Z(n3552) );
  XOR U3876 ( .A(n3554), .B(n3268), .Z(out[176]) );
  XOR U3877 ( .A(round_reg[649]), .B(n2064), .Z(n3268) );
  ANDN U3878 ( .B(n3555), .A(n2908), .Z(n3554) );
  XOR U3879 ( .A(n3556), .B(n3270), .Z(out[175]) );
  IV U3880 ( .A(n3455), .Z(n3270) );
  XNOR U3881 ( .A(round_reg[648]), .B(n2066), .Z(n3455) );
  NOR U3882 ( .A(n3454), .B(n2932), .Z(n3556) );
  XOR U3883 ( .A(n3557), .B(n3272), .Z(out[174]) );
  XOR U3884 ( .A(round_reg[647]), .B(n2070), .Z(n3272) );
  ANDN U3885 ( .B(n3558), .A(n2956), .Z(n3557) );
  XOR U3886 ( .A(n3559), .B(n3274), .Z(out[173]) );
  XOR U3887 ( .A(round_reg[646]), .B(n2072), .Z(n3274) );
  ANDN U3888 ( .B(n3560), .A(n2980), .Z(n3559) );
  XOR U3889 ( .A(n3561), .B(n3276), .Z(out[172]) );
  XOR U3890 ( .A(round_reg[645]), .B(n2074), .Z(n3276) );
  ANDN U3891 ( .B(n3562), .A(n3007), .Z(n3561) );
  XOR U3892 ( .A(n3563), .B(n3284), .Z(out[171]) );
  XOR U3893 ( .A(round_reg[644]), .B(n2076), .Z(n3284) );
  ANDN U3894 ( .B(n3564), .A(n3023), .Z(n3563) );
  XOR U3895 ( .A(n3565), .B(n3286), .Z(out[170]) );
  XOR U3896 ( .A(round_reg[643]), .B(n2078), .Z(n3286) );
  ANDN U3897 ( .B(n3566), .A(n3042), .Z(n3565) );
  XNOR U3898 ( .A(n3567), .B(n1787), .Z(out[16]) );
  ANDN U3899 ( .B(n3364), .A(n3365), .Z(n3567) );
  XOR U3900 ( .A(round_reg[1049]), .B(n1759), .Z(n3365) );
  XNOR U3901 ( .A(round_reg[1426]), .B(n2282), .Z(n3364) );
  XOR U3902 ( .A(n3568), .B(n3288), .Z(out[169]) );
  XOR U3903 ( .A(round_reg[642]), .B(n2080), .Z(n3288) );
  ANDN U3904 ( .B(n3569), .A(n3065), .Z(n3568) );
  XOR U3905 ( .A(n3570), .B(n3290), .Z(out[168]) );
  XOR U3906 ( .A(round_reg[641]), .B(n2082), .Z(n3290) );
  ANDN U3907 ( .B(n3571), .A(n3083), .Z(n3570) );
  XOR U3908 ( .A(n3572), .B(n3292), .Z(out[167]) );
  XOR U3909 ( .A(round_reg[640]), .B(n2084), .Z(n3292) );
  ANDN U3910 ( .B(n3573), .A(n3108), .Z(n3572) );
  XOR U3911 ( .A(n3574), .B(n3294), .Z(out[166]) );
  XNOR U3912 ( .A(round_reg[703]), .B(n2086), .Z(n3294) );
  ANDN U3913 ( .B(n3575), .A(n3128), .Z(n3574) );
  XOR U3914 ( .A(n3576), .B(n3296), .Z(out[165]) );
  XOR U3915 ( .A(round_reg[702]), .B(n2088), .Z(n3296) );
  ANDN U3916 ( .B(n3577), .A(n3142), .Z(n3576) );
  XOR U3917 ( .A(n3578), .B(n3298), .Z(out[164]) );
  XOR U3918 ( .A(round_reg[701]), .B(n2094), .Z(n3298) );
  ANDN U3919 ( .B(n3579), .A(n3156), .Z(n3578) );
  XOR U3920 ( .A(n3580), .B(n3300), .Z(out[163]) );
  XOR U3921 ( .A(round_reg[700]), .B(n2096), .Z(n3300) );
  ANDN U3922 ( .B(n1058), .A(n1056), .Z(n3580) );
  XOR U3923 ( .A(round_reg[634]), .B(n2333), .Z(n1056) );
  XOR U3924 ( .A(round_reg[225]), .B(n2239), .Z(n1058) );
  XOR U3925 ( .A(n3581), .B(n3302), .Z(out[162]) );
  XOR U3926 ( .A(round_reg[699]), .B(n2098), .Z(n3302) );
  ANDN U3927 ( .B(n1102), .A(n1100), .Z(n3581) );
  XOR U3928 ( .A(round_reg[633]), .B(n2337), .Z(n1100) );
  XNOR U3929 ( .A(round_reg[224]), .B(n2243), .Z(n1102) );
  XOR U3930 ( .A(n3582), .B(n3307), .Z(out[161]) );
  XOR U3931 ( .A(round_reg[698]), .B(n2100), .Z(n3307) );
  NOR U3932 ( .A(n1146), .B(n1144), .Z(n3582) );
  XOR U3933 ( .A(round_reg[632]), .B(n2341), .Z(n1144) );
  XOR U3934 ( .A(round_reg[223]), .B(n2247), .Z(n1146) );
  XOR U3935 ( .A(n3583), .B(n3309), .Z(out[160]) );
  XOR U3936 ( .A(round_reg[697]), .B(n2102), .Z(n3309) );
  ANDN U3937 ( .B(n1188), .A(n1190), .Z(n3583) );
  XOR U3938 ( .A(round_reg[222]), .B(n2251), .Z(n1190) );
  XNOR U3939 ( .A(round_reg[631]), .B(n2349), .Z(n1188) );
  XNOR U3940 ( .A(n3584), .B(n1825), .Z(out[15]) );
  ANDN U3941 ( .B(n3368), .A(n3369), .Z(n3584) );
  XOR U3942 ( .A(round_reg[1048]), .B(n1762), .Z(n3369) );
  XNOR U3943 ( .A(round_reg[1425]), .B(n2286), .Z(n3368) );
  XOR U3944 ( .A(n3585), .B(n3311), .Z(out[159]) );
  XOR U3945 ( .A(round_reg[696]), .B(n2104), .Z(n3311) );
  ANDN U3946 ( .B(n1232), .A(n1234), .Z(n3585) );
  XOR U3947 ( .A(round_reg[221]), .B(n2255), .Z(n1234) );
  XNOR U3948 ( .A(round_reg[630]), .B(n2353), .Z(n1232) );
  XOR U3949 ( .A(n3586), .B(n3587), .Z(out[1599]) );
  XOR U3950 ( .A(n3588), .B(n3589), .Z(n3587) );
  NAND U3951 ( .A(n3590), .B(n3591), .Z(n3589) );
  AND U3952 ( .A(n3592), .B(n3593), .Z(n3591) );
  NOR U3953 ( .A(rc_i[2]), .B(rc_i[3]), .Z(n3593) );
  NOR U3954 ( .A(rc_i[17]), .B(rc_i[19]), .Z(n3592) );
  AND U3955 ( .A(n3594), .B(n3595), .Z(n3590) );
  NOR U3956 ( .A(rc_i[16]), .B(n3596), .Z(n3595) );
  ANDN U3957 ( .B(n3597), .A(n3598), .Z(n3594) );
  XOR U3958 ( .A(n3601), .B(n3602), .Z(out[1598]) );
  AND U3959 ( .A(n3603), .B(n3604), .Z(n3601) );
  XOR U3960 ( .A(n3605), .B(n3606), .Z(out[1597]) );
  AND U3961 ( .A(n3607), .B(n3608), .Z(n3605) );
  XOR U3962 ( .A(n3609), .B(n3610), .Z(out[1596]) );
  AND U3963 ( .A(n3611), .B(n3612), .Z(n3609) );
  XOR U3964 ( .A(n3613), .B(n3614), .Z(out[1595]) );
  AND U3965 ( .A(n3615), .B(n3616), .Z(n3613) );
  XOR U3966 ( .A(n3617), .B(n3618), .Z(out[1594]) );
  AND U3967 ( .A(n3619), .B(n3620), .Z(n3617) );
  XOR U3968 ( .A(n3621), .B(n3622), .Z(out[1593]) );
  AND U3969 ( .A(n3623), .B(n3624), .Z(n3621) );
  XOR U3970 ( .A(n3625), .B(n3626), .Z(out[1592]) );
  AND U3971 ( .A(n3627), .B(n3628), .Z(n3625) );
  XOR U3972 ( .A(n3629), .B(n3630), .Z(out[1591]) );
  AND U3973 ( .A(n3631), .B(n3632), .Z(n3629) );
  XOR U3974 ( .A(n3633), .B(n3634), .Z(out[1590]) );
  AND U3975 ( .A(n3635), .B(n3636), .Z(n3633) );
  XOR U3976 ( .A(n3637), .B(n3313), .Z(out[158]) );
  XOR U3977 ( .A(round_reg[695]), .B(n1936), .Z(n3313) );
  ANDN U3978 ( .B(n1276), .A(n1277), .Z(n3637) );
  XOR U3979 ( .A(round_reg[220]), .B(n2263), .Z(n1277) );
  XNOR U3980 ( .A(round_reg[629]), .B(n2357), .Z(n1276) );
  XOR U3981 ( .A(n3638), .B(n3639), .Z(out[1589]) );
  AND U3982 ( .A(n3640), .B(n3641), .Z(n3638) );
  XOR U3983 ( .A(n3642), .B(n3643), .Z(out[1588]) );
  AND U3984 ( .A(n3644), .B(n3645), .Z(n3642) );
  XOR U3985 ( .A(n3646), .B(n3647), .Z(out[1587]) );
  XOR U3986 ( .A(n3650), .B(n3651), .Z(out[1586]) );
  AND U3987 ( .A(n3652), .B(n3653), .Z(n3650) );
  XOR U3988 ( .A(n3654), .B(n3655), .Z(out[1585]) );
  AND U3989 ( .A(n3656), .B(n3657), .Z(n3654) );
  XOR U3990 ( .A(n3658), .B(n3659), .Z(out[1584]) );
  AND U3991 ( .A(n3660), .B(n3661), .Z(n3658) );
  XOR U3992 ( .A(n3662), .B(n3663), .Z(out[1583]) );
  AND U3993 ( .A(n3664), .B(n3665), .Z(n3662) );
  XOR U3994 ( .A(n3666), .B(n3667), .Z(out[1582]) );
  AND U3995 ( .A(n3668), .B(n3669), .Z(n3666) );
  XOR U3996 ( .A(n3670), .B(n3671), .Z(out[1581]) );
  AND U3997 ( .A(n3672), .B(n3673), .Z(n3670) );
  XOR U3998 ( .A(n3674), .B(n3675), .Z(out[1580]) );
  AND U3999 ( .A(n3676), .B(n3677), .Z(n3674) );
  XOR U4000 ( .A(n3678), .B(n3315), .Z(out[157]) );
  XOR U4001 ( .A(round_reg[694]), .B(n1938), .Z(n3315) );
  ANDN U4002 ( .B(n1320), .A(n1321), .Z(n3678) );
  XNOR U4003 ( .A(round_reg[219]), .B(n2267), .Z(n1321) );
  XNOR U4004 ( .A(round_reg[628]), .B(n2361), .Z(n1320) );
  XOR U4005 ( .A(n3679), .B(n3680), .Z(out[1579]) );
  AND U4006 ( .A(n3681), .B(n3682), .Z(n3679) );
  XOR U4007 ( .A(n3683), .B(n3684), .Z(out[1578]) );
  ANDN U4008 ( .B(n3685), .A(n3686), .Z(n3683) );
  XOR U4009 ( .A(n3687), .B(n3688), .Z(out[1577]) );
  AND U4010 ( .A(n3689), .B(n3690), .Z(n3687) );
  XOR U4011 ( .A(n3691), .B(n3692), .Z(out[1576]) );
  XOR U4012 ( .A(n3695), .B(n3696), .Z(out[1575]) );
  XOR U4013 ( .A(n3699), .B(n3700), .Z(out[1574]) );
  AND U4014 ( .A(n3701), .B(n3702), .Z(n3699) );
  XOR U4015 ( .A(n3703), .B(n3704), .Z(out[1573]) );
  AND U4016 ( .A(n3705), .B(n3706), .Z(n3703) );
  XNOR U4017 ( .A(n3707), .B(n3708), .Z(out[1572]) );
  AND U4018 ( .A(n3709), .B(n3710), .Z(n3707) );
  XOR U4019 ( .A(n3711), .B(n3712), .Z(out[1571]) );
  AND U4020 ( .A(n3713), .B(n3714), .Z(n3711) );
  XOR U4021 ( .A(n3715), .B(n3716), .Z(out[1570]) );
  AND U4022 ( .A(n3717), .B(n3718), .Z(n3715) );
  XOR U4023 ( .A(n3719), .B(n3317), .Z(out[156]) );
  XOR U4024 ( .A(round_reg[693]), .B(n1940), .Z(n3317) );
  ANDN U4025 ( .B(n1364), .A(n1365), .Z(n3719) );
  XNOR U4026 ( .A(round_reg[218]), .B(n2271), .Z(n1365) );
  XNOR U4027 ( .A(round_reg[627]), .B(n2365), .Z(n1364) );
  XNOR U4028 ( .A(n3720), .B(n3721), .Z(out[1569]) );
  AND U4029 ( .A(n3722), .B(n3723), .Z(n3720) );
  XNOR U4030 ( .A(n3724), .B(n3725), .Z(out[1568]) );
  AND U4031 ( .A(n3726), .B(n3727), .Z(n3724) );
  XNOR U4032 ( .A(n3728), .B(n3729), .Z(out[1567]) );
  XOR U4033 ( .A(n3730), .B(n3731), .Z(n3729) );
  NAND U4034 ( .A(n3732), .B(n3733), .Z(n3731) );
  AND U4035 ( .A(n3734), .B(n3735), .Z(n3733) );
  ANDN U4036 ( .B(n3736), .A(rc_i[3]), .Z(n3735) );
  NOR U4037 ( .A(rc_i[5]), .B(rc_i[6]), .Z(n3736) );
  NOR U4038 ( .A(rc_i[23]), .B(rc_i[22]), .Z(n3734) );
  AND U4039 ( .A(n3737), .B(n3738), .Z(n3732) );
  AND U4040 ( .A(n3739), .B(n3740), .Z(n3738) );
  NOR U4041 ( .A(rc_i[20]), .B(rc_i[19]), .Z(n3739) );
  NOR U4042 ( .A(rc_i[10]), .B(rc_i[11]), .Z(n3737) );
  AND U4043 ( .A(n3741), .B(n3742), .Z(n3730) );
  XNOR U4044 ( .A(n3743), .B(n3744), .Z(out[1566]) );
  AND U4045 ( .A(n3745), .B(n3746), .Z(n3743) );
  XNOR U4046 ( .A(n3747), .B(n3748), .Z(out[1565]) );
  AND U4047 ( .A(n3749), .B(n3750), .Z(n3747) );
  XNOR U4048 ( .A(n3751), .B(n3752), .Z(out[1564]) );
  AND U4049 ( .A(n3753), .B(n3754), .Z(n3751) );
  XNOR U4050 ( .A(n3755), .B(n3756), .Z(out[1563]) );
  AND U4051 ( .A(n3757), .B(n3758), .Z(n3755) );
  XNOR U4052 ( .A(n3759), .B(n3760), .Z(out[1562]) );
  AND U4053 ( .A(n3761), .B(n3762), .Z(n3759) );
  XOR U4054 ( .A(n3763), .B(n3764), .Z(out[1561]) );
  XOR U4055 ( .A(n3767), .B(n3768), .Z(out[1560]) );
  XOR U4056 ( .A(n3771), .B(n3320), .Z(out[155]) );
  XOR U4057 ( .A(round_reg[692]), .B(n1942), .Z(n3320) );
  ANDN U4058 ( .B(n1408), .A(n1409), .Z(n3771) );
  XNOR U4059 ( .A(round_reg[217]), .B(n2275), .Z(n1409) );
  XNOR U4060 ( .A(round_reg[626]), .B(n2369), .Z(n1408) );
  XOR U4061 ( .A(n3772), .B(n3773), .Z(out[1559]) );
  XOR U4062 ( .A(n3776), .B(n3777), .Z(out[1558]) );
  XNOR U4063 ( .A(n3780), .B(n3781), .Z(out[1557]) );
  XNOR U4064 ( .A(n3784), .B(n3785), .Z(out[1556]) );
  XNOR U4065 ( .A(n3788), .B(n3789), .Z(out[1555]) );
  XNOR U4066 ( .A(n3792), .B(n3793), .Z(out[1554]) );
  XOR U4067 ( .A(n3796), .B(n3797), .Z(out[1553]) );
  XNOR U4068 ( .A(n3800), .B(n3801), .Z(out[1552]) );
  XNOR U4069 ( .A(n3804), .B(n3805), .Z(out[1551]) );
  XOR U4070 ( .A(n3806), .B(n3807), .Z(n3805) );
  NAND U4071 ( .A(n3808), .B(n3809), .Z(n3807) );
  AND U4072 ( .A(n3810), .B(n3811), .Z(n3809) );
  ANDN U4073 ( .B(n3812), .A(rc_i[18]), .Z(n3811) );
  NOR U4074 ( .A(rc_i[3]), .B(rc_i[4]), .Z(n3812) );
  NOR U4075 ( .A(rc_i[16]), .B(n3813), .Z(n3810) );
  AND U4076 ( .A(n3814), .B(n3815), .Z(n3808) );
  ANDN U4077 ( .B(n3597), .A(n3596), .Z(n3815) );
  NANDN U4078 ( .A(rc_i[20]), .B(n3816), .Z(n3596) );
  NOR U4079 ( .A(rc_i[23]), .B(rc_i[21]), .Z(n3816) );
  NOR U4080 ( .A(n3817), .B(n3818), .Z(n3814) );
  XNOR U4081 ( .A(n3821), .B(n3822), .Z(out[1550]) );
  XOR U4082 ( .A(n3825), .B(n3324), .Z(out[154]) );
  XOR U4083 ( .A(round_reg[691]), .B(n1945), .Z(n3324) );
  ANDN U4084 ( .B(n1452), .A(n1453), .Z(n3825) );
  XNOR U4085 ( .A(round_reg[216]), .B(n2279), .Z(n1453) );
  XNOR U4086 ( .A(round_reg[625]), .B(n2373), .Z(n1452) );
  XNOR U4087 ( .A(n3826), .B(n3827), .Z(out[1549]) );
  XOR U4088 ( .A(n3830), .B(n3831), .Z(out[1548]) );
  XNOR U4089 ( .A(n3834), .B(n3835), .Z(out[1547]) );
  XOR U4090 ( .A(n3838), .B(n3839), .Z(out[1546]) );
  XOR U4091 ( .A(n3842), .B(n3843), .Z(out[1545]) );
  XOR U4092 ( .A(n3846), .B(n3847), .Z(out[1544]) );
  XOR U4093 ( .A(n3850), .B(n3851), .Z(out[1543]) );
  XOR U4094 ( .A(n3852), .B(n3853), .Z(n3851) );
  NAND U4095 ( .A(n3854), .B(n3855), .Z(n3853) );
  AND U4096 ( .A(n3856), .B(n3857), .Z(n3855) );
  ANDN U4097 ( .B(n3858), .A(rc_i[6]), .Z(n3857) );
  ANDN U4098 ( .B(n3859), .A(rc_i[9]), .Z(n3858) );
  NOR U4099 ( .A(rc_i[20]), .B(rc_i[21]), .Z(n3856) );
  AND U4100 ( .A(n3860), .B(n3861), .Z(n3854) );
  ANDN U4101 ( .B(n3862), .A(rc_i[13]), .Z(n3861) );
  NOR U4102 ( .A(rc_i[17]), .B(rc_i[14]), .Z(n3862) );
  ANDN U4103 ( .B(n3740), .A(n3863), .Z(n3860) );
  XOR U4104 ( .A(n3866), .B(n3867), .Z(out[1542]) );
  XOR U4105 ( .A(n3870), .B(n3871), .Z(out[1541]) );
  XOR U4106 ( .A(n3874), .B(n3875), .Z(out[1540]) );
  XOR U4107 ( .A(n3878), .B(n3328), .Z(out[153]) );
  XOR U4108 ( .A(round_reg[690]), .B(n1948), .Z(n3328) );
  ANDN U4109 ( .B(n1500), .A(n1501), .Z(n3878) );
  XNOR U4110 ( .A(round_reg[215]), .B(n2283), .Z(n1501) );
  XNOR U4111 ( .A(round_reg[624]), .B(n2377), .Z(n1500) );
  XOR U4112 ( .A(n3879), .B(n3880), .Z(out[1539]) );
  XOR U4113 ( .A(n3881), .B(n3882), .Z(n3880) );
  NAND U4114 ( .A(n3883), .B(n3884), .Z(n3882) );
  AND U4115 ( .A(n3885), .B(n3886), .Z(n3884) );
  AND U4116 ( .A(n3887), .B(n3888), .Z(n3886) );
  NOR U4117 ( .A(rc_i[8]), .B(rc_i[9]), .Z(n3888) );
  NOR U4118 ( .A(rc_i[4]), .B(rc_i[7]), .Z(n3887) );
  ANDN U4119 ( .B(n3889), .A(rc_i[19]), .Z(n3885) );
  NOR U4120 ( .A(rc_i[23]), .B(rc_i[2]), .Z(n3889) );
  AND U4121 ( .A(n3890), .B(n3891), .Z(n3883) );
  ANDN U4122 ( .B(n3892), .A(rc_i[13]), .Z(n3891) );
  NOR U4123 ( .A(rc_i[18]), .B(rc_i[14]), .Z(n3892) );
  ANDN U4124 ( .B(n3893), .A(rc_i[10]), .Z(n3890) );
  ANDN U4125 ( .B(n3740), .A(rc_i[11]), .Z(n3893) );
  IV U4126 ( .A(rc_i[12]), .Z(n3740) );
  XOR U4127 ( .A(n3896), .B(n3897), .Z(out[1538]) );
  XOR U4128 ( .A(n3900), .B(n3901), .Z(out[1537]) );
  XOR U4129 ( .A(n3902), .B(n3903), .Z(n3901) );
  NAND U4130 ( .A(n3904), .B(n3905), .Z(n3903) );
  AND U4131 ( .A(n3906), .B(n3907), .Z(n3905) );
  ANDN U4132 ( .B(n3908), .A(rc_i[18]), .Z(n3907) );
  ANDN U4133 ( .B(n3859), .A(rc_i[19]), .Z(n3908) );
  IV U4134 ( .A(rc_i[8]), .Z(n3859) );
  NOR U4135 ( .A(rc_i[16]), .B(rc_i[15]), .Z(n3906) );
  AND U4136 ( .A(n3909), .B(n3910), .Z(n3904) );
  NOR U4137 ( .A(rc_i[12]), .B(rc_i[13]), .Z(n3910) );
  NOR U4138 ( .A(n3863), .B(rc_i[11]), .Z(n3909) );
  OR U4139 ( .A(n3818), .B(rc_i[4]), .Z(n3863) );
  OR U4140 ( .A(rc_i[1]), .B(rc_i[2]), .Z(n3818) );
  XOR U4141 ( .A(n3913), .B(n3914), .Z(out[1536]) );
  XOR U4142 ( .A(n3915), .B(n3916), .Z(n3914) );
  NAND U4143 ( .A(n3917), .B(n3918), .Z(n3916) );
  AND U4144 ( .A(n3919), .B(n3920), .Z(n3918) );
  NOR U4145 ( .A(rc_i[5]), .B(rc_i[4]), .Z(n3920) );
  NOR U4146 ( .A(rc_i[20]), .B(rc_i[22]), .Z(n3919) );
  AND U4147 ( .A(n3921), .B(n3922), .Z(n3917) );
  ANDN U4148 ( .B(n3597), .A(rc_i[0]), .Z(n3922) );
  NOR U4149 ( .A(rc_i[7]), .B(rc_i[6]), .Z(n3597) );
  NOR U4150 ( .A(n3817), .B(n3598), .Z(n3921) );
  OR U4151 ( .A(n3813), .B(rc_i[13]), .Z(n3598) );
  OR U4152 ( .A(rc_i[15]), .B(rc_i[14]), .Z(n3813) );
  OR U4153 ( .A(rc_i[10]), .B(rc_i[12]), .Z(n3817) );
  XOR U4154 ( .A(n3925), .B(n3600), .Z(out[1535]) );
  ANDN U4155 ( .B(n3926), .A(n3599), .Z(n3925) );
  XNOR U4156 ( .A(n3927), .B(n3604), .Z(out[1534]) );
  ANDN U4157 ( .B(n3928), .A(n3603), .Z(n3927) );
  XNOR U4158 ( .A(n3929), .B(n3608), .Z(out[1533]) );
  ANDN U4159 ( .B(n3930), .A(n3607), .Z(n3929) );
  XNOR U4160 ( .A(n3931), .B(n3612), .Z(out[1532]) );
  ANDN U4161 ( .B(n3932), .A(n3611), .Z(n3931) );
  XNOR U4162 ( .A(n3933), .B(n3616), .Z(out[1531]) );
  ANDN U4163 ( .B(n3934), .A(n3615), .Z(n3933) );
  XNOR U4164 ( .A(n3935), .B(n3620), .Z(out[1530]) );
  ANDN U4165 ( .B(n3936), .A(n3619), .Z(n3935) );
  XOR U4166 ( .A(n3937), .B(n3332), .Z(out[152]) );
  XOR U4167 ( .A(round_reg[689]), .B(n1951), .Z(n3332) );
  ANDN U4168 ( .B(n1534), .A(n1535), .Z(n3937) );
  XNOR U4169 ( .A(round_reg[214]), .B(n2287), .Z(n1535) );
  XNOR U4170 ( .A(round_reg[623]), .B(n2381), .Z(n1534) );
  XNOR U4171 ( .A(n3938), .B(n3624), .Z(out[1529]) );
  ANDN U4172 ( .B(n3939), .A(n3623), .Z(n3938) );
  XNOR U4173 ( .A(n3940), .B(n3628), .Z(out[1528]) );
  ANDN U4174 ( .B(n3941), .A(n3627), .Z(n3940) );
  XNOR U4175 ( .A(n3942), .B(n3632), .Z(out[1527]) );
  ANDN U4176 ( .B(n3943), .A(n3631), .Z(n3942) );
  XNOR U4177 ( .A(n3944), .B(n3636), .Z(out[1526]) );
  ANDN U4178 ( .B(n3945), .A(n3635), .Z(n3944) );
  XNOR U4179 ( .A(n3946), .B(n3641), .Z(out[1525]) );
  ANDN U4180 ( .B(n3947), .A(n3640), .Z(n3946) );
  XNOR U4181 ( .A(n3948), .B(n3645), .Z(out[1524]) );
  ANDN U4182 ( .B(n3949), .A(n3644), .Z(n3948) );
  XOR U4183 ( .A(n3950), .B(n3649), .Z(out[1523]) );
  ANDN U4184 ( .B(n3951), .A(n3648), .Z(n3950) );
  XNOR U4185 ( .A(n3952), .B(n3653), .Z(out[1522]) );
  ANDN U4186 ( .B(n3953), .A(n3652), .Z(n3952) );
  XNOR U4187 ( .A(n3954), .B(n3657), .Z(out[1521]) );
  ANDN U4188 ( .B(n3955), .A(n3656), .Z(n3954) );
  XNOR U4189 ( .A(n3956), .B(n3661), .Z(out[1520]) );
  ANDN U4190 ( .B(n3957), .A(n3660), .Z(n3956) );
  XOR U4191 ( .A(n3958), .B(n3337), .Z(out[151]) );
  XOR U4192 ( .A(round_reg[688]), .B(n1954), .Z(n3337) );
  ANDN U4193 ( .B(n1564), .A(n1565), .Z(n3958) );
  XNOR U4194 ( .A(round_reg[213]), .B(n2291), .Z(n1565) );
  XNOR U4195 ( .A(round_reg[622]), .B(n2385), .Z(n1564) );
  XNOR U4196 ( .A(n3959), .B(n3665), .Z(out[1519]) );
  ANDN U4197 ( .B(n3960), .A(n3664), .Z(n3959) );
  XNOR U4198 ( .A(n3961), .B(n3669), .Z(out[1518]) );
  ANDN U4199 ( .B(n3962), .A(n3668), .Z(n3961) );
  XNOR U4200 ( .A(n3963), .B(n3673), .Z(out[1517]) );
  ANDN U4201 ( .B(n3964), .A(n3672), .Z(n3963) );
  XNOR U4202 ( .A(n3965), .B(n3677), .Z(out[1516]) );
  ANDN U4203 ( .B(n3966), .A(n3676), .Z(n3965) );
  XNOR U4204 ( .A(n3967), .B(n3682), .Z(out[1515]) );
  ANDN U4205 ( .B(n3968), .A(n3681), .Z(n3967) );
  XOR U4206 ( .A(n3969), .B(n3686), .Z(out[1514]) );
  ANDN U4207 ( .B(n3970), .A(n3685), .Z(n3969) );
  XNOR U4208 ( .A(n3971), .B(n3690), .Z(out[1513]) );
  ANDN U4209 ( .B(n3972), .A(n3689), .Z(n3971) );
  XOR U4210 ( .A(n3973), .B(n3694), .Z(out[1512]) );
  ANDN U4211 ( .B(n3974), .A(n3693), .Z(n3973) );
  XOR U4212 ( .A(n3975), .B(n3698), .Z(out[1511]) );
  ANDN U4213 ( .B(n3976), .A(n3697), .Z(n3975) );
  XNOR U4214 ( .A(n3977), .B(n3702), .Z(out[1510]) );
  ANDN U4215 ( .B(n3978), .A(n3701), .Z(n3977) );
  XOR U4216 ( .A(n3979), .B(n3341), .Z(out[150]) );
  XOR U4217 ( .A(round_reg[687]), .B(n1961), .Z(n3341) );
  ANDN U4218 ( .B(n1589), .A(n1590), .Z(n3979) );
  XNOR U4219 ( .A(round_reg[212]), .B(n2295), .Z(n1590) );
  XNOR U4220 ( .A(round_reg[621]), .B(n2106), .Z(n1589) );
  XNOR U4221 ( .A(n3980), .B(n3706), .Z(out[1509]) );
  ANDN U4222 ( .B(n3981), .A(n3705), .Z(n3980) );
  XNOR U4223 ( .A(n3982), .B(n3710), .Z(out[1508]) );
  ANDN U4224 ( .B(n3983), .A(n3709), .Z(n3982) );
  XNOR U4225 ( .A(n3984), .B(n3714), .Z(out[1507]) );
  ANDN U4226 ( .B(n3985), .A(n3713), .Z(n3984) );
  XNOR U4227 ( .A(n3986), .B(n3717), .Z(out[1506]) );
  AND U4228 ( .A(n3987), .B(n3988), .Z(n3986) );
  IV U4229 ( .A(n3718), .Z(n3988) );
  XNOR U4230 ( .A(n3989), .B(n3722), .Z(out[1505]) );
  AND U4231 ( .A(n3990), .B(n3991), .Z(n3989) );
  IV U4232 ( .A(n3723), .Z(n3991) );
  XNOR U4233 ( .A(n3992), .B(n3726), .Z(out[1504]) );
  XNOR U4234 ( .A(n3994), .B(n3742), .Z(out[1503]) );
  ANDN U4235 ( .B(n3995), .A(n3741), .Z(n3994) );
  XNOR U4236 ( .A(n3996), .B(n3746), .Z(out[1502]) );
  ANDN U4237 ( .B(n3997), .A(n3745), .Z(n3996) );
  XNOR U4238 ( .A(n3998), .B(n3750), .Z(out[1501]) );
  ANDN U4239 ( .B(n3999), .A(n3749), .Z(n3998) );
  XNOR U4240 ( .A(n4000), .B(n3754), .Z(out[1500]) );
  ANDN U4241 ( .B(n4001), .A(n3753), .Z(n4000) );
  XNOR U4242 ( .A(n4002), .B(n1859), .Z(out[14]) );
  ANDN U4243 ( .B(n3372), .A(n3373), .Z(n4002) );
  XOR U4244 ( .A(round_reg[1047]), .B(n1765), .Z(n3373) );
  XNOR U4245 ( .A(round_reg[1424]), .B(n2290), .Z(n3372) );
  XOR U4246 ( .A(n4003), .B(n3345), .Z(out[149]) );
  XOR U4247 ( .A(round_reg[686]), .B(n1964), .Z(n3345) );
  ANDN U4248 ( .B(n1622), .A(n1623), .Z(n4003) );
  XNOR U4249 ( .A(round_reg[211]), .B(n2299), .Z(n1623) );
  XNOR U4250 ( .A(round_reg[620]), .B(n2110), .Z(n1622) );
  XNOR U4251 ( .A(n4004), .B(n3758), .Z(out[1499]) );
  ANDN U4252 ( .B(n4005), .A(n3757), .Z(n4004) );
  XNOR U4253 ( .A(n4006), .B(n3762), .Z(out[1498]) );
  ANDN U4254 ( .B(n4007), .A(n3761), .Z(n4006) );
  XOR U4255 ( .A(n4008), .B(n3766), .Z(out[1497]) );
  ANDN U4256 ( .B(n4009), .A(n3765), .Z(n4008) );
  XOR U4257 ( .A(n4010), .B(n3770), .Z(out[1496]) );
  ANDN U4258 ( .B(n4011), .A(n3769), .Z(n4010) );
  XOR U4259 ( .A(n4012), .B(n3775), .Z(out[1495]) );
  ANDN U4260 ( .B(n4013), .A(n3774), .Z(n4012) );
  XOR U4261 ( .A(n4014), .B(n3779), .Z(out[1494]) );
  ANDN U4262 ( .B(n4015), .A(n3778), .Z(n4014) );
  XOR U4263 ( .A(n4016), .B(n3783), .Z(out[1493]) );
  ANDN U4264 ( .B(n4017), .A(n3782), .Z(n4016) );
  XOR U4265 ( .A(n4018), .B(n3787), .Z(out[1492]) );
  ANDN U4266 ( .B(n4019), .A(n3786), .Z(n4018) );
  XOR U4267 ( .A(n4020), .B(n3791), .Z(out[1491]) );
  ANDN U4268 ( .B(n4021), .A(n3790), .Z(n4020) );
  XOR U4269 ( .A(n4022), .B(n3795), .Z(out[1490]) );
  ANDN U4270 ( .B(n4023), .A(n3794), .Z(n4022) );
  XOR U4271 ( .A(n4024), .B(n3349), .Z(out[148]) );
  XOR U4272 ( .A(round_reg[685]), .B(n1967), .Z(n3349) );
  ANDN U4273 ( .B(n1656), .A(n1657), .Z(n4024) );
  XNOR U4274 ( .A(round_reg[210]), .B(n2307), .Z(n1657) );
  XNOR U4275 ( .A(round_reg[619]), .B(n2114), .Z(n1656) );
  IV U4276 ( .A(n4025), .Z(n2114) );
  XOR U4277 ( .A(n4026), .B(n3799), .Z(out[1489]) );
  ANDN U4278 ( .B(n4027), .A(n3798), .Z(n4026) );
  XOR U4279 ( .A(n4028), .B(n3803), .Z(out[1488]) );
  ANDN U4280 ( .B(n4029), .A(n3802), .Z(n4028) );
  XOR U4281 ( .A(n4030), .B(n3820), .Z(out[1487]) );
  ANDN U4282 ( .B(n4031), .A(n3819), .Z(n4030) );
  XOR U4283 ( .A(n4032), .B(n3824), .Z(out[1486]) );
  ANDN U4284 ( .B(n4033), .A(n3823), .Z(n4032) );
  XOR U4285 ( .A(n4034), .B(n3829), .Z(out[1485]) );
  ANDN U4286 ( .B(n4035), .A(n3828), .Z(n4034) );
  XOR U4287 ( .A(n4036), .B(n3833), .Z(out[1484]) );
  ANDN U4288 ( .B(n4037), .A(n3832), .Z(n4036) );
  XOR U4289 ( .A(n4038), .B(n3837), .Z(out[1483]) );
  ANDN U4290 ( .B(n4039), .A(n3836), .Z(n4038) );
  XOR U4291 ( .A(n4040), .B(n3841), .Z(out[1482]) );
  ANDN U4292 ( .B(n4041), .A(n3840), .Z(n4040) );
  XOR U4293 ( .A(n4042), .B(n3845), .Z(out[1481]) );
  ANDN U4294 ( .B(n4043), .A(n3844), .Z(n4042) );
  XOR U4295 ( .A(n4044), .B(n3849), .Z(out[1480]) );
  ANDN U4296 ( .B(n4045), .A(n3848), .Z(n4044) );
  XOR U4297 ( .A(n4046), .B(n3353), .Z(out[147]) );
  XOR U4298 ( .A(round_reg[684]), .B(n1970), .Z(n3353) );
  ANDN U4299 ( .B(n1690), .A(n1691), .Z(n4046) );
  XNOR U4300 ( .A(round_reg[209]), .B(n2311), .Z(n1691) );
  XNOR U4301 ( .A(round_reg[618]), .B(n2118), .Z(n1690) );
  IV U4302 ( .A(n4047), .Z(n2118) );
  XOR U4303 ( .A(n4048), .B(n3865), .Z(out[1479]) );
  ANDN U4304 ( .B(n4049), .A(n3864), .Z(n4048) );
  XOR U4305 ( .A(n4050), .B(n3869), .Z(out[1478]) );
  ANDN U4306 ( .B(n4051), .A(n3868), .Z(n4050) );
  XOR U4307 ( .A(n4052), .B(n3873), .Z(out[1477]) );
  ANDN U4308 ( .B(n4053), .A(n3872), .Z(n4052) );
  XOR U4309 ( .A(n4054), .B(n3877), .Z(out[1476]) );
  ANDN U4310 ( .B(n4055), .A(n3876), .Z(n4054) );
  XOR U4311 ( .A(n4056), .B(n3895), .Z(out[1475]) );
  ANDN U4312 ( .B(n4057), .A(n3894), .Z(n4056) );
  XOR U4313 ( .A(n4058), .B(n3899), .Z(out[1474]) );
  ANDN U4314 ( .B(n4059), .A(n3898), .Z(n4058) );
  XOR U4315 ( .A(n4060), .B(n3912), .Z(out[1473]) );
  ANDN U4316 ( .B(n4061), .A(n3911), .Z(n4060) );
  XOR U4317 ( .A(n4062), .B(n3924), .Z(out[1472]) );
  ANDN U4318 ( .B(n4063), .A(n3923), .Z(n4062) );
  XOR U4319 ( .A(n4064), .B(n3599), .Z(out[1471]) );
  XOR U4320 ( .A(round_reg[788]), .B(n2274), .Z(n3599) );
  ANDN U4321 ( .B(n4065), .A(n3926), .Z(n4064) );
  XOR U4322 ( .A(n4066), .B(n3603), .Z(out[1470]) );
  XOR U4323 ( .A(round_reg[787]), .B(n2278), .Z(n3603) );
  ANDN U4324 ( .B(n4067), .A(n3928), .Z(n4066) );
  XOR U4325 ( .A(n4068), .B(n3358), .Z(out[146]) );
  XOR U4326 ( .A(round_reg[683]), .B(n1973), .Z(n3358) );
  ANDN U4327 ( .B(n1718), .A(n1719), .Z(n4068) );
  XNOR U4328 ( .A(round_reg[208]), .B(n2315), .Z(n1719) );
  XNOR U4329 ( .A(round_reg[617]), .B(n2129), .Z(n1718) );
  IV U4330 ( .A(n4069), .Z(n2129) );
  XOR U4331 ( .A(n4070), .B(n3607), .Z(out[1469]) );
  XOR U4332 ( .A(round_reg[786]), .B(n2282), .Z(n3607) );
  ANDN U4333 ( .B(n4071), .A(n3930), .Z(n4070) );
  XOR U4334 ( .A(n4072), .B(n3611), .Z(out[1468]) );
  XOR U4335 ( .A(round_reg[785]), .B(n2286), .Z(n3611) );
  ANDN U4336 ( .B(n4073), .A(n3932), .Z(n4072) );
  XOR U4337 ( .A(n4074), .B(n3615), .Z(out[1467]) );
  XOR U4338 ( .A(round_reg[784]), .B(n2290), .Z(n3615) );
  ANDN U4339 ( .B(n4075), .A(n3934), .Z(n4074) );
  XOR U4340 ( .A(n4076), .B(n3619), .Z(out[1466]) );
  XOR U4341 ( .A(round_reg[783]), .B(n2294), .Z(n3619) );
  ANDN U4342 ( .B(n4077), .A(n3936), .Z(n4076) );
  XOR U4343 ( .A(n4078), .B(n3623), .Z(out[1465]) );
  XOR U4344 ( .A(round_reg[782]), .B(n2298), .Z(n3623) );
  ANDN U4345 ( .B(n4079), .A(n3939), .Z(n4078) );
  XOR U4346 ( .A(n4080), .B(n3627), .Z(out[1464]) );
  XOR U4347 ( .A(round_reg[781]), .B(n2306), .Z(n3627) );
  ANDN U4348 ( .B(n4081), .A(n3941), .Z(n4080) );
  XOR U4349 ( .A(n4082), .B(n3631), .Z(out[1463]) );
  XOR U4350 ( .A(round_reg[780]), .B(n2310), .Z(n3631) );
  ANDN U4351 ( .B(n4083), .A(n3943), .Z(n4082) );
  XOR U4352 ( .A(n4084), .B(n3635), .Z(out[1462]) );
  XOR U4353 ( .A(round_reg[779]), .B(n2314), .Z(n3635) );
  ANDN U4354 ( .B(n4085), .A(n3945), .Z(n4084) );
  XOR U4355 ( .A(n4086), .B(n3640), .Z(out[1461]) );
  XOR U4356 ( .A(round_reg[778]), .B(n2318), .Z(n3640) );
  ANDN U4357 ( .B(n4087), .A(n3947), .Z(n4086) );
  XOR U4358 ( .A(n4088), .B(n3644), .Z(out[1460]) );
  XOR U4359 ( .A(round_reg[777]), .B(n2322), .Z(n3644) );
  ANDN U4360 ( .B(n4089), .A(n3949), .Z(n4088) );
  XOR U4361 ( .A(n4090), .B(n3362), .Z(out[145]) );
  XOR U4362 ( .A(round_reg[682]), .B(n1975), .Z(n3362) );
  ANDN U4363 ( .B(n1752), .A(n1753), .Z(n4090) );
  XNOR U4364 ( .A(round_reg[207]), .B(n2319), .Z(n1753) );
  XNOR U4365 ( .A(round_reg[616]), .B(n2133), .Z(n1752) );
  IV U4366 ( .A(n4091), .Z(n2133) );
  XOR U4367 ( .A(n4092), .B(n3648), .Z(out[1459]) );
  XOR U4368 ( .A(round_reg[776]), .B(n2326), .Z(n3648) );
  ANDN U4369 ( .B(n4093), .A(n3951), .Z(n4092) );
  XOR U4370 ( .A(n4094), .B(n3652), .Z(out[1458]) );
  XOR U4371 ( .A(round_reg[775]), .B(n2330), .Z(n3652) );
  ANDN U4372 ( .B(n4095), .A(n3953), .Z(n4094) );
  XOR U4373 ( .A(n4096), .B(n3656), .Z(out[1457]) );
  XOR U4374 ( .A(round_reg[774]), .B(n2334), .Z(n3656) );
  ANDN U4375 ( .B(n4097), .A(n3955), .Z(n4096) );
  XOR U4376 ( .A(n4098), .B(n3660), .Z(out[1456]) );
  XOR U4377 ( .A(round_reg[773]), .B(n2338), .Z(n3660) );
  ANDN U4378 ( .B(n4099), .A(n3957), .Z(n4098) );
  XOR U4379 ( .A(n4100), .B(n3664), .Z(out[1455]) );
  XOR U4380 ( .A(round_reg[772]), .B(n2342), .Z(n3664) );
  ANDN U4381 ( .B(n4101), .A(n3960), .Z(n4100) );
  XOR U4382 ( .A(n4102), .B(n3668), .Z(out[1454]) );
  XOR U4383 ( .A(round_reg[771]), .B(n2350), .Z(n3668) );
  ANDN U4384 ( .B(n4103), .A(n3962), .Z(n4102) );
  XOR U4385 ( .A(n4104), .B(n3672), .Z(out[1453]) );
  XOR U4386 ( .A(round_reg[770]), .B(n2354), .Z(n3672) );
  ANDN U4387 ( .B(n4105), .A(n3964), .Z(n4104) );
  XOR U4388 ( .A(n4106), .B(n3676), .Z(out[1452]) );
  XOR U4389 ( .A(round_reg[769]), .B(n2358), .Z(n3676) );
  ANDN U4390 ( .B(n4107), .A(n3966), .Z(n4106) );
  XOR U4391 ( .A(n4108), .B(n3681), .Z(out[1451]) );
  XOR U4392 ( .A(round_reg[768]), .B(n2362), .Z(n3681) );
  ANDN U4393 ( .B(n4109), .A(n3968), .Z(n4108) );
  XOR U4394 ( .A(n4110), .B(n3685), .Z(out[1450]) );
  XOR U4395 ( .A(round_reg[831]), .B(n2366), .Z(n3685) );
  ANDN U4396 ( .B(n4111), .A(n3970), .Z(n4110) );
  XOR U4397 ( .A(n4112), .B(n3366), .Z(out[144]) );
  IV U4398 ( .A(n3501), .Z(n3366) );
  XNOR U4399 ( .A(round_reg[681]), .B(n1977), .Z(n3501) );
  ANDN U4400 ( .B(n1786), .A(n1787), .Z(n4112) );
  XNOR U4401 ( .A(round_reg[206]), .B(n2323), .Z(n1787) );
  XNOR U4402 ( .A(round_reg[615]), .B(n2137), .Z(n1786) );
  IV U4403 ( .A(n4113), .Z(n2137) );
  XOR U4404 ( .A(n4114), .B(n3689), .Z(out[1449]) );
  XOR U4405 ( .A(round_reg[830]), .B(n2370), .Z(n3689) );
  ANDN U4406 ( .B(n4115), .A(n3972), .Z(n4114) );
  XOR U4407 ( .A(n4116), .B(n3693), .Z(out[1448]) );
  XOR U4408 ( .A(round_reg[829]), .B(n2374), .Z(n3693) );
  ANDN U4409 ( .B(n4117), .A(n3974), .Z(n4116) );
  XOR U4410 ( .A(n4118), .B(n3697), .Z(out[1447]) );
  XOR U4411 ( .A(round_reg[828]), .B(n2378), .Z(n3697) );
  ANDN U4412 ( .B(n4119), .A(n3976), .Z(n4118) );
  XOR U4413 ( .A(n4120), .B(n3701), .Z(out[1446]) );
  XOR U4414 ( .A(round_reg[827]), .B(n2382), .Z(n3701) );
  XOR U4415 ( .A(n4122), .B(n3705), .Z(out[1445]) );
  XOR U4416 ( .A(round_reg[826]), .B(n2386), .Z(n3705) );
  XOR U4417 ( .A(n4124), .B(n3709), .Z(out[1444]) );
  XNOR U4418 ( .A(round_reg[825]), .B(n4125), .Z(n3709) );
  AND U4419 ( .A(n4126), .B(n4127), .Z(n4124) );
  IV U4420 ( .A(n3983), .Z(n4127) );
  XOR U4421 ( .A(n4128), .B(n3713), .Z(out[1443]) );
  XNOR U4422 ( .A(round_reg[824]), .B(n4129), .Z(n3713) );
  AND U4423 ( .A(n4130), .B(n4131), .Z(n4128) );
  IV U4424 ( .A(n3985), .Z(n4131) );
  XOR U4425 ( .A(n4132), .B(n3718), .Z(out[1442]) );
  XOR U4426 ( .A(round_reg[823]), .B(n2116), .Z(n3718) );
  AND U4427 ( .A(n4133), .B(n4134), .Z(n4132) );
  IV U4428 ( .A(n3987), .Z(n4134) );
  XOR U4429 ( .A(n4135), .B(n3723), .Z(out[1441]) );
  XOR U4430 ( .A(round_reg[822]), .B(n2120), .Z(n3723) );
  XOR U4431 ( .A(n4137), .B(n3727), .Z(out[1440]) );
  XOR U4432 ( .A(round_reg[821]), .B(n2131), .Z(n3727) );
  ANDN U4433 ( .B(n4138), .A(n3993), .Z(n4137) );
  XOR U4434 ( .A(n4139), .B(n3370), .Z(out[143]) );
  IV U4435 ( .A(n3503), .Z(n3370) );
  XNOR U4436 ( .A(round_reg[680]), .B(n1980), .Z(n3503) );
  ANDN U4437 ( .B(n1824), .A(n1825), .Z(n4139) );
  XNOR U4438 ( .A(round_reg[205]), .B(n2327), .Z(n1825) );
  XNOR U4439 ( .A(round_reg[614]), .B(n2141), .Z(n1824) );
  IV U4440 ( .A(n4140), .Z(n2141) );
  XOR U4441 ( .A(n4141), .B(n3741), .Z(out[1439]) );
  XOR U4442 ( .A(round_reg[820]), .B(n2134), .Z(n3741) );
  ANDN U4443 ( .B(n4142), .A(n3995), .Z(n4141) );
  XOR U4444 ( .A(n4143), .B(n3745), .Z(out[1438]) );
  XOR U4445 ( .A(round_reg[819]), .B(n2138), .Z(n3745) );
  ANDN U4446 ( .B(n4144), .A(n3997), .Z(n4143) );
  XOR U4447 ( .A(n4145), .B(n3749), .Z(out[1437]) );
  XOR U4448 ( .A(round_reg[818]), .B(n2142), .Z(n3749) );
  ANDN U4449 ( .B(n4146), .A(n3999), .Z(n4145) );
  XOR U4450 ( .A(n4147), .B(n3753), .Z(out[1436]) );
  XOR U4451 ( .A(round_reg[817]), .B(n2146), .Z(n3753) );
  ANDN U4452 ( .B(n4148), .A(n4001), .Z(n4147) );
  XOR U4453 ( .A(n4149), .B(n3757), .Z(out[1435]) );
  XOR U4454 ( .A(round_reg[816]), .B(n2150), .Z(n3757) );
  ANDN U4455 ( .B(n4150), .A(n4005), .Z(n4149) );
  XOR U4456 ( .A(n4151), .B(n3761), .Z(out[1434]) );
  XOR U4457 ( .A(round_reg[815]), .B(n2154), .Z(n3761) );
  ANDN U4458 ( .B(n4152), .A(n4007), .Z(n4151) );
  XOR U4459 ( .A(n4153), .B(n3765), .Z(out[1433]) );
  XOR U4460 ( .A(round_reg[814]), .B(n2158), .Z(n3765) );
  ANDN U4461 ( .B(n4154), .A(n4009), .Z(n4153) );
  XOR U4462 ( .A(n4155), .B(n3769), .Z(out[1432]) );
  XOR U4463 ( .A(round_reg[813]), .B(n2162), .Z(n3769) );
  ANDN U4464 ( .B(n4156), .A(n4011), .Z(n4155) );
  XOR U4465 ( .A(n4157), .B(n3774), .Z(out[1431]) );
  XOR U4466 ( .A(round_reg[812]), .B(n2166), .Z(n3774) );
  ANDN U4467 ( .B(n4158), .A(n4013), .Z(n4157) );
  XOR U4468 ( .A(n4159), .B(n3778), .Z(out[1430]) );
  XOR U4469 ( .A(round_reg[811]), .B(n2174), .Z(n3778) );
  ANDN U4470 ( .B(n4160), .A(n4015), .Z(n4159) );
  XOR U4471 ( .A(n4161), .B(n3374), .Z(out[142]) );
  IV U4472 ( .A(n3505), .Z(n3374) );
  XNOR U4473 ( .A(round_reg[679]), .B(n1983), .Z(n3505) );
  ANDN U4474 ( .B(n1858), .A(n1859), .Z(n4161) );
  XNOR U4475 ( .A(round_reg[204]), .B(n2331), .Z(n1859) );
  XNOR U4476 ( .A(round_reg[613]), .B(n2145), .Z(n1858) );
  IV U4477 ( .A(n4162), .Z(n2145) );
  XOR U4478 ( .A(n4163), .B(n3782), .Z(out[1429]) );
  XOR U4479 ( .A(round_reg[810]), .B(n2178), .Z(n3782) );
  ANDN U4480 ( .B(n4164), .A(n4017), .Z(n4163) );
  XOR U4481 ( .A(n4165), .B(n3786), .Z(out[1428]) );
  XOR U4482 ( .A(round_reg[809]), .B(n2182), .Z(n3786) );
  ANDN U4483 ( .B(n4166), .A(n4019), .Z(n4165) );
  XOR U4484 ( .A(n4167), .B(n3790), .Z(out[1427]) );
  XOR U4485 ( .A(round_reg[808]), .B(n2186), .Z(n3790) );
  ANDN U4486 ( .B(n4168), .A(n4021), .Z(n4167) );
  XOR U4487 ( .A(n4169), .B(n3794), .Z(out[1426]) );
  XOR U4488 ( .A(round_reg[807]), .B(n2190), .Z(n3794) );
  ANDN U4489 ( .B(n4170), .A(n4023), .Z(n4169) );
  XOR U4490 ( .A(n4171), .B(n3798), .Z(out[1425]) );
  XOR U4491 ( .A(round_reg[806]), .B(n2194), .Z(n3798) );
  ANDN U4492 ( .B(n4172), .A(n4027), .Z(n4171) );
  XOR U4493 ( .A(n4173), .B(n3802), .Z(out[1424]) );
  XOR U4494 ( .A(round_reg[805]), .B(n2198), .Z(n3802) );
  ANDN U4495 ( .B(n4174), .A(n4029), .Z(n4173) );
  XOR U4496 ( .A(n4175), .B(n3819), .Z(out[1423]) );
  XOR U4497 ( .A(round_reg[804]), .B(n2202), .Z(n3819) );
  ANDN U4498 ( .B(n4176), .A(n4031), .Z(n4175) );
  XOR U4499 ( .A(n4177), .B(n3823), .Z(out[1422]) );
  XNOR U4500 ( .A(round_reg[803]), .B(n3032), .Z(n3823) );
  ANDN U4501 ( .B(n4178), .A(n4033), .Z(n4177) );
  XOR U4502 ( .A(n4179), .B(n3828), .Z(out[1421]) );
  XOR U4503 ( .A(round_reg[802]), .B(n2210), .Z(n3828) );
  ANDN U4504 ( .B(n4180), .A(n4035), .Z(n4179) );
  XOR U4505 ( .A(n4181), .B(n3832), .Z(out[1420]) );
  XOR U4506 ( .A(round_reg[801]), .B(n2218), .Z(n3832) );
  ANDN U4507 ( .B(n4182), .A(n4037), .Z(n4181) );
  XOR U4508 ( .A(n4183), .B(n3379), .Z(out[141]) );
  IV U4509 ( .A(n3507), .Z(n3379) );
  XNOR U4510 ( .A(round_reg[678]), .B(n1986), .Z(n3507) );
  AND U4511 ( .A(n1892), .B(n1894), .Z(n4183) );
  XNOR U4512 ( .A(round_reg[612]), .B(n2149), .Z(n1892) );
  XOR U4513 ( .A(n4184), .B(n3836), .Z(out[1419]) );
  XOR U4514 ( .A(round_reg[800]), .B(n2222), .Z(n3836) );
  ANDN U4515 ( .B(n4185), .A(n4039), .Z(n4184) );
  XOR U4516 ( .A(n4186), .B(n3840), .Z(out[1418]) );
  XOR U4517 ( .A(round_reg[799]), .B(n2226), .Z(n3840) );
  ANDN U4518 ( .B(n4187), .A(n4041), .Z(n4186) );
  XOR U4519 ( .A(n4188), .B(n3844), .Z(out[1417]) );
  XOR U4520 ( .A(round_reg[798]), .B(n2230), .Z(n3844) );
  ANDN U4521 ( .B(n4189), .A(n4043), .Z(n4188) );
  XOR U4522 ( .A(n4190), .B(n3848), .Z(out[1416]) );
  XOR U4523 ( .A(round_reg[797]), .B(n2234), .Z(n3848) );
  ANDN U4524 ( .B(n4191), .A(n4045), .Z(n4190) );
  XOR U4525 ( .A(n4192), .B(n3864), .Z(out[1415]) );
  XOR U4526 ( .A(round_reg[796]), .B(n2238), .Z(n3864) );
  ANDN U4527 ( .B(n4193), .A(n4049), .Z(n4192) );
  XOR U4528 ( .A(n4194), .B(n3868), .Z(out[1414]) );
  XOR U4529 ( .A(round_reg[795]), .B(n2242), .Z(n3868) );
  ANDN U4530 ( .B(n4195), .A(n4051), .Z(n4194) );
  XOR U4531 ( .A(n4196), .B(n3872), .Z(out[1413]) );
  XOR U4532 ( .A(round_reg[794]), .B(n2246), .Z(n3872) );
  ANDN U4533 ( .B(n4197), .A(n4053), .Z(n4196) );
  XOR U4534 ( .A(n4198), .B(n3876), .Z(out[1412]) );
  XOR U4535 ( .A(round_reg[793]), .B(n2250), .Z(n3876) );
  ANDN U4536 ( .B(n4199), .A(n4055), .Z(n4198) );
  XOR U4537 ( .A(n4200), .B(n3894), .Z(out[1411]) );
  XOR U4538 ( .A(round_reg[792]), .B(n2254), .Z(n3894) );
  ANDN U4539 ( .B(n4201), .A(n4057), .Z(n4200) );
  XOR U4540 ( .A(n4202), .B(n3898), .Z(out[1410]) );
  XOR U4541 ( .A(round_reg[791]), .B(n2262), .Z(n3898) );
  ANDN U4542 ( .B(n4203), .A(n4059), .Z(n4202) );
  XOR U4543 ( .A(n4204), .B(n3383), .Z(out[140]) );
  IV U4544 ( .A(n3509), .Z(n3383) );
  XNOR U4545 ( .A(round_reg[677]), .B(n1993), .Z(n3509) );
  AND U4546 ( .A(n1926), .B(n1928), .Z(n4204) );
  XNOR U4547 ( .A(round_reg[611]), .B(n2153), .Z(n1926) );
  IV U4548 ( .A(n4205), .Z(n2153) );
  XOR U4549 ( .A(n4206), .B(n3911), .Z(out[1409]) );
  XOR U4550 ( .A(round_reg[790]), .B(n2266), .Z(n3911) );
  ANDN U4551 ( .B(n4207), .A(n4061), .Z(n4206) );
  XOR U4552 ( .A(n4208), .B(n3923), .Z(out[1408]) );
  XOR U4553 ( .A(round_reg[789]), .B(n2270), .Z(n3923) );
  ANDN U4554 ( .B(n4209), .A(n4063), .Z(n4208) );
  XOR U4555 ( .A(n4210), .B(n3926), .Z(out[1407]) );
  XNOR U4556 ( .A(round_reg[426]), .B(n1920), .Z(n3926) );
  ANDN U4557 ( .B(n3586), .A(n4065), .Z(n4210) );
  XOR U4558 ( .A(n4211), .B(n3928), .Z(out[1406]) );
  XNOR U4559 ( .A(round_reg[425]), .B(n1923), .Z(n3928) );
  ANDN U4560 ( .B(n3602), .A(n4067), .Z(n4211) );
  XOR U4561 ( .A(n4212), .B(n3930), .Z(out[1405]) );
  XNOR U4562 ( .A(round_reg[424]), .B(n1930), .Z(n3930) );
  ANDN U4563 ( .B(n3606), .A(n4071), .Z(n4212) );
  XOR U4564 ( .A(n4213), .B(n3932), .Z(out[1404]) );
  XNOR U4565 ( .A(round_reg[423]), .B(n1933), .Z(n3932) );
  ANDN U4566 ( .B(n3610), .A(n4073), .Z(n4213) );
  XOR U4567 ( .A(n4214), .B(n3934), .Z(out[1403]) );
  XNOR U4568 ( .A(round_reg[422]), .B(n1712), .Z(n3934) );
  ANDN U4569 ( .B(n3614), .A(n4075), .Z(n4214) );
  XOR U4570 ( .A(n4215), .B(n3936), .Z(out[1402]) );
  XNOR U4571 ( .A(round_reg[421]), .B(n1715), .Z(n3936) );
  ANDN U4572 ( .B(n3618), .A(n4077), .Z(n4215) );
  XOR U4573 ( .A(n4216), .B(n3939), .Z(out[1401]) );
  XNOR U4574 ( .A(round_reg[420]), .B(n1722), .Z(n3939) );
  XOR U4575 ( .A(n4217), .B(n3941), .Z(out[1400]) );
  XNOR U4576 ( .A(round_reg[419]), .B(n1725), .Z(n3941) );
  XOR U4577 ( .A(n4218), .B(n1894), .Z(out[13]) );
  XOR U4578 ( .A(round_reg[203]), .B(n2335), .Z(n1894) );
  ANDN U4579 ( .B(n3377), .A(n3378), .Z(n4218) );
  XOR U4580 ( .A(round_reg[1046]), .B(n1768), .Z(n3378) );
  XNOR U4581 ( .A(round_reg[1423]), .B(n2294), .Z(n3377) );
  XOR U4582 ( .A(n4219), .B(n3387), .Z(out[139]) );
  IV U4583 ( .A(n3511), .Z(n3387) );
  XNOR U4584 ( .A(round_reg[676]), .B(n1996), .Z(n3511) );
  AND U4585 ( .A(n1957), .B(n1959), .Z(n4219) );
  XNOR U4586 ( .A(round_reg[610]), .B(n2157), .Z(n1957) );
  IV U4587 ( .A(n4220), .Z(n2157) );
  XOR U4588 ( .A(n4221), .B(n3943), .Z(out[1399]) );
  XOR U4589 ( .A(round_reg[418]), .B(n1728), .Z(n3943) );
  ANDN U4590 ( .B(n3630), .A(n4083), .Z(n4221) );
  XOR U4591 ( .A(n4222), .B(n3945), .Z(out[1398]) );
  XOR U4592 ( .A(round_reg[417]), .B(n1731), .Z(n3945) );
  ANDN U4593 ( .B(n3634), .A(n4085), .Z(n4222) );
  XOR U4594 ( .A(n4223), .B(n3947), .Z(out[1397]) );
  XOR U4595 ( .A(round_reg[416]), .B(n1734), .Z(n3947) );
  ANDN U4596 ( .B(n3639), .A(n4087), .Z(n4223) );
  XOR U4597 ( .A(n4224), .B(n3949), .Z(out[1396]) );
  XOR U4598 ( .A(round_reg[415]), .B(n1737), .Z(n3949) );
  ANDN U4599 ( .B(n3643), .A(n4089), .Z(n4224) );
  XOR U4600 ( .A(n4225), .B(n3951), .Z(out[1395]) );
  XOR U4601 ( .A(round_reg[414]), .B(n1740), .Z(n3951) );
  ANDN U4602 ( .B(n3647), .A(n4093), .Z(n4225) );
  XOR U4603 ( .A(n4226), .B(n3953), .Z(out[1394]) );
  XOR U4604 ( .A(round_reg[413]), .B(n1743), .Z(n3953) );
  ANDN U4605 ( .B(n3651), .A(n4095), .Z(n4226) );
  XOR U4606 ( .A(n4227), .B(n3955), .Z(out[1393]) );
  XOR U4607 ( .A(round_reg[412]), .B(n1746), .Z(n3955) );
  ANDN U4608 ( .B(n3655), .A(n4097), .Z(n4227) );
  XOR U4609 ( .A(n4228), .B(n3957), .Z(out[1392]) );
  XOR U4610 ( .A(round_reg[411]), .B(n1749), .Z(n3957) );
  ANDN U4611 ( .B(n3659), .A(n4099), .Z(n4228) );
  XOR U4612 ( .A(n4229), .B(n3960), .Z(out[1391]) );
  XNOR U4613 ( .A(round_reg[410]), .B(n1756), .Z(n3960) );
  AND U4614 ( .A(n3663), .B(n4230), .Z(n4229) );
  IV U4615 ( .A(n4101), .Z(n4230) );
  XOR U4616 ( .A(n4231), .B(n3962), .Z(out[1390]) );
  XNOR U4617 ( .A(round_reg[409]), .B(n1759), .Z(n3962) );
  AND U4618 ( .A(n3667), .B(n4232), .Z(n4231) );
  IV U4619 ( .A(n4103), .Z(n4232) );
  XOR U4620 ( .A(n4233), .B(n3391), .Z(out[138]) );
  IV U4621 ( .A(n3513), .Z(n3391) );
  XNOR U4622 ( .A(round_reg[675]), .B(n1999), .Z(n3513) );
  AND U4623 ( .A(n1989), .B(n1991), .Z(n4233) );
  XNOR U4624 ( .A(round_reg[609]), .B(n2161), .Z(n1989) );
  XOR U4625 ( .A(n4234), .B(n3964), .Z(out[1389]) );
  XNOR U4626 ( .A(round_reg[408]), .B(n1762), .Z(n3964) );
  AND U4627 ( .A(n3671), .B(n4235), .Z(n4234) );
  IV U4628 ( .A(n4105), .Z(n4235) );
  XOR U4629 ( .A(n4236), .B(n3966), .Z(out[1388]) );
  XNOR U4630 ( .A(round_reg[407]), .B(n1765), .Z(n3966) );
  XOR U4631 ( .A(n4237), .B(n3968), .Z(out[1387]) );
  XNOR U4632 ( .A(round_reg[406]), .B(n1768), .Z(n3968) );
  XOR U4633 ( .A(n4238), .B(n3970), .Z(out[1386]) );
  XNOR U4634 ( .A(round_reg[405]), .B(n1771), .Z(n3970) );
  ANDN U4635 ( .B(n3684), .A(n4111), .Z(n4238) );
  XOR U4636 ( .A(n4239), .B(n3972), .Z(out[1385]) );
  XNOR U4637 ( .A(round_reg[404]), .B(n1774), .Z(n3972) );
  ANDN U4638 ( .B(n3688), .A(n4115), .Z(n4239) );
  XOR U4639 ( .A(n4240), .B(n3974), .Z(out[1384]) );
  XNOR U4640 ( .A(round_reg[403]), .B(n1777), .Z(n3974) );
  ANDN U4641 ( .B(n3692), .A(n4117), .Z(n4240) );
  XOR U4642 ( .A(n4241), .B(n3976), .Z(out[1383]) );
  XOR U4643 ( .A(round_reg[402]), .B(n1780), .Z(n3976) );
  ANDN U4644 ( .B(n3696), .A(n4119), .Z(n4241) );
  XOR U4645 ( .A(n4242), .B(n3978), .Z(out[1382]) );
  XOR U4646 ( .A(round_reg[401]), .B(n1783), .Z(n3978) );
  IV U4647 ( .A(n4243), .Z(n1783) );
  ANDN U4648 ( .B(n3700), .A(n4121), .Z(n4242) );
  XOR U4649 ( .A(n4244), .B(n3981), .Z(out[1381]) );
  XOR U4650 ( .A(round_reg[400]), .B(n1790), .Z(n3981) );
  IV U4651 ( .A(n4245), .Z(n1790) );
  ANDN U4652 ( .B(n3704), .A(n4123), .Z(n4244) );
  XOR U4653 ( .A(n4246), .B(n3983), .Z(out[1380]) );
  XOR U4654 ( .A(round_reg[399]), .B(n1793), .Z(n3983) );
  IV U4655 ( .A(n4247), .Z(n1793) );
  NOR U4656 ( .A(n4126), .B(n3708), .Z(n4246) );
  XOR U4657 ( .A(n4248), .B(n3515), .Z(out[137]) );
  XOR U4658 ( .A(round_reg[674]), .B(n2002), .Z(n3515) );
  IV U4659 ( .A(n4249), .Z(n2002) );
  AND U4660 ( .A(n2017), .B(n1052), .Z(n4248) );
  IV U4661 ( .A(n2018), .Z(n1052) );
  XNOR U4662 ( .A(round_reg[199]), .B(n2355), .Z(n2018) );
  XNOR U4663 ( .A(round_reg[608]), .B(n2165), .Z(n2017) );
  XOR U4664 ( .A(n4250), .B(n3985), .Z(out[1379]) );
  XOR U4665 ( .A(round_reg[398]), .B(n1796), .Z(n3985) );
  IV U4666 ( .A(n4251), .Z(n1796) );
  ANDN U4667 ( .B(n3712), .A(n4130), .Z(n4250) );
  XOR U4668 ( .A(n4252), .B(n3987), .Z(out[1378]) );
  XOR U4669 ( .A(round_reg[397]), .B(n1799), .Z(n3987) );
  IV U4670 ( .A(n4253), .Z(n1799) );
  ANDN U4671 ( .B(n3716), .A(n4133), .Z(n4252) );
  XOR U4672 ( .A(n4254), .B(n3990), .Z(out[1377]) );
  XOR U4673 ( .A(round_reg[396]), .B(n1802), .Z(n3990) );
  IV U4674 ( .A(n4255), .Z(n1802) );
  NOR U4675 ( .A(n4136), .B(n3721), .Z(n4254) );
  XOR U4676 ( .A(n4256), .B(n3993), .Z(out[1376]) );
  XOR U4677 ( .A(round_reg[395]), .B(n1805), .Z(n3993) );
  NOR U4678 ( .A(n3725), .B(n4138), .Z(n4256) );
  XOR U4679 ( .A(n4257), .B(n3995), .Z(out[1375]) );
  XOR U4680 ( .A(round_reg[394]), .B(n1808), .Z(n3995) );
  NOR U4681 ( .A(n4142), .B(n3728), .Z(n4257) );
  XOR U4682 ( .A(n4258), .B(n3997), .Z(out[1374]) );
  XOR U4683 ( .A(round_reg[393]), .B(n1811), .Z(n3997) );
  NOR U4684 ( .A(n4144), .B(n3744), .Z(n4258) );
  XOR U4685 ( .A(n4259), .B(n3999), .Z(out[1373]) );
  XOR U4686 ( .A(round_reg[392]), .B(n1814), .Z(n3999) );
  NOR U4687 ( .A(n4146), .B(n3748), .Z(n4259) );
  XOR U4688 ( .A(n4260), .B(n4001), .Z(out[1372]) );
  XOR U4689 ( .A(round_reg[391]), .B(n1817), .Z(n4001) );
  NOR U4690 ( .A(n4148), .B(n3752), .Z(n4260) );
  XOR U4691 ( .A(n4261), .B(n4005), .Z(out[1371]) );
  XOR U4692 ( .A(round_reg[390]), .B(n1828), .Z(n4005) );
  NOR U4693 ( .A(n4150), .B(n3756), .Z(n4261) );
  XOR U4694 ( .A(n4262), .B(n4007), .Z(out[1370]) );
  XOR U4695 ( .A(round_reg[389]), .B(n1831), .Z(n4007) );
  NOR U4696 ( .A(n4152), .B(n3760), .Z(n4262) );
  XOR U4697 ( .A(n4263), .B(n3395), .Z(out[136]) );
  XOR U4698 ( .A(round_reg[673]), .B(n2004), .Z(n3395) );
  ANDN U4699 ( .B(n2046), .A(n1496), .Z(n4263) );
  XNOR U4700 ( .A(round_reg[198]), .B(n2359), .Z(n1496) );
  XNOR U4701 ( .A(round_reg[607]), .B(n2173), .Z(n2046) );
  XOR U4702 ( .A(n4264), .B(n4009), .Z(out[1369]) );
  XOR U4703 ( .A(round_reg[388]), .B(n1834), .Z(n4009) );
  ANDN U4704 ( .B(n3764), .A(n4154), .Z(n4264) );
  XOR U4705 ( .A(n4265), .B(n4011), .Z(out[1368]) );
  XOR U4706 ( .A(round_reg[387]), .B(n1837), .Z(n4011) );
  ANDN U4707 ( .B(n3768), .A(n4156), .Z(n4265) );
  XOR U4708 ( .A(n4266), .B(n4013), .Z(out[1367]) );
  XOR U4709 ( .A(round_reg[386]), .B(n1840), .Z(n4013) );
  ANDN U4710 ( .B(n3773), .A(n4158), .Z(n4266) );
  XOR U4711 ( .A(n4267), .B(n4015), .Z(out[1366]) );
  XOR U4712 ( .A(round_reg[385]), .B(n1843), .Z(n4015) );
  ANDN U4713 ( .B(n3777), .A(n4160), .Z(n4267) );
  XOR U4714 ( .A(n4268), .B(n4017), .Z(out[1365]) );
  XOR U4715 ( .A(round_reg[384]), .B(n1846), .Z(n4017) );
  NOR U4716 ( .A(n4164), .B(n3781), .Z(n4268) );
  XOR U4717 ( .A(n4269), .B(n4019), .Z(out[1364]) );
  XOR U4718 ( .A(round_reg[447]), .B(n1849), .Z(n4019) );
  NOR U4719 ( .A(n4166), .B(n3785), .Z(n4269) );
  XOR U4720 ( .A(n4270), .B(n4021), .Z(out[1363]) );
  XOR U4721 ( .A(round_reg[446]), .B(n1852), .Z(n4021) );
  NOR U4722 ( .A(n4168), .B(n3789), .Z(n4270) );
  XOR U4723 ( .A(n4271), .B(n4023), .Z(out[1362]) );
  XOR U4724 ( .A(round_reg[445]), .B(n1855), .Z(n4023) );
  NOR U4725 ( .A(n4170), .B(n3793), .Z(n4271) );
  XOR U4726 ( .A(n4272), .B(n4027), .Z(out[1361]) );
  XOR U4727 ( .A(round_reg[444]), .B(n1862), .Z(n4027) );
  ANDN U4728 ( .B(n3797), .A(n4172), .Z(n4272) );
  XOR U4729 ( .A(n4273), .B(n4029), .Z(out[1360]) );
  XOR U4730 ( .A(round_reg[443]), .B(n1865), .Z(n4029) );
  NOR U4731 ( .A(n4174), .B(n3801), .Z(n4273) );
  XOR U4732 ( .A(n4274), .B(n3398), .Z(out[135]) );
  XOR U4733 ( .A(round_reg[672]), .B(n2006), .Z(n3398) );
  ANDN U4734 ( .B(n2068), .A(n1820), .Z(n4274) );
  XNOR U4735 ( .A(round_reg[197]), .B(n2363), .Z(n1820) );
  XNOR U4736 ( .A(round_reg[606]), .B(n2177), .Z(n2068) );
  XOR U4737 ( .A(n4275), .B(n4031), .Z(out[1359]) );
  XOR U4738 ( .A(round_reg[442]), .B(n1868), .Z(n4031) );
  NOR U4739 ( .A(n4176), .B(n3804), .Z(n4275) );
  XOR U4740 ( .A(n4276), .B(n4033), .Z(out[1358]) );
  XOR U4741 ( .A(round_reg[441]), .B(n1871), .Z(n4033) );
  NOR U4742 ( .A(n4178), .B(n3822), .Z(n4276) );
  XOR U4743 ( .A(n4277), .B(n4035), .Z(out[1357]) );
  XOR U4744 ( .A(round_reg[440]), .B(n1874), .Z(n4035) );
  NOR U4745 ( .A(n4180), .B(n3827), .Z(n4277) );
  XOR U4746 ( .A(n4278), .B(n4037), .Z(out[1356]) );
  XOR U4747 ( .A(round_reg[439]), .B(n1877), .Z(n4037) );
  ANDN U4748 ( .B(n3831), .A(n4182), .Z(n4278) );
  XOR U4749 ( .A(n4279), .B(n4039), .Z(out[1355]) );
  XOR U4750 ( .A(round_reg[438]), .B(n1880), .Z(n4039) );
  NOR U4751 ( .A(n4185), .B(n3835), .Z(n4279) );
  XOR U4752 ( .A(n4280), .B(n4041), .Z(out[1354]) );
  XOR U4753 ( .A(round_reg[437]), .B(n1883), .Z(n4041) );
  ANDN U4754 ( .B(n3839), .A(n4187), .Z(n4280) );
  XOR U4755 ( .A(n4281), .B(n4043), .Z(out[1353]) );
  XOR U4756 ( .A(round_reg[436]), .B(n1886), .Z(n4043) );
  ANDN U4757 ( .B(n3843), .A(n4189), .Z(n4281) );
  XOR U4758 ( .A(n4282), .B(n4045), .Z(out[1352]) );
  XOR U4759 ( .A(round_reg[435]), .B(n1889), .Z(n4045) );
  ANDN U4760 ( .B(n3847), .A(n4191), .Z(n4282) );
  XOR U4761 ( .A(n4283), .B(n4049), .Z(out[1351]) );
  XOR U4762 ( .A(round_reg[434]), .B(n1896), .Z(n4049) );
  ANDN U4763 ( .B(n3850), .A(n4193), .Z(n4283) );
  XOR U4764 ( .A(n4284), .B(n4051), .Z(out[1350]) );
  XOR U4765 ( .A(round_reg[433]), .B(n1899), .Z(n4051) );
  ANDN U4766 ( .B(n3867), .A(n4195), .Z(n4284) );
  XOR U4767 ( .A(n4285), .B(n3401), .Z(out[134]) );
  XOR U4768 ( .A(round_reg[671]), .B(n2008), .Z(n3401) );
  ANDN U4769 ( .B(n2090), .A(n2091), .Z(n4285) );
  XNOR U4770 ( .A(round_reg[196]), .B(n2367), .Z(n2091) );
  XNOR U4771 ( .A(round_reg[605]), .B(n2181), .Z(n2090) );
  XOR U4772 ( .A(n4286), .B(n4053), .Z(out[1349]) );
  XOR U4773 ( .A(round_reg[432]), .B(n1902), .Z(n4053) );
  ANDN U4774 ( .B(n3871), .A(n4197), .Z(n4286) );
  XOR U4775 ( .A(n4287), .B(n4055), .Z(out[1348]) );
  XOR U4776 ( .A(round_reg[431]), .B(n1905), .Z(n4055) );
  ANDN U4777 ( .B(n3875), .A(n4199), .Z(n4287) );
  XOR U4778 ( .A(n4288), .B(n4057), .Z(out[1347]) );
  XOR U4779 ( .A(round_reg[430]), .B(n1908), .Z(n4057) );
  ANDN U4780 ( .B(n3879), .A(n4201), .Z(n4288) );
  XOR U4781 ( .A(n4289), .B(n4059), .Z(out[1346]) );
  XOR U4782 ( .A(round_reg[429]), .B(n1911), .Z(n4059) );
  ANDN U4783 ( .B(n3897), .A(n4203), .Z(n4289) );
  XOR U4784 ( .A(n4290), .B(n4061), .Z(out[1345]) );
  XNOR U4785 ( .A(round_reg[428]), .B(n1914), .Z(n4061) );
  ANDN U4786 ( .B(n3900), .A(n4207), .Z(n4290) );
  XOR U4787 ( .A(n4291), .B(n4063), .Z(out[1344]) );
  XNOR U4788 ( .A(round_reg[427]), .B(n1917), .Z(n4063) );
  ANDN U4789 ( .B(n3913), .A(n4209), .Z(n4291) );
  XOR U4790 ( .A(n4292), .B(n4065), .Z(out[1343]) );
  XOR U4791 ( .A(round_reg[49]), .B(n1951), .Z(n4065) );
  ANDN U4792 ( .B(n3600), .A(n3586), .Z(n4292) );
  XOR U4793 ( .A(round_reg[1599]), .B(n2313), .Z(n3586) );
  XOR U4794 ( .A(round_reg[1171]), .B(n2299), .Z(n3600) );
  XOR U4795 ( .A(n4293), .B(n4067), .Z(out[1342]) );
  XOR U4796 ( .A(round_reg[48]), .B(n1954), .Z(n4067) );
  NOR U4797 ( .A(n3604), .B(n3602), .Z(n4293) );
  XOR U4798 ( .A(round_reg[1598]), .B(n2317), .Z(n3602) );
  XNOR U4799 ( .A(round_reg[1170]), .B(n2307), .Z(n3604) );
  IV U4800 ( .A(n4294), .Z(n2307) );
  XOR U4801 ( .A(n4295), .B(n4071), .Z(out[1341]) );
  XOR U4802 ( .A(round_reg[47]), .B(n1961), .Z(n4071) );
  NOR U4803 ( .A(n3608), .B(n3606), .Z(n4295) );
  XOR U4804 ( .A(round_reg[1597]), .B(n2321), .Z(n3606) );
  XNOR U4805 ( .A(round_reg[1169]), .B(n2311), .Z(n3608) );
  IV U4806 ( .A(n4296), .Z(n2311) );
  XOR U4807 ( .A(n4297), .B(n4073), .Z(out[1340]) );
  XOR U4808 ( .A(round_reg[46]), .B(n1964), .Z(n4073) );
  NOR U4809 ( .A(n3612), .B(n3610), .Z(n4297) );
  XOR U4810 ( .A(round_reg[1596]), .B(n2325), .Z(n3610) );
  XNOR U4811 ( .A(round_reg[1168]), .B(n2315), .Z(n3612) );
  IV U4812 ( .A(n4298), .Z(n2315) );
  XOR U4813 ( .A(n4299), .B(n3403), .Z(out[133]) );
  XOR U4814 ( .A(round_reg[670]), .B(n2010), .Z(n3403) );
  ANDN U4815 ( .B(n2125), .A(n2126), .Z(n4299) );
  XNOR U4816 ( .A(round_reg[195]), .B(n2371), .Z(n2126) );
  XNOR U4817 ( .A(round_reg[604]), .B(n2185), .Z(n2125) );
  XOR U4818 ( .A(n4300), .B(n4075), .Z(out[1339]) );
  XOR U4819 ( .A(round_reg[45]), .B(n1967), .Z(n4075) );
  NOR U4820 ( .A(n3616), .B(n3614), .Z(n4300) );
  XOR U4821 ( .A(round_reg[1595]), .B(n2329), .Z(n3614) );
  XNOR U4822 ( .A(round_reg[1167]), .B(n2319), .Z(n3616) );
  IV U4823 ( .A(n4301), .Z(n2319) );
  XOR U4824 ( .A(n4302), .B(n4077), .Z(out[1338]) );
  XOR U4825 ( .A(round_reg[44]), .B(n1970), .Z(n4077) );
  NOR U4826 ( .A(n3620), .B(n3618), .Z(n4302) );
  XOR U4827 ( .A(round_reg[1594]), .B(n2333), .Z(n3618) );
  XNOR U4828 ( .A(round_reg[1166]), .B(n2323), .Z(n3620) );
  IV U4829 ( .A(n4303), .Z(n2323) );
  XOR U4830 ( .A(n4304), .B(n4079), .Z(out[1337]) );
  XOR U4831 ( .A(round_reg[43]), .B(n1973), .Z(n4079) );
  IV U4832 ( .A(n4305), .Z(n1973) );
  NOR U4833 ( .A(n3624), .B(n3622), .Z(n4304) );
  XOR U4834 ( .A(round_reg[1593]), .B(n2337), .Z(n3622) );
  XNOR U4835 ( .A(round_reg[1165]), .B(n2327), .Z(n3624) );
  IV U4836 ( .A(n4306), .Z(n2327) );
  XOR U4837 ( .A(n4307), .B(n4081), .Z(out[1336]) );
  XOR U4838 ( .A(round_reg[42]), .B(n1975), .Z(n4081) );
  IV U4839 ( .A(n4308), .Z(n1975) );
  NOR U4840 ( .A(n3628), .B(n3626), .Z(n4307) );
  XOR U4841 ( .A(round_reg[1592]), .B(n2341), .Z(n3626) );
  XNOR U4842 ( .A(round_reg[1164]), .B(n2331), .Z(n3628) );
  IV U4843 ( .A(n4309), .Z(n2331) );
  XOR U4844 ( .A(n4310), .B(n4083), .Z(out[1335]) );
  XOR U4845 ( .A(round_reg[41]), .B(n1977), .Z(n4083) );
  NOR U4846 ( .A(n3632), .B(n3630), .Z(n4310) );
  XOR U4847 ( .A(round_reg[1591]), .B(n2349), .Z(n3630) );
  XNOR U4848 ( .A(round_reg[1163]), .B(n2335), .Z(n3632) );
  IV U4849 ( .A(n4311), .Z(n2335) );
  XOR U4850 ( .A(n4312), .B(n4085), .Z(out[1334]) );
  XOR U4851 ( .A(round_reg[40]), .B(n1980), .Z(n4085) );
  NOR U4852 ( .A(n3636), .B(n3634), .Z(n4312) );
  XOR U4853 ( .A(round_reg[1590]), .B(n2353), .Z(n3634) );
  XNOR U4854 ( .A(round_reg[1162]), .B(n2339), .Z(n3636) );
  XOR U4855 ( .A(n4313), .B(n4087), .Z(out[1333]) );
  XOR U4856 ( .A(round_reg[39]), .B(n1983), .Z(n4087) );
  NOR U4857 ( .A(n3641), .B(n3639), .Z(n4313) );
  XOR U4858 ( .A(round_reg[1589]), .B(n2357), .Z(n3639) );
  XNOR U4859 ( .A(round_reg[1161]), .B(n2343), .Z(n3641) );
  XOR U4860 ( .A(n4314), .B(n4089), .Z(out[1332]) );
  XOR U4861 ( .A(round_reg[38]), .B(n1986), .Z(n4089) );
  NOR U4862 ( .A(n3645), .B(n3643), .Z(n4314) );
  XOR U4863 ( .A(round_reg[1588]), .B(n2361), .Z(n3643) );
  XNOR U4864 ( .A(round_reg[1160]), .B(n2351), .Z(n3645) );
  XOR U4865 ( .A(n4315), .B(n4093), .Z(out[1331]) );
  XOR U4866 ( .A(round_reg[37]), .B(n1993), .Z(n4093) );
  ANDN U4867 ( .B(n3649), .A(n3647), .Z(n4315) );
  XOR U4868 ( .A(round_reg[1587]), .B(n2365), .Z(n3647) );
  XOR U4869 ( .A(round_reg[1159]), .B(n2355), .Z(n3649) );
  XOR U4870 ( .A(n4316), .B(n4095), .Z(out[1330]) );
  XOR U4871 ( .A(round_reg[36]), .B(n1996), .Z(n4095) );
  NOR U4872 ( .A(n3653), .B(n3651), .Z(n4316) );
  XOR U4873 ( .A(round_reg[1586]), .B(n2369), .Z(n3651) );
  XNOR U4874 ( .A(round_reg[1158]), .B(n2359), .Z(n3653) );
  IV U4875 ( .A(n4317), .Z(n2359) );
  XOR U4876 ( .A(n4318), .B(n3405), .Z(out[132]) );
  XOR U4877 ( .A(round_reg[669]), .B(n2012), .Z(n3405) );
  ANDN U4878 ( .B(n2169), .A(n2170), .Z(n4318) );
  XNOR U4879 ( .A(round_reg[194]), .B(n2375), .Z(n2170) );
  XNOR U4880 ( .A(round_reg[603]), .B(n2189), .Z(n2169) );
  XOR U4881 ( .A(n4319), .B(n4097), .Z(out[1329]) );
  XOR U4882 ( .A(round_reg[35]), .B(n1999), .Z(n4097) );
  NOR U4883 ( .A(n3657), .B(n3655), .Z(n4319) );
  XOR U4884 ( .A(round_reg[1585]), .B(n2373), .Z(n3655) );
  XNOR U4885 ( .A(round_reg[1157]), .B(n2363), .Z(n3657) );
  IV U4886 ( .A(n4320), .Z(n2363) );
  XOR U4887 ( .A(n4321), .B(n4099), .Z(out[1328]) );
  XNOR U4888 ( .A(round_reg[34]), .B(n4249), .Z(n4099) );
  NOR U4889 ( .A(n3661), .B(n3659), .Z(n4321) );
  XOR U4890 ( .A(round_reg[1584]), .B(n2377), .Z(n3659) );
  XNOR U4891 ( .A(round_reg[1156]), .B(n2367), .Z(n3661) );
  IV U4892 ( .A(n4322), .Z(n2367) );
  XOR U4893 ( .A(n4323), .B(n4101), .Z(out[1327]) );
  XOR U4894 ( .A(round_reg[33]), .B(n2004), .Z(n4101) );
  IV U4895 ( .A(n4324), .Z(n2004) );
  NOR U4896 ( .A(n3665), .B(n3663), .Z(n4323) );
  XOR U4897 ( .A(round_reg[1583]), .B(n2381), .Z(n3663) );
  XNOR U4898 ( .A(round_reg[1155]), .B(n2371), .Z(n3665) );
  IV U4899 ( .A(n4325), .Z(n2371) );
  XOR U4900 ( .A(n4326), .B(n4103), .Z(out[1326]) );
  XOR U4901 ( .A(round_reg[32]), .B(n2006), .Z(n4103) );
  IV U4902 ( .A(n4327), .Z(n2006) );
  NOR U4903 ( .A(n3669), .B(n3667), .Z(n4326) );
  XOR U4904 ( .A(round_reg[1582]), .B(n2385), .Z(n3667) );
  XNOR U4905 ( .A(round_reg[1154]), .B(n2375), .Z(n3669) );
  IV U4906 ( .A(n4328), .Z(n2375) );
  XOR U4907 ( .A(n4329), .B(n4105), .Z(out[1325]) );
  XOR U4908 ( .A(round_reg[31]), .B(n2008), .Z(n4105) );
  IV U4909 ( .A(n4330), .Z(n2008) );
  NOR U4910 ( .A(n3673), .B(n3671), .Z(n4329) );
  XOR U4911 ( .A(round_reg[1581]), .B(n2106), .Z(n3671) );
  XNOR U4912 ( .A(round_reg[1153]), .B(n2379), .Z(n3673) );
  XOR U4913 ( .A(n4331), .B(n4107), .Z(out[1324]) );
  XOR U4914 ( .A(round_reg[30]), .B(n2010), .Z(n4107) );
  IV U4915 ( .A(n4332), .Z(n2010) );
  NOR U4916 ( .A(n3677), .B(n3675), .Z(n4331) );
  XOR U4917 ( .A(round_reg[1580]), .B(n2110), .Z(n3675) );
  XNOR U4918 ( .A(round_reg[1152]), .B(n2383), .Z(n3677) );
  XOR U4919 ( .A(n4333), .B(n4109), .Z(out[1323]) );
  XOR U4920 ( .A(round_reg[29]), .B(n2012), .Z(n4109) );
  IV U4921 ( .A(n4334), .Z(n2012) );
  NOR U4922 ( .A(n3682), .B(n3680), .Z(n4333) );
  XNOR U4923 ( .A(round_reg[1579]), .B(n4025), .Z(n3680) );
  XNOR U4924 ( .A(round_reg[1215]), .B(n2387), .Z(n3682) );
  XOR U4925 ( .A(n4335), .B(n4111), .Z(out[1322]) );
  XOR U4926 ( .A(round_reg[28]), .B(n2014), .Z(n4111) );
  ANDN U4927 ( .B(n3686), .A(n3684), .Z(n4335) );
  XNOR U4928 ( .A(round_reg[1578]), .B(n4047), .Z(n3684) );
  XNOR U4929 ( .A(round_reg[1214]), .B(n2107), .Z(n3686) );
  XOR U4930 ( .A(n4336), .B(n4115), .Z(out[1321]) );
  XOR U4931 ( .A(round_reg[27]), .B(n2020), .Z(n4115) );
  NOR U4932 ( .A(n3690), .B(n3688), .Z(n4336) );
  XNOR U4933 ( .A(round_reg[1577]), .B(n4069), .Z(n3688) );
  XNOR U4934 ( .A(round_reg[1213]), .B(n2993), .Z(n3690) );
  XOR U4935 ( .A(n4337), .B(n4117), .Z(out[1320]) );
  XOR U4936 ( .A(round_reg[26]), .B(n2022), .Z(n4117) );
  ANDN U4937 ( .B(n3694), .A(n3692), .Z(n4337) );
  XNOR U4938 ( .A(round_reg[1576]), .B(n4091), .Z(n3692) );
  XOR U4939 ( .A(round_reg[1212]), .B(n2115), .Z(n3694) );
  XOR U4940 ( .A(n4338), .B(n3408), .Z(out[131]) );
  XOR U4941 ( .A(round_reg[668]), .B(n2014), .Z(n3408) );
  ANDN U4942 ( .B(n2213), .A(n2214), .Z(n4338) );
  XNOR U4943 ( .A(round_reg[193]), .B(n2379), .Z(n2214) );
  IV U4944 ( .A(n4339), .Z(n2379) );
  XNOR U4945 ( .A(round_reg[602]), .B(n2193), .Z(n2213) );
  XOR U4946 ( .A(n4340), .B(n4119), .Z(out[1319]) );
  XOR U4947 ( .A(round_reg[25]), .B(n2025), .Z(n4119) );
  ANDN U4948 ( .B(n3698), .A(n3696), .Z(n4340) );
  XNOR U4949 ( .A(round_reg[1575]), .B(n4113), .Z(n3696) );
  XOR U4950 ( .A(round_reg[1211]), .B(n2119), .Z(n3698) );
  XOR U4951 ( .A(n4341), .B(n4121), .Z(out[1318]) );
  XOR U4952 ( .A(round_reg[24]), .B(n2028), .Z(n4121) );
  NOR U4953 ( .A(n3702), .B(n3700), .Z(n4341) );
  XNOR U4954 ( .A(round_reg[1574]), .B(n4140), .Z(n3700) );
  XNOR U4955 ( .A(round_reg[1210]), .B(n3000), .Z(n3702) );
  XOR U4956 ( .A(n4342), .B(n4123), .Z(out[1317]) );
  XOR U4957 ( .A(round_reg[23]), .B(n2031), .Z(n4123) );
  NOR U4958 ( .A(n3706), .B(n3704), .Z(n4342) );
  XNOR U4959 ( .A(round_reg[1573]), .B(n4162), .Z(n3704) );
  XNOR U4960 ( .A(round_reg[1209]), .B(n2135), .Z(n3706) );
  XOR U4961 ( .A(n4343), .B(n4126), .Z(out[1316]) );
  XOR U4962 ( .A(round_reg[22]), .B(n2034), .Z(n4126) );
  ANDN U4963 ( .B(n3708), .A(n3710), .Z(n4343) );
  XNOR U4964 ( .A(round_reg[1208]), .B(n2139), .Z(n3710) );
  XNOR U4965 ( .A(round_reg[1572]), .B(n2149), .Z(n3708) );
  IV U4966 ( .A(n4344), .Z(n2149) );
  XOR U4967 ( .A(n4345), .B(n4130), .Z(out[1315]) );
  XOR U4968 ( .A(round_reg[21]), .B(n2037), .Z(n4130) );
  NOR U4969 ( .A(n3714), .B(n3712), .Z(n4345) );
  XNOR U4970 ( .A(round_reg[1571]), .B(n4205), .Z(n3712) );
  XNOR U4971 ( .A(round_reg[1207]), .B(n2143), .Z(n3714) );
  XOR U4972 ( .A(n4346), .B(n4133), .Z(out[1314]) );
  XOR U4973 ( .A(round_reg[20]), .B(n2040), .Z(n4133) );
  NOR U4974 ( .A(n3717), .B(n3716), .Z(n4346) );
  XNOR U4975 ( .A(round_reg[1570]), .B(n4220), .Z(n3716) );
  XNOR U4976 ( .A(round_reg[1206]), .B(n2147), .Z(n3717) );
  XOR U4977 ( .A(n4347), .B(n4136), .Z(out[1313]) );
  XOR U4978 ( .A(round_reg[19]), .B(n2042), .Z(n4136) );
  ANDN U4979 ( .B(n3721), .A(n3722), .Z(n4347) );
  XNOR U4980 ( .A(round_reg[1205]), .B(n2151), .Z(n3722) );
  XNOR U4981 ( .A(round_reg[1569]), .B(n2161), .Z(n3721) );
  IV U4982 ( .A(n4348), .Z(n2161) );
  XOR U4983 ( .A(n4349), .B(n4138), .Z(out[1312]) );
  XOR U4984 ( .A(round_reg[18]), .B(n2044), .Z(n4138) );
  ANDN U4985 ( .B(n3725), .A(n3726), .Z(n4349) );
  XNOR U4986 ( .A(round_reg[1204]), .B(n2155), .Z(n3726) );
  XNOR U4987 ( .A(round_reg[1568]), .B(n2165), .Z(n3725) );
  IV U4988 ( .A(n4350), .Z(n2165) );
  XOR U4989 ( .A(n4351), .B(n4142), .Z(out[1311]) );
  XOR U4990 ( .A(round_reg[17]), .B(n2048), .Z(n4142) );
  ANDN U4991 ( .B(n3728), .A(n3742), .Z(n4351) );
  XNOR U4992 ( .A(round_reg[1203]), .B(n2159), .Z(n3742) );
  XNOR U4993 ( .A(round_reg[1567]), .B(n2173), .Z(n3728) );
  IV U4994 ( .A(n4352), .Z(n2173) );
  XOR U4995 ( .A(n4353), .B(n4144), .Z(out[1310]) );
  XOR U4996 ( .A(round_reg[16]), .B(n2050), .Z(n4144) );
  ANDN U4997 ( .B(n3744), .A(n3746), .Z(n4353) );
  XNOR U4998 ( .A(round_reg[1202]), .B(n2163), .Z(n3746) );
  XNOR U4999 ( .A(round_reg[1566]), .B(n2177), .Z(n3744) );
  IV U5000 ( .A(n4354), .Z(n2177) );
  XOR U5001 ( .A(n4355), .B(n3410), .Z(out[130]) );
  IV U5002 ( .A(n3525), .Z(n3410) );
  XNOR U5003 ( .A(round_reg[667]), .B(n2020), .Z(n3525) );
  ANDN U5004 ( .B(n2257), .A(n2258), .Z(n4355) );
  XNOR U5005 ( .A(round_reg[192]), .B(n2383), .Z(n2258) );
  IV U5006 ( .A(n4356), .Z(n2383) );
  XNOR U5007 ( .A(round_reg[601]), .B(n2197), .Z(n2257) );
  IV U5008 ( .A(n4357), .Z(n2197) );
  XOR U5009 ( .A(n4358), .B(n4146), .Z(out[1309]) );
  XOR U5010 ( .A(round_reg[15]), .B(n2052), .Z(n4146) );
  ANDN U5011 ( .B(n3748), .A(n3750), .Z(n4358) );
  XNOR U5012 ( .A(round_reg[1201]), .B(n2167), .Z(n3750) );
  XNOR U5013 ( .A(round_reg[1565]), .B(n2181), .Z(n3748) );
  IV U5014 ( .A(n4359), .Z(n2181) );
  XOR U5015 ( .A(n4360), .B(n4148), .Z(out[1308]) );
  XOR U5016 ( .A(round_reg[14]), .B(n2054), .Z(n4148) );
  ANDN U5017 ( .B(n3752), .A(n3754), .Z(n4360) );
  XNOR U5018 ( .A(round_reg[1200]), .B(n2175), .Z(n3754) );
  XNOR U5019 ( .A(round_reg[1564]), .B(n2185), .Z(n3752) );
  IV U5020 ( .A(n4361), .Z(n2185) );
  XOR U5021 ( .A(n4362), .B(n4150), .Z(out[1307]) );
  XOR U5022 ( .A(round_reg[13]), .B(n2056), .Z(n4150) );
  ANDN U5023 ( .B(n3756), .A(n3758), .Z(n4362) );
  XNOR U5024 ( .A(round_reg[1199]), .B(n2179), .Z(n3758) );
  XNOR U5025 ( .A(round_reg[1563]), .B(n2189), .Z(n3756) );
  IV U5026 ( .A(n4363), .Z(n2189) );
  XOR U5027 ( .A(n4364), .B(n4152), .Z(out[1306]) );
  XOR U5028 ( .A(round_reg[12]), .B(n2058), .Z(n4152) );
  ANDN U5029 ( .B(n3760), .A(n3762), .Z(n4364) );
  XNOR U5030 ( .A(round_reg[1198]), .B(n2183), .Z(n3762) );
  XNOR U5031 ( .A(round_reg[1562]), .B(n2193), .Z(n3760) );
  IV U5032 ( .A(n4365), .Z(n2193) );
  XOR U5033 ( .A(n4366), .B(n4154), .Z(out[1305]) );
  XOR U5034 ( .A(round_reg[11]), .B(n2060), .Z(n4154) );
  ANDN U5035 ( .B(n3766), .A(n3764), .Z(n4366) );
  XNOR U5036 ( .A(round_reg[1561]), .B(n4357), .Z(n3764) );
  XOR U5037 ( .A(round_reg[1197]), .B(n2187), .Z(n3766) );
  XOR U5038 ( .A(n4367), .B(n4156), .Z(out[1304]) );
  XOR U5039 ( .A(round_reg[10]), .B(n2062), .Z(n4156) );
  ANDN U5040 ( .B(n3770), .A(n3768), .Z(n4367) );
  XNOR U5041 ( .A(round_reg[1560]), .B(n4368), .Z(n3768) );
  XOR U5042 ( .A(round_reg[1196]), .B(n2191), .Z(n3770) );
  XOR U5043 ( .A(n4369), .B(n4158), .Z(out[1303]) );
  XOR U5044 ( .A(round_reg[9]), .B(n2064), .Z(n4158) );
  ANDN U5045 ( .B(n3775), .A(n3773), .Z(n4369) );
  XNOR U5046 ( .A(round_reg[1559]), .B(n4370), .Z(n3773) );
  XOR U5047 ( .A(round_reg[1195]), .B(n2195), .Z(n3775) );
  XOR U5048 ( .A(n4371), .B(n4160), .Z(out[1302]) );
  XOR U5049 ( .A(round_reg[8]), .B(n2066), .Z(n4160) );
  ANDN U5050 ( .B(n3779), .A(n3777), .Z(n4371) );
  XNOR U5051 ( .A(round_reg[1558]), .B(n4372), .Z(n3777) );
  XOR U5052 ( .A(round_reg[1194]), .B(n2199), .Z(n3779) );
  XOR U5053 ( .A(n4373), .B(n4164), .Z(out[1301]) );
  XOR U5054 ( .A(round_reg[7]), .B(n2070), .Z(n4164) );
  AND U5055 ( .A(n3781), .B(n3783), .Z(n4373) );
  XOR U5056 ( .A(round_reg[1193]), .B(n2203), .Z(n3783) );
  XNOR U5057 ( .A(round_reg[1557]), .B(n2217), .Z(n3781) );
  XOR U5058 ( .A(n4374), .B(n4166), .Z(out[1300]) );
  XOR U5059 ( .A(round_reg[6]), .B(n2072), .Z(n4166) );
  AND U5060 ( .A(n3785), .B(n3787), .Z(n4374) );
  XOR U5061 ( .A(round_reg[1192]), .B(n2207), .Z(n3787) );
  XNOR U5062 ( .A(round_reg[1556]), .B(n2221), .Z(n3785) );
  XOR U5063 ( .A(n4375), .B(n1928), .Z(out[12]) );
  XOR U5064 ( .A(round_reg[202]), .B(n2339), .Z(n1928) );
  IV U5065 ( .A(n4376), .Z(n2339) );
  ANDN U5066 ( .B(n3381), .A(n3382), .Z(n4375) );
  XOR U5067 ( .A(round_reg[1045]), .B(n1771), .Z(n3382) );
  XNOR U5068 ( .A(round_reg[1422]), .B(n2298), .Z(n3381) );
  XOR U5069 ( .A(n4377), .B(n3413), .Z(out[129]) );
  XOR U5070 ( .A(round_reg[666]), .B(n2022), .Z(n3413) );
  ANDN U5071 ( .B(n2301), .A(n2302), .Z(n4377) );
  XNOR U5072 ( .A(round_reg[255]), .B(n2387), .Z(n2302) );
  IV U5073 ( .A(n4378), .Z(n2387) );
  XNOR U5074 ( .A(round_reg[600]), .B(n2201), .Z(n2301) );
  IV U5075 ( .A(n4368), .Z(n2201) );
  XOR U5076 ( .A(n4379), .B(n4168), .Z(out[1299]) );
  XOR U5077 ( .A(round_reg[5]), .B(n2074), .Z(n4168) );
  AND U5078 ( .A(n3789), .B(n3791), .Z(n4379) );
  XOR U5079 ( .A(round_reg[1191]), .B(n2211), .Z(n3791) );
  XNOR U5080 ( .A(round_reg[1555]), .B(n2225), .Z(n3789) );
  XOR U5081 ( .A(n4380), .B(n4170), .Z(out[1298]) );
  XOR U5082 ( .A(round_reg[4]), .B(n2076), .Z(n4170) );
  AND U5083 ( .A(n3793), .B(n3795), .Z(n4380) );
  XOR U5084 ( .A(round_reg[1190]), .B(n2219), .Z(n3795) );
  XNOR U5085 ( .A(round_reg[1554]), .B(n2229), .Z(n3793) );
  XOR U5086 ( .A(n4381), .B(n4172), .Z(out[1297]) );
  XOR U5087 ( .A(round_reg[3]), .B(n2078), .Z(n4172) );
  ANDN U5088 ( .B(n3799), .A(n3797), .Z(n4381) );
  XOR U5089 ( .A(round_reg[1553]), .B(n2233), .Z(n3797) );
  XOR U5090 ( .A(round_reg[1189]), .B(n2223), .Z(n3799) );
  XOR U5091 ( .A(n4382), .B(n4174), .Z(out[1296]) );
  XOR U5092 ( .A(round_reg[2]), .B(n2080), .Z(n4174) );
  AND U5093 ( .A(n3801), .B(n3803), .Z(n4382) );
  XOR U5094 ( .A(round_reg[1188]), .B(n2227), .Z(n3803) );
  XNOR U5095 ( .A(round_reg[1552]), .B(n2237), .Z(n3801) );
  XOR U5096 ( .A(n4383), .B(n4176), .Z(out[1295]) );
  XOR U5097 ( .A(round_reg[1]), .B(n2082), .Z(n4176) );
  AND U5098 ( .A(n3804), .B(n3820), .Z(n4383) );
  XOR U5099 ( .A(round_reg[1187]), .B(n2231), .Z(n3820) );
  XNOR U5100 ( .A(round_reg[1551]), .B(n2241), .Z(n3804) );
  XOR U5101 ( .A(n4384), .B(n4178), .Z(out[1294]) );
  XOR U5102 ( .A(round_reg[0]), .B(n2084), .Z(n4178) );
  AND U5103 ( .A(n3822), .B(n3824), .Z(n4384) );
  XOR U5104 ( .A(round_reg[1186]), .B(n2235), .Z(n3824) );
  XNOR U5105 ( .A(round_reg[1550]), .B(n2245), .Z(n3822) );
  XOR U5106 ( .A(n4385), .B(n4180), .Z(out[1293]) );
  XNOR U5107 ( .A(round_reg[63]), .B(n2086), .Z(n4180) );
  AND U5108 ( .A(n3827), .B(n3829), .Z(n4385) );
  XOR U5109 ( .A(round_reg[1185]), .B(n2239), .Z(n3829) );
  XNOR U5110 ( .A(round_reg[1549]), .B(n2249), .Z(n3827) );
  XOR U5111 ( .A(n4386), .B(n4182), .Z(out[1292]) );
  XOR U5112 ( .A(round_reg[62]), .B(n2088), .Z(n4182) );
  ANDN U5113 ( .B(n3833), .A(n3831), .Z(n4386) );
  XNOR U5114 ( .A(round_reg[1548]), .B(n4387), .Z(n3831) );
  XNOR U5115 ( .A(round_reg[1184]), .B(n2243), .Z(n3833) );
  XOR U5116 ( .A(n4388), .B(n4185), .Z(out[1291]) );
  XOR U5117 ( .A(round_reg[61]), .B(n2094), .Z(n4185) );
  AND U5118 ( .A(n3835), .B(n3837), .Z(n4388) );
  XNOR U5119 ( .A(round_reg[1183]), .B(n2247), .Z(n3837) );
  XNOR U5120 ( .A(round_reg[1547]), .B(n2261), .Z(n3835) );
  XOR U5121 ( .A(n4389), .B(n4187), .Z(out[1290]) );
  XOR U5122 ( .A(round_reg[60]), .B(n2096), .Z(n4187) );
  ANDN U5123 ( .B(n3841), .A(n3839), .Z(n4389) );
  XOR U5124 ( .A(round_reg[1546]), .B(n2265), .Z(n3839) );
  XNOR U5125 ( .A(round_reg[1182]), .B(n2251), .Z(n3841) );
  XOR U5126 ( .A(n4390), .B(n3417), .Z(out[128]) );
  XOR U5127 ( .A(round_reg[665]), .B(n2025), .Z(n3417) );
  AND U5128 ( .A(n2345), .B(n2347), .Z(n4390) );
  XNOR U5129 ( .A(round_reg[599]), .B(n2205), .Z(n2345) );
  IV U5130 ( .A(n4370), .Z(n2205) );
  XOR U5131 ( .A(n4391), .B(n4189), .Z(out[1289]) );
  XOR U5132 ( .A(round_reg[59]), .B(n2098), .Z(n4189) );
  ANDN U5133 ( .B(n3845), .A(n3843), .Z(n4391) );
  XOR U5134 ( .A(round_reg[1545]), .B(n2269), .Z(n3843) );
  XNOR U5135 ( .A(round_reg[1181]), .B(n2255), .Z(n3845) );
  XOR U5136 ( .A(n4392), .B(n4191), .Z(out[1288]) );
  XOR U5137 ( .A(round_reg[58]), .B(n2100), .Z(n4191) );
  ANDN U5138 ( .B(n3849), .A(n3847), .Z(n4392) );
  XOR U5139 ( .A(round_reg[1544]), .B(n2273), .Z(n3847) );
  XNOR U5140 ( .A(round_reg[1180]), .B(n2263), .Z(n3849) );
  XOR U5141 ( .A(n4393), .B(n4193), .Z(out[1287]) );
  XOR U5142 ( .A(round_reg[57]), .B(n2102), .Z(n4193) );
  ANDN U5143 ( .B(n3865), .A(n3850), .Z(n4393) );
  XOR U5144 ( .A(round_reg[1543]), .B(n2277), .Z(n3850) );
  XOR U5145 ( .A(round_reg[1179]), .B(n2267), .Z(n3865) );
  XOR U5146 ( .A(n4394), .B(n4195), .Z(out[1286]) );
  XNOR U5147 ( .A(round_reg[56]), .B(n4395), .Z(n4195) );
  ANDN U5148 ( .B(n3869), .A(n3867), .Z(n4394) );
  XOR U5149 ( .A(round_reg[1542]), .B(n2281), .Z(n3867) );
  XOR U5150 ( .A(round_reg[1178]), .B(n2271), .Z(n3869) );
  XOR U5151 ( .A(n4396), .B(n4197), .Z(out[1285]) );
  XNOR U5152 ( .A(round_reg[55]), .B(n4397), .Z(n4197) );
  ANDN U5153 ( .B(n3873), .A(n3871), .Z(n4396) );
  XOR U5154 ( .A(round_reg[1541]), .B(n2285), .Z(n3871) );
  XOR U5155 ( .A(round_reg[1177]), .B(n2275), .Z(n3873) );
  XOR U5156 ( .A(n4398), .B(n4199), .Z(out[1284]) );
  XNOR U5157 ( .A(round_reg[54]), .B(n4399), .Z(n4199) );
  ANDN U5158 ( .B(n3877), .A(n3875), .Z(n4398) );
  XOR U5159 ( .A(round_reg[1540]), .B(n2289), .Z(n3875) );
  XOR U5160 ( .A(round_reg[1176]), .B(n2279), .Z(n3877) );
  XOR U5161 ( .A(n4400), .B(n4201), .Z(out[1283]) );
  XNOR U5162 ( .A(round_reg[53]), .B(n4401), .Z(n4201) );
  ANDN U5163 ( .B(n3895), .A(n3879), .Z(n4400) );
  XOR U5164 ( .A(round_reg[1539]), .B(n2293), .Z(n3879) );
  XOR U5165 ( .A(round_reg[1175]), .B(n2283), .Z(n3895) );
  XOR U5166 ( .A(n4402), .B(n4203), .Z(out[1282]) );
  XOR U5167 ( .A(round_reg[52]), .B(n1942), .Z(n4203) );
  ANDN U5168 ( .B(n3899), .A(n3897), .Z(n4402) );
  XOR U5169 ( .A(round_reg[1538]), .B(n2297), .Z(n3897) );
  XOR U5170 ( .A(round_reg[1174]), .B(n2287), .Z(n3899) );
  XOR U5171 ( .A(n4403), .B(n4207), .Z(out[1281]) );
  XOR U5172 ( .A(round_reg[51]), .B(n1945), .Z(n4207) );
  ANDN U5173 ( .B(n3912), .A(n3900), .Z(n4403) );
  XOR U5174 ( .A(round_reg[1537]), .B(n2305), .Z(n3900) );
  XOR U5175 ( .A(round_reg[1173]), .B(n2291), .Z(n3912) );
  XOR U5176 ( .A(n4404), .B(n4209), .Z(out[1280]) );
  XOR U5177 ( .A(round_reg[50]), .B(n1948), .Z(n4209) );
  ANDN U5178 ( .B(n3924), .A(n3913), .Z(n4404) );
  XOR U5179 ( .A(round_reg[1536]), .B(n2309), .Z(n3913) );
  XOR U5180 ( .A(round_reg[1172]), .B(n2295), .Z(n3924) );
  XOR U5181 ( .A(n4405), .B(n3529), .Z(out[127]) );
  XOR U5182 ( .A(round_reg[598]), .B(n2209), .Z(n3529) );
  IV U5183 ( .A(n4372), .Z(n2209) );
  ANDN U5184 ( .B(n2389), .A(n2390), .Z(n4405) );
  XNOR U5185 ( .A(round_reg[1409]), .B(n2358), .Z(n2390) );
  XNOR U5186 ( .A(round_reg[253]), .B(n2993), .Z(n2389) );
  IV U5187 ( .A(n2111), .Z(n2993) );
  XOR U5188 ( .A(n4406), .B(n4407), .Z(out[1279]) );
  ANDN U5189 ( .B(n4408), .A(n4409), .Z(n4406) );
  XOR U5190 ( .A(n4410), .B(n4411), .Z(out[1278]) );
  ANDN U5191 ( .B(n4412), .A(n4413), .Z(n4410) );
  XOR U5192 ( .A(n4414), .B(n4415), .Z(out[1277]) );
  XOR U5193 ( .A(n4418), .B(n4419), .Z(out[1276]) );
  XOR U5194 ( .A(n4422), .B(n4423), .Z(out[1275]) );
  XOR U5195 ( .A(n4426), .B(n4427), .Z(out[1274]) );
  XOR U5196 ( .A(n4430), .B(n4431), .Z(out[1273]) );
  XOR U5197 ( .A(n4434), .B(n4435), .Z(out[1272]) );
  XOR U5198 ( .A(n4438), .B(n4439), .Z(out[1271]) );
  XOR U5199 ( .A(n4442), .B(n4443), .Z(out[1270]) );
  ANDN U5200 ( .B(n4444), .A(n4445), .Z(n4442) );
  XOR U5201 ( .A(n4446), .B(n3531), .Z(out[126]) );
  XOR U5202 ( .A(round_reg[597]), .B(n2217), .Z(n3531) );
  IV U5203 ( .A(n4447), .Z(n2217) );
  ANDN U5204 ( .B(n2433), .A(n2434), .Z(n4446) );
  XNOR U5205 ( .A(round_reg[1408]), .B(n2362), .Z(n2434) );
  XNOR U5206 ( .A(round_reg[252]), .B(n2115), .Z(n2433) );
  XOR U5207 ( .A(n4448), .B(n4449), .Z(out[1269]) );
  ANDN U5208 ( .B(n4450), .A(n4451), .Z(n4448) );
  XOR U5209 ( .A(n4452), .B(n4453), .Z(out[1268]) );
  ANDN U5210 ( .B(n4454), .A(n4455), .Z(n4452) );
  XOR U5211 ( .A(n4456), .B(n4457), .Z(out[1267]) );
  ANDN U5212 ( .B(n4458), .A(n4459), .Z(n4456) );
  XOR U5213 ( .A(n4460), .B(n4461), .Z(out[1266]) );
  ANDN U5214 ( .B(n4462), .A(n4463), .Z(n4460) );
  XOR U5215 ( .A(n4464), .B(n4465), .Z(out[1265]) );
  ANDN U5216 ( .B(n4466), .A(n4467), .Z(n4464) );
  XOR U5217 ( .A(n4468), .B(n4469), .Z(out[1264]) );
  XOR U5218 ( .A(n4472), .B(n4473), .Z(out[1263]) );
  XOR U5219 ( .A(n4476), .B(n4477), .Z(out[1262]) );
  XOR U5220 ( .A(n4480), .B(n4481), .Z(out[1261]) );
  XOR U5221 ( .A(n4484), .B(n4485), .Z(out[1260]) );
  XOR U5222 ( .A(n4488), .B(n3534), .Z(out[125]) );
  XOR U5223 ( .A(round_reg[596]), .B(n2221), .Z(n3534) );
  IV U5224 ( .A(n4489), .Z(n2221) );
  ANDN U5225 ( .B(n2477), .A(n2478), .Z(n4488) );
  XNOR U5226 ( .A(round_reg[1471]), .B(n2366), .Z(n2478) );
  XNOR U5227 ( .A(round_reg[251]), .B(n2119), .Z(n2477) );
  XOR U5228 ( .A(n4490), .B(n4491), .Z(out[1259]) );
  XOR U5229 ( .A(n4494), .B(n4495), .Z(out[1258]) );
  XOR U5230 ( .A(n4498), .B(n4499), .Z(out[1257]) );
  XOR U5231 ( .A(n4502), .B(n4503), .Z(out[1256]) );
  XOR U5232 ( .A(n4506), .B(n1062), .Z(out[1255]) );
  ANDN U5233 ( .B(n4507), .A(n1061), .Z(n4506) );
  XNOR U5234 ( .A(n4508), .B(n1066), .Z(out[1254]) );
  ANDN U5235 ( .B(n4509), .A(n1065), .Z(n4508) );
  XOR U5236 ( .A(n4510), .B(n1070), .Z(out[1253]) );
  ANDN U5237 ( .B(n4511), .A(n1069), .Z(n4510) );
  XOR U5238 ( .A(n4512), .B(n1074), .Z(out[1252]) );
  ANDN U5239 ( .B(n4513), .A(n1073), .Z(n4512) );
  XOR U5240 ( .A(n4514), .B(n1078), .Z(out[1251]) );
  ANDN U5241 ( .B(n4515), .A(n1077), .Z(n4514) );
  XOR U5242 ( .A(n4516), .B(n1082), .Z(out[1250]) );
  ANDN U5243 ( .B(n4517), .A(n1081), .Z(n4516) );
  XOR U5244 ( .A(n4518), .B(n3536), .Z(out[124]) );
  XOR U5245 ( .A(round_reg[595]), .B(n2225), .Z(n3536) );
  IV U5246 ( .A(n4519), .Z(n2225) );
  ANDN U5247 ( .B(n2521), .A(n2522), .Z(n4518) );
  XNOR U5248 ( .A(round_reg[1470]), .B(n2370), .Z(n2522) );
  XNOR U5249 ( .A(round_reg[250]), .B(n3000), .Z(n2521) );
  IV U5250 ( .A(n2130), .Z(n3000) );
  XOR U5251 ( .A(n4520), .B(n1086), .Z(out[1249]) );
  ANDN U5252 ( .B(n4521), .A(n1085), .Z(n4520) );
  XOR U5253 ( .A(n4522), .B(n1090), .Z(out[1248]) );
  ANDN U5254 ( .B(n4523), .A(n1089), .Z(n4522) );
  XOR U5255 ( .A(n4524), .B(n1094), .Z(out[1247]) );
  ANDN U5256 ( .B(n4525), .A(n1093), .Z(n4524) );
  XOR U5257 ( .A(n4526), .B(n1098), .Z(out[1246]) );
  ANDN U5258 ( .B(n4527), .A(n1097), .Z(n4526) );
  XOR U5259 ( .A(n4528), .B(n1106), .Z(out[1245]) );
  ANDN U5260 ( .B(n4529), .A(n1105), .Z(n4528) );
  XOR U5261 ( .A(n4530), .B(n1110), .Z(out[1244]) );
  ANDN U5262 ( .B(n4531), .A(n1109), .Z(n4530) );
  XOR U5263 ( .A(n4532), .B(n1114), .Z(out[1243]) );
  ANDN U5264 ( .B(n4533), .A(n1113), .Z(n4532) );
  XOR U5265 ( .A(n4534), .B(n1118), .Z(out[1242]) );
  ANDN U5266 ( .B(n4535), .A(n1117), .Z(n4534) );
  XOR U5267 ( .A(n4536), .B(n1122), .Z(out[1241]) );
  ANDN U5268 ( .B(n4537), .A(n1121), .Z(n4536) );
  XOR U5269 ( .A(n4538), .B(n1126), .Z(out[1240]) );
  ANDN U5270 ( .B(n4539), .A(n1125), .Z(n4538) );
  XOR U5271 ( .A(n4540), .B(n3538), .Z(out[123]) );
  XOR U5272 ( .A(round_reg[594]), .B(n2229), .Z(n3538) );
  IV U5273 ( .A(n4541), .Z(n2229) );
  ANDN U5274 ( .B(n2568), .A(n2569), .Z(n4540) );
  XNOR U5275 ( .A(round_reg[1469]), .B(n2374), .Z(n2569) );
  XNOR U5276 ( .A(round_reg[249]), .B(n2135), .Z(n2568) );
  IV U5277 ( .A(n4542), .Z(n2135) );
  XOR U5278 ( .A(n4543), .B(n1130), .Z(out[1239]) );
  ANDN U5279 ( .B(n4544), .A(n1129), .Z(n4543) );
  XOR U5280 ( .A(n4545), .B(n1134), .Z(out[1238]) );
  ANDN U5281 ( .B(n4546), .A(n1133), .Z(n4545) );
  XOR U5282 ( .A(n4547), .B(n1138), .Z(out[1237]) );
  ANDN U5283 ( .B(n4548), .A(n1137), .Z(n4547) );
  XOR U5284 ( .A(n4549), .B(n1142), .Z(out[1236]) );
  ANDN U5285 ( .B(n4550), .A(n1141), .Z(n4549) );
  XOR U5286 ( .A(n4551), .B(n1150), .Z(out[1235]) );
  AND U5287 ( .A(n4552), .B(n1149), .Z(n4551) );
  IV U5288 ( .A(n4553), .Z(n1149) );
  XOR U5289 ( .A(n4554), .B(n1154), .Z(out[1234]) );
  ANDN U5290 ( .B(n4555), .A(n1153), .Z(n4554) );
  XOR U5291 ( .A(n4556), .B(n1158), .Z(out[1233]) );
  ANDN U5292 ( .B(n4557), .A(n1157), .Z(n4556) );
  XOR U5293 ( .A(n4558), .B(n1162), .Z(out[1232]) );
  ANDN U5294 ( .B(n4559), .A(n1161), .Z(n4558) );
  XOR U5295 ( .A(n4560), .B(n1166), .Z(out[1231]) );
  ANDN U5296 ( .B(n4561), .A(n1165), .Z(n4560) );
  XOR U5297 ( .A(n4562), .B(n1170), .Z(out[1230]) );
  ANDN U5298 ( .B(n4563), .A(n1169), .Z(n4562) );
  XOR U5299 ( .A(n4564), .B(n3430), .Z(out[122]) );
  IV U5300 ( .A(n3540), .Z(n3430) );
  XNOR U5301 ( .A(round_reg[593]), .B(n2233), .Z(n3540) );
  ANDN U5302 ( .B(n2612), .A(n2613), .Z(n4564) );
  XNOR U5303 ( .A(round_reg[1468]), .B(n2378), .Z(n2613) );
  XNOR U5304 ( .A(round_reg[248]), .B(n2139), .Z(n2612) );
  IV U5305 ( .A(n4565), .Z(n2139) );
  XOR U5306 ( .A(n4566), .B(n1174), .Z(out[1229]) );
  ANDN U5307 ( .B(n4567), .A(n1173), .Z(n4566) );
  XOR U5308 ( .A(n4568), .B(n1178), .Z(out[1228]) );
  AND U5309 ( .A(n4569), .B(n1177), .Z(n4568) );
  IV U5310 ( .A(n4570), .Z(n1177) );
  XOR U5311 ( .A(n4571), .B(n1182), .Z(out[1227]) );
  AND U5312 ( .A(n4572), .B(n1181), .Z(n4571) );
  IV U5313 ( .A(n4573), .Z(n1181) );
  XOR U5314 ( .A(n4574), .B(n1186), .Z(out[1226]) );
  AND U5315 ( .A(n4575), .B(n1185), .Z(n4574) );
  IV U5316 ( .A(n4576), .Z(n1185) );
  XOR U5317 ( .A(n4577), .B(n1194), .Z(out[1225]) );
  AND U5318 ( .A(n4578), .B(n1193), .Z(n4577) );
  IV U5319 ( .A(n4579), .Z(n1193) );
  XOR U5320 ( .A(n4580), .B(n1198), .Z(out[1224]) );
  ANDN U5321 ( .B(n4581), .A(n1197), .Z(n4580) );
  XOR U5322 ( .A(n4582), .B(n1202), .Z(out[1223]) );
  ANDN U5323 ( .B(n4583), .A(n1201), .Z(n4582) );
  XOR U5324 ( .A(n4584), .B(n1206), .Z(out[1222]) );
  ANDN U5325 ( .B(n4585), .A(n1205), .Z(n4584) );
  XNOR U5326 ( .A(n4586), .B(n1209), .Z(out[1221]) );
  AND U5327 ( .A(n4587), .B(n4588), .Z(n4586) );
  XNOR U5328 ( .A(n4589), .B(n1213), .Z(out[1220]) );
  AND U5329 ( .A(n4590), .B(n4591), .Z(n4589) );
  XOR U5330 ( .A(n4592), .B(n3433), .Z(out[121]) );
  XOR U5331 ( .A(round_reg[592]), .B(n2237), .Z(n3433) );
  IV U5332 ( .A(n4593), .Z(n2237) );
  ANDN U5333 ( .B(n2656), .A(n2657), .Z(n4592) );
  XNOR U5334 ( .A(round_reg[1467]), .B(n2382), .Z(n2657) );
  XNOR U5335 ( .A(round_reg[247]), .B(n2143), .Z(n2656) );
  IV U5336 ( .A(n4594), .Z(n2143) );
  XNOR U5337 ( .A(n4595), .B(n1217), .Z(out[1219]) );
  AND U5338 ( .A(n4596), .B(n4597), .Z(n4595) );
  XNOR U5339 ( .A(n4598), .B(n1221), .Z(out[1218]) );
  AND U5340 ( .A(n4599), .B(n4600), .Z(n4598) );
  XNOR U5341 ( .A(n4601), .B(n1225), .Z(out[1217]) );
  AND U5342 ( .A(n4602), .B(n4603), .Z(n4601) );
  XNOR U5343 ( .A(n4604), .B(n1229), .Z(out[1216]) );
  AND U5344 ( .A(n4605), .B(n4606), .Z(n4604) );
  XOR U5345 ( .A(n4607), .B(n4409), .Z(out[1215]) );
  ANDN U5346 ( .B(n4608), .A(n4408), .Z(n4607) );
  XOR U5347 ( .A(n4609), .B(n4413), .Z(out[1214]) );
  ANDN U5348 ( .B(n4610), .A(n4412), .Z(n4609) );
  XOR U5349 ( .A(n4611), .B(n4417), .Z(out[1213]) );
  ANDN U5350 ( .B(n4612), .A(n4416), .Z(n4611) );
  XOR U5351 ( .A(n4613), .B(n4421), .Z(out[1212]) );
  ANDN U5352 ( .B(n4614), .A(n4420), .Z(n4613) );
  XOR U5353 ( .A(n4615), .B(n4425), .Z(out[1211]) );
  ANDN U5354 ( .B(n4616), .A(n4424), .Z(n4615) );
  XOR U5355 ( .A(n4617), .B(n4429), .Z(out[1210]) );
  ANDN U5356 ( .B(n4618), .A(n4428), .Z(n4617) );
  XOR U5357 ( .A(n4619), .B(n3435), .Z(out[120]) );
  XOR U5358 ( .A(round_reg[591]), .B(n2241), .Z(n3435) );
  IV U5359 ( .A(n4620), .Z(n2241) );
  ANDN U5360 ( .B(n2688), .A(n2689), .Z(n4619) );
  XNOR U5361 ( .A(round_reg[1466]), .B(n2386), .Z(n2689) );
  XNOR U5362 ( .A(round_reg[246]), .B(n2147), .Z(n2688) );
  IV U5363 ( .A(n4621), .Z(n2147) );
  XOR U5364 ( .A(n4622), .B(n4433), .Z(out[1209]) );
  ANDN U5365 ( .B(n4623), .A(n4432), .Z(n4622) );
  XOR U5366 ( .A(n4624), .B(n4437), .Z(out[1208]) );
  ANDN U5367 ( .B(n4625), .A(n4436), .Z(n4624) );
  XOR U5368 ( .A(n4626), .B(n4441), .Z(out[1207]) );
  ANDN U5369 ( .B(n4627), .A(n4440), .Z(n4626) );
  XOR U5370 ( .A(n4628), .B(n4445), .Z(out[1206]) );
  ANDN U5371 ( .B(n4629), .A(n4444), .Z(n4628) );
  XOR U5372 ( .A(n4630), .B(n4451), .Z(out[1205]) );
  ANDN U5373 ( .B(n4631), .A(n4450), .Z(n4630) );
  XOR U5374 ( .A(n4632), .B(n4455), .Z(out[1204]) );
  ANDN U5375 ( .B(n4633), .A(n4454), .Z(n4632) );
  XOR U5376 ( .A(n4634), .B(n4459), .Z(out[1203]) );
  ANDN U5377 ( .B(n4635), .A(n4458), .Z(n4634) );
  XOR U5378 ( .A(n4636), .B(n4463), .Z(out[1202]) );
  ANDN U5379 ( .B(n4637), .A(n4462), .Z(n4636) );
  XOR U5380 ( .A(n4638), .B(n4467), .Z(out[1201]) );
  ANDN U5381 ( .B(n4639), .A(n4466), .Z(n4638) );
  XOR U5382 ( .A(n4640), .B(n4471), .Z(out[1200]) );
  ANDN U5383 ( .B(n4641), .A(n4470), .Z(n4640) );
  XOR U5384 ( .A(n4642), .B(n1959), .Z(out[11]) );
  XOR U5385 ( .A(round_reg[201]), .B(n2343), .Z(n1959) );
  IV U5386 ( .A(n4643), .Z(n2343) );
  ANDN U5387 ( .B(n3385), .A(n3386), .Z(n4642) );
  XOR U5388 ( .A(round_reg[1044]), .B(n1774), .Z(n3386) );
  XNOR U5389 ( .A(round_reg[1421]), .B(n2306), .Z(n3385) );
  XOR U5390 ( .A(n4644), .B(n3437), .Z(out[119]) );
  XOR U5391 ( .A(round_reg[590]), .B(n2245), .Z(n3437) );
  IV U5392 ( .A(n4645), .Z(n2245) );
  ANDN U5393 ( .B(n2720), .A(n2721), .Z(n4644) );
  XNOR U5394 ( .A(round_reg[1465]), .B(n2108), .Z(n2721) );
  IV U5395 ( .A(n4125), .Z(n2108) );
  XNOR U5396 ( .A(round_reg[245]), .B(n2151), .Z(n2720) );
  IV U5397 ( .A(n4646), .Z(n2151) );
  XOR U5398 ( .A(n4647), .B(n4475), .Z(out[1199]) );
  ANDN U5399 ( .B(n4648), .A(n4474), .Z(n4647) );
  XOR U5400 ( .A(n4649), .B(n4479), .Z(out[1198]) );
  ANDN U5401 ( .B(n4650), .A(n4478), .Z(n4649) );
  XOR U5402 ( .A(n4651), .B(n4483), .Z(out[1197]) );
  ANDN U5403 ( .B(n4652), .A(n4482), .Z(n4651) );
  XOR U5404 ( .A(n4653), .B(n4487), .Z(out[1196]) );
  ANDN U5405 ( .B(n4654), .A(n4486), .Z(n4653) );
  XOR U5406 ( .A(n4655), .B(n4493), .Z(out[1195]) );
  ANDN U5407 ( .B(n4656), .A(n4492), .Z(n4655) );
  XOR U5408 ( .A(n4657), .B(n4497), .Z(out[1194]) );
  ANDN U5409 ( .B(n4658), .A(n4496), .Z(n4657) );
  XOR U5410 ( .A(n4659), .B(n4501), .Z(out[1193]) );
  ANDN U5411 ( .B(n4660), .A(n4500), .Z(n4659) );
  XOR U5412 ( .A(n4661), .B(n4505), .Z(out[1192]) );
  ANDN U5413 ( .B(n4662), .A(n4504), .Z(n4661) );
  XOR U5414 ( .A(n4663), .B(n1061), .Z(out[1191]) );
  XOR U5415 ( .A(round_reg[979]), .B(n2042), .Z(n1061) );
  XOR U5416 ( .A(n4664), .B(n4665), .Z(n2042) );
  ANDN U5417 ( .B(n4666), .A(n4507), .Z(n4663) );
  XOR U5418 ( .A(n4667), .B(n1065), .Z(out[1190]) );
  XOR U5419 ( .A(round_reg[978]), .B(n2044), .Z(n1065) );
  XOR U5420 ( .A(n4668), .B(n4669), .Z(n2044) );
  ANDN U5421 ( .B(n4670), .A(n4509), .Z(n4667) );
  XOR U5422 ( .A(n4671), .B(n3439), .Z(out[118]) );
  XOR U5423 ( .A(round_reg[589]), .B(n2249), .Z(n3439) );
  IV U5424 ( .A(n4672), .Z(n2249) );
  ANDN U5425 ( .B(n2749), .A(n2750), .Z(n4671) );
  XNOR U5426 ( .A(round_reg[1464]), .B(n2112), .Z(n2750) );
  IV U5427 ( .A(n4129), .Z(n2112) );
  XNOR U5428 ( .A(round_reg[244]), .B(n2155), .Z(n2749) );
  IV U5429 ( .A(n4673), .Z(n2155) );
  XOR U5430 ( .A(n4674), .B(n1069), .Z(out[1189]) );
  XOR U5431 ( .A(round_reg[977]), .B(n2048), .Z(n1069) );
  XOR U5432 ( .A(n4675), .B(n4676), .Z(n2048) );
  ANDN U5433 ( .B(n4677), .A(n4511), .Z(n4674) );
  XOR U5434 ( .A(n4678), .B(n1073), .Z(out[1188]) );
  XOR U5435 ( .A(round_reg[976]), .B(n2050), .Z(n1073) );
  XOR U5436 ( .A(n4679), .B(n4680), .Z(n2050) );
  ANDN U5437 ( .B(n4681), .A(n4513), .Z(n4678) );
  XOR U5438 ( .A(n4682), .B(n1077), .Z(out[1187]) );
  XOR U5439 ( .A(round_reg[975]), .B(n2052), .Z(n1077) );
  XOR U5440 ( .A(n4683), .B(n4684), .Z(n2052) );
  ANDN U5441 ( .B(n4685), .A(n4515), .Z(n4682) );
  XOR U5442 ( .A(n4686), .B(n1081), .Z(out[1186]) );
  XOR U5443 ( .A(round_reg[974]), .B(n2054), .Z(n1081) );
  XOR U5444 ( .A(n4687), .B(n4688), .Z(n2054) );
  ANDN U5445 ( .B(n4689), .A(n4517), .Z(n4686) );
  XOR U5446 ( .A(n4690), .B(n1085), .Z(out[1185]) );
  XOR U5447 ( .A(round_reg[973]), .B(n2056), .Z(n1085) );
  XNOR U5448 ( .A(n4691), .B(n4692), .Z(n2056) );
  ANDN U5449 ( .B(n4693), .A(n4521), .Z(n4690) );
  XOR U5450 ( .A(n4694), .B(n1089), .Z(out[1184]) );
  XOR U5451 ( .A(round_reg[972]), .B(n2058), .Z(n1089) );
  XNOR U5452 ( .A(n4695), .B(n4696), .Z(n2058) );
  ANDN U5453 ( .B(n4697), .A(n4523), .Z(n4694) );
  XOR U5454 ( .A(n4698), .B(n1093), .Z(out[1183]) );
  XOR U5455 ( .A(round_reg[971]), .B(n2060), .Z(n1093) );
  XNOR U5456 ( .A(n4699), .B(n4700), .Z(n2060) );
  ANDN U5457 ( .B(n4701), .A(n4525), .Z(n4698) );
  XOR U5458 ( .A(n4702), .B(n1097), .Z(out[1182]) );
  XOR U5459 ( .A(round_reg[970]), .B(n2062), .Z(n1097) );
  XNOR U5460 ( .A(n4703), .B(n4704), .Z(n2062) );
  ANDN U5461 ( .B(n4705), .A(n4527), .Z(n4702) );
  XOR U5462 ( .A(n4706), .B(n1105), .Z(out[1181]) );
  XOR U5463 ( .A(round_reg[969]), .B(n2064), .Z(n1105) );
  XNOR U5464 ( .A(n4707), .B(n4708), .Z(n2064) );
  ANDN U5465 ( .B(n4709), .A(n4529), .Z(n4706) );
  XOR U5466 ( .A(n4710), .B(n1109), .Z(out[1180]) );
  XOR U5467 ( .A(round_reg[968]), .B(n2066), .Z(n1109) );
  XOR U5468 ( .A(n4711), .B(n4712), .Z(n2066) );
  ANDN U5469 ( .B(n4713), .A(n4531), .Z(n4710) );
  XOR U5470 ( .A(n4714), .B(n3441), .Z(out[117]) );
  XOR U5471 ( .A(round_reg[588]), .B(n2253), .Z(n3441) );
  IV U5472 ( .A(n4387), .Z(n2253) );
  ANDN U5473 ( .B(n2782), .A(n2783), .Z(n4714) );
  XNOR U5474 ( .A(round_reg[1463]), .B(n2116), .Z(n2783) );
  IV U5475 ( .A(n4715), .Z(n2116) );
  XNOR U5476 ( .A(round_reg[243]), .B(n2159), .Z(n2782) );
  IV U5477 ( .A(n4716), .Z(n2159) );
  XOR U5478 ( .A(n4717), .B(n1113), .Z(out[1179]) );
  XOR U5479 ( .A(round_reg[967]), .B(n2070), .Z(n1113) );
  XNOR U5480 ( .A(n4718), .B(n4719), .Z(n2070) );
  ANDN U5481 ( .B(n4720), .A(n4533), .Z(n4717) );
  XOR U5482 ( .A(n4721), .B(n1117), .Z(out[1178]) );
  XOR U5483 ( .A(round_reg[966]), .B(n2072), .Z(n1117) );
  XNOR U5484 ( .A(n4722), .B(n4723), .Z(n2072) );
  ANDN U5485 ( .B(n4724), .A(n4535), .Z(n4721) );
  XOR U5486 ( .A(n4725), .B(n1121), .Z(out[1177]) );
  XOR U5487 ( .A(round_reg[965]), .B(n2074), .Z(n1121) );
  XNOR U5488 ( .A(n4726), .B(n4727), .Z(n2074) );
  ANDN U5489 ( .B(n4728), .A(n4537), .Z(n4725) );
  XOR U5490 ( .A(n4729), .B(n1125), .Z(out[1176]) );
  XOR U5491 ( .A(round_reg[964]), .B(n2076), .Z(n1125) );
  XNOR U5492 ( .A(n4730), .B(n4731), .Z(n2076) );
  ANDN U5493 ( .B(n4732), .A(n4539), .Z(n4729) );
  XOR U5494 ( .A(n4733), .B(n1129), .Z(out[1175]) );
  XOR U5495 ( .A(round_reg[963]), .B(n2078), .Z(n1129) );
  XNOR U5496 ( .A(n4734), .B(n4735), .Z(n2078) );
  ANDN U5497 ( .B(n4736), .A(n4544), .Z(n4733) );
  XOR U5498 ( .A(n4737), .B(n1133), .Z(out[1174]) );
  XOR U5499 ( .A(round_reg[962]), .B(n2080), .Z(n1133) );
  XNOR U5500 ( .A(n4738), .B(n4739), .Z(n2080) );
  ANDN U5501 ( .B(n4740), .A(n4546), .Z(n4737) );
  XOR U5502 ( .A(n4741), .B(n1137), .Z(out[1173]) );
  XOR U5503 ( .A(round_reg[961]), .B(n2082), .Z(n1137) );
  XNOR U5504 ( .A(n4742), .B(n4743), .Z(n2082) );
  ANDN U5505 ( .B(n4744), .A(n4548), .Z(n4741) );
  XOR U5506 ( .A(n4745), .B(n1141), .Z(out[1172]) );
  XOR U5507 ( .A(round_reg[960]), .B(n2084), .Z(n1141) );
  XNOR U5508 ( .A(n4746), .B(n4747), .Z(n2084) );
  ANDN U5509 ( .B(n4748), .A(n4550), .Z(n4745) );
  XOR U5510 ( .A(n4749), .B(n4553), .Z(out[1171]) );
  XNOR U5511 ( .A(round_reg[1023]), .B(n2086), .Z(n4553) );
  ANDN U5512 ( .B(n4752), .A(n4552), .Z(n4749) );
  XOR U5513 ( .A(n4753), .B(n1153), .Z(out[1170]) );
  XOR U5514 ( .A(round_reg[1022]), .B(n2088), .Z(n1153) );
  XNOR U5515 ( .A(n4754), .B(n4755), .Z(n2088) );
  ANDN U5516 ( .B(n4756), .A(n4555), .Z(n4753) );
  XOR U5517 ( .A(n4757), .B(n3443), .Z(out[116]) );
  XOR U5518 ( .A(round_reg[587]), .B(n2261), .Z(n3443) );
  IV U5519 ( .A(n4758), .Z(n2261) );
  ANDN U5520 ( .B(n2806), .A(n2807), .Z(n4757) );
  XNOR U5521 ( .A(round_reg[1462]), .B(n2120), .Z(n2807) );
  IV U5522 ( .A(n4759), .Z(n2120) );
  XNOR U5523 ( .A(round_reg[242]), .B(n2163), .Z(n2806) );
  IV U5524 ( .A(n4760), .Z(n2163) );
  XOR U5525 ( .A(n4761), .B(n1157), .Z(out[1169]) );
  XOR U5526 ( .A(round_reg[1021]), .B(n2094), .Z(n1157) );
  XNOR U5527 ( .A(n4762), .B(n4763), .Z(n2094) );
  ANDN U5528 ( .B(n4764), .A(n4557), .Z(n4761) );
  XOR U5529 ( .A(n4765), .B(n1161), .Z(out[1168]) );
  XOR U5530 ( .A(round_reg[1020]), .B(n2096), .Z(n1161) );
  XNOR U5531 ( .A(n4766), .B(n4767), .Z(n2096) );
  ANDN U5532 ( .B(n4768), .A(n4559), .Z(n4765) );
  XOR U5533 ( .A(n4769), .B(n1165), .Z(out[1167]) );
  XOR U5534 ( .A(round_reg[1019]), .B(n2098), .Z(n1165) );
  XNOR U5535 ( .A(n4770), .B(n4771), .Z(n2098) );
  ANDN U5536 ( .B(n4772), .A(n4561), .Z(n4769) );
  XOR U5537 ( .A(n4773), .B(n1169), .Z(out[1166]) );
  XOR U5538 ( .A(round_reg[1018]), .B(n2100), .Z(n1169) );
  XNOR U5539 ( .A(n4774), .B(n4775), .Z(n2100) );
  ANDN U5540 ( .B(n4776), .A(n4563), .Z(n4773) );
  XOR U5541 ( .A(n4777), .B(n1173), .Z(out[1165]) );
  XOR U5542 ( .A(round_reg[1017]), .B(n2102), .Z(n1173) );
  XNOR U5543 ( .A(n4778), .B(n4779), .Z(n2102) );
  ANDN U5544 ( .B(n4780), .A(n4567), .Z(n4777) );
  XOR U5545 ( .A(n4781), .B(n4570), .Z(out[1164]) );
  XOR U5546 ( .A(round_reg[1016]), .B(n2104), .Z(n4570) );
  IV U5547 ( .A(n4395), .Z(n2104) );
  ANDN U5548 ( .B(n4784), .A(n4569), .Z(n4781) );
  XOR U5549 ( .A(n4785), .B(n4573), .Z(out[1163]) );
  XOR U5550 ( .A(round_reg[1015]), .B(n1936), .Z(n4573) );
  IV U5551 ( .A(n4397), .Z(n1936) );
  ANDN U5552 ( .B(n4788), .A(n4572), .Z(n4785) );
  XOR U5553 ( .A(n4789), .B(n4576), .Z(out[1162]) );
  XOR U5554 ( .A(round_reg[1014]), .B(n1938), .Z(n4576) );
  IV U5555 ( .A(n4399), .Z(n1938) );
  ANDN U5556 ( .B(n4792), .A(n4575), .Z(n4789) );
  XOR U5557 ( .A(n4793), .B(n4579), .Z(out[1161]) );
  XOR U5558 ( .A(round_reg[1013]), .B(n1940), .Z(n4579) );
  IV U5559 ( .A(n4401), .Z(n1940) );
  ANDN U5560 ( .B(n4796), .A(n4578), .Z(n4793) );
  XOR U5561 ( .A(n4797), .B(n1197), .Z(out[1160]) );
  XOR U5562 ( .A(round_reg[1012]), .B(n1942), .Z(n1197) );
  XNOR U5563 ( .A(n4798), .B(n4799), .Z(n1942) );
  ANDN U5564 ( .B(n4800), .A(n4581), .Z(n4797) );
  XOR U5565 ( .A(n4801), .B(n3445), .Z(out[115]) );
  IV U5566 ( .A(n3549), .Z(n3445) );
  XNOR U5567 ( .A(round_reg[586]), .B(n2265), .Z(n3549) );
  ANDN U5568 ( .B(n2831), .A(n2832), .Z(n4801) );
  XNOR U5569 ( .A(round_reg[1461]), .B(n2131), .Z(n2832) );
  IV U5570 ( .A(n4802), .Z(n2131) );
  XNOR U5571 ( .A(round_reg[241]), .B(n2167), .Z(n2831) );
  IV U5572 ( .A(n4803), .Z(n2167) );
  XOR U5573 ( .A(n4804), .B(n1201), .Z(out[1159]) );
  XOR U5574 ( .A(round_reg[1011]), .B(n1945), .Z(n1201) );
  XNOR U5575 ( .A(n4805), .B(n4806), .Z(n1945) );
  ANDN U5576 ( .B(n4807), .A(n4583), .Z(n4804) );
  XOR U5577 ( .A(n4808), .B(n1205), .Z(out[1158]) );
  XOR U5578 ( .A(round_reg[1010]), .B(n1948), .Z(n1205) );
  XNOR U5579 ( .A(n4809), .B(n4810), .Z(n1948) );
  ANDN U5580 ( .B(n4811), .A(n4585), .Z(n4808) );
  XOR U5581 ( .A(n4812), .B(n1210), .Z(out[1157]) );
  IV U5582 ( .A(n4588), .Z(n1210) );
  XNOR U5583 ( .A(round_reg[1009]), .B(n1951), .Z(n4588) );
  XNOR U5584 ( .A(n4813), .B(n4814), .Z(n1951) );
  ANDN U5585 ( .B(n4815), .A(n4587), .Z(n4812) );
  XOR U5586 ( .A(n4816), .B(n1214), .Z(out[1156]) );
  IV U5587 ( .A(n4591), .Z(n1214) );
  XNOR U5588 ( .A(round_reg[1008]), .B(n1954), .Z(n4591) );
  XNOR U5589 ( .A(n4817), .B(n4818), .Z(n1954) );
  ANDN U5590 ( .B(n4819), .A(n4590), .Z(n4816) );
  XOR U5591 ( .A(n4820), .B(n1218), .Z(out[1155]) );
  IV U5592 ( .A(n4597), .Z(n1218) );
  XNOR U5593 ( .A(round_reg[1007]), .B(n1961), .Z(n4597) );
  XNOR U5594 ( .A(n4821), .B(n4822), .Z(n1961) );
  ANDN U5595 ( .B(n4823), .A(n4596), .Z(n4820) );
  XOR U5596 ( .A(n4824), .B(n1222), .Z(out[1154]) );
  IV U5597 ( .A(n4600), .Z(n1222) );
  XNOR U5598 ( .A(round_reg[1006]), .B(n1964), .Z(n4600) );
  XNOR U5599 ( .A(n4825), .B(n4826), .Z(n1964) );
  ANDN U5600 ( .B(n4827), .A(n4599), .Z(n4824) );
  XOR U5601 ( .A(n4828), .B(n1226), .Z(out[1153]) );
  IV U5602 ( .A(n4603), .Z(n1226) );
  XNOR U5603 ( .A(round_reg[1005]), .B(n1967), .Z(n4603) );
  XNOR U5604 ( .A(n4829), .B(n4830), .Z(n1967) );
  ANDN U5605 ( .B(n4831), .A(n4602), .Z(n4828) );
  XOR U5606 ( .A(n4832), .B(n1230), .Z(out[1152]) );
  IV U5607 ( .A(n4606), .Z(n1230) );
  XNOR U5608 ( .A(round_reg[1004]), .B(n1970), .Z(n4606) );
  XNOR U5609 ( .A(n4833), .B(n4834), .Z(n1970) );
  ANDN U5610 ( .B(n4835), .A(n4605), .Z(n4832) );
  XOR U5611 ( .A(n4836), .B(n4408), .Z(out[1151]) );
  XOR U5612 ( .A(round_reg[956]), .B(n2325), .Z(n4408) );
  ANDN U5613 ( .B(n4837), .A(n4608), .Z(n4836) );
  XOR U5614 ( .A(n4838), .B(n4412), .Z(out[1150]) );
  XOR U5615 ( .A(round_reg[955]), .B(n2329), .Z(n4412) );
  ANDN U5616 ( .B(n4839), .A(n4610), .Z(n4838) );
  XOR U5617 ( .A(n4840), .B(n3447), .Z(out[114]) );
  IV U5618 ( .A(n3551), .Z(n3447) );
  XNOR U5619 ( .A(round_reg[585]), .B(n2269), .Z(n3551) );
  ANDN U5620 ( .B(n2857), .A(n2858), .Z(n4840) );
  XNOR U5621 ( .A(round_reg[1460]), .B(n2134), .Z(n2858) );
  XNOR U5622 ( .A(round_reg[240]), .B(n2175), .Z(n2857) );
  IV U5623 ( .A(n4841), .Z(n2175) );
  XOR U5624 ( .A(n4842), .B(n4416), .Z(out[1149]) );
  XOR U5625 ( .A(round_reg[954]), .B(n2333), .Z(n4416) );
  XOR U5626 ( .A(n4843), .B(n4844), .Z(n2333) );
  ANDN U5627 ( .B(n4845), .A(n4612), .Z(n4842) );
  XOR U5628 ( .A(n4846), .B(n4420), .Z(out[1148]) );
  XOR U5629 ( .A(round_reg[953]), .B(n2337), .Z(n4420) );
  XOR U5630 ( .A(n4847), .B(n4848), .Z(n2337) );
  ANDN U5631 ( .B(n4849), .A(n4614), .Z(n4846) );
  XOR U5632 ( .A(n4850), .B(n4424), .Z(out[1147]) );
  XOR U5633 ( .A(round_reg[952]), .B(n2341), .Z(n4424) );
  XOR U5634 ( .A(n4851), .B(n4852), .Z(n2341) );
  ANDN U5635 ( .B(n4853), .A(n4616), .Z(n4850) );
  XOR U5636 ( .A(n4854), .B(n4428), .Z(out[1146]) );
  XOR U5637 ( .A(round_reg[951]), .B(n2349), .Z(n4428) );
  XOR U5638 ( .A(n4855), .B(n4856), .Z(n2349) );
  ANDN U5639 ( .B(n4857), .A(n4618), .Z(n4854) );
  XOR U5640 ( .A(n4858), .B(n4432), .Z(out[1145]) );
  XOR U5641 ( .A(round_reg[950]), .B(n2353), .Z(n4432) );
  XNOR U5642 ( .A(n4859), .B(n4860), .Z(n2353) );
  ANDN U5643 ( .B(n4861), .A(n4623), .Z(n4858) );
  XOR U5644 ( .A(n4862), .B(n4436), .Z(out[1144]) );
  XOR U5645 ( .A(round_reg[949]), .B(n2357), .Z(n4436) );
  XNOR U5646 ( .A(n4863), .B(n4864), .Z(n2357) );
  ANDN U5647 ( .B(n4865), .A(n4625), .Z(n4862) );
  XOR U5648 ( .A(n4866), .B(n4440), .Z(out[1143]) );
  XOR U5649 ( .A(round_reg[948]), .B(n2361), .Z(n4440) );
  XNOR U5650 ( .A(n4867), .B(n4868), .Z(n2361) );
  ANDN U5651 ( .B(n4869), .A(n4627), .Z(n4866) );
  XOR U5652 ( .A(n4870), .B(n4444), .Z(out[1142]) );
  XOR U5653 ( .A(round_reg[947]), .B(n2365), .Z(n4444) );
  XNOR U5654 ( .A(n4871), .B(n4872), .Z(n2365) );
  ANDN U5655 ( .B(n4873), .A(n4629), .Z(n4870) );
  XOR U5656 ( .A(n4874), .B(n4450), .Z(out[1141]) );
  XOR U5657 ( .A(round_reg[946]), .B(n2369), .Z(n4450) );
  XNOR U5658 ( .A(n4875), .B(n4876), .Z(n2369) );
  ANDN U5659 ( .B(n4877), .A(n4631), .Z(n4874) );
  XOR U5660 ( .A(n4878), .B(n4454), .Z(out[1140]) );
  XOR U5661 ( .A(round_reg[945]), .B(n2373), .Z(n4454) );
  XNOR U5662 ( .A(n4879), .B(n4880), .Z(n2373) );
  ANDN U5663 ( .B(n4881), .A(n4633), .Z(n4878) );
  XOR U5664 ( .A(n4882), .B(n3449), .Z(out[113]) );
  IV U5665 ( .A(n3553), .Z(n3449) );
  XNOR U5666 ( .A(round_reg[584]), .B(n2273), .Z(n3553) );
  ANDN U5667 ( .B(n2884), .A(n2885), .Z(n4882) );
  XNOR U5668 ( .A(round_reg[1459]), .B(n2138), .Z(n2885) );
  XNOR U5669 ( .A(round_reg[239]), .B(n2179), .Z(n2884) );
  IV U5670 ( .A(n4883), .Z(n2179) );
  XOR U5671 ( .A(n4884), .B(n4458), .Z(out[1139]) );
  XOR U5672 ( .A(round_reg[944]), .B(n2377), .Z(n4458) );
  XNOR U5673 ( .A(n4885), .B(n4886), .Z(n2377) );
  ANDN U5674 ( .B(n4887), .A(n4635), .Z(n4884) );
  XOR U5675 ( .A(n4888), .B(n4462), .Z(out[1138]) );
  XOR U5676 ( .A(round_reg[943]), .B(n2381), .Z(n4462) );
  XNOR U5677 ( .A(n4889), .B(n4890), .Z(n2381) );
  ANDN U5678 ( .B(n4891), .A(n4637), .Z(n4888) );
  XOR U5679 ( .A(n4892), .B(n4466), .Z(out[1137]) );
  XOR U5680 ( .A(round_reg[942]), .B(n2385), .Z(n4466) );
  XNOR U5681 ( .A(n4893), .B(n4894), .Z(n2385) );
  ANDN U5682 ( .B(n4895), .A(n4639), .Z(n4892) );
  XOR U5683 ( .A(n4896), .B(n4470), .Z(out[1136]) );
  XOR U5684 ( .A(round_reg[941]), .B(n2106), .Z(n4470) );
  XNOR U5685 ( .A(n4897), .B(n4898), .Z(n2106) );
  ANDN U5686 ( .B(n4899), .A(n4641), .Z(n4896) );
  XOR U5687 ( .A(n4900), .B(n4474), .Z(out[1135]) );
  XOR U5688 ( .A(round_reg[940]), .B(n2110), .Z(n4474) );
  XNOR U5689 ( .A(n4901), .B(n4902), .Z(n2110) );
  ANDN U5690 ( .B(n4903), .A(n4648), .Z(n4900) );
  XOR U5691 ( .A(n4904), .B(n4478), .Z(out[1134]) );
  XNOR U5692 ( .A(round_reg[939]), .B(n4025), .Z(n4478) );
  XOR U5693 ( .A(n4905), .B(n4906), .Z(n4025) );
  ANDN U5694 ( .B(n4907), .A(n4650), .Z(n4904) );
  XOR U5695 ( .A(n4908), .B(n4482), .Z(out[1133]) );
  XNOR U5696 ( .A(round_reg[938]), .B(n4047), .Z(n4482) );
  XOR U5697 ( .A(n4909), .B(n4910), .Z(n4047) );
  ANDN U5698 ( .B(n4911), .A(n4652), .Z(n4908) );
  XOR U5699 ( .A(n4912), .B(n4486), .Z(out[1132]) );
  XNOR U5700 ( .A(round_reg[937]), .B(n4069), .Z(n4486) );
  XOR U5701 ( .A(n4913), .B(n4914), .Z(n4069) );
  ANDN U5702 ( .B(n4915), .A(n4654), .Z(n4912) );
  XOR U5703 ( .A(n4916), .B(n4492), .Z(out[1131]) );
  XNOR U5704 ( .A(round_reg[936]), .B(n4091), .Z(n4492) );
  XOR U5705 ( .A(n4917), .B(n4918), .Z(n4091) );
  ANDN U5706 ( .B(n4919), .A(n4656), .Z(n4916) );
  XOR U5707 ( .A(n4920), .B(n4496), .Z(out[1130]) );
  XNOR U5708 ( .A(round_reg[935]), .B(n4113), .Z(n4496) );
  XOR U5709 ( .A(n4921), .B(n4922), .Z(n4113) );
  ANDN U5710 ( .B(n4923), .A(n4658), .Z(n4920) );
  XOR U5711 ( .A(n4924), .B(n3451), .Z(out[112]) );
  IV U5712 ( .A(n3555), .Z(n3451) );
  XNOR U5713 ( .A(round_reg[583]), .B(n2277), .Z(n3555) );
  ANDN U5714 ( .B(n2908), .A(n2910), .Z(n4924) );
  XNOR U5715 ( .A(round_reg[1458]), .B(n2142), .Z(n2910) );
  XNOR U5716 ( .A(round_reg[238]), .B(n2183), .Z(n2908) );
  IV U5717 ( .A(n4925), .Z(n2183) );
  XOR U5718 ( .A(n4926), .B(n4500), .Z(out[1129]) );
  XNOR U5719 ( .A(round_reg[934]), .B(n4140), .Z(n4500) );
  XOR U5720 ( .A(n4927), .B(n4928), .Z(n4140) );
  ANDN U5721 ( .B(n4929), .A(n4660), .Z(n4926) );
  XOR U5722 ( .A(n4930), .B(n4504), .Z(out[1128]) );
  XNOR U5723 ( .A(round_reg[933]), .B(n4162), .Z(n4504) );
  XOR U5724 ( .A(n4931), .B(n4932), .Z(n4162) );
  ANDN U5725 ( .B(n4933), .A(n4662), .Z(n4930) );
  XOR U5726 ( .A(n4934), .B(n4507), .Z(out[1127]) );
  XNOR U5727 ( .A(round_reg[932]), .B(n4344), .Z(n4507) );
  XOR U5728 ( .A(n4935), .B(n4936), .Z(n4344) );
  ANDN U5729 ( .B(n1060), .A(n4666), .Z(n4934) );
  XOR U5730 ( .A(n4937), .B(n4509), .Z(out[1126]) );
  XNOR U5731 ( .A(round_reg[931]), .B(n4205), .Z(n4509) );
  XOR U5732 ( .A(n4938), .B(n4939), .Z(n4205) );
  ANDN U5733 ( .B(n1064), .A(n4670), .Z(n4937) );
  XOR U5734 ( .A(n4940), .B(n4511), .Z(out[1125]) );
  XNOR U5735 ( .A(round_reg[930]), .B(n4220), .Z(n4511) );
  XOR U5736 ( .A(n4941), .B(n4942), .Z(n4220) );
  ANDN U5737 ( .B(n1068), .A(n4677), .Z(n4940) );
  XOR U5738 ( .A(n4943), .B(n4513), .Z(out[1124]) );
  XNOR U5739 ( .A(round_reg[929]), .B(n4348), .Z(n4513) );
  XOR U5740 ( .A(n4944), .B(n4945), .Z(n4348) );
  ANDN U5741 ( .B(n1072), .A(n4681), .Z(n4943) );
  XOR U5742 ( .A(n4946), .B(n4515), .Z(out[1123]) );
  XNOR U5743 ( .A(round_reg[928]), .B(n4350), .Z(n4515) );
  XOR U5744 ( .A(n4947), .B(n4948), .Z(n4350) );
  ANDN U5745 ( .B(n1076), .A(n4685), .Z(n4946) );
  XOR U5746 ( .A(n4949), .B(n4517), .Z(out[1122]) );
  XNOR U5747 ( .A(round_reg[927]), .B(n4352), .Z(n4517) );
  XOR U5748 ( .A(n4950), .B(n4951), .Z(n4352) );
  ANDN U5749 ( .B(n1080), .A(n4689), .Z(n4949) );
  XOR U5750 ( .A(n4952), .B(n4521), .Z(out[1121]) );
  XNOR U5751 ( .A(round_reg[926]), .B(n4354), .Z(n4521) );
  XOR U5752 ( .A(n4953), .B(n4954), .Z(n4354) );
  ANDN U5753 ( .B(n1084), .A(n4693), .Z(n4952) );
  XOR U5754 ( .A(n4955), .B(n4523), .Z(out[1120]) );
  XNOR U5755 ( .A(round_reg[925]), .B(n4359), .Z(n4523) );
  XOR U5756 ( .A(n4956), .B(n4957), .Z(n4359) );
  ANDN U5757 ( .B(n1088), .A(n4697), .Z(n4955) );
  XOR U5758 ( .A(n4958), .B(n3454), .Z(out[111]) );
  XOR U5759 ( .A(round_reg[582]), .B(n2281), .Z(n3454) );
  ANDN U5760 ( .B(n2932), .A(n2934), .Z(n4958) );
  XNOR U5761 ( .A(round_reg[1457]), .B(n2146), .Z(n2934) );
  XNOR U5762 ( .A(round_reg[237]), .B(n2187), .Z(n2932) );
  XOR U5763 ( .A(n4959), .B(n4525), .Z(out[1119]) );
  XNOR U5764 ( .A(round_reg[924]), .B(n4361), .Z(n4525) );
  XOR U5765 ( .A(n4960), .B(n4961), .Z(n4361) );
  ANDN U5766 ( .B(n1092), .A(n4701), .Z(n4959) );
  XOR U5767 ( .A(n4962), .B(n4527), .Z(out[1118]) );
  XNOR U5768 ( .A(round_reg[923]), .B(n4363), .Z(n4527) );
  XOR U5769 ( .A(n4963), .B(n4964), .Z(n4363) );
  ANDN U5770 ( .B(n1096), .A(n4705), .Z(n4962) );
  XOR U5771 ( .A(n4965), .B(n4529), .Z(out[1117]) );
  XNOR U5772 ( .A(round_reg[922]), .B(n4365), .Z(n4529) );
  XOR U5773 ( .A(n4966), .B(n4967), .Z(n4365) );
  NOR U5774 ( .A(n1104), .B(n4709), .Z(n4965) );
  XOR U5775 ( .A(n4968), .B(n4531), .Z(out[1116]) );
  XNOR U5776 ( .A(round_reg[921]), .B(n4357), .Z(n4531) );
  XOR U5777 ( .A(n4969), .B(n4970), .Z(n4357) );
  NOR U5778 ( .A(n1108), .B(n4713), .Z(n4968) );
  XOR U5779 ( .A(n4971), .B(n4533), .Z(out[1115]) );
  XNOR U5780 ( .A(round_reg[920]), .B(n4368), .Z(n4533) );
  XOR U5781 ( .A(n4972), .B(n4973), .Z(n4368) );
  ANDN U5782 ( .B(n1112), .A(n4720), .Z(n4971) );
  XOR U5783 ( .A(n4974), .B(n4535), .Z(out[1114]) );
  XNOR U5784 ( .A(round_reg[919]), .B(n4370), .Z(n4535) );
  XOR U5785 ( .A(n4975), .B(n4976), .Z(n4370) );
  ANDN U5786 ( .B(n1116), .A(n4724), .Z(n4974) );
  XOR U5787 ( .A(n4977), .B(n4537), .Z(out[1113]) );
  XNOR U5788 ( .A(round_reg[918]), .B(n4372), .Z(n4537) );
  XOR U5789 ( .A(n4978), .B(n4979), .Z(n4372) );
  ANDN U5790 ( .B(n1120), .A(n4728), .Z(n4977) );
  XOR U5791 ( .A(n4980), .B(n4539), .Z(out[1112]) );
  XNOR U5792 ( .A(round_reg[917]), .B(n4447), .Z(n4539) );
  XOR U5793 ( .A(n4981), .B(n4982), .Z(n4447) );
  ANDN U5794 ( .B(n1124), .A(n4732), .Z(n4980) );
  XOR U5795 ( .A(n4983), .B(n4544), .Z(out[1111]) );
  XNOR U5796 ( .A(round_reg[916]), .B(n4489), .Z(n4544) );
  XOR U5797 ( .A(n4984), .B(n4985), .Z(n4489) );
  ANDN U5798 ( .B(n1128), .A(n4736), .Z(n4983) );
  XOR U5799 ( .A(n4986), .B(n4546), .Z(out[1110]) );
  XNOR U5800 ( .A(round_reg[915]), .B(n4519), .Z(n4546) );
  XOR U5801 ( .A(n4987), .B(n4988), .Z(n4519) );
  ANDN U5802 ( .B(n1132), .A(n4740), .Z(n4986) );
  XOR U5803 ( .A(n4989), .B(n3457), .Z(out[110]) );
  IV U5804 ( .A(n3558), .Z(n3457) );
  XNOR U5805 ( .A(round_reg[581]), .B(n2285), .Z(n3558) );
  ANDN U5806 ( .B(n2956), .A(n2958), .Z(n4989) );
  XNOR U5807 ( .A(round_reg[1456]), .B(n2150), .Z(n2958) );
  XNOR U5808 ( .A(round_reg[236]), .B(n2191), .Z(n2956) );
  XOR U5809 ( .A(n4990), .B(n4548), .Z(out[1109]) );
  XNOR U5810 ( .A(round_reg[914]), .B(n4541), .Z(n4548) );
  XOR U5811 ( .A(n4991), .B(n4992), .Z(n4541) );
  ANDN U5812 ( .B(n1136), .A(n4744), .Z(n4990) );
  XOR U5813 ( .A(n4993), .B(n4550), .Z(out[1108]) );
  XOR U5814 ( .A(round_reg[913]), .B(n2233), .Z(n4550) );
  XNOR U5815 ( .A(n4994), .B(n4995), .Z(n2233) );
  ANDN U5816 ( .B(n1140), .A(n4748), .Z(n4993) );
  XOR U5817 ( .A(n4996), .B(n4552), .Z(out[1107]) );
  XNOR U5818 ( .A(round_reg[912]), .B(n4593), .Z(n4552) );
  XOR U5819 ( .A(n4997), .B(n4998), .Z(n4593) );
  ANDN U5820 ( .B(n1148), .A(n4752), .Z(n4996) );
  XOR U5821 ( .A(n4999), .B(n4555), .Z(out[1106]) );
  XNOR U5822 ( .A(round_reg[911]), .B(n4620), .Z(n4555) );
  XOR U5823 ( .A(n5000), .B(n5001), .Z(n4620) );
  ANDN U5824 ( .B(n1152), .A(n4756), .Z(n4999) );
  XOR U5825 ( .A(n5002), .B(n4557), .Z(out[1105]) );
  XNOR U5826 ( .A(round_reg[910]), .B(n4645), .Z(n4557) );
  XOR U5827 ( .A(n5003), .B(n5004), .Z(n4645) );
  ANDN U5828 ( .B(n1156), .A(n4764), .Z(n5002) );
  XOR U5829 ( .A(n5005), .B(n4559), .Z(out[1104]) );
  XNOR U5830 ( .A(round_reg[909]), .B(n4672), .Z(n4559) );
  XOR U5831 ( .A(n5006), .B(n5007), .Z(n4672) );
  ANDN U5832 ( .B(n1160), .A(n4768), .Z(n5005) );
  XOR U5833 ( .A(n5008), .B(n4561), .Z(out[1103]) );
  XNOR U5834 ( .A(round_reg[908]), .B(n4387), .Z(n4561) );
  XOR U5835 ( .A(n5009), .B(n5010), .Z(n4387) );
  NOR U5836 ( .A(n1164), .B(n4772), .Z(n5008) );
  XOR U5837 ( .A(n5011), .B(n4563), .Z(out[1102]) );
  XNOR U5838 ( .A(round_reg[907]), .B(n4758), .Z(n4563) );
  XOR U5839 ( .A(n5012), .B(n5013), .Z(n4758) );
  ANDN U5840 ( .B(n1168), .A(n4776), .Z(n5011) );
  XOR U5841 ( .A(n5014), .B(n4567), .Z(out[1101]) );
  XOR U5842 ( .A(round_reg[906]), .B(n2265), .Z(n4567) );
  XNOR U5843 ( .A(n5015), .B(n5016), .Z(n2265) );
  ANDN U5844 ( .B(n1172), .A(n4780), .Z(n5014) );
  XOR U5845 ( .A(n5017), .B(n4569), .Z(out[1100]) );
  XOR U5846 ( .A(round_reg[905]), .B(n2269), .Z(n4569) );
  XNOR U5847 ( .A(n5018), .B(n5019), .Z(n2269) );
  ANDN U5848 ( .B(n1176), .A(n4784), .Z(n5017) );
  XOR U5849 ( .A(n5020), .B(n1991), .Z(out[10]) );
  XOR U5850 ( .A(round_reg[200]), .B(n2351), .Z(n1991) );
  IV U5851 ( .A(n5021), .Z(n2351) );
  ANDN U5852 ( .B(n3389), .A(n3390), .Z(n5020) );
  XOR U5853 ( .A(round_reg[1043]), .B(n1777), .Z(n3390) );
  XNOR U5854 ( .A(round_reg[1420]), .B(n2310), .Z(n3389) );
  XOR U5855 ( .A(n5022), .B(n3459), .Z(out[109]) );
  IV U5856 ( .A(n3560), .Z(n3459) );
  XNOR U5857 ( .A(round_reg[580]), .B(n2289), .Z(n3560) );
  ANDN U5858 ( .B(n2980), .A(n2982), .Z(n5022) );
  XNOR U5859 ( .A(round_reg[1455]), .B(n2154), .Z(n2982) );
  XNOR U5860 ( .A(round_reg[235]), .B(n2195), .Z(n2980) );
  XOR U5861 ( .A(n5023), .B(n4572), .Z(out[1099]) );
  XOR U5862 ( .A(round_reg[904]), .B(n2273), .Z(n4572) );
  XNOR U5863 ( .A(n5024), .B(n5025), .Z(n2273) );
  ANDN U5864 ( .B(n1180), .A(n4788), .Z(n5023) );
  XOR U5865 ( .A(n5026), .B(n4575), .Z(out[1098]) );
  XOR U5866 ( .A(round_reg[903]), .B(n2277), .Z(n4575) );
  XNOR U5867 ( .A(n5027), .B(n5028), .Z(n2277) );
  ANDN U5868 ( .B(n1184), .A(n4792), .Z(n5026) );
  XOR U5869 ( .A(n5029), .B(n4578), .Z(out[1097]) );
  XOR U5870 ( .A(round_reg[902]), .B(n2281), .Z(n4578) );
  XNOR U5871 ( .A(n5030), .B(n5031), .Z(n2281) );
  ANDN U5872 ( .B(n1192), .A(n4796), .Z(n5029) );
  XOR U5873 ( .A(n5032), .B(n4581), .Z(out[1096]) );
  XOR U5874 ( .A(round_reg[901]), .B(n2285), .Z(n4581) );
  XNOR U5875 ( .A(n5033), .B(n5034), .Z(n2285) );
  NOR U5876 ( .A(n1196), .B(n4800), .Z(n5032) );
  XOR U5877 ( .A(n5035), .B(n4583), .Z(out[1095]) );
  XOR U5878 ( .A(round_reg[900]), .B(n2289), .Z(n4583) );
  XNOR U5879 ( .A(n5036), .B(n5037), .Z(n2289) );
  NOR U5880 ( .A(n1200), .B(n4807), .Z(n5035) );
  XOR U5881 ( .A(n5038), .B(n4585), .Z(out[1094]) );
  XOR U5882 ( .A(round_reg[899]), .B(n2293), .Z(n4585) );
  NOR U5883 ( .A(n1204), .B(n4811), .Z(n5038) );
  XOR U5884 ( .A(n5039), .B(n4587), .Z(out[1093]) );
  XOR U5885 ( .A(round_reg[898]), .B(n2297), .Z(n4587) );
  NOR U5886 ( .A(n1208), .B(n4815), .Z(n5039) );
  XOR U5887 ( .A(n5040), .B(n4590), .Z(out[1092]) );
  XOR U5888 ( .A(round_reg[897]), .B(n2305), .Z(n4590) );
  NOR U5889 ( .A(n1212), .B(n4819), .Z(n5040) );
  XOR U5890 ( .A(n5041), .B(n4596), .Z(out[1091]) );
  XOR U5891 ( .A(round_reg[896]), .B(n2309), .Z(n4596) );
  NOR U5892 ( .A(n1216), .B(n4823), .Z(n5041) );
  XOR U5893 ( .A(n5042), .B(n4599), .Z(out[1090]) );
  XOR U5894 ( .A(round_reg[959]), .B(n2313), .Z(n4599) );
  NOR U5895 ( .A(n1220), .B(n4827), .Z(n5042) );
  XOR U5896 ( .A(n5043), .B(n3461), .Z(out[108]) );
  IV U5897 ( .A(n3562), .Z(n3461) );
  XNOR U5898 ( .A(round_reg[579]), .B(n2293), .Z(n3562) );
  XNOR U5899 ( .A(n5044), .B(n5045), .Z(n2293) );
  ANDN U5900 ( .B(n3007), .A(n3009), .Z(n5043) );
  XNOR U5901 ( .A(round_reg[1454]), .B(n2158), .Z(n3009) );
  XNOR U5902 ( .A(round_reg[234]), .B(n2199), .Z(n3007) );
  XOR U5903 ( .A(n5046), .B(n4602), .Z(out[1089]) );
  XOR U5904 ( .A(round_reg[958]), .B(n2317), .Z(n4602) );
  NOR U5905 ( .A(n1224), .B(n4831), .Z(n5046) );
  XOR U5906 ( .A(n5047), .B(n4605), .Z(out[1088]) );
  XOR U5907 ( .A(round_reg[957]), .B(n2321), .Z(n4605) );
  NOR U5908 ( .A(n1228), .B(n4835), .Z(n5047) );
  XOR U5909 ( .A(n5048), .B(n4608), .Z(out[1087]) );
  XNOR U5910 ( .A(round_reg[530]), .B(n4294), .Z(n4608) );
  XOR U5911 ( .A(n4664), .B(n5049), .Z(n4294) );
  XOR U5912 ( .A(n5050), .B(n5051), .Z(n4664) );
  XNOR U5913 ( .A(round_reg[1554]), .B(round_reg[1234]), .Z(n5051) );
  XOR U5914 ( .A(round_reg[274]), .B(n5052), .Z(n5050) );
  XOR U5915 ( .A(round_reg[914]), .B(round_reg[594]), .Z(n5052) );
  ANDN U5916 ( .B(n4407), .A(n4837), .Z(n5048) );
  XOR U5917 ( .A(n5053), .B(n4610), .Z(out[1086]) );
  XNOR U5918 ( .A(round_reg[529]), .B(n4296), .Z(n4610) );
  XOR U5919 ( .A(n4668), .B(n5054), .Z(n4296) );
  XOR U5920 ( .A(n5055), .B(n5056), .Z(n4668) );
  XNOR U5921 ( .A(round_reg[1553]), .B(round_reg[1233]), .Z(n5056) );
  XOR U5922 ( .A(round_reg[273]), .B(n5057), .Z(n5055) );
  XOR U5923 ( .A(round_reg[913]), .B(round_reg[593]), .Z(n5057) );
  ANDN U5924 ( .B(n4411), .A(n4839), .Z(n5053) );
  XOR U5925 ( .A(n5058), .B(n4612), .Z(out[1085]) );
  XNOR U5926 ( .A(round_reg[528]), .B(n4298), .Z(n4612) );
  XOR U5927 ( .A(n4675), .B(n5059), .Z(n4298) );
  XOR U5928 ( .A(n5060), .B(n5061), .Z(n4675) );
  XNOR U5929 ( .A(round_reg[1552]), .B(round_reg[1232]), .Z(n5061) );
  XOR U5930 ( .A(round_reg[272]), .B(n5062), .Z(n5060) );
  XOR U5931 ( .A(round_reg[912]), .B(round_reg[592]), .Z(n5062) );
  ANDN U5932 ( .B(n4415), .A(n4845), .Z(n5058) );
  XOR U5933 ( .A(n5063), .B(n4614), .Z(out[1084]) );
  XNOR U5934 ( .A(round_reg[527]), .B(n4301), .Z(n4614) );
  XOR U5935 ( .A(n4679), .B(n5064), .Z(n4301) );
  XOR U5936 ( .A(n5065), .B(n5066), .Z(n4679) );
  XNOR U5937 ( .A(round_reg[1551]), .B(round_reg[1231]), .Z(n5066) );
  XOR U5938 ( .A(round_reg[271]), .B(n5067), .Z(n5065) );
  XOR U5939 ( .A(round_reg[911]), .B(round_reg[591]), .Z(n5067) );
  ANDN U5940 ( .B(n4419), .A(n4849), .Z(n5063) );
  XOR U5941 ( .A(n5068), .B(n4616), .Z(out[1083]) );
  XNOR U5942 ( .A(round_reg[526]), .B(n4303), .Z(n4616) );
  XOR U5943 ( .A(n4683), .B(n5069), .Z(n4303) );
  XOR U5944 ( .A(n5070), .B(n5071), .Z(n4683) );
  XNOR U5945 ( .A(round_reg[1550]), .B(round_reg[1230]), .Z(n5071) );
  XOR U5946 ( .A(round_reg[270]), .B(n5072), .Z(n5070) );
  XOR U5947 ( .A(round_reg[910]), .B(round_reg[590]), .Z(n5072) );
  ANDN U5948 ( .B(n4423), .A(n4853), .Z(n5068) );
  XOR U5949 ( .A(n5073), .B(n4618), .Z(out[1082]) );
  XNOR U5950 ( .A(round_reg[525]), .B(n4306), .Z(n4618) );
  XOR U5951 ( .A(n4687), .B(n5074), .Z(n4306) );
  XOR U5952 ( .A(n5075), .B(n5076), .Z(n4687) );
  XNOR U5953 ( .A(round_reg[1549]), .B(round_reg[1229]), .Z(n5076) );
  XOR U5954 ( .A(round_reg[269]), .B(n5077), .Z(n5075) );
  XOR U5955 ( .A(round_reg[909]), .B(round_reg[589]), .Z(n5077) );
  ANDN U5956 ( .B(n4427), .A(n4857), .Z(n5073) );
  XOR U5957 ( .A(n5078), .B(n4623), .Z(out[1081]) );
  XNOR U5958 ( .A(round_reg[524]), .B(n4309), .Z(n4623) );
  XOR U5959 ( .A(n5079), .B(n4692), .Z(n4309) );
  XNOR U5960 ( .A(n5080), .B(n5081), .Z(n4692) );
  XNOR U5961 ( .A(round_reg[1548]), .B(round_reg[1228]), .Z(n5081) );
  XOR U5962 ( .A(round_reg[268]), .B(n5082), .Z(n5080) );
  XOR U5963 ( .A(round_reg[908]), .B(round_reg[588]), .Z(n5082) );
  ANDN U5964 ( .B(n4431), .A(n4861), .Z(n5078) );
  XOR U5965 ( .A(n5083), .B(n4625), .Z(out[1080]) );
  XNOR U5966 ( .A(round_reg[523]), .B(n4311), .Z(n4625) );
  XOR U5967 ( .A(n5084), .B(n4696), .Z(n4311) );
  XNOR U5968 ( .A(n5085), .B(n5086), .Z(n4696) );
  XNOR U5969 ( .A(round_reg[1547]), .B(round_reg[1227]), .Z(n5086) );
  XOR U5970 ( .A(round_reg[267]), .B(n5087), .Z(n5085) );
  XOR U5971 ( .A(round_reg[907]), .B(round_reg[587]), .Z(n5087) );
  ANDN U5972 ( .B(n4435), .A(n4865), .Z(n5083) );
  XOR U5973 ( .A(n5088), .B(n3463), .Z(out[107]) );
  IV U5974 ( .A(n3564), .Z(n3463) );
  XNOR U5975 ( .A(round_reg[578]), .B(n2297), .Z(n3564) );
  XNOR U5976 ( .A(n5089), .B(n5090), .Z(n2297) );
  ANDN U5977 ( .B(n3023), .A(n3025), .Z(n5088) );
  XNOR U5978 ( .A(round_reg[1453]), .B(n2162), .Z(n3025) );
  XNOR U5979 ( .A(round_reg[233]), .B(n2203), .Z(n3023) );
  XOR U5980 ( .A(n5091), .B(n4627), .Z(out[1079]) );
  XNOR U5981 ( .A(round_reg[522]), .B(n4376), .Z(n4627) );
  XOR U5982 ( .A(n5092), .B(n4700), .Z(n4376) );
  XNOR U5983 ( .A(n5093), .B(n5094), .Z(n4700) );
  XNOR U5984 ( .A(round_reg[1546]), .B(round_reg[1226]), .Z(n5094) );
  XOR U5985 ( .A(round_reg[266]), .B(n5095), .Z(n5093) );
  XOR U5986 ( .A(round_reg[906]), .B(round_reg[586]), .Z(n5095) );
  ANDN U5987 ( .B(n4439), .A(n4869), .Z(n5091) );
  XOR U5988 ( .A(n5096), .B(n4629), .Z(out[1078]) );
  XNOR U5989 ( .A(round_reg[521]), .B(n4643), .Z(n4629) );
  XOR U5990 ( .A(n5097), .B(n4704), .Z(n4643) );
  XNOR U5991 ( .A(n5098), .B(n5099), .Z(n4704) );
  XNOR U5992 ( .A(round_reg[1545]), .B(round_reg[1225]), .Z(n5099) );
  XOR U5993 ( .A(round_reg[265]), .B(n5100), .Z(n5098) );
  XOR U5994 ( .A(round_reg[905]), .B(round_reg[585]), .Z(n5100) );
  ANDN U5995 ( .B(n4443), .A(n4873), .Z(n5096) );
  XOR U5996 ( .A(n5101), .B(n4631), .Z(out[1077]) );
  XNOR U5997 ( .A(round_reg[520]), .B(n5021), .Z(n4631) );
  XOR U5998 ( .A(n5102), .B(n4708), .Z(n5021) );
  XNOR U5999 ( .A(n5103), .B(n5104), .Z(n4708) );
  XNOR U6000 ( .A(round_reg[1544]), .B(round_reg[1224]), .Z(n5104) );
  XOR U6001 ( .A(round_reg[264]), .B(n5105), .Z(n5103) );
  XOR U6002 ( .A(round_reg[904]), .B(round_reg[584]), .Z(n5105) );
  ANDN U6003 ( .B(n4449), .A(n4877), .Z(n5101) );
  XOR U6004 ( .A(n5106), .B(n4633), .Z(out[1076]) );
  XOR U6005 ( .A(round_reg[519]), .B(n2355), .Z(n4633) );
  XOR U6006 ( .A(n4711), .B(n5107), .Z(n2355) );
  XOR U6007 ( .A(n5108), .B(n5109), .Z(n4711) );
  XNOR U6008 ( .A(round_reg[1543]), .B(round_reg[1223]), .Z(n5109) );
  XOR U6009 ( .A(round_reg[263]), .B(n5110), .Z(n5108) );
  XOR U6010 ( .A(round_reg[903]), .B(round_reg[583]), .Z(n5110) );
  ANDN U6011 ( .B(n4453), .A(n4881), .Z(n5106) );
  XOR U6012 ( .A(n5111), .B(n4635), .Z(out[1075]) );
  XNOR U6013 ( .A(round_reg[518]), .B(n4317), .Z(n4635) );
  XOR U6014 ( .A(n5112), .B(n4719), .Z(n4317) );
  XNOR U6015 ( .A(n5113), .B(n5114), .Z(n4719) );
  XNOR U6016 ( .A(round_reg[1542]), .B(round_reg[1222]), .Z(n5114) );
  XOR U6017 ( .A(round_reg[262]), .B(n5115), .Z(n5113) );
  XOR U6018 ( .A(round_reg[902]), .B(round_reg[582]), .Z(n5115) );
  ANDN U6019 ( .B(n4457), .A(n4887), .Z(n5111) );
  XOR U6020 ( .A(n5116), .B(n4637), .Z(out[1074]) );
  XNOR U6021 ( .A(round_reg[517]), .B(n4320), .Z(n4637) );
  XOR U6022 ( .A(n5117), .B(n4723), .Z(n4320) );
  XNOR U6023 ( .A(n5118), .B(n5119), .Z(n4723) );
  XNOR U6024 ( .A(round_reg[1541]), .B(round_reg[1221]), .Z(n5119) );
  XOR U6025 ( .A(round_reg[261]), .B(n5120), .Z(n5118) );
  XOR U6026 ( .A(round_reg[901]), .B(round_reg[581]), .Z(n5120) );
  ANDN U6027 ( .B(n4461), .A(n4891), .Z(n5116) );
  XOR U6028 ( .A(n5121), .B(n4639), .Z(out[1073]) );
  XNOR U6029 ( .A(round_reg[516]), .B(n4322), .Z(n4639) );
  XOR U6030 ( .A(n5122), .B(n4727), .Z(n4322) );
  XNOR U6031 ( .A(n5123), .B(n5124), .Z(n4727) );
  XNOR U6032 ( .A(round_reg[1540]), .B(round_reg[1220]), .Z(n5124) );
  XOR U6033 ( .A(round_reg[260]), .B(n5125), .Z(n5123) );
  XOR U6034 ( .A(round_reg[900]), .B(round_reg[580]), .Z(n5125) );
  ANDN U6035 ( .B(n4465), .A(n4895), .Z(n5121) );
  XOR U6036 ( .A(n5126), .B(n4641), .Z(out[1072]) );
  XNOR U6037 ( .A(round_reg[515]), .B(n4325), .Z(n4641) );
  XOR U6038 ( .A(n5127), .B(n4731), .Z(n4325) );
  XNOR U6039 ( .A(n5128), .B(n5129), .Z(n4731) );
  XNOR U6040 ( .A(round_reg[1539]), .B(round_reg[1219]), .Z(n5129) );
  XOR U6041 ( .A(round_reg[259]), .B(n5130), .Z(n5128) );
  XOR U6042 ( .A(round_reg[899]), .B(round_reg[579]), .Z(n5130) );
  ANDN U6043 ( .B(n4469), .A(n4899), .Z(n5126) );
  XOR U6044 ( .A(n5131), .B(n4648), .Z(out[1071]) );
  XNOR U6045 ( .A(round_reg[514]), .B(n4328), .Z(n4648) );
  XOR U6046 ( .A(n5132), .B(n4735), .Z(n4328) );
  XNOR U6047 ( .A(n5133), .B(n5134), .Z(n4735) );
  XNOR U6048 ( .A(round_reg[1538]), .B(round_reg[1218]), .Z(n5134) );
  XOR U6049 ( .A(round_reg[258]), .B(n5135), .Z(n5133) );
  XOR U6050 ( .A(round_reg[898]), .B(round_reg[578]), .Z(n5135) );
  ANDN U6051 ( .B(n4473), .A(n4903), .Z(n5131) );
  XOR U6052 ( .A(n5136), .B(n4650), .Z(out[1070]) );
  XNOR U6053 ( .A(round_reg[513]), .B(n4339), .Z(n4650) );
  XOR U6054 ( .A(n5137), .B(n4739), .Z(n4339) );
  XNOR U6055 ( .A(n5138), .B(n5139), .Z(n4739) );
  XNOR U6056 ( .A(round_reg[1537]), .B(round_reg[1217]), .Z(n5139) );
  XOR U6057 ( .A(round_reg[257]), .B(n5140), .Z(n5138) );
  XOR U6058 ( .A(round_reg[897]), .B(round_reg[577]), .Z(n5140) );
  ANDN U6059 ( .B(n4477), .A(n4907), .Z(n5136) );
  XOR U6060 ( .A(n5141), .B(n3465), .Z(out[106]) );
  IV U6061 ( .A(n3566), .Z(n3465) );
  XNOR U6062 ( .A(round_reg[577]), .B(n2305), .Z(n3566) );
  XNOR U6063 ( .A(n5142), .B(n5143), .Z(n2305) );
  ANDN U6064 ( .B(n3042), .A(n3044), .Z(n5141) );
  XNOR U6065 ( .A(round_reg[1452]), .B(n2166), .Z(n3044) );
  XNOR U6066 ( .A(round_reg[232]), .B(n2207), .Z(n3042) );
  XOR U6067 ( .A(n5144), .B(n4652), .Z(out[1069]) );
  XNOR U6068 ( .A(round_reg[512]), .B(n4356), .Z(n4652) );
  XOR U6069 ( .A(n5145), .B(n4743), .Z(n4356) );
  XNOR U6070 ( .A(n5146), .B(n5147), .Z(n4743) );
  XNOR U6071 ( .A(round_reg[1536]), .B(round_reg[1216]), .Z(n5147) );
  XOR U6072 ( .A(round_reg[256]), .B(n5148), .Z(n5146) );
  XOR U6073 ( .A(round_reg[896]), .B(round_reg[576]), .Z(n5148) );
  ANDN U6074 ( .B(n4481), .A(n4911), .Z(n5144) );
  XOR U6075 ( .A(n5149), .B(n4654), .Z(out[1068]) );
  XNOR U6076 ( .A(round_reg[575]), .B(n4378), .Z(n4654) );
  XOR U6077 ( .A(n5150), .B(n4747), .Z(n4378) );
  XNOR U6078 ( .A(n5151), .B(n5152), .Z(n4747) );
  XNOR U6079 ( .A(round_reg[1599]), .B(round_reg[1279]), .Z(n5152) );
  XOR U6080 ( .A(round_reg[319]), .B(n5153), .Z(n5151) );
  XOR U6081 ( .A(round_reg[959]), .B(round_reg[639]), .Z(n5153) );
  ANDN U6082 ( .B(n4485), .A(n4915), .Z(n5149) );
  XOR U6083 ( .A(n5154), .B(n4656), .Z(out[1067]) );
  XNOR U6084 ( .A(round_reg[574]), .B(n2107), .Z(n4656) );
  ANDN U6085 ( .B(n4491), .A(n4919), .Z(n5154) );
  XOR U6086 ( .A(n5155), .B(n4658), .Z(out[1066]) );
  XNOR U6087 ( .A(round_reg[573]), .B(n2111), .Z(n4658) );
  XOR U6088 ( .A(n5156), .B(n4755), .Z(n2111) );
  XNOR U6089 ( .A(n5157), .B(n5158), .Z(n4755) );
  XNOR U6090 ( .A(round_reg[1597]), .B(round_reg[1277]), .Z(n5158) );
  XOR U6091 ( .A(round_reg[317]), .B(n5159), .Z(n5157) );
  XOR U6092 ( .A(round_reg[957]), .B(round_reg[637]), .Z(n5159) );
  ANDN U6093 ( .B(n4495), .A(n4923), .Z(n5155) );
  XOR U6094 ( .A(n5160), .B(n4660), .Z(out[1065]) );
  XOR U6095 ( .A(round_reg[572]), .B(n2115), .Z(n4660) );
  XNOR U6096 ( .A(n5161), .B(n4763), .Z(n2115) );
  XNOR U6097 ( .A(n5162), .B(n5163), .Z(n4763) );
  XNOR U6098 ( .A(round_reg[1596]), .B(round_reg[1276]), .Z(n5163) );
  XOR U6099 ( .A(round_reg[316]), .B(n5164), .Z(n5162) );
  XOR U6100 ( .A(round_reg[956]), .B(round_reg[636]), .Z(n5164) );
  ANDN U6101 ( .B(n4499), .A(n4929), .Z(n5160) );
  XOR U6102 ( .A(n5165), .B(n4662), .Z(out[1064]) );
  XOR U6103 ( .A(round_reg[571]), .B(n2119), .Z(n4662) );
  XNOR U6104 ( .A(n5166), .B(n4767), .Z(n2119) );
  XNOR U6105 ( .A(n5167), .B(n5168), .Z(n4767) );
  XNOR U6106 ( .A(round_reg[1595]), .B(round_reg[1275]), .Z(n5168) );
  XOR U6107 ( .A(round_reg[315]), .B(n5169), .Z(n5167) );
  XOR U6108 ( .A(round_reg[955]), .B(round_reg[635]), .Z(n5169) );
  ANDN U6109 ( .B(n4503), .A(n4933), .Z(n5165) );
  XOR U6110 ( .A(n5170), .B(n4666), .Z(out[1063]) );
  XNOR U6111 ( .A(round_reg[570]), .B(n2130), .Z(n4666) );
  XOR U6112 ( .A(n5171), .B(n4771), .Z(n2130) );
  XNOR U6113 ( .A(n5172), .B(n5173), .Z(n4771) );
  XNOR U6114 ( .A(round_reg[1594]), .B(round_reg[1274]), .Z(n5173) );
  XOR U6115 ( .A(round_reg[314]), .B(n5174), .Z(n5172) );
  XOR U6116 ( .A(round_reg[954]), .B(round_reg[634]), .Z(n5174) );
  ANDN U6117 ( .B(n1062), .A(n1060), .Z(n5170) );
  XOR U6118 ( .A(round_reg[170]), .B(n2178), .Z(n1060) );
  XOR U6119 ( .A(round_reg[1355]), .B(n1805), .Z(n1062) );
  XOR U6120 ( .A(n5079), .B(n5015), .Z(n1805) );
  XOR U6121 ( .A(n5175), .B(n5176), .Z(n5015) );
  XNOR U6122 ( .A(round_reg[1290]), .B(round_reg[10]), .Z(n5176) );
  XOR U6123 ( .A(round_reg[330]), .B(n5177), .Z(n5175) );
  XOR U6124 ( .A(round_reg[970]), .B(round_reg[650]), .Z(n5177) );
  XOR U6125 ( .A(n5178), .B(n5179), .Z(n5079) );
  XNOR U6126 ( .A(round_reg[139]), .B(round_reg[1099]), .Z(n5179) );
  XOR U6127 ( .A(round_reg[1419]), .B(n5180), .Z(n5178) );
  XOR U6128 ( .A(round_reg[779]), .B(round_reg[459]), .Z(n5180) );
  XOR U6129 ( .A(n5181), .B(n4670), .Z(out[1062]) );
  XNOR U6130 ( .A(round_reg[569]), .B(n4542), .Z(n4670) );
  XOR U6131 ( .A(n5182), .B(n4775), .Z(n4542) );
  XNOR U6132 ( .A(n5183), .B(n5184), .Z(n4775) );
  XNOR U6133 ( .A(round_reg[1593]), .B(round_reg[1273]), .Z(n5184) );
  XOR U6134 ( .A(round_reg[313]), .B(n5185), .Z(n5183) );
  XOR U6135 ( .A(round_reg[953]), .B(round_reg[633]), .Z(n5185) );
  NOR U6136 ( .A(n1066), .B(n1064), .Z(n5181) );
  XOR U6137 ( .A(round_reg[169]), .B(n2182), .Z(n1064) );
  XNOR U6138 ( .A(round_reg[1354]), .B(n1808), .Z(n1066) );
  XOR U6139 ( .A(n5084), .B(n5018), .Z(n1808) );
  XOR U6140 ( .A(n5186), .B(n5187), .Z(n5018) );
  XNOR U6141 ( .A(round_reg[329]), .B(round_reg[1289]), .Z(n5187) );
  XOR U6142 ( .A(round_reg[649]), .B(n5188), .Z(n5186) );
  XOR U6143 ( .A(round_reg[9]), .B(round_reg[969]), .Z(n5188) );
  XOR U6144 ( .A(n5189), .B(n5190), .Z(n5084) );
  XNOR U6145 ( .A(round_reg[138]), .B(round_reg[1098]), .Z(n5190) );
  XOR U6146 ( .A(round_reg[1418]), .B(n5191), .Z(n5189) );
  XOR U6147 ( .A(round_reg[778]), .B(round_reg[458]), .Z(n5191) );
  XOR U6148 ( .A(n5192), .B(n4677), .Z(out[1061]) );
  XNOR U6149 ( .A(round_reg[568]), .B(n4565), .Z(n4677) );
  XOR U6150 ( .A(n5193), .B(n4779), .Z(n4565) );
  XNOR U6151 ( .A(n5194), .B(n5195), .Z(n4779) );
  XNOR U6152 ( .A(round_reg[1592]), .B(round_reg[1272]), .Z(n5195) );
  XOR U6153 ( .A(round_reg[312]), .B(n5196), .Z(n5194) );
  XOR U6154 ( .A(round_reg[952]), .B(round_reg[632]), .Z(n5196) );
  ANDN U6155 ( .B(n1070), .A(n1068), .Z(n5192) );
  XOR U6156 ( .A(round_reg[168]), .B(n2186), .Z(n1068) );
  XOR U6157 ( .A(round_reg[1353]), .B(n1811), .Z(n1070) );
  XOR U6158 ( .A(n5197), .B(n4681), .Z(out[1060]) );
  XNOR U6159 ( .A(round_reg[567]), .B(n4594), .Z(n4681) );
  XOR U6160 ( .A(n5198), .B(n4782), .Z(n4594) );
  XNOR U6161 ( .A(n5199), .B(n5200), .Z(n4782) );
  XNOR U6162 ( .A(round_reg[1591]), .B(round_reg[1271]), .Z(n5200) );
  XOR U6163 ( .A(round_reg[311]), .B(n5201), .Z(n5199) );
  XOR U6164 ( .A(round_reg[951]), .B(round_reg[631]), .Z(n5201) );
  ANDN U6165 ( .B(n1074), .A(n1072), .Z(n5197) );
  XOR U6166 ( .A(round_reg[167]), .B(n2190), .Z(n1072) );
  XOR U6167 ( .A(round_reg[1352]), .B(n1814), .Z(n1074) );
  XOR U6168 ( .A(n5097), .B(n5027), .Z(n1814) );
  XOR U6169 ( .A(n5202), .B(n5203), .Z(n5027) );
  XNOR U6170 ( .A(round_reg[327]), .B(round_reg[1287]), .Z(n5203) );
  XOR U6171 ( .A(round_reg[647]), .B(n5204), .Z(n5202) );
  XOR U6172 ( .A(round_reg[967]), .B(round_reg[7]), .Z(n5204) );
  XOR U6173 ( .A(n5205), .B(n5206), .Z(n5097) );
  XNOR U6174 ( .A(round_reg[136]), .B(round_reg[1096]), .Z(n5206) );
  XOR U6175 ( .A(round_reg[1416]), .B(n5207), .Z(n5205) );
  XOR U6176 ( .A(round_reg[776]), .B(round_reg[456]), .Z(n5207) );
  XOR U6177 ( .A(n5208), .B(n3467), .Z(out[105]) );
  IV U6178 ( .A(n3569), .Z(n3467) );
  XNOR U6179 ( .A(round_reg[576]), .B(n2309), .Z(n3569) );
  XNOR U6180 ( .A(n5209), .B(n5210), .Z(n2309) );
  ANDN U6181 ( .B(n3065), .A(n3067), .Z(n5208) );
  XNOR U6182 ( .A(round_reg[1451]), .B(n2174), .Z(n3067) );
  XNOR U6183 ( .A(round_reg[231]), .B(n2211), .Z(n3065) );
  XOR U6184 ( .A(n5211), .B(n4685), .Z(out[1059]) );
  XNOR U6185 ( .A(round_reg[566]), .B(n4621), .Z(n4685) );
  XOR U6186 ( .A(n5212), .B(n4786), .Z(n4621) );
  XNOR U6187 ( .A(n5213), .B(n5214), .Z(n4786) );
  XNOR U6188 ( .A(round_reg[1590]), .B(round_reg[1270]), .Z(n5214) );
  XOR U6189 ( .A(round_reg[310]), .B(n5215), .Z(n5213) );
  XOR U6190 ( .A(round_reg[950]), .B(round_reg[630]), .Z(n5215) );
  ANDN U6191 ( .B(n1078), .A(n1076), .Z(n5211) );
  XOR U6192 ( .A(round_reg[166]), .B(n2194), .Z(n1076) );
  XOR U6193 ( .A(round_reg[1351]), .B(n1817), .Z(n1078) );
  XOR U6194 ( .A(n5102), .B(n5030), .Z(n1817) );
  XOR U6195 ( .A(n5216), .B(n5217), .Z(n5030) );
  XNOR U6196 ( .A(round_reg[326]), .B(round_reg[1286]), .Z(n5217) );
  XOR U6197 ( .A(round_reg[646]), .B(n5218), .Z(n5216) );
  XOR U6198 ( .A(round_reg[966]), .B(round_reg[6]), .Z(n5218) );
  XOR U6199 ( .A(n5219), .B(n5220), .Z(n5102) );
  XNOR U6200 ( .A(round_reg[135]), .B(round_reg[1095]), .Z(n5220) );
  XOR U6201 ( .A(round_reg[1415]), .B(n5221), .Z(n5219) );
  XOR U6202 ( .A(round_reg[775]), .B(round_reg[455]), .Z(n5221) );
  XOR U6203 ( .A(n5222), .B(n4689), .Z(out[1058]) );
  XNOR U6204 ( .A(round_reg[565]), .B(n4646), .Z(n4689) );
  XOR U6205 ( .A(n5223), .B(n4790), .Z(n4646) );
  XNOR U6206 ( .A(n5224), .B(n5225), .Z(n4790) );
  XNOR U6207 ( .A(round_reg[1589]), .B(round_reg[1269]), .Z(n5225) );
  XOR U6208 ( .A(round_reg[309]), .B(n5226), .Z(n5224) );
  XOR U6209 ( .A(round_reg[949]), .B(round_reg[629]), .Z(n5226) );
  ANDN U6210 ( .B(n1082), .A(n1080), .Z(n5222) );
  XOR U6211 ( .A(round_reg[165]), .B(n2198), .Z(n1080) );
  XOR U6212 ( .A(n4927), .B(n5227), .Z(n2198) );
  XOR U6213 ( .A(n5228), .B(n5229), .Z(n4927) );
  XNOR U6214 ( .A(round_reg[1509]), .B(round_reg[1189]), .Z(n5229) );
  XOR U6215 ( .A(round_reg[229]), .B(n5230), .Z(n5228) );
  XOR U6216 ( .A(round_reg[869]), .B(round_reg[549]), .Z(n5230) );
  XOR U6217 ( .A(round_reg[1350]), .B(n1828), .Z(n1082) );
  XOR U6218 ( .A(n5107), .B(n5033), .Z(n1828) );
  XOR U6219 ( .A(n5231), .B(n5232), .Z(n5033) );
  XNOR U6220 ( .A(round_reg[325]), .B(round_reg[1285]), .Z(n5232) );
  XOR U6221 ( .A(round_reg[5]), .B(n5233), .Z(n5231) );
  XOR U6222 ( .A(round_reg[965]), .B(round_reg[645]), .Z(n5233) );
  XOR U6223 ( .A(n5234), .B(n5235), .Z(n5107) );
  XNOR U6224 ( .A(round_reg[134]), .B(round_reg[1094]), .Z(n5235) );
  XOR U6225 ( .A(round_reg[1414]), .B(n5236), .Z(n5234) );
  XOR U6226 ( .A(round_reg[774]), .B(round_reg[454]), .Z(n5236) );
  XOR U6227 ( .A(n5237), .B(n4693), .Z(out[1057]) );
  XNOR U6228 ( .A(round_reg[564]), .B(n4673), .Z(n4693) );
  XOR U6229 ( .A(n5238), .B(n4794), .Z(n4673) );
  XNOR U6230 ( .A(n5239), .B(n5240), .Z(n4794) );
  XNOR U6231 ( .A(round_reg[1588]), .B(round_reg[1268]), .Z(n5240) );
  XOR U6232 ( .A(round_reg[308]), .B(n5241), .Z(n5239) );
  XOR U6233 ( .A(round_reg[948]), .B(round_reg[628]), .Z(n5241) );
  ANDN U6234 ( .B(n1086), .A(n1084), .Z(n5237) );
  XOR U6235 ( .A(round_reg[164]), .B(n2202), .Z(n1084) );
  XOR U6236 ( .A(n4931), .B(n5242), .Z(n2202) );
  XOR U6237 ( .A(n5243), .B(n5244), .Z(n4931) );
  XNOR U6238 ( .A(round_reg[1508]), .B(round_reg[1188]), .Z(n5244) );
  XOR U6239 ( .A(round_reg[228]), .B(n5245), .Z(n5243) );
  XOR U6240 ( .A(round_reg[868]), .B(round_reg[548]), .Z(n5245) );
  XOR U6241 ( .A(round_reg[1349]), .B(n1831), .Z(n1086) );
  XOR U6242 ( .A(n5112), .B(n5036), .Z(n1831) );
  XOR U6243 ( .A(n5246), .B(n5247), .Z(n5036) );
  XNOR U6244 ( .A(round_reg[324]), .B(round_reg[1284]), .Z(n5247) );
  XOR U6245 ( .A(round_reg[4]), .B(n5248), .Z(n5246) );
  XOR U6246 ( .A(round_reg[964]), .B(round_reg[644]), .Z(n5248) );
  XOR U6247 ( .A(n5249), .B(n5250), .Z(n5112) );
  XNOR U6248 ( .A(round_reg[133]), .B(round_reg[1093]), .Z(n5250) );
  XOR U6249 ( .A(round_reg[1413]), .B(n5251), .Z(n5249) );
  XOR U6250 ( .A(round_reg[773]), .B(round_reg[453]), .Z(n5251) );
  XOR U6251 ( .A(n5252), .B(n4697), .Z(out[1056]) );
  XNOR U6252 ( .A(round_reg[563]), .B(n4716), .Z(n4697) );
  XOR U6253 ( .A(n5253), .B(n4799), .Z(n4716) );
  XNOR U6254 ( .A(n5254), .B(n5255), .Z(n4799) );
  XNOR U6255 ( .A(round_reg[1587]), .B(round_reg[1267]), .Z(n5255) );
  XOR U6256 ( .A(round_reg[307]), .B(n5256), .Z(n5254) );
  XOR U6257 ( .A(round_reg[947]), .B(round_reg[627]), .Z(n5256) );
  ANDN U6258 ( .B(n1090), .A(n1088), .Z(n5252) );
  XNOR U6259 ( .A(round_reg[163]), .B(n3032), .Z(n1088) );
  IV U6260 ( .A(n2206), .Z(n3032) );
  XOR U6261 ( .A(n5257), .B(n5258), .Z(n4935) );
  XNOR U6262 ( .A(round_reg[1507]), .B(round_reg[1187]), .Z(n5258) );
  XOR U6263 ( .A(round_reg[227]), .B(n5259), .Z(n5257) );
  XOR U6264 ( .A(round_reg[867]), .B(round_reg[547]), .Z(n5259) );
  XOR U6265 ( .A(round_reg[1348]), .B(n1834), .Z(n1090) );
  XOR U6266 ( .A(n5117), .B(n5044), .Z(n1834) );
  XOR U6267 ( .A(n5261), .B(n5262), .Z(n5044) );
  XNOR U6268 ( .A(round_reg[323]), .B(round_reg[1283]), .Z(n5262) );
  XOR U6269 ( .A(round_reg[3]), .B(n5263), .Z(n5261) );
  XOR U6270 ( .A(round_reg[963]), .B(round_reg[643]), .Z(n5263) );
  XOR U6271 ( .A(n5264), .B(n5265), .Z(n5117) );
  XNOR U6272 ( .A(round_reg[132]), .B(round_reg[1092]), .Z(n5265) );
  XOR U6273 ( .A(round_reg[1412]), .B(n5266), .Z(n5264) );
  XOR U6274 ( .A(round_reg[772]), .B(round_reg[452]), .Z(n5266) );
  XOR U6275 ( .A(n5267), .B(n4701), .Z(out[1055]) );
  XNOR U6276 ( .A(round_reg[562]), .B(n4760), .Z(n4701) );
  XOR U6277 ( .A(n5268), .B(n4806), .Z(n4760) );
  XNOR U6278 ( .A(n5269), .B(n5270), .Z(n4806) );
  XNOR U6279 ( .A(round_reg[1586]), .B(round_reg[1266]), .Z(n5270) );
  XOR U6280 ( .A(round_reg[306]), .B(n5271), .Z(n5269) );
  XOR U6281 ( .A(round_reg[946]), .B(round_reg[626]), .Z(n5271) );
  ANDN U6282 ( .B(n1094), .A(n1092), .Z(n5267) );
  XOR U6283 ( .A(round_reg[162]), .B(n2210), .Z(n1092) );
  XOR U6284 ( .A(n4938), .B(n5272), .Z(n2210) );
  XOR U6285 ( .A(n5273), .B(n5274), .Z(n4938) );
  XNOR U6286 ( .A(round_reg[1506]), .B(round_reg[1186]), .Z(n5274) );
  XOR U6287 ( .A(round_reg[226]), .B(n5275), .Z(n5273) );
  XOR U6288 ( .A(round_reg[866]), .B(round_reg[546]), .Z(n5275) );
  XOR U6289 ( .A(round_reg[1347]), .B(n1837), .Z(n1094) );
  XOR U6290 ( .A(n5122), .B(n5089), .Z(n1837) );
  XOR U6291 ( .A(n5276), .B(n5277), .Z(n5089) );
  XNOR U6292 ( .A(round_reg[2]), .B(round_reg[1282]), .Z(n5277) );
  XOR U6293 ( .A(round_reg[322]), .B(n5278), .Z(n5276) );
  XOR U6294 ( .A(round_reg[962]), .B(round_reg[642]), .Z(n5278) );
  XOR U6295 ( .A(n5279), .B(n5280), .Z(n5122) );
  XNOR U6296 ( .A(round_reg[131]), .B(round_reg[1091]), .Z(n5280) );
  XOR U6297 ( .A(round_reg[1411]), .B(n5281), .Z(n5279) );
  XOR U6298 ( .A(round_reg[771]), .B(round_reg[451]), .Z(n5281) );
  XOR U6299 ( .A(n5282), .B(n4705), .Z(out[1054]) );
  XNOR U6300 ( .A(round_reg[561]), .B(n4803), .Z(n4705) );
  XOR U6301 ( .A(n5283), .B(n4810), .Z(n4803) );
  XNOR U6302 ( .A(n5284), .B(n5285), .Z(n4810) );
  XNOR U6303 ( .A(round_reg[1585]), .B(round_reg[1265]), .Z(n5285) );
  XOR U6304 ( .A(round_reg[305]), .B(n5286), .Z(n5284) );
  XOR U6305 ( .A(round_reg[945]), .B(round_reg[625]), .Z(n5286) );
  ANDN U6306 ( .B(n1098), .A(n1096), .Z(n5282) );
  XOR U6307 ( .A(round_reg[161]), .B(n2218), .Z(n1096) );
  XOR U6308 ( .A(n4941), .B(n5287), .Z(n2218) );
  XOR U6309 ( .A(n5288), .B(n5289), .Z(n4941) );
  XNOR U6310 ( .A(round_reg[1505]), .B(round_reg[1185]), .Z(n5289) );
  XOR U6311 ( .A(round_reg[225]), .B(n5290), .Z(n5288) );
  XOR U6312 ( .A(round_reg[865]), .B(round_reg[545]), .Z(n5290) );
  XOR U6313 ( .A(round_reg[1346]), .B(n1840), .Z(n1098) );
  XOR U6314 ( .A(n5127), .B(n5142), .Z(n1840) );
  XOR U6315 ( .A(n5291), .B(n5292), .Z(n5142) );
  XNOR U6316 ( .A(round_reg[1]), .B(round_reg[1281]), .Z(n5292) );
  XOR U6317 ( .A(round_reg[321]), .B(n5293), .Z(n5291) );
  XOR U6318 ( .A(round_reg[961]), .B(round_reg[641]), .Z(n5293) );
  XOR U6319 ( .A(n5294), .B(n5295), .Z(n5127) );
  XNOR U6320 ( .A(round_reg[130]), .B(round_reg[1090]), .Z(n5295) );
  XOR U6321 ( .A(round_reg[1410]), .B(n5296), .Z(n5294) );
  XOR U6322 ( .A(round_reg[770]), .B(round_reg[450]), .Z(n5296) );
  XOR U6323 ( .A(n5297), .B(n4709), .Z(out[1053]) );
  XNOR U6324 ( .A(round_reg[560]), .B(n4841), .Z(n4709) );
  XOR U6325 ( .A(n5298), .B(n4814), .Z(n4841) );
  XNOR U6326 ( .A(n5299), .B(n5300), .Z(n4814) );
  XNOR U6327 ( .A(round_reg[1584]), .B(round_reg[1264]), .Z(n5300) );
  XOR U6328 ( .A(round_reg[304]), .B(n5301), .Z(n5299) );
  XOR U6329 ( .A(round_reg[944]), .B(round_reg[624]), .Z(n5301) );
  AND U6330 ( .A(n1106), .B(n1104), .Z(n5297) );
  XNOR U6331 ( .A(round_reg[160]), .B(n2222), .Z(n1104) );
  XOR U6332 ( .A(n4944), .B(n5302), .Z(n2222) );
  XOR U6333 ( .A(n5303), .B(n5304), .Z(n4944) );
  XNOR U6334 ( .A(round_reg[1504]), .B(round_reg[1184]), .Z(n5304) );
  XOR U6335 ( .A(round_reg[224]), .B(n5305), .Z(n5303) );
  XOR U6336 ( .A(round_reg[864]), .B(round_reg[544]), .Z(n5305) );
  XOR U6337 ( .A(round_reg[1345]), .B(n1843), .Z(n1106) );
  XOR U6338 ( .A(n5132), .B(n5209), .Z(n1843) );
  XOR U6339 ( .A(n5306), .B(n5307), .Z(n5209) );
  XNOR U6340 ( .A(round_reg[1280]), .B(round_reg[0]), .Z(n5307) );
  XOR U6341 ( .A(round_reg[320]), .B(n5308), .Z(n5306) );
  XOR U6342 ( .A(round_reg[960]), .B(round_reg[640]), .Z(n5308) );
  XOR U6343 ( .A(n5309), .B(n5310), .Z(n5132) );
  XNOR U6344 ( .A(round_reg[129]), .B(round_reg[1089]), .Z(n5310) );
  XOR U6345 ( .A(round_reg[1409]), .B(n5311), .Z(n5309) );
  XOR U6346 ( .A(round_reg[769]), .B(round_reg[449]), .Z(n5311) );
  XOR U6347 ( .A(n5312), .B(n4713), .Z(out[1052]) );
  XNOR U6348 ( .A(round_reg[559]), .B(n4883), .Z(n4713) );
  XOR U6349 ( .A(n5313), .B(n4818), .Z(n4883) );
  XNOR U6350 ( .A(n5314), .B(n5315), .Z(n4818) );
  XNOR U6351 ( .A(round_reg[1583]), .B(round_reg[1263]), .Z(n5315) );
  XOR U6352 ( .A(round_reg[303]), .B(n5316), .Z(n5314) );
  XOR U6353 ( .A(round_reg[943]), .B(round_reg[623]), .Z(n5316) );
  AND U6354 ( .A(n1110), .B(n1108), .Z(n5312) );
  XNOR U6355 ( .A(round_reg[159]), .B(n2226), .Z(n1108) );
  XOR U6356 ( .A(n4947), .B(n5317), .Z(n2226) );
  XOR U6357 ( .A(n5318), .B(n5319), .Z(n4947) );
  XNOR U6358 ( .A(round_reg[1503]), .B(round_reg[1183]), .Z(n5319) );
  XOR U6359 ( .A(round_reg[223]), .B(n5320), .Z(n5318) );
  XOR U6360 ( .A(round_reg[863]), .B(round_reg[543]), .Z(n5320) );
  XOR U6361 ( .A(round_reg[1344]), .B(n1846), .Z(n1110) );
  XOR U6362 ( .A(n5137), .B(n5321), .Z(n1846) );
  XOR U6363 ( .A(n5322), .B(n5323), .Z(n5137) );
  XNOR U6364 ( .A(round_reg[128]), .B(round_reg[1088]), .Z(n5323) );
  XOR U6365 ( .A(round_reg[1408]), .B(n5324), .Z(n5322) );
  XOR U6366 ( .A(round_reg[768]), .B(round_reg[448]), .Z(n5324) );
  XOR U6367 ( .A(n5325), .B(n4720), .Z(out[1051]) );
  XNOR U6368 ( .A(round_reg[558]), .B(n4925), .Z(n4720) );
  XOR U6369 ( .A(n5326), .B(n4822), .Z(n4925) );
  XNOR U6370 ( .A(n5327), .B(n5328), .Z(n4822) );
  XNOR U6371 ( .A(round_reg[1582]), .B(round_reg[1262]), .Z(n5328) );
  XOR U6372 ( .A(round_reg[302]), .B(n5329), .Z(n5327) );
  XOR U6373 ( .A(round_reg[942]), .B(round_reg[622]), .Z(n5329) );
  ANDN U6374 ( .B(n1114), .A(n1112), .Z(n5325) );
  XOR U6375 ( .A(round_reg[158]), .B(n2230), .Z(n1112) );
  XOR U6376 ( .A(n4950), .B(n5330), .Z(n2230) );
  XOR U6377 ( .A(n5331), .B(n5332), .Z(n4950) );
  XNOR U6378 ( .A(round_reg[1502]), .B(round_reg[1182]), .Z(n5332) );
  XOR U6379 ( .A(round_reg[222]), .B(n5333), .Z(n5331) );
  XOR U6380 ( .A(round_reg[862]), .B(round_reg[542]), .Z(n5333) );
  XOR U6381 ( .A(round_reg[1407]), .B(n1849), .Z(n1114) );
  XOR U6382 ( .A(n5145), .B(n5334), .Z(n1849) );
  XOR U6383 ( .A(n5335), .B(n5336), .Z(n5145) );
  XNOR U6384 ( .A(round_reg[1471]), .B(round_reg[1151]), .Z(n5336) );
  XOR U6385 ( .A(round_reg[191]), .B(n5337), .Z(n5335) );
  XOR U6386 ( .A(round_reg[831]), .B(round_reg[511]), .Z(n5337) );
  XOR U6387 ( .A(n5338), .B(n4724), .Z(out[1050]) );
  XOR U6388 ( .A(round_reg[557]), .B(n2187), .Z(n4724) );
  XNOR U6389 ( .A(n5339), .B(n4826), .Z(n2187) );
  XNOR U6390 ( .A(n5340), .B(n5341), .Z(n4826) );
  XNOR U6391 ( .A(round_reg[1581]), .B(round_reg[1261]), .Z(n5341) );
  XOR U6392 ( .A(round_reg[301]), .B(n5342), .Z(n5340) );
  XOR U6393 ( .A(round_reg[941]), .B(round_reg[621]), .Z(n5342) );
  ANDN U6394 ( .B(n1118), .A(n1116), .Z(n5338) );
  XOR U6395 ( .A(round_reg[157]), .B(n2234), .Z(n1116) );
  XOR U6396 ( .A(n4953), .B(n5343), .Z(n2234) );
  XOR U6397 ( .A(n5344), .B(n5345), .Z(n4953) );
  XNOR U6398 ( .A(round_reg[1501]), .B(round_reg[1181]), .Z(n5345) );
  XOR U6399 ( .A(round_reg[221]), .B(n5346), .Z(n5344) );
  XOR U6400 ( .A(round_reg[861]), .B(round_reg[541]), .Z(n5346) );
  XOR U6401 ( .A(round_reg[1406]), .B(n1852), .Z(n1118) );
  XOR U6402 ( .A(n5150), .B(n5347), .Z(n1852) );
  XOR U6403 ( .A(n5348), .B(n5349), .Z(n5150) );
  XNOR U6404 ( .A(round_reg[1470]), .B(round_reg[1150]), .Z(n5349) );
  XOR U6405 ( .A(round_reg[190]), .B(n5350), .Z(n5348) );
  XOR U6406 ( .A(round_reg[830]), .B(round_reg[510]), .Z(n5350) );
  XOR U6407 ( .A(n5351), .B(n3469), .Z(out[104]) );
  IV U6408 ( .A(n3571), .Z(n3469) );
  XNOR U6409 ( .A(round_reg[639]), .B(n2313), .Z(n3571) );
  XNOR U6410 ( .A(n5321), .B(n5352), .Z(n2313) );
  XOR U6411 ( .A(n5353), .B(n5354), .Z(n5321) );
  XNOR U6412 ( .A(round_reg[1343]), .B(round_reg[1023]), .Z(n5354) );
  XOR U6413 ( .A(round_reg[383]), .B(n5355), .Z(n5353) );
  XOR U6414 ( .A(round_reg[703]), .B(round_reg[63]), .Z(n5355) );
  AND U6415 ( .A(n3083), .B(n3085), .Z(n5351) );
  XOR U6416 ( .A(round_reg[1450]), .B(n2178), .Z(n3085) );
  XOR U6417 ( .A(n4905), .B(n5356), .Z(n2178) );
  XOR U6418 ( .A(n5357), .B(n5358), .Z(n4905) );
  XNOR U6419 ( .A(round_reg[1514]), .B(round_reg[1194]), .Z(n5358) );
  XOR U6420 ( .A(round_reg[234]), .B(n5359), .Z(n5357) );
  XOR U6421 ( .A(round_reg[874]), .B(round_reg[554]), .Z(n5359) );
  XNOR U6422 ( .A(round_reg[230]), .B(n2219), .Z(n3083) );
  XOR U6423 ( .A(n5360), .B(n4728), .Z(out[1049]) );
  XOR U6424 ( .A(round_reg[556]), .B(n2191), .Z(n4728) );
  XNOR U6425 ( .A(n5361), .B(n4830), .Z(n2191) );
  XNOR U6426 ( .A(n5362), .B(n5363), .Z(n4830) );
  XNOR U6427 ( .A(round_reg[1580]), .B(round_reg[1260]), .Z(n5363) );
  XOR U6428 ( .A(round_reg[300]), .B(n5364), .Z(n5362) );
  XOR U6429 ( .A(round_reg[940]), .B(round_reg[620]), .Z(n5364) );
  ANDN U6430 ( .B(n1122), .A(n1120), .Z(n5360) );
  XOR U6431 ( .A(round_reg[156]), .B(n2238), .Z(n1120) );
  XOR U6432 ( .A(n4956), .B(n5365), .Z(n2238) );
  XOR U6433 ( .A(n5366), .B(n5367), .Z(n4956) );
  XNOR U6434 ( .A(round_reg[1500]), .B(round_reg[1180]), .Z(n5367) );
  XOR U6435 ( .A(round_reg[220]), .B(n5368), .Z(n5366) );
  XOR U6436 ( .A(round_reg[860]), .B(round_reg[540]), .Z(n5368) );
  XOR U6437 ( .A(round_reg[1405]), .B(n1855), .Z(n1122) );
  XOR U6438 ( .A(n5369), .B(n5370), .Z(n1855) );
  XOR U6439 ( .A(n5371), .B(n4732), .Z(out[1048]) );
  XOR U6440 ( .A(round_reg[555]), .B(n2195), .Z(n4732) );
  XNOR U6441 ( .A(n5372), .B(n4834), .Z(n2195) );
  XNOR U6442 ( .A(n5373), .B(n5374), .Z(n4834) );
  XNOR U6443 ( .A(round_reg[1579]), .B(round_reg[1259]), .Z(n5374) );
  XOR U6444 ( .A(round_reg[299]), .B(n5375), .Z(n5373) );
  XOR U6445 ( .A(round_reg[939]), .B(round_reg[619]), .Z(n5375) );
  ANDN U6446 ( .B(n1126), .A(n1124), .Z(n5371) );
  XOR U6447 ( .A(round_reg[155]), .B(n2242), .Z(n1124) );
  XOR U6448 ( .A(n4960), .B(n5376), .Z(n2242) );
  XOR U6449 ( .A(n5377), .B(n5378), .Z(n4960) );
  XNOR U6450 ( .A(round_reg[1499]), .B(round_reg[1179]), .Z(n5378) );
  XOR U6451 ( .A(round_reg[219]), .B(n5379), .Z(n5377) );
  XOR U6452 ( .A(round_reg[859]), .B(round_reg[539]), .Z(n5379) );
  XOR U6453 ( .A(round_reg[1404]), .B(n1862), .Z(n1126) );
  XOR U6454 ( .A(n5156), .B(n5380), .Z(n1862) );
  XOR U6455 ( .A(n5381), .B(n5382), .Z(n5156) );
  XNOR U6456 ( .A(round_reg[1468]), .B(round_reg[1148]), .Z(n5382) );
  XOR U6457 ( .A(round_reg[188]), .B(n5383), .Z(n5381) );
  XOR U6458 ( .A(round_reg[828]), .B(round_reg[508]), .Z(n5383) );
  XOR U6459 ( .A(n5384), .B(n4736), .Z(out[1047]) );
  XOR U6460 ( .A(round_reg[554]), .B(n2199), .Z(n4736) );
  XNOR U6461 ( .A(n5385), .B(n5386), .Z(n2199) );
  ANDN U6462 ( .B(n1130), .A(n1128), .Z(n5384) );
  XOR U6463 ( .A(round_reg[154]), .B(n2246), .Z(n1128) );
  XOR U6464 ( .A(n4963), .B(n5387), .Z(n2246) );
  XOR U6465 ( .A(n5388), .B(n5389), .Z(n4963) );
  XNOR U6466 ( .A(round_reg[1498]), .B(round_reg[1178]), .Z(n5389) );
  XOR U6467 ( .A(round_reg[218]), .B(n5390), .Z(n5388) );
  XOR U6468 ( .A(round_reg[858]), .B(round_reg[538]), .Z(n5390) );
  XOR U6469 ( .A(round_reg[1403]), .B(n1865), .Z(n1130) );
  XOR U6470 ( .A(n4844), .B(n5161), .Z(n1865) );
  XOR U6471 ( .A(n5391), .B(n5392), .Z(n5161) );
  XNOR U6472 ( .A(round_reg[1467]), .B(round_reg[1147]), .Z(n5392) );
  XOR U6473 ( .A(round_reg[187]), .B(n5393), .Z(n5391) );
  XOR U6474 ( .A(round_reg[827]), .B(round_reg[507]), .Z(n5393) );
  XOR U6475 ( .A(n5394), .B(n5395), .Z(n4844) );
  XNOR U6476 ( .A(round_reg[1338]), .B(round_reg[1018]), .Z(n5395) );
  XOR U6477 ( .A(round_reg[378]), .B(n5396), .Z(n5394) );
  XOR U6478 ( .A(round_reg[698]), .B(round_reg[58]), .Z(n5396) );
  XOR U6479 ( .A(n5397), .B(n4740), .Z(out[1046]) );
  XOR U6480 ( .A(round_reg[553]), .B(n2203), .Z(n4740) );
  XNOR U6481 ( .A(n5398), .B(n5399), .Z(n2203) );
  ANDN U6482 ( .B(n1134), .A(n1132), .Z(n5397) );
  XOR U6483 ( .A(round_reg[153]), .B(n2250), .Z(n1132) );
  XOR U6484 ( .A(n4966), .B(n5400), .Z(n2250) );
  XOR U6485 ( .A(n5401), .B(n5402), .Z(n4966) );
  XNOR U6486 ( .A(round_reg[1497]), .B(round_reg[1177]), .Z(n5402) );
  XOR U6487 ( .A(round_reg[217]), .B(n5403), .Z(n5401) );
  XOR U6488 ( .A(round_reg[857]), .B(round_reg[537]), .Z(n5403) );
  XOR U6489 ( .A(round_reg[1402]), .B(n1868), .Z(n1134) );
  XOR U6490 ( .A(n4848), .B(n5166), .Z(n1868) );
  XOR U6491 ( .A(n5404), .B(n5405), .Z(n5166) );
  XNOR U6492 ( .A(round_reg[1466]), .B(round_reg[1146]), .Z(n5405) );
  XOR U6493 ( .A(round_reg[186]), .B(n5406), .Z(n5404) );
  XOR U6494 ( .A(round_reg[826]), .B(round_reg[506]), .Z(n5406) );
  XOR U6495 ( .A(n5407), .B(n5408), .Z(n4848) );
  XNOR U6496 ( .A(round_reg[1337]), .B(round_reg[1017]), .Z(n5408) );
  XOR U6497 ( .A(round_reg[377]), .B(n5409), .Z(n5407) );
  XOR U6498 ( .A(round_reg[697]), .B(round_reg[57]), .Z(n5409) );
  XOR U6499 ( .A(n5410), .B(n4744), .Z(out[1045]) );
  XOR U6500 ( .A(round_reg[552]), .B(n2207), .Z(n4744) );
  XNOR U6501 ( .A(n5411), .B(n5412), .Z(n2207) );
  ANDN U6502 ( .B(n1138), .A(n1136), .Z(n5410) );
  XOR U6503 ( .A(round_reg[152]), .B(n2254), .Z(n1136) );
  XOR U6504 ( .A(n4969), .B(n5413), .Z(n2254) );
  XOR U6505 ( .A(n5414), .B(n5415), .Z(n4969) );
  XNOR U6506 ( .A(round_reg[1496]), .B(round_reg[1176]), .Z(n5415) );
  XOR U6507 ( .A(round_reg[216]), .B(n5416), .Z(n5414) );
  XOR U6508 ( .A(round_reg[856]), .B(round_reg[536]), .Z(n5416) );
  XOR U6509 ( .A(round_reg[1401]), .B(n1871), .Z(n1138) );
  XOR U6510 ( .A(n5171), .B(n4851), .Z(n1871) );
  XOR U6511 ( .A(n5417), .B(n5418), .Z(n4851) );
  XNOR U6512 ( .A(round_reg[1336]), .B(round_reg[1016]), .Z(n5418) );
  XOR U6513 ( .A(round_reg[376]), .B(n5419), .Z(n5417) );
  XOR U6514 ( .A(round_reg[696]), .B(round_reg[56]), .Z(n5419) );
  XOR U6515 ( .A(n5420), .B(n5421), .Z(n5171) );
  XNOR U6516 ( .A(round_reg[1465]), .B(round_reg[1145]), .Z(n5421) );
  XOR U6517 ( .A(round_reg[185]), .B(n5422), .Z(n5420) );
  XOR U6518 ( .A(round_reg[825]), .B(round_reg[505]), .Z(n5422) );
  XOR U6519 ( .A(n5423), .B(n4748), .Z(out[1044]) );
  XOR U6520 ( .A(round_reg[551]), .B(n2211), .Z(n4748) );
  XNOR U6521 ( .A(n5424), .B(n5425), .Z(n2211) );
  ANDN U6522 ( .B(n1142), .A(n1140), .Z(n5423) );
  XOR U6523 ( .A(round_reg[151]), .B(n2262), .Z(n1140) );
  XOR U6524 ( .A(n4972), .B(n5426), .Z(n2262) );
  XOR U6525 ( .A(n5427), .B(n5428), .Z(n4972) );
  XNOR U6526 ( .A(round_reg[1495]), .B(round_reg[1175]), .Z(n5428) );
  XOR U6527 ( .A(round_reg[215]), .B(n5429), .Z(n5427) );
  XOR U6528 ( .A(round_reg[855]), .B(round_reg[535]), .Z(n5429) );
  XOR U6529 ( .A(round_reg[1400]), .B(n1874), .Z(n1142) );
  XOR U6530 ( .A(n5182), .B(n4855), .Z(n1874) );
  XOR U6531 ( .A(n5430), .B(n5431), .Z(n4855) );
  XNOR U6532 ( .A(round_reg[1335]), .B(round_reg[1015]), .Z(n5431) );
  XOR U6533 ( .A(round_reg[375]), .B(n5432), .Z(n5430) );
  XOR U6534 ( .A(round_reg[695]), .B(round_reg[55]), .Z(n5432) );
  XOR U6535 ( .A(n5433), .B(n5434), .Z(n5182) );
  XNOR U6536 ( .A(round_reg[1464]), .B(round_reg[1144]), .Z(n5434) );
  XOR U6537 ( .A(round_reg[184]), .B(n5435), .Z(n5433) );
  XOR U6538 ( .A(round_reg[824]), .B(round_reg[504]), .Z(n5435) );
  XOR U6539 ( .A(n5436), .B(n4752), .Z(out[1043]) );
  XOR U6540 ( .A(round_reg[550]), .B(n2219), .Z(n4752) );
  XNOR U6541 ( .A(n5437), .B(n5438), .Z(n2219) );
  ANDN U6542 ( .B(n1150), .A(n1148), .Z(n5436) );
  XOR U6543 ( .A(round_reg[150]), .B(n2266), .Z(n1148) );
  XOR U6544 ( .A(n4975), .B(n5439), .Z(n2266) );
  XOR U6545 ( .A(n5440), .B(n5441), .Z(n4975) );
  XNOR U6546 ( .A(round_reg[1494]), .B(round_reg[1174]), .Z(n5441) );
  XOR U6547 ( .A(round_reg[214]), .B(n5442), .Z(n5440) );
  XOR U6548 ( .A(round_reg[854]), .B(round_reg[534]), .Z(n5442) );
  XOR U6549 ( .A(round_reg[1399]), .B(n1877), .Z(n1150) );
  XOR U6550 ( .A(n5193), .B(n4859), .Z(n1877) );
  XOR U6551 ( .A(n5443), .B(n5444), .Z(n4859) );
  XNOR U6552 ( .A(round_reg[1334]), .B(round_reg[1014]), .Z(n5444) );
  XOR U6553 ( .A(round_reg[374]), .B(n5445), .Z(n5443) );
  XOR U6554 ( .A(round_reg[694]), .B(round_reg[54]), .Z(n5445) );
  XOR U6555 ( .A(n5446), .B(n5447), .Z(n5193) );
  XNOR U6556 ( .A(round_reg[1463]), .B(round_reg[1143]), .Z(n5447) );
  XOR U6557 ( .A(round_reg[183]), .B(n5448), .Z(n5446) );
  XOR U6558 ( .A(round_reg[823]), .B(round_reg[503]), .Z(n5448) );
  XOR U6559 ( .A(n5449), .B(n4756), .Z(out[1042]) );
  XOR U6560 ( .A(round_reg[549]), .B(n2223), .Z(n4756) );
  ANDN U6561 ( .B(n1154), .A(n1152), .Z(n5449) );
  XOR U6562 ( .A(round_reg[149]), .B(n2270), .Z(n1152) );
  XOR U6563 ( .A(n4978), .B(n5450), .Z(n2270) );
  XOR U6564 ( .A(n5451), .B(n5452), .Z(n4978) );
  XNOR U6565 ( .A(round_reg[1493]), .B(round_reg[1173]), .Z(n5452) );
  XOR U6566 ( .A(round_reg[213]), .B(n5453), .Z(n5451) );
  XOR U6567 ( .A(round_reg[853]), .B(round_reg[533]), .Z(n5453) );
  XOR U6568 ( .A(round_reg[1398]), .B(n1880), .Z(n1154) );
  XOR U6569 ( .A(n5198), .B(n4863), .Z(n1880) );
  XOR U6570 ( .A(n5454), .B(n5455), .Z(n4863) );
  XNOR U6571 ( .A(round_reg[1333]), .B(round_reg[1013]), .Z(n5455) );
  XOR U6572 ( .A(round_reg[373]), .B(n5456), .Z(n5454) );
  XOR U6573 ( .A(round_reg[693]), .B(round_reg[53]), .Z(n5456) );
  XOR U6574 ( .A(n5457), .B(n5458), .Z(n5198) );
  XNOR U6575 ( .A(round_reg[1462]), .B(round_reg[1142]), .Z(n5458) );
  XOR U6576 ( .A(round_reg[182]), .B(n5459), .Z(n5457) );
  XOR U6577 ( .A(round_reg[822]), .B(round_reg[502]), .Z(n5459) );
  XOR U6578 ( .A(n5460), .B(n4764), .Z(out[1041]) );
  XOR U6579 ( .A(round_reg[548]), .B(n2227), .Z(n4764) );
  ANDN U6580 ( .B(n1158), .A(n1156), .Z(n5460) );
  XOR U6581 ( .A(round_reg[148]), .B(n2274), .Z(n1156) );
  XOR U6582 ( .A(n4665), .B(n4981), .Z(n2274) );
  XOR U6583 ( .A(n5461), .B(n5462), .Z(n4981) );
  XNOR U6584 ( .A(round_reg[1492]), .B(round_reg[1172]), .Z(n5462) );
  XOR U6585 ( .A(round_reg[212]), .B(n5463), .Z(n5461) );
  XOR U6586 ( .A(round_reg[852]), .B(round_reg[532]), .Z(n5463) );
  XOR U6587 ( .A(n5464), .B(n5465), .Z(n4665) );
  XNOR U6588 ( .A(round_reg[1363]), .B(round_reg[1043]), .Z(n5465) );
  XOR U6589 ( .A(round_reg[403]), .B(n5466), .Z(n5464) );
  XOR U6590 ( .A(round_reg[83]), .B(round_reg[723]), .Z(n5466) );
  XOR U6591 ( .A(round_reg[1397]), .B(n1883), .Z(n1158) );
  XOR U6592 ( .A(n5212), .B(n4867), .Z(n1883) );
  XOR U6593 ( .A(n5467), .B(n5468), .Z(n4867) );
  XNOR U6594 ( .A(round_reg[1332]), .B(round_reg[1012]), .Z(n5468) );
  XOR U6595 ( .A(round_reg[372]), .B(n5469), .Z(n5467) );
  XOR U6596 ( .A(round_reg[692]), .B(round_reg[52]), .Z(n5469) );
  XOR U6597 ( .A(n5470), .B(n5471), .Z(n5212) );
  XNOR U6598 ( .A(round_reg[1461]), .B(round_reg[1141]), .Z(n5471) );
  XOR U6599 ( .A(round_reg[181]), .B(n5472), .Z(n5470) );
  XOR U6600 ( .A(round_reg[821]), .B(round_reg[501]), .Z(n5472) );
  XOR U6601 ( .A(n5473), .B(n4768), .Z(out[1040]) );
  XOR U6602 ( .A(round_reg[547]), .B(n2231), .Z(n4768) );
  ANDN U6603 ( .B(n1162), .A(n1160), .Z(n5473) );
  XOR U6604 ( .A(round_reg[147]), .B(n2278), .Z(n1160) );
  XOR U6605 ( .A(n4669), .B(n4984), .Z(n2278) );
  XOR U6606 ( .A(n5474), .B(n5475), .Z(n4984) );
  XNOR U6607 ( .A(round_reg[1491]), .B(round_reg[1171]), .Z(n5475) );
  XOR U6608 ( .A(round_reg[211]), .B(n5476), .Z(n5474) );
  XOR U6609 ( .A(round_reg[851]), .B(round_reg[531]), .Z(n5476) );
  XOR U6610 ( .A(n5477), .B(n5478), .Z(n4669) );
  XNOR U6611 ( .A(round_reg[1362]), .B(round_reg[1042]), .Z(n5478) );
  XOR U6612 ( .A(round_reg[402]), .B(n5479), .Z(n5477) );
  XOR U6613 ( .A(round_reg[82]), .B(round_reg[722]), .Z(n5479) );
  XOR U6614 ( .A(round_reg[1396]), .B(n1886), .Z(n1162) );
  XOR U6615 ( .A(n5223), .B(n4871), .Z(n1886) );
  XOR U6616 ( .A(n5480), .B(n5481), .Z(n4871) );
  XNOR U6617 ( .A(round_reg[1331]), .B(round_reg[1011]), .Z(n5481) );
  XOR U6618 ( .A(round_reg[371]), .B(n5482), .Z(n5480) );
  XOR U6619 ( .A(round_reg[691]), .B(round_reg[51]), .Z(n5482) );
  XOR U6620 ( .A(n5483), .B(n5484), .Z(n5223) );
  XNOR U6621 ( .A(round_reg[1460]), .B(round_reg[1140]), .Z(n5484) );
  XOR U6622 ( .A(round_reg[180]), .B(n5485), .Z(n5483) );
  XOR U6623 ( .A(round_reg[820]), .B(round_reg[500]), .Z(n5485) );
  XOR U6624 ( .A(n5486), .B(n3471), .Z(out[103]) );
  IV U6625 ( .A(n3573), .Z(n3471) );
  XNOR U6626 ( .A(round_reg[638]), .B(n2317), .Z(n3573) );
  XNOR U6627 ( .A(n5334), .B(n5487), .Z(n2317) );
  XOR U6628 ( .A(n5488), .B(n5489), .Z(n5334) );
  XNOR U6629 ( .A(round_reg[1342]), .B(round_reg[1022]), .Z(n5489) );
  XOR U6630 ( .A(round_reg[382]), .B(n5490), .Z(n5488) );
  XOR U6631 ( .A(round_reg[702]), .B(round_reg[62]), .Z(n5490) );
  AND U6632 ( .A(n3108), .B(n3110), .Z(n5486) );
  XOR U6633 ( .A(round_reg[1449]), .B(n2182), .Z(n3110) );
  XOR U6634 ( .A(n4909), .B(n5491), .Z(n2182) );
  XOR U6635 ( .A(n5492), .B(n5493), .Z(n4909) );
  XNOR U6636 ( .A(round_reg[1513]), .B(round_reg[1193]), .Z(n5493) );
  XOR U6637 ( .A(round_reg[233]), .B(n5494), .Z(n5492) );
  XOR U6638 ( .A(round_reg[873]), .B(round_reg[553]), .Z(n5494) );
  XNOR U6639 ( .A(round_reg[229]), .B(n2223), .Z(n3108) );
  XNOR U6640 ( .A(n5495), .B(n5496), .Z(n2223) );
  XOR U6641 ( .A(n5497), .B(n4772), .Z(out[1039]) );
  XOR U6642 ( .A(round_reg[546]), .B(n2235), .Z(n4772) );
  AND U6643 ( .A(n1166), .B(n1164), .Z(n5497) );
  XNOR U6644 ( .A(round_reg[146]), .B(n2282), .Z(n1164) );
  XOR U6645 ( .A(n4676), .B(n4987), .Z(n2282) );
  XOR U6646 ( .A(n5498), .B(n5499), .Z(n4987) );
  XNOR U6647 ( .A(round_reg[1490]), .B(round_reg[1170]), .Z(n5499) );
  XOR U6648 ( .A(round_reg[210]), .B(n5500), .Z(n5498) );
  XOR U6649 ( .A(round_reg[850]), .B(round_reg[530]), .Z(n5500) );
  XOR U6650 ( .A(n5501), .B(n5502), .Z(n4676) );
  XNOR U6651 ( .A(round_reg[1361]), .B(round_reg[1041]), .Z(n5502) );
  XOR U6652 ( .A(round_reg[401]), .B(n5503), .Z(n5501) );
  XOR U6653 ( .A(round_reg[81]), .B(round_reg[721]), .Z(n5503) );
  XOR U6654 ( .A(round_reg[1395]), .B(n1889), .Z(n1166) );
  XOR U6655 ( .A(n5238), .B(n4875), .Z(n1889) );
  XOR U6656 ( .A(n5504), .B(n5505), .Z(n4875) );
  XNOR U6657 ( .A(round_reg[1330]), .B(round_reg[1010]), .Z(n5505) );
  XOR U6658 ( .A(round_reg[370]), .B(n5506), .Z(n5504) );
  XOR U6659 ( .A(round_reg[690]), .B(round_reg[50]), .Z(n5506) );
  XOR U6660 ( .A(n5507), .B(n5508), .Z(n5238) );
  XNOR U6661 ( .A(round_reg[1459]), .B(round_reg[1139]), .Z(n5508) );
  XOR U6662 ( .A(round_reg[179]), .B(n5509), .Z(n5507) );
  XOR U6663 ( .A(round_reg[819]), .B(round_reg[499]), .Z(n5509) );
  XOR U6664 ( .A(n5510), .B(n4776), .Z(out[1038]) );
  XOR U6665 ( .A(round_reg[545]), .B(n2239), .Z(n4776) );
  XOR U6666 ( .A(n5511), .B(n5512), .Z(n2239) );
  ANDN U6667 ( .B(n1170), .A(n1168), .Z(n5510) );
  XOR U6668 ( .A(round_reg[145]), .B(n2286), .Z(n1168) );
  XOR U6669 ( .A(n4680), .B(n4991), .Z(n2286) );
  XOR U6670 ( .A(n5513), .B(n5514), .Z(n4991) );
  XNOR U6671 ( .A(round_reg[1489]), .B(round_reg[1169]), .Z(n5514) );
  XOR U6672 ( .A(round_reg[209]), .B(n5515), .Z(n5513) );
  XOR U6673 ( .A(round_reg[849]), .B(round_reg[529]), .Z(n5515) );
  XOR U6674 ( .A(n5516), .B(n5517), .Z(n4680) );
  XNOR U6675 ( .A(round_reg[1360]), .B(round_reg[1040]), .Z(n5517) );
  XOR U6676 ( .A(round_reg[400]), .B(n5518), .Z(n5516) );
  XOR U6677 ( .A(round_reg[80]), .B(round_reg[720]), .Z(n5518) );
  XOR U6678 ( .A(round_reg[1394]), .B(n1896), .Z(n1170) );
  XOR U6679 ( .A(n5253), .B(n4879), .Z(n1896) );
  XOR U6680 ( .A(n5519), .B(n5520), .Z(n4879) );
  XNOR U6681 ( .A(round_reg[1329]), .B(round_reg[1009]), .Z(n5520) );
  XOR U6682 ( .A(round_reg[369]), .B(n5521), .Z(n5519) );
  XOR U6683 ( .A(round_reg[689]), .B(round_reg[49]), .Z(n5521) );
  XOR U6684 ( .A(n5522), .B(n5523), .Z(n5253) );
  XNOR U6685 ( .A(round_reg[1458]), .B(round_reg[1138]), .Z(n5523) );
  XOR U6686 ( .A(round_reg[178]), .B(n5524), .Z(n5522) );
  XOR U6687 ( .A(round_reg[818]), .B(round_reg[498]), .Z(n5524) );
  XOR U6688 ( .A(n5525), .B(n4780), .Z(out[1037]) );
  XNOR U6689 ( .A(round_reg[544]), .B(n2243), .Z(n4780) );
  ANDN U6690 ( .B(n1174), .A(n1172), .Z(n5525) );
  XOR U6691 ( .A(round_reg[144]), .B(n2290), .Z(n1172) );
  XNOR U6692 ( .A(n4684), .B(n4995), .Z(n2290) );
  XNOR U6693 ( .A(n5528), .B(n5529), .Z(n4995) );
  XNOR U6694 ( .A(round_reg[1488]), .B(round_reg[1168]), .Z(n5529) );
  XOR U6695 ( .A(round_reg[208]), .B(n5530), .Z(n5528) );
  XOR U6696 ( .A(round_reg[848]), .B(round_reg[528]), .Z(n5530) );
  XOR U6697 ( .A(n5531), .B(n5532), .Z(n4684) );
  XNOR U6698 ( .A(round_reg[1359]), .B(round_reg[1039]), .Z(n5532) );
  XOR U6699 ( .A(round_reg[399]), .B(n5533), .Z(n5531) );
  XOR U6700 ( .A(round_reg[79]), .B(round_reg[719]), .Z(n5533) );
  XOR U6701 ( .A(round_reg[1393]), .B(n1899), .Z(n1174) );
  XOR U6702 ( .A(n5268), .B(n4885), .Z(n1899) );
  XOR U6703 ( .A(n5534), .B(n5535), .Z(n4885) );
  XNOR U6704 ( .A(round_reg[1328]), .B(round_reg[1008]), .Z(n5535) );
  XOR U6705 ( .A(round_reg[368]), .B(n5536), .Z(n5534) );
  XOR U6706 ( .A(round_reg[688]), .B(round_reg[48]), .Z(n5536) );
  XOR U6707 ( .A(n5537), .B(n5538), .Z(n5268) );
  XNOR U6708 ( .A(round_reg[1457]), .B(round_reg[1137]), .Z(n5538) );
  XOR U6709 ( .A(round_reg[177]), .B(n5539), .Z(n5537) );
  XOR U6710 ( .A(round_reg[817]), .B(round_reg[497]), .Z(n5539) );
  XOR U6711 ( .A(n5540), .B(n4784), .Z(out[1036]) );
  XNOR U6712 ( .A(round_reg[543]), .B(n2247), .Z(n4784) );
  ANDN U6713 ( .B(n1178), .A(n1176), .Z(n5540) );
  XOR U6714 ( .A(round_reg[143]), .B(n2294), .Z(n1176) );
  XOR U6715 ( .A(n4688), .B(n4997), .Z(n2294) );
  XOR U6716 ( .A(n5543), .B(n5544), .Z(n4997) );
  XNOR U6717 ( .A(round_reg[1487]), .B(round_reg[1167]), .Z(n5544) );
  XOR U6718 ( .A(round_reg[207]), .B(n5545), .Z(n5543) );
  XOR U6719 ( .A(round_reg[847]), .B(round_reg[527]), .Z(n5545) );
  XOR U6720 ( .A(n5546), .B(n5547), .Z(n4688) );
  XNOR U6721 ( .A(round_reg[1358]), .B(round_reg[1038]), .Z(n5547) );
  XOR U6722 ( .A(round_reg[398]), .B(n5548), .Z(n5546) );
  XOR U6723 ( .A(round_reg[78]), .B(round_reg[718]), .Z(n5548) );
  XOR U6724 ( .A(round_reg[1392]), .B(n1902), .Z(n1178) );
  XOR U6725 ( .A(n5283), .B(n4889), .Z(n1902) );
  XOR U6726 ( .A(n5549), .B(n5550), .Z(n4889) );
  XNOR U6727 ( .A(round_reg[1327]), .B(round_reg[1007]), .Z(n5550) );
  XOR U6728 ( .A(round_reg[367]), .B(n5551), .Z(n5549) );
  XOR U6729 ( .A(round_reg[687]), .B(round_reg[47]), .Z(n5551) );
  XOR U6730 ( .A(n5552), .B(n5553), .Z(n5283) );
  XNOR U6731 ( .A(round_reg[1456]), .B(round_reg[1136]), .Z(n5553) );
  XOR U6732 ( .A(round_reg[176]), .B(n5554), .Z(n5552) );
  XOR U6733 ( .A(round_reg[816]), .B(round_reg[496]), .Z(n5554) );
  XOR U6734 ( .A(n5555), .B(n4788), .Z(out[1035]) );
  XNOR U6735 ( .A(round_reg[542]), .B(n2251), .Z(n4788) );
  ANDN U6736 ( .B(n1182), .A(n1180), .Z(n5555) );
  XOR U6737 ( .A(round_reg[142]), .B(n2298), .Z(n1180) );
  XOR U6738 ( .A(n4691), .B(n5000), .Z(n2298) );
  XOR U6739 ( .A(n5558), .B(n5559), .Z(n5000) );
  XNOR U6740 ( .A(round_reg[1486]), .B(round_reg[1166]), .Z(n5559) );
  XOR U6741 ( .A(round_reg[206]), .B(n5560), .Z(n5558) );
  XOR U6742 ( .A(round_reg[846]), .B(round_reg[526]), .Z(n5560) );
  XOR U6743 ( .A(n5561), .B(n5562), .Z(n4691) );
  XNOR U6744 ( .A(round_reg[1357]), .B(round_reg[1037]), .Z(n5562) );
  XOR U6745 ( .A(round_reg[397]), .B(n5563), .Z(n5561) );
  XOR U6746 ( .A(round_reg[77]), .B(round_reg[717]), .Z(n5563) );
  XOR U6747 ( .A(round_reg[1391]), .B(n1905), .Z(n1182) );
  XOR U6748 ( .A(n5298), .B(n4893), .Z(n1905) );
  XOR U6749 ( .A(n5564), .B(n5565), .Z(n4893) );
  XNOR U6750 ( .A(round_reg[1326]), .B(round_reg[1006]), .Z(n5565) );
  XOR U6751 ( .A(round_reg[366]), .B(n5566), .Z(n5564) );
  XOR U6752 ( .A(round_reg[686]), .B(round_reg[46]), .Z(n5566) );
  XOR U6753 ( .A(n5567), .B(n5568), .Z(n5298) );
  XNOR U6754 ( .A(round_reg[1455]), .B(round_reg[1135]), .Z(n5568) );
  XOR U6755 ( .A(round_reg[175]), .B(n5569), .Z(n5567) );
  XOR U6756 ( .A(round_reg[815]), .B(round_reg[495]), .Z(n5569) );
  XOR U6757 ( .A(n5570), .B(n4792), .Z(out[1034]) );
  XNOR U6758 ( .A(round_reg[541]), .B(n2255), .Z(n4792) );
  ANDN U6759 ( .B(n1186), .A(n1184), .Z(n5570) );
  XOR U6760 ( .A(round_reg[141]), .B(n2306), .Z(n1184) );
  XOR U6761 ( .A(n4695), .B(n5003), .Z(n2306) );
  XOR U6762 ( .A(n5573), .B(n5574), .Z(n5003) );
  XNOR U6763 ( .A(round_reg[1485]), .B(round_reg[1165]), .Z(n5574) );
  XOR U6764 ( .A(round_reg[205]), .B(n5575), .Z(n5573) );
  XOR U6765 ( .A(round_reg[845]), .B(round_reg[525]), .Z(n5575) );
  XOR U6766 ( .A(n5576), .B(n5577), .Z(n4695) );
  XNOR U6767 ( .A(round_reg[1356]), .B(round_reg[1036]), .Z(n5577) );
  XOR U6768 ( .A(round_reg[396]), .B(n5578), .Z(n5576) );
  XOR U6769 ( .A(round_reg[76]), .B(round_reg[716]), .Z(n5578) );
  XOR U6770 ( .A(round_reg[1390]), .B(n1908), .Z(n1186) );
  XOR U6771 ( .A(n5313), .B(n4897), .Z(n1908) );
  XOR U6772 ( .A(n5579), .B(n5580), .Z(n4897) );
  XNOR U6773 ( .A(round_reg[1325]), .B(round_reg[1005]), .Z(n5580) );
  XOR U6774 ( .A(round_reg[365]), .B(n5581), .Z(n5579) );
  XOR U6775 ( .A(round_reg[685]), .B(round_reg[45]), .Z(n5581) );
  XOR U6776 ( .A(n5582), .B(n5583), .Z(n5313) );
  XNOR U6777 ( .A(round_reg[1454]), .B(round_reg[1134]), .Z(n5583) );
  XOR U6778 ( .A(round_reg[174]), .B(n5584), .Z(n5582) );
  XOR U6779 ( .A(round_reg[814]), .B(round_reg[494]), .Z(n5584) );
  XOR U6780 ( .A(n5585), .B(n4796), .Z(out[1033]) );
  XNOR U6781 ( .A(round_reg[540]), .B(n2263), .Z(n4796) );
  ANDN U6782 ( .B(n1194), .A(n1192), .Z(n5585) );
  XOR U6783 ( .A(round_reg[140]), .B(n2310), .Z(n1192) );
  XOR U6784 ( .A(n4699), .B(n5006), .Z(n2310) );
  XOR U6785 ( .A(n5588), .B(n5589), .Z(n5006) );
  XNOR U6786 ( .A(round_reg[1484]), .B(round_reg[1164]), .Z(n5589) );
  XOR U6787 ( .A(round_reg[204]), .B(n5590), .Z(n5588) );
  XOR U6788 ( .A(round_reg[844]), .B(round_reg[524]), .Z(n5590) );
  XOR U6789 ( .A(n5591), .B(n5592), .Z(n4699) );
  XNOR U6790 ( .A(round_reg[1355]), .B(round_reg[1035]), .Z(n5592) );
  XOR U6791 ( .A(round_reg[395]), .B(n5593), .Z(n5591) );
  XOR U6792 ( .A(round_reg[75]), .B(round_reg[715]), .Z(n5593) );
  XOR U6793 ( .A(round_reg[1389]), .B(n1911), .Z(n1194) );
  XOR U6794 ( .A(n5326), .B(n4901), .Z(n1911) );
  XOR U6795 ( .A(n5594), .B(n5595), .Z(n4901) );
  XNOR U6796 ( .A(round_reg[1324]), .B(round_reg[1004]), .Z(n5595) );
  XOR U6797 ( .A(round_reg[364]), .B(n5596), .Z(n5594) );
  XOR U6798 ( .A(round_reg[684]), .B(round_reg[44]), .Z(n5596) );
  XOR U6799 ( .A(n5597), .B(n5598), .Z(n5326) );
  XNOR U6800 ( .A(round_reg[1453]), .B(round_reg[1133]), .Z(n5598) );
  XOR U6801 ( .A(round_reg[173]), .B(n5599), .Z(n5597) );
  XOR U6802 ( .A(round_reg[813]), .B(round_reg[493]), .Z(n5599) );
  XOR U6803 ( .A(n5600), .B(n4800), .Z(out[1032]) );
  XOR U6804 ( .A(round_reg[539]), .B(n2267), .Z(n4800) );
  XNOR U6805 ( .A(n5601), .B(n5602), .Z(n2267) );
  AND U6806 ( .A(n1198), .B(n1196), .Z(n5600) );
  XNOR U6807 ( .A(round_reg[139]), .B(n2314), .Z(n1196) );
  XOR U6808 ( .A(n5009), .B(n4703), .Z(n2314) );
  XOR U6809 ( .A(n5603), .B(n5604), .Z(n4703) );
  XNOR U6810 ( .A(round_reg[1354]), .B(round_reg[1034]), .Z(n5604) );
  XOR U6811 ( .A(round_reg[394]), .B(n5605), .Z(n5603) );
  XOR U6812 ( .A(round_reg[74]), .B(round_reg[714]), .Z(n5605) );
  XOR U6813 ( .A(n5606), .B(n5607), .Z(n5009) );
  XNOR U6814 ( .A(round_reg[1483]), .B(round_reg[1163]), .Z(n5607) );
  XOR U6815 ( .A(round_reg[203]), .B(n5608), .Z(n5606) );
  XOR U6816 ( .A(round_reg[843]), .B(round_reg[523]), .Z(n5608) );
  XNOR U6817 ( .A(round_reg[1388]), .B(n1914), .Z(n1198) );
  XOR U6818 ( .A(n5609), .B(n5610), .Z(n5339) );
  XNOR U6819 ( .A(round_reg[1452]), .B(round_reg[1132]), .Z(n5610) );
  XOR U6820 ( .A(round_reg[172]), .B(n5611), .Z(n5609) );
  XOR U6821 ( .A(round_reg[812]), .B(round_reg[492]), .Z(n5611) );
  XNOR U6822 ( .A(n5612), .B(n5613), .Z(n4906) );
  XNOR U6823 ( .A(round_reg[1323]), .B(round_reg[1003]), .Z(n5613) );
  XOR U6824 ( .A(round_reg[363]), .B(n5614), .Z(n5612) );
  XOR U6825 ( .A(round_reg[683]), .B(round_reg[43]), .Z(n5614) );
  XOR U6826 ( .A(n5615), .B(n4807), .Z(out[1031]) );
  XOR U6827 ( .A(round_reg[538]), .B(n2271), .Z(n4807) );
  XNOR U6828 ( .A(n5616), .B(n5617), .Z(n2271) );
  AND U6829 ( .A(n1202), .B(n1200), .Z(n5615) );
  XNOR U6830 ( .A(round_reg[138]), .B(n2318), .Z(n1200) );
  XOR U6831 ( .A(n4707), .B(n5012), .Z(n2318) );
  XOR U6832 ( .A(n5618), .B(n5619), .Z(n5012) );
  XNOR U6833 ( .A(round_reg[1482]), .B(round_reg[1162]), .Z(n5619) );
  XOR U6834 ( .A(round_reg[202]), .B(n5620), .Z(n5618) );
  XOR U6835 ( .A(round_reg[842]), .B(round_reg[522]), .Z(n5620) );
  XOR U6836 ( .A(n5621), .B(n5622), .Z(n4707) );
  XNOR U6837 ( .A(round_reg[1353]), .B(round_reg[1033]), .Z(n5622) );
  XOR U6838 ( .A(round_reg[393]), .B(n5623), .Z(n5621) );
  XOR U6839 ( .A(round_reg[73]), .B(round_reg[713]), .Z(n5623) );
  XNOR U6840 ( .A(round_reg[1387]), .B(n1917), .Z(n1202) );
  XOR U6841 ( .A(n5624), .B(n5625), .Z(n5361) );
  XNOR U6842 ( .A(round_reg[1451]), .B(round_reg[1131]), .Z(n5625) );
  XOR U6843 ( .A(round_reg[171]), .B(n5626), .Z(n5624) );
  XOR U6844 ( .A(round_reg[811]), .B(round_reg[491]), .Z(n5626) );
  XNOR U6845 ( .A(n5627), .B(n5628), .Z(n4910) );
  XNOR U6846 ( .A(round_reg[1322]), .B(round_reg[1002]), .Z(n5628) );
  XOR U6847 ( .A(round_reg[362]), .B(n5629), .Z(n5627) );
  XOR U6848 ( .A(round_reg[682]), .B(round_reg[42]), .Z(n5629) );
  XOR U6849 ( .A(n5630), .B(n4811), .Z(out[1030]) );
  XOR U6850 ( .A(round_reg[537]), .B(n2275), .Z(n4811) );
  XNOR U6851 ( .A(n5631), .B(n5632), .Z(n2275) );
  AND U6852 ( .A(n1206), .B(n1204), .Z(n5630) );
  XNOR U6853 ( .A(round_reg[137]), .B(n2322), .Z(n1204) );
  XNOR U6854 ( .A(n4712), .B(n5016), .Z(n2322) );
  XNOR U6855 ( .A(n5633), .B(n5634), .Z(n5016) );
  XNOR U6856 ( .A(round_reg[1481]), .B(round_reg[1161]), .Z(n5634) );
  XOR U6857 ( .A(round_reg[201]), .B(n5635), .Z(n5633) );
  XOR U6858 ( .A(round_reg[841]), .B(round_reg[521]), .Z(n5635) );
  XOR U6859 ( .A(n5636), .B(n5637), .Z(n4712) );
  XNOR U6860 ( .A(round_reg[1352]), .B(round_reg[1032]), .Z(n5637) );
  XOR U6861 ( .A(round_reg[392]), .B(n5638), .Z(n5636) );
  XOR U6862 ( .A(round_reg[72]), .B(round_reg[712]), .Z(n5638) );
  XNOR U6863 ( .A(round_reg[1386]), .B(n1920), .Z(n1206) );
  XOR U6864 ( .A(n5639), .B(n5640), .Z(n5372) );
  XNOR U6865 ( .A(round_reg[1450]), .B(round_reg[1130]), .Z(n5640) );
  XOR U6866 ( .A(round_reg[170]), .B(n5641), .Z(n5639) );
  XOR U6867 ( .A(round_reg[810]), .B(round_reg[490]), .Z(n5641) );
  XNOR U6868 ( .A(n5642), .B(n5643), .Z(n4914) );
  XNOR U6869 ( .A(round_reg[1321]), .B(round_reg[1001]), .Z(n5643) );
  XOR U6870 ( .A(round_reg[361]), .B(n5644), .Z(n5642) );
  XOR U6871 ( .A(round_reg[681]), .B(round_reg[41]), .Z(n5644) );
  XOR U6872 ( .A(n5645), .B(n3473), .Z(out[102]) );
  IV U6873 ( .A(n3575), .Z(n3473) );
  XNOR U6874 ( .A(round_reg[637]), .B(n2321), .Z(n3575) );
  XNOR U6875 ( .A(n5347), .B(n5646), .Z(n2321) );
  XOR U6876 ( .A(n5647), .B(n5648), .Z(n5347) );
  XNOR U6877 ( .A(round_reg[1341]), .B(round_reg[1021]), .Z(n5648) );
  XOR U6878 ( .A(round_reg[381]), .B(n5649), .Z(n5647) );
  XOR U6879 ( .A(round_reg[701]), .B(round_reg[61]), .Z(n5649) );
  AND U6880 ( .A(n3128), .B(n3130), .Z(n5645) );
  XOR U6881 ( .A(round_reg[1448]), .B(n2186), .Z(n3130) );
  XOR U6882 ( .A(n4913), .B(n5650), .Z(n2186) );
  XOR U6883 ( .A(n5651), .B(n5652), .Z(n4913) );
  XNOR U6884 ( .A(round_reg[1512]), .B(round_reg[1192]), .Z(n5652) );
  XOR U6885 ( .A(round_reg[232]), .B(n5653), .Z(n5651) );
  XOR U6886 ( .A(round_reg[872]), .B(round_reg[552]), .Z(n5653) );
  XNOR U6887 ( .A(round_reg[228]), .B(n2227), .Z(n3128) );
  XNOR U6888 ( .A(n5654), .B(n5655), .Z(n2227) );
  XOR U6889 ( .A(n5656), .B(n4815), .Z(out[1029]) );
  XOR U6890 ( .A(round_reg[536]), .B(n2279), .Z(n4815) );
  XNOR U6891 ( .A(n5657), .B(n5658), .Z(n2279) );
  ANDN U6892 ( .B(n1208), .A(n1209), .Z(n5656) );
  XOR U6893 ( .A(round_reg[1385]), .B(n1923), .Z(n1209) );
  XOR U6894 ( .A(n5659), .B(n5660), .Z(n5385) );
  XNOR U6895 ( .A(round_reg[1449]), .B(round_reg[1129]), .Z(n5660) );
  XOR U6896 ( .A(round_reg[169]), .B(n5661), .Z(n5659) );
  XOR U6897 ( .A(round_reg[809]), .B(round_reg[489]), .Z(n5661) );
  XNOR U6898 ( .A(n5662), .B(n5663), .Z(n4918) );
  XNOR U6899 ( .A(round_reg[1320]), .B(round_reg[1000]), .Z(n5663) );
  XOR U6900 ( .A(round_reg[360]), .B(n5664), .Z(n5662) );
  XOR U6901 ( .A(round_reg[680]), .B(round_reg[40]), .Z(n5664) );
  XNOR U6902 ( .A(round_reg[136]), .B(n2326), .Z(n1208) );
  XNOR U6903 ( .A(n4718), .B(n5019), .Z(n2326) );
  XNOR U6904 ( .A(n5665), .B(n5666), .Z(n5019) );
  XNOR U6905 ( .A(round_reg[1480]), .B(round_reg[1160]), .Z(n5666) );
  XOR U6906 ( .A(round_reg[200]), .B(n5667), .Z(n5665) );
  XOR U6907 ( .A(round_reg[840]), .B(round_reg[520]), .Z(n5667) );
  XOR U6908 ( .A(n5668), .B(n5669), .Z(n4718) );
  XNOR U6909 ( .A(round_reg[1351]), .B(round_reg[1031]), .Z(n5669) );
  XOR U6910 ( .A(round_reg[391]), .B(n5670), .Z(n5668) );
  XOR U6911 ( .A(round_reg[71]), .B(round_reg[711]), .Z(n5670) );
  XOR U6912 ( .A(n5671), .B(n4819), .Z(out[1028]) );
  XOR U6913 ( .A(round_reg[535]), .B(n2283), .Z(n4819) );
  XNOR U6914 ( .A(n5672), .B(n5673), .Z(n2283) );
  ANDN U6915 ( .B(n1212), .A(n1213), .Z(n5671) );
  XOR U6916 ( .A(round_reg[1384]), .B(n1930), .Z(n1213) );
  XOR U6917 ( .A(n5674), .B(n5675), .Z(n5398) );
  XNOR U6918 ( .A(round_reg[1448]), .B(round_reg[1128]), .Z(n5675) );
  XOR U6919 ( .A(round_reg[168]), .B(n5676), .Z(n5674) );
  XOR U6920 ( .A(round_reg[808]), .B(round_reg[488]), .Z(n5676) );
  XNOR U6921 ( .A(n5677), .B(n5678), .Z(n4922) );
  XNOR U6922 ( .A(round_reg[359]), .B(round_reg[1319]), .Z(n5678) );
  XOR U6923 ( .A(round_reg[39]), .B(n5679), .Z(n5677) );
  XOR U6924 ( .A(round_reg[999]), .B(round_reg[679]), .Z(n5679) );
  XNOR U6925 ( .A(round_reg[135]), .B(n2330), .Z(n1212) );
  XNOR U6926 ( .A(n4722), .B(n5025), .Z(n2330) );
  XNOR U6927 ( .A(n5680), .B(n5681), .Z(n5025) );
  XNOR U6928 ( .A(round_reg[1479]), .B(round_reg[1159]), .Z(n5681) );
  XOR U6929 ( .A(round_reg[199]), .B(n5682), .Z(n5680) );
  XOR U6930 ( .A(round_reg[839]), .B(round_reg[519]), .Z(n5682) );
  XOR U6931 ( .A(n5683), .B(n5684), .Z(n4722) );
  XNOR U6932 ( .A(round_reg[1350]), .B(round_reg[1030]), .Z(n5684) );
  XOR U6933 ( .A(round_reg[390]), .B(n5685), .Z(n5683) );
  XOR U6934 ( .A(round_reg[710]), .B(round_reg[70]), .Z(n5685) );
  XOR U6935 ( .A(n5686), .B(n4823), .Z(out[1027]) );
  XOR U6936 ( .A(round_reg[534]), .B(n2287), .Z(n4823) );
  XNOR U6937 ( .A(n5687), .B(n5688), .Z(n2287) );
  ANDN U6938 ( .B(n1216), .A(n1217), .Z(n5686) );
  XOR U6939 ( .A(round_reg[1383]), .B(n1933), .Z(n1217) );
  XOR U6940 ( .A(n5689), .B(n5690), .Z(n5411) );
  XNOR U6941 ( .A(round_reg[1447]), .B(round_reg[1127]), .Z(n5690) );
  XOR U6942 ( .A(round_reg[167]), .B(n5691), .Z(n5689) );
  XOR U6943 ( .A(round_reg[807]), .B(round_reg[487]), .Z(n5691) );
  XNOR U6944 ( .A(n5692), .B(n5693), .Z(n4928) );
  XNOR U6945 ( .A(round_reg[358]), .B(round_reg[1318]), .Z(n5693) );
  XOR U6946 ( .A(round_reg[38]), .B(n5694), .Z(n5692) );
  XOR U6947 ( .A(round_reg[998]), .B(round_reg[678]), .Z(n5694) );
  XNOR U6948 ( .A(round_reg[134]), .B(n2334), .Z(n1216) );
  XNOR U6949 ( .A(n4726), .B(n5028), .Z(n2334) );
  XNOR U6950 ( .A(n5695), .B(n5696), .Z(n5028) );
  XNOR U6951 ( .A(round_reg[1478]), .B(round_reg[1158]), .Z(n5696) );
  XOR U6952 ( .A(round_reg[198]), .B(n5697), .Z(n5695) );
  XOR U6953 ( .A(round_reg[838]), .B(round_reg[518]), .Z(n5697) );
  XOR U6954 ( .A(n5698), .B(n5699), .Z(n4726) );
  XNOR U6955 ( .A(round_reg[1349]), .B(round_reg[1029]), .Z(n5699) );
  XOR U6956 ( .A(round_reg[389]), .B(n5700), .Z(n5698) );
  XOR U6957 ( .A(round_reg[709]), .B(round_reg[69]), .Z(n5700) );
  XOR U6958 ( .A(n5701), .B(n4827), .Z(out[1026]) );
  XOR U6959 ( .A(round_reg[533]), .B(n2291), .Z(n4827) );
  XNOR U6960 ( .A(n5702), .B(n5703), .Z(n2291) );
  ANDN U6961 ( .B(n1220), .A(n1221), .Z(n5701) );
  XOR U6962 ( .A(round_reg[1382]), .B(n1712), .Z(n1221) );
  XOR U6963 ( .A(n5704), .B(n5705), .Z(n5424) );
  XNOR U6964 ( .A(round_reg[1446]), .B(round_reg[1126]), .Z(n5705) );
  XOR U6965 ( .A(round_reg[166]), .B(n5706), .Z(n5704) );
  XOR U6966 ( .A(round_reg[806]), .B(round_reg[486]), .Z(n5706) );
  XNOR U6967 ( .A(n5707), .B(n5708), .Z(n4932) );
  XNOR U6968 ( .A(round_reg[357]), .B(round_reg[1317]), .Z(n5708) );
  XOR U6969 ( .A(round_reg[37]), .B(n5709), .Z(n5707) );
  XOR U6970 ( .A(round_reg[997]), .B(round_reg[677]), .Z(n5709) );
  XNOR U6971 ( .A(round_reg[133]), .B(n2338), .Z(n1220) );
  XNOR U6972 ( .A(n4730), .B(n5031), .Z(n2338) );
  XNOR U6973 ( .A(n5710), .B(n5711), .Z(n5031) );
  XNOR U6974 ( .A(round_reg[1477]), .B(round_reg[1157]), .Z(n5711) );
  XOR U6975 ( .A(round_reg[197]), .B(n5712), .Z(n5710) );
  XOR U6976 ( .A(round_reg[837]), .B(round_reg[517]), .Z(n5712) );
  XOR U6977 ( .A(n5713), .B(n5714), .Z(n4730) );
  XNOR U6978 ( .A(round_reg[1348]), .B(round_reg[1028]), .Z(n5714) );
  XOR U6979 ( .A(round_reg[388]), .B(n5715), .Z(n5713) );
  XOR U6980 ( .A(round_reg[708]), .B(round_reg[68]), .Z(n5715) );
  XOR U6981 ( .A(n5716), .B(n4831), .Z(out[1025]) );
  XOR U6982 ( .A(round_reg[532]), .B(n2295), .Z(n4831) );
  XNOR U6983 ( .A(n5717), .B(n5718), .Z(n2295) );
  ANDN U6984 ( .B(n1224), .A(n1225), .Z(n5716) );
  XOR U6985 ( .A(round_reg[1381]), .B(n1715), .Z(n1225) );
  XOR U6986 ( .A(n5719), .B(n5720), .Z(n5437) );
  XNOR U6987 ( .A(round_reg[1445]), .B(round_reg[1125]), .Z(n5720) );
  XOR U6988 ( .A(round_reg[165]), .B(n5721), .Z(n5719) );
  XOR U6989 ( .A(round_reg[805]), .B(round_reg[485]), .Z(n5721) );
  XNOR U6990 ( .A(n5722), .B(n5723), .Z(n4936) );
  XNOR U6991 ( .A(round_reg[356]), .B(round_reg[1316]), .Z(n5723) );
  XOR U6992 ( .A(round_reg[36]), .B(n5724), .Z(n5722) );
  XOR U6993 ( .A(round_reg[996]), .B(round_reg[676]), .Z(n5724) );
  XNOR U6994 ( .A(round_reg[132]), .B(n2342), .Z(n1224) );
  XNOR U6995 ( .A(n4734), .B(n5034), .Z(n2342) );
  XNOR U6996 ( .A(n5725), .B(n5726), .Z(n5034) );
  XNOR U6997 ( .A(round_reg[1476]), .B(round_reg[1156]), .Z(n5726) );
  XOR U6998 ( .A(round_reg[196]), .B(n5727), .Z(n5725) );
  XOR U6999 ( .A(round_reg[836]), .B(round_reg[516]), .Z(n5727) );
  XOR U7000 ( .A(n5728), .B(n5729), .Z(n4734) );
  XNOR U7001 ( .A(round_reg[1347]), .B(round_reg[1027]), .Z(n5729) );
  XOR U7002 ( .A(round_reg[387]), .B(n5730), .Z(n5728) );
  XOR U7003 ( .A(round_reg[707]), .B(round_reg[67]), .Z(n5730) );
  XOR U7004 ( .A(n5731), .B(n4835), .Z(out[1024]) );
  XOR U7005 ( .A(round_reg[531]), .B(n2299), .Z(n4835) );
  XNOR U7006 ( .A(n5732), .B(n5733), .Z(n2299) );
  ANDN U7007 ( .B(n1228), .A(n1229), .Z(n5731) );
  XOR U7008 ( .A(round_reg[1380]), .B(n1722), .Z(n1229) );
  XOR U7009 ( .A(n5734), .B(n5735), .Z(n5495) );
  XNOR U7010 ( .A(round_reg[1444]), .B(round_reg[1124]), .Z(n5735) );
  XOR U7011 ( .A(round_reg[164]), .B(n5736), .Z(n5734) );
  XOR U7012 ( .A(round_reg[804]), .B(round_reg[484]), .Z(n5736) );
  XNOR U7013 ( .A(n5737), .B(n5738), .Z(n4939) );
  XNOR U7014 ( .A(round_reg[355]), .B(round_reg[1315]), .Z(n5738) );
  XOR U7015 ( .A(round_reg[35]), .B(n5739), .Z(n5737) );
  XOR U7016 ( .A(round_reg[995]), .B(round_reg[675]), .Z(n5739) );
  XNOR U7017 ( .A(round_reg[131]), .B(n2350), .Z(n1228) );
  XNOR U7018 ( .A(n4738), .B(n5037), .Z(n2350) );
  XNOR U7019 ( .A(n5740), .B(n5741), .Z(n5037) );
  XNOR U7020 ( .A(round_reg[1475]), .B(round_reg[1155]), .Z(n5741) );
  XOR U7021 ( .A(round_reg[195]), .B(n5742), .Z(n5740) );
  XOR U7022 ( .A(round_reg[835]), .B(round_reg[515]), .Z(n5742) );
  XOR U7023 ( .A(n5743), .B(n5744), .Z(n4738) );
  XNOR U7024 ( .A(round_reg[1346]), .B(round_reg[1026]), .Z(n5744) );
  XOR U7025 ( .A(round_reg[386]), .B(n5745), .Z(n5743) );
  XOR U7026 ( .A(round_reg[706]), .B(round_reg[66]), .Z(n5745) );
  XOR U7027 ( .A(n5746), .B(n4837), .Z(out[1023]) );
  XOR U7028 ( .A(round_reg[130]), .B(n2354), .Z(n4837) );
  ANDN U7029 ( .B(n4409), .A(n4407), .Z(n5746) );
  XNOR U7030 ( .A(round_reg[1379]), .B(n1725), .Z(n4407) );
  XOR U7031 ( .A(n5747), .B(n5748), .Z(n5654) );
  XNOR U7032 ( .A(round_reg[1443]), .B(round_reg[1123]), .Z(n5748) );
  XOR U7033 ( .A(round_reg[163]), .B(n5749), .Z(n5747) );
  XOR U7034 ( .A(round_reg[803]), .B(round_reg[483]), .Z(n5749) );
  XNOR U7035 ( .A(n5750), .B(n5751), .Z(n4942) );
  XNOR U7036 ( .A(round_reg[34]), .B(round_reg[1314]), .Z(n5751) );
  XOR U7037 ( .A(round_reg[354]), .B(n5752), .Z(n5750) );
  XOR U7038 ( .A(round_reg[994]), .B(round_reg[674]), .Z(n5752) );
  XNOR U7039 ( .A(round_reg[1003]), .B(n4305), .Z(n4409) );
  XOR U7040 ( .A(n5753), .B(n5386), .Z(n4305) );
  XNOR U7041 ( .A(n5754), .B(n5755), .Z(n5386) );
  XNOR U7042 ( .A(round_reg[1578]), .B(round_reg[1258]), .Z(n5755) );
  XOR U7043 ( .A(round_reg[298]), .B(n5756), .Z(n5754) );
  XOR U7044 ( .A(round_reg[938]), .B(round_reg[618]), .Z(n5756) );
  XOR U7045 ( .A(n5757), .B(n4839), .Z(out[1022]) );
  XOR U7046 ( .A(round_reg[129]), .B(n2358), .Z(n4839) );
  XNOR U7047 ( .A(n4746), .B(n5090), .Z(n2358) );
  XNOR U7048 ( .A(n5758), .B(n5759), .Z(n5090) );
  XNOR U7049 ( .A(round_reg[1473]), .B(round_reg[1153]), .Z(n5759) );
  XOR U7050 ( .A(round_reg[193]), .B(n5760), .Z(n5758) );
  XOR U7051 ( .A(round_reg[833]), .B(round_reg[513]), .Z(n5760) );
  XOR U7052 ( .A(n5761), .B(n5762), .Z(n4746) );
  XNOR U7053 ( .A(round_reg[1344]), .B(round_reg[1024]), .Z(n5762) );
  XOR U7054 ( .A(round_reg[384]), .B(n5763), .Z(n5761) );
  XOR U7055 ( .A(round_reg[704]), .B(round_reg[64]), .Z(n5763) );
  ANDN U7056 ( .B(n4413), .A(n4411), .Z(n5757) );
  XOR U7057 ( .A(round_reg[1378]), .B(n1728), .Z(n4411) );
  XNOR U7058 ( .A(n5764), .B(n4945), .Z(n1728) );
  XNOR U7059 ( .A(n5765), .B(n5766), .Z(n4945) );
  XNOR U7060 ( .A(round_reg[33]), .B(round_reg[1313]), .Z(n5766) );
  XOR U7061 ( .A(round_reg[353]), .B(n5767), .Z(n5765) );
  XOR U7062 ( .A(round_reg[993]), .B(round_reg[673]), .Z(n5767) );
  XNOR U7063 ( .A(round_reg[1002]), .B(n4308), .Z(n4413) );
  XOR U7064 ( .A(n5768), .B(n5399), .Z(n4308) );
  XNOR U7065 ( .A(n5769), .B(n5770), .Z(n5399) );
  XNOR U7066 ( .A(round_reg[1577]), .B(round_reg[1257]), .Z(n5770) );
  XOR U7067 ( .A(round_reg[297]), .B(n5771), .Z(n5769) );
  XOR U7068 ( .A(round_reg[937]), .B(round_reg[617]), .Z(n5771) );
  XOR U7069 ( .A(n5772), .B(n4845), .Z(out[1021]) );
  XOR U7070 ( .A(round_reg[128]), .B(n2362), .Z(n4845) );
  XNOR U7071 ( .A(n4750), .B(n5143), .Z(n2362) );
  XNOR U7072 ( .A(n5773), .B(n5774), .Z(n5143) );
  XNOR U7073 ( .A(round_reg[1472]), .B(round_reg[1152]), .Z(n5774) );
  XOR U7074 ( .A(round_reg[192]), .B(n5775), .Z(n5773) );
  XOR U7075 ( .A(round_reg[832]), .B(round_reg[512]), .Z(n5775) );
  XOR U7076 ( .A(n5776), .B(n5777), .Z(n4750) );
  XNOR U7077 ( .A(round_reg[127]), .B(round_reg[1087]), .Z(n5777) );
  XOR U7078 ( .A(round_reg[1407]), .B(n5778), .Z(n5776) );
  XOR U7079 ( .A(round_reg[767]), .B(round_reg[447]), .Z(n5778) );
  ANDN U7080 ( .B(n4417), .A(n4415), .Z(n5772) );
  XOR U7081 ( .A(round_reg[1377]), .B(n1731), .Z(n4415) );
  XNOR U7082 ( .A(n5779), .B(n4948), .Z(n1731) );
  XNOR U7083 ( .A(n5780), .B(n5781), .Z(n4948) );
  XNOR U7084 ( .A(round_reg[32]), .B(round_reg[1312]), .Z(n5781) );
  XOR U7085 ( .A(round_reg[352]), .B(n5782), .Z(n5780) );
  XOR U7086 ( .A(round_reg[992]), .B(round_reg[672]), .Z(n5782) );
  XOR U7087 ( .A(round_reg[1001]), .B(n1977), .Z(n4417) );
  XNOR U7088 ( .A(n5356), .B(n5412), .Z(n1977) );
  XNOR U7089 ( .A(n5783), .B(n5784), .Z(n5412) );
  XNOR U7090 ( .A(round_reg[1576]), .B(round_reg[1256]), .Z(n5784) );
  XOR U7091 ( .A(round_reg[296]), .B(n5785), .Z(n5783) );
  XOR U7092 ( .A(round_reg[936]), .B(round_reg[616]), .Z(n5785) );
  XOR U7093 ( .A(n5786), .B(n5787), .Z(n5356) );
  XNOR U7094 ( .A(round_reg[1065]), .B(round_reg[105]), .Z(n5787) );
  XOR U7095 ( .A(round_reg[1385]), .B(n5788), .Z(n5786) );
  XOR U7096 ( .A(round_reg[745]), .B(round_reg[425]), .Z(n5788) );
  XOR U7097 ( .A(n5789), .B(n4849), .Z(out[1020]) );
  XOR U7098 ( .A(round_reg[191]), .B(n2366), .Z(n4849) );
  XNOR U7099 ( .A(n4754), .B(n5210), .Z(n2366) );
  XNOR U7100 ( .A(n5790), .B(n5791), .Z(n5210) );
  XNOR U7101 ( .A(round_reg[1535]), .B(round_reg[1215]), .Z(n5791) );
  XOR U7102 ( .A(round_reg[255]), .B(n5792), .Z(n5790) );
  XOR U7103 ( .A(round_reg[895]), .B(round_reg[575]), .Z(n5792) );
  XOR U7104 ( .A(n5793), .B(n5794), .Z(n4754) );
  XNOR U7105 ( .A(round_reg[126]), .B(round_reg[1086]), .Z(n5794) );
  XOR U7106 ( .A(round_reg[1406]), .B(n5795), .Z(n5793) );
  XOR U7107 ( .A(round_reg[766]), .B(round_reg[446]), .Z(n5795) );
  ANDN U7108 ( .B(n4421), .A(n4419), .Z(n5789) );
  XOR U7109 ( .A(round_reg[1376]), .B(n1734), .Z(n4419) );
  XNOR U7110 ( .A(n5512), .B(n4951), .Z(n1734) );
  XNOR U7111 ( .A(n5796), .B(n5797), .Z(n4951) );
  XNOR U7112 ( .A(round_reg[31]), .B(round_reg[1311]), .Z(n5797) );
  XOR U7113 ( .A(round_reg[351]), .B(n5798), .Z(n5796) );
  XOR U7114 ( .A(round_reg[991]), .B(round_reg[671]), .Z(n5798) );
  XOR U7115 ( .A(n5799), .B(n5800), .Z(n5512) );
  XNOR U7116 ( .A(round_reg[1440]), .B(round_reg[1120]), .Z(n5800) );
  XOR U7117 ( .A(round_reg[160]), .B(n5801), .Z(n5799) );
  XOR U7118 ( .A(round_reg[800]), .B(round_reg[480]), .Z(n5801) );
  XOR U7119 ( .A(round_reg[1000]), .B(n1980), .Z(n4421) );
  XNOR U7120 ( .A(n5491), .B(n5425), .Z(n1980) );
  XNOR U7121 ( .A(n5802), .B(n5803), .Z(n5425) );
  XNOR U7122 ( .A(round_reg[1575]), .B(round_reg[1255]), .Z(n5803) );
  XOR U7123 ( .A(round_reg[295]), .B(n5804), .Z(n5802) );
  XOR U7124 ( .A(round_reg[935]), .B(round_reg[615]), .Z(n5804) );
  XOR U7125 ( .A(n5805), .B(n5806), .Z(n5491) );
  XNOR U7126 ( .A(round_reg[1064]), .B(round_reg[104]), .Z(n5806) );
  XOR U7127 ( .A(round_reg[1384]), .B(n5807), .Z(n5805) );
  XOR U7128 ( .A(round_reg[744]), .B(round_reg[424]), .Z(n5807) );
  XOR U7129 ( .A(n5808), .B(n3476), .Z(out[101]) );
  IV U7130 ( .A(n3577), .Z(n3476) );
  XNOR U7131 ( .A(round_reg[636]), .B(n2325), .Z(n3577) );
  XNOR U7132 ( .A(n5370), .B(n5809), .Z(n2325) );
  XOR U7133 ( .A(n5810), .B(n5811), .Z(n5370) );
  XNOR U7134 ( .A(round_reg[1340]), .B(round_reg[1020]), .Z(n5811) );
  XOR U7135 ( .A(round_reg[380]), .B(n5812), .Z(n5810) );
  XOR U7136 ( .A(round_reg[700]), .B(round_reg[60]), .Z(n5812) );
  AND U7137 ( .A(n3142), .B(n3144), .Z(n5808) );
  XOR U7138 ( .A(round_reg[1447]), .B(n2190), .Z(n3144) );
  XOR U7139 ( .A(n4917), .B(n5813), .Z(n2190) );
  XOR U7140 ( .A(n5814), .B(n5815), .Z(n4917) );
  XNOR U7141 ( .A(round_reg[1511]), .B(round_reg[1191]), .Z(n5815) );
  XOR U7142 ( .A(round_reg[231]), .B(n5816), .Z(n5814) );
  XOR U7143 ( .A(round_reg[871]), .B(round_reg[551]), .Z(n5816) );
  XNOR U7144 ( .A(round_reg[227]), .B(n2231), .Z(n3142) );
  XNOR U7145 ( .A(n5764), .B(n5817), .Z(n2231) );
  XOR U7146 ( .A(n5818), .B(n5819), .Z(n5764) );
  XNOR U7147 ( .A(round_reg[1442]), .B(round_reg[1122]), .Z(n5819) );
  XOR U7148 ( .A(round_reg[162]), .B(n5820), .Z(n5818) );
  XOR U7149 ( .A(round_reg[802]), .B(round_reg[482]), .Z(n5820) );
  XOR U7150 ( .A(n5821), .B(n4853), .Z(out[1019]) );
  XOR U7151 ( .A(round_reg[190]), .B(n2370), .Z(n4853) );
  XNOR U7152 ( .A(n4762), .B(n5352), .Z(n2370) );
  XNOR U7153 ( .A(n5822), .B(n5823), .Z(n5352) );
  XNOR U7154 ( .A(round_reg[1534]), .B(round_reg[1214]), .Z(n5823) );
  XOR U7155 ( .A(round_reg[254]), .B(n5824), .Z(n5822) );
  XOR U7156 ( .A(round_reg[894]), .B(round_reg[574]), .Z(n5824) );
  XOR U7157 ( .A(n5825), .B(n5826), .Z(n4762) );
  XNOR U7158 ( .A(round_reg[125]), .B(round_reg[1085]), .Z(n5826) );
  XOR U7159 ( .A(round_reg[1405]), .B(n5827), .Z(n5825) );
  XOR U7160 ( .A(round_reg[765]), .B(round_reg[445]), .Z(n5827) );
  ANDN U7161 ( .B(n4425), .A(n4423), .Z(n5821) );
  XOR U7162 ( .A(round_reg[1375]), .B(n1737), .Z(n4423) );
  XNOR U7163 ( .A(n5526), .B(n4954), .Z(n1737) );
  XNOR U7164 ( .A(n5828), .B(n5829), .Z(n4954) );
  XNOR U7165 ( .A(round_reg[30]), .B(round_reg[1310]), .Z(n5829) );
  XOR U7166 ( .A(round_reg[350]), .B(n5830), .Z(n5828) );
  XOR U7167 ( .A(round_reg[990]), .B(round_reg[670]), .Z(n5830) );
  XOR U7168 ( .A(n5831), .B(n5832), .Z(n5526) );
  XNOR U7169 ( .A(round_reg[1439]), .B(round_reg[1119]), .Z(n5832) );
  XOR U7170 ( .A(round_reg[159]), .B(n5833), .Z(n5831) );
  XOR U7171 ( .A(round_reg[799]), .B(round_reg[479]), .Z(n5833) );
  XOR U7172 ( .A(round_reg[999]), .B(n1983), .Z(n4425) );
  XNOR U7173 ( .A(n5650), .B(n5438), .Z(n1983) );
  XNOR U7174 ( .A(n5834), .B(n5835), .Z(n5438) );
  XNOR U7175 ( .A(round_reg[1574]), .B(round_reg[1254]), .Z(n5835) );
  XOR U7176 ( .A(round_reg[294]), .B(n5836), .Z(n5834) );
  XOR U7177 ( .A(round_reg[934]), .B(round_reg[614]), .Z(n5836) );
  XOR U7178 ( .A(n5837), .B(n5838), .Z(n5650) );
  XNOR U7179 ( .A(round_reg[1063]), .B(round_reg[103]), .Z(n5838) );
  XOR U7180 ( .A(round_reg[1383]), .B(n5839), .Z(n5837) );
  XOR U7181 ( .A(round_reg[743]), .B(round_reg[423]), .Z(n5839) );
  XOR U7182 ( .A(n5840), .B(n4857), .Z(out[1018]) );
  XOR U7183 ( .A(round_reg[189]), .B(n2374), .Z(n4857) );
  XNOR U7184 ( .A(n4766), .B(n5487), .Z(n2374) );
  XNOR U7185 ( .A(n5841), .B(n5842), .Z(n5487) );
  XNOR U7186 ( .A(round_reg[1533]), .B(round_reg[1213]), .Z(n5842) );
  XOR U7187 ( .A(round_reg[253]), .B(n5843), .Z(n5841) );
  XOR U7188 ( .A(round_reg[893]), .B(round_reg[573]), .Z(n5843) );
  XOR U7189 ( .A(n5844), .B(n5845), .Z(n4766) );
  XNOR U7190 ( .A(round_reg[124]), .B(round_reg[1084]), .Z(n5845) );
  XOR U7191 ( .A(round_reg[1404]), .B(n5846), .Z(n5844) );
  XOR U7192 ( .A(round_reg[764]), .B(round_reg[444]), .Z(n5846) );
  ANDN U7193 ( .B(n4429), .A(n4427), .Z(n5840) );
  XOR U7194 ( .A(round_reg[1374]), .B(n1740), .Z(n4427) );
  XNOR U7195 ( .A(n5541), .B(n4957), .Z(n1740) );
  XNOR U7196 ( .A(n5847), .B(n5848), .Z(n4957) );
  XNOR U7197 ( .A(round_reg[29]), .B(round_reg[1309]), .Z(n5848) );
  XOR U7198 ( .A(round_reg[349]), .B(n5849), .Z(n5847) );
  XOR U7199 ( .A(round_reg[989]), .B(round_reg[669]), .Z(n5849) );
  XOR U7200 ( .A(n5850), .B(n5851), .Z(n5541) );
  XNOR U7201 ( .A(round_reg[1438]), .B(round_reg[1118]), .Z(n5851) );
  XOR U7202 ( .A(round_reg[158]), .B(n5852), .Z(n5850) );
  XOR U7203 ( .A(round_reg[798]), .B(round_reg[478]), .Z(n5852) );
  XOR U7204 ( .A(round_reg[998]), .B(n1986), .Z(n4429) );
  XNOR U7205 ( .A(n5813), .B(n5496), .Z(n1986) );
  XNOR U7206 ( .A(n5853), .B(n5854), .Z(n5496) );
  XNOR U7207 ( .A(round_reg[1573]), .B(round_reg[1253]), .Z(n5854) );
  XOR U7208 ( .A(round_reg[293]), .B(n5855), .Z(n5853) );
  XOR U7209 ( .A(round_reg[933]), .B(round_reg[613]), .Z(n5855) );
  XOR U7210 ( .A(n5856), .B(n5857), .Z(n5813) );
  XNOR U7211 ( .A(round_reg[1062]), .B(round_reg[102]), .Z(n5857) );
  XOR U7212 ( .A(round_reg[1382]), .B(n5858), .Z(n5856) );
  XOR U7213 ( .A(round_reg[742]), .B(round_reg[422]), .Z(n5858) );
  XOR U7214 ( .A(n5859), .B(n4861), .Z(out[1017]) );
  XOR U7215 ( .A(round_reg[188]), .B(n2378), .Z(n4861) );
  XNOR U7216 ( .A(n4770), .B(n5646), .Z(n2378) );
  XNOR U7217 ( .A(n5860), .B(n5861), .Z(n5646) );
  XNOR U7218 ( .A(round_reg[1532]), .B(round_reg[1212]), .Z(n5861) );
  XOR U7219 ( .A(round_reg[252]), .B(n5862), .Z(n5860) );
  XOR U7220 ( .A(round_reg[892]), .B(round_reg[572]), .Z(n5862) );
  XOR U7221 ( .A(n5863), .B(n5864), .Z(n4770) );
  XNOR U7222 ( .A(round_reg[123]), .B(round_reg[1083]), .Z(n5864) );
  XOR U7223 ( .A(round_reg[1403]), .B(n5865), .Z(n5863) );
  XOR U7224 ( .A(round_reg[763]), .B(round_reg[443]), .Z(n5865) );
  ANDN U7225 ( .B(n4433), .A(n4431), .Z(n5859) );
  XOR U7226 ( .A(round_reg[1373]), .B(n1743), .Z(n4431) );
  XNOR U7227 ( .A(n5556), .B(n4961), .Z(n1743) );
  XNOR U7228 ( .A(n5866), .B(n5867), .Z(n4961) );
  XNOR U7229 ( .A(round_reg[28]), .B(round_reg[1308]), .Z(n5867) );
  XOR U7230 ( .A(round_reg[348]), .B(n5868), .Z(n5866) );
  XOR U7231 ( .A(round_reg[988]), .B(round_reg[668]), .Z(n5868) );
  XOR U7232 ( .A(n5869), .B(n5870), .Z(n5556) );
  XNOR U7233 ( .A(round_reg[1437]), .B(round_reg[1117]), .Z(n5870) );
  XOR U7234 ( .A(round_reg[157]), .B(n5871), .Z(n5869) );
  XOR U7235 ( .A(round_reg[797]), .B(round_reg[477]), .Z(n5871) );
  XOR U7236 ( .A(round_reg[997]), .B(n1993), .Z(n4433) );
  XNOR U7237 ( .A(n5872), .B(n5655), .Z(n1993) );
  XNOR U7238 ( .A(n5873), .B(n5874), .Z(n5655) );
  XNOR U7239 ( .A(round_reg[1572]), .B(round_reg[1252]), .Z(n5874) );
  XOR U7240 ( .A(round_reg[292]), .B(n5875), .Z(n5873) );
  XOR U7241 ( .A(round_reg[932]), .B(round_reg[612]), .Z(n5875) );
  XOR U7242 ( .A(n5876), .B(n4865), .Z(out[1016]) );
  XOR U7243 ( .A(round_reg[187]), .B(n2382), .Z(n4865) );
  XNOR U7244 ( .A(n4774), .B(n5809), .Z(n2382) );
  XNOR U7245 ( .A(n5877), .B(n5878), .Z(n5809) );
  XNOR U7246 ( .A(round_reg[1531]), .B(round_reg[1211]), .Z(n5878) );
  XOR U7247 ( .A(round_reg[251]), .B(n5879), .Z(n5877) );
  XOR U7248 ( .A(round_reg[891]), .B(round_reg[571]), .Z(n5879) );
  XOR U7249 ( .A(n5880), .B(n5881), .Z(n4774) );
  XNOR U7250 ( .A(round_reg[122]), .B(round_reg[1082]), .Z(n5881) );
  XOR U7251 ( .A(round_reg[1402]), .B(n5882), .Z(n5880) );
  XOR U7252 ( .A(round_reg[762]), .B(round_reg[442]), .Z(n5882) );
  ANDN U7253 ( .B(n4437), .A(n4435), .Z(n5876) );
  XOR U7254 ( .A(round_reg[1372]), .B(n1746), .Z(n4435) );
  XNOR U7255 ( .A(n5571), .B(n4964), .Z(n1746) );
  XNOR U7256 ( .A(n5883), .B(n5884), .Z(n4964) );
  XNOR U7257 ( .A(round_reg[27]), .B(round_reg[1307]), .Z(n5884) );
  XOR U7258 ( .A(round_reg[347]), .B(n5885), .Z(n5883) );
  XOR U7259 ( .A(round_reg[987]), .B(round_reg[667]), .Z(n5885) );
  XOR U7260 ( .A(n5886), .B(n5887), .Z(n5571) );
  XNOR U7261 ( .A(round_reg[1436]), .B(round_reg[1116]), .Z(n5887) );
  XOR U7262 ( .A(round_reg[156]), .B(n5888), .Z(n5886) );
  XOR U7263 ( .A(round_reg[796]), .B(round_reg[476]), .Z(n5888) );
  XOR U7264 ( .A(round_reg[996]), .B(n1996), .Z(n4437) );
  XNOR U7265 ( .A(n5227), .B(n5817), .Z(n1996) );
  XNOR U7266 ( .A(n5889), .B(n5890), .Z(n5817) );
  XNOR U7267 ( .A(round_reg[1571]), .B(round_reg[1251]), .Z(n5890) );
  XOR U7268 ( .A(round_reg[291]), .B(n5891), .Z(n5889) );
  XOR U7269 ( .A(round_reg[931]), .B(round_reg[611]), .Z(n5891) );
  XOR U7270 ( .A(n5892), .B(n5893), .Z(n5227) );
  XNOR U7271 ( .A(round_reg[1060]), .B(round_reg[100]), .Z(n5893) );
  XOR U7272 ( .A(round_reg[1380]), .B(n5894), .Z(n5892) );
  XOR U7273 ( .A(round_reg[740]), .B(round_reg[420]), .Z(n5894) );
  XOR U7274 ( .A(n5895), .B(n4869), .Z(out[1015]) );
  XOR U7275 ( .A(round_reg[186]), .B(n2386), .Z(n4869) );
  XNOR U7276 ( .A(n4778), .B(n5896), .Z(n2386) );
  XOR U7277 ( .A(n5897), .B(n5898), .Z(n4778) );
  XNOR U7278 ( .A(round_reg[121]), .B(round_reg[1081]), .Z(n5898) );
  XOR U7279 ( .A(round_reg[1401]), .B(n5899), .Z(n5897) );
  XOR U7280 ( .A(round_reg[761]), .B(round_reg[441]), .Z(n5899) );
  ANDN U7281 ( .B(n4441), .A(n4439), .Z(n5895) );
  XOR U7282 ( .A(round_reg[1371]), .B(n1749), .Z(n4439) );
  XNOR U7283 ( .A(n5586), .B(n4967), .Z(n1749) );
  XNOR U7284 ( .A(n5900), .B(n5901), .Z(n4967) );
  XNOR U7285 ( .A(round_reg[26]), .B(round_reg[1306]), .Z(n5901) );
  XOR U7286 ( .A(round_reg[346]), .B(n5902), .Z(n5900) );
  XOR U7287 ( .A(round_reg[986]), .B(round_reg[666]), .Z(n5902) );
  XOR U7288 ( .A(n5903), .B(n5904), .Z(n5586) );
  XNOR U7289 ( .A(round_reg[1435]), .B(round_reg[1115]), .Z(n5904) );
  XOR U7290 ( .A(round_reg[155]), .B(n5905), .Z(n5903) );
  XOR U7291 ( .A(round_reg[795]), .B(round_reg[475]), .Z(n5905) );
  XOR U7292 ( .A(round_reg[995]), .B(n1999), .Z(n4441) );
  XNOR U7293 ( .A(n5242), .B(n5906), .Z(n1999) );
  XOR U7294 ( .A(n5907), .B(n5908), .Z(n5242) );
  XNOR U7295 ( .A(round_reg[1379]), .B(round_reg[1059]), .Z(n5908) );
  XOR U7296 ( .A(round_reg[419]), .B(n5909), .Z(n5907) );
  XOR U7297 ( .A(round_reg[99]), .B(round_reg[739]), .Z(n5909) );
  XOR U7298 ( .A(n5910), .B(n4873), .Z(out[1014]) );
  XNOR U7299 ( .A(round_reg[185]), .B(n4125), .Z(n4873) );
  XOR U7300 ( .A(n4843), .B(n4783), .Z(n4125) );
  XNOR U7301 ( .A(n5911), .B(n5912), .Z(n4783) );
  XNOR U7302 ( .A(round_reg[120]), .B(round_reg[1080]), .Z(n5912) );
  XOR U7303 ( .A(round_reg[1400]), .B(n5913), .Z(n5911) );
  XOR U7304 ( .A(round_reg[760]), .B(round_reg[440]), .Z(n5913) );
  XOR U7305 ( .A(n5914), .B(n5915), .Z(n4843) );
  XNOR U7306 ( .A(round_reg[1529]), .B(round_reg[1209]), .Z(n5915) );
  XOR U7307 ( .A(round_reg[249]), .B(n5916), .Z(n5914) );
  XOR U7308 ( .A(round_reg[889]), .B(round_reg[569]), .Z(n5916) );
  ANDN U7309 ( .B(n4445), .A(n4443), .Z(n5910) );
  XNOR U7310 ( .A(round_reg[1370]), .B(n1756), .Z(n4443) );
  XOR U7311 ( .A(n5917), .B(n5918), .Z(n5601) );
  XNOR U7312 ( .A(round_reg[1434]), .B(round_reg[1114]), .Z(n5918) );
  XOR U7313 ( .A(round_reg[154]), .B(n5919), .Z(n5917) );
  XOR U7314 ( .A(round_reg[794]), .B(round_reg[474]), .Z(n5919) );
  XNOR U7315 ( .A(n5920), .B(n5921), .Z(n4970) );
  XNOR U7316 ( .A(round_reg[25]), .B(round_reg[1305]), .Z(n5921) );
  XOR U7317 ( .A(round_reg[345]), .B(n5922), .Z(n5920) );
  XOR U7318 ( .A(round_reg[985]), .B(round_reg[665]), .Z(n5922) );
  XNOR U7319 ( .A(round_reg[994]), .B(n4249), .Z(n4445) );
  XOR U7320 ( .A(n5511), .B(n5260), .Z(n4249) );
  XNOR U7321 ( .A(n5923), .B(n5924), .Z(n5260) );
  XNOR U7322 ( .A(round_reg[1378]), .B(round_reg[1058]), .Z(n5924) );
  XOR U7323 ( .A(round_reg[418]), .B(n5925), .Z(n5923) );
  XOR U7324 ( .A(round_reg[98]), .B(round_reg[738]), .Z(n5925) );
  XOR U7325 ( .A(n5926), .B(n5927), .Z(n5511) );
  XNOR U7326 ( .A(round_reg[1569]), .B(round_reg[1249]), .Z(n5927) );
  XOR U7327 ( .A(round_reg[289]), .B(n5928), .Z(n5926) );
  XOR U7328 ( .A(round_reg[929]), .B(round_reg[609]), .Z(n5928) );
  XOR U7329 ( .A(n5929), .B(n4877), .Z(out[1013]) );
  XNOR U7330 ( .A(round_reg[184]), .B(n4129), .Z(n4877) );
  XOR U7331 ( .A(n4847), .B(n4787), .Z(n4129) );
  XNOR U7332 ( .A(n5930), .B(n5931), .Z(n4787) );
  XNOR U7333 ( .A(round_reg[119]), .B(round_reg[1079]), .Z(n5931) );
  XOR U7334 ( .A(round_reg[1399]), .B(n5932), .Z(n5930) );
  XOR U7335 ( .A(round_reg[759]), .B(round_reg[439]), .Z(n5932) );
  XOR U7336 ( .A(n5933), .B(n5934), .Z(n4847) );
  XNOR U7337 ( .A(round_reg[1528]), .B(round_reg[1208]), .Z(n5934) );
  XOR U7338 ( .A(round_reg[248]), .B(n5935), .Z(n5933) );
  XOR U7339 ( .A(round_reg[888]), .B(round_reg[568]), .Z(n5935) );
  ANDN U7340 ( .B(n4451), .A(n4449), .Z(n5929) );
  XNOR U7341 ( .A(round_reg[1369]), .B(n1759), .Z(n4449) );
  XOR U7342 ( .A(n5936), .B(n5937), .Z(n5616) );
  XNOR U7343 ( .A(round_reg[1433]), .B(round_reg[1113]), .Z(n5937) );
  XOR U7344 ( .A(round_reg[153]), .B(n5938), .Z(n5936) );
  XOR U7345 ( .A(round_reg[793]), .B(round_reg[473]), .Z(n5938) );
  XNOR U7346 ( .A(n5939), .B(n5940), .Z(n4973) );
  XNOR U7347 ( .A(round_reg[24]), .B(round_reg[1304]), .Z(n5940) );
  XOR U7348 ( .A(round_reg[344]), .B(n5941), .Z(n5939) );
  XOR U7349 ( .A(round_reg[984]), .B(round_reg[664]), .Z(n5941) );
  XNOR U7350 ( .A(round_reg[993]), .B(n4324), .Z(n4451) );
  XOR U7351 ( .A(n5272), .B(n5527), .Z(n4324) );
  XNOR U7352 ( .A(n5942), .B(n5943), .Z(n5527) );
  XNOR U7353 ( .A(round_reg[1568]), .B(round_reg[1248]), .Z(n5943) );
  XOR U7354 ( .A(round_reg[288]), .B(n5944), .Z(n5942) );
  XOR U7355 ( .A(round_reg[928]), .B(round_reg[608]), .Z(n5944) );
  XOR U7356 ( .A(n5945), .B(n5946), .Z(n5272) );
  XNOR U7357 ( .A(round_reg[1377]), .B(round_reg[1057]), .Z(n5946) );
  XOR U7358 ( .A(round_reg[417]), .B(n5947), .Z(n5945) );
  XOR U7359 ( .A(round_reg[97]), .B(round_reg[737]), .Z(n5947) );
  XOR U7360 ( .A(n5948), .B(n4881), .Z(out[1012]) );
  XNOR U7361 ( .A(round_reg[183]), .B(n4715), .Z(n4881) );
  XOR U7362 ( .A(n4852), .B(n4791), .Z(n4715) );
  XNOR U7363 ( .A(n5949), .B(n5950), .Z(n4791) );
  XNOR U7364 ( .A(round_reg[118]), .B(round_reg[1078]), .Z(n5950) );
  XOR U7365 ( .A(round_reg[1398]), .B(n5951), .Z(n5949) );
  XOR U7366 ( .A(round_reg[758]), .B(round_reg[438]), .Z(n5951) );
  XOR U7367 ( .A(n5952), .B(n5953), .Z(n4852) );
  XNOR U7368 ( .A(round_reg[1527]), .B(round_reg[1207]), .Z(n5953) );
  XOR U7369 ( .A(round_reg[247]), .B(n5954), .Z(n5952) );
  XOR U7370 ( .A(round_reg[887]), .B(round_reg[567]), .Z(n5954) );
  ANDN U7371 ( .B(n4455), .A(n4453), .Z(n5948) );
  XNOR U7372 ( .A(round_reg[1368]), .B(n1762), .Z(n4453) );
  XOR U7373 ( .A(n5955), .B(n5956), .Z(n5631) );
  XNOR U7374 ( .A(round_reg[1432]), .B(round_reg[1112]), .Z(n5956) );
  XOR U7375 ( .A(round_reg[152]), .B(n5957), .Z(n5955) );
  XOR U7376 ( .A(round_reg[792]), .B(round_reg[472]), .Z(n5957) );
  XNOR U7377 ( .A(n5958), .B(n5959), .Z(n4976) );
  XNOR U7378 ( .A(round_reg[23]), .B(round_reg[1303]), .Z(n5959) );
  XOR U7379 ( .A(round_reg[343]), .B(n5960), .Z(n5958) );
  XOR U7380 ( .A(round_reg[983]), .B(round_reg[663]), .Z(n5960) );
  XNOR U7381 ( .A(round_reg[992]), .B(n4327), .Z(n4455) );
  XOR U7382 ( .A(n5287), .B(n5542), .Z(n4327) );
  XNOR U7383 ( .A(n5961), .B(n5962), .Z(n5542) );
  XNOR U7384 ( .A(round_reg[1567]), .B(round_reg[1247]), .Z(n5962) );
  XOR U7385 ( .A(round_reg[287]), .B(n5963), .Z(n5961) );
  XOR U7386 ( .A(round_reg[927]), .B(round_reg[607]), .Z(n5963) );
  XOR U7387 ( .A(n5964), .B(n5965), .Z(n5287) );
  XNOR U7388 ( .A(round_reg[1376]), .B(round_reg[1056]), .Z(n5965) );
  XOR U7389 ( .A(round_reg[416]), .B(n5966), .Z(n5964) );
  XOR U7390 ( .A(round_reg[96]), .B(round_reg[736]), .Z(n5966) );
  XOR U7391 ( .A(n5967), .B(n4887), .Z(out[1011]) );
  XNOR U7392 ( .A(round_reg[182]), .B(n4759), .Z(n4887) );
  XOR U7393 ( .A(n4856), .B(n4795), .Z(n4759) );
  XNOR U7394 ( .A(n5968), .B(n5969), .Z(n4795) );
  XNOR U7395 ( .A(round_reg[117]), .B(round_reg[1077]), .Z(n5969) );
  XOR U7396 ( .A(round_reg[1397]), .B(n5970), .Z(n5968) );
  XOR U7397 ( .A(round_reg[757]), .B(round_reg[437]), .Z(n5970) );
  XOR U7398 ( .A(n5971), .B(n5972), .Z(n4856) );
  XNOR U7399 ( .A(round_reg[1526]), .B(round_reg[1206]), .Z(n5972) );
  XOR U7400 ( .A(round_reg[246]), .B(n5973), .Z(n5971) );
  XOR U7401 ( .A(round_reg[886]), .B(round_reg[566]), .Z(n5973) );
  ANDN U7402 ( .B(n4459), .A(n4457), .Z(n5967) );
  XNOR U7403 ( .A(round_reg[1367]), .B(n1765), .Z(n4457) );
  XOR U7404 ( .A(n5974), .B(n5975), .Z(n5657) );
  XNOR U7405 ( .A(round_reg[1431]), .B(round_reg[1111]), .Z(n5975) );
  XOR U7406 ( .A(round_reg[151]), .B(n5976), .Z(n5974) );
  XOR U7407 ( .A(round_reg[791]), .B(round_reg[471]), .Z(n5976) );
  XNOR U7408 ( .A(n5977), .B(n5978), .Z(n4979) );
  XNOR U7409 ( .A(round_reg[22]), .B(round_reg[1302]), .Z(n5978) );
  XOR U7410 ( .A(round_reg[342]), .B(n5979), .Z(n5977) );
  XOR U7411 ( .A(round_reg[982]), .B(round_reg[662]), .Z(n5979) );
  XNOR U7412 ( .A(round_reg[991]), .B(n4330), .Z(n4459) );
  XOR U7413 ( .A(n5302), .B(n5557), .Z(n4330) );
  XNOR U7414 ( .A(n5980), .B(n5981), .Z(n5557) );
  XNOR U7415 ( .A(round_reg[1566]), .B(round_reg[1246]), .Z(n5981) );
  XOR U7416 ( .A(round_reg[286]), .B(n5982), .Z(n5980) );
  XOR U7417 ( .A(round_reg[926]), .B(round_reg[606]), .Z(n5982) );
  XOR U7418 ( .A(n5983), .B(n5984), .Z(n5302) );
  XNOR U7419 ( .A(round_reg[1375]), .B(round_reg[1055]), .Z(n5984) );
  XOR U7420 ( .A(round_reg[415]), .B(n5985), .Z(n5983) );
  XOR U7421 ( .A(round_reg[95]), .B(round_reg[735]), .Z(n5985) );
  XOR U7422 ( .A(n5986), .B(n4891), .Z(out[1010]) );
  XNOR U7423 ( .A(round_reg[181]), .B(n4802), .Z(n4891) );
  XOR U7424 ( .A(n4798), .B(n4860), .Z(n4802) );
  XNOR U7425 ( .A(n5987), .B(n5988), .Z(n4860) );
  XNOR U7426 ( .A(round_reg[1525]), .B(round_reg[1205]), .Z(n5988) );
  XOR U7427 ( .A(round_reg[245]), .B(n5989), .Z(n5987) );
  XOR U7428 ( .A(round_reg[885]), .B(round_reg[565]), .Z(n5989) );
  XOR U7429 ( .A(n5990), .B(n5991), .Z(n4798) );
  XNOR U7430 ( .A(round_reg[116]), .B(round_reg[1076]), .Z(n5991) );
  XOR U7431 ( .A(round_reg[1396]), .B(n5992), .Z(n5990) );
  XOR U7432 ( .A(round_reg[756]), .B(round_reg[436]), .Z(n5992) );
  ANDN U7433 ( .B(n4463), .A(n4461), .Z(n5986) );
  XNOR U7434 ( .A(round_reg[1366]), .B(n1768), .Z(n4461) );
  XOR U7435 ( .A(n5993), .B(n5994), .Z(n5672) );
  XNOR U7436 ( .A(round_reg[1430]), .B(round_reg[1110]), .Z(n5994) );
  XOR U7437 ( .A(round_reg[150]), .B(n5995), .Z(n5993) );
  XOR U7438 ( .A(round_reg[790]), .B(round_reg[470]), .Z(n5995) );
  XNOR U7439 ( .A(n5996), .B(n5997), .Z(n4982) );
  XNOR U7440 ( .A(round_reg[21]), .B(round_reg[1301]), .Z(n5997) );
  XOR U7441 ( .A(round_reg[341]), .B(n5998), .Z(n5996) );
  XOR U7442 ( .A(round_reg[981]), .B(round_reg[661]), .Z(n5998) );
  XNOR U7443 ( .A(round_reg[990]), .B(n4332), .Z(n4463) );
  XOR U7444 ( .A(n5317), .B(n5572), .Z(n4332) );
  XNOR U7445 ( .A(n5999), .B(n6000), .Z(n5572) );
  XNOR U7446 ( .A(round_reg[1565]), .B(round_reg[1245]), .Z(n6000) );
  XOR U7447 ( .A(round_reg[285]), .B(n6001), .Z(n5999) );
  XOR U7448 ( .A(round_reg[925]), .B(round_reg[605]), .Z(n6001) );
  XOR U7449 ( .A(n6002), .B(n6003), .Z(n5317) );
  XNOR U7450 ( .A(round_reg[1374]), .B(round_reg[1054]), .Z(n6003) );
  XOR U7451 ( .A(round_reg[414]), .B(n6004), .Z(n6002) );
  XOR U7452 ( .A(round_reg[94]), .B(round_reg[734]), .Z(n6004) );
  XOR U7453 ( .A(n6005), .B(n3478), .Z(out[100]) );
  IV U7454 ( .A(n3579), .Z(n3478) );
  XNOR U7455 ( .A(round_reg[635]), .B(n2329), .Z(n3579) );
  XNOR U7456 ( .A(n5380), .B(n5896), .Z(n2329) );
  XNOR U7457 ( .A(n6006), .B(n6007), .Z(n5896) );
  XNOR U7458 ( .A(round_reg[1530]), .B(round_reg[1210]), .Z(n6007) );
  XOR U7459 ( .A(round_reg[250]), .B(n6008), .Z(n6006) );
  XOR U7460 ( .A(round_reg[890]), .B(round_reg[570]), .Z(n6008) );
  XOR U7461 ( .A(n6009), .B(n6010), .Z(n5380) );
  XNOR U7462 ( .A(round_reg[1339]), .B(round_reg[1019]), .Z(n6010) );
  XOR U7463 ( .A(round_reg[379]), .B(n6011), .Z(n6009) );
  XOR U7464 ( .A(round_reg[699]), .B(round_reg[59]), .Z(n6011) );
  AND U7465 ( .A(n3156), .B(n3158), .Z(n6005) );
  XOR U7466 ( .A(round_reg[1446]), .B(n2194), .Z(n3158) );
  XOR U7467 ( .A(n4921), .B(n5872), .Z(n2194) );
  XOR U7468 ( .A(n6012), .B(n6013), .Z(n5872) );
  XNOR U7469 ( .A(round_reg[1061]), .B(round_reg[101]), .Z(n6013) );
  XOR U7470 ( .A(round_reg[1381]), .B(n6014), .Z(n6012) );
  XOR U7471 ( .A(round_reg[741]), .B(round_reg[421]), .Z(n6014) );
  XOR U7472 ( .A(n6015), .B(n6016), .Z(n4921) );
  XNOR U7473 ( .A(round_reg[1510]), .B(round_reg[1190]), .Z(n6016) );
  XOR U7474 ( .A(round_reg[230]), .B(n6017), .Z(n6015) );
  XOR U7475 ( .A(round_reg[870]), .B(round_reg[550]), .Z(n6017) );
  XNOR U7476 ( .A(round_reg[226]), .B(n2235), .Z(n3156) );
  XNOR U7477 ( .A(n5779), .B(n5906), .Z(n2235) );
  XNOR U7478 ( .A(n6018), .B(n6019), .Z(n5906) );
  XNOR U7479 ( .A(round_reg[1570]), .B(round_reg[1250]), .Z(n6019) );
  XOR U7480 ( .A(round_reg[290]), .B(n6020), .Z(n6018) );
  XOR U7481 ( .A(round_reg[930]), .B(round_reg[610]), .Z(n6020) );
  XOR U7482 ( .A(n6021), .B(n6022), .Z(n5779) );
  XNOR U7483 ( .A(round_reg[1441]), .B(round_reg[1121]), .Z(n6022) );
  XOR U7484 ( .A(round_reg[161]), .B(n6023), .Z(n6021) );
  XOR U7485 ( .A(round_reg[801]), .B(round_reg[481]), .Z(n6023) );
  XOR U7486 ( .A(n6024), .B(n4895), .Z(out[1009]) );
  XOR U7487 ( .A(round_reg[180]), .B(n2134), .Z(n4895) );
  XNOR U7488 ( .A(n4805), .B(n4864), .Z(n2134) );
  XNOR U7489 ( .A(n6025), .B(n6026), .Z(n4864) );
  XNOR U7490 ( .A(round_reg[1524]), .B(round_reg[1204]), .Z(n6026) );
  XOR U7491 ( .A(round_reg[244]), .B(n6027), .Z(n6025) );
  XOR U7492 ( .A(round_reg[884]), .B(round_reg[564]), .Z(n6027) );
  XOR U7493 ( .A(n6028), .B(n6029), .Z(n4805) );
  XNOR U7494 ( .A(round_reg[115]), .B(round_reg[1075]), .Z(n6029) );
  XOR U7495 ( .A(round_reg[1395]), .B(n6030), .Z(n6028) );
  XOR U7496 ( .A(round_reg[755]), .B(round_reg[435]), .Z(n6030) );
  ANDN U7497 ( .B(n4467), .A(n4465), .Z(n6024) );
  XNOR U7498 ( .A(round_reg[1365]), .B(n1771), .Z(n4465) );
  XOR U7499 ( .A(n6031), .B(n6032), .Z(n5687) );
  XNOR U7500 ( .A(round_reg[1429]), .B(round_reg[1109]), .Z(n6032) );
  XOR U7501 ( .A(round_reg[149]), .B(n6033), .Z(n6031) );
  XOR U7502 ( .A(round_reg[789]), .B(round_reg[469]), .Z(n6033) );
  XNOR U7503 ( .A(n6034), .B(n6035), .Z(n4985) );
  XNOR U7504 ( .A(round_reg[20]), .B(round_reg[1300]), .Z(n6035) );
  XOR U7505 ( .A(round_reg[340]), .B(n6036), .Z(n6034) );
  XOR U7506 ( .A(round_reg[980]), .B(round_reg[660]), .Z(n6036) );
  XNOR U7507 ( .A(round_reg[989]), .B(n4334), .Z(n4467) );
  XOR U7508 ( .A(n5330), .B(n5587), .Z(n4334) );
  XNOR U7509 ( .A(n6037), .B(n6038), .Z(n5587) );
  XNOR U7510 ( .A(round_reg[1564]), .B(round_reg[1244]), .Z(n6038) );
  XOR U7511 ( .A(round_reg[284]), .B(n6039), .Z(n6037) );
  XOR U7512 ( .A(round_reg[924]), .B(round_reg[604]), .Z(n6039) );
  XOR U7513 ( .A(n6040), .B(n6041), .Z(n5330) );
  XNOR U7514 ( .A(round_reg[1373]), .B(round_reg[1053]), .Z(n6041) );
  XOR U7515 ( .A(round_reg[413]), .B(n6042), .Z(n6040) );
  XOR U7516 ( .A(round_reg[93]), .B(round_reg[733]), .Z(n6042) );
  XOR U7517 ( .A(n6043), .B(n4899), .Z(out[1008]) );
  XOR U7518 ( .A(round_reg[179]), .B(n2138), .Z(n4899) );
  XNOR U7519 ( .A(n4809), .B(n4868), .Z(n2138) );
  XNOR U7520 ( .A(n6044), .B(n6045), .Z(n4868) );
  XNOR U7521 ( .A(round_reg[1523]), .B(round_reg[1203]), .Z(n6045) );
  XOR U7522 ( .A(round_reg[243]), .B(n6046), .Z(n6044) );
  XOR U7523 ( .A(round_reg[883]), .B(round_reg[563]), .Z(n6046) );
  XOR U7524 ( .A(n6047), .B(n6048), .Z(n4809) );
  XNOR U7525 ( .A(round_reg[114]), .B(round_reg[1074]), .Z(n6048) );
  XOR U7526 ( .A(round_reg[1394]), .B(n6049), .Z(n6047) );
  XOR U7527 ( .A(round_reg[754]), .B(round_reg[434]), .Z(n6049) );
  ANDN U7528 ( .B(n4471), .A(n4469), .Z(n6043) );
  XNOR U7529 ( .A(round_reg[1364]), .B(n1774), .Z(n4469) );
  XOR U7530 ( .A(n6050), .B(n6051), .Z(n5702) );
  XNOR U7531 ( .A(round_reg[1428]), .B(round_reg[1108]), .Z(n6051) );
  XOR U7532 ( .A(round_reg[148]), .B(n6052), .Z(n6050) );
  XOR U7533 ( .A(round_reg[788]), .B(round_reg[468]), .Z(n6052) );
  XNOR U7534 ( .A(n6053), .B(n6054), .Z(n4988) );
  XNOR U7535 ( .A(round_reg[19]), .B(round_reg[1299]), .Z(n6054) );
  XOR U7536 ( .A(round_reg[339]), .B(n6055), .Z(n6053) );
  XOR U7537 ( .A(round_reg[979]), .B(round_reg[659]), .Z(n6055) );
  XOR U7538 ( .A(round_reg[988]), .B(n2014), .Z(n4471) );
  XNOR U7539 ( .A(n5343), .B(n5602), .Z(n2014) );
  XNOR U7540 ( .A(n6056), .B(n6057), .Z(n5602) );
  XNOR U7541 ( .A(round_reg[1563]), .B(round_reg[1243]), .Z(n6057) );
  XOR U7542 ( .A(round_reg[283]), .B(n6058), .Z(n6056) );
  XOR U7543 ( .A(round_reg[923]), .B(round_reg[603]), .Z(n6058) );
  XOR U7544 ( .A(n6059), .B(n6060), .Z(n5343) );
  XNOR U7545 ( .A(round_reg[1372]), .B(round_reg[1052]), .Z(n6060) );
  XOR U7546 ( .A(round_reg[412]), .B(n6061), .Z(n6059) );
  XOR U7547 ( .A(round_reg[92]), .B(round_reg[732]), .Z(n6061) );
  XOR U7548 ( .A(n6062), .B(n4903), .Z(out[1007]) );
  XOR U7549 ( .A(round_reg[178]), .B(n2142), .Z(n4903) );
  XNOR U7550 ( .A(n4813), .B(n4872), .Z(n2142) );
  XNOR U7551 ( .A(n6063), .B(n6064), .Z(n4872) );
  XNOR U7552 ( .A(round_reg[1522]), .B(round_reg[1202]), .Z(n6064) );
  XOR U7553 ( .A(round_reg[242]), .B(n6065), .Z(n6063) );
  XOR U7554 ( .A(round_reg[882]), .B(round_reg[562]), .Z(n6065) );
  XOR U7555 ( .A(n6066), .B(n6067), .Z(n4813) );
  XNOR U7556 ( .A(round_reg[113]), .B(round_reg[1073]), .Z(n6067) );
  XOR U7557 ( .A(round_reg[1393]), .B(n6068), .Z(n6066) );
  XOR U7558 ( .A(round_reg[753]), .B(round_reg[433]), .Z(n6068) );
  ANDN U7559 ( .B(n4475), .A(n4473), .Z(n6062) );
  XNOR U7560 ( .A(round_reg[1363]), .B(n1777), .Z(n4473) );
  XOR U7561 ( .A(n6069), .B(n6070), .Z(n5717) );
  XNOR U7562 ( .A(round_reg[1427]), .B(round_reg[1107]), .Z(n6070) );
  XOR U7563 ( .A(round_reg[147]), .B(n6071), .Z(n6069) );
  XOR U7564 ( .A(round_reg[787]), .B(round_reg[467]), .Z(n6071) );
  XNOR U7565 ( .A(n6072), .B(n6073), .Z(n4992) );
  XNOR U7566 ( .A(round_reg[18]), .B(round_reg[1298]), .Z(n6073) );
  XOR U7567 ( .A(round_reg[338]), .B(n6074), .Z(n6072) );
  XOR U7568 ( .A(round_reg[978]), .B(round_reg[658]), .Z(n6074) );
  XOR U7569 ( .A(round_reg[987]), .B(n2020), .Z(n4475) );
  XNOR U7570 ( .A(n5365), .B(n5617), .Z(n2020) );
  XNOR U7571 ( .A(n6075), .B(n6076), .Z(n5617) );
  XNOR U7572 ( .A(round_reg[1562]), .B(round_reg[1242]), .Z(n6076) );
  XOR U7573 ( .A(round_reg[282]), .B(n6077), .Z(n6075) );
  XOR U7574 ( .A(round_reg[922]), .B(round_reg[602]), .Z(n6077) );
  XOR U7575 ( .A(n6078), .B(n6079), .Z(n5365) );
  XNOR U7576 ( .A(round_reg[1371]), .B(round_reg[1051]), .Z(n6079) );
  XOR U7577 ( .A(round_reg[411]), .B(n6080), .Z(n6078) );
  XOR U7578 ( .A(round_reg[91]), .B(round_reg[731]), .Z(n6080) );
  XOR U7579 ( .A(n6081), .B(n4907), .Z(out[1006]) );
  XOR U7580 ( .A(round_reg[177]), .B(n2146), .Z(n4907) );
  XNOR U7581 ( .A(n4817), .B(n4876), .Z(n2146) );
  XNOR U7582 ( .A(n6082), .B(n6083), .Z(n4876) );
  XNOR U7583 ( .A(round_reg[1521]), .B(round_reg[1201]), .Z(n6083) );
  XOR U7584 ( .A(round_reg[241]), .B(n6084), .Z(n6082) );
  XOR U7585 ( .A(round_reg[881]), .B(round_reg[561]), .Z(n6084) );
  XOR U7586 ( .A(n6085), .B(n6086), .Z(n4817) );
  XNOR U7587 ( .A(round_reg[112]), .B(round_reg[1072]), .Z(n6086) );
  XOR U7588 ( .A(round_reg[1392]), .B(n6087), .Z(n6085) );
  XOR U7589 ( .A(round_reg[752]), .B(round_reg[432]), .Z(n6087) );
  ANDN U7590 ( .B(n4479), .A(n4477), .Z(n6081) );
  XOR U7591 ( .A(round_reg[1362]), .B(n1780), .Z(n4477) );
  XOR U7592 ( .A(n5732), .B(n4994), .Z(n1780) );
  XOR U7593 ( .A(n6088), .B(n6089), .Z(n4994) );
  XNOR U7594 ( .A(round_reg[17]), .B(round_reg[1297]), .Z(n6089) );
  XOR U7595 ( .A(round_reg[337]), .B(n6090), .Z(n6088) );
  XOR U7596 ( .A(round_reg[977]), .B(round_reg[657]), .Z(n6090) );
  XOR U7597 ( .A(n6091), .B(n6092), .Z(n5732) );
  XNOR U7598 ( .A(round_reg[1426]), .B(round_reg[1106]), .Z(n6092) );
  XOR U7599 ( .A(round_reg[146]), .B(n6093), .Z(n6091) );
  XOR U7600 ( .A(round_reg[786]), .B(round_reg[466]), .Z(n6093) );
  XOR U7601 ( .A(round_reg[986]), .B(n2022), .Z(n4479) );
  XNOR U7602 ( .A(n5376), .B(n5632), .Z(n2022) );
  XNOR U7603 ( .A(n6094), .B(n6095), .Z(n5632) );
  XNOR U7604 ( .A(round_reg[1561]), .B(round_reg[1241]), .Z(n6095) );
  XOR U7605 ( .A(round_reg[281]), .B(n6096), .Z(n6094) );
  XOR U7606 ( .A(round_reg[921]), .B(round_reg[601]), .Z(n6096) );
  XOR U7607 ( .A(n6097), .B(n6098), .Z(n5376) );
  XNOR U7608 ( .A(round_reg[1370]), .B(round_reg[1050]), .Z(n6098) );
  XOR U7609 ( .A(round_reg[410]), .B(n6099), .Z(n6097) );
  XOR U7610 ( .A(round_reg[90]), .B(round_reg[730]), .Z(n6099) );
  XOR U7611 ( .A(n6100), .B(n4911), .Z(out[1005]) );
  XOR U7612 ( .A(round_reg[176]), .B(n2150), .Z(n4911) );
  XNOR U7613 ( .A(n4821), .B(n4880), .Z(n2150) );
  XNOR U7614 ( .A(n6101), .B(n6102), .Z(n4880) );
  XNOR U7615 ( .A(round_reg[1520]), .B(round_reg[1200]), .Z(n6102) );
  XOR U7616 ( .A(round_reg[240]), .B(n6103), .Z(n6101) );
  XOR U7617 ( .A(round_reg[880]), .B(round_reg[560]), .Z(n6103) );
  XOR U7618 ( .A(n6104), .B(n6105), .Z(n4821) );
  XNOR U7619 ( .A(round_reg[111]), .B(round_reg[1071]), .Z(n6105) );
  XOR U7620 ( .A(round_reg[1391]), .B(n6106), .Z(n6104) );
  XOR U7621 ( .A(round_reg[751]), .B(round_reg[431]), .Z(n6106) );
  ANDN U7622 ( .B(n4483), .A(n4481), .Z(n6100) );
  XNOR U7623 ( .A(round_reg[1361]), .B(n4243), .Z(n4481) );
  XNOR U7624 ( .A(n6107), .B(n6108), .Z(n5049) );
  XNOR U7625 ( .A(round_reg[1425]), .B(round_reg[1105]), .Z(n6108) );
  XOR U7626 ( .A(round_reg[145]), .B(n6109), .Z(n6107) );
  XOR U7627 ( .A(round_reg[785]), .B(round_reg[465]), .Z(n6109) );
  XNOR U7628 ( .A(n6110), .B(n6111), .Z(n4998) );
  XNOR U7629 ( .A(round_reg[16]), .B(round_reg[1296]), .Z(n6111) );
  XOR U7630 ( .A(round_reg[336]), .B(n6112), .Z(n6110) );
  XOR U7631 ( .A(round_reg[976]), .B(round_reg[656]), .Z(n6112) );
  XOR U7632 ( .A(round_reg[985]), .B(n2025), .Z(n4483) );
  XNOR U7633 ( .A(n5387), .B(n5658), .Z(n2025) );
  XNOR U7634 ( .A(n6113), .B(n6114), .Z(n5658) );
  XNOR U7635 ( .A(round_reg[1560]), .B(round_reg[1240]), .Z(n6114) );
  XOR U7636 ( .A(round_reg[280]), .B(n6115), .Z(n6113) );
  XOR U7637 ( .A(round_reg[920]), .B(round_reg[600]), .Z(n6115) );
  XOR U7638 ( .A(n6116), .B(n6117), .Z(n5387) );
  XNOR U7639 ( .A(round_reg[1369]), .B(round_reg[1049]), .Z(n6117) );
  XOR U7640 ( .A(round_reg[409]), .B(n6118), .Z(n6116) );
  XOR U7641 ( .A(round_reg[89]), .B(round_reg[729]), .Z(n6118) );
  XOR U7642 ( .A(n6119), .B(n4915), .Z(out[1004]) );
  XOR U7643 ( .A(round_reg[175]), .B(n2154), .Z(n4915) );
  XNOR U7644 ( .A(n4825), .B(n4886), .Z(n2154) );
  XNOR U7645 ( .A(n6120), .B(n6121), .Z(n4886) );
  XNOR U7646 ( .A(round_reg[1519]), .B(round_reg[1199]), .Z(n6121) );
  XOR U7647 ( .A(round_reg[239]), .B(n6122), .Z(n6120) );
  XOR U7648 ( .A(round_reg[879]), .B(round_reg[559]), .Z(n6122) );
  XOR U7649 ( .A(n6123), .B(n6124), .Z(n4825) );
  XNOR U7650 ( .A(round_reg[110]), .B(round_reg[1070]), .Z(n6124) );
  XOR U7651 ( .A(round_reg[1390]), .B(n6125), .Z(n6123) );
  XOR U7652 ( .A(round_reg[750]), .B(round_reg[430]), .Z(n6125) );
  ANDN U7653 ( .B(n4487), .A(n4485), .Z(n6119) );
  XNOR U7654 ( .A(round_reg[1360]), .B(n4245), .Z(n4485) );
  XOR U7655 ( .A(n6126), .B(n5054), .Z(n4245) );
  XNOR U7656 ( .A(n6127), .B(n6128), .Z(n5054) );
  XNOR U7657 ( .A(round_reg[1424]), .B(round_reg[1104]), .Z(n6128) );
  XOR U7658 ( .A(round_reg[144]), .B(n6129), .Z(n6127) );
  XOR U7659 ( .A(round_reg[784]), .B(round_reg[464]), .Z(n6129) );
  IV U7660 ( .A(n5001), .Z(n6126) );
  XNOR U7661 ( .A(n6130), .B(n6131), .Z(n5001) );
  XNOR U7662 ( .A(round_reg[15]), .B(round_reg[1295]), .Z(n6131) );
  XOR U7663 ( .A(round_reg[335]), .B(n6132), .Z(n6130) );
  XOR U7664 ( .A(round_reg[975]), .B(round_reg[655]), .Z(n6132) );
  XOR U7665 ( .A(round_reg[984]), .B(n2028), .Z(n4487) );
  XNOR U7666 ( .A(n5400), .B(n5673), .Z(n2028) );
  XNOR U7667 ( .A(n6133), .B(n6134), .Z(n5673) );
  XNOR U7668 ( .A(round_reg[1559]), .B(round_reg[1239]), .Z(n6134) );
  XOR U7669 ( .A(round_reg[279]), .B(n6135), .Z(n6133) );
  XOR U7670 ( .A(round_reg[919]), .B(round_reg[599]), .Z(n6135) );
  XOR U7671 ( .A(n6136), .B(n6137), .Z(n5400) );
  XNOR U7672 ( .A(round_reg[1368]), .B(round_reg[1048]), .Z(n6137) );
  XOR U7673 ( .A(round_reg[408]), .B(n6138), .Z(n6136) );
  XOR U7674 ( .A(round_reg[88]), .B(round_reg[728]), .Z(n6138) );
  XOR U7675 ( .A(n6139), .B(n4919), .Z(out[1003]) );
  XOR U7676 ( .A(round_reg[174]), .B(n2158), .Z(n4919) );
  XNOR U7677 ( .A(n4829), .B(n4890), .Z(n2158) );
  XNOR U7678 ( .A(n6140), .B(n6141), .Z(n4890) );
  XNOR U7679 ( .A(round_reg[1518]), .B(round_reg[1198]), .Z(n6141) );
  XOR U7680 ( .A(round_reg[238]), .B(n6142), .Z(n6140) );
  XOR U7681 ( .A(round_reg[878]), .B(round_reg[558]), .Z(n6142) );
  XOR U7682 ( .A(n6143), .B(n6144), .Z(n4829) );
  XNOR U7683 ( .A(round_reg[109]), .B(round_reg[1069]), .Z(n6144) );
  XOR U7684 ( .A(round_reg[1389]), .B(n6145), .Z(n6143) );
  XOR U7685 ( .A(round_reg[749]), .B(round_reg[429]), .Z(n6145) );
  ANDN U7686 ( .B(n4493), .A(n4491), .Z(n6139) );
  XNOR U7687 ( .A(round_reg[1359]), .B(n4247), .Z(n4491) );
  XOR U7688 ( .A(n6146), .B(n5059), .Z(n4247) );
  XNOR U7689 ( .A(n6147), .B(n6148), .Z(n5059) );
  XNOR U7690 ( .A(round_reg[1423]), .B(round_reg[1103]), .Z(n6148) );
  XOR U7691 ( .A(round_reg[143]), .B(n6149), .Z(n6147) );
  XOR U7692 ( .A(round_reg[783]), .B(round_reg[463]), .Z(n6149) );
  IV U7693 ( .A(n5004), .Z(n6146) );
  XNOR U7694 ( .A(n6150), .B(n6151), .Z(n5004) );
  XNOR U7695 ( .A(round_reg[14]), .B(round_reg[1294]), .Z(n6151) );
  XOR U7696 ( .A(round_reg[334]), .B(n6152), .Z(n6150) );
  XOR U7697 ( .A(round_reg[974]), .B(round_reg[654]), .Z(n6152) );
  XOR U7698 ( .A(round_reg[983]), .B(n2031), .Z(n4493) );
  XNOR U7699 ( .A(n5413), .B(n5688), .Z(n2031) );
  XNOR U7700 ( .A(n6153), .B(n6154), .Z(n5688) );
  XNOR U7701 ( .A(round_reg[1558]), .B(round_reg[1238]), .Z(n6154) );
  XOR U7702 ( .A(round_reg[278]), .B(n6155), .Z(n6153) );
  XOR U7703 ( .A(round_reg[918]), .B(round_reg[598]), .Z(n6155) );
  XOR U7704 ( .A(n6156), .B(n6157), .Z(n5413) );
  XNOR U7705 ( .A(round_reg[1367]), .B(round_reg[1047]), .Z(n6157) );
  XOR U7706 ( .A(round_reg[407]), .B(n6158), .Z(n6156) );
  XOR U7707 ( .A(round_reg[87]), .B(round_reg[727]), .Z(n6158) );
  XOR U7708 ( .A(n6159), .B(n4923), .Z(out[1002]) );
  XOR U7709 ( .A(round_reg[173]), .B(n2162), .Z(n4923) );
  XNOR U7710 ( .A(n4833), .B(n4894), .Z(n2162) );
  XNOR U7711 ( .A(n6160), .B(n6161), .Z(n4894) );
  XNOR U7712 ( .A(round_reg[1517]), .B(round_reg[1197]), .Z(n6161) );
  XOR U7713 ( .A(round_reg[237]), .B(n6162), .Z(n6160) );
  XOR U7714 ( .A(round_reg[877]), .B(round_reg[557]), .Z(n6162) );
  XOR U7715 ( .A(n6163), .B(n6164), .Z(n4833) );
  XNOR U7716 ( .A(round_reg[108]), .B(round_reg[1068]), .Z(n6164) );
  XOR U7717 ( .A(round_reg[1388]), .B(n6165), .Z(n6163) );
  XOR U7718 ( .A(round_reg[748]), .B(round_reg[428]), .Z(n6165) );
  ANDN U7719 ( .B(n4497), .A(n4495), .Z(n6159) );
  XNOR U7720 ( .A(round_reg[1358]), .B(n4251), .Z(n4495) );
  XOR U7721 ( .A(n6166), .B(n5064), .Z(n4251) );
  XNOR U7722 ( .A(n6167), .B(n6168), .Z(n5064) );
  XNOR U7723 ( .A(round_reg[1422]), .B(round_reg[1102]), .Z(n6168) );
  XOR U7724 ( .A(round_reg[142]), .B(n6169), .Z(n6167) );
  XOR U7725 ( .A(round_reg[782]), .B(round_reg[462]), .Z(n6169) );
  IV U7726 ( .A(n5007), .Z(n6166) );
  XNOR U7727 ( .A(n6170), .B(n6171), .Z(n5007) );
  XNOR U7728 ( .A(round_reg[13]), .B(round_reg[1293]), .Z(n6171) );
  XOR U7729 ( .A(round_reg[333]), .B(n6172), .Z(n6170) );
  XOR U7730 ( .A(round_reg[973]), .B(round_reg[653]), .Z(n6172) );
  XOR U7731 ( .A(round_reg[982]), .B(n2034), .Z(n4497) );
  XNOR U7732 ( .A(n5426), .B(n5703), .Z(n2034) );
  XNOR U7733 ( .A(n6173), .B(n6174), .Z(n5703) );
  XNOR U7734 ( .A(round_reg[1557]), .B(round_reg[1237]), .Z(n6174) );
  XOR U7735 ( .A(round_reg[277]), .B(n6175), .Z(n6173) );
  XOR U7736 ( .A(round_reg[917]), .B(round_reg[597]), .Z(n6175) );
  XOR U7737 ( .A(n6176), .B(n6177), .Z(n5426) );
  XNOR U7738 ( .A(round_reg[1366]), .B(round_reg[1046]), .Z(n6177) );
  XOR U7739 ( .A(round_reg[406]), .B(n6178), .Z(n6176) );
  XOR U7740 ( .A(round_reg[86]), .B(round_reg[726]), .Z(n6178) );
  XOR U7741 ( .A(n6179), .B(n4929), .Z(out[1001]) );
  XOR U7742 ( .A(round_reg[172]), .B(n2166), .Z(n4929) );
  XNOR U7743 ( .A(n5753), .B(n4898), .Z(n2166) );
  XNOR U7744 ( .A(n6180), .B(n6181), .Z(n4898) );
  XNOR U7745 ( .A(round_reg[1516]), .B(round_reg[1196]), .Z(n6181) );
  XOR U7746 ( .A(round_reg[236]), .B(n6182), .Z(n6180) );
  XOR U7747 ( .A(round_reg[876]), .B(round_reg[556]), .Z(n6182) );
  XOR U7748 ( .A(n6183), .B(n6184), .Z(n5753) );
  XNOR U7749 ( .A(round_reg[107]), .B(round_reg[1067]), .Z(n6184) );
  XOR U7750 ( .A(round_reg[1387]), .B(n6185), .Z(n6183) );
  XOR U7751 ( .A(round_reg[747]), .B(round_reg[427]), .Z(n6185) );
  ANDN U7752 ( .B(n4501), .A(n4499), .Z(n6179) );
  XNOR U7753 ( .A(round_reg[1357]), .B(n4253), .Z(n4499) );
  XOR U7754 ( .A(n6186), .B(n5069), .Z(n4253) );
  XNOR U7755 ( .A(n6187), .B(n6188), .Z(n5069) );
  XNOR U7756 ( .A(round_reg[141]), .B(round_reg[1101]), .Z(n6188) );
  XOR U7757 ( .A(round_reg[1421]), .B(n6189), .Z(n6187) );
  XOR U7758 ( .A(round_reg[781]), .B(round_reg[461]), .Z(n6189) );
  IV U7759 ( .A(n5010), .Z(n6186) );
  XNOR U7760 ( .A(n6190), .B(n6191), .Z(n5010) );
  XNOR U7761 ( .A(round_reg[12]), .B(round_reg[1292]), .Z(n6191) );
  XOR U7762 ( .A(round_reg[332]), .B(n6192), .Z(n6190) );
  XOR U7763 ( .A(round_reg[972]), .B(round_reg[652]), .Z(n6192) );
  XOR U7764 ( .A(round_reg[981]), .B(n2037), .Z(n4501) );
  XNOR U7765 ( .A(n5439), .B(n5718), .Z(n2037) );
  XNOR U7766 ( .A(n6193), .B(n6194), .Z(n5718) );
  XNOR U7767 ( .A(round_reg[1556]), .B(round_reg[1236]), .Z(n6194) );
  XOR U7768 ( .A(round_reg[276]), .B(n6195), .Z(n6193) );
  XOR U7769 ( .A(round_reg[916]), .B(round_reg[596]), .Z(n6195) );
  XOR U7770 ( .A(n6196), .B(n6197), .Z(n5439) );
  XNOR U7771 ( .A(round_reg[1365]), .B(round_reg[1045]), .Z(n6197) );
  XOR U7772 ( .A(round_reg[405]), .B(n6198), .Z(n6196) );
  XOR U7773 ( .A(round_reg[85]), .B(round_reg[725]), .Z(n6198) );
  XOR U7774 ( .A(n6199), .B(n4933), .Z(out[1000]) );
  XOR U7775 ( .A(round_reg[171]), .B(n2174), .Z(n4933) );
  XNOR U7776 ( .A(n5768), .B(n4902), .Z(n2174) );
  XNOR U7777 ( .A(n6200), .B(n6201), .Z(n4902) );
  XNOR U7778 ( .A(round_reg[1515]), .B(round_reg[1195]), .Z(n6201) );
  XOR U7779 ( .A(round_reg[235]), .B(n6202), .Z(n6200) );
  XOR U7780 ( .A(round_reg[875]), .B(round_reg[555]), .Z(n6202) );
  XOR U7781 ( .A(n6203), .B(n6204), .Z(n5768) );
  XNOR U7782 ( .A(round_reg[106]), .B(round_reg[1066]), .Z(n6204) );
  XOR U7783 ( .A(round_reg[1386]), .B(n6205), .Z(n6203) );
  XOR U7784 ( .A(round_reg[746]), .B(round_reg[426]), .Z(n6205) );
  ANDN U7785 ( .B(n4505), .A(n4503), .Z(n6199) );
  XNOR U7786 ( .A(round_reg[1356]), .B(n4255), .Z(n4503) );
  XOR U7787 ( .A(n6206), .B(n5074), .Z(n4255) );
  XNOR U7788 ( .A(n6207), .B(n6208), .Z(n5074) );
  XNOR U7789 ( .A(round_reg[140]), .B(round_reg[1100]), .Z(n6208) );
  XOR U7790 ( .A(round_reg[1420]), .B(n6209), .Z(n6207) );
  XOR U7791 ( .A(round_reg[780]), .B(round_reg[460]), .Z(n6209) );
  IV U7792 ( .A(n5013), .Z(n6206) );
  XNOR U7793 ( .A(n6210), .B(n6211), .Z(n5013) );
  XNOR U7794 ( .A(round_reg[1291]), .B(round_reg[11]), .Z(n6211) );
  XOR U7795 ( .A(round_reg[331]), .B(n6212), .Z(n6210) );
  XOR U7796 ( .A(round_reg[971]), .B(round_reg[651]), .Z(n6212) );
  XOR U7797 ( .A(round_reg[980]), .B(n2040), .Z(n4505) );
  XNOR U7798 ( .A(n5450), .B(n5733), .Z(n2040) );
  XNOR U7799 ( .A(n6213), .B(n6214), .Z(n5733) );
  XNOR U7800 ( .A(round_reg[1555]), .B(round_reg[1235]), .Z(n6214) );
  XOR U7801 ( .A(round_reg[275]), .B(n6215), .Z(n6213) );
  XOR U7802 ( .A(round_reg[915]), .B(round_reg[595]), .Z(n6215) );
  XOR U7803 ( .A(n6216), .B(n6217), .Z(n5450) );
  XNOR U7804 ( .A(round_reg[1364]), .B(round_reg[1044]), .Z(n6217) );
  XOR U7805 ( .A(round_reg[404]), .B(n6218), .Z(n6216) );
  XOR U7806 ( .A(round_reg[84]), .B(round_reg[724]), .Z(n6218) );
  XOR U7807 ( .A(n6219), .B(n2347), .Z(out[0]) );
  XOR U7808 ( .A(round_reg[254]), .B(n2990), .Z(n2347) );
  IV U7809 ( .A(n2107), .Z(n2990) );
  XOR U7810 ( .A(n5369), .B(n4751), .Z(n2107) );
  XNOR U7811 ( .A(n6220), .B(n6221), .Z(n4751) );
  XNOR U7812 ( .A(round_reg[1598]), .B(round_reg[1278]), .Z(n6221) );
  XOR U7813 ( .A(round_reg[318]), .B(n6222), .Z(n6220) );
  XOR U7814 ( .A(round_reg[958]), .B(round_reg[638]), .Z(n6222) );
  XOR U7815 ( .A(n6223), .B(n6224), .Z(n5369) );
  XNOR U7816 ( .A(round_reg[1469]), .B(round_reg[1149]), .Z(n6224) );
  XOR U7817 ( .A(round_reg[189]), .B(n6225), .Z(n6223) );
  XOR U7818 ( .A(round_reg[829]), .B(round_reg[509]), .Z(n6225) );
  AND U7819 ( .A(n3418), .B(n3416), .Z(n6219) );
  XNOR U7820 ( .A(round_reg[1410]), .B(n2354), .Z(n3416) );
  XNOR U7821 ( .A(n4742), .B(n5045), .Z(n2354) );
  XNOR U7822 ( .A(n6226), .B(n6227), .Z(n5045) );
  XNOR U7823 ( .A(round_reg[1474]), .B(round_reg[1154]), .Z(n6227) );
  XOR U7824 ( .A(round_reg[194]), .B(n6228), .Z(n6226) );
  XOR U7825 ( .A(round_reg[834]), .B(round_reg[514]), .Z(n6228) );
  XOR U7826 ( .A(n6229), .B(n6230), .Z(n4742) );
  XNOR U7827 ( .A(round_reg[1345]), .B(round_reg[1025]), .Z(n6230) );
  XOR U7828 ( .A(round_reg[385]), .B(n6231), .Z(n6229) );
  XOR U7829 ( .A(round_reg[705]), .B(round_reg[65]), .Z(n6231) );
  XOR U7830 ( .A(round_reg[1033]), .B(n1811), .Z(n3418) );
  XOR U7831 ( .A(n5092), .B(n5024), .Z(n1811) );
  XOR U7832 ( .A(n6232), .B(n6233), .Z(n5024) );
  XNOR U7833 ( .A(round_reg[328]), .B(round_reg[1288]), .Z(n6233) );
  XOR U7834 ( .A(round_reg[648]), .B(n6234), .Z(n6232) );
  XOR U7835 ( .A(round_reg[968]), .B(round_reg[8]), .Z(n6234) );
  XOR U7836 ( .A(n6235), .B(n6236), .Z(n5092) );
  XNOR U7837 ( .A(round_reg[137]), .B(round_reg[1097]), .Z(n6236) );
  XOR U7838 ( .A(round_reg[1417]), .B(n6237), .Z(n6235) );
  XOR U7839 ( .A(round_reg[777]), .B(round_reg[457]), .Z(n6237) );
  IV U7840 ( .A(init), .Z(n1050) );
endmodule

