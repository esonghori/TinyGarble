
module sha3_seq_CC24 ( clk, rst, g_init, e_init, o );
  input [287:0] g_init;
  input [287:0] e_init;
  output [1599:0] o;
  input clk, rst;
  wire   init, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257;
  wire   [23:0] rc_i;
  wire   [1599:0] round_reg;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .I(1'b0), .Q(init) );
  DFF \rc_i_reg[0]  ( .D(n1050), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[0])
         );
  DFF \rc_i_reg[1]  ( .D(rc_i[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[1])
         );
  DFF \rc_i_reg[2]  ( .D(rc_i[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[2])
         );
  DFF \rc_i_reg[3]  ( .D(rc_i[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[3])
         );
  DFF \rc_i_reg[4]  ( .D(rc_i[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[4])
         );
  DFF \rc_i_reg[5]  ( .D(rc_i[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[5])
         );
  DFF \rc_i_reg[6]  ( .D(rc_i[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[6])
         );
  DFF \rc_i_reg[7]  ( .D(rc_i[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[7])
         );
  DFF \rc_i_reg[8]  ( .D(rc_i[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[8])
         );
  DFF \rc_i_reg[9]  ( .D(rc_i[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(rc_i[9])
         );
  DFF \rc_i_reg[10]  ( .D(rc_i[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[10]) );
  DFF \rc_i_reg[11]  ( .D(rc_i[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[11]) );
  DFF \rc_i_reg[12]  ( .D(rc_i[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[12]) );
  DFF \rc_i_reg[13]  ( .D(rc_i[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[13]) );
  DFF \rc_i_reg[14]  ( .D(rc_i[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[14]) );
  DFF \rc_i_reg[15]  ( .D(rc_i[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[15]) );
  DFF \rc_i_reg[16]  ( .D(rc_i[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[16]) );
  DFF \rc_i_reg[17]  ( .D(rc_i[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[17]) );
  DFF \rc_i_reg[18]  ( .D(rc_i[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[18]) );
  DFF \rc_i_reg[19]  ( .D(rc_i[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[19]) );
  DFF \rc_i_reg[20]  ( .D(rc_i[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[20]) );
  DFF \rc_i_reg[21]  ( .D(rc_i[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[21]) );
  DFF \rc_i_reg[22]  ( .D(rc_i[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[22]) );
  DFF \rc_i_reg[23]  ( .D(rc_i[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        rc_i[23]) );
  DFF \round_reg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .I(g_init[0]), .Q(
        round_reg[0]) );
  DFF \round_reg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .I(g_init[1]), .Q(
        round_reg[1]) );
  DFF \round_reg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .I(g_init[2]), .Q(
        round_reg[2]) );
  DFF \round_reg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .I(g_init[3]), .Q(
        round_reg[3]) );
  DFF \round_reg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .I(g_init[4]), .Q(
        round_reg[4]) );
  DFF \round_reg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .I(g_init[5]), .Q(
        round_reg[5]) );
  DFF \round_reg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .I(g_init[6]), .Q(
        round_reg[6]) );
  DFF \round_reg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .I(g_init[7]), .Q(
        round_reg[7]) );
  DFF \round_reg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .I(g_init[8]), .Q(
        round_reg[8]) );
  DFF \round_reg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .I(g_init[9]), .Q(
        round_reg[9]) );
  DFF \round_reg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .I(g_init[10]), 
        .Q(round_reg[10]) );
  DFF \round_reg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .I(g_init[11]), 
        .Q(round_reg[11]) );
  DFF \round_reg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .I(g_init[12]), 
        .Q(round_reg[12]) );
  DFF \round_reg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .I(g_init[13]), 
        .Q(round_reg[13]) );
  DFF \round_reg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .I(g_init[14]), 
        .Q(round_reg[14]) );
  DFF \round_reg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .I(g_init[15]), 
        .Q(round_reg[15]) );
  DFF \round_reg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .I(g_init[16]), 
        .Q(round_reg[16]) );
  DFF \round_reg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .I(g_init[17]), 
        .Q(round_reg[17]) );
  DFF \round_reg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .I(g_init[18]), 
        .Q(round_reg[18]) );
  DFF \round_reg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .I(g_init[19]), 
        .Q(round_reg[19]) );
  DFF \round_reg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .I(g_init[20]), 
        .Q(round_reg[20]) );
  DFF \round_reg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .I(g_init[21]), 
        .Q(round_reg[21]) );
  DFF \round_reg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .I(g_init[22]), 
        .Q(round_reg[22]) );
  DFF \round_reg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .I(g_init[23]), 
        .Q(round_reg[23]) );
  DFF \round_reg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .I(g_init[24]), 
        .Q(round_reg[24]) );
  DFF \round_reg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .I(g_init[25]), 
        .Q(round_reg[25]) );
  DFF \round_reg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .I(g_init[26]), 
        .Q(round_reg[26]) );
  DFF \round_reg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .I(g_init[27]), 
        .Q(round_reg[27]) );
  DFF \round_reg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .I(g_init[28]), 
        .Q(round_reg[28]) );
  DFF \round_reg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .I(g_init[29]), 
        .Q(round_reg[29]) );
  DFF \round_reg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .I(g_init[30]), 
        .Q(round_reg[30]) );
  DFF \round_reg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .I(g_init[31]), 
        .Q(round_reg[31]) );
  DFF \round_reg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .I(g_init[32]), 
        .Q(round_reg[32]) );
  DFF \round_reg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .I(g_init[33]), 
        .Q(round_reg[33]) );
  DFF \round_reg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .I(g_init[34]), 
        .Q(round_reg[34]) );
  DFF \round_reg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .I(g_init[35]), 
        .Q(round_reg[35]) );
  DFF \round_reg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .I(g_init[36]), 
        .Q(round_reg[36]) );
  DFF \round_reg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .I(g_init[37]), 
        .Q(round_reg[37]) );
  DFF \round_reg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .I(g_init[38]), 
        .Q(round_reg[38]) );
  DFF \round_reg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .I(g_init[39]), 
        .Q(round_reg[39]) );
  DFF \round_reg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .I(g_init[40]), 
        .Q(round_reg[40]) );
  DFF \round_reg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .I(g_init[41]), 
        .Q(round_reg[41]) );
  DFF \round_reg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .I(g_init[42]), 
        .Q(round_reg[42]) );
  DFF \round_reg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .I(g_init[43]), 
        .Q(round_reg[43]) );
  DFF \round_reg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .I(g_init[44]), 
        .Q(round_reg[44]) );
  DFF \round_reg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .I(g_init[45]), 
        .Q(round_reg[45]) );
  DFF \round_reg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .I(g_init[46]), 
        .Q(round_reg[46]) );
  DFF \round_reg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .I(g_init[47]), 
        .Q(round_reg[47]) );
  DFF \round_reg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .I(g_init[48]), 
        .Q(round_reg[48]) );
  DFF \round_reg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .I(g_init[49]), 
        .Q(round_reg[49]) );
  DFF \round_reg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .I(g_init[50]), 
        .Q(round_reg[50]) );
  DFF \round_reg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .I(g_init[51]), 
        .Q(round_reg[51]) );
  DFF \round_reg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .I(g_init[52]), 
        .Q(round_reg[52]) );
  DFF \round_reg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .I(g_init[53]), 
        .Q(round_reg[53]) );
  DFF \round_reg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .I(g_init[54]), 
        .Q(round_reg[54]) );
  DFF \round_reg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .I(g_init[55]), 
        .Q(round_reg[55]) );
  DFF \round_reg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .I(g_init[56]), 
        .Q(round_reg[56]) );
  DFF \round_reg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .I(g_init[57]), 
        .Q(round_reg[57]) );
  DFF \round_reg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .I(g_init[58]), 
        .Q(round_reg[58]) );
  DFF \round_reg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .I(g_init[59]), 
        .Q(round_reg[59]) );
  DFF \round_reg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .I(g_init[60]), 
        .Q(round_reg[60]) );
  DFF \round_reg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .I(g_init[61]), 
        .Q(round_reg[61]) );
  DFF \round_reg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .I(g_init[62]), 
        .Q(round_reg[62]) );
  DFF \round_reg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .I(g_init[63]), 
        .Q(round_reg[63]) );
  DFF \round_reg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .I(g_init[64]), 
        .Q(round_reg[64]) );
  DFF \round_reg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .I(g_init[65]), 
        .Q(round_reg[65]) );
  DFF \round_reg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .I(g_init[66]), 
        .Q(round_reg[66]) );
  DFF \round_reg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .I(g_init[67]), 
        .Q(round_reg[67]) );
  DFF \round_reg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .I(g_init[68]), 
        .Q(round_reg[68]) );
  DFF \round_reg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .I(g_init[69]), 
        .Q(round_reg[69]) );
  DFF \round_reg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .I(g_init[70]), 
        .Q(round_reg[70]) );
  DFF \round_reg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .I(g_init[71]), 
        .Q(round_reg[71]) );
  DFF \round_reg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .I(g_init[72]), 
        .Q(round_reg[72]) );
  DFF \round_reg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .I(g_init[73]), 
        .Q(round_reg[73]) );
  DFF \round_reg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .I(g_init[74]), 
        .Q(round_reg[74]) );
  DFF \round_reg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .I(g_init[75]), 
        .Q(round_reg[75]) );
  DFF \round_reg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .I(g_init[76]), 
        .Q(round_reg[76]) );
  DFF \round_reg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .I(g_init[77]), 
        .Q(round_reg[77]) );
  DFF \round_reg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .I(g_init[78]), 
        .Q(round_reg[78]) );
  DFF \round_reg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .I(g_init[79]), 
        .Q(round_reg[79]) );
  DFF \round_reg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .I(g_init[80]), 
        .Q(round_reg[80]) );
  DFF \round_reg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .I(g_init[81]), 
        .Q(round_reg[81]) );
  DFF \round_reg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .I(g_init[82]), 
        .Q(round_reg[82]) );
  DFF \round_reg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .I(g_init[83]), 
        .Q(round_reg[83]) );
  DFF \round_reg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .I(g_init[84]), 
        .Q(round_reg[84]) );
  DFF \round_reg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .I(g_init[85]), 
        .Q(round_reg[85]) );
  DFF \round_reg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .I(g_init[86]), 
        .Q(round_reg[86]) );
  DFF \round_reg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .I(g_init[87]), 
        .Q(round_reg[87]) );
  DFF \round_reg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .I(g_init[88]), 
        .Q(round_reg[88]) );
  DFF \round_reg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .I(g_init[89]), 
        .Q(round_reg[89]) );
  DFF \round_reg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .I(g_init[90]), 
        .Q(round_reg[90]) );
  DFF \round_reg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .I(g_init[91]), 
        .Q(round_reg[91]) );
  DFF \round_reg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .I(g_init[92]), 
        .Q(round_reg[92]) );
  DFF \round_reg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .I(g_init[93]), 
        .Q(round_reg[93]) );
  DFF \round_reg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .I(g_init[94]), 
        .Q(round_reg[94]) );
  DFF \round_reg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .I(g_init[95]), 
        .Q(round_reg[95]) );
  DFF \round_reg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .I(g_init[96]), 
        .Q(round_reg[96]) );
  DFF \round_reg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .I(g_init[97]), 
        .Q(round_reg[97]) );
  DFF \round_reg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .I(g_init[98]), 
        .Q(round_reg[98]) );
  DFF \round_reg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .I(g_init[99]), 
        .Q(round_reg[99]) );
  DFF \round_reg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .I(g_init[100]), 
        .Q(round_reg[100]) );
  DFF \round_reg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .I(g_init[101]), 
        .Q(round_reg[101]) );
  DFF \round_reg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .I(g_init[102]), 
        .Q(round_reg[102]) );
  DFF \round_reg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .I(g_init[103]), 
        .Q(round_reg[103]) );
  DFF \round_reg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .I(g_init[104]), 
        .Q(round_reg[104]) );
  DFF \round_reg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .I(g_init[105]), 
        .Q(round_reg[105]) );
  DFF \round_reg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .I(g_init[106]), 
        .Q(round_reg[106]) );
  DFF \round_reg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .I(g_init[107]), 
        .Q(round_reg[107]) );
  DFF \round_reg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .I(g_init[108]), 
        .Q(round_reg[108]) );
  DFF \round_reg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .I(g_init[109]), 
        .Q(round_reg[109]) );
  DFF \round_reg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .I(g_init[110]), 
        .Q(round_reg[110]) );
  DFF \round_reg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .I(g_init[111]), 
        .Q(round_reg[111]) );
  DFF \round_reg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .I(g_init[112]), 
        .Q(round_reg[112]) );
  DFF \round_reg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .I(g_init[113]), 
        .Q(round_reg[113]) );
  DFF \round_reg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .I(g_init[114]), 
        .Q(round_reg[114]) );
  DFF \round_reg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .I(g_init[115]), 
        .Q(round_reg[115]) );
  DFF \round_reg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .I(g_init[116]), 
        .Q(round_reg[116]) );
  DFF \round_reg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .I(g_init[117]), 
        .Q(round_reg[117]) );
  DFF \round_reg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .I(g_init[118]), 
        .Q(round_reg[118]) );
  DFF \round_reg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .I(g_init[119]), 
        .Q(round_reg[119]) );
  DFF \round_reg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .I(g_init[120]), 
        .Q(round_reg[120]) );
  DFF \round_reg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .I(g_init[121]), 
        .Q(round_reg[121]) );
  DFF \round_reg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .I(g_init[122]), 
        .Q(round_reg[122]) );
  DFF \round_reg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .I(g_init[123]), 
        .Q(round_reg[123]) );
  DFF \round_reg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .I(g_init[124]), 
        .Q(round_reg[124]) );
  DFF \round_reg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .I(g_init[125]), 
        .Q(round_reg[125]) );
  DFF \round_reg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .I(g_init[126]), 
        .Q(round_reg[126]) );
  DFF \round_reg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .I(g_init[127]), 
        .Q(round_reg[127]) );
  DFF \round_reg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .I(g_init[128]), 
        .Q(round_reg[128]) );
  DFF \round_reg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .I(g_init[129]), 
        .Q(round_reg[129]) );
  DFF \round_reg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .I(g_init[130]), 
        .Q(round_reg[130]) );
  DFF \round_reg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .I(g_init[131]), 
        .Q(round_reg[131]) );
  DFF \round_reg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .I(g_init[132]), 
        .Q(round_reg[132]) );
  DFF \round_reg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .I(g_init[133]), 
        .Q(round_reg[133]) );
  DFF \round_reg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .I(g_init[134]), 
        .Q(round_reg[134]) );
  DFF \round_reg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .I(g_init[135]), 
        .Q(round_reg[135]) );
  DFF \round_reg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .I(g_init[136]), 
        .Q(round_reg[136]) );
  DFF \round_reg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .I(g_init[137]), 
        .Q(round_reg[137]) );
  DFF \round_reg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .I(g_init[138]), 
        .Q(round_reg[138]) );
  DFF \round_reg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .I(g_init[139]), 
        .Q(round_reg[139]) );
  DFF \round_reg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .I(g_init[140]), 
        .Q(round_reg[140]) );
  DFF \round_reg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .I(g_init[141]), 
        .Q(round_reg[141]) );
  DFF \round_reg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .I(g_init[142]), 
        .Q(round_reg[142]) );
  DFF \round_reg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .I(g_init[143]), 
        .Q(round_reg[143]) );
  DFF \round_reg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .I(g_init[144]), 
        .Q(round_reg[144]) );
  DFF \round_reg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .I(g_init[145]), 
        .Q(round_reg[145]) );
  DFF \round_reg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .I(g_init[146]), 
        .Q(round_reg[146]) );
  DFF \round_reg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .I(g_init[147]), 
        .Q(round_reg[147]) );
  DFF \round_reg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .I(g_init[148]), 
        .Q(round_reg[148]) );
  DFF \round_reg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .I(g_init[149]), 
        .Q(round_reg[149]) );
  DFF \round_reg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .I(g_init[150]), 
        .Q(round_reg[150]) );
  DFF \round_reg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .I(g_init[151]), 
        .Q(round_reg[151]) );
  DFF \round_reg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .I(g_init[152]), 
        .Q(round_reg[152]) );
  DFF \round_reg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .I(g_init[153]), 
        .Q(round_reg[153]) );
  DFF \round_reg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .I(g_init[154]), 
        .Q(round_reg[154]) );
  DFF \round_reg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .I(g_init[155]), 
        .Q(round_reg[155]) );
  DFF \round_reg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .I(g_init[156]), 
        .Q(round_reg[156]) );
  DFF \round_reg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .I(g_init[157]), 
        .Q(round_reg[157]) );
  DFF \round_reg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .I(g_init[158]), 
        .Q(round_reg[158]) );
  DFF \round_reg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .I(g_init[159]), 
        .Q(round_reg[159]) );
  DFF \round_reg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .I(g_init[160]), 
        .Q(round_reg[160]) );
  DFF \round_reg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .I(g_init[161]), 
        .Q(round_reg[161]) );
  DFF \round_reg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .I(g_init[162]), 
        .Q(round_reg[162]) );
  DFF \round_reg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .I(g_init[163]), 
        .Q(round_reg[163]) );
  DFF \round_reg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .I(g_init[164]), 
        .Q(round_reg[164]) );
  DFF \round_reg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .I(g_init[165]), 
        .Q(round_reg[165]) );
  DFF \round_reg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .I(g_init[166]), 
        .Q(round_reg[166]) );
  DFF \round_reg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .I(g_init[167]), 
        .Q(round_reg[167]) );
  DFF \round_reg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .I(g_init[168]), 
        .Q(round_reg[168]) );
  DFF \round_reg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .I(g_init[169]), 
        .Q(round_reg[169]) );
  DFF \round_reg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .I(g_init[170]), 
        .Q(round_reg[170]) );
  DFF \round_reg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .I(g_init[171]), 
        .Q(round_reg[171]) );
  DFF \round_reg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .I(g_init[172]), 
        .Q(round_reg[172]) );
  DFF \round_reg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .I(g_init[173]), 
        .Q(round_reg[173]) );
  DFF \round_reg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .I(g_init[174]), 
        .Q(round_reg[174]) );
  DFF \round_reg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .I(g_init[175]), 
        .Q(round_reg[175]) );
  DFF \round_reg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .I(g_init[176]), 
        .Q(round_reg[176]) );
  DFF \round_reg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .I(g_init[177]), 
        .Q(round_reg[177]) );
  DFF \round_reg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .I(g_init[178]), 
        .Q(round_reg[178]) );
  DFF \round_reg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .I(g_init[179]), 
        .Q(round_reg[179]) );
  DFF \round_reg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .I(g_init[180]), 
        .Q(round_reg[180]) );
  DFF \round_reg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .I(g_init[181]), 
        .Q(round_reg[181]) );
  DFF \round_reg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .I(g_init[182]), 
        .Q(round_reg[182]) );
  DFF \round_reg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .I(g_init[183]), 
        .Q(round_reg[183]) );
  DFF \round_reg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .I(g_init[184]), 
        .Q(round_reg[184]) );
  DFF \round_reg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .I(g_init[185]), 
        .Q(round_reg[185]) );
  DFF \round_reg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .I(g_init[186]), 
        .Q(round_reg[186]) );
  DFF \round_reg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .I(g_init[187]), 
        .Q(round_reg[187]) );
  DFF \round_reg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .I(g_init[188]), 
        .Q(round_reg[188]) );
  DFF \round_reg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .I(g_init[189]), 
        .Q(round_reg[189]) );
  DFF \round_reg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .I(g_init[190]), 
        .Q(round_reg[190]) );
  DFF \round_reg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .I(g_init[191]), 
        .Q(round_reg[191]) );
  DFF \round_reg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .I(g_init[192]), 
        .Q(round_reg[192]) );
  DFF \round_reg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .I(g_init[193]), 
        .Q(round_reg[193]) );
  DFF \round_reg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .I(g_init[194]), 
        .Q(round_reg[194]) );
  DFF \round_reg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .I(g_init[195]), 
        .Q(round_reg[195]) );
  DFF \round_reg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .I(g_init[196]), 
        .Q(round_reg[196]) );
  DFF \round_reg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .I(g_init[197]), 
        .Q(round_reg[197]) );
  DFF \round_reg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .I(g_init[198]), 
        .Q(round_reg[198]) );
  DFF \round_reg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .I(g_init[199]), 
        .Q(round_reg[199]) );
  DFF \round_reg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .I(g_init[200]), 
        .Q(round_reg[200]) );
  DFF \round_reg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .I(g_init[201]), 
        .Q(round_reg[201]) );
  DFF \round_reg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .I(g_init[202]), 
        .Q(round_reg[202]) );
  DFF \round_reg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .I(g_init[203]), 
        .Q(round_reg[203]) );
  DFF \round_reg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .I(g_init[204]), 
        .Q(round_reg[204]) );
  DFF \round_reg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .I(g_init[205]), 
        .Q(round_reg[205]) );
  DFF \round_reg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .I(g_init[206]), 
        .Q(round_reg[206]) );
  DFF \round_reg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .I(g_init[207]), 
        .Q(round_reg[207]) );
  DFF \round_reg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .I(g_init[208]), 
        .Q(round_reg[208]) );
  DFF \round_reg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .I(g_init[209]), 
        .Q(round_reg[209]) );
  DFF \round_reg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .I(g_init[210]), 
        .Q(round_reg[210]) );
  DFF \round_reg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .I(g_init[211]), 
        .Q(round_reg[211]) );
  DFF \round_reg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .I(g_init[212]), 
        .Q(round_reg[212]) );
  DFF \round_reg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .I(g_init[213]), 
        .Q(round_reg[213]) );
  DFF \round_reg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .I(g_init[214]), 
        .Q(round_reg[214]) );
  DFF \round_reg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .I(g_init[215]), 
        .Q(round_reg[215]) );
  DFF \round_reg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .I(g_init[216]), 
        .Q(round_reg[216]) );
  DFF \round_reg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .I(g_init[217]), 
        .Q(round_reg[217]) );
  DFF \round_reg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .I(g_init[218]), 
        .Q(round_reg[218]) );
  DFF \round_reg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .I(g_init[219]), 
        .Q(round_reg[219]) );
  DFF \round_reg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .I(g_init[220]), 
        .Q(round_reg[220]) );
  DFF \round_reg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .I(g_init[221]), 
        .Q(round_reg[221]) );
  DFF \round_reg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .I(g_init[222]), 
        .Q(round_reg[222]) );
  DFF \round_reg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .I(g_init[223]), 
        .Q(round_reg[223]) );
  DFF \round_reg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .I(g_init[224]), 
        .Q(round_reg[224]) );
  DFF \round_reg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .I(g_init[225]), 
        .Q(round_reg[225]) );
  DFF \round_reg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .I(g_init[226]), 
        .Q(round_reg[226]) );
  DFF \round_reg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .I(g_init[227]), 
        .Q(round_reg[227]) );
  DFF \round_reg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .I(g_init[228]), 
        .Q(round_reg[228]) );
  DFF \round_reg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .I(g_init[229]), 
        .Q(round_reg[229]) );
  DFF \round_reg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .I(g_init[230]), 
        .Q(round_reg[230]) );
  DFF \round_reg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .I(g_init[231]), 
        .Q(round_reg[231]) );
  DFF \round_reg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .I(g_init[232]), 
        .Q(round_reg[232]) );
  DFF \round_reg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .I(g_init[233]), 
        .Q(round_reg[233]) );
  DFF \round_reg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .I(g_init[234]), 
        .Q(round_reg[234]) );
  DFF \round_reg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .I(g_init[235]), 
        .Q(round_reg[235]) );
  DFF \round_reg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .I(g_init[236]), 
        .Q(round_reg[236]) );
  DFF \round_reg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .I(g_init[237]), 
        .Q(round_reg[237]) );
  DFF \round_reg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .I(g_init[238]), 
        .Q(round_reg[238]) );
  DFF \round_reg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .I(g_init[239]), 
        .Q(round_reg[239]) );
  DFF \round_reg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .I(g_init[240]), 
        .Q(round_reg[240]) );
  DFF \round_reg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .I(g_init[241]), 
        .Q(round_reg[241]) );
  DFF \round_reg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .I(g_init[242]), 
        .Q(round_reg[242]) );
  DFF \round_reg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .I(g_init[243]), 
        .Q(round_reg[243]) );
  DFF \round_reg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .I(g_init[244]), 
        .Q(round_reg[244]) );
  DFF \round_reg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .I(g_init[245]), 
        .Q(round_reg[245]) );
  DFF \round_reg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .I(g_init[246]), 
        .Q(round_reg[246]) );
  DFF \round_reg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .I(g_init[247]), 
        .Q(round_reg[247]) );
  DFF \round_reg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .I(g_init[248]), 
        .Q(round_reg[248]) );
  DFF \round_reg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .I(g_init[249]), 
        .Q(round_reg[249]) );
  DFF \round_reg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .I(g_init[250]), 
        .Q(round_reg[250]) );
  DFF \round_reg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .I(g_init[251]), 
        .Q(round_reg[251]) );
  DFF \round_reg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .I(g_init[252]), 
        .Q(round_reg[252]) );
  DFF \round_reg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .I(g_init[253]), 
        .Q(round_reg[253]) );
  DFF \round_reg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .I(g_init[254]), 
        .Q(round_reg[254]) );
  DFF \round_reg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .I(g_init[255]), 
        .Q(round_reg[255]) );
  DFF \round_reg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(rst), .I(g_init[256]), 
        .Q(round_reg[256]) );
  DFF \round_reg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(rst), .I(g_init[257]), 
        .Q(round_reg[257]) );
  DFF \round_reg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(rst), .I(g_init[258]), 
        .Q(round_reg[258]) );
  DFF \round_reg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(rst), .I(g_init[259]), 
        .Q(round_reg[259]) );
  DFF \round_reg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(rst), .I(g_init[260]), 
        .Q(round_reg[260]) );
  DFF \round_reg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(rst), .I(g_init[261]), 
        .Q(round_reg[261]) );
  DFF \round_reg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(rst), .I(g_init[262]), 
        .Q(round_reg[262]) );
  DFF \round_reg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(rst), .I(g_init[263]), 
        .Q(round_reg[263]) );
  DFF \round_reg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(rst), .I(g_init[264]), 
        .Q(round_reg[264]) );
  DFF \round_reg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(rst), .I(g_init[265]), 
        .Q(round_reg[265]) );
  DFF \round_reg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(rst), .I(g_init[266]), 
        .Q(round_reg[266]) );
  DFF \round_reg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(rst), .I(g_init[267]), 
        .Q(round_reg[267]) );
  DFF \round_reg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(rst), .I(g_init[268]), 
        .Q(round_reg[268]) );
  DFF \round_reg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(rst), .I(g_init[269]), 
        .Q(round_reg[269]) );
  DFF \round_reg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(rst), .I(g_init[270]), 
        .Q(round_reg[270]) );
  DFF \round_reg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(rst), .I(g_init[271]), 
        .Q(round_reg[271]) );
  DFF \round_reg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(rst), .I(g_init[272]), 
        .Q(round_reg[272]) );
  DFF \round_reg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(rst), .I(g_init[273]), 
        .Q(round_reg[273]) );
  DFF \round_reg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(rst), .I(g_init[274]), 
        .Q(round_reg[274]) );
  DFF \round_reg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(rst), .I(g_init[275]), 
        .Q(round_reg[275]) );
  DFF \round_reg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(rst), .I(g_init[276]), 
        .Q(round_reg[276]) );
  DFF \round_reg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(rst), .I(g_init[277]), 
        .Q(round_reg[277]) );
  DFF \round_reg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(rst), .I(g_init[278]), 
        .Q(round_reg[278]) );
  DFF \round_reg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(rst), .I(g_init[279]), 
        .Q(round_reg[279]) );
  DFF \round_reg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(rst), .I(g_init[280]), 
        .Q(round_reg[280]) );
  DFF \round_reg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(rst), .I(g_init[281]), 
        .Q(round_reg[281]) );
  DFF \round_reg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(rst), .I(g_init[282]), 
        .Q(round_reg[282]) );
  DFF \round_reg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(rst), .I(g_init[283]), 
        .Q(round_reg[283]) );
  DFF \round_reg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(rst), .I(g_init[284]), 
        .Q(round_reg[284]) );
  DFF \round_reg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(rst), .I(g_init[285]), 
        .Q(round_reg[285]) );
  DFF \round_reg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(rst), .I(g_init[286]), 
        .Q(round_reg[286]) );
  DFF \round_reg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(rst), .I(g_init[287]), 
        .Q(round_reg[287]) );
  DFF \round_reg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(rst), .I(e_init[0]), 
        .Q(round_reg[288]) );
  DFF \round_reg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(rst), .I(e_init[1]), 
        .Q(round_reg[289]) );
  DFF \round_reg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(rst), .I(e_init[2]), 
        .Q(round_reg[290]) );
  DFF \round_reg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(rst), .I(e_init[3]), 
        .Q(round_reg[291]) );
  DFF \round_reg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(rst), .I(e_init[4]), 
        .Q(round_reg[292]) );
  DFF \round_reg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(rst), .I(e_init[5]), 
        .Q(round_reg[293]) );
  DFF \round_reg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(rst), .I(e_init[6]), 
        .Q(round_reg[294]) );
  DFF \round_reg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(rst), .I(e_init[7]), 
        .Q(round_reg[295]) );
  DFF \round_reg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(rst), .I(e_init[8]), 
        .Q(round_reg[296]) );
  DFF \round_reg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(rst), .I(e_init[9]), 
        .Q(round_reg[297]) );
  DFF \round_reg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(rst), .I(e_init[10]), 
        .Q(round_reg[298]) );
  DFF \round_reg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(rst), .I(e_init[11]), 
        .Q(round_reg[299]) );
  DFF \round_reg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(rst), .I(e_init[12]), 
        .Q(round_reg[300]) );
  DFF \round_reg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(rst), .I(e_init[13]), 
        .Q(round_reg[301]) );
  DFF \round_reg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(rst), .I(e_init[14]), 
        .Q(round_reg[302]) );
  DFF \round_reg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(rst), .I(e_init[15]), 
        .Q(round_reg[303]) );
  DFF \round_reg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(rst), .I(e_init[16]), 
        .Q(round_reg[304]) );
  DFF \round_reg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(rst), .I(e_init[17]), 
        .Q(round_reg[305]) );
  DFF \round_reg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(rst), .I(e_init[18]), 
        .Q(round_reg[306]) );
  DFF \round_reg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(rst), .I(e_init[19]), 
        .Q(round_reg[307]) );
  DFF \round_reg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(rst), .I(e_init[20]), 
        .Q(round_reg[308]) );
  DFF \round_reg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(rst), .I(e_init[21]), 
        .Q(round_reg[309]) );
  DFF \round_reg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(rst), .I(e_init[22]), 
        .Q(round_reg[310]) );
  DFF \round_reg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(rst), .I(e_init[23]), 
        .Q(round_reg[311]) );
  DFF \round_reg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(rst), .I(e_init[24]), 
        .Q(round_reg[312]) );
  DFF \round_reg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(rst), .I(e_init[25]), 
        .Q(round_reg[313]) );
  DFF \round_reg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(rst), .I(e_init[26]), 
        .Q(round_reg[314]) );
  DFF \round_reg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(rst), .I(e_init[27]), 
        .Q(round_reg[315]) );
  DFF \round_reg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(rst), .I(e_init[28]), 
        .Q(round_reg[316]) );
  DFF \round_reg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(rst), .I(e_init[29]), 
        .Q(round_reg[317]) );
  DFF \round_reg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(rst), .I(e_init[30]), 
        .Q(round_reg[318]) );
  DFF \round_reg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(rst), .I(e_init[31]), 
        .Q(round_reg[319]) );
  DFF \round_reg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(rst), .I(e_init[32]), 
        .Q(round_reg[320]) );
  DFF \round_reg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(rst), .I(e_init[33]), 
        .Q(round_reg[321]) );
  DFF \round_reg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(rst), .I(e_init[34]), 
        .Q(round_reg[322]) );
  DFF \round_reg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(rst), .I(e_init[35]), 
        .Q(round_reg[323]) );
  DFF \round_reg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(rst), .I(e_init[36]), 
        .Q(round_reg[324]) );
  DFF \round_reg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(rst), .I(e_init[37]), 
        .Q(round_reg[325]) );
  DFF \round_reg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(rst), .I(e_init[38]), 
        .Q(round_reg[326]) );
  DFF \round_reg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(rst), .I(e_init[39]), 
        .Q(round_reg[327]) );
  DFF \round_reg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(rst), .I(e_init[40]), 
        .Q(round_reg[328]) );
  DFF \round_reg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(rst), .I(e_init[41]), 
        .Q(round_reg[329]) );
  DFF \round_reg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(rst), .I(e_init[42]), 
        .Q(round_reg[330]) );
  DFF \round_reg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(rst), .I(e_init[43]), 
        .Q(round_reg[331]) );
  DFF \round_reg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(rst), .I(e_init[44]), 
        .Q(round_reg[332]) );
  DFF \round_reg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(rst), .I(e_init[45]), 
        .Q(round_reg[333]) );
  DFF \round_reg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(rst), .I(e_init[46]), 
        .Q(round_reg[334]) );
  DFF \round_reg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(rst), .I(e_init[47]), 
        .Q(round_reg[335]) );
  DFF \round_reg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(rst), .I(e_init[48]), 
        .Q(round_reg[336]) );
  DFF \round_reg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(rst), .I(e_init[49]), 
        .Q(round_reg[337]) );
  DFF \round_reg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(rst), .I(e_init[50]), 
        .Q(round_reg[338]) );
  DFF \round_reg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(rst), .I(e_init[51]), 
        .Q(round_reg[339]) );
  DFF \round_reg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(rst), .I(e_init[52]), 
        .Q(round_reg[340]) );
  DFF \round_reg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(rst), .I(e_init[53]), 
        .Q(round_reg[341]) );
  DFF \round_reg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(rst), .I(e_init[54]), 
        .Q(round_reg[342]) );
  DFF \round_reg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(rst), .I(e_init[55]), 
        .Q(round_reg[343]) );
  DFF \round_reg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(rst), .I(e_init[56]), 
        .Q(round_reg[344]) );
  DFF \round_reg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(rst), .I(e_init[57]), 
        .Q(round_reg[345]) );
  DFF \round_reg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(rst), .I(e_init[58]), 
        .Q(round_reg[346]) );
  DFF \round_reg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(rst), .I(e_init[59]), 
        .Q(round_reg[347]) );
  DFF \round_reg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(rst), .I(e_init[60]), 
        .Q(round_reg[348]) );
  DFF \round_reg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(rst), .I(e_init[61]), 
        .Q(round_reg[349]) );
  DFF \round_reg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(rst), .I(e_init[62]), 
        .Q(round_reg[350]) );
  DFF \round_reg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(rst), .I(e_init[63]), 
        .Q(round_reg[351]) );
  DFF \round_reg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(rst), .I(e_init[64]), 
        .Q(round_reg[352]) );
  DFF \round_reg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(rst), .I(e_init[65]), 
        .Q(round_reg[353]) );
  DFF \round_reg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(rst), .I(e_init[66]), 
        .Q(round_reg[354]) );
  DFF \round_reg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(rst), .I(e_init[67]), 
        .Q(round_reg[355]) );
  DFF \round_reg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(rst), .I(e_init[68]), 
        .Q(round_reg[356]) );
  DFF \round_reg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(rst), .I(e_init[69]), 
        .Q(round_reg[357]) );
  DFF \round_reg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(rst), .I(e_init[70]), 
        .Q(round_reg[358]) );
  DFF \round_reg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(rst), .I(e_init[71]), 
        .Q(round_reg[359]) );
  DFF \round_reg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(rst), .I(e_init[72]), 
        .Q(round_reg[360]) );
  DFF \round_reg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(rst), .I(e_init[73]), 
        .Q(round_reg[361]) );
  DFF \round_reg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(rst), .I(e_init[74]), 
        .Q(round_reg[362]) );
  DFF \round_reg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(rst), .I(e_init[75]), 
        .Q(round_reg[363]) );
  DFF \round_reg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(rst), .I(e_init[76]), 
        .Q(round_reg[364]) );
  DFF \round_reg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(rst), .I(e_init[77]), 
        .Q(round_reg[365]) );
  DFF \round_reg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(rst), .I(e_init[78]), 
        .Q(round_reg[366]) );
  DFF \round_reg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(rst), .I(e_init[79]), 
        .Q(round_reg[367]) );
  DFF \round_reg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(rst), .I(e_init[80]), 
        .Q(round_reg[368]) );
  DFF \round_reg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(rst), .I(e_init[81]), 
        .Q(round_reg[369]) );
  DFF \round_reg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(rst), .I(e_init[82]), 
        .Q(round_reg[370]) );
  DFF \round_reg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(rst), .I(e_init[83]), 
        .Q(round_reg[371]) );
  DFF \round_reg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(rst), .I(e_init[84]), 
        .Q(round_reg[372]) );
  DFF \round_reg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(rst), .I(e_init[85]), 
        .Q(round_reg[373]) );
  DFF \round_reg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(rst), .I(e_init[86]), 
        .Q(round_reg[374]) );
  DFF \round_reg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(rst), .I(e_init[87]), 
        .Q(round_reg[375]) );
  DFF \round_reg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(rst), .I(e_init[88]), 
        .Q(round_reg[376]) );
  DFF \round_reg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(rst), .I(e_init[89]), 
        .Q(round_reg[377]) );
  DFF \round_reg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(rst), .I(e_init[90]), 
        .Q(round_reg[378]) );
  DFF \round_reg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(rst), .I(e_init[91]), 
        .Q(round_reg[379]) );
  DFF \round_reg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(rst), .I(e_init[92]), 
        .Q(round_reg[380]) );
  DFF \round_reg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(rst), .I(e_init[93]), 
        .Q(round_reg[381]) );
  DFF \round_reg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(rst), .I(e_init[94]), 
        .Q(round_reg[382]) );
  DFF \round_reg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(rst), .I(e_init[95]), 
        .Q(round_reg[383]) );
  DFF \round_reg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(rst), .I(e_init[96]), 
        .Q(round_reg[384]) );
  DFF \round_reg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(rst), .I(e_init[97]), 
        .Q(round_reg[385]) );
  DFF \round_reg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(rst), .I(e_init[98]), 
        .Q(round_reg[386]) );
  DFF \round_reg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(rst), .I(e_init[99]), 
        .Q(round_reg[387]) );
  DFF \round_reg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(rst), .I(e_init[100]), 
        .Q(round_reg[388]) );
  DFF \round_reg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(rst), .I(e_init[101]), 
        .Q(round_reg[389]) );
  DFF \round_reg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(rst), .I(e_init[102]), 
        .Q(round_reg[390]) );
  DFF \round_reg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(rst), .I(e_init[103]), 
        .Q(round_reg[391]) );
  DFF \round_reg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(rst), .I(e_init[104]), 
        .Q(round_reg[392]) );
  DFF \round_reg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(rst), .I(e_init[105]), 
        .Q(round_reg[393]) );
  DFF \round_reg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(rst), .I(e_init[106]), 
        .Q(round_reg[394]) );
  DFF \round_reg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(rst), .I(e_init[107]), 
        .Q(round_reg[395]) );
  DFF \round_reg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(rst), .I(e_init[108]), 
        .Q(round_reg[396]) );
  DFF \round_reg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(rst), .I(e_init[109]), 
        .Q(round_reg[397]) );
  DFF \round_reg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(rst), .I(e_init[110]), 
        .Q(round_reg[398]) );
  DFF \round_reg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(rst), .I(e_init[111]), 
        .Q(round_reg[399]) );
  DFF \round_reg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(rst), .I(e_init[112]), 
        .Q(round_reg[400]) );
  DFF \round_reg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(rst), .I(e_init[113]), 
        .Q(round_reg[401]) );
  DFF \round_reg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(rst), .I(e_init[114]), 
        .Q(round_reg[402]) );
  DFF \round_reg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(rst), .I(e_init[115]), 
        .Q(round_reg[403]) );
  DFF \round_reg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(rst), .I(e_init[116]), 
        .Q(round_reg[404]) );
  DFF \round_reg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(rst), .I(e_init[117]), 
        .Q(round_reg[405]) );
  DFF \round_reg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(rst), .I(e_init[118]), 
        .Q(round_reg[406]) );
  DFF \round_reg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(rst), .I(e_init[119]), 
        .Q(round_reg[407]) );
  DFF \round_reg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(rst), .I(e_init[120]), 
        .Q(round_reg[408]) );
  DFF \round_reg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(rst), .I(e_init[121]), 
        .Q(round_reg[409]) );
  DFF \round_reg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(rst), .I(e_init[122]), 
        .Q(round_reg[410]) );
  DFF \round_reg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(rst), .I(e_init[123]), 
        .Q(round_reg[411]) );
  DFF \round_reg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(rst), .I(e_init[124]), 
        .Q(round_reg[412]) );
  DFF \round_reg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(rst), .I(e_init[125]), 
        .Q(round_reg[413]) );
  DFF \round_reg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(rst), .I(e_init[126]), 
        .Q(round_reg[414]) );
  DFF \round_reg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(rst), .I(e_init[127]), 
        .Q(round_reg[415]) );
  DFF \round_reg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(rst), .I(e_init[128]), 
        .Q(round_reg[416]) );
  DFF \round_reg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(rst), .I(e_init[129]), 
        .Q(round_reg[417]) );
  DFF \round_reg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(rst), .I(e_init[130]), 
        .Q(round_reg[418]) );
  DFF \round_reg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(rst), .I(e_init[131]), 
        .Q(round_reg[419]) );
  DFF \round_reg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(rst), .I(e_init[132]), 
        .Q(round_reg[420]) );
  DFF \round_reg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(rst), .I(e_init[133]), 
        .Q(round_reg[421]) );
  DFF \round_reg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(rst), .I(e_init[134]), 
        .Q(round_reg[422]) );
  DFF \round_reg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(rst), .I(e_init[135]), 
        .Q(round_reg[423]) );
  DFF \round_reg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(rst), .I(e_init[136]), 
        .Q(round_reg[424]) );
  DFF \round_reg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(rst), .I(e_init[137]), 
        .Q(round_reg[425]) );
  DFF \round_reg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(rst), .I(e_init[138]), 
        .Q(round_reg[426]) );
  DFF \round_reg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(rst), .I(e_init[139]), 
        .Q(round_reg[427]) );
  DFF \round_reg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(rst), .I(e_init[140]), 
        .Q(round_reg[428]) );
  DFF \round_reg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(rst), .I(e_init[141]), 
        .Q(round_reg[429]) );
  DFF \round_reg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(rst), .I(e_init[142]), 
        .Q(round_reg[430]) );
  DFF \round_reg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(rst), .I(e_init[143]), 
        .Q(round_reg[431]) );
  DFF \round_reg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(rst), .I(e_init[144]), 
        .Q(round_reg[432]) );
  DFF \round_reg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(rst), .I(e_init[145]), 
        .Q(round_reg[433]) );
  DFF \round_reg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(rst), .I(e_init[146]), 
        .Q(round_reg[434]) );
  DFF \round_reg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(rst), .I(e_init[147]), 
        .Q(round_reg[435]) );
  DFF \round_reg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(rst), .I(e_init[148]), 
        .Q(round_reg[436]) );
  DFF \round_reg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(rst), .I(e_init[149]), 
        .Q(round_reg[437]) );
  DFF \round_reg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(rst), .I(e_init[150]), 
        .Q(round_reg[438]) );
  DFF \round_reg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(rst), .I(e_init[151]), 
        .Q(round_reg[439]) );
  DFF \round_reg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(rst), .I(e_init[152]), 
        .Q(round_reg[440]) );
  DFF \round_reg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(rst), .I(e_init[153]), 
        .Q(round_reg[441]) );
  DFF \round_reg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(rst), .I(e_init[154]), 
        .Q(round_reg[442]) );
  DFF \round_reg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(rst), .I(e_init[155]), 
        .Q(round_reg[443]) );
  DFF \round_reg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(rst), .I(e_init[156]), 
        .Q(round_reg[444]) );
  DFF \round_reg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(rst), .I(e_init[157]), 
        .Q(round_reg[445]) );
  DFF \round_reg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(rst), .I(e_init[158]), 
        .Q(round_reg[446]) );
  DFF \round_reg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(rst), .I(e_init[159]), 
        .Q(round_reg[447]) );
  DFF \round_reg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(rst), .I(e_init[160]), 
        .Q(round_reg[448]) );
  DFF \round_reg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(rst), .I(e_init[161]), 
        .Q(round_reg[449]) );
  DFF \round_reg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(rst), .I(e_init[162]), 
        .Q(round_reg[450]) );
  DFF \round_reg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(rst), .I(e_init[163]), 
        .Q(round_reg[451]) );
  DFF \round_reg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(rst), .I(e_init[164]), 
        .Q(round_reg[452]) );
  DFF \round_reg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(rst), .I(e_init[165]), 
        .Q(round_reg[453]) );
  DFF \round_reg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(rst), .I(e_init[166]), 
        .Q(round_reg[454]) );
  DFF \round_reg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(rst), .I(e_init[167]), 
        .Q(round_reg[455]) );
  DFF \round_reg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(rst), .I(e_init[168]), 
        .Q(round_reg[456]) );
  DFF \round_reg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(rst), .I(e_init[169]), 
        .Q(round_reg[457]) );
  DFF \round_reg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(rst), .I(e_init[170]), 
        .Q(round_reg[458]) );
  DFF \round_reg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(rst), .I(e_init[171]), 
        .Q(round_reg[459]) );
  DFF \round_reg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(rst), .I(e_init[172]), 
        .Q(round_reg[460]) );
  DFF \round_reg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(rst), .I(e_init[173]), 
        .Q(round_reg[461]) );
  DFF \round_reg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(rst), .I(e_init[174]), 
        .Q(round_reg[462]) );
  DFF \round_reg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(rst), .I(e_init[175]), 
        .Q(round_reg[463]) );
  DFF \round_reg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(rst), .I(e_init[176]), 
        .Q(round_reg[464]) );
  DFF \round_reg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(rst), .I(e_init[177]), 
        .Q(round_reg[465]) );
  DFF \round_reg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(rst), .I(e_init[178]), 
        .Q(round_reg[466]) );
  DFF \round_reg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(rst), .I(e_init[179]), 
        .Q(round_reg[467]) );
  DFF \round_reg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(rst), .I(e_init[180]), 
        .Q(round_reg[468]) );
  DFF \round_reg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(rst), .I(e_init[181]), 
        .Q(round_reg[469]) );
  DFF \round_reg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(rst), .I(e_init[182]), 
        .Q(round_reg[470]) );
  DFF \round_reg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(rst), .I(e_init[183]), 
        .Q(round_reg[471]) );
  DFF \round_reg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(rst), .I(e_init[184]), 
        .Q(round_reg[472]) );
  DFF \round_reg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(rst), .I(e_init[185]), 
        .Q(round_reg[473]) );
  DFF \round_reg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(rst), .I(e_init[186]), 
        .Q(round_reg[474]) );
  DFF \round_reg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(rst), .I(e_init[187]), 
        .Q(round_reg[475]) );
  DFF \round_reg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(rst), .I(e_init[188]), 
        .Q(round_reg[476]) );
  DFF \round_reg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(rst), .I(e_init[189]), 
        .Q(round_reg[477]) );
  DFF \round_reg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(rst), .I(e_init[190]), 
        .Q(round_reg[478]) );
  DFF \round_reg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(rst), .I(e_init[191]), 
        .Q(round_reg[479]) );
  DFF \round_reg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(rst), .I(e_init[192]), 
        .Q(round_reg[480]) );
  DFF \round_reg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(rst), .I(e_init[193]), 
        .Q(round_reg[481]) );
  DFF \round_reg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(rst), .I(e_init[194]), 
        .Q(round_reg[482]) );
  DFF \round_reg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(rst), .I(e_init[195]), 
        .Q(round_reg[483]) );
  DFF \round_reg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(rst), .I(e_init[196]), 
        .Q(round_reg[484]) );
  DFF \round_reg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(rst), .I(e_init[197]), 
        .Q(round_reg[485]) );
  DFF \round_reg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(rst), .I(e_init[198]), 
        .Q(round_reg[486]) );
  DFF \round_reg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(rst), .I(e_init[199]), 
        .Q(round_reg[487]) );
  DFF \round_reg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(rst), .I(e_init[200]), 
        .Q(round_reg[488]) );
  DFF \round_reg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(rst), .I(e_init[201]), 
        .Q(round_reg[489]) );
  DFF \round_reg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(rst), .I(e_init[202]), 
        .Q(round_reg[490]) );
  DFF \round_reg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(rst), .I(e_init[203]), 
        .Q(round_reg[491]) );
  DFF \round_reg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(rst), .I(e_init[204]), 
        .Q(round_reg[492]) );
  DFF \round_reg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(rst), .I(e_init[205]), 
        .Q(round_reg[493]) );
  DFF \round_reg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(rst), .I(e_init[206]), 
        .Q(round_reg[494]) );
  DFF \round_reg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(rst), .I(e_init[207]), 
        .Q(round_reg[495]) );
  DFF \round_reg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(rst), .I(e_init[208]), 
        .Q(round_reg[496]) );
  DFF \round_reg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(rst), .I(e_init[209]), 
        .Q(round_reg[497]) );
  DFF \round_reg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(rst), .I(e_init[210]), 
        .Q(round_reg[498]) );
  DFF \round_reg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(rst), .I(e_init[211]), 
        .Q(round_reg[499]) );
  DFF \round_reg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(rst), .I(e_init[212]), 
        .Q(round_reg[500]) );
  DFF \round_reg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(rst), .I(e_init[213]), 
        .Q(round_reg[501]) );
  DFF \round_reg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(rst), .I(e_init[214]), 
        .Q(round_reg[502]) );
  DFF \round_reg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(rst), .I(e_init[215]), 
        .Q(round_reg[503]) );
  DFF \round_reg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(rst), .I(e_init[216]), 
        .Q(round_reg[504]) );
  DFF \round_reg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(rst), .I(e_init[217]), 
        .Q(round_reg[505]) );
  DFF \round_reg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(rst), .I(e_init[218]), 
        .Q(round_reg[506]) );
  DFF \round_reg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(rst), .I(e_init[219]), 
        .Q(round_reg[507]) );
  DFF \round_reg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(rst), .I(e_init[220]), 
        .Q(round_reg[508]) );
  DFF \round_reg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(rst), .I(e_init[221]), 
        .Q(round_reg[509]) );
  DFF \round_reg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(rst), .I(e_init[222]), 
        .Q(round_reg[510]) );
  DFF \round_reg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(rst), .I(e_init[223]), 
        .Q(round_reg[511]) );
  DFF \round_reg_reg[512]  ( .D(o[512]), .CLK(clk), .RST(rst), .I(e_init[224]), 
        .Q(round_reg[512]) );
  DFF \round_reg_reg[513]  ( .D(o[513]), .CLK(clk), .RST(rst), .I(e_init[225]), 
        .Q(round_reg[513]) );
  DFF \round_reg_reg[514]  ( .D(o[514]), .CLK(clk), .RST(rst), .I(e_init[226]), 
        .Q(round_reg[514]) );
  DFF \round_reg_reg[515]  ( .D(o[515]), .CLK(clk), .RST(rst), .I(e_init[227]), 
        .Q(round_reg[515]) );
  DFF \round_reg_reg[516]  ( .D(o[516]), .CLK(clk), .RST(rst), .I(e_init[228]), 
        .Q(round_reg[516]) );
  DFF \round_reg_reg[517]  ( .D(o[517]), .CLK(clk), .RST(rst), .I(e_init[229]), 
        .Q(round_reg[517]) );
  DFF \round_reg_reg[518]  ( .D(o[518]), .CLK(clk), .RST(rst), .I(e_init[230]), 
        .Q(round_reg[518]) );
  DFF \round_reg_reg[519]  ( .D(o[519]), .CLK(clk), .RST(rst), .I(e_init[231]), 
        .Q(round_reg[519]) );
  DFF \round_reg_reg[520]  ( .D(o[520]), .CLK(clk), .RST(rst), .I(e_init[232]), 
        .Q(round_reg[520]) );
  DFF \round_reg_reg[521]  ( .D(o[521]), .CLK(clk), .RST(rst), .I(e_init[233]), 
        .Q(round_reg[521]) );
  DFF \round_reg_reg[522]  ( .D(o[522]), .CLK(clk), .RST(rst), .I(e_init[234]), 
        .Q(round_reg[522]) );
  DFF \round_reg_reg[523]  ( .D(o[523]), .CLK(clk), .RST(rst), .I(e_init[235]), 
        .Q(round_reg[523]) );
  DFF \round_reg_reg[524]  ( .D(o[524]), .CLK(clk), .RST(rst), .I(e_init[236]), 
        .Q(round_reg[524]) );
  DFF \round_reg_reg[525]  ( .D(o[525]), .CLK(clk), .RST(rst), .I(e_init[237]), 
        .Q(round_reg[525]) );
  DFF \round_reg_reg[526]  ( .D(o[526]), .CLK(clk), .RST(rst), .I(e_init[238]), 
        .Q(round_reg[526]) );
  DFF \round_reg_reg[527]  ( .D(o[527]), .CLK(clk), .RST(rst), .I(e_init[239]), 
        .Q(round_reg[527]) );
  DFF \round_reg_reg[528]  ( .D(o[528]), .CLK(clk), .RST(rst), .I(e_init[240]), 
        .Q(round_reg[528]) );
  DFF \round_reg_reg[529]  ( .D(o[529]), .CLK(clk), .RST(rst), .I(e_init[241]), 
        .Q(round_reg[529]) );
  DFF \round_reg_reg[530]  ( .D(o[530]), .CLK(clk), .RST(rst), .I(e_init[242]), 
        .Q(round_reg[530]) );
  DFF \round_reg_reg[531]  ( .D(o[531]), .CLK(clk), .RST(rst), .I(e_init[243]), 
        .Q(round_reg[531]) );
  DFF \round_reg_reg[532]  ( .D(o[532]), .CLK(clk), .RST(rst), .I(e_init[244]), 
        .Q(round_reg[532]) );
  DFF \round_reg_reg[533]  ( .D(o[533]), .CLK(clk), .RST(rst), .I(e_init[245]), 
        .Q(round_reg[533]) );
  DFF \round_reg_reg[534]  ( .D(o[534]), .CLK(clk), .RST(rst), .I(e_init[246]), 
        .Q(round_reg[534]) );
  DFF \round_reg_reg[535]  ( .D(o[535]), .CLK(clk), .RST(rst), .I(e_init[247]), 
        .Q(round_reg[535]) );
  DFF \round_reg_reg[536]  ( .D(o[536]), .CLK(clk), .RST(rst), .I(e_init[248]), 
        .Q(round_reg[536]) );
  DFF \round_reg_reg[537]  ( .D(o[537]), .CLK(clk), .RST(rst), .I(e_init[249]), 
        .Q(round_reg[537]) );
  DFF \round_reg_reg[538]  ( .D(o[538]), .CLK(clk), .RST(rst), .I(e_init[250]), 
        .Q(round_reg[538]) );
  DFF \round_reg_reg[539]  ( .D(o[539]), .CLK(clk), .RST(rst), .I(e_init[251]), 
        .Q(round_reg[539]) );
  DFF \round_reg_reg[540]  ( .D(o[540]), .CLK(clk), .RST(rst), .I(e_init[252]), 
        .Q(round_reg[540]) );
  DFF \round_reg_reg[541]  ( .D(o[541]), .CLK(clk), .RST(rst), .I(e_init[253]), 
        .Q(round_reg[541]) );
  DFF \round_reg_reg[542]  ( .D(o[542]), .CLK(clk), .RST(rst), .I(e_init[254]), 
        .Q(round_reg[542]) );
  DFF \round_reg_reg[543]  ( .D(o[543]), .CLK(clk), .RST(rst), .I(e_init[255]), 
        .Q(round_reg[543]) );
  DFF \round_reg_reg[544]  ( .D(o[544]), .CLK(clk), .RST(rst), .I(e_init[256]), 
        .Q(round_reg[544]) );
  DFF \round_reg_reg[545]  ( .D(o[545]), .CLK(clk), .RST(rst), .I(e_init[257]), 
        .Q(round_reg[545]) );
  DFF \round_reg_reg[546]  ( .D(o[546]), .CLK(clk), .RST(rst), .I(e_init[258]), 
        .Q(round_reg[546]) );
  DFF \round_reg_reg[547]  ( .D(o[547]), .CLK(clk), .RST(rst), .I(e_init[259]), 
        .Q(round_reg[547]) );
  DFF \round_reg_reg[548]  ( .D(o[548]), .CLK(clk), .RST(rst), .I(e_init[260]), 
        .Q(round_reg[548]) );
  DFF \round_reg_reg[549]  ( .D(o[549]), .CLK(clk), .RST(rst), .I(e_init[261]), 
        .Q(round_reg[549]) );
  DFF \round_reg_reg[550]  ( .D(o[550]), .CLK(clk), .RST(rst), .I(e_init[262]), 
        .Q(round_reg[550]) );
  DFF \round_reg_reg[551]  ( .D(o[551]), .CLK(clk), .RST(rst), .I(e_init[263]), 
        .Q(round_reg[551]) );
  DFF \round_reg_reg[552]  ( .D(o[552]), .CLK(clk), .RST(rst), .I(e_init[264]), 
        .Q(round_reg[552]) );
  DFF \round_reg_reg[553]  ( .D(o[553]), .CLK(clk), .RST(rst), .I(e_init[265]), 
        .Q(round_reg[553]) );
  DFF \round_reg_reg[554]  ( .D(o[554]), .CLK(clk), .RST(rst), .I(e_init[266]), 
        .Q(round_reg[554]) );
  DFF \round_reg_reg[555]  ( .D(o[555]), .CLK(clk), .RST(rst), .I(e_init[267]), 
        .Q(round_reg[555]) );
  DFF \round_reg_reg[556]  ( .D(o[556]), .CLK(clk), .RST(rst), .I(e_init[268]), 
        .Q(round_reg[556]) );
  DFF \round_reg_reg[557]  ( .D(o[557]), .CLK(clk), .RST(rst), .I(e_init[269]), 
        .Q(round_reg[557]) );
  DFF \round_reg_reg[558]  ( .D(o[558]), .CLK(clk), .RST(rst), .I(e_init[270]), 
        .Q(round_reg[558]) );
  DFF \round_reg_reg[559]  ( .D(o[559]), .CLK(clk), .RST(rst), .I(e_init[271]), 
        .Q(round_reg[559]) );
  DFF \round_reg_reg[560]  ( .D(o[560]), .CLK(clk), .RST(rst), .I(e_init[272]), 
        .Q(round_reg[560]) );
  DFF \round_reg_reg[561]  ( .D(o[561]), .CLK(clk), .RST(rst), .I(e_init[273]), 
        .Q(round_reg[561]) );
  DFF \round_reg_reg[562]  ( .D(o[562]), .CLK(clk), .RST(rst), .I(e_init[274]), 
        .Q(round_reg[562]) );
  DFF \round_reg_reg[563]  ( .D(o[563]), .CLK(clk), .RST(rst), .I(e_init[275]), 
        .Q(round_reg[563]) );
  DFF \round_reg_reg[564]  ( .D(o[564]), .CLK(clk), .RST(rst), .I(e_init[276]), 
        .Q(round_reg[564]) );
  DFF \round_reg_reg[565]  ( .D(o[565]), .CLK(clk), .RST(rst), .I(e_init[277]), 
        .Q(round_reg[565]) );
  DFF \round_reg_reg[566]  ( .D(o[566]), .CLK(clk), .RST(rst), .I(e_init[278]), 
        .Q(round_reg[566]) );
  DFF \round_reg_reg[567]  ( .D(o[567]), .CLK(clk), .RST(rst), .I(e_init[279]), 
        .Q(round_reg[567]) );
  DFF \round_reg_reg[568]  ( .D(o[568]), .CLK(clk), .RST(rst), .I(e_init[280]), 
        .Q(round_reg[568]) );
  DFF \round_reg_reg[569]  ( .D(o[569]), .CLK(clk), .RST(rst), .I(e_init[281]), 
        .Q(round_reg[569]) );
  DFF \round_reg_reg[570]  ( .D(o[570]), .CLK(clk), .RST(rst), .I(e_init[282]), 
        .Q(round_reg[570]) );
  DFF \round_reg_reg[571]  ( .D(o[571]), .CLK(clk), .RST(rst), .I(e_init[283]), 
        .Q(round_reg[571]) );
  DFF \round_reg_reg[572]  ( .D(o[572]), .CLK(clk), .RST(rst), .I(e_init[284]), 
        .Q(round_reg[572]) );
  DFF \round_reg_reg[573]  ( .D(o[573]), .CLK(clk), .RST(rst), .I(e_init[285]), 
        .Q(round_reg[573]) );
  DFF \round_reg_reg[574]  ( .D(o[574]), .CLK(clk), .RST(rst), .I(e_init[286]), 
        .Q(round_reg[574]) );
  DFF \round_reg_reg[575]  ( .D(o[575]), .CLK(clk), .RST(rst), .I(e_init[287]), 
        .Q(round_reg[575]) );
  DFF \round_reg_reg[576]  ( .D(o[576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[576]) );
  DFF \round_reg_reg[577]  ( .D(o[577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[577]) );
  DFF \round_reg_reg[578]  ( .D(o[578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[578]) );
  DFF \round_reg_reg[579]  ( .D(o[579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[579]) );
  DFF \round_reg_reg[580]  ( .D(o[580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[580]) );
  DFF \round_reg_reg[581]  ( .D(o[581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[581]) );
  DFF \round_reg_reg[582]  ( .D(o[582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[582]) );
  DFF \round_reg_reg[583]  ( .D(o[583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[583]) );
  DFF \round_reg_reg[584]  ( .D(o[584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[584]) );
  DFF \round_reg_reg[585]  ( .D(o[585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[585]) );
  DFF \round_reg_reg[586]  ( .D(o[586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[586]) );
  DFF \round_reg_reg[587]  ( .D(o[587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[587]) );
  DFF \round_reg_reg[588]  ( .D(o[588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[588]) );
  DFF \round_reg_reg[589]  ( .D(o[589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[589]) );
  DFF \round_reg_reg[590]  ( .D(o[590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[590]) );
  DFF \round_reg_reg[591]  ( .D(o[591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[591]) );
  DFF \round_reg_reg[592]  ( .D(o[592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[592]) );
  DFF \round_reg_reg[593]  ( .D(o[593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[593]) );
  DFF \round_reg_reg[594]  ( .D(o[594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[594]) );
  DFF \round_reg_reg[595]  ( .D(o[595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[595]) );
  DFF \round_reg_reg[596]  ( .D(o[596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[596]) );
  DFF \round_reg_reg[597]  ( .D(o[597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[597]) );
  DFF \round_reg_reg[598]  ( .D(o[598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[598]) );
  DFF \round_reg_reg[599]  ( .D(o[599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[599]) );
  DFF \round_reg_reg[600]  ( .D(o[600]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[600]) );
  DFF \round_reg_reg[601]  ( .D(o[601]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[601]) );
  DFF \round_reg_reg[602]  ( .D(o[602]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[602]) );
  DFF \round_reg_reg[603]  ( .D(o[603]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[603]) );
  DFF \round_reg_reg[604]  ( .D(o[604]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[604]) );
  DFF \round_reg_reg[605]  ( .D(o[605]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[605]) );
  DFF \round_reg_reg[606]  ( .D(o[606]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[606]) );
  DFF \round_reg_reg[607]  ( .D(o[607]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[607]) );
  DFF \round_reg_reg[608]  ( .D(o[608]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[608]) );
  DFF \round_reg_reg[609]  ( .D(o[609]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[609]) );
  DFF \round_reg_reg[610]  ( .D(o[610]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[610]) );
  DFF \round_reg_reg[611]  ( .D(o[611]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[611]) );
  DFF \round_reg_reg[612]  ( .D(o[612]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[612]) );
  DFF \round_reg_reg[613]  ( .D(o[613]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[613]) );
  DFF \round_reg_reg[614]  ( .D(o[614]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[614]) );
  DFF \round_reg_reg[615]  ( .D(o[615]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[615]) );
  DFF \round_reg_reg[616]  ( .D(o[616]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[616]) );
  DFF \round_reg_reg[617]  ( .D(o[617]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[617]) );
  DFF \round_reg_reg[618]  ( .D(o[618]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[618]) );
  DFF \round_reg_reg[619]  ( .D(o[619]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[619]) );
  DFF \round_reg_reg[620]  ( .D(o[620]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[620]) );
  DFF \round_reg_reg[621]  ( .D(o[621]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[621]) );
  DFF \round_reg_reg[622]  ( .D(o[622]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[622]) );
  DFF \round_reg_reg[623]  ( .D(o[623]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[623]) );
  DFF \round_reg_reg[624]  ( .D(o[624]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[624]) );
  DFF \round_reg_reg[625]  ( .D(o[625]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[625]) );
  DFF \round_reg_reg[626]  ( .D(o[626]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[626]) );
  DFF \round_reg_reg[627]  ( .D(o[627]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[627]) );
  DFF \round_reg_reg[628]  ( .D(o[628]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[628]) );
  DFF \round_reg_reg[629]  ( .D(o[629]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[629]) );
  DFF \round_reg_reg[630]  ( .D(o[630]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[630]) );
  DFF \round_reg_reg[631]  ( .D(o[631]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[631]) );
  DFF \round_reg_reg[632]  ( .D(o[632]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[632]) );
  DFF \round_reg_reg[633]  ( .D(o[633]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[633]) );
  DFF \round_reg_reg[634]  ( .D(o[634]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[634]) );
  DFF \round_reg_reg[635]  ( .D(o[635]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[635]) );
  DFF \round_reg_reg[636]  ( .D(o[636]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[636]) );
  DFF \round_reg_reg[637]  ( .D(o[637]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[637]) );
  DFF \round_reg_reg[638]  ( .D(o[638]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[638]) );
  DFF \round_reg_reg[639]  ( .D(o[639]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[639]) );
  DFF \round_reg_reg[640]  ( .D(o[640]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[640]) );
  DFF \round_reg_reg[641]  ( .D(o[641]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[641]) );
  DFF \round_reg_reg[642]  ( .D(o[642]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[642]) );
  DFF \round_reg_reg[643]  ( .D(o[643]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[643]) );
  DFF \round_reg_reg[644]  ( .D(o[644]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[644]) );
  DFF \round_reg_reg[645]  ( .D(o[645]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[645]) );
  DFF \round_reg_reg[646]  ( .D(o[646]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[646]) );
  DFF \round_reg_reg[647]  ( .D(o[647]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[647]) );
  DFF \round_reg_reg[648]  ( .D(o[648]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[648]) );
  DFF \round_reg_reg[649]  ( .D(o[649]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[649]) );
  DFF \round_reg_reg[650]  ( .D(o[650]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[650]) );
  DFF \round_reg_reg[651]  ( .D(o[651]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[651]) );
  DFF \round_reg_reg[652]  ( .D(o[652]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[652]) );
  DFF \round_reg_reg[653]  ( .D(o[653]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[653]) );
  DFF \round_reg_reg[654]  ( .D(o[654]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[654]) );
  DFF \round_reg_reg[655]  ( .D(o[655]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[655]) );
  DFF \round_reg_reg[656]  ( .D(o[656]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[656]) );
  DFF \round_reg_reg[657]  ( .D(o[657]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[657]) );
  DFF \round_reg_reg[658]  ( .D(o[658]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[658]) );
  DFF \round_reg_reg[659]  ( .D(o[659]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[659]) );
  DFF \round_reg_reg[660]  ( .D(o[660]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[660]) );
  DFF \round_reg_reg[661]  ( .D(o[661]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[661]) );
  DFF \round_reg_reg[662]  ( .D(o[662]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[662]) );
  DFF \round_reg_reg[663]  ( .D(o[663]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[663]) );
  DFF \round_reg_reg[664]  ( .D(o[664]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[664]) );
  DFF \round_reg_reg[665]  ( .D(o[665]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[665]) );
  DFF \round_reg_reg[666]  ( .D(o[666]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[666]) );
  DFF \round_reg_reg[667]  ( .D(o[667]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[667]) );
  DFF \round_reg_reg[668]  ( .D(o[668]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[668]) );
  DFF \round_reg_reg[669]  ( .D(o[669]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[669]) );
  DFF \round_reg_reg[670]  ( .D(o[670]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[670]) );
  DFF \round_reg_reg[671]  ( .D(o[671]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[671]) );
  DFF \round_reg_reg[672]  ( .D(o[672]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[672]) );
  DFF \round_reg_reg[673]  ( .D(o[673]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[673]) );
  DFF \round_reg_reg[674]  ( .D(o[674]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[674]) );
  DFF \round_reg_reg[675]  ( .D(o[675]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[675]) );
  DFF \round_reg_reg[676]  ( .D(o[676]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[676]) );
  DFF \round_reg_reg[677]  ( .D(o[677]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[677]) );
  DFF \round_reg_reg[678]  ( .D(o[678]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[678]) );
  DFF \round_reg_reg[679]  ( .D(o[679]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[679]) );
  DFF \round_reg_reg[680]  ( .D(o[680]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[680]) );
  DFF \round_reg_reg[681]  ( .D(o[681]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[681]) );
  DFF \round_reg_reg[682]  ( .D(o[682]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[682]) );
  DFF \round_reg_reg[683]  ( .D(o[683]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[683]) );
  DFF \round_reg_reg[684]  ( .D(o[684]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[684]) );
  DFF \round_reg_reg[685]  ( .D(o[685]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[685]) );
  DFF \round_reg_reg[686]  ( .D(o[686]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[686]) );
  DFF \round_reg_reg[687]  ( .D(o[687]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[687]) );
  DFF \round_reg_reg[688]  ( .D(o[688]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[688]) );
  DFF \round_reg_reg[689]  ( .D(o[689]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[689]) );
  DFF \round_reg_reg[690]  ( .D(o[690]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[690]) );
  DFF \round_reg_reg[691]  ( .D(o[691]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[691]) );
  DFF \round_reg_reg[692]  ( .D(o[692]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[692]) );
  DFF \round_reg_reg[693]  ( .D(o[693]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[693]) );
  DFF \round_reg_reg[694]  ( .D(o[694]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[694]) );
  DFF \round_reg_reg[695]  ( .D(o[695]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[695]) );
  DFF \round_reg_reg[696]  ( .D(o[696]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[696]) );
  DFF \round_reg_reg[697]  ( .D(o[697]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[697]) );
  DFF \round_reg_reg[698]  ( .D(o[698]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[698]) );
  DFF \round_reg_reg[699]  ( .D(o[699]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[699]) );
  DFF \round_reg_reg[700]  ( .D(o[700]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[700]) );
  DFF \round_reg_reg[701]  ( .D(o[701]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[701]) );
  DFF \round_reg_reg[702]  ( .D(o[702]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[702]) );
  DFF \round_reg_reg[703]  ( .D(o[703]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[703]) );
  DFF \round_reg_reg[704]  ( .D(o[704]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[704]) );
  DFF \round_reg_reg[705]  ( .D(o[705]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[705]) );
  DFF \round_reg_reg[706]  ( .D(o[706]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[706]) );
  DFF \round_reg_reg[707]  ( .D(o[707]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[707]) );
  DFF \round_reg_reg[708]  ( .D(o[708]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[708]) );
  DFF \round_reg_reg[709]  ( .D(o[709]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[709]) );
  DFF \round_reg_reg[710]  ( .D(o[710]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[710]) );
  DFF \round_reg_reg[711]  ( .D(o[711]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[711]) );
  DFF \round_reg_reg[712]  ( .D(o[712]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[712]) );
  DFF \round_reg_reg[713]  ( .D(o[713]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[713]) );
  DFF \round_reg_reg[714]  ( .D(o[714]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[714]) );
  DFF \round_reg_reg[715]  ( .D(o[715]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[715]) );
  DFF \round_reg_reg[716]  ( .D(o[716]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[716]) );
  DFF \round_reg_reg[717]  ( .D(o[717]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[717]) );
  DFF \round_reg_reg[718]  ( .D(o[718]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[718]) );
  DFF \round_reg_reg[719]  ( .D(o[719]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[719]) );
  DFF \round_reg_reg[720]  ( .D(o[720]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[720]) );
  DFF \round_reg_reg[721]  ( .D(o[721]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[721]) );
  DFF \round_reg_reg[722]  ( .D(o[722]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[722]) );
  DFF \round_reg_reg[723]  ( .D(o[723]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[723]) );
  DFF \round_reg_reg[724]  ( .D(o[724]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[724]) );
  DFF \round_reg_reg[725]  ( .D(o[725]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[725]) );
  DFF \round_reg_reg[726]  ( .D(o[726]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[726]) );
  DFF \round_reg_reg[727]  ( .D(o[727]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[727]) );
  DFF \round_reg_reg[728]  ( .D(o[728]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[728]) );
  DFF \round_reg_reg[729]  ( .D(o[729]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[729]) );
  DFF \round_reg_reg[730]  ( .D(o[730]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[730]) );
  DFF \round_reg_reg[731]  ( .D(o[731]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[731]) );
  DFF \round_reg_reg[732]  ( .D(o[732]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[732]) );
  DFF \round_reg_reg[733]  ( .D(o[733]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[733]) );
  DFF \round_reg_reg[734]  ( .D(o[734]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[734]) );
  DFF \round_reg_reg[735]  ( .D(o[735]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[735]) );
  DFF \round_reg_reg[736]  ( .D(o[736]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[736]) );
  DFF \round_reg_reg[737]  ( .D(o[737]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[737]) );
  DFF \round_reg_reg[738]  ( .D(o[738]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[738]) );
  DFF \round_reg_reg[739]  ( .D(o[739]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[739]) );
  DFF \round_reg_reg[740]  ( .D(o[740]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[740]) );
  DFF \round_reg_reg[741]  ( .D(o[741]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[741]) );
  DFF \round_reg_reg[742]  ( .D(o[742]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[742]) );
  DFF \round_reg_reg[743]  ( .D(o[743]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[743]) );
  DFF \round_reg_reg[744]  ( .D(o[744]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[744]) );
  DFF \round_reg_reg[745]  ( .D(o[745]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[745]) );
  DFF \round_reg_reg[746]  ( .D(o[746]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[746]) );
  DFF \round_reg_reg[747]  ( .D(o[747]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[747]) );
  DFF \round_reg_reg[748]  ( .D(o[748]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[748]) );
  DFF \round_reg_reg[749]  ( .D(o[749]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[749]) );
  DFF \round_reg_reg[750]  ( .D(o[750]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[750]) );
  DFF \round_reg_reg[751]  ( .D(o[751]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[751]) );
  DFF \round_reg_reg[752]  ( .D(o[752]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[752]) );
  DFF \round_reg_reg[753]  ( .D(o[753]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[753]) );
  DFF \round_reg_reg[754]  ( .D(o[754]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[754]) );
  DFF \round_reg_reg[755]  ( .D(o[755]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[755]) );
  DFF \round_reg_reg[756]  ( .D(o[756]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[756]) );
  DFF \round_reg_reg[757]  ( .D(o[757]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[757]) );
  DFF \round_reg_reg[758]  ( .D(o[758]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[758]) );
  DFF \round_reg_reg[759]  ( .D(o[759]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[759]) );
  DFF \round_reg_reg[760]  ( .D(o[760]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[760]) );
  DFF \round_reg_reg[761]  ( .D(o[761]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[761]) );
  DFF \round_reg_reg[762]  ( .D(o[762]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[762]) );
  DFF \round_reg_reg[763]  ( .D(o[763]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[763]) );
  DFF \round_reg_reg[764]  ( .D(o[764]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[764]) );
  DFF \round_reg_reg[765]  ( .D(o[765]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[765]) );
  DFF \round_reg_reg[766]  ( .D(o[766]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[766]) );
  DFF \round_reg_reg[767]  ( .D(o[767]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[767]) );
  DFF \round_reg_reg[768]  ( .D(o[768]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[768]) );
  DFF \round_reg_reg[769]  ( .D(o[769]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[769]) );
  DFF \round_reg_reg[770]  ( .D(o[770]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[770]) );
  DFF \round_reg_reg[771]  ( .D(o[771]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[771]) );
  DFF \round_reg_reg[772]  ( .D(o[772]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[772]) );
  DFF \round_reg_reg[773]  ( .D(o[773]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[773]) );
  DFF \round_reg_reg[774]  ( .D(o[774]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[774]) );
  DFF \round_reg_reg[775]  ( .D(o[775]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[775]) );
  DFF \round_reg_reg[776]  ( .D(o[776]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[776]) );
  DFF \round_reg_reg[777]  ( .D(o[777]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[777]) );
  DFF \round_reg_reg[778]  ( .D(o[778]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[778]) );
  DFF \round_reg_reg[779]  ( .D(o[779]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[779]) );
  DFF \round_reg_reg[780]  ( .D(o[780]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[780]) );
  DFF \round_reg_reg[781]  ( .D(o[781]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[781]) );
  DFF \round_reg_reg[782]  ( .D(o[782]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[782]) );
  DFF \round_reg_reg[783]  ( .D(o[783]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[783]) );
  DFF \round_reg_reg[784]  ( .D(o[784]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[784]) );
  DFF \round_reg_reg[785]  ( .D(o[785]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[785]) );
  DFF \round_reg_reg[786]  ( .D(o[786]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[786]) );
  DFF \round_reg_reg[787]  ( .D(o[787]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[787]) );
  DFF \round_reg_reg[788]  ( .D(o[788]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[788]) );
  DFF \round_reg_reg[789]  ( .D(o[789]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[789]) );
  DFF \round_reg_reg[790]  ( .D(o[790]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[790]) );
  DFF \round_reg_reg[791]  ( .D(o[791]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[791]) );
  DFF \round_reg_reg[792]  ( .D(o[792]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[792]) );
  DFF \round_reg_reg[793]  ( .D(o[793]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[793]) );
  DFF \round_reg_reg[794]  ( .D(o[794]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[794]) );
  DFF \round_reg_reg[795]  ( .D(o[795]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[795]) );
  DFF \round_reg_reg[796]  ( .D(o[796]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[796]) );
  DFF \round_reg_reg[797]  ( .D(o[797]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[797]) );
  DFF \round_reg_reg[798]  ( .D(o[798]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[798]) );
  DFF \round_reg_reg[799]  ( .D(o[799]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[799]) );
  DFF \round_reg_reg[800]  ( .D(o[800]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[800]) );
  DFF \round_reg_reg[801]  ( .D(o[801]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[801]) );
  DFF \round_reg_reg[802]  ( .D(o[802]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[802]) );
  DFF \round_reg_reg[803]  ( .D(o[803]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[803]) );
  DFF \round_reg_reg[804]  ( .D(o[804]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[804]) );
  DFF \round_reg_reg[805]  ( .D(o[805]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[805]) );
  DFF \round_reg_reg[806]  ( .D(o[806]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[806]) );
  DFF \round_reg_reg[807]  ( .D(o[807]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[807]) );
  DFF \round_reg_reg[808]  ( .D(o[808]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[808]) );
  DFF \round_reg_reg[809]  ( .D(o[809]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[809]) );
  DFF \round_reg_reg[810]  ( .D(o[810]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[810]) );
  DFF \round_reg_reg[811]  ( .D(o[811]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[811]) );
  DFF \round_reg_reg[812]  ( .D(o[812]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[812]) );
  DFF \round_reg_reg[813]  ( .D(o[813]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[813]) );
  DFF \round_reg_reg[814]  ( .D(o[814]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[814]) );
  DFF \round_reg_reg[815]  ( .D(o[815]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[815]) );
  DFF \round_reg_reg[816]  ( .D(o[816]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[816]) );
  DFF \round_reg_reg[817]  ( .D(o[817]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[817]) );
  DFF \round_reg_reg[818]  ( .D(o[818]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[818]) );
  DFF \round_reg_reg[819]  ( .D(o[819]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[819]) );
  DFF \round_reg_reg[820]  ( .D(o[820]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[820]) );
  DFF \round_reg_reg[821]  ( .D(o[821]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[821]) );
  DFF \round_reg_reg[822]  ( .D(o[822]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[822]) );
  DFF \round_reg_reg[823]  ( .D(o[823]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[823]) );
  DFF \round_reg_reg[824]  ( .D(o[824]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[824]) );
  DFF \round_reg_reg[825]  ( .D(o[825]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[825]) );
  DFF \round_reg_reg[826]  ( .D(o[826]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[826]) );
  DFF \round_reg_reg[827]  ( .D(o[827]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[827]) );
  DFF \round_reg_reg[828]  ( .D(o[828]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[828]) );
  DFF \round_reg_reg[829]  ( .D(o[829]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[829]) );
  DFF \round_reg_reg[830]  ( .D(o[830]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[830]) );
  DFF \round_reg_reg[831]  ( .D(o[831]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[831]) );
  DFF \round_reg_reg[832]  ( .D(o[832]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[832]) );
  DFF \round_reg_reg[833]  ( .D(o[833]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[833]) );
  DFF \round_reg_reg[834]  ( .D(o[834]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[834]) );
  DFF \round_reg_reg[835]  ( .D(o[835]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[835]) );
  DFF \round_reg_reg[836]  ( .D(o[836]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[836]) );
  DFF \round_reg_reg[837]  ( .D(o[837]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[837]) );
  DFF \round_reg_reg[838]  ( .D(o[838]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[838]) );
  DFF \round_reg_reg[839]  ( .D(o[839]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[839]) );
  DFF \round_reg_reg[840]  ( .D(o[840]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[840]) );
  DFF \round_reg_reg[841]  ( .D(o[841]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[841]) );
  DFF \round_reg_reg[842]  ( .D(o[842]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[842]) );
  DFF \round_reg_reg[843]  ( .D(o[843]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[843]) );
  DFF \round_reg_reg[844]  ( .D(o[844]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[844]) );
  DFF \round_reg_reg[845]  ( .D(o[845]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[845]) );
  DFF \round_reg_reg[846]  ( .D(o[846]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[846]) );
  DFF \round_reg_reg[847]  ( .D(o[847]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[847]) );
  DFF \round_reg_reg[848]  ( .D(o[848]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[848]) );
  DFF \round_reg_reg[849]  ( .D(o[849]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[849]) );
  DFF \round_reg_reg[850]  ( .D(o[850]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[850]) );
  DFF \round_reg_reg[851]  ( .D(o[851]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[851]) );
  DFF \round_reg_reg[852]  ( .D(o[852]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[852]) );
  DFF \round_reg_reg[853]  ( .D(o[853]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[853]) );
  DFF \round_reg_reg[854]  ( .D(o[854]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[854]) );
  DFF \round_reg_reg[855]  ( .D(o[855]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[855]) );
  DFF \round_reg_reg[856]  ( .D(o[856]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[856]) );
  DFF \round_reg_reg[857]  ( .D(o[857]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[857]) );
  DFF \round_reg_reg[858]  ( .D(o[858]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[858]) );
  DFF \round_reg_reg[859]  ( .D(o[859]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[859]) );
  DFF \round_reg_reg[860]  ( .D(o[860]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[860]) );
  DFF \round_reg_reg[861]  ( .D(o[861]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[861]) );
  DFF \round_reg_reg[862]  ( .D(o[862]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[862]) );
  DFF \round_reg_reg[863]  ( .D(o[863]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[863]) );
  DFF \round_reg_reg[864]  ( .D(o[864]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[864]) );
  DFF \round_reg_reg[865]  ( .D(o[865]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[865]) );
  DFF \round_reg_reg[866]  ( .D(o[866]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[866]) );
  DFF \round_reg_reg[867]  ( .D(o[867]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[867]) );
  DFF \round_reg_reg[868]  ( .D(o[868]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[868]) );
  DFF \round_reg_reg[869]  ( .D(o[869]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[869]) );
  DFF \round_reg_reg[870]  ( .D(o[870]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[870]) );
  DFF \round_reg_reg[871]  ( .D(o[871]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[871]) );
  DFF \round_reg_reg[872]  ( .D(o[872]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[872]) );
  DFF \round_reg_reg[873]  ( .D(o[873]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[873]) );
  DFF \round_reg_reg[874]  ( .D(o[874]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[874]) );
  DFF \round_reg_reg[875]  ( .D(o[875]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[875]) );
  DFF \round_reg_reg[876]  ( .D(o[876]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[876]) );
  DFF \round_reg_reg[877]  ( .D(o[877]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[877]) );
  DFF \round_reg_reg[878]  ( .D(o[878]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[878]) );
  DFF \round_reg_reg[879]  ( .D(o[879]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[879]) );
  DFF \round_reg_reg[880]  ( .D(o[880]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[880]) );
  DFF \round_reg_reg[881]  ( .D(o[881]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[881]) );
  DFF \round_reg_reg[882]  ( .D(o[882]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[882]) );
  DFF \round_reg_reg[883]  ( .D(o[883]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[883]) );
  DFF \round_reg_reg[884]  ( .D(o[884]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[884]) );
  DFF \round_reg_reg[885]  ( .D(o[885]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[885]) );
  DFF \round_reg_reg[886]  ( .D(o[886]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[886]) );
  DFF \round_reg_reg[887]  ( .D(o[887]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[887]) );
  DFF \round_reg_reg[888]  ( .D(o[888]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[888]) );
  DFF \round_reg_reg[889]  ( .D(o[889]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[889]) );
  DFF \round_reg_reg[890]  ( .D(o[890]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[890]) );
  DFF \round_reg_reg[891]  ( .D(o[891]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[891]) );
  DFF \round_reg_reg[892]  ( .D(o[892]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[892]) );
  DFF \round_reg_reg[893]  ( .D(o[893]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[893]) );
  DFF \round_reg_reg[894]  ( .D(o[894]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[894]) );
  DFF \round_reg_reg[895]  ( .D(o[895]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[895]) );
  DFF \round_reg_reg[896]  ( .D(o[896]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[896]) );
  DFF \round_reg_reg[897]  ( .D(o[897]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[897]) );
  DFF \round_reg_reg[898]  ( .D(o[898]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[898]) );
  DFF \round_reg_reg[899]  ( .D(o[899]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[899]) );
  DFF \round_reg_reg[900]  ( .D(o[900]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[900]) );
  DFF \round_reg_reg[901]  ( .D(o[901]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[901]) );
  DFF \round_reg_reg[902]  ( .D(o[902]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[902]) );
  DFF \round_reg_reg[903]  ( .D(o[903]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[903]) );
  DFF \round_reg_reg[904]  ( .D(o[904]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[904]) );
  DFF \round_reg_reg[905]  ( .D(o[905]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[905]) );
  DFF \round_reg_reg[906]  ( .D(o[906]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[906]) );
  DFF \round_reg_reg[907]  ( .D(o[907]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[907]) );
  DFF \round_reg_reg[908]  ( .D(o[908]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[908]) );
  DFF \round_reg_reg[909]  ( .D(o[909]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[909]) );
  DFF \round_reg_reg[910]  ( .D(o[910]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[910]) );
  DFF \round_reg_reg[911]  ( .D(o[911]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[911]) );
  DFF \round_reg_reg[912]  ( .D(o[912]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[912]) );
  DFF \round_reg_reg[913]  ( .D(o[913]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[913]) );
  DFF \round_reg_reg[914]  ( .D(o[914]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[914]) );
  DFF \round_reg_reg[915]  ( .D(o[915]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[915]) );
  DFF \round_reg_reg[916]  ( .D(o[916]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[916]) );
  DFF \round_reg_reg[917]  ( .D(o[917]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[917]) );
  DFF \round_reg_reg[918]  ( .D(o[918]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[918]) );
  DFF \round_reg_reg[919]  ( .D(o[919]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[919]) );
  DFF \round_reg_reg[920]  ( .D(o[920]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[920]) );
  DFF \round_reg_reg[921]  ( .D(o[921]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[921]) );
  DFF \round_reg_reg[922]  ( .D(o[922]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[922]) );
  DFF \round_reg_reg[923]  ( .D(o[923]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[923]) );
  DFF \round_reg_reg[924]  ( .D(o[924]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[924]) );
  DFF \round_reg_reg[925]  ( .D(o[925]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[925]) );
  DFF \round_reg_reg[926]  ( .D(o[926]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[926]) );
  DFF \round_reg_reg[927]  ( .D(o[927]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[927]) );
  DFF \round_reg_reg[928]  ( .D(o[928]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[928]) );
  DFF \round_reg_reg[929]  ( .D(o[929]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[929]) );
  DFF \round_reg_reg[930]  ( .D(o[930]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[930]) );
  DFF \round_reg_reg[931]  ( .D(o[931]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[931]) );
  DFF \round_reg_reg[932]  ( .D(o[932]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[932]) );
  DFF \round_reg_reg[933]  ( .D(o[933]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[933]) );
  DFF \round_reg_reg[934]  ( .D(o[934]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[934]) );
  DFF \round_reg_reg[935]  ( .D(o[935]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[935]) );
  DFF \round_reg_reg[936]  ( .D(o[936]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[936]) );
  DFF \round_reg_reg[937]  ( .D(o[937]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[937]) );
  DFF \round_reg_reg[938]  ( .D(o[938]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[938]) );
  DFF \round_reg_reg[939]  ( .D(o[939]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[939]) );
  DFF \round_reg_reg[940]  ( .D(o[940]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[940]) );
  DFF \round_reg_reg[941]  ( .D(o[941]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[941]) );
  DFF \round_reg_reg[942]  ( .D(o[942]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[942]) );
  DFF \round_reg_reg[943]  ( .D(o[943]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[943]) );
  DFF \round_reg_reg[944]  ( .D(o[944]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[944]) );
  DFF \round_reg_reg[945]  ( .D(o[945]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[945]) );
  DFF \round_reg_reg[946]  ( .D(o[946]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[946]) );
  DFF \round_reg_reg[947]  ( .D(o[947]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[947]) );
  DFF \round_reg_reg[948]  ( .D(o[948]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[948]) );
  DFF \round_reg_reg[949]  ( .D(o[949]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[949]) );
  DFF \round_reg_reg[950]  ( .D(o[950]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[950]) );
  DFF \round_reg_reg[951]  ( .D(o[951]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[951]) );
  DFF \round_reg_reg[952]  ( .D(o[952]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[952]) );
  DFF \round_reg_reg[953]  ( .D(o[953]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[953]) );
  DFF \round_reg_reg[954]  ( .D(o[954]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[954]) );
  DFF \round_reg_reg[955]  ( .D(o[955]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[955]) );
  DFF \round_reg_reg[956]  ( .D(o[956]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[956]) );
  DFF \round_reg_reg[957]  ( .D(o[957]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[957]) );
  DFF \round_reg_reg[958]  ( .D(o[958]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[958]) );
  DFF \round_reg_reg[959]  ( .D(o[959]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[959]) );
  DFF \round_reg_reg[960]  ( .D(o[960]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[960]) );
  DFF \round_reg_reg[961]  ( .D(o[961]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[961]) );
  DFF \round_reg_reg[962]  ( .D(o[962]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[962]) );
  DFF \round_reg_reg[963]  ( .D(o[963]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[963]) );
  DFF \round_reg_reg[964]  ( .D(o[964]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[964]) );
  DFF \round_reg_reg[965]  ( .D(o[965]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[965]) );
  DFF \round_reg_reg[966]  ( .D(o[966]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[966]) );
  DFF \round_reg_reg[967]  ( .D(o[967]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[967]) );
  DFF \round_reg_reg[968]  ( .D(o[968]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[968]) );
  DFF \round_reg_reg[969]  ( .D(o[969]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[969]) );
  DFF \round_reg_reg[970]  ( .D(o[970]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[970]) );
  DFF \round_reg_reg[971]  ( .D(o[971]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[971]) );
  DFF \round_reg_reg[972]  ( .D(o[972]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[972]) );
  DFF \round_reg_reg[973]  ( .D(o[973]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[973]) );
  DFF \round_reg_reg[974]  ( .D(o[974]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[974]) );
  DFF \round_reg_reg[975]  ( .D(o[975]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[975]) );
  DFF \round_reg_reg[976]  ( .D(o[976]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[976]) );
  DFF \round_reg_reg[977]  ( .D(o[977]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[977]) );
  DFF \round_reg_reg[978]  ( .D(o[978]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[978]) );
  DFF \round_reg_reg[979]  ( .D(o[979]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[979]) );
  DFF \round_reg_reg[980]  ( .D(o[980]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[980]) );
  DFF \round_reg_reg[981]  ( .D(o[981]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[981]) );
  DFF \round_reg_reg[982]  ( .D(o[982]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[982]) );
  DFF \round_reg_reg[983]  ( .D(o[983]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[983]) );
  DFF \round_reg_reg[984]  ( .D(o[984]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[984]) );
  DFF \round_reg_reg[985]  ( .D(o[985]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[985]) );
  DFF \round_reg_reg[986]  ( .D(o[986]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[986]) );
  DFF \round_reg_reg[987]  ( .D(o[987]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[987]) );
  DFF \round_reg_reg[988]  ( .D(o[988]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[988]) );
  DFF \round_reg_reg[989]  ( .D(o[989]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[989]) );
  DFF \round_reg_reg[990]  ( .D(o[990]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[990]) );
  DFF \round_reg_reg[991]  ( .D(o[991]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[991]) );
  DFF \round_reg_reg[992]  ( .D(o[992]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[992]) );
  DFF \round_reg_reg[993]  ( .D(o[993]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[993]) );
  DFF \round_reg_reg[994]  ( .D(o[994]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[994]) );
  DFF \round_reg_reg[995]  ( .D(o[995]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[995]) );
  DFF \round_reg_reg[996]  ( .D(o[996]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[996]) );
  DFF \round_reg_reg[997]  ( .D(o[997]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[997]) );
  DFF \round_reg_reg[998]  ( .D(o[998]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[998]) );
  DFF \round_reg_reg[999]  ( .D(o[999]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[999]) );
  DFF \round_reg_reg[1000]  ( .D(o[1000]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1000]) );
  DFF \round_reg_reg[1001]  ( .D(o[1001]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1001]) );
  DFF \round_reg_reg[1002]  ( .D(o[1002]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1002]) );
  DFF \round_reg_reg[1003]  ( .D(o[1003]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1003]) );
  DFF \round_reg_reg[1004]  ( .D(o[1004]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1004]) );
  DFF \round_reg_reg[1005]  ( .D(o[1005]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1005]) );
  DFF \round_reg_reg[1006]  ( .D(o[1006]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1006]) );
  DFF \round_reg_reg[1007]  ( .D(o[1007]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1007]) );
  DFF \round_reg_reg[1008]  ( .D(o[1008]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1008]) );
  DFF \round_reg_reg[1009]  ( .D(o[1009]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1009]) );
  DFF \round_reg_reg[1010]  ( .D(o[1010]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1010]) );
  DFF \round_reg_reg[1011]  ( .D(o[1011]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1011]) );
  DFF \round_reg_reg[1012]  ( .D(o[1012]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1012]) );
  DFF \round_reg_reg[1013]  ( .D(o[1013]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1013]) );
  DFF \round_reg_reg[1014]  ( .D(o[1014]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1014]) );
  DFF \round_reg_reg[1015]  ( .D(o[1015]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1015]) );
  DFF \round_reg_reg[1016]  ( .D(o[1016]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1016]) );
  DFF \round_reg_reg[1017]  ( .D(o[1017]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1017]) );
  DFF \round_reg_reg[1018]  ( .D(o[1018]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1018]) );
  DFF \round_reg_reg[1019]  ( .D(o[1019]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1019]) );
  DFF \round_reg_reg[1020]  ( .D(o[1020]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1020]) );
  DFF \round_reg_reg[1021]  ( .D(o[1021]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1021]) );
  DFF \round_reg_reg[1022]  ( .D(o[1022]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1022]) );
  DFF \round_reg_reg[1023]  ( .D(o[1023]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1023]) );
  DFF \round_reg_reg[1024]  ( .D(o[1024]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1024]) );
  DFF \round_reg_reg[1025]  ( .D(o[1025]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1025]) );
  DFF \round_reg_reg[1026]  ( .D(o[1026]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1026]) );
  DFF \round_reg_reg[1027]  ( .D(o[1027]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1027]) );
  DFF \round_reg_reg[1028]  ( .D(o[1028]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1028]) );
  DFF \round_reg_reg[1029]  ( .D(o[1029]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1029]) );
  DFF \round_reg_reg[1030]  ( .D(o[1030]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1030]) );
  DFF \round_reg_reg[1031]  ( .D(o[1031]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1031]) );
  DFF \round_reg_reg[1032]  ( .D(o[1032]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1032]) );
  DFF \round_reg_reg[1033]  ( .D(o[1033]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1033]) );
  DFF \round_reg_reg[1034]  ( .D(o[1034]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1034]) );
  DFF \round_reg_reg[1035]  ( .D(o[1035]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1035]) );
  DFF \round_reg_reg[1036]  ( .D(o[1036]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1036]) );
  DFF \round_reg_reg[1037]  ( .D(o[1037]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1037]) );
  DFF \round_reg_reg[1038]  ( .D(o[1038]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1038]) );
  DFF \round_reg_reg[1039]  ( .D(o[1039]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1039]) );
  DFF \round_reg_reg[1040]  ( .D(o[1040]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1040]) );
  DFF \round_reg_reg[1041]  ( .D(o[1041]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1041]) );
  DFF \round_reg_reg[1042]  ( .D(o[1042]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1042]) );
  DFF \round_reg_reg[1043]  ( .D(o[1043]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1043]) );
  DFF \round_reg_reg[1044]  ( .D(o[1044]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1044]) );
  DFF \round_reg_reg[1045]  ( .D(o[1045]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1045]) );
  DFF \round_reg_reg[1046]  ( .D(o[1046]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1046]) );
  DFF \round_reg_reg[1047]  ( .D(o[1047]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1047]) );
  DFF \round_reg_reg[1048]  ( .D(o[1048]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1048]) );
  DFF \round_reg_reg[1049]  ( .D(o[1049]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1049]) );
  DFF \round_reg_reg[1050]  ( .D(o[1050]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1050]) );
  DFF \round_reg_reg[1051]  ( .D(o[1051]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1051]) );
  DFF \round_reg_reg[1052]  ( .D(o[1052]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1052]) );
  DFF \round_reg_reg[1053]  ( .D(o[1053]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1053]) );
  DFF \round_reg_reg[1054]  ( .D(o[1054]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1054]) );
  DFF \round_reg_reg[1055]  ( .D(o[1055]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1055]) );
  DFF \round_reg_reg[1056]  ( .D(o[1056]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1056]) );
  DFF \round_reg_reg[1057]  ( .D(o[1057]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1057]) );
  DFF \round_reg_reg[1058]  ( .D(o[1058]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1058]) );
  DFF \round_reg_reg[1059]  ( .D(o[1059]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1059]) );
  DFF \round_reg_reg[1060]  ( .D(o[1060]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1060]) );
  DFF \round_reg_reg[1061]  ( .D(o[1061]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1061]) );
  DFF \round_reg_reg[1062]  ( .D(o[1062]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1062]) );
  DFF \round_reg_reg[1063]  ( .D(o[1063]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1063]) );
  DFF \round_reg_reg[1064]  ( .D(o[1064]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1064]) );
  DFF \round_reg_reg[1065]  ( .D(o[1065]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1065]) );
  DFF \round_reg_reg[1066]  ( .D(o[1066]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1066]) );
  DFF \round_reg_reg[1067]  ( .D(o[1067]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1067]) );
  DFF \round_reg_reg[1068]  ( .D(o[1068]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1068]) );
  DFF \round_reg_reg[1069]  ( .D(o[1069]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1069]) );
  DFF \round_reg_reg[1070]  ( .D(o[1070]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1070]) );
  DFF \round_reg_reg[1071]  ( .D(o[1071]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1071]) );
  DFF \round_reg_reg[1072]  ( .D(o[1072]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1072]) );
  DFF \round_reg_reg[1073]  ( .D(o[1073]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1073]) );
  DFF \round_reg_reg[1074]  ( .D(o[1074]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1074]) );
  DFF \round_reg_reg[1075]  ( .D(o[1075]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1075]) );
  DFF \round_reg_reg[1076]  ( .D(o[1076]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1076]) );
  DFF \round_reg_reg[1077]  ( .D(o[1077]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1077]) );
  DFF \round_reg_reg[1078]  ( .D(o[1078]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1078]) );
  DFF \round_reg_reg[1079]  ( .D(o[1079]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1079]) );
  DFF \round_reg_reg[1080]  ( .D(o[1080]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1080]) );
  DFF \round_reg_reg[1081]  ( .D(o[1081]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1081]) );
  DFF \round_reg_reg[1082]  ( .D(o[1082]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1082]) );
  DFF \round_reg_reg[1083]  ( .D(o[1083]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1083]) );
  DFF \round_reg_reg[1084]  ( .D(o[1084]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1084]) );
  DFF \round_reg_reg[1085]  ( .D(o[1085]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1085]) );
  DFF \round_reg_reg[1086]  ( .D(o[1086]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1086]) );
  DFF \round_reg_reg[1087]  ( .D(o[1087]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1087]) );
  DFF \round_reg_reg[1088]  ( .D(o[1088]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1088]) );
  DFF \round_reg_reg[1089]  ( .D(o[1089]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1089]) );
  DFF \round_reg_reg[1090]  ( .D(o[1090]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1090]) );
  DFF \round_reg_reg[1091]  ( .D(o[1091]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1091]) );
  DFF \round_reg_reg[1092]  ( .D(o[1092]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1092]) );
  DFF \round_reg_reg[1093]  ( .D(o[1093]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1093]) );
  DFF \round_reg_reg[1094]  ( .D(o[1094]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1094]) );
  DFF \round_reg_reg[1095]  ( .D(o[1095]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1095]) );
  DFF \round_reg_reg[1096]  ( .D(o[1096]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1096]) );
  DFF \round_reg_reg[1097]  ( .D(o[1097]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1097]) );
  DFF \round_reg_reg[1098]  ( .D(o[1098]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1098]) );
  DFF \round_reg_reg[1099]  ( .D(o[1099]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1099]) );
  DFF \round_reg_reg[1100]  ( .D(o[1100]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1100]) );
  DFF \round_reg_reg[1101]  ( .D(o[1101]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1101]) );
  DFF \round_reg_reg[1102]  ( .D(o[1102]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1102]) );
  DFF \round_reg_reg[1103]  ( .D(o[1103]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1103]) );
  DFF \round_reg_reg[1104]  ( .D(o[1104]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1104]) );
  DFF \round_reg_reg[1105]  ( .D(o[1105]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1105]) );
  DFF \round_reg_reg[1106]  ( .D(o[1106]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1106]) );
  DFF \round_reg_reg[1107]  ( .D(o[1107]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1107]) );
  DFF \round_reg_reg[1108]  ( .D(o[1108]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1108]) );
  DFF \round_reg_reg[1109]  ( .D(o[1109]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1109]) );
  DFF \round_reg_reg[1110]  ( .D(o[1110]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1110]) );
  DFF \round_reg_reg[1111]  ( .D(o[1111]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1111]) );
  DFF \round_reg_reg[1112]  ( .D(o[1112]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1112]) );
  DFF \round_reg_reg[1113]  ( .D(o[1113]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1113]) );
  DFF \round_reg_reg[1114]  ( .D(o[1114]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1114]) );
  DFF \round_reg_reg[1115]  ( .D(o[1115]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1115]) );
  DFF \round_reg_reg[1116]  ( .D(o[1116]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1116]) );
  DFF \round_reg_reg[1117]  ( .D(o[1117]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1117]) );
  DFF \round_reg_reg[1118]  ( .D(o[1118]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1118]) );
  DFF \round_reg_reg[1119]  ( .D(o[1119]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1119]) );
  DFF \round_reg_reg[1120]  ( .D(o[1120]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1120]) );
  DFF \round_reg_reg[1121]  ( .D(o[1121]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1121]) );
  DFF \round_reg_reg[1122]  ( .D(o[1122]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1122]) );
  DFF \round_reg_reg[1123]  ( .D(o[1123]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1123]) );
  DFF \round_reg_reg[1124]  ( .D(o[1124]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1124]) );
  DFF \round_reg_reg[1125]  ( .D(o[1125]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1125]) );
  DFF \round_reg_reg[1126]  ( .D(o[1126]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1126]) );
  DFF \round_reg_reg[1127]  ( .D(o[1127]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1127]) );
  DFF \round_reg_reg[1128]  ( .D(o[1128]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1128]) );
  DFF \round_reg_reg[1129]  ( .D(o[1129]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1129]) );
  DFF \round_reg_reg[1130]  ( .D(o[1130]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1130]) );
  DFF \round_reg_reg[1131]  ( .D(o[1131]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1131]) );
  DFF \round_reg_reg[1132]  ( .D(o[1132]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1132]) );
  DFF \round_reg_reg[1133]  ( .D(o[1133]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1133]) );
  DFF \round_reg_reg[1134]  ( .D(o[1134]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1134]) );
  DFF \round_reg_reg[1135]  ( .D(o[1135]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1135]) );
  DFF \round_reg_reg[1136]  ( .D(o[1136]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1136]) );
  DFF \round_reg_reg[1137]  ( .D(o[1137]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1137]) );
  DFF \round_reg_reg[1138]  ( .D(o[1138]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1138]) );
  DFF \round_reg_reg[1139]  ( .D(o[1139]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1139]) );
  DFF \round_reg_reg[1140]  ( .D(o[1140]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1140]) );
  DFF \round_reg_reg[1141]  ( .D(o[1141]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1141]) );
  DFF \round_reg_reg[1142]  ( .D(o[1142]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1142]) );
  DFF \round_reg_reg[1143]  ( .D(o[1143]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1143]) );
  DFF \round_reg_reg[1144]  ( .D(o[1144]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1144]) );
  DFF \round_reg_reg[1145]  ( .D(o[1145]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1145]) );
  DFF \round_reg_reg[1146]  ( .D(o[1146]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1146]) );
  DFF \round_reg_reg[1147]  ( .D(o[1147]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1147]) );
  DFF \round_reg_reg[1148]  ( .D(o[1148]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1148]) );
  DFF \round_reg_reg[1149]  ( .D(o[1149]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1149]) );
  DFF \round_reg_reg[1150]  ( .D(o[1150]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1150]) );
  DFF \round_reg_reg[1151]  ( .D(o[1151]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1151]) );
  DFF \round_reg_reg[1152]  ( .D(o[1152]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1152]) );
  DFF \round_reg_reg[1153]  ( .D(o[1153]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1153]) );
  DFF \round_reg_reg[1154]  ( .D(o[1154]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1154]) );
  DFF \round_reg_reg[1155]  ( .D(o[1155]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1155]) );
  DFF \round_reg_reg[1156]  ( .D(o[1156]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1156]) );
  DFF \round_reg_reg[1157]  ( .D(o[1157]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1157]) );
  DFF \round_reg_reg[1158]  ( .D(o[1158]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1158]) );
  DFF \round_reg_reg[1159]  ( .D(o[1159]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1159]) );
  DFF \round_reg_reg[1160]  ( .D(o[1160]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1160]) );
  DFF \round_reg_reg[1161]  ( .D(o[1161]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1161]) );
  DFF \round_reg_reg[1162]  ( .D(o[1162]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1162]) );
  DFF \round_reg_reg[1163]  ( .D(o[1163]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1163]) );
  DFF \round_reg_reg[1164]  ( .D(o[1164]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1164]) );
  DFF \round_reg_reg[1165]  ( .D(o[1165]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1165]) );
  DFF \round_reg_reg[1166]  ( .D(o[1166]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1166]) );
  DFF \round_reg_reg[1167]  ( .D(o[1167]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1167]) );
  DFF \round_reg_reg[1168]  ( .D(o[1168]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1168]) );
  DFF \round_reg_reg[1169]  ( .D(o[1169]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1169]) );
  DFF \round_reg_reg[1170]  ( .D(o[1170]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1170]) );
  DFF \round_reg_reg[1171]  ( .D(o[1171]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1171]) );
  DFF \round_reg_reg[1172]  ( .D(o[1172]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1172]) );
  DFF \round_reg_reg[1173]  ( .D(o[1173]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1173]) );
  DFF \round_reg_reg[1174]  ( .D(o[1174]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1174]) );
  DFF \round_reg_reg[1175]  ( .D(o[1175]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1175]) );
  DFF \round_reg_reg[1176]  ( .D(o[1176]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1176]) );
  DFF \round_reg_reg[1177]  ( .D(o[1177]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1177]) );
  DFF \round_reg_reg[1178]  ( .D(o[1178]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1178]) );
  DFF \round_reg_reg[1179]  ( .D(o[1179]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1179]) );
  DFF \round_reg_reg[1180]  ( .D(o[1180]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1180]) );
  DFF \round_reg_reg[1181]  ( .D(o[1181]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1181]) );
  DFF \round_reg_reg[1182]  ( .D(o[1182]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1182]) );
  DFF \round_reg_reg[1183]  ( .D(o[1183]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1183]) );
  DFF \round_reg_reg[1184]  ( .D(o[1184]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1184]) );
  DFF \round_reg_reg[1185]  ( .D(o[1185]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1185]) );
  DFF \round_reg_reg[1186]  ( .D(o[1186]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1186]) );
  DFF \round_reg_reg[1187]  ( .D(o[1187]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1187]) );
  DFF \round_reg_reg[1188]  ( .D(o[1188]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1188]) );
  DFF \round_reg_reg[1189]  ( .D(o[1189]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1189]) );
  DFF \round_reg_reg[1190]  ( .D(o[1190]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1190]) );
  DFF \round_reg_reg[1191]  ( .D(o[1191]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1191]) );
  DFF \round_reg_reg[1192]  ( .D(o[1192]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1192]) );
  DFF \round_reg_reg[1193]  ( .D(o[1193]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1193]) );
  DFF \round_reg_reg[1194]  ( .D(o[1194]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1194]) );
  DFF \round_reg_reg[1195]  ( .D(o[1195]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1195]) );
  DFF \round_reg_reg[1196]  ( .D(o[1196]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1196]) );
  DFF \round_reg_reg[1197]  ( .D(o[1197]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1197]) );
  DFF \round_reg_reg[1198]  ( .D(o[1198]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1198]) );
  DFF \round_reg_reg[1199]  ( .D(o[1199]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1199]) );
  DFF \round_reg_reg[1200]  ( .D(o[1200]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1200]) );
  DFF \round_reg_reg[1201]  ( .D(o[1201]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1201]) );
  DFF \round_reg_reg[1202]  ( .D(o[1202]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1202]) );
  DFF \round_reg_reg[1203]  ( .D(o[1203]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1203]) );
  DFF \round_reg_reg[1204]  ( .D(o[1204]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1204]) );
  DFF \round_reg_reg[1205]  ( .D(o[1205]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1205]) );
  DFF \round_reg_reg[1206]  ( .D(o[1206]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1206]) );
  DFF \round_reg_reg[1207]  ( .D(o[1207]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1207]) );
  DFF \round_reg_reg[1208]  ( .D(o[1208]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1208]) );
  DFF \round_reg_reg[1209]  ( .D(o[1209]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1209]) );
  DFF \round_reg_reg[1210]  ( .D(o[1210]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1210]) );
  DFF \round_reg_reg[1211]  ( .D(o[1211]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1211]) );
  DFF \round_reg_reg[1212]  ( .D(o[1212]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1212]) );
  DFF \round_reg_reg[1213]  ( .D(o[1213]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1213]) );
  DFF \round_reg_reg[1214]  ( .D(o[1214]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1214]) );
  DFF \round_reg_reg[1215]  ( .D(o[1215]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1215]) );
  DFF \round_reg_reg[1216]  ( .D(o[1216]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1216]) );
  DFF \round_reg_reg[1217]  ( .D(o[1217]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1217]) );
  DFF \round_reg_reg[1218]  ( .D(o[1218]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1218]) );
  DFF \round_reg_reg[1219]  ( .D(o[1219]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1219]) );
  DFF \round_reg_reg[1220]  ( .D(o[1220]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1220]) );
  DFF \round_reg_reg[1221]  ( .D(o[1221]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1221]) );
  DFF \round_reg_reg[1222]  ( .D(o[1222]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1222]) );
  DFF \round_reg_reg[1223]  ( .D(o[1223]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1223]) );
  DFF \round_reg_reg[1224]  ( .D(o[1224]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1224]) );
  DFF \round_reg_reg[1225]  ( .D(o[1225]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1225]) );
  DFF \round_reg_reg[1226]  ( .D(o[1226]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1226]) );
  DFF \round_reg_reg[1227]  ( .D(o[1227]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1227]) );
  DFF \round_reg_reg[1228]  ( .D(o[1228]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1228]) );
  DFF \round_reg_reg[1229]  ( .D(o[1229]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1229]) );
  DFF \round_reg_reg[1230]  ( .D(o[1230]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1230]) );
  DFF \round_reg_reg[1231]  ( .D(o[1231]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1231]) );
  DFF \round_reg_reg[1232]  ( .D(o[1232]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1232]) );
  DFF \round_reg_reg[1233]  ( .D(o[1233]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1233]) );
  DFF \round_reg_reg[1234]  ( .D(o[1234]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1234]) );
  DFF \round_reg_reg[1235]  ( .D(o[1235]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1235]) );
  DFF \round_reg_reg[1236]  ( .D(o[1236]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1236]) );
  DFF \round_reg_reg[1237]  ( .D(o[1237]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1237]) );
  DFF \round_reg_reg[1238]  ( .D(o[1238]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1238]) );
  DFF \round_reg_reg[1239]  ( .D(o[1239]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1239]) );
  DFF \round_reg_reg[1240]  ( .D(o[1240]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1240]) );
  DFF \round_reg_reg[1241]  ( .D(o[1241]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1241]) );
  DFF \round_reg_reg[1242]  ( .D(o[1242]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1242]) );
  DFF \round_reg_reg[1243]  ( .D(o[1243]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1243]) );
  DFF \round_reg_reg[1244]  ( .D(o[1244]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1244]) );
  DFF \round_reg_reg[1245]  ( .D(o[1245]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1245]) );
  DFF \round_reg_reg[1246]  ( .D(o[1246]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1246]) );
  DFF \round_reg_reg[1247]  ( .D(o[1247]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1247]) );
  DFF \round_reg_reg[1248]  ( .D(o[1248]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1248]) );
  DFF \round_reg_reg[1249]  ( .D(o[1249]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1249]) );
  DFF \round_reg_reg[1250]  ( .D(o[1250]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1250]) );
  DFF \round_reg_reg[1251]  ( .D(o[1251]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1251]) );
  DFF \round_reg_reg[1252]  ( .D(o[1252]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1252]) );
  DFF \round_reg_reg[1253]  ( .D(o[1253]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1253]) );
  DFF \round_reg_reg[1254]  ( .D(o[1254]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1254]) );
  DFF \round_reg_reg[1255]  ( .D(o[1255]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1255]) );
  DFF \round_reg_reg[1256]  ( .D(o[1256]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1256]) );
  DFF \round_reg_reg[1257]  ( .D(o[1257]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1257]) );
  DFF \round_reg_reg[1258]  ( .D(o[1258]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1258]) );
  DFF \round_reg_reg[1259]  ( .D(o[1259]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1259]) );
  DFF \round_reg_reg[1260]  ( .D(o[1260]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1260]) );
  DFF \round_reg_reg[1261]  ( .D(o[1261]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1261]) );
  DFF \round_reg_reg[1262]  ( .D(o[1262]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1262]) );
  DFF \round_reg_reg[1263]  ( .D(o[1263]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1263]) );
  DFF \round_reg_reg[1264]  ( .D(o[1264]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1264]) );
  DFF \round_reg_reg[1265]  ( .D(o[1265]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1265]) );
  DFF \round_reg_reg[1266]  ( .D(o[1266]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1266]) );
  DFF \round_reg_reg[1267]  ( .D(o[1267]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1267]) );
  DFF \round_reg_reg[1268]  ( .D(o[1268]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1268]) );
  DFF \round_reg_reg[1269]  ( .D(o[1269]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1269]) );
  DFF \round_reg_reg[1270]  ( .D(o[1270]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1270]) );
  DFF \round_reg_reg[1271]  ( .D(o[1271]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1271]) );
  DFF \round_reg_reg[1272]  ( .D(o[1272]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1272]) );
  DFF \round_reg_reg[1273]  ( .D(o[1273]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1273]) );
  DFF \round_reg_reg[1274]  ( .D(o[1274]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1274]) );
  DFF \round_reg_reg[1275]  ( .D(o[1275]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1275]) );
  DFF \round_reg_reg[1276]  ( .D(o[1276]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1276]) );
  DFF \round_reg_reg[1277]  ( .D(o[1277]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1277]) );
  DFF \round_reg_reg[1278]  ( .D(o[1278]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1278]) );
  DFF \round_reg_reg[1279]  ( .D(o[1279]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1279]) );
  DFF \round_reg_reg[1280]  ( .D(o[1280]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1280]) );
  DFF \round_reg_reg[1281]  ( .D(o[1281]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1281]) );
  DFF \round_reg_reg[1282]  ( .D(o[1282]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1282]) );
  DFF \round_reg_reg[1283]  ( .D(o[1283]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1283]) );
  DFF \round_reg_reg[1284]  ( .D(o[1284]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1284]) );
  DFF \round_reg_reg[1285]  ( .D(o[1285]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1285]) );
  DFF \round_reg_reg[1286]  ( .D(o[1286]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1286]) );
  DFF \round_reg_reg[1287]  ( .D(o[1287]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1287]) );
  DFF \round_reg_reg[1288]  ( .D(o[1288]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1288]) );
  DFF \round_reg_reg[1289]  ( .D(o[1289]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1289]) );
  DFF \round_reg_reg[1290]  ( .D(o[1290]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1290]) );
  DFF \round_reg_reg[1291]  ( .D(o[1291]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1291]) );
  DFF \round_reg_reg[1292]  ( .D(o[1292]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1292]) );
  DFF \round_reg_reg[1293]  ( .D(o[1293]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1293]) );
  DFF \round_reg_reg[1294]  ( .D(o[1294]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1294]) );
  DFF \round_reg_reg[1295]  ( .D(o[1295]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1295]) );
  DFF \round_reg_reg[1296]  ( .D(o[1296]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1296]) );
  DFF \round_reg_reg[1297]  ( .D(o[1297]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1297]) );
  DFF \round_reg_reg[1298]  ( .D(o[1298]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1298]) );
  DFF \round_reg_reg[1299]  ( .D(o[1299]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1299]) );
  DFF \round_reg_reg[1300]  ( .D(o[1300]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1300]) );
  DFF \round_reg_reg[1301]  ( .D(o[1301]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1301]) );
  DFF \round_reg_reg[1302]  ( .D(o[1302]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1302]) );
  DFF \round_reg_reg[1303]  ( .D(o[1303]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1303]) );
  DFF \round_reg_reg[1304]  ( .D(o[1304]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1304]) );
  DFF \round_reg_reg[1305]  ( .D(o[1305]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1305]) );
  DFF \round_reg_reg[1306]  ( .D(o[1306]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1306]) );
  DFF \round_reg_reg[1307]  ( .D(o[1307]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1307]) );
  DFF \round_reg_reg[1308]  ( .D(o[1308]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1308]) );
  DFF \round_reg_reg[1309]  ( .D(o[1309]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1309]) );
  DFF \round_reg_reg[1310]  ( .D(o[1310]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1310]) );
  DFF \round_reg_reg[1311]  ( .D(o[1311]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1311]) );
  DFF \round_reg_reg[1312]  ( .D(o[1312]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1312]) );
  DFF \round_reg_reg[1313]  ( .D(o[1313]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1313]) );
  DFF \round_reg_reg[1314]  ( .D(o[1314]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1314]) );
  DFF \round_reg_reg[1315]  ( .D(o[1315]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1315]) );
  DFF \round_reg_reg[1316]  ( .D(o[1316]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1316]) );
  DFF \round_reg_reg[1317]  ( .D(o[1317]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1317]) );
  DFF \round_reg_reg[1318]  ( .D(o[1318]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1318]) );
  DFF \round_reg_reg[1319]  ( .D(o[1319]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1319]) );
  DFF \round_reg_reg[1320]  ( .D(o[1320]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1320]) );
  DFF \round_reg_reg[1321]  ( .D(o[1321]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1321]) );
  DFF \round_reg_reg[1322]  ( .D(o[1322]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1322]) );
  DFF \round_reg_reg[1323]  ( .D(o[1323]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1323]) );
  DFF \round_reg_reg[1324]  ( .D(o[1324]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1324]) );
  DFF \round_reg_reg[1325]  ( .D(o[1325]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1325]) );
  DFF \round_reg_reg[1326]  ( .D(o[1326]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1326]) );
  DFF \round_reg_reg[1327]  ( .D(o[1327]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1327]) );
  DFF \round_reg_reg[1328]  ( .D(o[1328]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1328]) );
  DFF \round_reg_reg[1329]  ( .D(o[1329]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1329]) );
  DFF \round_reg_reg[1330]  ( .D(o[1330]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1330]) );
  DFF \round_reg_reg[1331]  ( .D(o[1331]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1331]) );
  DFF \round_reg_reg[1332]  ( .D(o[1332]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1332]) );
  DFF \round_reg_reg[1333]  ( .D(o[1333]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1333]) );
  DFF \round_reg_reg[1334]  ( .D(o[1334]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1334]) );
  DFF \round_reg_reg[1335]  ( .D(o[1335]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1335]) );
  DFF \round_reg_reg[1336]  ( .D(o[1336]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1336]) );
  DFF \round_reg_reg[1337]  ( .D(o[1337]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1337]) );
  DFF \round_reg_reg[1338]  ( .D(o[1338]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1338]) );
  DFF \round_reg_reg[1339]  ( .D(o[1339]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1339]) );
  DFF \round_reg_reg[1340]  ( .D(o[1340]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1340]) );
  DFF \round_reg_reg[1341]  ( .D(o[1341]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1341]) );
  DFF \round_reg_reg[1342]  ( .D(o[1342]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1342]) );
  DFF \round_reg_reg[1343]  ( .D(o[1343]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1343]) );
  DFF \round_reg_reg[1344]  ( .D(o[1344]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1344]) );
  DFF \round_reg_reg[1345]  ( .D(o[1345]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1345]) );
  DFF \round_reg_reg[1346]  ( .D(o[1346]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1346]) );
  DFF \round_reg_reg[1347]  ( .D(o[1347]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1347]) );
  DFF \round_reg_reg[1348]  ( .D(o[1348]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1348]) );
  DFF \round_reg_reg[1349]  ( .D(o[1349]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1349]) );
  DFF \round_reg_reg[1350]  ( .D(o[1350]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1350]) );
  DFF \round_reg_reg[1351]  ( .D(o[1351]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1351]) );
  DFF \round_reg_reg[1352]  ( .D(o[1352]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1352]) );
  DFF \round_reg_reg[1353]  ( .D(o[1353]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1353]) );
  DFF \round_reg_reg[1354]  ( .D(o[1354]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1354]) );
  DFF \round_reg_reg[1355]  ( .D(o[1355]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1355]) );
  DFF \round_reg_reg[1356]  ( .D(o[1356]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1356]) );
  DFF \round_reg_reg[1357]  ( .D(o[1357]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1357]) );
  DFF \round_reg_reg[1358]  ( .D(o[1358]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1358]) );
  DFF \round_reg_reg[1359]  ( .D(o[1359]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1359]) );
  DFF \round_reg_reg[1360]  ( .D(o[1360]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1360]) );
  DFF \round_reg_reg[1361]  ( .D(o[1361]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1361]) );
  DFF \round_reg_reg[1362]  ( .D(o[1362]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1362]) );
  DFF \round_reg_reg[1363]  ( .D(o[1363]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1363]) );
  DFF \round_reg_reg[1364]  ( .D(o[1364]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1364]) );
  DFF \round_reg_reg[1365]  ( .D(o[1365]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1365]) );
  DFF \round_reg_reg[1366]  ( .D(o[1366]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1366]) );
  DFF \round_reg_reg[1367]  ( .D(o[1367]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1367]) );
  DFF \round_reg_reg[1368]  ( .D(o[1368]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1368]) );
  DFF \round_reg_reg[1369]  ( .D(o[1369]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1369]) );
  DFF \round_reg_reg[1370]  ( .D(o[1370]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1370]) );
  DFF \round_reg_reg[1371]  ( .D(o[1371]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1371]) );
  DFF \round_reg_reg[1372]  ( .D(o[1372]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1372]) );
  DFF \round_reg_reg[1373]  ( .D(o[1373]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1373]) );
  DFF \round_reg_reg[1374]  ( .D(o[1374]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1374]) );
  DFF \round_reg_reg[1375]  ( .D(o[1375]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1375]) );
  DFF \round_reg_reg[1376]  ( .D(o[1376]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1376]) );
  DFF \round_reg_reg[1377]  ( .D(o[1377]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1377]) );
  DFF \round_reg_reg[1378]  ( .D(o[1378]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1378]) );
  DFF \round_reg_reg[1379]  ( .D(o[1379]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1379]) );
  DFF \round_reg_reg[1380]  ( .D(o[1380]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1380]) );
  DFF \round_reg_reg[1381]  ( .D(o[1381]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1381]) );
  DFF \round_reg_reg[1382]  ( .D(o[1382]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1382]) );
  DFF \round_reg_reg[1383]  ( .D(o[1383]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1383]) );
  DFF \round_reg_reg[1384]  ( .D(o[1384]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1384]) );
  DFF \round_reg_reg[1385]  ( .D(o[1385]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1385]) );
  DFF \round_reg_reg[1386]  ( .D(o[1386]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1386]) );
  DFF \round_reg_reg[1387]  ( .D(o[1387]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1387]) );
  DFF \round_reg_reg[1388]  ( .D(o[1388]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1388]) );
  DFF \round_reg_reg[1389]  ( .D(o[1389]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1389]) );
  DFF \round_reg_reg[1390]  ( .D(o[1390]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1390]) );
  DFF \round_reg_reg[1391]  ( .D(o[1391]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1391]) );
  DFF \round_reg_reg[1392]  ( .D(o[1392]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1392]) );
  DFF \round_reg_reg[1393]  ( .D(o[1393]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1393]) );
  DFF \round_reg_reg[1394]  ( .D(o[1394]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1394]) );
  DFF \round_reg_reg[1395]  ( .D(o[1395]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1395]) );
  DFF \round_reg_reg[1396]  ( .D(o[1396]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1396]) );
  DFF \round_reg_reg[1397]  ( .D(o[1397]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1397]) );
  DFF \round_reg_reg[1398]  ( .D(o[1398]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1398]) );
  DFF \round_reg_reg[1399]  ( .D(o[1399]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1399]) );
  DFF \round_reg_reg[1400]  ( .D(o[1400]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1400]) );
  DFF \round_reg_reg[1401]  ( .D(o[1401]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1401]) );
  DFF \round_reg_reg[1402]  ( .D(o[1402]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1402]) );
  DFF \round_reg_reg[1403]  ( .D(o[1403]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1403]) );
  DFF \round_reg_reg[1404]  ( .D(o[1404]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1404]) );
  DFF \round_reg_reg[1405]  ( .D(o[1405]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1405]) );
  DFF \round_reg_reg[1406]  ( .D(o[1406]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1406]) );
  DFF \round_reg_reg[1407]  ( .D(o[1407]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1407]) );
  DFF \round_reg_reg[1408]  ( .D(o[1408]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1408]) );
  DFF \round_reg_reg[1409]  ( .D(o[1409]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1409]) );
  DFF \round_reg_reg[1410]  ( .D(o[1410]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1410]) );
  DFF \round_reg_reg[1411]  ( .D(o[1411]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1411]) );
  DFF \round_reg_reg[1412]  ( .D(o[1412]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1412]) );
  DFF \round_reg_reg[1413]  ( .D(o[1413]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1413]) );
  DFF \round_reg_reg[1414]  ( .D(o[1414]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1414]) );
  DFF \round_reg_reg[1415]  ( .D(o[1415]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1415]) );
  DFF \round_reg_reg[1416]  ( .D(o[1416]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1416]) );
  DFF \round_reg_reg[1417]  ( .D(o[1417]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1417]) );
  DFF \round_reg_reg[1418]  ( .D(o[1418]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1418]) );
  DFF \round_reg_reg[1419]  ( .D(o[1419]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1419]) );
  DFF \round_reg_reg[1420]  ( .D(o[1420]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1420]) );
  DFF \round_reg_reg[1421]  ( .D(o[1421]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1421]) );
  DFF \round_reg_reg[1422]  ( .D(o[1422]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1422]) );
  DFF \round_reg_reg[1423]  ( .D(o[1423]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1423]) );
  DFF \round_reg_reg[1424]  ( .D(o[1424]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1424]) );
  DFF \round_reg_reg[1425]  ( .D(o[1425]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1425]) );
  DFF \round_reg_reg[1426]  ( .D(o[1426]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1426]) );
  DFF \round_reg_reg[1427]  ( .D(o[1427]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1427]) );
  DFF \round_reg_reg[1428]  ( .D(o[1428]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1428]) );
  DFF \round_reg_reg[1429]  ( .D(o[1429]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1429]) );
  DFF \round_reg_reg[1430]  ( .D(o[1430]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1430]) );
  DFF \round_reg_reg[1431]  ( .D(o[1431]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1431]) );
  DFF \round_reg_reg[1432]  ( .D(o[1432]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1432]) );
  DFF \round_reg_reg[1433]  ( .D(o[1433]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1433]) );
  DFF \round_reg_reg[1434]  ( .D(o[1434]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1434]) );
  DFF \round_reg_reg[1435]  ( .D(o[1435]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1435]) );
  DFF \round_reg_reg[1436]  ( .D(o[1436]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1436]) );
  DFF \round_reg_reg[1437]  ( .D(o[1437]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1437]) );
  DFF \round_reg_reg[1438]  ( .D(o[1438]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1438]) );
  DFF \round_reg_reg[1439]  ( .D(o[1439]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1439]) );
  DFF \round_reg_reg[1440]  ( .D(o[1440]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1440]) );
  DFF \round_reg_reg[1441]  ( .D(o[1441]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1441]) );
  DFF \round_reg_reg[1442]  ( .D(o[1442]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1442]) );
  DFF \round_reg_reg[1443]  ( .D(o[1443]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1443]) );
  DFF \round_reg_reg[1444]  ( .D(o[1444]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1444]) );
  DFF \round_reg_reg[1445]  ( .D(o[1445]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1445]) );
  DFF \round_reg_reg[1446]  ( .D(o[1446]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1446]) );
  DFF \round_reg_reg[1447]  ( .D(o[1447]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1447]) );
  DFF \round_reg_reg[1448]  ( .D(o[1448]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1448]) );
  DFF \round_reg_reg[1449]  ( .D(o[1449]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1449]) );
  DFF \round_reg_reg[1450]  ( .D(o[1450]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1450]) );
  DFF \round_reg_reg[1451]  ( .D(o[1451]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1451]) );
  DFF \round_reg_reg[1452]  ( .D(o[1452]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1452]) );
  DFF \round_reg_reg[1453]  ( .D(o[1453]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1453]) );
  DFF \round_reg_reg[1454]  ( .D(o[1454]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1454]) );
  DFF \round_reg_reg[1455]  ( .D(o[1455]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1455]) );
  DFF \round_reg_reg[1456]  ( .D(o[1456]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1456]) );
  DFF \round_reg_reg[1457]  ( .D(o[1457]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1457]) );
  DFF \round_reg_reg[1458]  ( .D(o[1458]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1458]) );
  DFF \round_reg_reg[1459]  ( .D(o[1459]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1459]) );
  DFF \round_reg_reg[1460]  ( .D(o[1460]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1460]) );
  DFF \round_reg_reg[1461]  ( .D(o[1461]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1461]) );
  DFF \round_reg_reg[1462]  ( .D(o[1462]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1462]) );
  DFF \round_reg_reg[1463]  ( .D(o[1463]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1463]) );
  DFF \round_reg_reg[1464]  ( .D(o[1464]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1464]) );
  DFF \round_reg_reg[1465]  ( .D(o[1465]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1465]) );
  DFF \round_reg_reg[1466]  ( .D(o[1466]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1466]) );
  DFF \round_reg_reg[1467]  ( .D(o[1467]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1467]) );
  DFF \round_reg_reg[1468]  ( .D(o[1468]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1468]) );
  DFF \round_reg_reg[1469]  ( .D(o[1469]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1469]) );
  DFF \round_reg_reg[1470]  ( .D(o[1470]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1470]) );
  DFF \round_reg_reg[1471]  ( .D(o[1471]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1471]) );
  DFF \round_reg_reg[1472]  ( .D(o[1472]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1472]) );
  DFF \round_reg_reg[1473]  ( .D(o[1473]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1473]) );
  DFF \round_reg_reg[1474]  ( .D(o[1474]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1474]) );
  DFF \round_reg_reg[1475]  ( .D(o[1475]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1475]) );
  DFF \round_reg_reg[1476]  ( .D(o[1476]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1476]) );
  DFF \round_reg_reg[1477]  ( .D(o[1477]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1477]) );
  DFF \round_reg_reg[1478]  ( .D(o[1478]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1478]) );
  DFF \round_reg_reg[1479]  ( .D(o[1479]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1479]) );
  DFF \round_reg_reg[1480]  ( .D(o[1480]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1480]) );
  DFF \round_reg_reg[1481]  ( .D(o[1481]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1481]) );
  DFF \round_reg_reg[1482]  ( .D(o[1482]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1482]) );
  DFF \round_reg_reg[1483]  ( .D(o[1483]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1483]) );
  DFF \round_reg_reg[1484]  ( .D(o[1484]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1484]) );
  DFF \round_reg_reg[1485]  ( .D(o[1485]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1485]) );
  DFF \round_reg_reg[1486]  ( .D(o[1486]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1486]) );
  DFF \round_reg_reg[1487]  ( .D(o[1487]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1487]) );
  DFF \round_reg_reg[1488]  ( .D(o[1488]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1488]) );
  DFF \round_reg_reg[1489]  ( .D(o[1489]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1489]) );
  DFF \round_reg_reg[1490]  ( .D(o[1490]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1490]) );
  DFF \round_reg_reg[1491]  ( .D(o[1491]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1491]) );
  DFF \round_reg_reg[1492]  ( .D(o[1492]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1492]) );
  DFF \round_reg_reg[1493]  ( .D(o[1493]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1493]) );
  DFF \round_reg_reg[1494]  ( .D(o[1494]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1494]) );
  DFF \round_reg_reg[1495]  ( .D(o[1495]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1495]) );
  DFF \round_reg_reg[1496]  ( .D(o[1496]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1496]) );
  DFF \round_reg_reg[1497]  ( .D(o[1497]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1497]) );
  DFF \round_reg_reg[1498]  ( .D(o[1498]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1498]) );
  DFF \round_reg_reg[1499]  ( .D(o[1499]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1499]) );
  DFF \round_reg_reg[1500]  ( .D(o[1500]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1500]) );
  DFF \round_reg_reg[1501]  ( .D(o[1501]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1501]) );
  DFF \round_reg_reg[1502]  ( .D(o[1502]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1502]) );
  DFF \round_reg_reg[1503]  ( .D(o[1503]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1503]) );
  DFF \round_reg_reg[1504]  ( .D(o[1504]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1504]) );
  DFF \round_reg_reg[1505]  ( .D(o[1505]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1505]) );
  DFF \round_reg_reg[1506]  ( .D(o[1506]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1506]) );
  DFF \round_reg_reg[1507]  ( .D(o[1507]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1507]) );
  DFF \round_reg_reg[1508]  ( .D(o[1508]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1508]) );
  DFF \round_reg_reg[1509]  ( .D(o[1509]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1509]) );
  DFF \round_reg_reg[1510]  ( .D(o[1510]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1510]) );
  DFF \round_reg_reg[1511]  ( .D(o[1511]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1511]) );
  DFF \round_reg_reg[1512]  ( .D(o[1512]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1512]) );
  DFF \round_reg_reg[1513]  ( .D(o[1513]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1513]) );
  DFF \round_reg_reg[1514]  ( .D(o[1514]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1514]) );
  DFF \round_reg_reg[1515]  ( .D(o[1515]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1515]) );
  DFF \round_reg_reg[1516]  ( .D(o[1516]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1516]) );
  DFF \round_reg_reg[1517]  ( .D(o[1517]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1517]) );
  DFF \round_reg_reg[1518]  ( .D(o[1518]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1518]) );
  DFF \round_reg_reg[1519]  ( .D(o[1519]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1519]) );
  DFF \round_reg_reg[1520]  ( .D(o[1520]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1520]) );
  DFF \round_reg_reg[1521]  ( .D(o[1521]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1521]) );
  DFF \round_reg_reg[1522]  ( .D(o[1522]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1522]) );
  DFF \round_reg_reg[1523]  ( .D(o[1523]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1523]) );
  DFF \round_reg_reg[1524]  ( .D(o[1524]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1524]) );
  DFF \round_reg_reg[1525]  ( .D(o[1525]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1525]) );
  DFF \round_reg_reg[1526]  ( .D(o[1526]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1526]) );
  DFF \round_reg_reg[1527]  ( .D(o[1527]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1527]) );
  DFF \round_reg_reg[1528]  ( .D(o[1528]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1528]) );
  DFF \round_reg_reg[1529]  ( .D(o[1529]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1529]) );
  DFF \round_reg_reg[1530]  ( .D(o[1530]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1530]) );
  DFF \round_reg_reg[1531]  ( .D(o[1531]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1531]) );
  DFF \round_reg_reg[1532]  ( .D(o[1532]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1532]) );
  DFF \round_reg_reg[1533]  ( .D(o[1533]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1533]) );
  DFF \round_reg_reg[1534]  ( .D(o[1534]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1534]) );
  DFF \round_reg_reg[1535]  ( .D(o[1535]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1535]) );
  DFF \round_reg_reg[1536]  ( .D(o[1536]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1536]) );
  DFF \round_reg_reg[1537]  ( .D(o[1537]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1537]) );
  DFF \round_reg_reg[1538]  ( .D(o[1538]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1538]) );
  DFF \round_reg_reg[1539]  ( .D(o[1539]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1539]) );
  DFF \round_reg_reg[1540]  ( .D(o[1540]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1540]) );
  DFF \round_reg_reg[1541]  ( .D(o[1541]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1541]) );
  DFF \round_reg_reg[1542]  ( .D(o[1542]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1542]) );
  DFF \round_reg_reg[1543]  ( .D(o[1543]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1543]) );
  DFF \round_reg_reg[1544]  ( .D(o[1544]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1544]) );
  DFF \round_reg_reg[1545]  ( .D(o[1545]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1545]) );
  DFF \round_reg_reg[1546]  ( .D(o[1546]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1546]) );
  DFF \round_reg_reg[1547]  ( .D(o[1547]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1547]) );
  DFF \round_reg_reg[1548]  ( .D(o[1548]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1548]) );
  DFF \round_reg_reg[1549]  ( .D(o[1549]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1549]) );
  DFF \round_reg_reg[1550]  ( .D(o[1550]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1550]) );
  DFF \round_reg_reg[1551]  ( .D(o[1551]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1551]) );
  DFF \round_reg_reg[1552]  ( .D(o[1552]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1552]) );
  DFF \round_reg_reg[1553]  ( .D(o[1553]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1553]) );
  DFF \round_reg_reg[1554]  ( .D(o[1554]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1554]) );
  DFF \round_reg_reg[1555]  ( .D(o[1555]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1555]) );
  DFF \round_reg_reg[1556]  ( .D(o[1556]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1556]) );
  DFF \round_reg_reg[1557]  ( .D(o[1557]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1557]) );
  DFF \round_reg_reg[1558]  ( .D(o[1558]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1558]) );
  DFF \round_reg_reg[1559]  ( .D(o[1559]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1559]) );
  DFF \round_reg_reg[1560]  ( .D(o[1560]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1560]) );
  DFF \round_reg_reg[1561]  ( .D(o[1561]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1561]) );
  DFF \round_reg_reg[1562]  ( .D(o[1562]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1562]) );
  DFF \round_reg_reg[1563]  ( .D(o[1563]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1563]) );
  DFF \round_reg_reg[1564]  ( .D(o[1564]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1564]) );
  DFF \round_reg_reg[1565]  ( .D(o[1565]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1565]) );
  DFF \round_reg_reg[1566]  ( .D(o[1566]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1566]) );
  DFF \round_reg_reg[1567]  ( .D(o[1567]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1567]) );
  DFF \round_reg_reg[1568]  ( .D(o[1568]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1568]) );
  DFF \round_reg_reg[1569]  ( .D(o[1569]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1569]) );
  DFF \round_reg_reg[1570]  ( .D(o[1570]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1570]) );
  DFF \round_reg_reg[1571]  ( .D(o[1571]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1571]) );
  DFF \round_reg_reg[1572]  ( .D(o[1572]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1572]) );
  DFF \round_reg_reg[1573]  ( .D(o[1573]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1573]) );
  DFF \round_reg_reg[1574]  ( .D(o[1574]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1574]) );
  DFF \round_reg_reg[1575]  ( .D(o[1575]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1575]) );
  DFF \round_reg_reg[1576]  ( .D(o[1576]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1576]) );
  DFF \round_reg_reg[1577]  ( .D(o[1577]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1577]) );
  DFF \round_reg_reg[1578]  ( .D(o[1578]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1578]) );
  DFF \round_reg_reg[1579]  ( .D(o[1579]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1579]) );
  DFF \round_reg_reg[1580]  ( .D(o[1580]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1580]) );
  DFF \round_reg_reg[1581]  ( .D(o[1581]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1581]) );
  DFF \round_reg_reg[1582]  ( .D(o[1582]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1582]) );
  DFF \round_reg_reg[1583]  ( .D(o[1583]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1583]) );
  DFF \round_reg_reg[1584]  ( .D(o[1584]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1584]) );
  DFF \round_reg_reg[1585]  ( .D(o[1585]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1585]) );
  DFF \round_reg_reg[1586]  ( .D(o[1586]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1586]) );
  DFF \round_reg_reg[1587]  ( .D(o[1587]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1587]) );
  DFF \round_reg_reg[1588]  ( .D(o[1588]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1588]) );
  DFF \round_reg_reg[1589]  ( .D(o[1589]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1589]) );
  DFF \round_reg_reg[1590]  ( .D(o[1590]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1590]) );
  DFF \round_reg_reg[1591]  ( .D(o[1591]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1591]) );
  DFF \round_reg_reg[1592]  ( .D(o[1592]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1592]) );
  DFF \round_reg_reg[1593]  ( .D(o[1593]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1593]) );
  DFF \round_reg_reg[1594]  ( .D(o[1594]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1594]) );
  DFF \round_reg_reg[1595]  ( .D(o[1595]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1595]) );
  DFF \round_reg_reg[1596]  ( .D(o[1596]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1596]) );
  DFF \round_reg_reg[1597]  ( .D(o[1597]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1597]) );
  DFF \round_reg_reg[1598]  ( .D(o[1598]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1598]) );
  DFF \round_reg_reg[1599]  ( .D(o[1599]), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        round_reg[1599]) );
  XNOR U1053 ( .A(n4796), .B(n4797), .Z(n4411) );
  XOR U1054 ( .A(n5784), .B(n4956), .Z(n1726) );
  XOR U1055 ( .A(n5708), .B(n4997), .Z(n1769) );
  XOR U1056 ( .A(n5723), .B(n5000), .Z(n1772) );
  XOR U1057 ( .A(n5738), .B(n5004), .Z(n1775) );
  ANDN U1058 ( .A(n3721), .B(n3722), .Z(n3719) );
  ANDN U1059 ( .A(n3738), .B(n3739), .Z(n3736) );
  ANDN U1060 ( .A(n3790), .B(n3791), .Z(n3788) );
  ANDN U1061 ( .A(n3798), .B(n3799), .Z(n3796) );
  ANDN U1062 ( .A(n3802), .B(n3803), .Z(n3800) );
  ANDN U1063 ( .A(n3806), .B(n3807), .Z(n3804) );
  ANDN U1064 ( .A(n3810), .B(n3811), .Z(n3808) );
  ANDN U1065 ( .A(n3814), .B(n3815), .Z(n3812) );
  ANDN U1066 ( .A(n3835), .B(n3836), .Z(n3833) );
  ANDN U1067 ( .A(n4133), .B(n3991), .Z(n4132) );
  NOR U1068 ( .A(n4131), .B(n3708), .Z(n4246) );
  NOR U1069 ( .A(n4135), .B(n3716), .Z(n4249) );
  ANDN U1070 ( .A(n1581), .B(n1338), .Z(n1580) );
  ANDN U1071 ( .A(n1583), .B(n1342), .Z(n1582) );
  ANDN U1072 ( .A(n1585), .B(n1346), .Z(n1584) );
  ANDN U1073 ( .A(n1591), .B(n1350), .Z(n1590) );
  XOR U1074 ( .A(n5693), .B(n4994), .Z(n1766) );
  ANDN U1075 ( .A(n3734), .B(n3735), .Z(n3732) );
  ANDN U1076 ( .A(n3786), .B(n3787), .Z(n3784) );
  ANDN U1077 ( .A(n3853), .B(n3854), .Z(n3851) );
  ANDN U1078 ( .A(n3857), .B(n3858), .Z(n3855) );
  ANDN U1079 ( .A(n3861), .B(n3862), .Z(n3859) );
  ANDN U1080 ( .A(n4009), .B(n3738), .Z(n4008) );
  NOR U1081 ( .A(n4097), .B(n3642), .Z(n4229) );
  NOR U1082 ( .A(n4103), .B(n3655), .Z(n4232) );
  NOR U1083 ( .A(n4106), .B(n3659), .Z(n4233) );
  NOR U1084 ( .A(n4108), .B(n3663), .Z(n4234) );
  NOR U1085 ( .A(n4110), .B(n3667), .Z(n4235) );
  NOR U1086 ( .A(n4124), .B(n3696), .Z(n4243) );
  NOR U1087 ( .A(n4127), .B(n3700), .Z(n4244) );
  NOR U1088 ( .A(n4129), .B(n3704), .Z(n4245) );
  NOR U1089 ( .A(n4133), .B(n3712), .Z(n4247) );
  ANDN U1090 ( .A(n1520), .B(n1238), .Z(n1519) );
  ANDN U1091 ( .A(n1522), .B(n1242), .Z(n1521) );
  ANDN U1092 ( .A(n1524), .B(n1246), .Z(n1523) );
  ANDN U1093 ( .A(n1579), .B(n1334), .Z(n1578) );
  ANDN U1094 ( .A(n1708), .B(n1518), .Z(n1707) );
  ANDN U1095 ( .A(n1792), .B(n1581), .Z(n1790) );
  ANDN U1096 ( .A(n1795), .B(n1583), .Z(n1793) );
  ANDN U1097 ( .A(n1798), .B(n1585), .Z(n1796) );
  ANDN U1098 ( .A(n1801), .B(n1591), .Z(n1799) );
  ANDN U1099 ( .A(n1813), .B(n1602), .Z(n1811) );
  ANDN U1100 ( .A(n1907), .B(n1692), .Z(n1905) );
  XOR U1101 ( .A(n5561), .B(n5562), .Z(n2253) );
  XOR U1102 ( .A(n5678), .B(n4991), .Z(n1763) );
  ANDN U1103 ( .A(n3765), .B(n3766), .Z(n3763) );
  ANDN U1104 ( .A(n3769), .B(n3770), .Z(n3767) );
  ANDN U1105 ( .A(n3781), .B(n3782), .Z(n3779) );
  ANDN U1106 ( .A(n3794), .B(n3795), .Z(n3792) );
  ANDN U1107 ( .A(n3646), .B(n4099), .Z(n4230) );
  ANDN U1108 ( .A(n4423), .B(n4424), .Z(n4421) );
  ANDN U1109 ( .A(n4427), .B(n4428), .Z(n4425) );
  ANDN U1110 ( .A(n1558), .B(n1298), .Z(n1557) );
  ANDN U1111 ( .A(n1566), .B(n1306), .Z(n1565) );
  ANDN U1112 ( .A(n1568), .B(n1310), .Z(n1567) );
  ANDN U1113 ( .A(n1570), .B(n1314), .Z(n1569) );
  ANDN U1114 ( .A(n1572), .B(n1318), .Z(n1571) );
  ANDN U1115 ( .A(n1577), .B(n1330), .Z(n1576) );
  ANDN U1116 ( .A(n1711), .B(n1520), .Z(n1709) );
  ANDN U1117 ( .A(n1714), .B(n1522), .Z(n1712) );
  ANDN U1118 ( .A(n1721), .B(n1524), .Z(n1719) );
  ANDN U1119 ( .A(n1779), .B(n1574), .Z(n1777) );
  ANDN U1120 ( .A(n1789), .B(n1579), .Z(n1787) );
  ANDN U1121 ( .A(n1804), .B(n1593), .Z(n1802) );
  ANDN U1122 ( .A(n1810), .B(n1599), .Z(n1808) );
  ANDN U1123 ( .A(n1816), .B(n1605), .Z(n1814) );
  ANDN U1124 ( .A(n1827), .B(n1608), .Z(n1825) );
  ANDN U1125 ( .A(n1830), .B(n1611), .Z(n1828) );
  ANDN U1126 ( .A(n1833), .B(n1614), .Z(n1831) );
  ANDN U1127 ( .A(n1836), .B(n1617), .Z(n1834) );
  ANDN U1128 ( .A(n1932), .B(n1708), .Z(n1930) );
  NOR U1129 ( .A(n1813), .B(n1368), .Z(n2015) );
  NOR U1130 ( .A(n1907), .B(n1480), .Z(n2085) );
  ANDN U1131 ( .A(n2862), .B(n2644), .Z(n2861) );
  ANDN U1132 ( .A(n3032), .B(n2868), .Z(n3031) );
  ANDN U1133 ( .A(n3034), .B(n2871), .Z(n3033) );
  ANDN U1134 ( .A(n3036), .B(n2874), .Z(n3035) );
  ANDN U1135 ( .A(n3038), .B(n2877), .Z(n3037) );
  XNOR U1136 ( .A(n4792), .B(n4793), .Z(n4409) );
  XNOR U1137 ( .A(n4800), .B(n4801), .Z(n4413) );
  XNOR U1138 ( .A(n4804), .B(n4805), .Z(n4415) );
  XOR U1139 ( .A(n5773), .B(n4909), .Z(n2172) );
  XOR U1140 ( .A(n5359), .B(n4917), .Z(n1912) );
  XOR U1141 ( .A(n5419), .B(n4933), .Z(n1928) );
  XOR U1142 ( .A(n5432), .B(n4939), .Z(n1931) );
  XOR U1143 ( .A(n5675), .B(n4953), .Z(n1723) );
  XOR U1144 ( .A(n5799), .B(n4959), .Z(n1729) );
  XOR U1145 ( .A(n5622), .B(n4982), .Z(n1754) );
  XOR U1146 ( .A(n5637), .B(n4985), .Z(n1757) );
  XOR U1147 ( .A(n5652), .B(n4988), .Z(n1760) );
  ANDN U1148 ( .A(n3652), .B(n3653), .Z(n3650) );
  ANDN U1149 ( .A(n3701), .B(n3702), .Z(n3699) );
  ANDN U1150 ( .A(n3705), .B(n3706), .Z(n3703) );
  ANDN U1151 ( .A(n3713), .B(n3714), .Z(n3711) );
  ANDN U1152 ( .A(n3744), .B(n3745), .Z(n3743) );
  ANDN U1153 ( .A(n3757), .B(n3758), .Z(n3755) );
  ANDN U1154 ( .A(n3881), .B(n3882), .Z(n3879) );
  ANDN U1155 ( .A(n3889), .B(n3890), .Z(n3887) );
  ANDN U1156 ( .A(n3896), .B(n3897), .Z(n3895) );
  ANDN U1157 ( .A(n3911), .B(n3912), .Z(n3909) );
  ANDN U1158 ( .A(n3930), .B(n3931), .Z(n3929) );
  ANDN U1159 ( .A(n1560), .B(n1302), .Z(n1559) );
  ANDN U1160 ( .A(n1767), .B(n1566), .Z(n1765) );
  ANDN U1161 ( .A(n1770), .B(n1568), .Z(n1768) );
  ANDN U1162 ( .A(n1773), .B(n1570), .Z(n1771) );
  ANDN U1163 ( .A(n1776), .B(n1572), .Z(n1774) );
  ANDN U1164 ( .A(n1782), .B(n1577), .Z(n1780) );
  ANDN U1165 ( .A(n1236), .B(n1711), .Z(n1933) );
  NOR U1166 ( .A(n1779), .B(n1324), .Z(n1992) );
  NOR U1167 ( .A(n1789), .B(n1332), .Z(n1996) );
  NOR U1168 ( .A(n1792), .B(n1336), .Z(n1998) );
  NOR U1169 ( .A(n1795), .B(n1340), .Z(n2000) );
  NOR U1170 ( .A(n1798), .B(n1344), .Z(n2002) );
  NOR U1171 ( .A(n1801), .B(n1348), .Z(n2004) );
  NOR U1172 ( .A(n1804), .B(n1352), .Z(n2006) );
  NOR U1173 ( .A(n1807), .B(n1356), .Z(n2011) );
  NOR U1174 ( .A(n1810), .B(n1360), .Z(n2013) );
  NOR U1175 ( .A(n1816), .B(n1372), .Z(n2017) );
  NOR U1176 ( .A(n1827), .B(n1376), .Z(n2019) );
  NOR U1177 ( .A(n1830), .B(n1380), .Z(n2021) );
  NOR U1178 ( .A(n1833), .B(n1384), .Z(n2023) );
  NOR U1179 ( .A(n1836), .B(n1388), .Z(n2025) );
  ANDN U1180 ( .A(n3030), .B(n2862), .Z(n3028) );
  NOR U1181 ( .A(n2985), .B(n2559), .Z(n3123) );
  NOR U1182 ( .A(n3032), .B(n2646), .Z(n3168) );
  NOR U1183 ( .A(n3034), .B(n2650), .Z(n3169) );
  NOR U1184 ( .A(n3036), .B(n2654), .Z(n3174) );
  NOR U1185 ( .A(n3038), .B(n2658), .Z(n3175) );
  ANDN U1186 ( .A(n3456), .B(n3457), .Z(n3454) );
  XNOR U1187 ( .A(n5069), .B(n5010), .Z(n4248) );
  XOR U1188 ( .A(n5788), .B(n4913), .Z(n2180) );
  XOR U1189 ( .A(n5381), .B(n4921), .Z(n1915) );
  XOR U1190 ( .A(n5392), .B(n4925), .Z(n1918) );
  XOR U1191 ( .A(n5406), .B(n4929), .Z(n1921) );
  XOR U1192 ( .A(n5445), .B(n4943), .Z(n1710) );
  XOR U1193 ( .A(n5458), .B(n4947), .Z(n1713) );
  XOR U1194 ( .A(n5516), .B(n4950), .Z(n1720) );
  ANDN U1195 ( .A(n3647), .B(n3648), .Z(n3645) );
  ANDN U1196 ( .A(n3656), .B(n3657), .Z(n3654) );
  ANDN U1197 ( .A(n3660), .B(n3661), .Z(n3658) );
  ANDN U1198 ( .A(n3672), .B(n3673), .Z(n3670) );
  ANDN U1199 ( .A(n3709), .B(n3710), .Z(n3707) );
  ANDN U1200 ( .A(n3717), .B(n3718), .Z(n3715) );
  ANDN U1201 ( .A(n3725), .B(n3726), .Z(n3723) );
  ANDN U1202 ( .A(n3729), .B(n3730), .Z(n3727) );
  ANDN U1203 ( .A(n3761), .B(n3762), .Z(n3759) );
  ANDN U1204 ( .A(n3773), .B(n3774), .Z(n3771) );
  ANDN U1205 ( .A(n3777), .B(n3778), .Z(n3775) );
  ANDN U1206 ( .A(n3820), .B(n3821), .Z(n3819) );
  ANDN U1207 ( .A(n3840), .B(n3841), .Z(n3838) );
  ANDN U1208 ( .A(n3849), .B(n3850), .Z(n3847) );
  ANDN U1209 ( .A(n3867), .B(n3868), .Z(n3866) );
  ANDN U1210 ( .A(n3885), .B(n3886), .Z(n3883) );
  ANDN U1211 ( .A(n3917), .B(n3918), .Z(n3916) );
  NOR U1212 ( .A(n4101), .B(n3651), .Z(n4231) );
  ANDN U1213 ( .A(n1526), .B(n1250), .Z(n1525) );
  ANDN U1214 ( .A(n1528), .B(n1254), .Z(n1527) );
  ANDN U1215 ( .A(n1530), .B(n1258), .Z(n1529) );
  ANDN U1216 ( .A(n1556), .B(n1294), .Z(n1555) );
  ANDN U1217 ( .A(n1706), .B(n1514), .Z(n1705) );
  ANDN U1218 ( .A(n1761), .B(n1558), .Z(n1759) );
  ANDN U1219 ( .A(n1764), .B(n1560), .Z(n1762) );
  ANDN U1220 ( .A(n1807), .B(n1596), .Z(n1805) );
  ANDN U1221 ( .A(n1240), .B(n1714), .Z(n1935) );
  ANDN U1222 ( .A(n1244), .B(n1721), .Z(n1937) );
  NOR U1223 ( .A(n1782), .B(n1328), .Z(n1994) );
  NOR U1224 ( .A(n1932), .B(n1516), .Z(n2109) );
  ANDN U1225 ( .A(n2753), .B(n2493), .Z(n2752) );
  ANDN U1226 ( .A(n2757), .B(n2501), .Z(n2756) );
  ANDN U1227 ( .A(n2759), .B(n2505), .Z(n2758) );
  ANDN U1228 ( .A(n2761), .B(n2509), .Z(n2760) );
  NOR U1229 ( .A(n2961), .B(n2515), .Z(n3101) );
  NOR U1230 ( .A(n2975), .B(n2539), .Z(n3114) );
  NOR U1231 ( .A(n3005), .B(n2598), .Z(n3142) );
  NOR U1232 ( .A(n3030), .B(n2642), .Z(n3167) );
  XNOR U1233 ( .A(n3419), .B(n1891), .Z(o[269]) );
  XNOR U1234 ( .A(n3422), .B(n1925), .Z(o[268]) );
  XNOR U1235 ( .A(n3425), .B(n1956), .Z(o[267]) );
  XNOR U1236 ( .A(n3428), .B(n1986), .Z(o[266]) );
  ANDN U1237 ( .A(n3440), .B(n2128), .Z(n3439) );
  ANDN U1238 ( .A(n3442), .B(n2571), .Z(n3441) );
  ANDN U1239 ( .A(n3444), .B(n2920), .Z(n3443) );
  ANDN U1240 ( .A(n3447), .B(n3148), .Z(n3446) );
  ANDN U1241 ( .A(n3452), .B(n3453), .Z(n3450) );
  ANDN U1242 ( .A(n3459), .B(n3263), .Z(n3458) );
  ANDN U1243 ( .A(n3461), .B(n3266), .Z(n3460) );
  ANDN U1244 ( .A(n3463), .B(n3269), .Z(n3462) );
  ANDN U1245 ( .A(n3465), .B(n3272), .Z(n3464) );
  ANDN U1246 ( .A(n3467), .B(n3275), .Z(n3466) );
  NOR U1247 ( .A(n3456), .B(n2351), .Z(n3559) );
  NOR U1248 ( .A(n3507), .B(n3125), .Z(n3587) );
  NOR U1249 ( .A(n3509), .B(n3151), .Z(n3588) );
  NOR U1250 ( .A(n3511), .B(n3171), .Z(n3589) );
  NOR U1251 ( .A(n3514), .B(n3185), .Z(n3590) );
  NOR U1252 ( .A(n3516), .B(n3199), .Z(n3591) );
  XOR U1253 ( .A(n4761), .B(n4762), .Z(n2086) );
  XOR U1254 ( .A(n5546), .B(n5547), .Z(n2249) );
  XOR U1255 ( .A(n4948), .B(n5277), .Z(n2212) );
  XOR U1256 ( .A(n5576), .B(n5577), .Z(n2257) );
  XOR U1257 ( .A(n5591), .B(n5592), .Z(n2261) );
  XOR U1258 ( .A(n5606), .B(n5607), .Z(n2269) );
  ANDN U1259 ( .A(n3602), .B(n3603), .Z(n3601) );
  ANDN U1260 ( .A(n3615), .B(n3616), .Z(n3613) );
  ANDN U1261 ( .A(n3619), .B(n3620), .Z(n3617) );
  ANDN U1262 ( .A(n3623), .B(n3624), .Z(n3621) );
  ANDN U1263 ( .A(n3627), .B(n3628), .Z(n3625) );
  ANDN U1264 ( .A(n3631), .B(n3632), .Z(n3629) );
  ANDN U1265 ( .A(n3635), .B(n3636), .Z(n3633) );
  ANDN U1266 ( .A(n3639), .B(n3640), .Z(n3637) );
  ANDN U1267 ( .A(n3643), .B(n3644), .Z(n3641) );
  ANDN U1268 ( .A(n3664), .B(n3665), .Z(n3662) );
  ANDN U1269 ( .A(n3668), .B(n3669), .Z(n3666) );
  ANDN U1270 ( .A(n3676), .B(n3677), .Z(n3674) );
  ANDN U1271 ( .A(n3680), .B(n3681), .Z(n3678) );
  ANDN U1272 ( .A(n3684), .B(n3685), .Z(n3682) );
  ANDN U1273 ( .A(n3688), .B(n3689), .Z(n3686) );
  ANDN U1274 ( .A(n3693), .B(n3694), .Z(n3691) );
  NOR U1275 ( .A(n4112), .B(n3671), .Z(n4236) );
  ANDN U1276 ( .A(n1554), .B(n1290), .Z(n1553) );
  ANDN U1277 ( .A(n1698), .B(n1490), .Z(n1697) );
  ANDN U1278 ( .A(n1700), .B(n1494), .Z(n1699) );
  ANDN U1279 ( .A(n1702), .B(n1506), .Z(n1701) );
  ANDN U1280 ( .A(n1704), .B(n1510), .Z(n1703) );
  ANDN U1281 ( .A(n2755), .B(n2497), .Z(n2754) );
  ANDN U1282 ( .A(n2904), .B(n2694), .Z(n2903) );
  ANDN U1283 ( .A(n2906), .B(n2697), .Z(n2905) );
  ANDN U1284 ( .A(n3363), .B(n3364), .Z(n3361) );
  ANDN U1285 ( .A(n3367), .B(n3368), .Z(n3365) );
  ANDN U1286 ( .A(n3371), .B(n3372), .Z(n3369) );
  ANDN U1287 ( .A(n3375), .B(n3376), .Z(n3373) );
  NOR U1288 ( .A(n3354), .B(n1232), .Z(n3521) );
  NOR U1289 ( .A(n3356), .B(n1276), .Z(n3522) );
  NOR U1290 ( .A(n3358), .B(n1320), .Z(n3523) );
  NOR U1291 ( .A(n3360), .B(n1364), .Z(n3524) );
  NOR U1292 ( .A(n3409), .B(n1784), .Z(n3540) );
  NOR U1293 ( .A(n3413), .B(n1822), .Z(n3541) );
  NOR U1294 ( .A(n3417), .B(n1856), .Z(n3542) );
  NOR U1295 ( .A(n3421), .B(n1890), .Z(n3543) );
  NOR U1296 ( .A(n3424), .B(n1924), .Z(n3544) );
  NOR U1297 ( .A(n3427), .B(n1955), .Z(n3545) );
  NOR U1298 ( .A(n3430), .B(n1985), .Z(n3546) );
  NOR U1299 ( .A(n3434), .B(n2034), .Z(n3549) );
  NOR U1300 ( .A(n3437), .B(n2065), .Z(n3552) );
  NOR U1301 ( .A(n3440), .B(n2091), .Z(n3553) );
  NOR U1302 ( .A(n3442), .B(n2131), .Z(n3554) );
  NOR U1303 ( .A(n3444), .B(n2175), .Z(n3555) );
  NOR U1304 ( .A(n3447), .B(n2219), .Z(n3556) );
  NOR U1305 ( .A(n3449), .B(n2263), .Z(n3557) );
  NOR U1306 ( .A(n3452), .B(n2307), .Z(n3558) );
  NOR U1307 ( .A(n3459), .B(n2395), .Z(n3560) );
  NOR U1308 ( .A(n3461), .B(n2439), .Z(n3561) );
  NOR U1309 ( .A(n3463), .B(n2483), .Z(n3563) );
  NOR U1310 ( .A(n3465), .B(n2527), .Z(n3564) );
  NOR U1311 ( .A(n3467), .B(n2574), .Z(n3565) );
  NOR U1312 ( .A(n3469), .B(n2618), .Z(n3566) );
  NOR U1313 ( .A(n3472), .B(n2662), .Z(n3567) );
  NOR U1314 ( .A(n3474), .B(n2700), .Z(n3568) );
  NOR U1315 ( .A(n3476), .B(n2734), .Z(n3569) );
  NOR U1316 ( .A(n3478), .B(n2763), .Z(n3570) );
  NOR U1317 ( .A(n3480), .B(n2797), .Z(n3571) );
  NOR U1318 ( .A(n3482), .B(n2831), .Z(n3572) );
  NOR U1319 ( .A(n3484), .B(n2864), .Z(n3574) );
  NOR U1320 ( .A(n3486), .B(n2896), .Z(n3575) );
  NOR U1321 ( .A(n3488), .B(n2923), .Z(n3576) );
  NOR U1322 ( .A(n3490), .B(n2947), .Z(n3577) );
  NOR U1323 ( .A(n3493), .B(n2971), .Z(n3578) );
  NOR U1324 ( .A(n3497), .B(n3019), .Z(n3581) );
  NOR U1325 ( .A(n3499), .B(n3044), .Z(n3582) );
  NOR U1326 ( .A(n3501), .B(n3060), .Z(n3583) );
  NOR U1327 ( .A(n3503), .B(n3080), .Z(n3584) );
  NOR U1328 ( .A(n3505), .B(n3103), .Z(n3586) );
  ANDN U1329 ( .A(n2352), .B(n2353), .Z(n2350) );
  ANDN U1330 ( .A(n3126), .B(n3127), .Z(n3124) );
  ANDN U1331 ( .A(n3152), .B(n3153), .Z(n3150) );
  ANDN U1332 ( .A(n3172), .B(n3173), .Z(n3170) );
  ANDN U1333 ( .A(n3186), .B(n3187), .Z(n3184) );
  ANDN U1334 ( .A(n3200), .B(n3201), .Z(n3198) );
  XOR U1335 ( .A(n1051), .B(n1052), .Z(o[9]) );
  ANDN U1336 ( .A(n1053), .B(n1054), .Z(n1051) );
  XOR U1337 ( .A(n1055), .B(n1056), .Z(o[99]) );
  ANDN U1338 ( .A(n1057), .B(n1058), .Z(n1055) );
  XOR U1339 ( .A(n1059), .B(n1060), .Z(o[999]) );
  ANDN U1340 ( .A(n1061), .B(n1062), .Z(n1059) );
  XOR U1341 ( .A(n1063), .B(n1064), .Z(o[998]) );
  AND U1342 ( .A(n1065), .B(n1066), .Z(n1063) );
  XOR U1343 ( .A(n1067), .B(n1068), .Z(o[997]) );
  ANDN U1344 ( .A(n1069), .B(n1070), .Z(n1067) );
  XOR U1345 ( .A(n1071), .B(n1072), .Z(o[996]) );
  ANDN U1346 ( .A(n1073), .B(n1074), .Z(n1071) );
  XOR U1347 ( .A(n1075), .B(n1076), .Z(o[995]) );
  ANDN U1348 ( .A(n1077), .B(n1078), .Z(n1075) );
  XOR U1349 ( .A(n1079), .B(n1080), .Z(o[994]) );
  ANDN U1350 ( .A(n1081), .B(n1082), .Z(n1079) );
  XOR U1351 ( .A(n1083), .B(n1084), .Z(o[993]) );
  ANDN U1352 ( .A(n1085), .B(n1086), .Z(n1083) );
  XOR U1353 ( .A(n1087), .B(n1088), .Z(o[992]) );
  ANDN U1354 ( .A(n1089), .B(n1090), .Z(n1087) );
  XOR U1355 ( .A(n1091), .B(n1092), .Z(o[991]) );
  ANDN U1356 ( .A(n1093), .B(n1094), .Z(n1091) );
  XOR U1357 ( .A(n1095), .B(n1096), .Z(o[990]) );
  ANDN U1358 ( .A(n1097), .B(n1098), .Z(n1095) );
  XOR U1359 ( .A(n1099), .B(n1100), .Z(o[98]) );
  ANDN U1360 ( .A(n1101), .B(n1102), .Z(n1099) );
  XNOR U1361 ( .A(n1103), .B(n1104), .Z(o[989]) );
  ANDN U1362 ( .A(n1105), .B(n1106), .Z(n1103) );
  XNOR U1363 ( .A(n1107), .B(n1108), .Z(o[988]) );
  ANDN U1364 ( .A(n1109), .B(n1110), .Z(n1107) );
  XOR U1365 ( .A(n1111), .B(n1112), .Z(o[987]) );
  ANDN U1366 ( .A(n1113), .B(n1114), .Z(n1111) );
  XOR U1367 ( .A(n1115), .B(n1116), .Z(o[986]) );
  ANDN U1368 ( .A(n1117), .B(n1118), .Z(n1115) );
  XOR U1369 ( .A(n1119), .B(n1120), .Z(o[985]) );
  ANDN U1370 ( .A(n1121), .B(n1122), .Z(n1119) );
  XOR U1371 ( .A(n1123), .B(n1124), .Z(o[984]) );
  ANDN U1372 ( .A(n1125), .B(n1126), .Z(n1123) );
  XOR U1373 ( .A(n1127), .B(n1128), .Z(o[983]) );
  ANDN U1374 ( .A(n1129), .B(n1130), .Z(n1127) );
  XOR U1375 ( .A(n1131), .B(n1132), .Z(o[982]) );
  ANDN U1376 ( .A(n1133), .B(n1134), .Z(n1131) );
  XOR U1377 ( .A(n1135), .B(n1136), .Z(o[981]) );
  ANDN U1378 ( .A(n1137), .B(n1138), .Z(n1135) );
  XOR U1379 ( .A(n1139), .B(n1140), .Z(o[980]) );
  ANDN U1380 ( .A(n1141), .B(n1142), .Z(n1139) );
  XOR U1381 ( .A(n1143), .B(n1144), .Z(o[97]) );
  AND U1382 ( .A(n1145), .B(n1146), .Z(n1143) );
  XOR U1383 ( .A(n1147), .B(n1148), .Z(o[979]) );
  NOR U1384 ( .A(n1149), .B(n1150), .Z(n1147) );
  XOR U1385 ( .A(n1151), .B(n1152), .Z(o[978]) );
  ANDN U1386 ( .A(n1153), .B(n1154), .Z(n1151) );
  XOR U1387 ( .A(n1155), .B(n1156), .Z(o[977]) );
  ANDN U1388 ( .A(n1157), .B(n1158), .Z(n1155) );
  XOR U1389 ( .A(n1159), .B(n1160), .Z(o[976]) );
  ANDN U1390 ( .A(n1161), .B(n1162), .Z(n1159) );
  XNOR U1391 ( .A(n1163), .B(n1164), .Z(o[975]) );
  ANDN U1392 ( .A(n1165), .B(n1166), .Z(n1163) );
  XOR U1393 ( .A(n1167), .B(n1168), .Z(o[974]) );
  ANDN U1394 ( .A(n1169), .B(n1170), .Z(n1167) );
  XOR U1395 ( .A(n1171), .B(n1172), .Z(o[973]) );
  ANDN U1396 ( .A(n1173), .B(n1174), .Z(n1171) );
  XOR U1397 ( .A(n1175), .B(n1176), .Z(o[972]) );
  NOR U1398 ( .A(n1177), .B(n1178), .Z(n1175) );
  XOR U1399 ( .A(n1179), .B(n1180), .Z(o[971]) );
  NOR U1400 ( .A(n1181), .B(n1182), .Z(n1179) );
  XOR U1401 ( .A(n1183), .B(n1184), .Z(o[970]) );
  NOR U1402 ( .A(n1185), .B(n1186), .Z(n1183) );
  XNOR U1403 ( .A(n1187), .B(n1188), .Z(o[96]) );
  AND U1404 ( .A(n1189), .B(n1190), .Z(n1187) );
  XOR U1405 ( .A(n1191), .B(n1192), .Z(o[969]) );
  NOR U1406 ( .A(n1193), .B(n1194), .Z(n1191) );
  XNOR U1407 ( .A(n1195), .B(n1196), .Z(o[968]) );
  ANDN U1408 ( .A(n1197), .B(n1198), .Z(n1195) );
  XNOR U1409 ( .A(n1199), .B(n1200), .Z(o[967]) );
  ANDN U1410 ( .A(n1201), .B(n1202), .Z(n1199) );
  XNOR U1411 ( .A(n1203), .B(n1204), .Z(o[966]) );
  ANDN U1412 ( .A(n1205), .B(n1206), .Z(n1203) );
  XNOR U1413 ( .A(n1207), .B(n1208), .Z(o[965]) );
  AND U1414 ( .A(n1209), .B(n1210), .Z(n1207) );
  XNOR U1415 ( .A(n1211), .B(n1212), .Z(o[964]) );
  AND U1416 ( .A(n1213), .B(n1214), .Z(n1211) );
  XNOR U1417 ( .A(n1215), .B(n1216), .Z(o[963]) );
  AND U1418 ( .A(n1217), .B(n1218), .Z(n1215) );
  XNOR U1419 ( .A(n1219), .B(n1220), .Z(o[962]) );
  AND U1420 ( .A(n1221), .B(n1222), .Z(n1219) );
  XNOR U1421 ( .A(n1223), .B(n1224), .Z(o[961]) );
  AND U1422 ( .A(n1225), .B(n1226), .Z(n1223) );
  XNOR U1423 ( .A(n1227), .B(n1228), .Z(o[960]) );
  AND U1424 ( .A(n1229), .B(n1230), .Z(n1227) );
  XNOR U1425 ( .A(n1231), .B(n1232), .Z(o[95]) );
  AND U1426 ( .A(n1233), .B(n1234), .Z(n1231) );
  XOR U1427 ( .A(n1235), .B(n1236), .Z(o[959]) );
  AND U1428 ( .A(n1237), .B(n1238), .Z(n1235) );
  XOR U1429 ( .A(n1239), .B(n1240), .Z(o[958]) );
  AND U1430 ( .A(n1241), .B(n1242), .Z(n1239) );
  XOR U1431 ( .A(n1243), .B(n1244), .Z(o[957]) );
  AND U1432 ( .A(n1245), .B(n1246), .Z(n1243) );
  XOR U1433 ( .A(n1247), .B(n1248), .Z(o[956]) );
  AND U1434 ( .A(n1249), .B(n1250), .Z(n1247) );
  XOR U1435 ( .A(n1251), .B(n1252), .Z(o[955]) );
  AND U1436 ( .A(n1253), .B(n1254), .Z(n1251) );
  XNOR U1437 ( .A(n1255), .B(n1256), .Z(o[954]) );
  AND U1438 ( .A(n1257), .B(n1258), .Z(n1255) );
  XNOR U1439 ( .A(n1259), .B(n1260), .Z(o[953]) );
  AND U1440 ( .A(n1261), .B(n1262), .Z(n1259) );
  XNOR U1441 ( .A(n1263), .B(n1264), .Z(o[952]) );
  AND U1442 ( .A(n1265), .B(n1266), .Z(n1263) );
  XNOR U1443 ( .A(n1267), .B(n1268), .Z(o[951]) );
  AND U1444 ( .A(n1269), .B(n1270), .Z(n1267) );
  XNOR U1445 ( .A(n1271), .B(n1272), .Z(o[950]) );
  AND U1446 ( .A(n1273), .B(n1274), .Z(n1271) );
  XNOR U1447 ( .A(n1275), .B(n1276), .Z(o[94]) );
  AND U1448 ( .A(n1277), .B(n1278), .Z(n1275) );
  XNOR U1449 ( .A(n1279), .B(n1280), .Z(o[949]) );
  AND U1450 ( .A(n1281), .B(n1282), .Z(n1279) );
  XNOR U1451 ( .A(n1283), .B(n1284), .Z(o[948]) );
  AND U1452 ( .A(n1285), .B(n1286), .Z(n1283) );
  XNOR U1453 ( .A(n1287), .B(n1288), .Z(o[947]) );
  AND U1454 ( .A(n1289), .B(n1290), .Z(n1287) );
  XNOR U1455 ( .A(n1291), .B(n1292), .Z(o[946]) );
  AND U1456 ( .A(n1293), .B(n1294), .Z(n1291) );
  XNOR U1457 ( .A(n1295), .B(n1296), .Z(o[945]) );
  AND U1458 ( .A(n1297), .B(n1298), .Z(n1295) );
  XNOR U1459 ( .A(n1299), .B(n1300), .Z(o[944]) );
  AND U1460 ( .A(n1301), .B(n1302), .Z(n1299) );
  XNOR U1461 ( .A(n1303), .B(n1304), .Z(o[943]) );
  AND U1462 ( .A(n1305), .B(n1306), .Z(n1303) );
  XNOR U1463 ( .A(n1307), .B(n1308), .Z(o[942]) );
  AND U1464 ( .A(n1309), .B(n1310), .Z(n1307) );
  XNOR U1465 ( .A(n1311), .B(n1312), .Z(o[941]) );
  AND U1466 ( .A(n1313), .B(n1314), .Z(n1311) );
  XNOR U1467 ( .A(n1315), .B(n1316), .Z(o[940]) );
  AND U1468 ( .A(n1317), .B(n1318), .Z(n1315) );
  XNOR U1469 ( .A(n1319), .B(n1320), .Z(o[93]) );
  AND U1470 ( .A(n1321), .B(n1322), .Z(n1319) );
  XNOR U1471 ( .A(n1323), .B(n1324), .Z(o[939]) );
  AND U1472 ( .A(n1325), .B(n1326), .Z(n1323) );
  XNOR U1473 ( .A(n1327), .B(n1328), .Z(o[938]) );
  AND U1474 ( .A(n1329), .B(n1330), .Z(n1327) );
  XNOR U1475 ( .A(n1331), .B(n1332), .Z(o[937]) );
  AND U1476 ( .A(n1333), .B(n1334), .Z(n1331) );
  XNOR U1477 ( .A(n1335), .B(n1336), .Z(o[936]) );
  AND U1478 ( .A(n1337), .B(n1338), .Z(n1335) );
  XNOR U1479 ( .A(n1339), .B(n1340), .Z(o[935]) );
  AND U1480 ( .A(n1341), .B(n1342), .Z(n1339) );
  XNOR U1481 ( .A(n1343), .B(n1344), .Z(o[934]) );
  AND U1482 ( .A(n1345), .B(n1346), .Z(n1343) );
  XNOR U1483 ( .A(n1347), .B(n1348), .Z(o[933]) );
  AND U1484 ( .A(n1349), .B(n1350), .Z(n1347) );
  XNOR U1485 ( .A(n1351), .B(n1352), .Z(o[932]) );
  AND U1486 ( .A(n1353), .B(n1354), .Z(n1351) );
  XNOR U1487 ( .A(n1355), .B(n1356), .Z(o[931]) );
  AND U1488 ( .A(n1357), .B(n1358), .Z(n1355) );
  XNOR U1489 ( .A(n1359), .B(n1360), .Z(o[930]) );
  AND U1490 ( .A(n1361), .B(n1362), .Z(n1359) );
  XNOR U1491 ( .A(n1363), .B(n1364), .Z(o[92]) );
  AND U1492 ( .A(n1365), .B(n1366), .Z(n1363) );
  XNOR U1493 ( .A(n1367), .B(n1368), .Z(o[929]) );
  AND U1494 ( .A(n1369), .B(n1370), .Z(n1367) );
  XNOR U1495 ( .A(n1371), .B(n1372), .Z(o[928]) );
  AND U1496 ( .A(n1373), .B(n1374), .Z(n1371) );
  XNOR U1497 ( .A(n1375), .B(n1376), .Z(o[927]) );
  AND U1498 ( .A(n1377), .B(n1378), .Z(n1375) );
  XNOR U1499 ( .A(n1379), .B(n1380), .Z(o[926]) );
  AND U1500 ( .A(n1381), .B(n1382), .Z(n1379) );
  XNOR U1501 ( .A(n1383), .B(n1384), .Z(o[925]) );
  AND U1502 ( .A(n1385), .B(n1386), .Z(n1383) );
  XNOR U1503 ( .A(n1387), .B(n1388), .Z(o[924]) );
  AND U1504 ( .A(n1389), .B(n1390), .Z(n1387) );
  XNOR U1505 ( .A(n1391), .B(n1392), .Z(o[923]) );
  AND U1506 ( .A(n1393), .B(n1394), .Z(n1391) );
  XNOR U1507 ( .A(n1395), .B(n1396), .Z(o[922]) );
  AND U1508 ( .A(n1397), .B(n1398), .Z(n1395) );
  XNOR U1509 ( .A(n1399), .B(n1400), .Z(o[921]) );
  AND U1510 ( .A(n1401), .B(n1402), .Z(n1399) );
  XNOR U1511 ( .A(n1403), .B(n1404), .Z(o[920]) );
  AND U1512 ( .A(n1405), .B(n1406), .Z(n1403) );
  XNOR U1513 ( .A(n1407), .B(n1408), .Z(o[91]) );
  AND U1514 ( .A(n1409), .B(n1410), .Z(n1407) );
  XNOR U1515 ( .A(n1411), .B(n1412), .Z(o[919]) );
  AND U1516 ( .A(n1413), .B(n1414), .Z(n1411) );
  XNOR U1517 ( .A(n1415), .B(n1416), .Z(o[918]) );
  AND U1518 ( .A(n1417), .B(n1418), .Z(n1415) );
  XNOR U1519 ( .A(n1419), .B(n1420), .Z(o[917]) );
  AND U1520 ( .A(n1421), .B(n1422), .Z(n1419) );
  XNOR U1521 ( .A(n1423), .B(n1424), .Z(o[916]) );
  AND U1522 ( .A(n1425), .B(n1426), .Z(n1423) );
  XNOR U1523 ( .A(n1427), .B(n1428), .Z(o[915]) );
  AND U1524 ( .A(n1429), .B(n1430), .Z(n1427) );
  XNOR U1525 ( .A(n1431), .B(n1432), .Z(o[914]) );
  AND U1526 ( .A(n1433), .B(n1434), .Z(n1431) );
  XNOR U1527 ( .A(n1435), .B(n1436), .Z(o[913]) );
  AND U1528 ( .A(n1437), .B(n1438), .Z(n1435) );
  XNOR U1529 ( .A(n1439), .B(n1440), .Z(o[912]) );
  AND U1530 ( .A(n1441), .B(n1442), .Z(n1439) );
  XNOR U1531 ( .A(n1443), .B(n1444), .Z(o[911]) );
  AND U1532 ( .A(n1445), .B(n1446), .Z(n1443) );
  XNOR U1533 ( .A(n1447), .B(n1448), .Z(o[910]) );
  AND U1534 ( .A(n1449), .B(n1450), .Z(n1447) );
  XNOR U1535 ( .A(n1451), .B(n1452), .Z(o[90]) );
  AND U1536 ( .A(n1453), .B(n1454), .Z(n1451) );
  XNOR U1537 ( .A(n1455), .B(n1456), .Z(o[909]) );
  AND U1538 ( .A(n1457), .B(n1458), .Z(n1455) );
  XNOR U1539 ( .A(n1459), .B(n1460), .Z(o[908]) );
  AND U1540 ( .A(n1461), .B(n1462), .Z(n1459) );
  XNOR U1541 ( .A(n1463), .B(n1464), .Z(o[907]) );
  AND U1542 ( .A(n1465), .B(n1466), .Z(n1463) );
  XNOR U1543 ( .A(n1467), .B(n1468), .Z(o[906]) );
  AND U1544 ( .A(n1469), .B(n1470), .Z(n1467) );
  XNOR U1545 ( .A(n1471), .B(n1472), .Z(o[905]) );
  AND U1546 ( .A(n1473), .B(n1474), .Z(n1471) );
  XNOR U1547 ( .A(n1475), .B(n1476), .Z(o[904]) );
  AND U1548 ( .A(n1477), .B(n1478), .Z(n1475) );
  XNOR U1549 ( .A(n1479), .B(n1480), .Z(o[903]) );
  AND U1550 ( .A(n1481), .B(n1482), .Z(n1479) );
  XNOR U1551 ( .A(n1483), .B(n1484), .Z(o[902]) );
  AND U1552 ( .A(n1485), .B(n1486), .Z(n1483) );
  XNOR U1553 ( .A(n1487), .B(n1488), .Z(o[901]) );
  AND U1554 ( .A(n1489), .B(n1490), .Z(n1487) );
  XNOR U1555 ( .A(n1491), .B(n1492), .Z(o[900]) );
  AND U1556 ( .A(n1493), .B(n1494), .Z(n1491) );
  XNOR U1557 ( .A(n1495), .B(n1496), .Z(o[8]) );
  NOR U1558 ( .A(n1497), .B(n1498), .Z(n1495) );
  XNOR U1559 ( .A(n1499), .B(n1500), .Z(o[89]) );
  AND U1560 ( .A(n1501), .B(n1502), .Z(n1499) );
  XNOR U1561 ( .A(n1503), .B(n1504), .Z(o[899]) );
  AND U1562 ( .A(n1505), .B(n1506), .Z(n1503) );
  XNOR U1563 ( .A(n1507), .B(n1508), .Z(o[898]) );
  AND U1564 ( .A(n1509), .B(n1510), .Z(n1507) );
  XNOR U1565 ( .A(n1511), .B(n1512), .Z(o[897]) );
  AND U1566 ( .A(n1513), .B(n1514), .Z(n1511) );
  XNOR U1567 ( .A(n1515), .B(n1516), .Z(o[896]) );
  AND U1568 ( .A(n1517), .B(n1518), .Z(n1515) );
  XNOR U1569 ( .A(n1519), .B(n1237), .Z(o[895]) );
  XNOR U1570 ( .A(n1521), .B(n1241), .Z(o[894]) );
  XNOR U1571 ( .A(n1523), .B(n1245), .Z(o[893]) );
  XNOR U1572 ( .A(n1525), .B(n1249), .Z(o[892]) );
  XNOR U1573 ( .A(n1527), .B(n1253), .Z(o[891]) );
  XNOR U1574 ( .A(n1529), .B(n1257), .Z(o[890]) );
  XNOR U1575 ( .A(n1531), .B(n1532), .Z(o[88]) );
  AND U1576 ( .A(n1533), .B(n1534), .Z(n1531) );
  XNOR U1577 ( .A(n1535), .B(n1261), .Z(o[889]) );
  AND U1578 ( .A(n1536), .B(n1537), .Z(n1535) );
  XNOR U1579 ( .A(n1538), .B(n1265), .Z(o[888]) );
  AND U1580 ( .A(n1539), .B(n1540), .Z(n1538) );
  XNOR U1581 ( .A(n1541), .B(n1269), .Z(o[887]) );
  AND U1582 ( .A(n1542), .B(n1543), .Z(n1541) );
  XNOR U1583 ( .A(n1544), .B(n1273), .Z(o[886]) );
  AND U1584 ( .A(n1545), .B(n1546), .Z(n1544) );
  XNOR U1585 ( .A(n1547), .B(n1281), .Z(o[885]) );
  AND U1586 ( .A(n1548), .B(n1549), .Z(n1547) );
  XNOR U1587 ( .A(n1550), .B(n1285), .Z(o[884]) );
  AND U1588 ( .A(n1551), .B(n1552), .Z(n1550) );
  XNOR U1589 ( .A(n1553), .B(n1289), .Z(o[883]) );
  XNOR U1590 ( .A(n1555), .B(n1293), .Z(o[882]) );
  XNOR U1591 ( .A(n1557), .B(n1297), .Z(o[881]) );
  XNOR U1592 ( .A(n1559), .B(n1301), .Z(o[880]) );
  XNOR U1593 ( .A(n1561), .B(n1562), .Z(o[87]) );
  AND U1594 ( .A(n1563), .B(n1564), .Z(n1561) );
  XNOR U1595 ( .A(n1565), .B(n1305), .Z(o[879]) );
  XNOR U1596 ( .A(n1567), .B(n1309), .Z(o[878]) );
  XNOR U1597 ( .A(n1569), .B(n1313), .Z(o[877]) );
  XNOR U1598 ( .A(n1571), .B(n1317), .Z(o[876]) );
  XNOR U1599 ( .A(n1573), .B(n1325), .Z(o[875]) );
  AND U1600 ( .A(n1574), .B(n1575), .Z(n1573) );
  XNOR U1601 ( .A(n1576), .B(n1329), .Z(o[874]) );
  XNOR U1602 ( .A(n1578), .B(n1333), .Z(o[873]) );
  XNOR U1603 ( .A(n1580), .B(n1337), .Z(o[872]) );
  XNOR U1604 ( .A(n1582), .B(n1341), .Z(o[871]) );
  XNOR U1605 ( .A(n1584), .B(n1345), .Z(o[870]) );
  XNOR U1606 ( .A(n1586), .B(n1587), .Z(o[86]) );
  AND U1607 ( .A(n1588), .B(n1589), .Z(n1586) );
  XNOR U1608 ( .A(n1590), .B(n1349), .Z(o[869]) );
  XNOR U1609 ( .A(n1592), .B(n1353), .Z(o[868]) );
  AND U1610 ( .A(n1593), .B(n1594), .Z(n1592) );
  XNOR U1611 ( .A(n1595), .B(n1357), .Z(o[867]) );
  AND U1612 ( .A(n1596), .B(n1597), .Z(n1595) );
  XNOR U1613 ( .A(n1598), .B(n1361), .Z(o[866]) );
  AND U1614 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1615 ( .A(n1601), .B(n1369), .Z(o[865]) );
  AND U1616 ( .A(n1602), .B(n1603), .Z(n1601) );
  XNOR U1617 ( .A(n1604), .B(n1373), .Z(o[864]) );
  AND U1618 ( .A(n1605), .B(n1606), .Z(n1604) );
  XNOR U1619 ( .A(n1607), .B(n1377), .Z(o[863]) );
  AND U1620 ( .A(n1608), .B(n1609), .Z(n1607) );
  XNOR U1621 ( .A(n1610), .B(n1381), .Z(o[862]) );
  AND U1622 ( .A(n1611), .B(n1612), .Z(n1610) );
  XNOR U1623 ( .A(n1613), .B(n1385), .Z(o[861]) );
  AND U1624 ( .A(n1614), .B(n1615), .Z(n1613) );
  XNOR U1625 ( .A(n1616), .B(n1389), .Z(o[860]) );
  AND U1626 ( .A(n1617), .B(n1618), .Z(n1616) );
  XNOR U1627 ( .A(n1619), .B(n1620), .Z(o[85]) );
  AND U1628 ( .A(n1621), .B(n1622), .Z(n1619) );
  XNOR U1629 ( .A(n1623), .B(n1393), .Z(o[859]) );
  AND U1630 ( .A(n1624), .B(n1625), .Z(n1623) );
  XNOR U1631 ( .A(n1626), .B(n1397), .Z(o[858]) );
  AND U1632 ( .A(n1627), .B(n1628), .Z(n1626) );
  XNOR U1633 ( .A(n1629), .B(n1401), .Z(o[857]) );
  AND U1634 ( .A(n1630), .B(n1631), .Z(n1629) );
  XNOR U1635 ( .A(n1632), .B(n1405), .Z(o[856]) );
  AND U1636 ( .A(n1633), .B(n1634), .Z(n1632) );
  XNOR U1637 ( .A(n1635), .B(n1413), .Z(o[855]) );
  AND U1638 ( .A(n1636), .B(n1637), .Z(n1635) );
  XNOR U1639 ( .A(n1638), .B(n1417), .Z(o[854]) );
  AND U1640 ( .A(n1639), .B(n1640), .Z(n1638) );
  XNOR U1641 ( .A(n1641), .B(n1421), .Z(o[853]) );
  AND U1642 ( .A(n1642), .B(n1643), .Z(n1641) );
  XNOR U1643 ( .A(n1644), .B(n1425), .Z(o[852]) );
  AND U1644 ( .A(n1645), .B(n1646), .Z(n1644) );
  XNOR U1645 ( .A(n1647), .B(n1429), .Z(o[851]) );
  AND U1646 ( .A(n1648), .B(n1649), .Z(n1647) );
  XNOR U1647 ( .A(n1650), .B(n1433), .Z(o[850]) );
  AND U1648 ( .A(n1651), .B(n1652), .Z(n1650) );
  XNOR U1649 ( .A(n1653), .B(n1654), .Z(o[84]) );
  AND U1650 ( .A(n1655), .B(n1656), .Z(n1653) );
  XNOR U1651 ( .A(n1657), .B(n1437), .Z(o[849]) );
  AND U1652 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1653 ( .A(n1660), .B(n1441), .Z(o[848]) );
  AND U1654 ( .A(n1661), .B(n1662), .Z(n1660) );
  XNOR U1655 ( .A(n1663), .B(n1445), .Z(o[847]) );
  AND U1656 ( .A(n1664), .B(n1665), .Z(n1663) );
  XNOR U1657 ( .A(n1666), .B(n1449), .Z(o[846]) );
  AND U1658 ( .A(n1667), .B(n1668), .Z(n1666) );
  XNOR U1659 ( .A(n1669), .B(n1457), .Z(o[845]) );
  AND U1660 ( .A(n1670), .B(n1671), .Z(n1669) );
  XNOR U1661 ( .A(n1672), .B(n1461), .Z(o[844]) );
  AND U1662 ( .A(n1673), .B(n1674), .Z(n1672) );
  XNOR U1663 ( .A(n1675), .B(n1465), .Z(o[843]) );
  AND U1664 ( .A(n1676), .B(n1677), .Z(n1675) );
  XNOR U1665 ( .A(n1678), .B(n1469), .Z(o[842]) );
  AND U1666 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1667 ( .A(n1681), .B(n1473), .Z(o[841]) );
  AND U1668 ( .A(n1682), .B(n1683), .Z(n1681) );
  XNOR U1669 ( .A(n1684), .B(n1477), .Z(o[840]) );
  AND U1670 ( .A(n1685), .B(n1686), .Z(n1684) );
  XNOR U1671 ( .A(n1687), .B(n1688), .Z(o[83]) );
  AND U1672 ( .A(n1689), .B(n1690), .Z(n1687) );
  XNOR U1673 ( .A(n1691), .B(n1481), .Z(o[839]) );
  AND U1674 ( .A(n1692), .B(n1693), .Z(n1691) );
  XNOR U1675 ( .A(n1694), .B(n1485), .Z(o[838]) );
  AND U1676 ( .A(n1695), .B(n1696), .Z(n1694) );
  XNOR U1677 ( .A(n1697), .B(n1489), .Z(o[837]) );
  XNOR U1678 ( .A(n1699), .B(n1493), .Z(o[836]) );
  XNOR U1679 ( .A(n1701), .B(n1505), .Z(o[835]) );
  XNOR U1680 ( .A(n1703), .B(n1509), .Z(o[834]) );
  XNOR U1681 ( .A(n1705), .B(n1513), .Z(o[833]) );
  XNOR U1682 ( .A(n1707), .B(n1517), .Z(o[832]) );
  XOR U1683 ( .A(n1709), .B(n1238), .Z(o[831]) );
  XNOR U1684 ( .A(n1710), .B(round_reg[742]), .Z(n1238) );
  XOR U1685 ( .A(n1712), .B(n1242), .Z(o[830]) );
  XNOR U1686 ( .A(n1713), .B(round_reg[741]), .Z(n1242) );
  XNOR U1687 ( .A(n1715), .B(n1716), .Z(o[82]) );
  AND U1688 ( .A(n1717), .B(n1718), .Z(n1715) );
  XOR U1689 ( .A(n1719), .B(n1246), .Z(o[829]) );
  XNOR U1690 ( .A(n1720), .B(round_reg[740]), .Z(n1246) );
  XOR U1691 ( .A(n1722), .B(n1250), .Z(o[828]) );
  XNOR U1692 ( .A(n1723), .B(round_reg[739]), .Z(n1250) );
  NOR U1693 ( .A(n1724), .B(n1526), .Z(n1722) );
  XOR U1694 ( .A(n1725), .B(n1254), .Z(o[827]) );
  XNOR U1695 ( .A(n1726), .B(round_reg[738]), .Z(n1254) );
  NOR U1696 ( .A(n1727), .B(n1528), .Z(n1725) );
  XOR U1697 ( .A(n1728), .B(n1258), .Z(o[826]) );
  XNOR U1698 ( .A(n1729), .B(round_reg[737]), .Z(n1258) );
  NOR U1699 ( .A(n1730), .B(n1530), .Z(n1728) );
  XOR U1700 ( .A(n1731), .B(n1262), .Z(o[825]) );
  IV U1701 ( .A(n1537), .Z(n1262) );
  XNOR U1702 ( .A(n1732), .B(round_reg[736]), .Z(n1537) );
  NOR U1703 ( .A(n1733), .B(n1536), .Z(n1731) );
  XOR U1704 ( .A(n1734), .B(n1266), .Z(o[824]) );
  IV U1705 ( .A(n1540), .Z(n1266) );
  XNOR U1706 ( .A(n1735), .B(round_reg[735]), .Z(n1540) );
  NOR U1707 ( .A(n1736), .B(n1539), .Z(n1734) );
  XOR U1708 ( .A(n1737), .B(n1270), .Z(o[823]) );
  IV U1709 ( .A(n1543), .Z(n1270) );
  XNOR U1710 ( .A(n1738), .B(round_reg[734]), .Z(n1543) );
  NOR U1711 ( .A(n1739), .B(n1542), .Z(n1737) );
  XOR U1712 ( .A(n1740), .B(n1274), .Z(o[822]) );
  IV U1713 ( .A(n1546), .Z(n1274) );
  XNOR U1714 ( .A(n1741), .B(round_reg[733]), .Z(n1546) );
  NOR U1715 ( .A(n1742), .B(n1545), .Z(n1740) );
  XOR U1716 ( .A(n1743), .B(n1282), .Z(o[821]) );
  IV U1717 ( .A(n1549), .Z(n1282) );
  XNOR U1718 ( .A(n1744), .B(round_reg[732]), .Z(n1549) );
  NOR U1719 ( .A(n1745), .B(n1548), .Z(n1743) );
  XOR U1720 ( .A(n1746), .B(n1286), .Z(o[820]) );
  IV U1721 ( .A(n1552), .Z(n1286) );
  XNOR U1722 ( .A(n1747), .B(round_reg[731]), .Z(n1552) );
  NOR U1723 ( .A(n1748), .B(n1551), .Z(n1746) );
  XNOR U1724 ( .A(n1749), .B(n1750), .Z(o[81]) );
  AND U1725 ( .A(n1751), .B(n1752), .Z(n1749) );
  XOR U1726 ( .A(n1753), .B(n1290), .Z(o[819]) );
  XNOR U1727 ( .A(n1754), .B(round_reg[730]), .Z(n1290) );
  NOR U1728 ( .A(n1755), .B(n1554), .Z(n1753) );
  XOR U1729 ( .A(n1756), .B(n1294), .Z(o[818]) );
  XNOR U1730 ( .A(n1757), .B(round_reg[729]), .Z(n1294) );
  NOR U1731 ( .A(n1758), .B(n1556), .Z(n1756) );
  XOR U1732 ( .A(n1759), .B(n1298), .Z(o[817]) );
  XNOR U1733 ( .A(n1760), .B(round_reg[728]), .Z(n1298) );
  XOR U1734 ( .A(n1762), .B(n1302), .Z(o[816]) );
  XNOR U1735 ( .A(n1763), .B(round_reg[727]), .Z(n1302) );
  XOR U1736 ( .A(n1765), .B(n1306), .Z(o[815]) );
  XNOR U1737 ( .A(n1766), .B(round_reg[726]), .Z(n1306) );
  XOR U1738 ( .A(n1768), .B(n1310), .Z(o[814]) );
  XNOR U1739 ( .A(n1769), .B(round_reg[725]), .Z(n1310) );
  XOR U1740 ( .A(n1771), .B(n1314), .Z(o[813]) );
  XNOR U1741 ( .A(n1772), .B(round_reg[724]), .Z(n1314) );
  XOR U1742 ( .A(n1774), .B(n1318), .Z(o[812]) );
  XNOR U1743 ( .A(n1775), .B(round_reg[723]), .Z(n1318) );
  XOR U1744 ( .A(n1777), .B(n1326), .Z(o[811]) );
  IV U1745 ( .A(n1575), .Z(n1326) );
  XNOR U1746 ( .A(n1778), .B(round_reg[722]), .Z(n1575) );
  XOR U1747 ( .A(n1780), .B(n1330), .Z(o[810]) );
  XOR U1748 ( .A(n1781), .B(round_reg[721]), .Z(n1330) );
  XNOR U1749 ( .A(n1783), .B(n1784), .Z(o[80]) );
  AND U1750 ( .A(n1785), .B(n1786), .Z(n1783) );
  XOR U1751 ( .A(n1787), .B(n1334), .Z(o[809]) );
  XOR U1752 ( .A(n1788), .B(round_reg[720]), .Z(n1334) );
  XOR U1753 ( .A(n1790), .B(n1338), .Z(o[808]) );
  XOR U1754 ( .A(n1791), .B(round_reg[719]), .Z(n1338) );
  XOR U1755 ( .A(n1793), .B(n1342), .Z(o[807]) );
  XOR U1756 ( .A(n1794), .B(round_reg[718]), .Z(n1342) );
  XOR U1757 ( .A(n1796), .B(n1346), .Z(o[806]) );
  XOR U1758 ( .A(n1797), .B(round_reg[717]), .Z(n1346) );
  XOR U1759 ( .A(n1799), .B(n1350), .Z(o[805]) );
  XOR U1760 ( .A(n1800), .B(round_reg[716]), .Z(n1350) );
  XOR U1761 ( .A(n1802), .B(n1354), .Z(o[804]) );
  IV U1762 ( .A(n1594), .Z(n1354) );
  XNOR U1763 ( .A(n1803), .B(round_reg[715]), .Z(n1594) );
  XOR U1764 ( .A(n1805), .B(n1358), .Z(o[803]) );
  IV U1765 ( .A(n1597), .Z(n1358) );
  XNOR U1766 ( .A(n1806), .B(round_reg[714]), .Z(n1597) );
  XOR U1767 ( .A(n1808), .B(n1362), .Z(o[802]) );
  IV U1768 ( .A(n1600), .Z(n1362) );
  XNOR U1769 ( .A(n1809), .B(round_reg[713]), .Z(n1600) );
  XOR U1770 ( .A(n1811), .B(n1370), .Z(o[801]) );
  IV U1771 ( .A(n1603), .Z(n1370) );
  XNOR U1772 ( .A(n1812), .B(round_reg[712]), .Z(n1603) );
  XOR U1773 ( .A(n1814), .B(n1374), .Z(o[800]) );
  IV U1774 ( .A(n1606), .Z(n1374) );
  XNOR U1775 ( .A(n1815), .B(round_reg[711]), .Z(n1606) );
  XNOR U1776 ( .A(n1817), .B(n1818), .Z(o[7]) );
  NOR U1777 ( .A(n1819), .B(n1820), .Z(n1817) );
  XNOR U1778 ( .A(n1821), .B(n1822), .Z(o[79]) );
  AND U1779 ( .A(n1823), .B(n1824), .Z(n1821) );
  XOR U1780 ( .A(n1825), .B(n1378), .Z(o[799]) );
  IV U1781 ( .A(n1609), .Z(n1378) );
  XNOR U1782 ( .A(n1826), .B(round_reg[710]), .Z(n1609) );
  XOR U1783 ( .A(n1828), .B(n1382), .Z(o[798]) );
  IV U1784 ( .A(n1612), .Z(n1382) );
  XNOR U1785 ( .A(n1829), .B(round_reg[709]), .Z(n1612) );
  XOR U1786 ( .A(n1831), .B(n1386), .Z(o[797]) );
  IV U1787 ( .A(n1615), .Z(n1386) );
  XNOR U1788 ( .A(n1832), .B(round_reg[708]), .Z(n1615) );
  XOR U1789 ( .A(n1834), .B(n1390), .Z(o[796]) );
  IV U1790 ( .A(n1618), .Z(n1390) );
  XNOR U1791 ( .A(n1835), .B(round_reg[707]), .Z(n1618) );
  XOR U1792 ( .A(n1837), .B(n1394), .Z(o[795]) );
  IV U1793 ( .A(n1625), .Z(n1394) );
  XNOR U1794 ( .A(n1838), .B(round_reg[706]), .Z(n1625) );
  NOR U1795 ( .A(n1839), .B(n1624), .Z(n1837) );
  XOR U1796 ( .A(n1840), .B(n1398), .Z(o[794]) );
  IV U1797 ( .A(n1628), .Z(n1398) );
  XNOR U1798 ( .A(n1841), .B(round_reg[705]), .Z(n1628) );
  NOR U1799 ( .A(n1842), .B(n1627), .Z(n1840) );
  XOR U1800 ( .A(n1843), .B(n1402), .Z(o[793]) );
  IV U1801 ( .A(n1631), .Z(n1402) );
  XNOR U1802 ( .A(n1844), .B(round_reg[704]), .Z(n1631) );
  NOR U1803 ( .A(n1845), .B(n1630), .Z(n1843) );
  XOR U1804 ( .A(n1846), .B(n1406), .Z(o[792]) );
  IV U1805 ( .A(n1634), .Z(n1406) );
  XNOR U1806 ( .A(n1847), .B(round_reg[767]), .Z(n1634) );
  NOR U1807 ( .A(n1848), .B(n1633), .Z(n1846) );
  XOR U1808 ( .A(n1849), .B(n1414), .Z(o[791]) );
  IV U1809 ( .A(n1637), .Z(n1414) );
  XNOR U1810 ( .A(n1850), .B(round_reg[766]), .Z(n1637) );
  ANDN U1811 ( .A(n1851), .B(n1636), .Z(n1849) );
  XOR U1812 ( .A(n1852), .B(n1418), .Z(o[790]) );
  IV U1813 ( .A(n1640), .Z(n1418) );
  XNOR U1814 ( .A(n1853), .B(round_reg[765]), .Z(n1640) );
  NOR U1815 ( .A(n1854), .B(n1639), .Z(n1852) );
  XNOR U1816 ( .A(n1855), .B(n1856), .Z(o[78]) );
  AND U1817 ( .A(n1857), .B(n1858), .Z(n1855) );
  XOR U1818 ( .A(n1859), .B(n1422), .Z(o[789]) );
  IV U1819 ( .A(n1643), .Z(n1422) );
  XNOR U1820 ( .A(n1860), .B(round_reg[764]), .Z(n1643) );
  NOR U1821 ( .A(n1861), .B(n1642), .Z(n1859) );
  XOR U1822 ( .A(n1862), .B(n1426), .Z(o[788]) );
  IV U1823 ( .A(n1646), .Z(n1426) );
  XNOR U1824 ( .A(n1863), .B(round_reg[763]), .Z(n1646) );
  NOR U1825 ( .A(n1864), .B(n1645), .Z(n1862) );
  XOR U1826 ( .A(n1865), .B(n1430), .Z(o[787]) );
  IV U1827 ( .A(n1649), .Z(n1430) );
  XNOR U1828 ( .A(n1866), .B(round_reg[762]), .Z(n1649) );
  NOR U1829 ( .A(n1867), .B(n1648), .Z(n1865) );
  XOR U1830 ( .A(n1868), .B(n1434), .Z(o[786]) );
  IV U1831 ( .A(n1652), .Z(n1434) );
  XNOR U1832 ( .A(n1869), .B(round_reg[761]), .Z(n1652) );
  NOR U1833 ( .A(n1870), .B(n1651), .Z(n1868) );
  XOR U1834 ( .A(n1871), .B(n1438), .Z(o[785]) );
  IV U1835 ( .A(n1659), .Z(n1438) );
  XNOR U1836 ( .A(n1872), .B(round_reg[760]), .Z(n1659) );
  NOR U1837 ( .A(n1873), .B(n1658), .Z(n1871) );
  XOR U1838 ( .A(n1874), .B(n1442), .Z(o[784]) );
  IV U1839 ( .A(n1662), .Z(n1442) );
  XNOR U1840 ( .A(n1875), .B(round_reg[759]), .Z(n1662) );
  NOR U1841 ( .A(n1876), .B(n1661), .Z(n1874) );
  XOR U1842 ( .A(n1877), .B(n1446), .Z(o[783]) );
  IV U1843 ( .A(n1665), .Z(n1446) );
  XNOR U1844 ( .A(n1878), .B(round_reg[758]), .Z(n1665) );
  NOR U1845 ( .A(n1879), .B(n1664), .Z(n1877) );
  XOR U1846 ( .A(n1880), .B(n1450), .Z(o[782]) );
  IV U1847 ( .A(n1668), .Z(n1450) );
  XNOR U1848 ( .A(n1881), .B(round_reg[757]), .Z(n1668) );
  NOR U1849 ( .A(n1882), .B(n1667), .Z(n1880) );
  XOR U1850 ( .A(n1883), .B(n1458), .Z(o[781]) );
  IV U1851 ( .A(n1671), .Z(n1458) );
  XNOR U1852 ( .A(n1884), .B(round_reg[756]), .Z(n1671) );
  NOR U1853 ( .A(n1885), .B(n1670), .Z(n1883) );
  XOR U1854 ( .A(n1886), .B(n1462), .Z(o[780]) );
  IV U1855 ( .A(n1674), .Z(n1462) );
  XNOR U1856 ( .A(n1887), .B(round_reg[755]), .Z(n1674) );
  ANDN U1857 ( .A(n1888), .B(n1673), .Z(n1886) );
  XNOR U1858 ( .A(n1889), .B(n1890), .Z(o[77]) );
  NOR U1859 ( .A(n1891), .B(n1892), .Z(n1889) );
  XOR U1860 ( .A(n1893), .B(n1466), .Z(o[779]) );
  IV U1861 ( .A(n1677), .Z(n1466) );
  XNOR U1862 ( .A(n1894), .B(round_reg[754]), .Z(n1677) );
  ANDN U1863 ( .A(n1895), .B(n1676), .Z(n1893) );
  XOR U1864 ( .A(n1896), .B(n1470), .Z(o[778]) );
  IV U1865 ( .A(n1680), .Z(n1470) );
  XNOR U1866 ( .A(n1897), .B(round_reg[753]), .Z(n1680) );
  ANDN U1867 ( .A(n1898), .B(n1679), .Z(n1896) );
  XOR U1868 ( .A(n1899), .B(n1474), .Z(o[777]) );
  IV U1869 ( .A(n1683), .Z(n1474) );
  XNOR U1870 ( .A(n1900), .B(round_reg[752]), .Z(n1683) );
  ANDN U1871 ( .A(n1901), .B(n1682), .Z(n1899) );
  XOR U1872 ( .A(n1902), .B(n1478), .Z(o[776]) );
  IV U1873 ( .A(n1686), .Z(n1478) );
  XNOR U1874 ( .A(n1903), .B(round_reg[751]), .Z(n1686) );
  ANDN U1875 ( .A(n1904), .B(n1685), .Z(n1902) );
  XOR U1876 ( .A(n1905), .B(n1482), .Z(o[775]) );
  IV U1877 ( .A(n1693), .Z(n1482) );
  XNOR U1878 ( .A(n1906), .B(round_reg[750]), .Z(n1693) );
  XOR U1879 ( .A(n1908), .B(n1486), .Z(o[774]) );
  IV U1880 ( .A(n1696), .Z(n1486) );
  XNOR U1881 ( .A(n1909), .B(round_reg[749]), .Z(n1696) );
  NOR U1882 ( .A(n1910), .B(n1695), .Z(n1908) );
  XOR U1883 ( .A(n1911), .B(n1490), .Z(o[773]) );
  XNOR U1884 ( .A(n1912), .B(round_reg[748]), .Z(n1490) );
  NOR U1885 ( .A(n1913), .B(n1698), .Z(n1911) );
  XOR U1886 ( .A(n1914), .B(n1494), .Z(o[772]) );
  XNOR U1887 ( .A(n1915), .B(round_reg[747]), .Z(n1494) );
  NOR U1888 ( .A(n1916), .B(n1700), .Z(n1914) );
  XOR U1889 ( .A(n1917), .B(n1506), .Z(o[771]) );
  XNOR U1890 ( .A(n1918), .B(round_reg[746]), .Z(n1506) );
  NOR U1891 ( .A(n1919), .B(n1702), .Z(n1917) );
  XOR U1892 ( .A(n1920), .B(n1510), .Z(o[770]) );
  XNOR U1893 ( .A(n1921), .B(round_reg[745]), .Z(n1510) );
  NOR U1894 ( .A(n1922), .B(n1704), .Z(n1920) );
  XNOR U1895 ( .A(n1923), .B(n1924), .Z(o[76]) );
  NOR U1896 ( .A(n1925), .B(n1926), .Z(n1923) );
  XOR U1897 ( .A(n1927), .B(n1514), .Z(o[769]) );
  XNOR U1898 ( .A(n1928), .B(round_reg[744]), .Z(n1514) );
  NOR U1899 ( .A(n1929), .B(n1706), .Z(n1927) );
  XOR U1900 ( .A(n1930), .B(n1518), .Z(o[768]) );
  XNOR U1901 ( .A(n1931), .B(round_reg[743]), .Z(n1518) );
  XOR U1902 ( .A(n1933), .B(n1520), .Z(o[767]) );
  XOR U1903 ( .A(n1934), .B(round_reg[375]), .Z(n1520) );
  XOR U1904 ( .A(n1935), .B(n1522), .Z(o[766]) );
  XOR U1905 ( .A(n1936), .B(round_reg[374]), .Z(n1522) );
  XOR U1906 ( .A(n1937), .B(n1524), .Z(o[765]) );
  XOR U1907 ( .A(n1938), .B(round_reg[373]), .Z(n1524) );
  XOR U1908 ( .A(n1939), .B(n1526), .Z(o[764]) );
  XOR U1909 ( .A(n1940), .B(round_reg[372]), .Z(n1526) );
  AND U1910 ( .A(n1248), .B(n1724), .Z(n1939) );
  IV U1911 ( .A(n1941), .Z(n1724) );
  XOR U1912 ( .A(n1942), .B(n1528), .Z(o[763]) );
  XOR U1913 ( .A(n1943), .B(round_reg[371]), .Z(n1528) );
  AND U1914 ( .A(n1252), .B(n1727), .Z(n1942) );
  IV U1915 ( .A(n1944), .Z(n1727) );
  XOR U1916 ( .A(n1945), .B(n1530), .Z(o[762]) );
  XOR U1917 ( .A(n1946), .B(round_reg[370]), .Z(n1530) );
  ANDN U1918 ( .A(n1730), .B(n1256), .Z(n1945) );
  IV U1919 ( .A(n1947), .Z(n1730) );
  XOR U1920 ( .A(n1948), .B(n1536), .Z(o[761]) );
  XOR U1921 ( .A(n1949), .B(round_reg[369]), .Z(n1536) );
  ANDN U1922 ( .A(n1733), .B(n1260), .Z(n1948) );
  IV U1923 ( .A(n1950), .Z(n1733) );
  XOR U1924 ( .A(n1951), .B(n1539), .Z(o[760]) );
  XOR U1925 ( .A(n1952), .B(round_reg[368]), .Z(n1539) );
  ANDN U1926 ( .A(n1736), .B(n1264), .Z(n1951) );
  IV U1927 ( .A(n1953), .Z(n1736) );
  XNOR U1928 ( .A(n1954), .B(n1955), .Z(o[75]) );
  NOR U1929 ( .A(n1956), .B(n1957), .Z(n1954) );
  XOR U1930 ( .A(n1958), .B(n1542), .Z(o[759]) );
  XOR U1931 ( .A(n1959), .B(round_reg[367]), .Z(n1542) );
  ANDN U1932 ( .A(n1739), .B(n1268), .Z(n1958) );
  IV U1933 ( .A(n1960), .Z(n1739) );
  XOR U1934 ( .A(n1961), .B(n1545), .Z(o[758]) );
  XOR U1935 ( .A(n1962), .B(round_reg[366]), .Z(n1545) );
  ANDN U1936 ( .A(n1742), .B(n1272), .Z(n1961) );
  IV U1937 ( .A(n1963), .Z(n1742) );
  XOR U1938 ( .A(n1964), .B(n1548), .Z(o[757]) );
  XOR U1939 ( .A(n1965), .B(round_reg[365]), .Z(n1548) );
  ANDN U1940 ( .A(n1745), .B(n1280), .Z(n1964) );
  IV U1941 ( .A(n1966), .Z(n1745) );
  XOR U1942 ( .A(n1967), .B(n1551), .Z(o[756]) );
  XOR U1943 ( .A(n1968), .B(round_reg[364]), .Z(n1551) );
  ANDN U1944 ( .A(n1748), .B(n1284), .Z(n1967) );
  IV U1945 ( .A(n1969), .Z(n1748) );
  XOR U1946 ( .A(n1970), .B(n1554), .Z(o[755]) );
  XOR U1947 ( .A(n1971), .B(round_reg[363]), .Z(n1554) );
  ANDN U1948 ( .A(n1755), .B(n1288), .Z(n1970) );
  IV U1949 ( .A(n1972), .Z(n1755) );
  XOR U1950 ( .A(n1973), .B(n1556), .Z(o[754]) );
  XOR U1951 ( .A(n1974), .B(round_reg[362]), .Z(n1556) );
  ANDN U1952 ( .A(n1758), .B(n1292), .Z(n1973) );
  IV U1953 ( .A(n1975), .Z(n1758) );
  XOR U1954 ( .A(n1976), .B(n1558), .Z(o[753]) );
  XOR U1955 ( .A(n1977), .B(round_reg[361]), .Z(n1558) );
  NOR U1956 ( .A(n1761), .B(n1296), .Z(n1976) );
  XOR U1957 ( .A(n1978), .B(n1560), .Z(o[752]) );
  XOR U1958 ( .A(n1979), .B(round_reg[360]), .Z(n1560) );
  NOR U1959 ( .A(n1764), .B(n1300), .Z(n1978) );
  XOR U1960 ( .A(n1980), .B(n1566), .Z(o[751]) );
  XOR U1961 ( .A(n1981), .B(round_reg[359]), .Z(n1566) );
  NOR U1962 ( .A(n1767), .B(n1304), .Z(n1980) );
  XOR U1963 ( .A(n1982), .B(n1568), .Z(o[750]) );
  XOR U1964 ( .A(n1983), .B(round_reg[358]), .Z(n1568) );
  NOR U1965 ( .A(n1770), .B(n1308), .Z(n1982) );
  XNOR U1966 ( .A(n1984), .B(n1985), .Z(o[74]) );
  NOR U1967 ( .A(n1986), .B(n1987), .Z(n1984) );
  XOR U1968 ( .A(n1988), .B(n1570), .Z(o[749]) );
  XOR U1969 ( .A(n1989), .B(round_reg[357]), .Z(n1570) );
  NOR U1970 ( .A(n1773), .B(n1312), .Z(n1988) );
  XOR U1971 ( .A(n1990), .B(n1572), .Z(o[748]) );
  XOR U1972 ( .A(n1991), .B(round_reg[356]), .Z(n1572) );
  NOR U1973 ( .A(n1776), .B(n1316), .Z(n1990) );
  XOR U1974 ( .A(n1992), .B(n1574), .Z(o[747]) );
  XOR U1975 ( .A(n1993), .B(round_reg[355]), .Z(n1574) );
  XOR U1976 ( .A(n1994), .B(n1577), .Z(o[746]) );
  XOR U1977 ( .A(n1995), .B(round_reg[354]), .Z(n1577) );
  XOR U1978 ( .A(n1996), .B(n1579), .Z(o[745]) );
  XOR U1979 ( .A(n1997), .B(round_reg[353]), .Z(n1579) );
  XOR U1980 ( .A(n1998), .B(n1581), .Z(o[744]) );
  XOR U1981 ( .A(n1999), .B(round_reg[352]), .Z(n1581) );
  XOR U1982 ( .A(n2000), .B(n1583), .Z(o[743]) );
  XOR U1983 ( .A(n2001), .B(round_reg[351]), .Z(n1583) );
  XOR U1984 ( .A(n2002), .B(n1585), .Z(o[742]) );
  XOR U1985 ( .A(n2003), .B(round_reg[350]), .Z(n1585) );
  XOR U1986 ( .A(n2004), .B(n1591), .Z(o[741]) );
  XOR U1987 ( .A(n2005), .B(round_reg[349]), .Z(n1591) );
  XOR U1988 ( .A(n2006), .B(n1593), .Z(o[740]) );
  XOR U1989 ( .A(n2007), .B(round_reg[348]), .Z(n1593) );
  XNOR U1990 ( .A(n2008), .B(n2009), .Z(o[73]) );
  AND U1991 ( .A(n1054), .B(n2010), .Z(n2008) );
  XOR U1992 ( .A(n2011), .B(n1596), .Z(o[739]) );
  XOR U1993 ( .A(n2012), .B(round_reg[347]), .Z(n1596) );
  XOR U1994 ( .A(n2013), .B(n1599), .Z(o[738]) );
  XOR U1995 ( .A(n2014), .B(round_reg[346]), .Z(n1599) );
  XOR U1996 ( .A(n2015), .B(n1602), .Z(o[737]) );
  XOR U1997 ( .A(n2016), .B(round_reg[345]), .Z(n1602) );
  XOR U1998 ( .A(n2017), .B(n1605), .Z(o[736]) );
  XOR U1999 ( .A(n2018), .B(round_reg[344]), .Z(n1605) );
  XOR U2000 ( .A(n2019), .B(n1608), .Z(o[735]) );
  XOR U2001 ( .A(n2020), .B(round_reg[343]), .Z(n1608) );
  XOR U2002 ( .A(n2021), .B(n1611), .Z(o[734]) );
  XOR U2003 ( .A(n2022), .B(round_reg[342]), .Z(n1611) );
  XOR U2004 ( .A(n2023), .B(n1614), .Z(o[733]) );
  XOR U2005 ( .A(n2024), .B(round_reg[341]), .Z(n1614) );
  XOR U2006 ( .A(n2025), .B(n1617), .Z(o[732]) );
  XOR U2007 ( .A(n2026), .B(round_reg[340]), .Z(n1617) );
  XOR U2008 ( .A(n2027), .B(n1624), .Z(o[731]) );
  XOR U2009 ( .A(n2028), .B(round_reg[339]), .Z(n1624) );
  ANDN U2010 ( .A(n1839), .B(n1392), .Z(n2027) );
  IV U2011 ( .A(n2029), .Z(n1839) );
  XOR U2012 ( .A(n2030), .B(n1627), .Z(o[730]) );
  XOR U2013 ( .A(n2031), .B(round_reg[338]), .Z(n1627) );
  ANDN U2014 ( .A(n1842), .B(n1396), .Z(n2030) );
  IV U2015 ( .A(n2032), .Z(n1842) );
  XNOR U2016 ( .A(n2033), .B(n2034), .Z(o[72]) );
  AND U2017 ( .A(n1498), .B(n1496), .Z(n2033) );
  XOR U2018 ( .A(n2035), .B(n1630), .Z(o[729]) );
  XOR U2019 ( .A(n2036), .B(round_reg[337]), .Z(n1630) );
  ANDN U2020 ( .A(n1845), .B(n1400), .Z(n2035) );
  IV U2021 ( .A(n2037), .Z(n1845) );
  XOR U2022 ( .A(n2038), .B(n1633), .Z(o[728]) );
  XOR U2023 ( .A(n2039), .B(round_reg[336]), .Z(n1633) );
  ANDN U2024 ( .A(n1848), .B(n1404), .Z(n2038) );
  IV U2025 ( .A(n2040), .Z(n1848) );
  XOR U2026 ( .A(n2041), .B(n1636), .Z(o[727]) );
  XOR U2027 ( .A(n2042), .B(round_reg[335]), .Z(n1636) );
  NOR U2028 ( .A(n1851), .B(n1412), .Z(n2041) );
  XOR U2029 ( .A(n2043), .B(n1639), .Z(o[726]) );
  XOR U2030 ( .A(n2044), .B(round_reg[334]), .Z(n1639) );
  ANDN U2031 ( .A(n1854), .B(n1416), .Z(n2043) );
  IV U2032 ( .A(n2045), .Z(n1854) );
  XOR U2033 ( .A(n2046), .B(n1642), .Z(o[725]) );
  XOR U2034 ( .A(n2047), .B(round_reg[333]), .Z(n1642) );
  ANDN U2035 ( .A(n1861), .B(n1420), .Z(n2046) );
  IV U2036 ( .A(n2048), .Z(n1861) );
  XOR U2037 ( .A(n2049), .B(n1645), .Z(o[724]) );
  XOR U2038 ( .A(n2050), .B(round_reg[332]), .Z(n1645) );
  ANDN U2039 ( .A(n1864), .B(n1424), .Z(n2049) );
  IV U2040 ( .A(n2051), .Z(n1864) );
  XOR U2041 ( .A(n2052), .B(n1648), .Z(o[723]) );
  XOR U2042 ( .A(n2053), .B(round_reg[331]), .Z(n1648) );
  ANDN U2043 ( .A(n1867), .B(n1428), .Z(n2052) );
  IV U2044 ( .A(n2054), .Z(n1867) );
  XOR U2045 ( .A(n2055), .B(n1651), .Z(o[722]) );
  XOR U2046 ( .A(n2056), .B(round_reg[330]), .Z(n1651) );
  ANDN U2047 ( .A(n1870), .B(n1432), .Z(n2055) );
  IV U2048 ( .A(n2057), .Z(n1870) );
  XOR U2049 ( .A(n2058), .B(n1658), .Z(o[721]) );
  XOR U2050 ( .A(n2059), .B(round_reg[329]), .Z(n1658) );
  ANDN U2051 ( .A(n1873), .B(n1436), .Z(n2058) );
  IV U2052 ( .A(n2060), .Z(n1873) );
  XOR U2053 ( .A(n2061), .B(n1661), .Z(o[720]) );
  XOR U2054 ( .A(n2062), .B(round_reg[328]), .Z(n1661) );
  ANDN U2055 ( .A(n1876), .B(n1440), .Z(n2061) );
  IV U2056 ( .A(n2063), .Z(n1876) );
  XNOR U2057 ( .A(n2064), .B(n2065), .Z(o[71]) );
  AND U2058 ( .A(n1820), .B(n1818), .Z(n2064) );
  XOR U2059 ( .A(n2066), .B(n1664), .Z(o[719]) );
  XOR U2060 ( .A(n2067), .B(round_reg[327]), .Z(n1664) );
  ANDN U2061 ( .A(n1879), .B(n1444), .Z(n2066) );
  IV U2062 ( .A(n2068), .Z(n1879) );
  XOR U2063 ( .A(n2069), .B(n1667), .Z(o[718]) );
  XOR U2064 ( .A(n2070), .B(round_reg[326]), .Z(n1667) );
  ANDN U2065 ( .A(n1882), .B(n1448), .Z(n2069) );
  IV U2066 ( .A(n2071), .Z(n1882) );
  XOR U2067 ( .A(n2072), .B(n1670), .Z(o[717]) );
  XOR U2068 ( .A(n2073), .B(round_reg[325]), .Z(n1670) );
  ANDN U2069 ( .A(n1885), .B(n1456), .Z(n2072) );
  IV U2070 ( .A(n2074), .Z(n1885) );
  XOR U2071 ( .A(n2075), .B(n1673), .Z(o[716]) );
  XOR U2072 ( .A(n2076), .B(round_reg[324]), .Z(n1673) );
  NOR U2073 ( .A(n1888), .B(n1460), .Z(n2075) );
  XOR U2074 ( .A(n2077), .B(n1676), .Z(o[715]) );
  XOR U2075 ( .A(n2078), .B(round_reg[323]), .Z(n1676) );
  NOR U2076 ( .A(n1895), .B(n1464), .Z(n2077) );
  XOR U2077 ( .A(n2079), .B(n1679), .Z(o[714]) );
  XOR U2078 ( .A(n2080), .B(round_reg[322]), .Z(n1679) );
  NOR U2079 ( .A(n1898), .B(n1468), .Z(n2079) );
  XOR U2080 ( .A(n2081), .B(n1682), .Z(o[713]) );
  XOR U2081 ( .A(n2082), .B(round_reg[321]), .Z(n1682) );
  NOR U2082 ( .A(n1901), .B(n1472), .Z(n2081) );
  XOR U2083 ( .A(n2083), .B(n1685), .Z(o[712]) );
  XOR U2084 ( .A(n2084), .B(round_reg[320]), .Z(n1685) );
  NOR U2085 ( .A(n1904), .B(n1476), .Z(n2083) );
  XOR U2086 ( .A(n2085), .B(n1692), .Z(o[711]) );
  XNOR U2087 ( .A(n2086), .B(round_reg[383]), .Z(n1692) );
  XOR U2088 ( .A(n2087), .B(n1695), .Z(o[710]) );
  XOR U2089 ( .A(n2088), .B(round_reg[382]), .Z(n1695) );
  ANDN U2090 ( .A(n1910), .B(n1484), .Z(n2087) );
  IV U2091 ( .A(n2089), .Z(n1910) );
  XNOR U2092 ( .A(n2090), .B(n2091), .Z(o[70]) );
  AND U2093 ( .A(n2092), .B(n2093), .Z(n2090) );
  XOR U2094 ( .A(n2094), .B(n1698), .Z(o[709]) );
  XOR U2095 ( .A(n2095), .B(round_reg[381]), .Z(n1698) );
  ANDN U2096 ( .A(n1913), .B(n1488), .Z(n2094) );
  IV U2097 ( .A(n2096), .Z(n1913) );
  XOR U2098 ( .A(n2097), .B(n1700), .Z(o[708]) );
  XOR U2099 ( .A(n2098), .B(round_reg[380]), .Z(n1700) );
  ANDN U2100 ( .A(n1916), .B(n1492), .Z(n2097) );
  IV U2101 ( .A(n2099), .Z(n1916) );
  XOR U2102 ( .A(n2100), .B(n1702), .Z(o[707]) );
  XOR U2103 ( .A(n2101), .B(round_reg[379]), .Z(n1702) );
  ANDN U2104 ( .A(n1919), .B(n1504), .Z(n2100) );
  IV U2105 ( .A(n2102), .Z(n1919) );
  XOR U2106 ( .A(n2103), .B(n1704), .Z(o[706]) );
  XOR U2107 ( .A(n2104), .B(round_reg[378]), .Z(n1704) );
  ANDN U2108 ( .A(n1922), .B(n1508), .Z(n2103) );
  IV U2109 ( .A(n2105), .Z(n1922) );
  XOR U2110 ( .A(n2106), .B(n1706), .Z(o[705]) );
  XOR U2111 ( .A(n2107), .B(round_reg[377]), .Z(n1706) );
  ANDN U2112 ( .A(n1929), .B(n1512), .Z(n2106) );
  IV U2113 ( .A(n2108), .Z(n1929) );
  XOR U2114 ( .A(n2109), .B(n1708), .Z(o[704]) );
  XOR U2115 ( .A(n2110), .B(round_reg[376]), .Z(n1708) );
  XOR U2116 ( .A(n2111), .B(n1711), .Z(o[703]) );
  XOR U2117 ( .A(n2112), .B(round_reg[301]), .Z(n1711) );
  NOR U2118 ( .A(n1237), .B(n1236), .Z(n2111) );
  XNOR U2119 ( .A(n2113), .B(round_reg[1534]), .Z(n1236) );
  XNOR U2120 ( .A(n2114), .B(round_reg[1145]), .Z(n1237) );
  XOR U2121 ( .A(n2115), .B(n1714), .Z(o[702]) );
  XOR U2122 ( .A(n2116), .B(round_reg[300]), .Z(n1714) );
  NOR U2123 ( .A(n1241), .B(n1240), .Z(n2115) );
  XOR U2124 ( .A(n2117), .B(round_reg[1533]), .Z(n1240) );
  XNOR U2125 ( .A(n2118), .B(round_reg[1144]), .Z(n1241) );
  XOR U2126 ( .A(n2119), .B(n1721), .Z(o[701]) );
  XOR U2127 ( .A(n2120), .B(round_reg[299]), .Z(n1721) );
  NOR U2128 ( .A(n1245), .B(n1244), .Z(n2119) );
  XOR U2129 ( .A(n2121), .B(round_reg[1532]), .Z(n1244) );
  XNOR U2130 ( .A(n2122), .B(round_reg[1143]), .Z(n1245) );
  XOR U2131 ( .A(n2123), .B(n1941), .Z(o[700]) );
  XOR U2132 ( .A(n2124), .B(round_reg[298]), .Z(n1941) );
  NOR U2133 ( .A(n1249), .B(n1248), .Z(n2123) );
  XOR U2134 ( .A(n2125), .B(round_reg[1531]), .Z(n1248) );
  XNOR U2135 ( .A(n2126), .B(round_reg[1142]), .Z(n1249) );
  XNOR U2136 ( .A(n2127), .B(n2092), .Z(o[6]) );
  AND U2137 ( .A(n2128), .B(n2129), .Z(n2127) );
  XNOR U2138 ( .A(n2130), .B(n2131), .Z(o[69]) );
  AND U2139 ( .A(n2132), .B(n2133), .Z(n2130) );
  XOR U2140 ( .A(n2134), .B(n1944), .Z(o[699]) );
  XOR U2141 ( .A(n2135), .B(round_reg[297]), .Z(n1944) );
  NOR U2142 ( .A(n1253), .B(n1252), .Z(n2134) );
  XOR U2143 ( .A(n2136), .B(round_reg[1530]), .Z(n1252) );
  XNOR U2144 ( .A(n2137), .B(round_reg[1141]), .Z(n1253) );
  XOR U2145 ( .A(n2138), .B(n1947), .Z(o[698]) );
  XOR U2146 ( .A(n2139), .B(round_reg[296]), .Z(n1947) );
  ANDN U2147 ( .A(n1256), .B(n1257), .Z(n2138) );
  XNOR U2148 ( .A(n2140), .B(round_reg[1140]), .Z(n1257) );
  XNOR U2149 ( .A(n2141), .B(round_reg[1529]), .Z(n1256) );
  XOR U2150 ( .A(n2142), .B(n1950), .Z(o[697]) );
  XOR U2151 ( .A(n2143), .B(round_reg[295]), .Z(n1950) );
  ANDN U2152 ( .A(n1260), .B(n1261), .Z(n2142) );
  XNOR U2153 ( .A(n2144), .B(round_reg[1139]), .Z(n1261) );
  XNOR U2154 ( .A(n2145), .B(round_reg[1528]), .Z(n1260) );
  XOR U2155 ( .A(n2146), .B(n1953), .Z(o[696]) );
  XOR U2156 ( .A(n2147), .B(round_reg[294]), .Z(n1953) );
  ANDN U2157 ( .A(n1264), .B(n1265), .Z(n2146) );
  XNOR U2158 ( .A(n2148), .B(round_reg[1138]), .Z(n1265) );
  XNOR U2159 ( .A(n2149), .B(round_reg[1527]), .Z(n1264) );
  XOR U2160 ( .A(n2150), .B(n1960), .Z(o[695]) );
  XOR U2161 ( .A(n2151), .B(round_reg[293]), .Z(n1960) );
  ANDN U2162 ( .A(n1268), .B(n1269), .Z(n2150) );
  XNOR U2163 ( .A(n2152), .B(round_reg[1137]), .Z(n1269) );
  XNOR U2164 ( .A(n2153), .B(round_reg[1526]), .Z(n1268) );
  XOR U2165 ( .A(n2154), .B(n1963), .Z(o[694]) );
  XOR U2166 ( .A(n2155), .B(round_reg[292]), .Z(n1963) );
  ANDN U2167 ( .A(n1272), .B(n1273), .Z(n2154) );
  XNOR U2168 ( .A(n2156), .B(round_reg[1136]), .Z(n1273) );
  XNOR U2169 ( .A(n2157), .B(round_reg[1525]), .Z(n1272) );
  XOR U2170 ( .A(n2158), .B(n1966), .Z(o[693]) );
  XOR U2171 ( .A(n2159), .B(round_reg[291]), .Z(n1966) );
  ANDN U2172 ( .A(n1280), .B(n1281), .Z(n2158) );
  XNOR U2173 ( .A(n2160), .B(round_reg[1135]), .Z(n1281) );
  XNOR U2174 ( .A(n2161), .B(round_reg[1524]), .Z(n1280) );
  XOR U2175 ( .A(n2162), .B(n1969), .Z(o[692]) );
  XOR U2176 ( .A(n2163), .B(round_reg[290]), .Z(n1969) );
  ANDN U2177 ( .A(n1284), .B(n1285), .Z(n2162) );
  XNOR U2178 ( .A(n2164), .B(round_reg[1134]), .Z(n1285) );
  XNOR U2179 ( .A(n2165), .B(round_reg[1523]), .Z(n1284) );
  XOR U2180 ( .A(n2166), .B(n1972), .Z(o[691]) );
  XOR U2181 ( .A(n2167), .B(round_reg[289]), .Z(n1972) );
  ANDN U2182 ( .A(n1288), .B(n1289), .Z(n2166) );
  XNOR U2183 ( .A(n2168), .B(round_reg[1133]), .Z(n1289) );
  XNOR U2184 ( .A(n2169), .B(round_reg[1522]), .Z(n1288) );
  XOR U2185 ( .A(n2170), .B(n1975), .Z(o[690]) );
  XOR U2186 ( .A(n2171), .B(round_reg[288]), .Z(n1975) );
  ANDN U2187 ( .A(n1292), .B(n1293), .Z(n2170) );
  XOR U2188 ( .A(n2172), .B(round_reg[1132]), .Z(n1293) );
  XNOR U2189 ( .A(n2173), .B(round_reg[1521]), .Z(n1292) );
  XNOR U2190 ( .A(n2174), .B(n2175), .Z(o[68]) );
  AND U2191 ( .A(n2176), .B(n2177), .Z(n2174) );
  XOR U2192 ( .A(n2178), .B(n1761), .Z(o[689]) );
  XOR U2193 ( .A(n2179), .B(round_reg[287]), .Z(n1761) );
  ANDN U2194 ( .A(n1296), .B(n1297), .Z(n2178) );
  XOR U2195 ( .A(n2180), .B(round_reg[1131]), .Z(n1297) );
  XNOR U2196 ( .A(n2181), .B(round_reg[1520]), .Z(n1296) );
  XOR U2197 ( .A(n2182), .B(n1764), .Z(o[688]) );
  XOR U2198 ( .A(n2183), .B(round_reg[286]), .Z(n1764) );
  ANDN U2199 ( .A(n1300), .B(n1301), .Z(n2182) );
  XNOR U2200 ( .A(n2184), .B(round_reg[1130]), .Z(n1301) );
  XNOR U2201 ( .A(n2185), .B(round_reg[1519]), .Z(n1300) );
  XOR U2202 ( .A(n2186), .B(n1767), .Z(o[687]) );
  XOR U2203 ( .A(n2187), .B(round_reg[285]), .Z(n1767) );
  ANDN U2204 ( .A(n1304), .B(n1305), .Z(n2186) );
  XNOR U2205 ( .A(n2188), .B(round_reg[1129]), .Z(n1305) );
  XNOR U2206 ( .A(n2189), .B(round_reg[1518]), .Z(n1304) );
  XOR U2207 ( .A(n2190), .B(n1770), .Z(o[686]) );
  XOR U2208 ( .A(n2191), .B(round_reg[284]), .Z(n1770) );
  ANDN U2209 ( .A(n1308), .B(n1309), .Z(n2190) );
  XNOR U2210 ( .A(n2192), .B(round_reg[1128]), .Z(n1309) );
  XNOR U2211 ( .A(n2193), .B(round_reg[1517]), .Z(n1308) );
  XOR U2212 ( .A(n2194), .B(n1773), .Z(o[685]) );
  XOR U2213 ( .A(n2195), .B(round_reg[283]), .Z(n1773) );
  ANDN U2214 ( .A(n1312), .B(n1313), .Z(n2194) );
  XNOR U2215 ( .A(n2196), .B(round_reg[1127]), .Z(n1313) );
  XNOR U2216 ( .A(n2197), .B(round_reg[1516]), .Z(n1312) );
  XOR U2217 ( .A(n2198), .B(n1776), .Z(o[684]) );
  XOR U2218 ( .A(n2199), .B(round_reg[282]), .Z(n1776) );
  ANDN U2219 ( .A(n1316), .B(n1317), .Z(n2198) );
  XNOR U2220 ( .A(n2200), .B(round_reg[1126]), .Z(n1317) );
  XNOR U2221 ( .A(n2201), .B(round_reg[1515]), .Z(n1316) );
  XOR U2222 ( .A(n2202), .B(n1779), .Z(o[683]) );
  XOR U2223 ( .A(n2203), .B(round_reg[281]), .Z(n1779) );
  ANDN U2224 ( .A(n1324), .B(n1325), .Z(n2202) );
  XNOR U2225 ( .A(n2204), .B(round_reg[1125]), .Z(n1325) );
  XNOR U2226 ( .A(n2205), .B(round_reg[1514]), .Z(n1324) );
  XOR U2227 ( .A(n2206), .B(n1782), .Z(o[682]) );
  XOR U2228 ( .A(n2207), .B(round_reg[280]), .Z(n1782) );
  ANDN U2229 ( .A(n1328), .B(n1329), .Z(n2206) );
  XNOR U2230 ( .A(n2208), .B(round_reg[1124]), .Z(n1329) );
  XNOR U2231 ( .A(n2209), .B(round_reg[1513]), .Z(n1328) );
  XOR U2232 ( .A(n2210), .B(n1789), .Z(o[681]) );
  XOR U2233 ( .A(n2211), .B(round_reg[279]), .Z(n1789) );
  ANDN U2234 ( .A(n1332), .B(n1333), .Z(n2210) );
  XOR U2235 ( .A(n2212), .B(round_reg[1123]), .Z(n1333) );
  XNOR U2236 ( .A(n2213), .B(round_reg[1512]), .Z(n1332) );
  XOR U2237 ( .A(n2214), .B(n1792), .Z(o[680]) );
  XOR U2238 ( .A(n2215), .B(round_reg[278]), .Z(n1792) );
  ANDN U2239 ( .A(n1336), .B(n1337), .Z(n2214) );
  XNOR U2240 ( .A(n2216), .B(round_reg[1122]), .Z(n1337) );
  XNOR U2241 ( .A(n2217), .B(round_reg[1511]), .Z(n1336) );
  XNOR U2242 ( .A(n2218), .B(n2219), .Z(o[67]) );
  AND U2243 ( .A(n2220), .B(n2221), .Z(n2218) );
  XOR U2244 ( .A(n2222), .B(n1795), .Z(o[679]) );
  XOR U2245 ( .A(n2223), .B(round_reg[277]), .Z(n1795) );
  ANDN U2246 ( .A(n1340), .B(n1341), .Z(n2222) );
  XNOR U2247 ( .A(n2224), .B(round_reg[1121]), .Z(n1341) );
  XNOR U2248 ( .A(n2225), .B(round_reg[1510]), .Z(n1340) );
  XOR U2249 ( .A(n2226), .B(n1798), .Z(o[678]) );
  XOR U2250 ( .A(n2227), .B(round_reg[276]), .Z(n1798) );
  ANDN U2251 ( .A(n1344), .B(n1345), .Z(n2226) );
  XNOR U2252 ( .A(n2228), .B(round_reg[1120]), .Z(n1345) );
  XNOR U2253 ( .A(n2229), .B(round_reg[1509]), .Z(n1344) );
  XOR U2254 ( .A(n2230), .B(n1801), .Z(o[677]) );
  XOR U2255 ( .A(n2231), .B(round_reg[275]), .Z(n1801) );
  ANDN U2256 ( .A(n1348), .B(n1349), .Z(n2230) );
  XNOR U2257 ( .A(n2232), .B(round_reg[1119]), .Z(n1349) );
  XNOR U2258 ( .A(n2233), .B(round_reg[1508]), .Z(n1348) );
  XOR U2259 ( .A(n2234), .B(n1804), .Z(o[676]) );
  XOR U2260 ( .A(n2235), .B(round_reg[274]), .Z(n1804) );
  ANDN U2261 ( .A(n1352), .B(n1353), .Z(n2234) );
  XNOR U2262 ( .A(n2236), .B(round_reg[1118]), .Z(n1353) );
  XNOR U2263 ( .A(n2237), .B(round_reg[1507]), .Z(n1352) );
  XOR U2264 ( .A(n2238), .B(n1807), .Z(o[675]) );
  XOR U2265 ( .A(n2239), .B(round_reg[273]), .Z(n1807) );
  ANDN U2266 ( .A(n1356), .B(n1357), .Z(n2238) );
  XNOR U2267 ( .A(n2240), .B(round_reg[1117]), .Z(n1357) );
  XNOR U2268 ( .A(n2241), .B(round_reg[1506]), .Z(n1356) );
  XOR U2269 ( .A(n2242), .B(n1810), .Z(o[674]) );
  XOR U2270 ( .A(n2243), .B(round_reg[272]), .Z(n1810) );
  ANDN U2271 ( .A(n1360), .B(n1361), .Z(n2242) );
  XNOR U2272 ( .A(n2244), .B(round_reg[1116]), .Z(n1361) );
  XNOR U2273 ( .A(n2245), .B(round_reg[1505]), .Z(n1360) );
  XOR U2274 ( .A(n2246), .B(n1813), .Z(o[673]) );
  XOR U2275 ( .A(n2247), .B(round_reg[271]), .Z(n1813) );
  ANDN U2276 ( .A(n1368), .B(n1369), .Z(n2246) );
  XNOR U2277 ( .A(n2248), .B(round_reg[1115]), .Z(n1369) );
  XOR U2278 ( .A(n2249), .B(round_reg[1504]), .Z(n1368) );
  XOR U2279 ( .A(n2250), .B(n1816), .Z(o[672]) );
  XOR U2280 ( .A(n2251), .B(round_reg[270]), .Z(n1816) );
  ANDN U2281 ( .A(n1372), .B(n1373), .Z(n2250) );
  XNOR U2282 ( .A(n2252), .B(round_reg[1114]), .Z(n1373) );
  XOR U2283 ( .A(n2253), .B(round_reg[1503]), .Z(n1372) );
  XOR U2284 ( .A(n2254), .B(n1827), .Z(o[671]) );
  XOR U2285 ( .A(n2255), .B(round_reg[269]), .Z(n1827) );
  ANDN U2286 ( .A(n1376), .B(n1377), .Z(n2254) );
  XNOR U2287 ( .A(n2256), .B(round_reg[1113]), .Z(n1377) );
  XOR U2288 ( .A(n2257), .B(round_reg[1502]), .Z(n1376) );
  XOR U2289 ( .A(n2258), .B(n1830), .Z(o[670]) );
  XOR U2290 ( .A(n2259), .B(round_reg[268]), .Z(n1830) );
  ANDN U2291 ( .A(n1380), .B(n1381), .Z(n2258) );
  XNOR U2292 ( .A(n2260), .B(round_reg[1112]), .Z(n1381) );
  XOR U2293 ( .A(n2261), .B(round_reg[1501]), .Z(n1380) );
  XNOR U2294 ( .A(n2262), .B(n2263), .Z(o[66]) );
  AND U2295 ( .A(n2264), .B(n2265), .Z(n2262) );
  XOR U2296 ( .A(n2266), .B(n1833), .Z(o[669]) );
  XOR U2297 ( .A(n2267), .B(round_reg[267]), .Z(n1833) );
  ANDN U2298 ( .A(n1384), .B(n1385), .Z(n2266) );
  XNOR U2299 ( .A(n2268), .B(round_reg[1111]), .Z(n1385) );
  XOR U2300 ( .A(n2269), .B(round_reg[1500]), .Z(n1384) );
  XOR U2301 ( .A(n2270), .B(n1836), .Z(o[668]) );
  XOR U2302 ( .A(n2271), .B(round_reg[266]), .Z(n1836) );
  ANDN U2303 ( .A(n1388), .B(n1389), .Z(n2270) );
  XNOR U2304 ( .A(n2272), .B(round_reg[1110]), .Z(n1389) );
  XNOR U2305 ( .A(n2273), .B(round_reg[1499]), .Z(n1388) );
  XOR U2306 ( .A(n2274), .B(n2029), .Z(o[667]) );
  XOR U2307 ( .A(n2275), .B(round_reg[265]), .Z(n2029) );
  ANDN U2308 ( .A(n1392), .B(n1393), .Z(n2274) );
  XNOR U2309 ( .A(n2276), .B(round_reg[1109]), .Z(n1393) );
  XNOR U2310 ( .A(n2277), .B(round_reg[1498]), .Z(n1392) );
  XOR U2311 ( .A(n2278), .B(n2032), .Z(o[666]) );
  XOR U2312 ( .A(n2279), .B(round_reg[264]), .Z(n2032) );
  ANDN U2313 ( .A(n1396), .B(n1397), .Z(n2278) );
  XNOR U2314 ( .A(n2280), .B(round_reg[1108]), .Z(n1397) );
  XNOR U2315 ( .A(n2281), .B(round_reg[1497]), .Z(n1396) );
  XOR U2316 ( .A(n2282), .B(n2037), .Z(o[665]) );
  XOR U2317 ( .A(n2283), .B(round_reg[263]), .Z(n2037) );
  ANDN U2318 ( .A(n1400), .B(n1401), .Z(n2282) );
  XNOR U2319 ( .A(n2284), .B(round_reg[1107]), .Z(n1401) );
  XNOR U2320 ( .A(n2285), .B(round_reg[1496]), .Z(n1400) );
  XOR U2321 ( .A(n2286), .B(n2040), .Z(o[664]) );
  XOR U2322 ( .A(n2287), .B(round_reg[262]), .Z(n2040) );
  ANDN U2323 ( .A(n1404), .B(n1405), .Z(n2286) );
  XNOR U2324 ( .A(n2288), .B(round_reg[1106]), .Z(n1405) );
  XNOR U2325 ( .A(n2289), .B(round_reg[1495]), .Z(n1404) );
  XOR U2326 ( .A(n2290), .B(n1851), .Z(o[663]) );
  XOR U2327 ( .A(n2291), .B(round_reg[261]), .Z(n1851) );
  ANDN U2328 ( .A(n1412), .B(n1413), .Z(n2290) );
  XNOR U2329 ( .A(n2292), .B(round_reg[1105]), .Z(n1413) );
  XNOR U2330 ( .A(n2293), .B(round_reg[1494]), .Z(n1412) );
  XOR U2331 ( .A(n2294), .B(n2045), .Z(o[662]) );
  XOR U2332 ( .A(n2295), .B(round_reg[260]), .Z(n2045) );
  ANDN U2333 ( .A(n1416), .B(n1417), .Z(n2294) );
  XNOR U2334 ( .A(n2296), .B(round_reg[1104]), .Z(n1417) );
  XNOR U2335 ( .A(n2297), .B(round_reg[1493]), .Z(n1416) );
  XOR U2336 ( .A(n2298), .B(n2048), .Z(o[661]) );
  XOR U2337 ( .A(n2299), .B(round_reg[259]), .Z(n2048) );
  ANDN U2338 ( .A(n1420), .B(n1421), .Z(n2298) );
  XNOR U2339 ( .A(n2300), .B(round_reg[1103]), .Z(n1421) );
  XNOR U2340 ( .A(n2301), .B(round_reg[1492]), .Z(n1420) );
  XOR U2341 ( .A(n2302), .B(n2051), .Z(o[660]) );
  XOR U2342 ( .A(n2303), .B(round_reg[258]), .Z(n2051) );
  ANDN U2343 ( .A(n1424), .B(n1425), .Z(n2302) );
  XNOR U2344 ( .A(n2304), .B(round_reg[1102]), .Z(n1425) );
  XNOR U2345 ( .A(n2305), .B(round_reg[1491]), .Z(n1424) );
  XNOR U2346 ( .A(n2306), .B(n2307), .Z(o[65]) );
  AND U2347 ( .A(n2308), .B(n2309), .Z(n2306) );
  XOR U2348 ( .A(n2310), .B(n2054), .Z(o[659]) );
  XOR U2349 ( .A(n2311), .B(round_reg[257]), .Z(n2054) );
  ANDN U2350 ( .A(n1428), .B(n1429), .Z(n2310) );
  XNOR U2351 ( .A(n2312), .B(round_reg[1101]), .Z(n1429) );
  XNOR U2352 ( .A(n2313), .B(round_reg[1490]), .Z(n1428) );
  XOR U2353 ( .A(n2314), .B(n2057), .Z(o[658]) );
  XOR U2354 ( .A(n2315), .B(round_reg[256]), .Z(n2057) );
  ANDN U2355 ( .A(n1432), .B(n1433), .Z(n2314) );
  XNOR U2356 ( .A(n2316), .B(round_reg[1100]), .Z(n1433) );
  XNOR U2357 ( .A(n2317), .B(round_reg[1489]), .Z(n1432) );
  XOR U2358 ( .A(n2318), .B(n2060), .Z(o[657]) );
  XOR U2359 ( .A(n2319), .B(round_reg[319]), .Z(n2060) );
  ANDN U2360 ( .A(n1436), .B(n1437), .Z(n2318) );
  XNOR U2361 ( .A(n2320), .B(round_reg[1099]), .Z(n1437) );
  XNOR U2362 ( .A(n2321), .B(round_reg[1488]), .Z(n1436) );
  XOR U2363 ( .A(n2322), .B(n2063), .Z(o[656]) );
  XOR U2364 ( .A(n2323), .B(round_reg[318]), .Z(n2063) );
  ANDN U2365 ( .A(n1440), .B(n1441), .Z(n2322) );
  XNOR U2366 ( .A(n2324), .B(round_reg[1098]), .Z(n1441) );
  XNOR U2367 ( .A(n2325), .B(round_reg[1487]), .Z(n1440) );
  XOR U2368 ( .A(n2326), .B(n2068), .Z(o[655]) );
  XOR U2369 ( .A(n2327), .B(round_reg[317]), .Z(n2068) );
  ANDN U2370 ( .A(n1444), .B(n1445), .Z(n2326) );
  XNOR U2371 ( .A(n2328), .B(round_reg[1097]), .Z(n1445) );
  XNOR U2372 ( .A(n2329), .B(round_reg[1486]), .Z(n1444) );
  XOR U2373 ( .A(n2330), .B(n2071), .Z(o[654]) );
  XOR U2374 ( .A(n2331), .B(round_reg[316]), .Z(n2071) );
  ANDN U2375 ( .A(n1448), .B(n1449), .Z(n2330) );
  XNOR U2376 ( .A(n2332), .B(round_reg[1096]), .Z(n1449) );
  XNOR U2377 ( .A(n2333), .B(round_reg[1485]), .Z(n1448) );
  XOR U2378 ( .A(n2334), .B(n2074), .Z(o[653]) );
  XOR U2379 ( .A(n2335), .B(round_reg[315]), .Z(n2074) );
  ANDN U2380 ( .A(n1456), .B(n1457), .Z(n2334) );
  XNOR U2381 ( .A(n2336), .B(round_reg[1095]), .Z(n1457) );
  XNOR U2382 ( .A(n2337), .B(round_reg[1484]), .Z(n1456) );
  XOR U2383 ( .A(n2338), .B(n1888), .Z(o[652]) );
  XOR U2384 ( .A(n2339), .B(round_reg[314]), .Z(n1888) );
  ANDN U2385 ( .A(n1460), .B(n1461), .Z(n2338) );
  XNOR U2386 ( .A(n2340), .B(round_reg[1094]), .Z(n1461) );
  XNOR U2387 ( .A(n2341), .B(round_reg[1483]), .Z(n1460) );
  XOR U2388 ( .A(n2342), .B(n1895), .Z(o[651]) );
  XOR U2389 ( .A(n2343), .B(round_reg[313]), .Z(n1895) );
  ANDN U2390 ( .A(n1464), .B(n1465), .Z(n2342) );
  XNOR U2391 ( .A(n2344), .B(round_reg[1093]), .Z(n1465) );
  XNOR U2392 ( .A(n2345), .B(round_reg[1482]), .Z(n1464) );
  XOR U2393 ( .A(n2346), .B(n1898), .Z(o[650]) );
  XOR U2394 ( .A(n2347), .B(round_reg[312]), .Z(n1898) );
  ANDN U2395 ( .A(n1468), .B(n1469), .Z(n2346) );
  XNOR U2396 ( .A(n2348), .B(round_reg[1092]), .Z(n1469) );
  XNOR U2397 ( .A(n2349), .B(round_reg[1481]), .Z(n1468) );
  XNOR U2398 ( .A(n2350), .B(n2351), .Z(o[64]) );
  XOR U2399 ( .A(n2354), .B(n1901), .Z(o[649]) );
  XOR U2400 ( .A(n2355), .B(round_reg[311]), .Z(n1901) );
  ANDN U2401 ( .A(n1472), .B(n1473), .Z(n2354) );
  XNOR U2402 ( .A(n2356), .B(round_reg[1091]), .Z(n1473) );
  XNOR U2403 ( .A(n2357), .B(round_reg[1480]), .Z(n1472) );
  XOR U2404 ( .A(n2358), .B(n1904), .Z(o[648]) );
  XOR U2405 ( .A(n2359), .B(round_reg[310]), .Z(n1904) );
  ANDN U2406 ( .A(n1476), .B(n1477), .Z(n2358) );
  XNOR U2407 ( .A(n2360), .B(round_reg[1090]), .Z(n1477) );
  XNOR U2408 ( .A(n2361), .B(round_reg[1479]), .Z(n1476) );
  XOR U2409 ( .A(n2362), .B(n1907), .Z(o[647]) );
  XOR U2410 ( .A(n2363), .B(round_reg[309]), .Z(n1907) );
  ANDN U2411 ( .A(n1480), .B(n1481), .Z(n2362) );
  XNOR U2412 ( .A(n2364), .B(round_reg[1089]), .Z(n1481) );
  XNOR U2413 ( .A(n2365), .B(round_reg[1478]), .Z(n1480) );
  XOR U2414 ( .A(n2366), .B(n2089), .Z(o[646]) );
  XOR U2415 ( .A(n2367), .B(round_reg[308]), .Z(n2089) );
  ANDN U2416 ( .A(n1484), .B(n1485), .Z(n2366) );
  XNOR U2417 ( .A(n2368), .B(round_reg[1088]), .Z(n1485) );
  XNOR U2418 ( .A(n2369), .B(round_reg[1477]), .Z(n1484) );
  XOR U2419 ( .A(n2370), .B(n2096), .Z(o[645]) );
  XOR U2420 ( .A(n2371), .B(round_reg[307]), .Z(n2096) );
  ANDN U2421 ( .A(n1488), .B(n1489), .Z(n2370) );
  XNOR U2422 ( .A(n2372), .B(round_reg[1151]), .Z(n1489) );
  XNOR U2423 ( .A(n2373), .B(round_reg[1476]), .Z(n1488) );
  XOR U2424 ( .A(n2374), .B(n2099), .Z(o[644]) );
  XOR U2425 ( .A(n2375), .B(round_reg[306]), .Z(n2099) );
  ANDN U2426 ( .A(n1492), .B(n1493), .Z(n2374) );
  XNOR U2427 ( .A(n2376), .B(round_reg[1150]), .Z(n1493) );
  XNOR U2428 ( .A(n2377), .B(round_reg[1475]), .Z(n1492) );
  XOR U2429 ( .A(n2378), .B(n2102), .Z(o[643]) );
  XOR U2430 ( .A(n2379), .B(round_reg[305]), .Z(n2102) );
  ANDN U2431 ( .A(n1504), .B(n1505), .Z(n2378) );
  XNOR U2432 ( .A(n2380), .B(round_reg[1149]), .Z(n1505) );
  XNOR U2433 ( .A(n2381), .B(round_reg[1474]), .Z(n1504) );
  XOR U2434 ( .A(n2382), .B(n2105), .Z(o[642]) );
  XOR U2435 ( .A(n2383), .B(round_reg[304]), .Z(n2105) );
  ANDN U2436 ( .A(n1508), .B(n1509), .Z(n2382) );
  XNOR U2437 ( .A(n2384), .B(round_reg[1148]), .Z(n1509) );
  XNOR U2438 ( .A(n2385), .B(round_reg[1473]), .Z(n1508) );
  XOR U2439 ( .A(n2386), .B(n2108), .Z(o[641]) );
  XOR U2440 ( .A(n2387), .B(round_reg[303]), .Z(n2108) );
  ANDN U2441 ( .A(n1512), .B(n1513), .Z(n2386) );
  XNOR U2442 ( .A(n2388), .B(round_reg[1147]), .Z(n1513) );
  XNOR U2443 ( .A(n2389), .B(round_reg[1472]), .Z(n1512) );
  XOR U2444 ( .A(n2390), .B(n1932), .Z(o[640]) );
  XOR U2445 ( .A(n2391), .B(round_reg[302]), .Z(n1932) );
  ANDN U2446 ( .A(n1516), .B(n1517), .Z(n2390) );
  XNOR U2447 ( .A(n2392), .B(round_reg[1146]), .Z(n1517) );
  XNOR U2448 ( .A(n2393), .B(round_reg[1535]), .Z(n1516) );
  XNOR U2449 ( .A(n2394), .B(n2395), .Z(o[63]) );
  AND U2450 ( .A(n2396), .B(n2397), .Z(n2394) );
  XNOR U2451 ( .A(n2398), .B(n2399), .Z(o[639]) );
  AND U2452 ( .A(n2400), .B(n2401), .Z(n2398) );
  XNOR U2453 ( .A(n2402), .B(n2403), .Z(o[638]) );
  AND U2454 ( .A(n2404), .B(n2405), .Z(n2402) );
  XNOR U2455 ( .A(n2406), .B(n2407), .Z(o[637]) );
  AND U2456 ( .A(n2408), .B(n2409), .Z(n2406) );
  XNOR U2457 ( .A(n2410), .B(n2411), .Z(o[636]) );
  AND U2458 ( .A(n2412), .B(n2413), .Z(n2410) );
  XNOR U2459 ( .A(n2414), .B(n2415), .Z(o[635]) );
  AND U2460 ( .A(n2416), .B(n2417), .Z(n2414) );
  XNOR U2461 ( .A(n2418), .B(n2419), .Z(o[634]) );
  AND U2462 ( .A(n2420), .B(n2421), .Z(n2418) );
  XNOR U2463 ( .A(n2422), .B(n2423), .Z(o[633]) );
  AND U2464 ( .A(n2424), .B(n2425), .Z(n2422) );
  XNOR U2465 ( .A(n2426), .B(n2427), .Z(o[632]) );
  AND U2466 ( .A(n2428), .B(n2429), .Z(n2426) );
  XNOR U2467 ( .A(n2430), .B(n2431), .Z(o[631]) );
  AND U2468 ( .A(n2432), .B(n2433), .Z(n2430) );
  XNOR U2469 ( .A(n2434), .B(n2435), .Z(o[630]) );
  AND U2470 ( .A(n2436), .B(n2437), .Z(n2434) );
  XNOR U2471 ( .A(n2438), .B(n2439), .Z(o[62]) );
  AND U2472 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR U2473 ( .A(n2442), .B(n2443), .Z(o[629]) );
  AND U2474 ( .A(n2444), .B(n2445), .Z(n2442) );
  XNOR U2475 ( .A(n2446), .B(n2447), .Z(o[628]) );
  AND U2476 ( .A(n2448), .B(n2449), .Z(n2446) );
  XNOR U2477 ( .A(n2450), .B(n2451), .Z(o[627]) );
  AND U2478 ( .A(n2452), .B(n2453), .Z(n2450) );
  XNOR U2479 ( .A(n2454), .B(n2455), .Z(o[626]) );
  AND U2480 ( .A(n2456), .B(n2457), .Z(n2454) );
  XNOR U2481 ( .A(n2458), .B(n2459), .Z(o[625]) );
  AND U2482 ( .A(n2460), .B(n2461), .Z(n2458) );
  XNOR U2483 ( .A(n2462), .B(n2463), .Z(o[624]) );
  AND U2484 ( .A(n2464), .B(n2465), .Z(n2462) );
  XNOR U2485 ( .A(n2466), .B(n2467), .Z(o[623]) );
  AND U2486 ( .A(n2468), .B(n2469), .Z(n2466) );
  XNOR U2487 ( .A(n2470), .B(n2471), .Z(o[622]) );
  AND U2488 ( .A(n2472), .B(n2473), .Z(n2470) );
  XNOR U2489 ( .A(n2474), .B(n2475), .Z(o[621]) );
  AND U2490 ( .A(n2476), .B(n2477), .Z(n2474) );
  XNOR U2491 ( .A(n2478), .B(n2479), .Z(o[620]) );
  AND U2492 ( .A(n2480), .B(n2481), .Z(n2478) );
  XNOR U2493 ( .A(n2482), .B(n2483), .Z(o[61]) );
  AND U2494 ( .A(n2484), .B(n2485), .Z(n2482) );
  XNOR U2495 ( .A(n2486), .B(n2487), .Z(o[619]) );
  AND U2496 ( .A(n2488), .B(n2489), .Z(n2486) );
  XNOR U2497 ( .A(n2490), .B(n2491), .Z(o[618]) );
  AND U2498 ( .A(n2492), .B(n2493), .Z(n2490) );
  XNOR U2499 ( .A(n2494), .B(n2495), .Z(o[617]) );
  AND U2500 ( .A(n2496), .B(n2497), .Z(n2494) );
  XNOR U2501 ( .A(n2498), .B(n2499), .Z(o[616]) );
  AND U2502 ( .A(n2500), .B(n2501), .Z(n2498) );
  XNOR U2503 ( .A(n2502), .B(n2503), .Z(o[615]) );
  AND U2504 ( .A(n2504), .B(n2505), .Z(n2502) );
  XNOR U2505 ( .A(n2506), .B(n2507), .Z(o[614]) );
  AND U2506 ( .A(n2508), .B(n2509), .Z(n2506) );
  XNOR U2507 ( .A(n2510), .B(n2511), .Z(o[613]) );
  AND U2508 ( .A(n2512), .B(n2513), .Z(n2510) );
  XNOR U2509 ( .A(n2514), .B(n2515), .Z(o[612]) );
  AND U2510 ( .A(n2516), .B(n2517), .Z(n2514) );
  XNOR U2511 ( .A(n2518), .B(n2519), .Z(o[611]) );
  AND U2512 ( .A(n2520), .B(n2521), .Z(n2518) );
  XNOR U2513 ( .A(n2522), .B(n2523), .Z(o[610]) );
  AND U2514 ( .A(n2524), .B(n2525), .Z(n2522) );
  XNOR U2515 ( .A(n2526), .B(n2527), .Z(o[60]) );
  AND U2516 ( .A(n2528), .B(n2529), .Z(n2526) );
  XNOR U2517 ( .A(n2530), .B(n2531), .Z(o[609]) );
  AND U2518 ( .A(n2532), .B(n2533), .Z(n2530) );
  XNOR U2519 ( .A(n2534), .B(n2535), .Z(o[608]) );
  AND U2520 ( .A(n2536), .B(n2537), .Z(n2534) );
  XNOR U2521 ( .A(n2538), .B(n2539), .Z(o[607]) );
  AND U2522 ( .A(n2540), .B(n2541), .Z(n2538) );
  XNOR U2523 ( .A(n2542), .B(n2543), .Z(o[606]) );
  AND U2524 ( .A(n2544), .B(n2545), .Z(n2542) );
  XNOR U2525 ( .A(n2546), .B(n2547), .Z(o[605]) );
  AND U2526 ( .A(n2548), .B(n2549), .Z(n2546) );
  XNOR U2527 ( .A(n2550), .B(n2551), .Z(o[604]) );
  AND U2528 ( .A(n2552), .B(n2553), .Z(n2550) );
  XNOR U2529 ( .A(n2554), .B(n2555), .Z(o[603]) );
  AND U2530 ( .A(n2556), .B(n2557), .Z(n2554) );
  XNOR U2531 ( .A(n2558), .B(n2559), .Z(o[602]) );
  AND U2532 ( .A(n2560), .B(n2561), .Z(n2558) );
  XNOR U2533 ( .A(n2562), .B(n2563), .Z(o[601]) );
  AND U2534 ( .A(n2564), .B(n2565), .Z(n2562) );
  XNOR U2535 ( .A(n2566), .B(n2567), .Z(o[600]) );
  AND U2536 ( .A(n2568), .B(n2569), .Z(n2566) );
  XNOR U2537 ( .A(n2570), .B(n2132), .Z(o[5]) );
  AND U2538 ( .A(n2571), .B(n2572), .Z(n2570) );
  XNOR U2539 ( .A(n2573), .B(n2574), .Z(o[59]) );
  AND U2540 ( .A(n2575), .B(n2576), .Z(n2573) );
  XNOR U2541 ( .A(n2577), .B(n2578), .Z(o[599]) );
  AND U2542 ( .A(n2579), .B(n2580), .Z(n2577) );
  XNOR U2543 ( .A(n2581), .B(n2582), .Z(o[598]) );
  AND U2544 ( .A(n2583), .B(n2584), .Z(n2581) );
  XNOR U2545 ( .A(n2585), .B(n2586), .Z(o[597]) );
  AND U2546 ( .A(n2587), .B(n2588), .Z(n2585) );
  XNOR U2547 ( .A(n2589), .B(n2590), .Z(o[596]) );
  AND U2548 ( .A(n2591), .B(n2592), .Z(n2589) );
  XNOR U2549 ( .A(n2593), .B(n2594), .Z(o[595]) );
  AND U2550 ( .A(n2595), .B(n2596), .Z(n2593) );
  XNOR U2551 ( .A(n2597), .B(n2598), .Z(o[594]) );
  AND U2552 ( .A(n2599), .B(n2600), .Z(n2597) );
  XNOR U2553 ( .A(n2601), .B(n2602), .Z(o[593]) );
  AND U2554 ( .A(n2603), .B(n2604), .Z(n2601) );
  XNOR U2555 ( .A(n2605), .B(n2606), .Z(o[592]) );
  AND U2556 ( .A(n2607), .B(n2608), .Z(n2605) );
  XNOR U2557 ( .A(n2609), .B(n2610), .Z(o[591]) );
  AND U2558 ( .A(n2611), .B(n2612), .Z(n2609) );
  XNOR U2559 ( .A(n2613), .B(n2614), .Z(o[590]) );
  AND U2560 ( .A(n2615), .B(n2616), .Z(n2613) );
  XNOR U2561 ( .A(n2617), .B(n2618), .Z(o[58]) );
  AND U2562 ( .A(n2619), .B(n2620), .Z(n2617) );
  XNOR U2563 ( .A(n2621), .B(n2622), .Z(o[589]) );
  AND U2564 ( .A(n2623), .B(n2624), .Z(n2621) );
  XNOR U2565 ( .A(n2625), .B(n2626), .Z(o[588]) );
  AND U2566 ( .A(n2627), .B(n2628), .Z(n2625) );
  XNOR U2567 ( .A(n2629), .B(n2630), .Z(o[587]) );
  AND U2568 ( .A(n2631), .B(n2632), .Z(n2629) );
  XNOR U2569 ( .A(n2633), .B(n2634), .Z(o[586]) );
  AND U2570 ( .A(n2635), .B(n2636), .Z(n2633) );
  XNOR U2571 ( .A(n2637), .B(n2638), .Z(o[585]) );
  AND U2572 ( .A(n2639), .B(n2640), .Z(n2637) );
  XNOR U2573 ( .A(n2641), .B(n2642), .Z(o[584]) );
  AND U2574 ( .A(n2643), .B(n2644), .Z(n2641) );
  XNOR U2575 ( .A(n2645), .B(n2646), .Z(o[583]) );
  AND U2576 ( .A(n2647), .B(n2648), .Z(n2645) );
  XNOR U2577 ( .A(n2649), .B(n2650), .Z(o[582]) );
  AND U2578 ( .A(n2651), .B(n2652), .Z(n2649) );
  XNOR U2579 ( .A(n2653), .B(n2654), .Z(o[581]) );
  AND U2580 ( .A(n2655), .B(n2656), .Z(n2653) );
  XNOR U2581 ( .A(n2657), .B(n2658), .Z(o[580]) );
  AND U2582 ( .A(n2659), .B(n2660), .Z(n2657) );
  XNOR U2583 ( .A(n2661), .B(n2662), .Z(o[57]) );
  AND U2584 ( .A(n2663), .B(n2664), .Z(n2661) );
  XNOR U2585 ( .A(n2665), .B(n2666), .Z(o[579]) );
  AND U2586 ( .A(n2667), .B(n2668), .Z(n2665) );
  XNOR U2587 ( .A(n2669), .B(n2670), .Z(o[578]) );
  AND U2588 ( .A(n2671), .B(n2672), .Z(n2669) );
  XNOR U2589 ( .A(n2673), .B(n2674), .Z(o[577]) );
  AND U2590 ( .A(n2675), .B(n2676), .Z(n2673) );
  XNOR U2591 ( .A(n2677), .B(n2678), .Z(o[576]) );
  AND U2592 ( .A(n2679), .B(n2680), .Z(n2677) );
  XNOR U2593 ( .A(n2681), .B(n2400), .Z(o[575]) );
  AND U2594 ( .A(n2682), .B(n2683), .Z(n2681) );
  XNOR U2595 ( .A(n2684), .B(n2404), .Z(o[574]) );
  AND U2596 ( .A(n2685), .B(n2686), .Z(n2684) );
  XNOR U2597 ( .A(n2687), .B(n2408), .Z(o[573]) );
  AND U2598 ( .A(n2688), .B(n2689), .Z(n2687) );
  XNOR U2599 ( .A(n2690), .B(n2412), .Z(o[572]) );
  AND U2600 ( .A(n2691), .B(n2692), .Z(n2690) );
  XNOR U2601 ( .A(n2693), .B(n2416), .Z(o[571]) );
  AND U2602 ( .A(n2694), .B(n2695), .Z(n2693) );
  XNOR U2603 ( .A(n2696), .B(n2420), .Z(o[570]) );
  AND U2604 ( .A(n2697), .B(n2698), .Z(n2696) );
  XNOR U2605 ( .A(n2699), .B(n2700), .Z(o[56]) );
  AND U2606 ( .A(n2701), .B(n2702), .Z(n2699) );
  XNOR U2607 ( .A(n2703), .B(n2424), .Z(o[569]) );
  AND U2608 ( .A(n2704), .B(n2705), .Z(n2703) );
  XNOR U2609 ( .A(n2706), .B(n2428), .Z(o[568]) );
  AND U2610 ( .A(n2707), .B(n2708), .Z(n2706) );
  XNOR U2611 ( .A(n2709), .B(n2432), .Z(o[567]) );
  AND U2612 ( .A(n2710), .B(n2711), .Z(n2709) );
  XNOR U2613 ( .A(n2712), .B(n2436), .Z(o[566]) );
  AND U2614 ( .A(n2713), .B(n2714), .Z(n2712) );
  XNOR U2615 ( .A(n2715), .B(n2444), .Z(o[565]) );
  AND U2616 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U2617 ( .A(n2718), .B(n2448), .Z(o[564]) );
  AND U2618 ( .A(n2719), .B(n2720), .Z(n2718) );
  XNOR U2619 ( .A(n2721), .B(n2452), .Z(o[563]) );
  AND U2620 ( .A(n2722), .B(n2723), .Z(n2721) );
  XNOR U2621 ( .A(n2724), .B(n2456), .Z(o[562]) );
  AND U2622 ( .A(n2725), .B(n2726), .Z(n2724) );
  XNOR U2623 ( .A(n2727), .B(n2460), .Z(o[561]) );
  AND U2624 ( .A(n2728), .B(n2729), .Z(n2727) );
  XNOR U2625 ( .A(n2730), .B(n2464), .Z(o[560]) );
  AND U2626 ( .A(n2731), .B(n2732), .Z(n2730) );
  XNOR U2627 ( .A(n2733), .B(n2734), .Z(o[55]) );
  AND U2628 ( .A(n2735), .B(n2736), .Z(n2733) );
  XNOR U2629 ( .A(n2737), .B(n2468), .Z(o[559]) );
  AND U2630 ( .A(n2738), .B(n2739), .Z(n2737) );
  XNOR U2631 ( .A(n2740), .B(n2472), .Z(o[558]) );
  AND U2632 ( .A(n2741), .B(n2742), .Z(n2740) );
  XNOR U2633 ( .A(n2743), .B(n2476), .Z(o[557]) );
  AND U2634 ( .A(n2744), .B(n2745), .Z(n2743) );
  XNOR U2635 ( .A(n2746), .B(n2480), .Z(o[556]) );
  AND U2636 ( .A(n2747), .B(n2748), .Z(n2746) );
  XNOR U2637 ( .A(n2749), .B(n2488), .Z(o[555]) );
  AND U2638 ( .A(n2750), .B(n2751), .Z(n2749) );
  XNOR U2639 ( .A(n2752), .B(n2492), .Z(o[554]) );
  XNOR U2640 ( .A(n2754), .B(n2496), .Z(o[553]) );
  XNOR U2641 ( .A(n2756), .B(n2500), .Z(o[552]) );
  XNOR U2642 ( .A(n2758), .B(n2504), .Z(o[551]) );
  XNOR U2643 ( .A(n2760), .B(n2508), .Z(o[550]) );
  XNOR U2644 ( .A(n2762), .B(n2763), .Z(o[54]) );
  AND U2645 ( .A(n2764), .B(n2765), .Z(n2762) );
  XNOR U2646 ( .A(n2766), .B(n2512), .Z(o[549]) );
  AND U2647 ( .A(n2767), .B(n2768), .Z(n2766) );
  XNOR U2648 ( .A(n2769), .B(n2516), .Z(o[548]) );
  AND U2649 ( .A(n2770), .B(n2771), .Z(n2769) );
  XNOR U2650 ( .A(n2772), .B(n2520), .Z(o[547]) );
  AND U2651 ( .A(n2773), .B(n2774), .Z(n2772) );
  XNOR U2652 ( .A(n2775), .B(n2524), .Z(o[546]) );
  AND U2653 ( .A(n2776), .B(n2777), .Z(n2775) );
  XNOR U2654 ( .A(n2778), .B(n2532), .Z(o[545]) );
  AND U2655 ( .A(n2779), .B(n2780), .Z(n2778) );
  XNOR U2656 ( .A(n2781), .B(n2536), .Z(o[544]) );
  AND U2657 ( .A(n2782), .B(n2783), .Z(n2781) );
  XNOR U2658 ( .A(n2784), .B(n2540), .Z(o[543]) );
  AND U2659 ( .A(n2785), .B(n2786), .Z(n2784) );
  XNOR U2660 ( .A(n2787), .B(n2544), .Z(o[542]) );
  AND U2661 ( .A(n2788), .B(n2789), .Z(n2787) );
  XNOR U2662 ( .A(n2790), .B(n2548), .Z(o[541]) );
  AND U2663 ( .A(n2791), .B(n2792), .Z(n2790) );
  XNOR U2664 ( .A(n2793), .B(n2552), .Z(o[540]) );
  AND U2665 ( .A(n2794), .B(n2795), .Z(n2793) );
  XNOR U2666 ( .A(n2796), .B(n2797), .Z(o[53]) );
  AND U2667 ( .A(n2798), .B(n2799), .Z(n2796) );
  XNOR U2668 ( .A(n2800), .B(n2556), .Z(o[539]) );
  AND U2669 ( .A(n2801), .B(n2802), .Z(n2800) );
  XNOR U2670 ( .A(n2803), .B(n2560), .Z(o[538]) );
  AND U2671 ( .A(n2804), .B(n2805), .Z(n2803) );
  XNOR U2672 ( .A(n2806), .B(n2564), .Z(o[537]) );
  AND U2673 ( .A(n2807), .B(n2808), .Z(n2806) );
  XNOR U2674 ( .A(n2809), .B(n2568), .Z(o[536]) );
  AND U2675 ( .A(n2810), .B(n2811), .Z(n2809) );
  XNOR U2676 ( .A(n2812), .B(n2579), .Z(o[535]) );
  AND U2677 ( .A(n2813), .B(n2814), .Z(n2812) );
  XNOR U2678 ( .A(n2815), .B(n2583), .Z(o[534]) );
  AND U2679 ( .A(n2816), .B(n2817), .Z(n2815) );
  XNOR U2680 ( .A(n2818), .B(n2587), .Z(o[533]) );
  AND U2681 ( .A(n2819), .B(n2820), .Z(n2818) );
  XNOR U2682 ( .A(n2821), .B(n2591), .Z(o[532]) );
  AND U2683 ( .A(n2822), .B(n2823), .Z(n2821) );
  XNOR U2684 ( .A(n2824), .B(n2595), .Z(o[531]) );
  AND U2685 ( .A(n2825), .B(n2826), .Z(n2824) );
  XNOR U2686 ( .A(n2827), .B(n2599), .Z(o[530]) );
  AND U2687 ( .A(n2828), .B(n2829), .Z(n2827) );
  XNOR U2688 ( .A(n2830), .B(n2831), .Z(o[52]) );
  AND U2689 ( .A(n2832), .B(n2833), .Z(n2830) );
  XNOR U2690 ( .A(n2834), .B(n2603), .Z(o[529]) );
  AND U2691 ( .A(n2835), .B(n2836), .Z(n2834) );
  XNOR U2692 ( .A(n2837), .B(n2607), .Z(o[528]) );
  AND U2693 ( .A(n2838), .B(n2839), .Z(n2837) );
  XNOR U2694 ( .A(n2840), .B(n2611), .Z(o[527]) );
  AND U2695 ( .A(n2841), .B(n2842), .Z(n2840) );
  XNOR U2696 ( .A(n2843), .B(n2615), .Z(o[526]) );
  AND U2697 ( .A(n2844), .B(n2845), .Z(n2843) );
  XNOR U2698 ( .A(n2846), .B(n2623), .Z(o[525]) );
  AND U2699 ( .A(n2847), .B(n2848), .Z(n2846) );
  XNOR U2700 ( .A(n2849), .B(n2627), .Z(o[524]) );
  AND U2701 ( .A(n2850), .B(n2851), .Z(n2849) );
  XNOR U2702 ( .A(n2852), .B(n2631), .Z(o[523]) );
  AND U2703 ( .A(n2853), .B(n2854), .Z(n2852) );
  XNOR U2704 ( .A(n2855), .B(n2635), .Z(o[522]) );
  AND U2705 ( .A(n2856), .B(n2857), .Z(n2855) );
  XNOR U2706 ( .A(n2858), .B(n2639), .Z(o[521]) );
  AND U2707 ( .A(n2859), .B(n2860), .Z(n2858) );
  XNOR U2708 ( .A(n2861), .B(n2643), .Z(o[520]) );
  XNOR U2709 ( .A(n2863), .B(n2864), .Z(o[51]) );
  AND U2710 ( .A(n2865), .B(n2866), .Z(n2863) );
  XNOR U2711 ( .A(n2867), .B(n2647), .Z(o[519]) );
  AND U2712 ( .A(n2868), .B(n2869), .Z(n2867) );
  XNOR U2713 ( .A(n2870), .B(n2651), .Z(o[518]) );
  AND U2714 ( .A(n2871), .B(n2872), .Z(n2870) );
  XNOR U2715 ( .A(n2873), .B(n2655), .Z(o[517]) );
  AND U2716 ( .A(n2874), .B(n2875), .Z(n2873) );
  XNOR U2717 ( .A(n2876), .B(n2659), .Z(o[516]) );
  AND U2718 ( .A(n2877), .B(n2878), .Z(n2876) );
  XNOR U2719 ( .A(n2879), .B(n2667), .Z(o[515]) );
  AND U2720 ( .A(n2880), .B(n2881), .Z(n2879) );
  XNOR U2721 ( .A(n2882), .B(n2671), .Z(o[514]) );
  AND U2722 ( .A(n2883), .B(n2884), .Z(n2882) );
  XNOR U2723 ( .A(n2885), .B(n2675), .Z(o[513]) );
  AND U2724 ( .A(n2886), .B(n2887), .Z(n2885) );
  XNOR U2725 ( .A(n2888), .B(n2679), .Z(o[512]) );
  AND U2726 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U2727 ( .A(n2891), .B(n2401), .Z(o[511]) );
  IV U2728 ( .A(n2683), .Z(n2401) );
  XNOR U2729 ( .A(n2157), .B(round_reg[885]), .Z(n2683) );
  ANDN U2730 ( .A(n2892), .B(n2682), .Z(n2891) );
  XOR U2731 ( .A(n2893), .B(n2405), .Z(o[510]) );
  IV U2732 ( .A(n2686), .Z(n2405) );
  XNOR U2733 ( .A(n2161), .B(round_reg[884]), .Z(n2686) );
  ANDN U2734 ( .A(n2894), .B(n2685), .Z(n2893) );
  XNOR U2735 ( .A(n2895), .B(n2896), .Z(o[50]) );
  AND U2736 ( .A(n2897), .B(n2898), .Z(n2895) );
  XOR U2737 ( .A(n2899), .B(n2409), .Z(o[509]) );
  IV U2738 ( .A(n2689), .Z(n2409) );
  XNOR U2739 ( .A(n2165), .B(round_reg[883]), .Z(n2689) );
  ANDN U2740 ( .A(n2900), .B(n2688), .Z(n2899) );
  XOR U2741 ( .A(n2901), .B(n2413), .Z(o[508]) );
  IV U2742 ( .A(n2692), .Z(n2413) );
  XNOR U2743 ( .A(n2169), .B(round_reg[882]), .Z(n2692) );
  ANDN U2744 ( .A(n2902), .B(n2691), .Z(n2901) );
  XOR U2745 ( .A(n2903), .B(n2417), .Z(o[507]) );
  IV U2746 ( .A(n2695), .Z(n2417) );
  XNOR U2747 ( .A(n2173), .B(round_reg[881]), .Z(n2695) );
  XOR U2748 ( .A(n2905), .B(n2421), .Z(o[506]) );
  IV U2749 ( .A(n2698), .Z(n2421) );
  XNOR U2750 ( .A(n2181), .B(round_reg[880]), .Z(n2698) );
  XOR U2751 ( .A(n2907), .B(n2425), .Z(o[505]) );
  IV U2752 ( .A(n2705), .Z(n2425) );
  XNOR U2753 ( .A(n2185), .B(round_reg[879]), .Z(n2705) );
  ANDN U2754 ( .A(n2908), .B(n2704), .Z(n2907) );
  XOR U2755 ( .A(n2909), .B(n2429), .Z(o[504]) );
  IV U2756 ( .A(n2708), .Z(n2429) );
  XNOR U2757 ( .A(n2189), .B(round_reg[878]), .Z(n2708) );
  ANDN U2758 ( .A(n2910), .B(n2707), .Z(n2909) );
  XOR U2759 ( .A(n2911), .B(n2433), .Z(o[503]) );
  IV U2760 ( .A(n2711), .Z(n2433) );
  XNOR U2761 ( .A(n2193), .B(round_reg[877]), .Z(n2711) );
  ANDN U2762 ( .A(n2912), .B(n2710), .Z(n2911) );
  XOR U2763 ( .A(n2913), .B(n2437), .Z(o[502]) );
  IV U2764 ( .A(n2714), .Z(n2437) );
  XNOR U2765 ( .A(n2197), .B(round_reg[876]), .Z(n2714) );
  ANDN U2766 ( .A(n2914), .B(n2713), .Z(n2913) );
  XOR U2767 ( .A(n2915), .B(n2445), .Z(o[501]) );
  IV U2768 ( .A(n2717), .Z(n2445) );
  XNOR U2769 ( .A(n2201), .B(round_reg[875]), .Z(n2717) );
  ANDN U2770 ( .A(n2916), .B(n2716), .Z(n2915) );
  XOR U2771 ( .A(n2917), .B(n2449), .Z(o[500]) );
  IV U2772 ( .A(n2720), .Z(n2449) );
  XNOR U2773 ( .A(n2205), .B(round_reg[874]), .Z(n2720) );
  ANDN U2774 ( .A(n2918), .B(n2719), .Z(n2917) );
  XNOR U2775 ( .A(n2919), .B(n2176), .Z(o[4]) );
  AND U2776 ( .A(n2920), .B(n2921), .Z(n2919) );
  XNOR U2777 ( .A(n2922), .B(n2923), .Z(o[49]) );
  AND U2778 ( .A(n2924), .B(n2925), .Z(n2922) );
  XOR U2779 ( .A(n2926), .B(n2453), .Z(o[499]) );
  IV U2780 ( .A(n2723), .Z(n2453) );
  XNOR U2781 ( .A(n2209), .B(round_reg[873]), .Z(n2723) );
  ANDN U2782 ( .A(n2927), .B(n2722), .Z(n2926) );
  XOR U2783 ( .A(n2928), .B(n2457), .Z(o[498]) );
  IV U2784 ( .A(n2726), .Z(n2457) );
  XNOR U2785 ( .A(n2213), .B(round_reg[872]), .Z(n2726) );
  ANDN U2786 ( .A(n2929), .B(n2725), .Z(n2928) );
  XOR U2787 ( .A(n2930), .B(n2461), .Z(o[497]) );
  IV U2788 ( .A(n2729), .Z(n2461) );
  XNOR U2789 ( .A(n2217), .B(round_reg[871]), .Z(n2729) );
  ANDN U2790 ( .A(n2931), .B(n2728), .Z(n2930) );
  XOR U2791 ( .A(n2932), .B(n2465), .Z(o[496]) );
  IV U2792 ( .A(n2732), .Z(n2465) );
  XNOR U2793 ( .A(n2225), .B(round_reg[870]), .Z(n2732) );
  ANDN U2794 ( .A(n2933), .B(n2731), .Z(n2932) );
  XOR U2795 ( .A(n2934), .B(n2469), .Z(o[495]) );
  IV U2796 ( .A(n2739), .Z(n2469) );
  XNOR U2797 ( .A(n2229), .B(round_reg[869]), .Z(n2739) );
  ANDN U2798 ( .A(n2935), .B(n2738), .Z(n2934) );
  XOR U2799 ( .A(n2936), .B(n2473), .Z(o[494]) );
  IV U2800 ( .A(n2742), .Z(n2473) );
  XNOR U2801 ( .A(n2233), .B(round_reg[868]), .Z(n2742) );
  ANDN U2802 ( .A(n2937), .B(n2741), .Z(n2936) );
  XOR U2803 ( .A(n2938), .B(n2477), .Z(o[493]) );
  IV U2804 ( .A(n2745), .Z(n2477) );
  XNOR U2805 ( .A(n2237), .B(round_reg[867]), .Z(n2745) );
  ANDN U2806 ( .A(n2939), .B(n2744), .Z(n2938) );
  XOR U2807 ( .A(n2940), .B(n2481), .Z(o[492]) );
  IV U2808 ( .A(n2748), .Z(n2481) );
  XNOR U2809 ( .A(n2241), .B(round_reg[866]), .Z(n2748) );
  ANDN U2810 ( .A(n2941), .B(n2747), .Z(n2940) );
  XOR U2811 ( .A(n2942), .B(n2489), .Z(o[491]) );
  IV U2812 ( .A(n2751), .Z(n2489) );
  XNOR U2813 ( .A(n2245), .B(round_reg[865]), .Z(n2751) );
  ANDN U2814 ( .A(n2943), .B(n2750), .Z(n2942) );
  XOR U2815 ( .A(n2944), .B(n2493), .Z(o[490]) );
  XNOR U2816 ( .A(n2249), .B(round_reg[864]), .Z(n2493) );
  ANDN U2817 ( .A(n2945), .B(n2753), .Z(n2944) );
  XNOR U2818 ( .A(n2946), .B(n2947), .Z(o[48]) );
  AND U2819 ( .A(n2948), .B(n2949), .Z(n2946) );
  XOR U2820 ( .A(n2950), .B(n2497), .Z(o[489]) );
  XNOR U2821 ( .A(n2253), .B(round_reg[863]), .Z(n2497) );
  ANDN U2822 ( .A(n2951), .B(n2755), .Z(n2950) );
  XOR U2823 ( .A(n2952), .B(n2501), .Z(o[488]) );
  XNOR U2824 ( .A(n2257), .B(round_reg[862]), .Z(n2501) );
  ANDN U2825 ( .A(n2953), .B(n2757), .Z(n2952) );
  XOR U2826 ( .A(n2954), .B(n2505), .Z(o[487]) );
  XNOR U2827 ( .A(n2261), .B(round_reg[861]), .Z(n2505) );
  ANDN U2828 ( .A(n2955), .B(n2759), .Z(n2954) );
  XOR U2829 ( .A(n2956), .B(n2509), .Z(o[486]) );
  XNOR U2830 ( .A(n2269), .B(round_reg[860]), .Z(n2509) );
  ANDN U2831 ( .A(n2957), .B(n2761), .Z(n2956) );
  XOR U2832 ( .A(n2958), .B(n2513), .Z(o[485]) );
  IV U2833 ( .A(n2768), .Z(n2513) );
  XNOR U2834 ( .A(n2273), .B(round_reg[859]), .Z(n2768) );
  ANDN U2835 ( .A(n2959), .B(n2767), .Z(n2958) );
  XOR U2836 ( .A(n2960), .B(n2517), .Z(o[484]) );
  IV U2837 ( .A(n2771), .Z(n2517) );
  XNOR U2838 ( .A(n2277), .B(round_reg[858]), .Z(n2771) );
  ANDN U2839 ( .A(n2961), .B(n2770), .Z(n2960) );
  XOR U2840 ( .A(n2962), .B(n2521), .Z(o[483]) );
  IV U2841 ( .A(n2774), .Z(n2521) );
  XNOR U2842 ( .A(n2281), .B(round_reg[857]), .Z(n2774) );
  NOR U2843 ( .A(n2963), .B(n2773), .Z(n2962) );
  XOR U2844 ( .A(n2964), .B(n2525), .Z(o[482]) );
  IV U2845 ( .A(n2777), .Z(n2525) );
  XNOR U2846 ( .A(n2285), .B(round_reg[856]), .Z(n2777) );
  NOR U2847 ( .A(n2965), .B(n2776), .Z(n2964) );
  XOR U2848 ( .A(n2966), .B(n2533), .Z(o[481]) );
  IV U2849 ( .A(n2780), .Z(n2533) );
  XNOR U2850 ( .A(n2289), .B(round_reg[855]), .Z(n2780) );
  NOR U2851 ( .A(n2967), .B(n2779), .Z(n2966) );
  XOR U2852 ( .A(n2968), .B(n2537), .Z(o[480]) );
  IV U2853 ( .A(n2783), .Z(n2537) );
  XNOR U2854 ( .A(n2293), .B(round_reg[854]), .Z(n2783) );
  NOR U2855 ( .A(n2969), .B(n2782), .Z(n2968) );
  XNOR U2856 ( .A(n2970), .B(n2971), .Z(o[47]) );
  AND U2857 ( .A(n2972), .B(n2973), .Z(n2970) );
  XOR U2858 ( .A(n2974), .B(n2541), .Z(o[479]) );
  IV U2859 ( .A(n2786), .Z(n2541) );
  XNOR U2860 ( .A(n2297), .B(round_reg[853]), .Z(n2786) );
  ANDN U2861 ( .A(n2975), .B(n2785), .Z(n2974) );
  XOR U2862 ( .A(n2976), .B(n2545), .Z(o[478]) );
  IV U2863 ( .A(n2789), .Z(n2545) );
  XNOR U2864 ( .A(n2301), .B(round_reg[852]), .Z(n2789) );
  NOR U2865 ( .A(n2977), .B(n2788), .Z(n2976) );
  XOR U2866 ( .A(n2978), .B(n2549), .Z(o[477]) );
  IV U2867 ( .A(n2792), .Z(n2549) );
  XNOR U2868 ( .A(n2305), .B(round_reg[851]), .Z(n2792) );
  NOR U2869 ( .A(n2979), .B(n2791), .Z(n2978) );
  XOR U2870 ( .A(n2980), .B(n2553), .Z(o[476]) );
  IV U2871 ( .A(n2795), .Z(n2553) );
  XNOR U2872 ( .A(n2313), .B(round_reg[850]), .Z(n2795) );
  NOR U2873 ( .A(n2981), .B(n2794), .Z(n2980) );
  XOR U2874 ( .A(n2982), .B(n2557), .Z(o[475]) );
  IV U2875 ( .A(n2802), .Z(n2557) );
  XNOR U2876 ( .A(n2317), .B(round_reg[849]), .Z(n2802) );
  NOR U2877 ( .A(n2983), .B(n2801), .Z(n2982) );
  XOR U2878 ( .A(n2984), .B(n2561), .Z(o[474]) );
  IV U2879 ( .A(n2805), .Z(n2561) );
  XNOR U2880 ( .A(n2321), .B(round_reg[848]), .Z(n2805) );
  ANDN U2881 ( .A(n2985), .B(n2804), .Z(n2984) );
  XOR U2882 ( .A(n2986), .B(n2565), .Z(o[473]) );
  IV U2883 ( .A(n2808), .Z(n2565) );
  XNOR U2884 ( .A(n2325), .B(round_reg[847]), .Z(n2808) );
  NOR U2885 ( .A(n2987), .B(n2807), .Z(n2986) );
  XOR U2886 ( .A(n2988), .B(n2569), .Z(o[472]) );
  IV U2887 ( .A(n2811), .Z(n2569) );
  XNOR U2888 ( .A(n2329), .B(round_reg[846]), .Z(n2811) );
  ANDN U2889 ( .A(n2989), .B(n2810), .Z(n2988) );
  XOR U2890 ( .A(n2990), .B(n2580), .Z(o[471]) );
  IV U2891 ( .A(n2814), .Z(n2580) );
  XNOR U2892 ( .A(n2333), .B(round_reg[845]), .Z(n2814) );
  ANDN U2893 ( .A(n2991), .B(n2813), .Z(n2990) );
  XOR U2894 ( .A(n2992), .B(n2584), .Z(o[470]) );
  IV U2895 ( .A(n2817), .Z(n2584) );
  XNOR U2896 ( .A(n2337), .B(round_reg[844]), .Z(n2817) );
  ANDN U2897 ( .A(n2993), .B(n2816), .Z(n2992) );
  XNOR U2898 ( .A(n2994), .B(n2995), .Z(o[46]) );
  AND U2899 ( .A(n2996), .B(n2997), .Z(n2994) );
  XOR U2900 ( .A(n2998), .B(n2588), .Z(o[469]) );
  IV U2901 ( .A(n2820), .Z(n2588) );
  XNOR U2902 ( .A(n2341), .B(round_reg[843]), .Z(n2820) );
  ANDN U2903 ( .A(n2999), .B(n2819), .Z(n2998) );
  XOR U2904 ( .A(n3000), .B(n2592), .Z(o[468]) );
  IV U2905 ( .A(n2823), .Z(n2592) );
  XNOR U2906 ( .A(n2345), .B(round_reg[842]), .Z(n2823) );
  ANDN U2907 ( .A(n3001), .B(n2822), .Z(n3000) );
  XOR U2908 ( .A(n3002), .B(n2596), .Z(o[467]) );
  IV U2909 ( .A(n2826), .Z(n2596) );
  XNOR U2910 ( .A(n2349), .B(round_reg[841]), .Z(n2826) );
  ANDN U2911 ( .A(n3003), .B(n2825), .Z(n3002) );
  XOR U2912 ( .A(n3004), .B(n2600), .Z(o[466]) );
  IV U2913 ( .A(n2829), .Z(n2600) );
  XNOR U2914 ( .A(n2357), .B(round_reg[840]), .Z(n2829) );
  ANDN U2915 ( .A(n3005), .B(n2828), .Z(n3004) );
  XOR U2916 ( .A(n3006), .B(n2604), .Z(o[465]) );
  IV U2917 ( .A(n2836), .Z(n2604) );
  XNOR U2918 ( .A(n2361), .B(round_reg[839]), .Z(n2836) );
  NOR U2919 ( .A(n3007), .B(n2835), .Z(n3006) );
  XOR U2920 ( .A(n3008), .B(n2608), .Z(o[464]) );
  IV U2921 ( .A(n2839), .Z(n2608) );
  XNOR U2922 ( .A(n2365), .B(round_reg[838]), .Z(n2839) );
  NOR U2923 ( .A(n3009), .B(n2838), .Z(n3008) );
  XOR U2924 ( .A(n3010), .B(n2612), .Z(o[463]) );
  IV U2925 ( .A(n2842), .Z(n2612) );
  XNOR U2926 ( .A(n2369), .B(round_reg[837]), .Z(n2842) );
  NOR U2927 ( .A(n3011), .B(n2841), .Z(n3010) );
  XOR U2928 ( .A(n3012), .B(n2616), .Z(o[462]) );
  IV U2929 ( .A(n2845), .Z(n2616) );
  XNOR U2930 ( .A(n2373), .B(round_reg[836]), .Z(n2845) );
  NOR U2931 ( .A(n3013), .B(n2844), .Z(n3012) );
  XOR U2932 ( .A(n3014), .B(n2624), .Z(o[461]) );
  IV U2933 ( .A(n2848), .Z(n2624) );
  XNOR U2934 ( .A(n2377), .B(round_reg[835]), .Z(n2848) );
  NOR U2935 ( .A(n3015), .B(n2847), .Z(n3014) );
  XOR U2936 ( .A(n3016), .B(n2628), .Z(o[460]) );
  IV U2937 ( .A(n2851), .Z(n2628) );
  XNOR U2938 ( .A(n2381), .B(round_reg[834]), .Z(n2851) );
  NOR U2939 ( .A(n3017), .B(n2850), .Z(n3016) );
  XNOR U2940 ( .A(n3018), .B(n3019), .Z(o[45]) );
  AND U2941 ( .A(n3020), .B(n3021), .Z(n3018) );
  XOR U2942 ( .A(n3022), .B(n2632), .Z(o[459]) );
  IV U2943 ( .A(n2854), .Z(n2632) );
  XNOR U2944 ( .A(n2385), .B(round_reg[833]), .Z(n2854) );
  NOR U2945 ( .A(n3023), .B(n2853), .Z(n3022) );
  XOR U2946 ( .A(n3024), .B(n2636), .Z(o[458]) );
  IV U2947 ( .A(n2857), .Z(n2636) );
  XNOR U2948 ( .A(n2389), .B(round_reg[832]), .Z(n2857) );
  ANDN U2949 ( .A(n3025), .B(n2856), .Z(n3024) );
  XOR U2950 ( .A(n3026), .B(n2640), .Z(o[457]) );
  IV U2951 ( .A(n2860), .Z(n2640) );
  XNOR U2952 ( .A(n2393), .B(round_reg[895]), .Z(n2860) );
  NOR U2953 ( .A(n3027), .B(n2859), .Z(n3026) );
  XOR U2954 ( .A(n3028), .B(n2644), .Z(o[456]) );
  XOR U2955 ( .A(n3029), .B(round_reg[894]), .Z(n2644) );
  XOR U2956 ( .A(n3031), .B(n2648), .Z(o[455]) );
  IV U2957 ( .A(n2869), .Z(n2648) );
  XNOR U2958 ( .A(n2117), .B(round_reg[893]), .Z(n2869) );
  XOR U2959 ( .A(n3033), .B(n2652), .Z(o[454]) );
  IV U2960 ( .A(n2872), .Z(n2652) );
  XNOR U2961 ( .A(n2121), .B(round_reg[892]), .Z(n2872) );
  XOR U2962 ( .A(n3035), .B(n2656), .Z(o[453]) );
  IV U2963 ( .A(n2875), .Z(n2656) );
  XNOR U2964 ( .A(n2125), .B(round_reg[891]), .Z(n2875) );
  XOR U2965 ( .A(n3037), .B(n2660), .Z(o[452]) );
  IV U2966 ( .A(n2878), .Z(n2660) );
  XNOR U2967 ( .A(n2136), .B(round_reg[890]), .Z(n2878) );
  XOR U2968 ( .A(n3039), .B(n2668), .Z(o[451]) );
  IV U2969 ( .A(n2881), .Z(n2668) );
  XNOR U2970 ( .A(n2141), .B(round_reg[889]), .Z(n2881) );
  ANDN U2971 ( .A(n3040), .B(n2880), .Z(n3039) );
  XOR U2972 ( .A(n3041), .B(n2672), .Z(o[450]) );
  IV U2973 ( .A(n2884), .Z(n2672) );
  XNOR U2974 ( .A(n2145), .B(round_reg[888]), .Z(n2884) );
  ANDN U2975 ( .A(n3042), .B(n2883), .Z(n3041) );
  XNOR U2976 ( .A(n3043), .B(n3044), .Z(o[44]) );
  AND U2977 ( .A(n3045), .B(n3046), .Z(n3043) );
  XOR U2978 ( .A(n3047), .B(n2676), .Z(o[449]) );
  IV U2979 ( .A(n2887), .Z(n2676) );
  XNOR U2980 ( .A(n2149), .B(round_reg[887]), .Z(n2887) );
  ANDN U2981 ( .A(n3048), .B(n2886), .Z(n3047) );
  XOR U2982 ( .A(n3049), .B(n2680), .Z(o[448]) );
  IV U2983 ( .A(n2890), .Z(n2680) );
  XNOR U2984 ( .A(n2153), .B(round_reg[886]), .Z(n2890) );
  ANDN U2985 ( .A(n3050), .B(n2889), .Z(n3049) );
  XOR U2986 ( .A(n3051), .B(n2682), .Z(o[447]) );
  XOR U2987 ( .A(n2156), .B(round_reg[496]), .Z(n2682) );
  NOR U2988 ( .A(n2892), .B(n2399), .Z(n3051) );
  XOR U2989 ( .A(n3052), .B(n2685), .Z(o[446]) );
  XOR U2990 ( .A(n2160), .B(round_reg[495]), .Z(n2685) );
  NOR U2991 ( .A(n2894), .B(n2403), .Z(n3052) );
  XOR U2992 ( .A(n3053), .B(n2688), .Z(o[445]) );
  XOR U2993 ( .A(n2164), .B(round_reg[494]), .Z(n2688) );
  NOR U2994 ( .A(n2900), .B(n2407), .Z(n3053) );
  XOR U2995 ( .A(n3054), .B(n2691), .Z(o[444]) );
  XOR U2996 ( .A(n2168), .B(round_reg[493]), .Z(n2691) );
  NOR U2997 ( .A(n2902), .B(n2411), .Z(n3054) );
  XOR U2998 ( .A(n3055), .B(n2694), .Z(o[443]) );
  XNOR U2999 ( .A(n2172), .B(round_reg[492]), .Z(n2694) );
  NOR U3000 ( .A(n2904), .B(n2415), .Z(n3055) );
  XOR U3001 ( .A(n3056), .B(n2697), .Z(o[442]) );
  XNOR U3002 ( .A(n2180), .B(round_reg[491]), .Z(n2697) );
  NOR U3003 ( .A(n2906), .B(n2419), .Z(n3056) );
  XOR U3004 ( .A(n3057), .B(n2704), .Z(o[441]) );
  XOR U3005 ( .A(n2184), .B(round_reg[490]), .Z(n2704) );
  NOR U3006 ( .A(n2908), .B(n2423), .Z(n3057) );
  XOR U3007 ( .A(n3058), .B(n2707), .Z(o[440]) );
  XOR U3008 ( .A(n2188), .B(round_reg[489]), .Z(n2707) );
  NOR U3009 ( .A(n2910), .B(n2427), .Z(n3058) );
  XNOR U3010 ( .A(n3059), .B(n3060), .Z(o[43]) );
  AND U3011 ( .A(n3061), .B(n3062), .Z(n3059) );
  XOR U3012 ( .A(n3063), .B(n2710), .Z(o[439]) );
  XOR U3013 ( .A(n2192), .B(round_reg[488]), .Z(n2710) );
  NOR U3014 ( .A(n2912), .B(n2431), .Z(n3063) );
  XOR U3015 ( .A(n3064), .B(n2713), .Z(o[438]) );
  XOR U3016 ( .A(n2196), .B(round_reg[487]), .Z(n2713) );
  NOR U3017 ( .A(n2914), .B(n2435), .Z(n3064) );
  XOR U3018 ( .A(n3065), .B(n2716), .Z(o[437]) );
  XOR U3019 ( .A(n2200), .B(round_reg[486]), .Z(n2716) );
  NOR U3020 ( .A(n2916), .B(n2443), .Z(n3065) );
  XOR U3021 ( .A(n3066), .B(n2719), .Z(o[436]) );
  XOR U3022 ( .A(n2204), .B(round_reg[485]), .Z(n2719) );
  NOR U3023 ( .A(n2447), .B(n2918), .Z(n3066) );
  XOR U3024 ( .A(n3067), .B(n2722), .Z(o[435]) );
  XOR U3025 ( .A(n2208), .B(round_reg[484]), .Z(n2722) );
  ANDN U3026 ( .A(n3068), .B(n2451), .Z(n3067) );
  XOR U3027 ( .A(n3069), .B(n2725), .Z(o[434]) );
  XNOR U3028 ( .A(n2212), .B(round_reg[483]), .Z(n2725) );
  ANDN U3029 ( .A(n3070), .B(n2455), .Z(n3069) );
  XOR U3030 ( .A(n3071), .B(n2728), .Z(o[433]) );
  XOR U3031 ( .A(n2216), .B(round_reg[482]), .Z(n2728) );
  ANDN U3032 ( .A(n3072), .B(n2459), .Z(n3071) );
  XOR U3033 ( .A(n3073), .B(n2731), .Z(o[432]) );
  XOR U3034 ( .A(n2224), .B(round_reg[481]), .Z(n2731) );
  ANDN U3035 ( .A(n3074), .B(n2463), .Z(n3073) );
  XOR U3036 ( .A(n3075), .B(n2738), .Z(o[431]) );
  XOR U3037 ( .A(n2228), .B(round_reg[480]), .Z(n2738) );
  ANDN U3038 ( .A(n3076), .B(n2467), .Z(n3075) );
  XOR U3039 ( .A(n3077), .B(n2741), .Z(o[430]) );
  XOR U3040 ( .A(n2232), .B(round_reg[479]), .Z(n2741) );
  ANDN U3041 ( .A(n3078), .B(n2471), .Z(n3077) );
  XNOR U3042 ( .A(n3079), .B(n3080), .Z(o[42]) );
  AND U3043 ( .A(n3081), .B(n3082), .Z(n3079) );
  XOR U3044 ( .A(n3083), .B(n2744), .Z(o[429]) );
  XOR U3045 ( .A(n2236), .B(round_reg[478]), .Z(n2744) );
  ANDN U3046 ( .A(n3084), .B(n2475), .Z(n3083) );
  XOR U3047 ( .A(n3085), .B(n2747), .Z(o[428]) );
  XOR U3048 ( .A(n2240), .B(round_reg[477]), .Z(n2747) );
  ANDN U3049 ( .A(n3086), .B(n2479), .Z(n3085) );
  XOR U3050 ( .A(n3087), .B(n2750), .Z(o[427]) );
  XOR U3051 ( .A(n2244), .B(round_reg[476]), .Z(n2750) );
  ANDN U3052 ( .A(n3088), .B(n2487), .Z(n3087) );
  XOR U3053 ( .A(n3089), .B(n2753), .Z(o[426]) );
  XOR U3054 ( .A(n2248), .B(round_reg[475]), .Z(n2753) );
  ANDN U3055 ( .A(n3090), .B(n2491), .Z(n3089) );
  XOR U3056 ( .A(n3091), .B(n2755), .Z(o[425]) );
  XOR U3057 ( .A(n2252), .B(round_reg[474]), .Z(n2755) );
  ANDN U3058 ( .A(n3092), .B(n2495), .Z(n3091) );
  XOR U3059 ( .A(n3093), .B(n2757), .Z(o[424]) );
  XOR U3060 ( .A(n2256), .B(round_reg[473]), .Z(n2757) );
  ANDN U3061 ( .A(n3094), .B(n2499), .Z(n3093) );
  XOR U3062 ( .A(n3095), .B(n2759), .Z(o[423]) );
  XOR U3063 ( .A(n2260), .B(round_reg[472]), .Z(n2759) );
  ANDN U3064 ( .A(n3096), .B(n2503), .Z(n3095) );
  XOR U3065 ( .A(n3097), .B(n2761), .Z(o[422]) );
  XOR U3066 ( .A(n2268), .B(round_reg[471]), .Z(n2761) );
  ANDN U3067 ( .A(n3098), .B(n2507), .Z(n3097) );
  XOR U3068 ( .A(n3099), .B(n2767), .Z(o[421]) );
  XOR U3069 ( .A(n2272), .B(round_reg[470]), .Z(n2767) );
  ANDN U3070 ( .A(n3100), .B(n2511), .Z(n3099) );
  XOR U3071 ( .A(n3101), .B(n2770), .Z(o[420]) );
  XOR U3072 ( .A(n2276), .B(round_reg[469]), .Z(n2770) );
  XNOR U3073 ( .A(n3102), .B(n3103), .Z(o[41]) );
  AND U3074 ( .A(n3104), .B(n3105), .Z(n3102) );
  XOR U3075 ( .A(n3106), .B(n2773), .Z(o[419]) );
  XOR U3076 ( .A(n2280), .B(round_reg[468]), .Z(n2773) );
  ANDN U3077 ( .A(n2963), .B(n2519), .Z(n3106) );
  IV U3078 ( .A(n3107), .Z(n2963) );
  XOR U3079 ( .A(n3108), .B(n2776), .Z(o[418]) );
  XOR U3080 ( .A(n2284), .B(round_reg[467]), .Z(n2776) );
  ANDN U3081 ( .A(n2965), .B(n2523), .Z(n3108) );
  IV U3082 ( .A(n3109), .Z(n2965) );
  XOR U3083 ( .A(n3110), .B(n2779), .Z(o[417]) );
  XOR U3084 ( .A(n2288), .B(round_reg[466]), .Z(n2779) );
  ANDN U3085 ( .A(n2967), .B(n2531), .Z(n3110) );
  IV U3086 ( .A(n3111), .Z(n2967) );
  XOR U3087 ( .A(n3112), .B(n2782), .Z(o[416]) );
  XOR U3088 ( .A(n2292), .B(round_reg[465]), .Z(n2782) );
  ANDN U3089 ( .A(n2969), .B(n2535), .Z(n3112) );
  IV U3090 ( .A(n3113), .Z(n2969) );
  XOR U3091 ( .A(n3114), .B(n2785), .Z(o[415]) );
  XOR U3092 ( .A(n2296), .B(round_reg[464]), .Z(n2785) );
  XOR U3093 ( .A(n3115), .B(n2788), .Z(o[414]) );
  XOR U3094 ( .A(n2300), .B(round_reg[463]), .Z(n2788) );
  ANDN U3095 ( .A(n2977), .B(n2543), .Z(n3115) );
  IV U3096 ( .A(n3116), .Z(n2977) );
  XOR U3097 ( .A(n3117), .B(n2791), .Z(o[413]) );
  XOR U3098 ( .A(n2304), .B(round_reg[462]), .Z(n2791) );
  ANDN U3099 ( .A(n2979), .B(n2547), .Z(n3117) );
  IV U3100 ( .A(n3118), .Z(n2979) );
  XOR U3101 ( .A(n3119), .B(n2794), .Z(o[412]) );
  XOR U3102 ( .A(n2312), .B(round_reg[461]), .Z(n2794) );
  ANDN U3103 ( .A(n2981), .B(n2551), .Z(n3119) );
  IV U3104 ( .A(n3120), .Z(n2981) );
  XOR U3105 ( .A(n3121), .B(n2801), .Z(o[411]) );
  XOR U3106 ( .A(n2316), .B(round_reg[460]), .Z(n2801) );
  ANDN U3107 ( .A(n2983), .B(n2555), .Z(n3121) );
  IV U3108 ( .A(n3122), .Z(n2983) );
  XOR U3109 ( .A(n3123), .B(n2804), .Z(o[410]) );
  XOR U3110 ( .A(n2320), .B(round_reg[459]), .Z(n2804) );
  XNOR U3111 ( .A(n3124), .B(n3125), .Z(o[40]) );
  XOR U3112 ( .A(n3128), .B(n2807), .Z(o[409]) );
  XOR U3113 ( .A(n2324), .B(round_reg[458]), .Z(n2807) );
  ANDN U3114 ( .A(n2987), .B(n2563), .Z(n3128) );
  IV U3115 ( .A(n3129), .Z(n2987) );
  XOR U3116 ( .A(n3130), .B(n2810), .Z(o[408]) );
  XOR U3117 ( .A(n2328), .B(round_reg[457]), .Z(n2810) );
  ANDN U3118 ( .A(n3131), .B(n2567), .Z(n3130) );
  XOR U3119 ( .A(n3132), .B(n2813), .Z(o[407]) );
  XOR U3120 ( .A(n2332), .B(round_reg[456]), .Z(n2813) );
  ANDN U3121 ( .A(n3133), .B(n2578), .Z(n3132) );
  XOR U3122 ( .A(n3134), .B(n2816), .Z(o[406]) );
  XOR U3123 ( .A(n2336), .B(round_reg[455]), .Z(n2816) );
  ANDN U3124 ( .A(n3135), .B(n2582), .Z(n3134) );
  XOR U3125 ( .A(n3136), .B(n2819), .Z(o[405]) );
  XOR U3126 ( .A(n2340), .B(round_reg[454]), .Z(n2819) );
  ANDN U3127 ( .A(n3137), .B(n2586), .Z(n3136) );
  XOR U3128 ( .A(n3138), .B(n2822), .Z(o[404]) );
  XOR U3129 ( .A(n2344), .B(round_reg[453]), .Z(n2822) );
  ANDN U3130 ( .A(n3139), .B(n2590), .Z(n3138) );
  XOR U3131 ( .A(n3140), .B(n2825), .Z(o[403]) );
  XOR U3132 ( .A(n2348), .B(round_reg[452]), .Z(n2825) );
  ANDN U3133 ( .A(n3141), .B(n2594), .Z(n3140) );
  XOR U3134 ( .A(n3142), .B(n2828), .Z(o[402]) );
  XOR U3135 ( .A(n2356), .B(round_reg[451]), .Z(n2828) );
  XOR U3136 ( .A(n3143), .B(n2835), .Z(o[401]) );
  XOR U3137 ( .A(n2360), .B(round_reg[450]), .Z(n2835) );
  ANDN U3138 ( .A(n3007), .B(n2602), .Z(n3143) );
  IV U3139 ( .A(n3144), .Z(n3007) );
  XOR U3140 ( .A(n3145), .B(n2838), .Z(o[400]) );
  XOR U3141 ( .A(n2364), .B(round_reg[449]), .Z(n2838) );
  ANDN U3142 ( .A(n3009), .B(n2606), .Z(n3145) );
  IV U3143 ( .A(n3146), .Z(n3009) );
  XNOR U3144 ( .A(n3147), .B(n2220), .Z(o[3]) );
  AND U3145 ( .A(n3148), .B(n3149), .Z(n3147) );
  XNOR U3146 ( .A(n3150), .B(n3151), .Z(o[39]) );
  XOR U3147 ( .A(n3154), .B(n2841), .Z(o[399]) );
  XOR U3148 ( .A(n2368), .B(round_reg[448]), .Z(n2841) );
  ANDN U3149 ( .A(n3011), .B(n2610), .Z(n3154) );
  IV U3150 ( .A(n3155), .Z(n3011) );
  XOR U3151 ( .A(n3156), .B(n2844), .Z(o[398]) );
  XOR U3152 ( .A(n2372), .B(round_reg[511]), .Z(n2844) );
  ANDN U3153 ( .A(n3013), .B(n2614), .Z(n3156) );
  IV U3154 ( .A(n3157), .Z(n3013) );
  XOR U3155 ( .A(n3158), .B(n2847), .Z(o[397]) );
  XOR U3156 ( .A(n2376), .B(round_reg[510]), .Z(n2847) );
  ANDN U3157 ( .A(n3015), .B(n2622), .Z(n3158) );
  IV U3158 ( .A(n3159), .Z(n3015) );
  XOR U3159 ( .A(n3160), .B(n2850), .Z(o[396]) );
  XOR U3160 ( .A(n2380), .B(round_reg[509]), .Z(n2850) );
  ANDN U3161 ( .A(n3017), .B(n2626), .Z(n3160) );
  IV U3162 ( .A(n3161), .Z(n3017) );
  XOR U3163 ( .A(n3162), .B(n2853), .Z(o[395]) );
  XOR U3164 ( .A(n2384), .B(round_reg[508]), .Z(n2853) );
  ANDN U3165 ( .A(n3023), .B(n2630), .Z(n3162) );
  IV U3166 ( .A(n3163), .Z(n3023) );
  XOR U3167 ( .A(n3164), .B(n2856), .Z(o[394]) );
  XOR U3168 ( .A(n2388), .B(round_reg[507]), .Z(n2856) );
  NOR U3169 ( .A(n3025), .B(n2634), .Z(n3164) );
  XOR U3170 ( .A(n3165), .B(n2859), .Z(o[393]) );
  XOR U3171 ( .A(n2392), .B(round_reg[506]), .Z(n2859) );
  ANDN U3172 ( .A(n3027), .B(n2638), .Z(n3165) );
  IV U3173 ( .A(n3166), .Z(n3027) );
  XOR U3174 ( .A(n3167), .B(n2862), .Z(o[392]) );
  XOR U3175 ( .A(n2114), .B(round_reg[505]), .Z(n2862) );
  XOR U3176 ( .A(n3168), .B(n2868), .Z(o[391]) );
  XOR U3177 ( .A(n2118), .B(round_reg[504]), .Z(n2868) );
  XOR U3178 ( .A(n3169), .B(n2871), .Z(o[390]) );
  XOR U3179 ( .A(n2122), .B(round_reg[503]), .Z(n2871) );
  XNOR U3180 ( .A(n3170), .B(n3171), .Z(o[38]) );
  XOR U3181 ( .A(n3174), .B(n2874), .Z(o[389]) );
  XOR U3182 ( .A(n2126), .B(round_reg[502]), .Z(n2874) );
  XOR U3183 ( .A(n3175), .B(n2877), .Z(o[388]) );
  XOR U3184 ( .A(n2137), .B(round_reg[501]), .Z(n2877) );
  XOR U3185 ( .A(n3176), .B(n2880), .Z(o[387]) );
  XOR U3186 ( .A(n2140), .B(round_reg[500]), .Z(n2880) );
  NOR U3187 ( .A(n3040), .B(n2666), .Z(n3176) );
  XOR U3188 ( .A(n3177), .B(n2883), .Z(o[386]) );
  XOR U3189 ( .A(n2144), .B(round_reg[499]), .Z(n2883) );
  NOR U3190 ( .A(n3042), .B(n2670), .Z(n3177) );
  XOR U3191 ( .A(n3178), .B(n2886), .Z(o[385]) );
  XOR U3192 ( .A(n2148), .B(round_reg[498]), .Z(n2886) );
  NOR U3193 ( .A(n3048), .B(n2674), .Z(n3178) );
  XOR U3194 ( .A(n3179), .B(n2889), .Z(o[384]) );
  XOR U3195 ( .A(n2152), .B(round_reg[497]), .Z(n2889) );
  NOR U3196 ( .A(n3050), .B(n2678), .Z(n3179) );
  XOR U3197 ( .A(n3180), .B(n2892), .Z(o[383]) );
  XOR U3198 ( .A(n1815), .B(round_reg[71]), .Z(n2892) );
  ANDN U3199 ( .A(n2399), .B(n2400), .Z(n3180) );
  XNOR U3200 ( .A(n2195), .B(round_reg[1243]), .Z(n2400) );
  XNOR U3201 ( .A(n1991), .B(round_reg[1316]), .Z(n2399) );
  XOR U3202 ( .A(n3181), .B(n2894), .Z(o[382]) );
  XOR U3203 ( .A(n1826), .B(round_reg[70]), .Z(n2894) );
  ANDN U3204 ( .A(n2403), .B(n2404), .Z(n3181) );
  XNOR U3205 ( .A(n2199), .B(round_reg[1242]), .Z(n2404) );
  XNOR U3206 ( .A(n1993), .B(round_reg[1315]), .Z(n2403) );
  XOR U3207 ( .A(n3182), .B(n2900), .Z(o[381]) );
  XOR U3208 ( .A(n1829), .B(round_reg[69]), .Z(n2900) );
  ANDN U3209 ( .A(n2407), .B(n2408), .Z(n3182) );
  XNOR U3210 ( .A(n2203), .B(round_reg[1241]), .Z(n2408) );
  XNOR U3211 ( .A(n1995), .B(round_reg[1314]), .Z(n2407) );
  XOR U3212 ( .A(n3183), .B(n2902), .Z(o[380]) );
  XOR U3213 ( .A(n1832), .B(round_reg[68]), .Z(n2902) );
  ANDN U3214 ( .A(n2411), .B(n2412), .Z(n3183) );
  XNOR U3215 ( .A(n2207), .B(round_reg[1240]), .Z(n2412) );
  XNOR U3216 ( .A(n1997), .B(round_reg[1313]), .Z(n2411) );
  XNOR U3217 ( .A(n3184), .B(n3185), .Z(o[37]) );
  XOR U3218 ( .A(n3188), .B(n2904), .Z(o[379]) );
  XOR U3219 ( .A(n1835), .B(round_reg[67]), .Z(n2904) );
  ANDN U3220 ( .A(n2415), .B(n2416), .Z(n3188) );
  XNOR U3221 ( .A(n2211), .B(round_reg[1239]), .Z(n2416) );
  XNOR U3222 ( .A(n1999), .B(round_reg[1312]), .Z(n2415) );
  XOR U3223 ( .A(n3189), .B(n2906), .Z(o[378]) );
  XOR U3224 ( .A(n1838), .B(round_reg[66]), .Z(n2906) );
  ANDN U3225 ( .A(n2419), .B(n2420), .Z(n3189) );
  XNOR U3226 ( .A(n2215), .B(round_reg[1238]), .Z(n2420) );
  XNOR U3227 ( .A(n2001), .B(round_reg[1311]), .Z(n2419) );
  XOR U3228 ( .A(n3190), .B(n2908), .Z(o[377]) );
  XOR U3229 ( .A(n1841), .B(round_reg[65]), .Z(n2908) );
  ANDN U3230 ( .A(n2423), .B(n2424), .Z(n3190) );
  XNOR U3231 ( .A(n2223), .B(round_reg[1237]), .Z(n2424) );
  XNOR U3232 ( .A(n2003), .B(round_reg[1310]), .Z(n2423) );
  XOR U3233 ( .A(n3191), .B(n2910), .Z(o[376]) );
  XOR U3234 ( .A(n1844), .B(round_reg[64]), .Z(n2910) );
  ANDN U3235 ( .A(n2427), .B(n2428), .Z(n3191) );
  XNOR U3236 ( .A(n2227), .B(round_reg[1236]), .Z(n2428) );
  XNOR U3237 ( .A(n2005), .B(round_reg[1309]), .Z(n2427) );
  XOR U3238 ( .A(n3192), .B(n2912), .Z(o[375]) );
  XOR U3239 ( .A(n1847), .B(round_reg[127]), .Z(n2912) );
  ANDN U3240 ( .A(n2431), .B(n2432), .Z(n3192) );
  XNOR U3241 ( .A(n2231), .B(round_reg[1235]), .Z(n2432) );
  XNOR U3242 ( .A(n2007), .B(round_reg[1308]), .Z(n2431) );
  XOR U3243 ( .A(n3193), .B(n2914), .Z(o[374]) );
  XOR U3244 ( .A(n1850), .B(round_reg[126]), .Z(n2914) );
  ANDN U3245 ( .A(n2435), .B(n2436), .Z(n3193) );
  XNOR U3246 ( .A(n2235), .B(round_reg[1234]), .Z(n2436) );
  XNOR U3247 ( .A(n2012), .B(round_reg[1307]), .Z(n2435) );
  XOR U3248 ( .A(n3194), .B(n2916), .Z(o[373]) );
  XOR U3249 ( .A(n1853), .B(round_reg[125]), .Z(n2916) );
  ANDN U3250 ( .A(n2443), .B(n2444), .Z(n3194) );
  XNOR U3251 ( .A(n2239), .B(round_reg[1233]), .Z(n2444) );
  XNOR U3252 ( .A(n2014), .B(round_reg[1306]), .Z(n2443) );
  XOR U3253 ( .A(n3195), .B(n2918), .Z(o[372]) );
  XOR U3254 ( .A(n1860), .B(round_reg[124]), .Z(n2918) );
  ANDN U3255 ( .A(n2447), .B(n2448), .Z(n3195) );
  XNOR U3256 ( .A(n2243), .B(round_reg[1232]), .Z(n2448) );
  XNOR U3257 ( .A(n2016), .B(round_reg[1305]), .Z(n2447) );
  XOR U3258 ( .A(n3196), .B(n2927), .Z(o[371]) );
  IV U3259 ( .A(n3068), .Z(n2927) );
  XNOR U3260 ( .A(n1863), .B(round_reg[123]), .Z(n3068) );
  ANDN U3261 ( .A(n2451), .B(n2452), .Z(n3196) );
  XNOR U3262 ( .A(n2247), .B(round_reg[1231]), .Z(n2452) );
  XNOR U3263 ( .A(n2018), .B(round_reg[1304]), .Z(n2451) );
  XOR U3264 ( .A(n3197), .B(n2929), .Z(o[370]) );
  IV U3265 ( .A(n3070), .Z(n2929) );
  XNOR U3266 ( .A(n1866), .B(round_reg[122]), .Z(n3070) );
  ANDN U3267 ( .A(n2455), .B(n2456), .Z(n3197) );
  XNOR U3268 ( .A(n2251), .B(round_reg[1230]), .Z(n2456) );
  XNOR U3269 ( .A(n2020), .B(round_reg[1303]), .Z(n2455) );
  XNOR U3270 ( .A(n3198), .B(n3199), .Z(o[36]) );
  XOR U3271 ( .A(n3202), .B(n2931), .Z(o[369]) );
  IV U3272 ( .A(n3072), .Z(n2931) );
  XNOR U3273 ( .A(n1869), .B(round_reg[121]), .Z(n3072) );
  ANDN U3274 ( .A(n2459), .B(n2460), .Z(n3202) );
  XNOR U3275 ( .A(n2255), .B(round_reg[1229]), .Z(n2460) );
  XNOR U3276 ( .A(n2022), .B(round_reg[1302]), .Z(n2459) );
  XOR U3277 ( .A(n3203), .B(n2933), .Z(o[368]) );
  IV U3278 ( .A(n3074), .Z(n2933) );
  XNOR U3279 ( .A(n1872), .B(round_reg[120]), .Z(n3074) );
  ANDN U3280 ( .A(n2463), .B(n2464), .Z(n3203) );
  XNOR U3281 ( .A(n2259), .B(round_reg[1228]), .Z(n2464) );
  XNOR U3282 ( .A(n2024), .B(round_reg[1301]), .Z(n2463) );
  XOR U3283 ( .A(n3204), .B(n2935), .Z(o[367]) );
  IV U3284 ( .A(n3076), .Z(n2935) );
  XNOR U3285 ( .A(n1875), .B(round_reg[119]), .Z(n3076) );
  ANDN U3286 ( .A(n2467), .B(n2468), .Z(n3204) );
  XNOR U3287 ( .A(n2267), .B(round_reg[1227]), .Z(n2468) );
  XNOR U3288 ( .A(n2026), .B(round_reg[1300]), .Z(n2467) );
  XOR U3289 ( .A(n3205), .B(n2937), .Z(o[366]) );
  IV U3290 ( .A(n3078), .Z(n2937) );
  XNOR U3291 ( .A(n1878), .B(round_reg[118]), .Z(n3078) );
  ANDN U3292 ( .A(n2471), .B(n2472), .Z(n3205) );
  XNOR U3293 ( .A(n2271), .B(round_reg[1226]), .Z(n2472) );
  XNOR U3294 ( .A(n2028), .B(round_reg[1299]), .Z(n2471) );
  XOR U3295 ( .A(n3206), .B(n2939), .Z(o[365]) );
  IV U3296 ( .A(n3084), .Z(n2939) );
  XNOR U3297 ( .A(n1881), .B(round_reg[117]), .Z(n3084) );
  ANDN U3298 ( .A(n2475), .B(n2476), .Z(n3206) );
  XNOR U3299 ( .A(n2275), .B(round_reg[1225]), .Z(n2476) );
  XNOR U3300 ( .A(n2031), .B(round_reg[1298]), .Z(n2475) );
  XOR U3301 ( .A(n3207), .B(n2941), .Z(o[364]) );
  IV U3302 ( .A(n3086), .Z(n2941) );
  XNOR U3303 ( .A(n1884), .B(round_reg[116]), .Z(n3086) );
  ANDN U3304 ( .A(n2479), .B(n2480), .Z(n3207) );
  XNOR U3305 ( .A(n2279), .B(round_reg[1224]), .Z(n2480) );
  XNOR U3306 ( .A(n2036), .B(round_reg[1297]), .Z(n2479) );
  XOR U3307 ( .A(n3208), .B(n2943), .Z(o[363]) );
  IV U3308 ( .A(n3088), .Z(n2943) );
  XNOR U3309 ( .A(n1887), .B(round_reg[115]), .Z(n3088) );
  ANDN U3310 ( .A(n2487), .B(n2488), .Z(n3208) );
  XNOR U3311 ( .A(n2283), .B(round_reg[1223]), .Z(n2488) );
  XNOR U3312 ( .A(n2039), .B(round_reg[1296]), .Z(n2487) );
  XOR U3313 ( .A(n3209), .B(n2945), .Z(o[362]) );
  IV U3314 ( .A(n3090), .Z(n2945) );
  XNOR U3315 ( .A(n1894), .B(round_reg[114]), .Z(n3090) );
  ANDN U3316 ( .A(n2491), .B(n2492), .Z(n3209) );
  XNOR U3317 ( .A(n2287), .B(round_reg[1222]), .Z(n2492) );
  XNOR U3318 ( .A(n2042), .B(round_reg[1295]), .Z(n2491) );
  XOR U3319 ( .A(n3210), .B(n2951), .Z(o[361]) );
  IV U3320 ( .A(n3092), .Z(n2951) );
  XNOR U3321 ( .A(n1897), .B(round_reg[113]), .Z(n3092) );
  ANDN U3322 ( .A(n2495), .B(n2496), .Z(n3210) );
  XNOR U3323 ( .A(n2291), .B(round_reg[1221]), .Z(n2496) );
  XNOR U3324 ( .A(n2044), .B(round_reg[1294]), .Z(n2495) );
  XOR U3325 ( .A(n3211), .B(n2953), .Z(o[360]) );
  IV U3326 ( .A(n3094), .Z(n2953) );
  XNOR U3327 ( .A(n1900), .B(round_reg[112]), .Z(n3094) );
  ANDN U3328 ( .A(n2499), .B(n2500), .Z(n3211) );
  XNOR U3329 ( .A(n2295), .B(round_reg[1220]), .Z(n2500) );
  XNOR U3330 ( .A(n2047), .B(round_reg[1293]), .Z(n2499) );
  XOR U3331 ( .A(n3212), .B(n1058), .Z(o[35]) );
  ANDN U3332 ( .A(n3213), .B(n1057), .Z(n3212) );
  XOR U3333 ( .A(n3214), .B(n2955), .Z(o[359]) );
  IV U3334 ( .A(n3096), .Z(n2955) );
  XNOR U3335 ( .A(n1903), .B(round_reg[111]), .Z(n3096) );
  ANDN U3336 ( .A(n2503), .B(n2504), .Z(n3214) );
  XNOR U3337 ( .A(n2299), .B(round_reg[1219]), .Z(n2504) );
  XNOR U3338 ( .A(n2050), .B(round_reg[1292]), .Z(n2503) );
  XOR U3339 ( .A(n3215), .B(n2957), .Z(o[358]) );
  IV U3340 ( .A(n3098), .Z(n2957) );
  XNOR U3341 ( .A(n1906), .B(round_reg[110]), .Z(n3098) );
  ANDN U3342 ( .A(n2507), .B(n2508), .Z(n3215) );
  XNOR U3343 ( .A(n2303), .B(round_reg[1218]), .Z(n2508) );
  XNOR U3344 ( .A(n2053), .B(round_reg[1291]), .Z(n2507) );
  XOR U3345 ( .A(n3216), .B(n2959), .Z(o[357]) );
  IV U3346 ( .A(n3100), .Z(n2959) );
  XNOR U3347 ( .A(n1909), .B(round_reg[109]), .Z(n3100) );
  ANDN U3348 ( .A(n2511), .B(n2512), .Z(n3216) );
  XNOR U3349 ( .A(n2311), .B(round_reg[1217]), .Z(n2512) );
  XNOR U3350 ( .A(n2056), .B(round_reg[1290]), .Z(n2511) );
  XOR U3351 ( .A(n3217), .B(n2961), .Z(o[356]) );
  XNOR U3352 ( .A(n1912), .B(round_reg[108]), .Z(n2961) );
  ANDN U3353 ( .A(n2515), .B(n2516), .Z(n3217) );
  XNOR U3354 ( .A(n2315), .B(round_reg[1216]), .Z(n2516) );
  XNOR U3355 ( .A(n2059), .B(round_reg[1289]), .Z(n2515) );
  XOR U3356 ( .A(n3218), .B(n3107), .Z(o[355]) );
  XNOR U3357 ( .A(n1915), .B(round_reg[107]), .Z(n3107) );
  ANDN U3358 ( .A(n2519), .B(n2520), .Z(n3218) );
  XNOR U3359 ( .A(n2319), .B(round_reg[1279]), .Z(n2520) );
  XNOR U3360 ( .A(n2062), .B(round_reg[1288]), .Z(n2519) );
  XOR U3361 ( .A(n3219), .B(n3109), .Z(o[354]) );
  XNOR U3362 ( .A(n1918), .B(round_reg[106]), .Z(n3109) );
  ANDN U3363 ( .A(n2523), .B(n2524), .Z(n3219) );
  XNOR U3364 ( .A(n2323), .B(round_reg[1278]), .Z(n2524) );
  XNOR U3365 ( .A(n2067), .B(round_reg[1287]), .Z(n2523) );
  XOR U3366 ( .A(n3220), .B(n3111), .Z(o[353]) );
  XNOR U3367 ( .A(n1921), .B(round_reg[105]), .Z(n3111) );
  ANDN U3368 ( .A(n2531), .B(n2532), .Z(n3220) );
  XNOR U3369 ( .A(n2327), .B(round_reg[1277]), .Z(n2532) );
  XNOR U3370 ( .A(n2070), .B(round_reg[1286]), .Z(n2531) );
  XOR U3371 ( .A(n3221), .B(n3113), .Z(o[352]) );
  XNOR U3372 ( .A(n1928), .B(round_reg[104]), .Z(n3113) );
  ANDN U3373 ( .A(n2535), .B(n2536), .Z(n3221) );
  XNOR U3374 ( .A(n2331), .B(round_reg[1276]), .Z(n2536) );
  XNOR U3375 ( .A(n2073), .B(round_reg[1285]), .Z(n2535) );
  XOR U3376 ( .A(n3222), .B(n2975), .Z(o[351]) );
  XNOR U3377 ( .A(n1931), .B(round_reg[103]), .Z(n2975) );
  ANDN U3378 ( .A(n2539), .B(n2540), .Z(n3222) );
  XNOR U3379 ( .A(n2335), .B(round_reg[1275]), .Z(n2540) );
  XNOR U3380 ( .A(n2076), .B(round_reg[1284]), .Z(n2539) );
  XOR U3381 ( .A(n3223), .B(n3116), .Z(o[350]) );
  XNOR U3382 ( .A(n1710), .B(round_reg[102]), .Z(n3116) );
  ANDN U3383 ( .A(n2543), .B(n2544), .Z(n3223) );
  XNOR U3384 ( .A(n2339), .B(round_reg[1274]), .Z(n2544) );
  XNOR U3385 ( .A(n2078), .B(round_reg[1283]), .Z(n2543) );
  XOR U3386 ( .A(n3224), .B(n1102), .Z(o[34]) );
  ANDN U3387 ( .A(n3225), .B(n1101), .Z(n3224) );
  XOR U3388 ( .A(n3226), .B(n3118), .Z(o[349]) );
  XNOR U3389 ( .A(n1713), .B(round_reg[101]), .Z(n3118) );
  ANDN U3390 ( .A(n2547), .B(n2548), .Z(n3226) );
  XNOR U3391 ( .A(n2343), .B(round_reg[1273]), .Z(n2548) );
  XNOR U3392 ( .A(n2080), .B(round_reg[1282]), .Z(n2547) );
  XOR U3393 ( .A(n3227), .B(n3120), .Z(o[348]) );
  XNOR U3394 ( .A(n1720), .B(round_reg[100]), .Z(n3120) );
  ANDN U3395 ( .A(n2551), .B(n2552), .Z(n3227) );
  XNOR U3396 ( .A(n2347), .B(round_reg[1272]), .Z(n2552) );
  XNOR U3397 ( .A(n2082), .B(round_reg[1281]), .Z(n2551) );
  XOR U3398 ( .A(n3228), .B(n3122), .Z(o[347]) );
  XNOR U3399 ( .A(n1723), .B(round_reg[99]), .Z(n3122) );
  ANDN U3400 ( .A(n2555), .B(n2556), .Z(n3228) );
  XNOR U3401 ( .A(n2355), .B(round_reg[1271]), .Z(n2556) );
  XNOR U3402 ( .A(n2084), .B(round_reg[1280]), .Z(n2555) );
  XOR U3403 ( .A(n3229), .B(n2985), .Z(o[346]) );
  XNOR U3404 ( .A(n1726), .B(round_reg[98]), .Z(n2985) );
  ANDN U3405 ( .A(n2559), .B(n2560), .Z(n3229) );
  XNOR U3406 ( .A(n2359), .B(round_reg[1270]), .Z(n2560) );
  XOR U3407 ( .A(n2086), .B(round_reg[1343]), .Z(n2559) );
  XOR U3408 ( .A(n3230), .B(n3129), .Z(o[345]) );
  XNOR U3409 ( .A(n1729), .B(round_reg[97]), .Z(n3129) );
  ANDN U3410 ( .A(n2563), .B(n2564), .Z(n3230) );
  XNOR U3411 ( .A(n2363), .B(round_reg[1269]), .Z(n2564) );
  XNOR U3412 ( .A(n2088), .B(round_reg[1342]), .Z(n2563) );
  XOR U3413 ( .A(n3231), .B(n2989), .Z(o[344]) );
  IV U3414 ( .A(n3131), .Z(n2989) );
  XNOR U3415 ( .A(n1732), .B(round_reg[96]), .Z(n3131) );
  ANDN U3416 ( .A(n2567), .B(n2568), .Z(n3231) );
  XNOR U3417 ( .A(n2367), .B(round_reg[1268]), .Z(n2568) );
  XNOR U3418 ( .A(n2095), .B(round_reg[1341]), .Z(n2567) );
  XOR U3419 ( .A(n3232), .B(n2991), .Z(o[343]) );
  IV U3420 ( .A(n3133), .Z(n2991) );
  XNOR U3421 ( .A(n1735), .B(round_reg[95]), .Z(n3133) );
  ANDN U3422 ( .A(n2578), .B(n2579), .Z(n3232) );
  XNOR U3423 ( .A(n2371), .B(round_reg[1267]), .Z(n2579) );
  XNOR U3424 ( .A(n2098), .B(round_reg[1340]), .Z(n2578) );
  XOR U3425 ( .A(n3233), .B(n2993), .Z(o[342]) );
  IV U3426 ( .A(n3135), .Z(n2993) );
  XNOR U3427 ( .A(n1738), .B(round_reg[94]), .Z(n3135) );
  ANDN U3428 ( .A(n2582), .B(n2583), .Z(n3233) );
  XNOR U3429 ( .A(n2375), .B(round_reg[1266]), .Z(n2583) );
  XNOR U3430 ( .A(n2101), .B(round_reg[1339]), .Z(n2582) );
  XOR U3431 ( .A(n3234), .B(n2999), .Z(o[341]) );
  IV U3432 ( .A(n3137), .Z(n2999) );
  XNOR U3433 ( .A(n1741), .B(round_reg[93]), .Z(n3137) );
  ANDN U3434 ( .A(n2586), .B(n2587), .Z(n3234) );
  XNOR U3435 ( .A(n2379), .B(round_reg[1265]), .Z(n2587) );
  XNOR U3436 ( .A(n2104), .B(round_reg[1338]), .Z(n2586) );
  XOR U3437 ( .A(n3235), .B(n3001), .Z(o[340]) );
  IV U3438 ( .A(n3139), .Z(n3001) );
  XNOR U3439 ( .A(n1744), .B(round_reg[92]), .Z(n3139) );
  ANDN U3440 ( .A(n2590), .B(n2591), .Z(n3235) );
  XNOR U3441 ( .A(n2383), .B(round_reg[1264]), .Z(n2591) );
  XNOR U3442 ( .A(n2107), .B(round_reg[1337]), .Z(n2590) );
  XNOR U3443 ( .A(n3236), .B(n1146), .Z(o[33]) );
  ANDN U3444 ( .A(n3237), .B(n1145), .Z(n3236) );
  XOR U3445 ( .A(n3238), .B(n3003), .Z(o[339]) );
  IV U3446 ( .A(n3141), .Z(n3003) );
  XNOR U3447 ( .A(n1747), .B(round_reg[91]), .Z(n3141) );
  ANDN U3448 ( .A(n2594), .B(n2595), .Z(n3238) );
  XNOR U3449 ( .A(n2387), .B(round_reg[1263]), .Z(n2595) );
  XNOR U3450 ( .A(n2110), .B(round_reg[1336]), .Z(n2594) );
  XOR U3451 ( .A(n3239), .B(n3005), .Z(o[338]) );
  XNOR U3452 ( .A(n1754), .B(round_reg[90]), .Z(n3005) );
  ANDN U3453 ( .A(n2598), .B(n2599), .Z(n3239) );
  XNOR U3454 ( .A(n2391), .B(round_reg[1262]), .Z(n2599) );
  XNOR U3455 ( .A(n1934), .B(round_reg[1335]), .Z(n2598) );
  XOR U3456 ( .A(n3240), .B(n3144), .Z(o[337]) );
  XNOR U3457 ( .A(n1757), .B(round_reg[89]), .Z(n3144) );
  ANDN U3458 ( .A(n2602), .B(n2603), .Z(n3240) );
  XNOR U3459 ( .A(n2112), .B(round_reg[1261]), .Z(n2603) );
  XNOR U3460 ( .A(n1936), .B(round_reg[1334]), .Z(n2602) );
  XOR U3461 ( .A(n3241), .B(n3146), .Z(o[336]) );
  XNOR U3462 ( .A(n1760), .B(round_reg[88]), .Z(n3146) );
  ANDN U3463 ( .A(n2606), .B(n2607), .Z(n3241) );
  XNOR U3464 ( .A(n2116), .B(round_reg[1260]), .Z(n2607) );
  XNOR U3465 ( .A(n1938), .B(round_reg[1333]), .Z(n2606) );
  XOR U3466 ( .A(n3242), .B(n3155), .Z(o[335]) );
  XNOR U3467 ( .A(n1763), .B(round_reg[87]), .Z(n3155) );
  ANDN U3468 ( .A(n2610), .B(n2611), .Z(n3242) );
  XNOR U3469 ( .A(n2120), .B(round_reg[1259]), .Z(n2611) );
  XNOR U3470 ( .A(n1940), .B(round_reg[1332]), .Z(n2610) );
  XOR U3471 ( .A(n3243), .B(n3157), .Z(o[334]) );
  XNOR U3472 ( .A(n1766), .B(round_reg[86]), .Z(n3157) );
  ANDN U3473 ( .A(n2614), .B(n2615), .Z(n3243) );
  XNOR U3474 ( .A(n2124), .B(round_reg[1258]), .Z(n2615) );
  XNOR U3475 ( .A(n1943), .B(round_reg[1331]), .Z(n2614) );
  XOR U3476 ( .A(n3244), .B(n3159), .Z(o[333]) );
  XNOR U3477 ( .A(n1769), .B(round_reg[85]), .Z(n3159) );
  ANDN U3478 ( .A(n2622), .B(n2623), .Z(n3244) );
  XNOR U3479 ( .A(n2135), .B(round_reg[1257]), .Z(n2623) );
  XNOR U3480 ( .A(n1946), .B(round_reg[1330]), .Z(n2622) );
  XOR U3481 ( .A(n3245), .B(n3161), .Z(o[332]) );
  XNOR U3482 ( .A(n1772), .B(round_reg[84]), .Z(n3161) );
  ANDN U3483 ( .A(n2626), .B(n2627), .Z(n3245) );
  XNOR U3484 ( .A(n2139), .B(round_reg[1256]), .Z(n2627) );
  XNOR U3485 ( .A(n1949), .B(round_reg[1329]), .Z(n2626) );
  XOR U3486 ( .A(n3246), .B(n3163), .Z(o[331]) );
  XNOR U3487 ( .A(n1775), .B(round_reg[83]), .Z(n3163) );
  ANDN U3488 ( .A(n2630), .B(n2631), .Z(n3246) );
  XNOR U3489 ( .A(n2143), .B(round_reg[1255]), .Z(n2631) );
  XNOR U3490 ( .A(n1952), .B(round_reg[1328]), .Z(n2630) );
  XOR U3491 ( .A(n3247), .B(n3025), .Z(o[330]) );
  XOR U3492 ( .A(n1778), .B(round_reg[82]), .Z(n3025) );
  ANDN U3493 ( .A(n2634), .B(n2635), .Z(n3247) );
  XNOR U3494 ( .A(n2147), .B(round_reg[1254]), .Z(n2635) );
  XNOR U3495 ( .A(n1959), .B(round_reg[1327]), .Z(n2634) );
  XNOR U3496 ( .A(n3248), .B(n1190), .Z(o[32]) );
  ANDN U3497 ( .A(n3249), .B(n1189), .Z(n3248) );
  XOR U3498 ( .A(n3250), .B(n3166), .Z(o[329]) );
  XOR U3499 ( .A(n1781), .B(round_reg[81]), .Z(n3166) );
  ANDN U3500 ( .A(n2638), .B(n2639), .Z(n3250) );
  XNOR U3501 ( .A(n2151), .B(round_reg[1253]), .Z(n2639) );
  XNOR U3502 ( .A(n1962), .B(round_reg[1326]), .Z(n2638) );
  XOR U3503 ( .A(n3251), .B(n3030), .Z(o[328]) );
  XOR U3504 ( .A(n1788), .B(round_reg[80]), .Z(n3030) );
  ANDN U3505 ( .A(n2642), .B(n2643), .Z(n3251) );
  XNOR U3506 ( .A(n2155), .B(round_reg[1252]), .Z(n2643) );
  XNOR U3507 ( .A(n1965), .B(round_reg[1325]), .Z(n2642) );
  XOR U3508 ( .A(n3252), .B(n3032), .Z(o[327]) );
  XOR U3509 ( .A(n1791), .B(round_reg[79]), .Z(n3032) );
  ANDN U3510 ( .A(n2646), .B(n2647), .Z(n3252) );
  XNOR U3511 ( .A(n2159), .B(round_reg[1251]), .Z(n2647) );
  XNOR U3512 ( .A(n1968), .B(round_reg[1324]), .Z(n2646) );
  XOR U3513 ( .A(n3253), .B(n3034), .Z(o[326]) );
  XOR U3514 ( .A(n1794), .B(round_reg[78]), .Z(n3034) );
  ANDN U3515 ( .A(n2650), .B(n2651), .Z(n3253) );
  XNOR U3516 ( .A(n2163), .B(round_reg[1250]), .Z(n2651) );
  XNOR U3517 ( .A(n1971), .B(round_reg[1323]), .Z(n2650) );
  XOR U3518 ( .A(n3254), .B(n3036), .Z(o[325]) );
  XOR U3519 ( .A(n1797), .B(round_reg[77]), .Z(n3036) );
  ANDN U3520 ( .A(n2654), .B(n2655), .Z(n3254) );
  XNOR U3521 ( .A(n2167), .B(round_reg[1249]), .Z(n2655) );
  XNOR U3522 ( .A(n1974), .B(round_reg[1322]), .Z(n2654) );
  XOR U3523 ( .A(n3255), .B(n3038), .Z(o[324]) );
  XOR U3524 ( .A(n1800), .B(round_reg[76]), .Z(n3038) );
  ANDN U3525 ( .A(n2658), .B(n2659), .Z(n3255) );
  XNOR U3526 ( .A(n2171), .B(round_reg[1248]), .Z(n2659) );
  XNOR U3527 ( .A(n1977), .B(round_reg[1321]), .Z(n2658) );
  XOR U3528 ( .A(n3256), .B(n3040), .Z(o[323]) );
  XOR U3529 ( .A(n1803), .B(round_reg[75]), .Z(n3040) );
  ANDN U3530 ( .A(n2666), .B(n2667), .Z(n3256) );
  XNOR U3531 ( .A(n2179), .B(round_reg[1247]), .Z(n2667) );
  XNOR U3532 ( .A(n1979), .B(round_reg[1320]), .Z(n2666) );
  XOR U3533 ( .A(n3257), .B(n3042), .Z(o[322]) );
  XOR U3534 ( .A(n1806), .B(round_reg[74]), .Z(n3042) );
  ANDN U3535 ( .A(n2670), .B(n2671), .Z(n3257) );
  XNOR U3536 ( .A(n2183), .B(round_reg[1246]), .Z(n2671) );
  XNOR U3537 ( .A(n1981), .B(round_reg[1319]), .Z(n2670) );
  XOR U3538 ( .A(n3258), .B(n3048), .Z(o[321]) );
  XOR U3539 ( .A(n1809), .B(round_reg[73]), .Z(n3048) );
  ANDN U3540 ( .A(n2674), .B(n2675), .Z(n3258) );
  XNOR U3541 ( .A(n2187), .B(round_reg[1245]), .Z(n2675) );
  XNOR U3542 ( .A(n1983), .B(round_reg[1318]), .Z(n2674) );
  XOR U3543 ( .A(n3259), .B(n3050), .Z(o[320]) );
  XOR U3544 ( .A(n1812), .B(round_reg[72]), .Z(n3050) );
  ANDN U3545 ( .A(n2678), .B(n2679), .Z(n3259) );
  XNOR U3546 ( .A(n2191), .B(round_reg[1244]), .Z(n2679) );
  XNOR U3547 ( .A(n1989), .B(round_reg[1317]), .Z(n2678) );
  XNOR U3548 ( .A(n3260), .B(n1234), .Z(o[31]) );
  ANDN U3549 ( .A(n3261), .B(n1233), .Z(n3260) );
  XNOR U3550 ( .A(n3262), .B(n2396), .Z(o[319]) );
  AND U3551 ( .A(n3263), .B(n3264), .Z(n3262) );
  XNOR U3552 ( .A(n3265), .B(n2440), .Z(o[318]) );
  AND U3553 ( .A(n3266), .B(n3267), .Z(n3265) );
  XNOR U3554 ( .A(n3268), .B(n2484), .Z(o[317]) );
  AND U3555 ( .A(n3269), .B(n3270), .Z(n3268) );
  XNOR U3556 ( .A(n3271), .B(n2528), .Z(o[316]) );
  AND U3557 ( .A(n3272), .B(n3273), .Z(n3271) );
  XNOR U3558 ( .A(n3274), .B(n2575), .Z(o[315]) );
  AND U3559 ( .A(n3275), .B(n3276), .Z(n3274) );
  XNOR U3560 ( .A(n3277), .B(n2619), .Z(o[314]) );
  AND U3561 ( .A(n3278), .B(n3279), .Z(n3277) );
  XNOR U3562 ( .A(n3280), .B(n2663), .Z(o[313]) );
  AND U3563 ( .A(n3281), .B(n3282), .Z(n3280) );
  XNOR U3564 ( .A(n3283), .B(n2701), .Z(o[312]) );
  AND U3565 ( .A(n3284), .B(n3285), .Z(n3283) );
  XNOR U3566 ( .A(n3286), .B(n2735), .Z(o[311]) );
  AND U3567 ( .A(n3287), .B(n3288), .Z(n3286) );
  XNOR U3568 ( .A(n3289), .B(n2764), .Z(o[310]) );
  AND U3569 ( .A(n3290), .B(n3291), .Z(n3289) );
  XNOR U3570 ( .A(n3292), .B(n1277), .Z(o[30]) );
  AND U3571 ( .A(n3293), .B(n3294), .Z(n3292) );
  XNOR U3572 ( .A(n3295), .B(n2798), .Z(o[309]) );
  AND U3573 ( .A(n3296), .B(n3297), .Z(n3295) );
  XNOR U3574 ( .A(n3298), .B(n2832), .Z(o[308]) );
  AND U3575 ( .A(n3299), .B(n3300), .Z(n3298) );
  XNOR U3576 ( .A(n3301), .B(n2865), .Z(o[307]) );
  AND U3577 ( .A(n3302), .B(n3303), .Z(n3301) );
  XNOR U3578 ( .A(n3304), .B(n2897), .Z(o[306]) );
  AND U3579 ( .A(n3305), .B(n3306), .Z(n3304) );
  XNOR U3580 ( .A(n3307), .B(n2924), .Z(o[305]) );
  AND U3581 ( .A(n3308), .B(n3309), .Z(n3307) );
  XNOR U3582 ( .A(n3310), .B(n2949), .Z(o[304]) );
  ANDN U3583 ( .A(n3311), .B(n2948), .Z(n3310) );
  XNOR U3584 ( .A(n3312), .B(n2973), .Z(o[303]) );
  ANDN U3585 ( .A(n3313), .B(n2972), .Z(n3312) );
  XNOR U3586 ( .A(n3314), .B(n2997), .Z(o[302]) );
  ANDN U3587 ( .A(n3315), .B(n2996), .Z(n3314) );
  XNOR U3588 ( .A(n3316), .B(n3021), .Z(o[301]) );
  ANDN U3589 ( .A(n3317), .B(n3020), .Z(n3316) );
  XNOR U3590 ( .A(n3318), .B(n3046), .Z(o[300]) );
  ANDN U3591 ( .A(n3319), .B(n3045), .Z(n3318) );
  XNOR U3592 ( .A(n3320), .B(n2264), .Z(o[2]) );
  AND U3593 ( .A(n3321), .B(n3322), .Z(n3320) );
  XNOR U3594 ( .A(n3323), .B(n1321), .Z(o[29]) );
  AND U3595 ( .A(n3324), .B(n3325), .Z(n3323) );
  XNOR U3596 ( .A(n3326), .B(n3062), .Z(o[299]) );
  ANDN U3597 ( .A(n3327), .B(n3061), .Z(n3326) );
  XNOR U3598 ( .A(n3328), .B(n3082), .Z(o[298]) );
  ANDN U3599 ( .A(n3329), .B(n3081), .Z(n3328) );
  XNOR U3600 ( .A(n3330), .B(n3105), .Z(o[297]) );
  ANDN U3601 ( .A(n3331), .B(n3104), .Z(n3330) );
  XOR U3602 ( .A(n3332), .B(n3127), .Z(o[296]) );
  ANDN U3603 ( .A(n3333), .B(n3126), .Z(n3332) );
  XOR U3604 ( .A(n3334), .B(n3153), .Z(o[295]) );
  ANDN U3605 ( .A(n3335), .B(n3152), .Z(n3334) );
  XOR U3606 ( .A(n3336), .B(n3173), .Z(o[294]) );
  ANDN U3607 ( .A(n3337), .B(n3172), .Z(n3336) );
  XOR U3608 ( .A(n3338), .B(n3187), .Z(o[293]) );
  ANDN U3609 ( .A(n3339), .B(n3186), .Z(n3338) );
  XOR U3610 ( .A(n3340), .B(n3201), .Z(o[292]) );
  ANDN U3611 ( .A(n3341), .B(n3200), .Z(n3340) );
  XOR U3612 ( .A(n3342), .B(n1057), .Z(o[291]) );
  XOR U3613 ( .A(n2204), .B(round_reg[1445]), .Z(n1057) );
  ANDN U3614 ( .A(n3343), .B(n3213), .Z(n3342) );
  XOR U3615 ( .A(n3344), .B(n1101), .Z(o[290]) );
  XOR U3616 ( .A(n2208), .B(round_reg[1444]), .Z(n1101) );
  ANDN U3617 ( .A(n3345), .B(n3225), .Z(n3344) );
  XNOR U3618 ( .A(n3346), .B(n1365), .Z(o[28]) );
  AND U3619 ( .A(n3347), .B(n3348), .Z(n3346) );
  XOR U3620 ( .A(n3349), .B(n1145), .Z(o[289]) );
  XNOR U3621 ( .A(n2212), .B(round_reg[1443]), .Z(n1145) );
  ANDN U3622 ( .A(n3350), .B(n3237), .Z(n3349) );
  XOR U3623 ( .A(n3351), .B(n1189), .Z(o[288]) );
  XOR U3624 ( .A(n2216), .B(round_reg[1442]), .Z(n1189) );
  ANDN U3625 ( .A(n3352), .B(n3249), .Z(n3351) );
  XOR U3626 ( .A(n3353), .B(n1233), .Z(o[287]) );
  XOR U3627 ( .A(n2224), .B(round_reg[1441]), .Z(n1233) );
  ANDN U3628 ( .A(n3354), .B(n3261), .Z(n3353) );
  XOR U3629 ( .A(n3355), .B(n1278), .Z(o[286]) );
  IV U3630 ( .A(n3294), .Z(n1278) );
  XNOR U3631 ( .A(n2228), .B(round_reg[1440]), .Z(n3294) );
  ANDN U3632 ( .A(n3356), .B(n3293), .Z(n3355) );
  XOR U3633 ( .A(n3357), .B(n1322), .Z(o[285]) );
  IV U3634 ( .A(n3325), .Z(n1322) );
  XNOR U3635 ( .A(n2232), .B(round_reg[1439]), .Z(n3325) );
  ANDN U3636 ( .A(n3358), .B(n3324), .Z(n3357) );
  XOR U3637 ( .A(n3359), .B(n1366), .Z(o[284]) );
  IV U3638 ( .A(n3348), .Z(n1366) );
  XNOR U3639 ( .A(n2236), .B(round_reg[1438]), .Z(n3348) );
  ANDN U3640 ( .A(n3360), .B(n3347), .Z(n3359) );
  XOR U3641 ( .A(n3361), .B(n1410), .Z(o[283]) );
  IV U3642 ( .A(n3362), .Z(n1410) );
  XOR U3643 ( .A(n3365), .B(n1454), .Z(o[282]) );
  IV U3644 ( .A(n3366), .Z(n1454) );
  XOR U3645 ( .A(n3369), .B(n1502), .Z(o[281]) );
  IV U3646 ( .A(n3370), .Z(n1502) );
  XOR U3647 ( .A(n3373), .B(n1534), .Z(o[280]) );
  IV U3648 ( .A(n3374), .Z(n1534) );
  XNOR U3649 ( .A(n3377), .B(n1409), .Z(o[27]) );
  AND U3650 ( .A(n3364), .B(n3362), .Z(n3377) );
  XNOR U3651 ( .A(n2240), .B(round_reg[1437]), .Z(n3362) );
  XOR U3652 ( .A(n3378), .B(n1564), .Z(o[279]) );
  IV U3653 ( .A(n3379), .Z(n1564) );
  ANDN U3654 ( .A(n3380), .B(n3381), .Z(n3378) );
  XOR U3655 ( .A(n3382), .B(n1589), .Z(o[278]) );
  IV U3656 ( .A(n3383), .Z(n1589) );
  ANDN U3657 ( .A(n3384), .B(n3385), .Z(n3382) );
  XOR U3658 ( .A(n3386), .B(n1622), .Z(o[277]) );
  IV U3659 ( .A(n3387), .Z(n1622) );
  ANDN U3660 ( .A(n3388), .B(n3389), .Z(n3386) );
  XOR U3661 ( .A(n3390), .B(n1656), .Z(o[276]) );
  IV U3662 ( .A(n3391), .Z(n1656) );
  AND U3663 ( .A(n3392), .B(n3393), .Z(n3390) );
  XOR U3664 ( .A(n3394), .B(n1690), .Z(o[275]) );
  IV U3665 ( .A(n3395), .Z(n1690) );
  AND U3666 ( .A(n3396), .B(n3397), .Z(n3394) );
  XOR U3667 ( .A(n3398), .B(n1718), .Z(o[274]) );
  IV U3668 ( .A(n3399), .Z(n1718) );
  AND U3669 ( .A(n3400), .B(n3401), .Z(n3398) );
  XOR U3670 ( .A(n3402), .B(n1752), .Z(o[273]) );
  IV U3671 ( .A(n3403), .Z(n1752) );
  AND U3672 ( .A(n3404), .B(n3405), .Z(n3402) );
  XOR U3673 ( .A(n3406), .B(n1786), .Z(o[272]) );
  IV U3674 ( .A(n3407), .Z(n1786) );
  AND U3675 ( .A(n3408), .B(n3409), .Z(n3406) );
  XOR U3676 ( .A(n3410), .B(n1824), .Z(o[271]) );
  IV U3677 ( .A(n3411), .Z(n1824) );
  AND U3678 ( .A(n3412), .B(n3413), .Z(n3410) );
  XOR U3679 ( .A(n3414), .B(n1858), .Z(o[270]) );
  IV U3680 ( .A(n3415), .Z(n1858) );
  AND U3681 ( .A(n3416), .B(n3417), .Z(n3414) );
  XNOR U3682 ( .A(n3418), .B(n1453), .Z(o[26]) );
  AND U3683 ( .A(n3368), .B(n3366), .Z(n3418) );
  XNOR U3684 ( .A(n2244), .B(round_reg[1436]), .Z(n3366) );
  AND U3685 ( .A(n3420), .B(n3421), .Z(n3419) );
  AND U3686 ( .A(n3423), .B(n3424), .Z(n3422) );
  AND U3687 ( .A(n3426), .B(n3427), .Z(n3425) );
  AND U3688 ( .A(n3429), .B(n3430), .Z(n3428) );
  XOR U3689 ( .A(n3431), .B(n1054), .Z(o[265]) );
  XOR U3690 ( .A(n2320), .B(round_reg[1419]), .Z(n1054) );
  NOR U3691 ( .A(n3432), .B(n1053), .Z(n3431) );
  XOR U3692 ( .A(n3433), .B(n1498), .Z(o[264]) );
  XOR U3693 ( .A(n2324), .B(round_reg[1418]), .Z(n1498) );
  AND U3694 ( .A(n3434), .B(n1497), .Z(n3433) );
  IV U3695 ( .A(n3435), .Z(n1497) );
  XOR U3696 ( .A(n3436), .B(n1820), .Z(o[263]) );
  XOR U3697 ( .A(n2328), .B(round_reg[1417]), .Z(n1820) );
  AND U3698 ( .A(n3437), .B(n1819), .Z(n3436) );
  IV U3699 ( .A(n3438), .Z(n1819) );
  XOR U3700 ( .A(n3439), .B(n2093), .Z(o[262]) );
  IV U3701 ( .A(n2129), .Z(n2093) );
  XNOR U3702 ( .A(n2332), .B(round_reg[1416]), .Z(n2129) );
  XOR U3703 ( .A(n3441), .B(n2133), .Z(o[261]) );
  IV U3704 ( .A(n2572), .Z(n2133) );
  XNOR U3705 ( .A(n2336), .B(round_reg[1415]), .Z(n2572) );
  XOR U3706 ( .A(n3443), .B(n2177), .Z(o[260]) );
  IV U3707 ( .A(n2921), .Z(n2177) );
  XNOR U3708 ( .A(n2340), .B(round_reg[1414]), .Z(n2921) );
  XNOR U3709 ( .A(n3445), .B(n1501), .Z(o[25]) );
  AND U3710 ( .A(n3372), .B(n3370), .Z(n3445) );
  XNOR U3711 ( .A(n2248), .B(round_reg[1435]), .Z(n3370) );
  XOR U3712 ( .A(n3446), .B(n2221), .Z(o[259]) );
  IV U3713 ( .A(n3149), .Z(n2221) );
  XNOR U3714 ( .A(n2344), .B(round_reg[1413]), .Z(n3149) );
  XOR U3715 ( .A(n3448), .B(n2265), .Z(o[258]) );
  IV U3716 ( .A(n3322), .Z(n2265) );
  XNOR U3717 ( .A(n2348), .B(round_reg[1412]), .Z(n3322) );
  ANDN U3718 ( .A(n3449), .B(n3321), .Z(n3448) );
  XOR U3719 ( .A(n3450), .B(n2309), .Z(o[257]) );
  IV U3720 ( .A(n3451), .Z(n2309) );
  XOR U3721 ( .A(n3454), .B(n2352), .Z(o[256]) );
  IV U3722 ( .A(n3455), .Z(n2352) );
  XOR U3723 ( .A(n3458), .B(n2397), .Z(o[255]) );
  IV U3724 ( .A(n3264), .Z(n2397) );
  XNOR U3725 ( .A(n1812), .B(round_reg[1032]), .Z(n3264) );
  XOR U3726 ( .A(n3460), .B(n2441), .Z(o[254]) );
  IV U3727 ( .A(n3267), .Z(n2441) );
  XNOR U3728 ( .A(n1815), .B(round_reg[1031]), .Z(n3267) );
  XOR U3729 ( .A(n3462), .B(n2485), .Z(o[253]) );
  IV U3730 ( .A(n3270), .Z(n2485) );
  XNOR U3731 ( .A(n1826), .B(round_reg[1030]), .Z(n3270) );
  XOR U3732 ( .A(n3464), .B(n2529), .Z(o[252]) );
  IV U3733 ( .A(n3273), .Z(n2529) );
  XNOR U3734 ( .A(n1829), .B(round_reg[1029]), .Z(n3273) );
  XOR U3735 ( .A(n3466), .B(n2576), .Z(o[251]) );
  IV U3736 ( .A(n3276), .Z(n2576) );
  XNOR U3737 ( .A(n1832), .B(round_reg[1028]), .Z(n3276) );
  XOR U3738 ( .A(n3468), .B(n2620), .Z(o[250]) );
  IV U3739 ( .A(n3279), .Z(n2620) );
  XNOR U3740 ( .A(n1835), .B(round_reg[1027]), .Z(n3279) );
  ANDN U3741 ( .A(n3469), .B(n3278), .Z(n3468) );
  XNOR U3742 ( .A(n3470), .B(n1533), .Z(o[24]) );
  AND U3743 ( .A(n3376), .B(n3374), .Z(n3470) );
  XNOR U3744 ( .A(n2252), .B(round_reg[1434]), .Z(n3374) );
  XOR U3745 ( .A(n3471), .B(n2664), .Z(o[249]) );
  IV U3746 ( .A(n3282), .Z(n2664) );
  XNOR U3747 ( .A(n1838), .B(round_reg[1026]), .Z(n3282) );
  ANDN U3748 ( .A(n3472), .B(n3281), .Z(n3471) );
  XOR U3749 ( .A(n3473), .B(n2702), .Z(o[248]) );
  IV U3750 ( .A(n3285), .Z(n2702) );
  XNOR U3751 ( .A(n1841), .B(round_reg[1025]), .Z(n3285) );
  ANDN U3752 ( .A(n3474), .B(n3284), .Z(n3473) );
  XOR U3753 ( .A(n3475), .B(n2736), .Z(o[247]) );
  IV U3754 ( .A(n3288), .Z(n2736) );
  XNOR U3755 ( .A(n1844), .B(round_reg[1024]), .Z(n3288) );
  ANDN U3756 ( .A(n3476), .B(n3287), .Z(n3475) );
  XOR U3757 ( .A(n3477), .B(n2765), .Z(o[246]) );
  IV U3758 ( .A(n3291), .Z(n2765) );
  XNOR U3759 ( .A(n1847), .B(round_reg[1087]), .Z(n3291) );
  ANDN U3760 ( .A(n3478), .B(n3290), .Z(n3477) );
  XOR U3761 ( .A(n3479), .B(n2799), .Z(o[245]) );
  IV U3762 ( .A(n3297), .Z(n2799) );
  XNOR U3763 ( .A(n1850), .B(round_reg[1086]), .Z(n3297) );
  ANDN U3764 ( .A(n3480), .B(n3296), .Z(n3479) );
  XOR U3765 ( .A(n3481), .B(n2833), .Z(o[244]) );
  IV U3766 ( .A(n3300), .Z(n2833) );
  XNOR U3767 ( .A(n1853), .B(round_reg[1085]), .Z(n3300) );
  ANDN U3768 ( .A(n3482), .B(n3299), .Z(n3481) );
  XOR U3769 ( .A(n3483), .B(n2866), .Z(o[243]) );
  IV U3770 ( .A(n3303), .Z(n2866) );
  XNOR U3771 ( .A(n1860), .B(round_reg[1084]), .Z(n3303) );
  ANDN U3772 ( .A(n3484), .B(n3302), .Z(n3483) );
  XOR U3773 ( .A(n3485), .B(n2898), .Z(o[242]) );
  IV U3774 ( .A(n3306), .Z(n2898) );
  XNOR U3775 ( .A(n1863), .B(round_reg[1083]), .Z(n3306) );
  ANDN U3776 ( .A(n3486), .B(n3305), .Z(n3485) );
  XOR U3777 ( .A(n3487), .B(n2925), .Z(o[241]) );
  IV U3778 ( .A(n3309), .Z(n2925) );
  XNOR U3779 ( .A(n1866), .B(round_reg[1082]), .Z(n3309) );
  ANDN U3780 ( .A(n3488), .B(n3308), .Z(n3487) );
  XOR U3781 ( .A(n3489), .B(n2948), .Z(o[240]) );
  XOR U3782 ( .A(n1869), .B(round_reg[1081]), .Z(n2948) );
  ANDN U3783 ( .A(n3490), .B(n3311), .Z(n3489) );
  XNOR U3784 ( .A(n3491), .B(n1563), .Z(o[23]) );
  AND U3785 ( .A(n3381), .B(n3379), .Z(n3491) );
  XNOR U3786 ( .A(n2256), .B(round_reg[1433]), .Z(n3379) );
  XOR U3787 ( .A(n3492), .B(n2972), .Z(o[239]) );
  XOR U3788 ( .A(n1872), .B(round_reg[1080]), .Z(n2972) );
  ANDN U3789 ( .A(n3493), .B(n3313), .Z(n3492) );
  XOR U3790 ( .A(n3494), .B(n2996), .Z(o[238]) );
  XOR U3791 ( .A(n1875), .B(round_reg[1079]), .Z(n2996) );
  ANDN U3792 ( .A(n3495), .B(n3315), .Z(n3494) );
  XOR U3793 ( .A(n3496), .B(n3020), .Z(o[237]) );
  XOR U3794 ( .A(n1878), .B(round_reg[1078]), .Z(n3020) );
  ANDN U3795 ( .A(n3497), .B(n3317), .Z(n3496) );
  XOR U3796 ( .A(n3498), .B(n3045), .Z(o[236]) );
  XOR U3797 ( .A(n1881), .B(round_reg[1077]), .Z(n3045) );
  ANDN U3798 ( .A(n3499), .B(n3319), .Z(n3498) );
  XOR U3799 ( .A(n3500), .B(n3061), .Z(o[235]) );
  XOR U3800 ( .A(n1884), .B(round_reg[1076]), .Z(n3061) );
  ANDN U3801 ( .A(n3501), .B(n3327), .Z(n3500) );
  XOR U3802 ( .A(n3502), .B(n3081), .Z(o[234]) );
  XOR U3803 ( .A(n1887), .B(round_reg[1075]), .Z(n3081) );
  ANDN U3804 ( .A(n3503), .B(n3329), .Z(n3502) );
  XOR U3805 ( .A(n3504), .B(n3104), .Z(o[233]) );
  XOR U3806 ( .A(n1894), .B(round_reg[1074]), .Z(n3104) );
  ANDN U3807 ( .A(n3505), .B(n3331), .Z(n3504) );
  XOR U3808 ( .A(n3506), .B(n3126), .Z(o[232]) );
  XOR U3809 ( .A(n1897), .B(round_reg[1073]), .Z(n3126) );
  ANDN U3810 ( .A(n3507), .B(n3333), .Z(n3506) );
  XOR U3811 ( .A(n3508), .B(n3152), .Z(o[231]) );
  XOR U3812 ( .A(n1900), .B(round_reg[1072]), .Z(n3152) );
  ANDN U3813 ( .A(n3509), .B(n3335), .Z(n3508) );
  XOR U3814 ( .A(n3510), .B(n3172), .Z(o[230]) );
  XOR U3815 ( .A(n1903), .B(round_reg[1071]), .Z(n3172) );
  ANDN U3816 ( .A(n3511), .B(n3337), .Z(n3510) );
  XNOR U3817 ( .A(n3512), .B(n1588), .Z(o[22]) );
  AND U3818 ( .A(n3385), .B(n3383), .Z(n3512) );
  XNOR U3819 ( .A(n2260), .B(round_reg[1432]), .Z(n3383) );
  XOR U3820 ( .A(n3513), .B(n3186), .Z(o[229]) );
  XOR U3821 ( .A(n1906), .B(round_reg[1070]), .Z(n3186) );
  ANDN U3822 ( .A(n3514), .B(n3339), .Z(n3513) );
  XOR U3823 ( .A(n3515), .B(n3200), .Z(o[228]) );
  XOR U3824 ( .A(n1909), .B(round_reg[1069]), .Z(n3200) );
  ANDN U3825 ( .A(n3516), .B(n3341), .Z(n3515) );
  XOR U3826 ( .A(n3517), .B(n3213), .Z(o[227]) );
  XNOR U3827 ( .A(n1912), .B(round_reg[1068]), .Z(n3213) );
  ANDN U3828 ( .A(n1056), .B(n3343), .Z(n3517) );
  XOR U3829 ( .A(n3518), .B(n3225), .Z(o[226]) );
  XNOR U3830 ( .A(n1915), .B(round_reg[1067]), .Z(n3225) );
  ANDN U3831 ( .A(n1100), .B(n3345), .Z(n3518) );
  XOR U3832 ( .A(n3519), .B(n3237), .Z(o[225]) );
  XNOR U3833 ( .A(n1918), .B(round_reg[1066]), .Z(n3237) );
  ANDN U3834 ( .A(n1144), .B(n3350), .Z(n3519) );
  XOR U3835 ( .A(n3520), .B(n3249), .Z(o[224]) );
  XNOR U3836 ( .A(n1921), .B(round_reg[1065]), .Z(n3249) );
  NOR U3837 ( .A(n1188), .B(n3352), .Z(n3520) );
  XOR U3838 ( .A(n3521), .B(n3261), .Z(o[223]) );
  XNOR U3839 ( .A(n1928), .B(round_reg[1064]), .Z(n3261) );
  XOR U3840 ( .A(n3522), .B(n3293), .Z(o[222]) );
  XNOR U3841 ( .A(n1931), .B(round_reg[1063]), .Z(n3293) );
  XOR U3842 ( .A(n3523), .B(n3324), .Z(o[221]) );
  XNOR U3843 ( .A(n1710), .B(round_reg[1062]), .Z(n3324) );
  XOR U3844 ( .A(n3524), .B(n3347), .Z(o[220]) );
  XNOR U3845 ( .A(n1713), .B(round_reg[1061]), .Z(n3347) );
  XNOR U3846 ( .A(n3525), .B(n1621), .Z(o[21]) );
  AND U3847 ( .A(n3389), .B(n3387), .Z(n3525) );
  XNOR U3848 ( .A(n2268), .B(round_reg[1431]), .Z(n3387) );
  XOR U3849 ( .A(n3526), .B(n3364), .Z(o[219]) );
  XNOR U3850 ( .A(n1720), .B(round_reg[1060]), .Z(n3364) );
  NOR U3851 ( .A(n3363), .B(n1408), .Z(n3526) );
  XOR U3852 ( .A(n3527), .B(n3368), .Z(o[218]) );
  XNOR U3853 ( .A(n1723), .B(round_reg[1059]), .Z(n3368) );
  NOR U3854 ( .A(n3367), .B(n1452), .Z(n3527) );
  XOR U3855 ( .A(n3528), .B(n3372), .Z(o[217]) );
  XNOR U3856 ( .A(n1726), .B(round_reg[1058]), .Z(n3372) );
  NOR U3857 ( .A(n3371), .B(n1500), .Z(n3528) );
  XOR U3858 ( .A(n3529), .B(n3376), .Z(o[216]) );
  XNOR U3859 ( .A(n1729), .B(round_reg[1057]), .Z(n3376) );
  NOR U3860 ( .A(n3375), .B(n1532), .Z(n3529) );
  XOR U3861 ( .A(n3530), .B(n3381), .Z(o[215]) );
  XOR U3862 ( .A(n1732), .B(round_reg[1056]), .Z(n3381) );
  NOR U3863 ( .A(n3380), .B(n1562), .Z(n3530) );
  XOR U3864 ( .A(n3531), .B(n3385), .Z(o[214]) );
  XOR U3865 ( .A(n1735), .B(round_reg[1055]), .Z(n3385) );
  NOR U3866 ( .A(n3384), .B(n1587), .Z(n3531) );
  XOR U3867 ( .A(n3532), .B(n3389), .Z(o[213]) );
  XOR U3868 ( .A(n1738), .B(round_reg[1054]), .Z(n3389) );
  NOR U3869 ( .A(n3388), .B(n1620), .Z(n3532) );
  XNOR U3870 ( .A(n3533), .B(n3393), .Z(o[212]) );
  NOR U3871 ( .A(n3392), .B(n1654), .Z(n3533) );
  XNOR U3872 ( .A(n3534), .B(n3397), .Z(o[211]) );
  NOR U3873 ( .A(n3396), .B(n1688), .Z(n3534) );
  XNOR U3874 ( .A(n3535), .B(n3400), .Z(o[210]) );
  ANDN U3875 ( .A(n3536), .B(n1716), .Z(n3535) );
  XNOR U3876 ( .A(n3537), .B(n1655), .Z(o[20]) );
  ANDN U3877 ( .A(n3391), .B(n3393), .Z(n3537) );
  XNOR U3878 ( .A(n1741), .B(round_reg[1053]), .Z(n3393) );
  XNOR U3879 ( .A(n2272), .B(round_reg[1430]), .Z(n3391) );
  XNOR U3880 ( .A(n3538), .B(n3404), .Z(o[209]) );
  ANDN U3881 ( .A(n3539), .B(n1750), .Z(n3538) );
  XNOR U3882 ( .A(n3540), .B(n3408), .Z(o[208]) );
  XNOR U3883 ( .A(n3541), .B(n3412), .Z(o[207]) );
  XNOR U3884 ( .A(n3542), .B(n3416), .Z(o[206]) );
  XNOR U3885 ( .A(n3543), .B(n3420), .Z(o[205]) );
  XNOR U3886 ( .A(n3544), .B(n3423), .Z(o[204]) );
  XNOR U3887 ( .A(n3545), .B(n3426), .Z(o[203]) );
  XNOR U3888 ( .A(n3546), .B(n3429), .Z(o[202]) );
  XOR U3889 ( .A(n3547), .B(n1053), .Z(o[201]) );
  XOR U3890 ( .A(n1778), .B(round_reg[1042]), .Z(n1053) );
  ANDN U3891 ( .A(n3432), .B(n2009), .Z(n3547) );
  IV U3892 ( .A(n3548), .Z(n3432) );
  XOR U3893 ( .A(n3549), .B(n3435), .Z(o[200]) );
  XOR U3894 ( .A(n1781), .B(round_reg[1041]), .Z(n3435) );
  XNOR U3895 ( .A(n3550), .B(n2308), .Z(o[1]) );
  AND U3896 ( .A(n3453), .B(n3451), .Z(n3550) );
  XNOR U3897 ( .A(n2356), .B(round_reg[1411]), .Z(n3451) );
  XNOR U3898 ( .A(n3551), .B(n1689), .Z(o[19]) );
  ANDN U3899 ( .A(n3395), .B(n3397), .Z(n3551) );
  XNOR U3900 ( .A(n1744), .B(round_reg[1052]), .Z(n3397) );
  XNOR U3901 ( .A(n2276), .B(round_reg[1429]), .Z(n3395) );
  XOR U3902 ( .A(n3552), .B(n3438), .Z(o[199]) );
  XOR U3903 ( .A(n1788), .B(round_reg[1040]), .Z(n3438) );
  XOR U3904 ( .A(n3553), .B(n2128), .Z(o[198]) );
  XOR U3905 ( .A(n1791), .B(round_reg[1039]), .Z(n2128) );
  XOR U3906 ( .A(n3554), .B(n2571), .Z(o[197]) );
  XOR U3907 ( .A(n1794), .B(round_reg[1038]), .Z(n2571) );
  XOR U3908 ( .A(n3555), .B(n2920), .Z(o[196]) );
  XOR U3909 ( .A(n1797), .B(round_reg[1037]), .Z(n2920) );
  XOR U3910 ( .A(n3556), .B(n3148), .Z(o[195]) );
  XOR U3911 ( .A(n1800), .B(round_reg[1036]), .Z(n3148) );
  XOR U3912 ( .A(n3557), .B(n3321), .Z(o[194]) );
  XOR U3913 ( .A(n1803), .B(round_reg[1035]), .Z(n3321) );
  XOR U3914 ( .A(n3558), .B(n3453), .Z(o[193]) );
  XOR U3915 ( .A(n1806), .B(round_reg[1034]), .Z(n3453) );
  XOR U3916 ( .A(n3559), .B(n3457), .Z(o[192]) );
  XOR U3917 ( .A(n3560), .B(n3263), .Z(o[191]) );
  XOR U3918 ( .A(n2018), .B(round_reg[664]), .Z(n3263) );
  XOR U3919 ( .A(n3561), .B(n3266), .Z(o[190]) );
  XOR U3920 ( .A(n2020), .B(round_reg[663]), .Z(n3266) );
  XNOR U3921 ( .A(n3562), .B(n1717), .Z(o[18]) );
  ANDN U3922 ( .A(n3399), .B(n3400), .Z(n3562) );
  XNOR U3923 ( .A(n1747), .B(round_reg[1051]), .Z(n3400) );
  XNOR U3924 ( .A(n2280), .B(round_reg[1428]), .Z(n3399) );
  XOR U3925 ( .A(n3563), .B(n3269), .Z(o[189]) );
  XOR U3926 ( .A(n2022), .B(round_reg[662]), .Z(n3269) );
  XOR U3927 ( .A(n3564), .B(n3272), .Z(o[188]) );
  XOR U3928 ( .A(n2024), .B(round_reg[661]), .Z(n3272) );
  XOR U3929 ( .A(n3565), .B(n3275), .Z(o[187]) );
  XOR U3930 ( .A(n2026), .B(round_reg[660]), .Z(n3275) );
  XOR U3931 ( .A(n3566), .B(n3278), .Z(o[186]) );
  XOR U3932 ( .A(n2028), .B(round_reg[659]), .Z(n3278) );
  XOR U3933 ( .A(n3567), .B(n3281), .Z(o[185]) );
  XOR U3934 ( .A(n2031), .B(round_reg[658]), .Z(n3281) );
  XOR U3935 ( .A(n3568), .B(n3284), .Z(o[184]) );
  XOR U3936 ( .A(n2036), .B(round_reg[657]), .Z(n3284) );
  XOR U3937 ( .A(n3569), .B(n3287), .Z(o[183]) );
  XOR U3938 ( .A(n2039), .B(round_reg[656]), .Z(n3287) );
  XOR U3939 ( .A(n3570), .B(n3290), .Z(o[182]) );
  XOR U3940 ( .A(n2042), .B(round_reg[655]), .Z(n3290) );
  XOR U3941 ( .A(n3571), .B(n3296), .Z(o[181]) );
  XOR U3942 ( .A(n2044), .B(round_reg[654]), .Z(n3296) );
  XOR U3943 ( .A(n3572), .B(n3299), .Z(o[180]) );
  XOR U3944 ( .A(n2047), .B(round_reg[653]), .Z(n3299) );
  XNOR U3945 ( .A(n3573), .B(n1751), .Z(o[17]) );
  ANDN U3946 ( .A(n3403), .B(n3404), .Z(n3573) );
  XOR U3947 ( .A(n1754), .B(round_reg[1050]), .Z(n3404) );
  XNOR U3948 ( .A(n2284), .B(round_reg[1427]), .Z(n3403) );
  XOR U3949 ( .A(n3574), .B(n3302), .Z(o[179]) );
  XOR U3950 ( .A(n2050), .B(round_reg[652]), .Z(n3302) );
  XOR U3951 ( .A(n3575), .B(n3305), .Z(o[178]) );
  XOR U3952 ( .A(n2053), .B(round_reg[651]), .Z(n3305) );
  XOR U3953 ( .A(n3576), .B(n3308), .Z(o[177]) );
  XOR U3954 ( .A(n2056), .B(round_reg[650]), .Z(n3308) );
  XOR U3955 ( .A(n3577), .B(n3311), .Z(o[176]) );
  XOR U3956 ( .A(n2059), .B(round_reg[649]), .Z(n3311) );
  XOR U3957 ( .A(n3578), .B(n3313), .Z(o[175]) );
  XOR U3958 ( .A(n2062), .B(round_reg[648]), .Z(n3313) );
  XOR U3959 ( .A(n3579), .B(n3315), .Z(o[174]) );
  XOR U3960 ( .A(n2067), .B(round_reg[647]), .Z(n3315) );
  ANDN U3961 ( .A(n3580), .B(n2995), .Z(n3579) );
  XOR U3962 ( .A(n3581), .B(n3317), .Z(o[173]) );
  XOR U3963 ( .A(n2070), .B(round_reg[646]), .Z(n3317) );
  XOR U3964 ( .A(n3582), .B(n3319), .Z(o[172]) );
  XOR U3965 ( .A(n2073), .B(round_reg[645]), .Z(n3319) );
  XOR U3966 ( .A(n3583), .B(n3327), .Z(o[171]) );
  XOR U3967 ( .A(n2076), .B(round_reg[644]), .Z(n3327) );
  XOR U3968 ( .A(n3584), .B(n3329), .Z(o[170]) );
  XOR U3969 ( .A(n2078), .B(round_reg[643]), .Z(n3329) );
  XNOR U3970 ( .A(n3585), .B(n1785), .Z(o[16]) );
  ANDN U3971 ( .A(n3407), .B(n3408), .Z(n3585) );
  XOR U3972 ( .A(n1757), .B(round_reg[1049]), .Z(n3408) );
  XNOR U3973 ( .A(n2288), .B(round_reg[1426]), .Z(n3407) );
  XOR U3974 ( .A(n3586), .B(n3331), .Z(o[169]) );
  XOR U3975 ( .A(n2080), .B(round_reg[642]), .Z(n3331) );
  XOR U3976 ( .A(n3587), .B(n3333), .Z(o[168]) );
  XOR U3977 ( .A(n2082), .B(round_reg[641]), .Z(n3333) );
  XOR U3978 ( .A(n3588), .B(n3335), .Z(o[167]) );
  XOR U3979 ( .A(n2084), .B(round_reg[640]), .Z(n3335) );
  XOR U3980 ( .A(n3589), .B(n3337), .Z(o[166]) );
  XNOR U3981 ( .A(n2086), .B(round_reg[703]), .Z(n3337) );
  XOR U3982 ( .A(n3590), .B(n3339), .Z(o[165]) );
  XOR U3983 ( .A(n2088), .B(round_reg[702]), .Z(n3339) );
  XOR U3984 ( .A(n3591), .B(n3341), .Z(o[164]) );
  XOR U3985 ( .A(n2095), .B(round_reg[701]), .Z(n3341) );
  XOR U3986 ( .A(n3592), .B(n3343), .Z(o[163]) );
  XOR U3987 ( .A(n2098), .B(round_reg[700]), .Z(n3343) );
  ANDN U3988 ( .A(n1058), .B(n1056), .Z(n3592) );
  XOR U3989 ( .A(n2339), .B(round_reg[634]), .Z(n1056) );
  XOR U3990 ( .A(n2245), .B(round_reg[225]), .Z(n1058) );
  XOR U3991 ( .A(n3593), .B(n3345), .Z(o[162]) );
  XOR U3992 ( .A(n2101), .B(round_reg[699]), .Z(n3345) );
  ANDN U3993 ( .A(n1102), .B(n1100), .Z(n3593) );
  XOR U3994 ( .A(n2343), .B(round_reg[633]), .Z(n1100) );
  XNOR U3995 ( .A(n2249), .B(round_reg[224]), .Z(n1102) );
  XOR U3996 ( .A(n3594), .B(n3350), .Z(o[161]) );
  XOR U3997 ( .A(n2104), .B(round_reg[698]), .Z(n3350) );
  NOR U3998 ( .A(n1146), .B(n1144), .Z(n3594) );
  XOR U3999 ( .A(n2347), .B(round_reg[632]), .Z(n1144) );
  XOR U4000 ( .A(n2253), .B(round_reg[223]), .Z(n1146) );
  XOR U4001 ( .A(n3595), .B(n3352), .Z(o[160]) );
  XOR U4002 ( .A(n2107), .B(round_reg[697]), .Z(n3352) );
  ANDN U4003 ( .A(n1188), .B(n1190), .Z(n3595) );
  XOR U4004 ( .A(n2257), .B(round_reg[222]), .Z(n1190) );
  XNOR U4005 ( .A(n2355), .B(round_reg[631]), .Z(n1188) );
  XNOR U4006 ( .A(n3596), .B(n1823), .Z(o[15]) );
  ANDN U4007 ( .A(n3411), .B(n3412), .Z(n3596) );
  XOR U4008 ( .A(n1760), .B(round_reg[1048]), .Z(n3412) );
  XNOR U4009 ( .A(n2292), .B(round_reg[1425]), .Z(n3411) );
  XOR U4010 ( .A(n3597), .B(n3354), .Z(o[159]) );
  XOR U4011 ( .A(n2110), .B(round_reg[696]), .Z(n3354) );
  ANDN U4012 ( .A(n1232), .B(n1234), .Z(n3597) );
  XOR U4013 ( .A(n2261), .B(round_reg[221]), .Z(n1234) );
  XNOR U4014 ( .A(n2359), .B(round_reg[630]), .Z(n1232) );
  XNOR U4015 ( .A(n3598), .B(n3599), .Z(o[1599]) );
  XOR U4016 ( .A(n3600), .B(n3601), .Z(n3598) );
  NAND U4017 ( .A(n3604), .B(n3605), .Z(n3600) );
  AND U4018 ( .A(n3606), .B(n3607), .Z(n3605) );
  NOR U4019 ( .A(rc_i[2]), .B(rc_i[3]), .Z(n3607) );
  NOR U4020 ( .A(rc_i[17]), .B(rc_i[19]), .Z(n3606) );
  AND U4021 ( .A(n3608), .B(n3609), .Z(n3604) );
  NOR U4022 ( .A(rc_i[16]), .B(n3610), .Z(n3609) );
  ANDN U4023 ( .A(n3611), .B(n3612), .Z(n3608) );
  XNOR U4024 ( .A(n3613), .B(n3614), .Z(o[1598]) );
  XNOR U4025 ( .A(n3617), .B(n3618), .Z(o[1597]) );
  XNOR U4026 ( .A(n3621), .B(n3622), .Z(o[1596]) );
  XNOR U4027 ( .A(n3625), .B(n3626), .Z(o[1595]) );
  XOR U4028 ( .A(n3629), .B(n3630), .Z(o[1594]) );
  XOR U4029 ( .A(n3633), .B(n3634), .Z(o[1593]) );
  XNOR U4030 ( .A(n3637), .B(n3638), .Z(o[1592]) );
  XNOR U4031 ( .A(n3641), .B(n3642), .Z(o[1591]) );
  XOR U4032 ( .A(n3645), .B(n3646), .Z(o[1590]) );
  XOR U4033 ( .A(n3649), .B(n3356), .Z(o[158]) );
  XOR U4034 ( .A(n1934), .B(round_reg[695]), .Z(n3356) );
  ANDN U4035 ( .A(n1276), .B(n1277), .Z(n3649) );
  XOR U4036 ( .A(n2269), .B(round_reg[220]), .Z(n1277) );
  XNOR U4037 ( .A(n2363), .B(round_reg[629]), .Z(n1276) );
  XNOR U4038 ( .A(n3650), .B(n3651), .Z(o[1589]) );
  XNOR U4039 ( .A(n3654), .B(n3655), .Z(o[1588]) );
  XNOR U4040 ( .A(n3658), .B(n3659), .Z(o[1587]) );
  XNOR U4041 ( .A(n3662), .B(n3663), .Z(o[1586]) );
  XNOR U4042 ( .A(n3666), .B(n3667), .Z(o[1585]) );
  XNOR U4043 ( .A(n3670), .B(n3671), .Z(o[1584]) );
  XNOR U4044 ( .A(n3674), .B(n3675), .Z(o[1583]) );
  XNOR U4045 ( .A(n3678), .B(n3679), .Z(o[1582]) );
  XOR U4046 ( .A(n3682), .B(n3683), .Z(o[1581]) );
  XOR U4047 ( .A(n3686), .B(n3687), .Z(o[1580]) );
  XOR U4048 ( .A(n3690), .B(n3358), .Z(o[157]) );
  XOR U4049 ( .A(n1936), .B(round_reg[694]), .Z(n3358) );
  ANDN U4050 ( .A(n1320), .B(n1321), .Z(n3690) );
  XNOR U4051 ( .A(n2273), .B(round_reg[219]), .Z(n1321) );
  XNOR U4052 ( .A(n2367), .B(round_reg[628]), .Z(n1320) );
  XNOR U4053 ( .A(n3691), .B(n3692), .Z(o[1579]) );
  XNOR U4054 ( .A(n3695), .B(n3696), .Z(o[1578]) );
  AND U4055 ( .A(n3697), .B(n3698), .Z(n3695) );
  XNOR U4056 ( .A(n3699), .B(n3700), .Z(o[1577]) );
  XNOR U4057 ( .A(n3703), .B(n3704), .Z(o[1576]) );
  XNOR U4058 ( .A(n3707), .B(n3708), .Z(o[1575]) );
  XNOR U4059 ( .A(n3711), .B(n3712), .Z(o[1574]) );
  XNOR U4060 ( .A(n3715), .B(n3716), .Z(o[1573]) );
  XNOR U4061 ( .A(n3719), .B(n3720), .Z(o[1572]) );
  XNOR U4062 ( .A(n3723), .B(n3724), .Z(o[1571]) );
  XNOR U4063 ( .A(n3727), .B(n3728), .Z(o[1570]) );
  XOR U4064 ( .A(n3731), .B(n3360), .Z(o[156]) );
  XOR U4065 ( .A(n1938), .B(round_reg[693]), .Z(n3360) );
  ANDN U4066 ( .A(n1364), .B(n1365), .Z(n3731) );
  XNOR U4067 ( .A(n2277), .B(round_reg[218]), .Z(n1365) );
  XNOR U4068 ( .A(n2371), .B(round_reg[627]), .Z(n1364) );
  XNOR U4069 ( .A(n3732), .B(n3733), .Z(o[1569]) );
  XNOR U4070 ( .A(n3736), .B(n3737), .Z(o[1568]) );
  XOR U4071 ( .A(n3740), .B(n3741), .Z(o[1567]) );
  XOR U4072 ( .A(n3742), .B(n3743), .Z(n3740) );
  NAND U4073 ( .A(n3746), .B(n3747), .Z(n3742) );
  AND U4074 ( .A(n3748), .B(n3749), .Z(n3747) );
  ANDN U4075 ( .A(n3750), .B(rc_i[3]), .Z(n3749) );
  NOR U4076 ( .A(rc_i[5]), .B(rc_i[6]), .Z(n3750) );
  NOR U4077 ( .A(rc_i[23]), .B(rc_i[22]), .Z(n3748) );
  AND U4078 ( .A(n3751), .B(n3752), .Z(n3746) );
  AND U4079 ( .A(n3753), .B(n3754), .Z(n3752) );
  NOR U4080 ( .A(rc_i[20]), .B(rc_i[19]), .Z(n3753) );
  NOR U4081 ( .A(rc_i[10]), .B(rc_i[11]), .Z(n3751) );
  XOR U4082 ( .A(n3755), .B(n3756), .Z(o[1566]) );
  XOR U4083 ( .A(n3759), .B(n3760), .Z(o[1565]) );
  XOR U4084 ( .A(n3763), .B(n3764), .Z(o[1564]) );
  XOR U4085 ( .A(n3767), .B(n3768), .Z(o[1563]) );
  XOR U4086 ( .A(n3771), .B(n3772), .Z(o[1562]) );
  XNOR U4087 ( .A(n3775), .B(n3776), .Z(o[1561]) );
  XNOR U4088 ( .A(n3779), .B(n3780), .Z(o[1560]) );
  XOR U4089 ( .A(n3783), .B(n3363), .Z(o[155]) );
  XOR U4090 ( .A(n1940), .B(round_reg[692]), .Z(n3363) );
  ANDN U4091 ( .A(n1408), .B(n1409), .Z(n3783) );
  XNOR U4092 ( .A(n2281), .B(round_reg[217]), .Z(n1409) );
  XNOR U4093 ( .A(n2375), .B(round_reg[626]), .Z(n1408) );
  XNOR U4094 ( .A(n3784), .B(n3785), .Z(o[1559]) );
  XNOR U4095 ( .A(n3788), .B(n3789), .Z(o[1558]) );
  XNOR U4096 ( .A(n3792), .B(n3793), .Z(o[1557]) );
  XNOR U4097 ( .A(n3796), .B(n3797), .Z(o[1556]) );
  XNOR U4098 ( .A(n3800), .B(n3801), .Z(o[1555]) );
  XNOR U4099 ( .A(n3804), .B(n3805), .Z(o[1554]) );
  XNOR U4100 ( .A(n3808), .B(n3809), .Z(o[1553]) );
  XNOR U4101 ( .A(n3812), .B(n3813), .Z(o[1552]) );
  XNOR U4102 ( .A(n3816), .B(n3817), .Z(o[1551]) );
  XOR U4103 ( .A(n3818), .B(n3819), .Z(n3816) );
  NAND U4104 ( .A(n3822), .B(n3823), .Z(n3818) );
  AND U4105 ( .A(n3824), .B(n3825), .Z(n3823) );
  ANDN U4106 ( .A(n3826), .B(rc_i[18]), .Z(n3825) );
  NOR U4107 ( .A(rc_i[3]), .B(rc_i[4]), .Z(n3826) );
  NOR U4108 ( .A(rc_i[16]), .B(n3827), .Z(n3824) );
  AND U4109 ( .A(n3828), .B(n3829), .Z(n3822) );
  ANDN U4110 ( .A(n3611), .B(n3610), .Z(n3829) );
  NANDN U4111 ( .B(rc_i[20]), .A(n3830), .Z(n3610) );
  NOR U4112 ( .A(rc_i[23]), .B(rc_i[21]), .Z(n3830) );
  NOR U4113 ( .A(n3831), .B(n3832), .Z(n3828) );
  XNOR U4114 ( .A(n3833), .B(n3834), .Z(o[1550]) );
  XOR U4115 ( .A(n3837), .B(n3367), .Z(o[154]) );
  XOR U4116 ( .A(n1943), .B(round_reg[691]), .Z(n3367) );
  ANDN U4117 ( .A(n1452), .B(n1453), .Z(n3837) );
  XNOR U4118 ( .A(n2285), .B(round_reg[216]), .Z(n1453) );
  XNOR U4119 ( .A(n2379), .B(round_reg[625]), .Z(n1452) );
  XNOR U4120 ( .A(n3838), .B(n3839), .Z(o[1549]) );
  XNOR U4121 ( .A(n3842), .B(n3843), .Z(o[1548]) );
  AND U4122 ( .A(n3844), .B(n3845), .Z(n3842) );
  IV U4123 ( .A(n3846), .Z(n3845) );
  XNOR U4124 ( .A(n3847), .B(n3848), .Z(o[1547]) );
  XNOR U4125 ( .A(n3851), .B(n3852), .Z(o[1546]) );
  XNOR U4126 ( .A(n3855), .B(n3856), .Z(o[1545]) );
  XNOR U4127 ( .A(n3859), .B(n3860), .Z(o[1544]) );
  XNOR U4128 ( .A(n3863), .B(n3864), .Z(o[1543]) );
  XOR U4129 ( .A(n3865), .B(n3866), .Z(n3863) );
  NAND U4130 ( .A(n3869), .B(n3870), .Z(n3865) );
  AND U4131 ( .A(n3871), .B(n3872), .Z(n3870) );
  ANDN U4132 ( .A(n3873), .B(rc_i[6]), .Z(n3872) );
  ANDN U4133 ( .A(n3874), .B(rc_i[9]), .Z(n3873) );
  NOR U4134 ( .A(rc_i[20]), .B(rc_i[21]), .Z(n3871) );
  AND U4135 ( .A(n3875), .B(n3876), .Z(n3869) );
  ANDN U4136 ( .A(n3877), .B(rc_i[13]), .Z(n3876) );
  NOR U4137 ( .A(rc_i[17]), .B(rc_i[14]), .Z(n3877) );
  ANDN U4138 ( .A(n3754), .B(n3878), .Z(n3875) );
  XNOR U4139 ( .A(n3879), .B(n3880), .Z(o[1542]) );
  XOR U4140 ( .A(n3883), .B(n3884), .Z(o[1541]) );
  XNOR U4141 ( .A(n3887), .B(n3888), .Z(o[1540]) );
  XOR U4142 ( .A(n3891), .B(n3371), .Z(o[153]) );
  XOR U4143 ( .A(n1946), .B(round_reg[690]), .Z(n3371) );
  ANDN U4144 ( .A(n1500), .B(n1501), .Z(n3891) );
  XNOR U4145 ( .A(n2289), .B(round_reg[215]), .Z(n1501) );
  XNOR U4146 ( .A(n2383), .B(round_reg[624]), .Z(n1500) );
  XNOR U4147 ( .A(n3892), .B(n3893), .Z(o[1539]) );
  XOR U4148 ( .A(n3894), .B(n3895), .Z(n3892) );
  NAND U4149 ( .A(n3898), .B(n3899), .Z(n3894) );
  AND U4150 ( .A(n3900), .B(n3901), .Z(n3899) );
  AND U4151 ( .A(n3902), .B(n3903), .Z(n3901) );
  NOR U4152 ( .A(rc_i[8]), .B(rc_i[9]), .Z(n3903) );
  NOR U4153 ( .A(rc_i[4]), .B(rc_i[7]), .Z(n3902) );
  ANDN U4154 ( .A(n3904), .B(rc_i[19]), .Z(n3900) );
  NOR U4155 ( .A(rc_i[23]), .B(rc_i[2]), .Z(n3904) );
  AND U4156 ( .A(n3905), .B(n3906), .Z(n3898) );
  ANDN U4157 ( .A(n3907), .B(rc_i[13]), .Z(n3906) );
  NOR U4158 ( .A(rc_i[18]), .B(rc_i[14]), .Z(n3907) );
  ANDN U4159 ( .A(n3908), .B(rc_i[10]), .Z(n3905) );
  ANDN U4160 ( .A(n3754), .B(rc_i[11]), .Z(n3908) );
  IV U4161 ( .A(rc_i[12]), .Z(n3754) );
  XNOR U4162 ( .A(n3909), .B(n3910), .Z(o[1538]) );
  XNOR U4163 ( .A(n3913), .B(n3914), .Z(o[1537]) );
  XOR U4164 ( .A(n3915), .B(n3916), .Z(n3913) );
  NAND U4165 ( .A(n3919), .B(n3920), .Z(n3915) );
  AND U4166 ( .A(n3921), .B(n3922), .Z(n3920) );
  ANDN U4167 ( .A(n3923), .B(rc_i[18]), .Z(n3922) );
  ANDN U4168 ( .A(n3874), .B(rc_i[19]), .Z(n3923) );
  IV U4169 ( .A(rc_i[8]), .Z(n3874) );
  NOR U4170 ( .A(rc_i[16]), .B(rc_i[15]), .Z(n3921) );
  AND U4171 ( .A(n3924), .B(n3925), .Z(n3919) );
  NOR U4172 ( .A(rc_i[12]), .B(rc_i[13]), .Z(n3925) );
  NOR U4173 ( .A(n3878), .B(rc_i[11]), .Z(n3924) );
  OR U4174 ( .A(n3832), .B(rc_i[4]), .Z(n3878) );
  OR U4175 ( .A(rc_i[1]), .B(rc_i[2]), .Z(n3832) );
  XNOR U4176 ( .A(n3926), .B(n3927), .Z(o[1536]) );
  XOR U4177 ( .A(n3928), .B(n3929), .Z(n3926) );
  NAND U4178 ( .A(n3932), .B(n3933), .Z(n3928) );
  AND U4179 ( .A(n3934), .B(n3935), .Z(n3933) );
  NOR U4180 ( .A(rc_i[5]), .B(rc_i[4]), .Z(n3935) );
  NOR U4181 ( .A(rc_i[20]), .B(rc_i[22]), .Z(n3934) );
  AND U4182 ( .A(n3936), .B(n3937), .Z(n3932) );
  ANDN U4183 ( .A(n3611), .B(rc_i[0]), .Z(n3937) );
  NOR U4184 ( .A(rc_i[7]), .B(rc_i[6]), .Z(n3611) );
  NOR U4185 ( .A(n3831), .B(n3612), .Z(n3936) );
  OR U4186 ( .A(n3827), .B(rc_i[13]), .Z(n3612) );
  OR U4187 ( .A(rc_i[15]), .B(rc_i[14]), .Z(n3827) );
  OR U4188 ( .A(rc_i[10]), .B(rc_i[12]), .Z(n3831) );
  XOR U4189 ( .A(n3938), .B(n3603), .Z(o[1535]) );
  ANDN U4190 ( .A(n3939), .B(n3602), .Z(n3938) );
  XOR U4191 ( .A(n3940), .B(n3616), .Z(o[1534]) );
  ANDN U4192 ( .A(n3941), .B(n3615), .Z(n3940) );
  XOR U4193 ( .A(n3942), .B(n3620), .Z(o[1533]) );
  ANDN U4194 ( .A(n3943), .B(n3619), .Z(n3942) );
  XOR U4195 ( .A(n3944), .B(n3624), .Z(o[1532]) );
  ANDN U4196 ( .A(n3945), .B(n3623), .Z(n3944) );
  XOR U4197 ( .A(n3946), .B(n3628), .Z(o[1531]) );
  ANDN U4198 ( .A(n3947), .B(n3627), .Z(n3946) );
  XOR U4199 ( .A(n3948), .B(n3632), .Z(o[1530]) );
  ANDN U4200 ( .A(n3949), .B(n3631), .Z(n3948) );
  XOR U4201 ( .A(n3950), .B(n3375), .Z(o[152]) );
  XOR U4202 ( .A(n1949), .B(round_reg[689]), .Z(n3375) );
  ANDN U4203 ( .A(n1532), .B(n1533), .Z(n3950) );
  XNOR U4204 ( .A(n2293), .B(round_reg[214]), .Z(n1533) );
  XNOR U4205 ( .A(n2387), .B(round_reg[623]), .Z(n1532) );
  XOR U4206 ( .A(n3951), .B(n3636), .Z(o[1529]) );
  ANDN U4207 ( .A(n3952), .B(n3635), .Z(n3951) );
  XOR U4208 ( .A(n3953), .B(n3640), .Z(o[1528]) );
  ANDN U4209 ( .A(n3954), .B(n3639), .Z(n3953) );
  XOR U4210 ( .A(n3955), .B(n3644), .Z(o[1527]) );
  ANDN U4211 ( .A(n3956), .B(n3643), .Z(n3955) );
  XOR U4212 ( .A(n3957), .B(n3648), .Z(o[1526]) );
  ANDN U4213 ( .A(n3958), .B(n3647), .Z(n3957) );
  XOR U4214 ( .A(n3959), .B(n3653), .Z(o[1525]) );
  ANDN U4215 ( .A(n3960), .B(n3652), .Z(n3959) );
  XOR U4216 ( .A(n3961), .B(n3657), .Z(o[1524]) );
  ANDN U4217 ( .A(n3962), .B(n3656), .Z(n3961) );
  XOR U4218 ( .A(n3963), .B(n3661), .Z(o[1523]) );
  ANDN U4219 ( .A(n3964), .B(n3660), .Z(n3963) );
  XOR U4220 ( .A(n3965), .B(n3665), .Z(o[1522]) );
  ANDN U4221 ( .A(n3966), .B(n3664), .Z(n3965) );
  XOR U4222 ( .A(n3967), .B(n3669), .Z(o[1521]) );
  ANDN U4223 ( .A(n3968), .B(n3668), .Z(n3967) );
  XOR U4224 ( .A(n3969), .B(n3673), .Z(o[1520]) );
  ANDN U4225 ( .A(n3970), .B(n3672), .Z(n3969) );
  XOR U4226 ( .A(n3971), .B(n3380), .Z(o[151]) );
  XOR U4227 ( .A(n1952), .B(round_reg[688]), .Z(n3380) );
  ANDN U4228 ( .A(n1562), .B(n1563), .Z(n3971) );
  XNOR U4229 ( .A(n2297), .B(round_reg[213]), .Z(n1563) );
  XNOR U4230 ( .A(n2391), .B(round_reg[622]), .Z(n1562) );
  XOR U4231 ( .A(n3972), .B(n3677), .Z(o[1519]) );
  ANDN U4232 ( .A(n3973), .B(n3676), .Z(n3972) );
  XOR U4233 ( .A(n3974), .B(n3681), .Z(o[1518]) );
  ANDN U4234 ( .A(n3975), .B(n3680), .Z(n3974) );
  XOR U4235 ( .A(n3976), .B(n3685), .Z(o[1517]) );
  ANDN U4236 ( .A(n3977), .B(n3684), .Z(n3976) );
  XOR U4237 ( .A(n3978), .B(n3689), .Z(o[1516]) );
  ANDN U4238 ( .A(n3979), .B(n3688), .Z(n3978) );
  XOR U4239 ( .A(n3980), .B(n3694), .Z(o[1515]) );
  ANDN U4240 ( .A(n3981), .B(n3693), .Z(n3980) );
  XNOR U4241 ( .A(n3982), .B(n3698), .Z(o[1514]) );
  ANDN U4242 ( .A(n3983), .B(n3697), .Z(n3982) );
  XOR U4243 ( .A(n3984), .B(n3702), .Z(o[1513]) );
  ANDN U4244 ( .A(n3985), .B(n3701), .Z(n3984) );
  XOR U4245 ( .A(n3986), .B(n3706), .Z(o[1512]) );
  ANDN U4246 ( .A(n3987), .B(n3705), .Z(n3986) );
  XOR U4247 ( .A(n3988), .B(n3710), .Z(o[1511]) );
  ANDN U4248 ( .A(n3989), .B(n3709), .Z(n3988) );
  XOR U4249 ( .A(n3990), .B(n3714), .Z(o[1510]) );
  ANDN U4250 ( .A(n3991), .B(n3713), .Z(n3990) );
  XOR U4251 ( .A(n3992), .B(n3384), .Z(o[150]) );
  XOR U4252 ( .A(n1959), .B(round_reg[687]), .Z(n3384) );
  ANDN U4253 ( .A(n1587), .B(n1588), .Z(n3992) );
  XNOR U4254 ( .A(n2301), .B(round_reg[212]), .Z(n1588) );
  XNOR U4255 ( .A(n2112), .B(round_reg[621]), .Z(n1587) );
  IV U4256 ( .A(n3993), .Z(n2112) );
  XOR U4257 ( .A(n3994), .B(n3718), .Z(o[1509]) );
  ANDN U4258 ( .A(n3995), .B(n3717), .Z(n3994) );
  XOR U4259 ( .A(n3996), .B(n3722), .Z(o[1508]) );
  AND U4260 ( .A(n3997), .B(n3998), .Z(n3996) );
  IV U4261 ( .A(n3721), .Z(n3998) );
  XOR U4262 ( .A(n3999), .B(n3726), .Z(o[1507]) );
  AND U4263 ( .A(n4000), .B(n4001), .Z(n3999) );
  IV U4264 ( .A(n3725), .Z(n4001) );
  XOR U4265 ( .A(n4002), .B(n3730), .Z(o[1506]) );
  AND U4266 ( .A(n4003), .B(n4004), .Z(n4002) );
  IV U4267 ( .A(n3729), .Z(n4004) );
  XOR U4268 ( .A(n4005), .B(n3735), .Z(o[1505]) );
  AND U4269 ( .A(n4006), .B(n4007), .Z(n4005) );
  IV U4270 ( .A(n3734), .Z(n4007) );
  XOR U4271 ( .A(n4008), .B(n3739), .Z(o[1504]) );
  XOR U4272 ( .A(n4010), .B(n3745), .Z(o[1503]) );
  ANDN U4273 ( .A(n4011), .B(n3744), .Z(n4010) );
  XOR U4274 ( .A(n4012), .B(n3758), .Z(o[1502]) );
  ANDN U4275 ( .A(n4013), .B(n3757), .Z(n4012) );
  XOR U4276 ( .A(n4014), .B(n3762), .Z(o[1501]) );
  ANDN U4277 ( .A(n4015), .B(n3761), .Z(n4014) );
  XOR U4278 ( .A(n4016), .B(n3766), .Z(o[1500]) );
  ANDN U4279 ( .A(n4017), .B(n3765), .Z(n4016) );
  XNOR U4280 ( .A(n4018), .B(n1857), .Z(o[14]) );
  ANDN U4281 ( .A(n3415), .B(n3416), .Z(n4018) );
  XOR U4282 ( .A(n1763), .B(round_reg[1047]), .Z(n3416) );
  XNOR U4283 ( .A(n2296), .B(round_reg[1424]), .Z(n3415) );
  XOR U4284 ( .A(n4019), .B(n3388), .Z(o[149]) );
  XOR U4285 ( .A(n1962), .B(round_reg[686]), .Z(n3388) );
  ANDN U4286 ( .A(n1620), .B(n1621), .Z(n4019) );
  XNOR U4287 ( .A(n2305), .B(round_reg[211]), .Z(n1621) );
  XNOR U4288 ( .A(n2116), .B(round_reg[620]), .Z(n1620) );
  IV U4289 ( .A(n4020), .Z(n2116) );
  XOR U4290 ( .A(n4021), .B(n3770), .Z(o[1499]) );
  ANDN U4291 ( .A(n4022), .B(n3769), .Z(n4021) );
  XOR U4292 ( .A(n4023), .B(n3774), .Z(o[1498]) );
  ANDN U4293 ( .A(n4024), .B(n3773), .Z(n4023) );
  XOR U4294 ( .A(n4025), .B(n3778), .Z(o[1497]) );
  ANDN U4295 ( .A(n4026), .B(n3777), .Z(n4025) );
  XOR U4296 ( .A(n4027), .B(n3782), .Z(o[1496]) );
  ANDN U4297 ( .A(n4028), .B(n3781), .Z(n4027) );
  XOR U4298 ( .A(n4029), .B(n3787), .Z(o[1495]) );
  ANDN U4299 ( .A(n4030), .B(n3786), .Z(n4029) );
  XOR U4300 ( .A(n4031), .B(n3791), .Z(o[1494]) );
  ANDN U4301 ( .A(n4032), .B(n3790), .Z(n4031) );
  XOR U4302 ( .A(n4033), .B(n3795), .Z(o[1493]) );
  ANDN U4303 ( .A(n4034), .B(n3794), .Z(n4033) );
  XOR U4304 ( .A(n4035), .B(n3799), .Z(o[1492]) );
  ANDN U4305 ( .A(n4036), .B(n3798), .Z(n4035) );
  XOR U4306 ( .A(n4037), .B(n3803), .Z(o[1491]) );
  ANDN U4307 ( .A(n4038), .B(n3802), .Z(n4037) );
  XOR U4308 ( .A(n4039), .B(n3807), .Z(o[1490]) );
  ANDN U4309 ( .A(n4040), .B(n3806), .Z(n4039) );
  XOR U4310 ( .A(n4041), .B(n3392), .Z(o[148]) );
  XOR U4311 ( .A(n1965), .B(round_reg[685]), .Z(n3392) );
  ANDN U4312 ( .A(n1654), .B(n1655), .Z(n4041) );
  XNOR U4313 ( .A(n2313), .B(round_reg[210]), .Z(n1655) );
  XNOR U4314 ( .A(n2120), .B(round_reg[619]), .Z(n1654) );
  XOR U4315 ( .A(n4042), .B(n3811), .Z(o[1489]) );
  ANDN U4316 ( .A(n4043), .B(n3810), .Z(n4042) );
  XOR U4317 ( .A(n4044), .B(n3815), .Z(o[1488]) );
  ANDN U4318 ( .A(n4045), .B(n3814), .Z(n4044) );
  XOR U4319 ( .A(n4046), .B(n3821), .Z(o[1487]) );
  ANDN U4320 ( .A(n4047), .B(n3820), .Z(n4046) );
  XOR U4321 ( .A(n4048), .B(n3836), .Z(o[1486]) );
  ANDN U4322 ( .A(n4049), .B(n3835), .Z(n4048) );
  XOR U4323 ( .A(n4050), .B(n3841), .Z(o[1485]) );
  ANDN U4324 ( .A(n4051), .B(n3840), .Z(n4050) );
  XOR U4325 ( .A(n4052), .B(n3846), .Z(o[1484]) );
  ANDN U4326 ( .A(n4053), .B(n3844), .Z(n4052) );
  XOR U4327 ( .A(n4054), .B(n3850), .Z(o[1483]) );
  ANDN U4328 ( .A(n4055), .B(n3849), .Z(n4054) );
  XOR U4329 ( .A(n4056), .B(n3854), .Z(o[1482]) );
  ANDN U4330 ( .A(n4057), .B(n3853), .Z(n4056) );
  XOR U4331 ( .A(n4058), .B(n3858), .Z(o[1481]) );
  ANDN U4332 ( .A(n4059), .B(n3857), .Z(n4058) );
  XOR U4333 ( .A(n4060), .B(n3862), .Z(o[1480]) );
  ANDN U4334 ( .A(n4061), .B(n3861), .Z(n4060) );
  XOR U4335 ( .A(n4062), .B(n3396), .Z(o[147]) );
  XOR U4336 ( .A(n1968), .B(round_reg[684]), .Z(n3396) );
  ANDN U4337 ( .A(n1688), .B(n1689), .Z(n4062) );
  XNOR U4338 ( .A(n2317), .B(round_reg[209]), .Z(n1689) );
  XNOR U4339 ( .A(n2124), .B(round_reg[618]), .Z(n1688) );
  XOR U4340 ( .A(n4063), .B(n3868), .Z(o[1479]) );
  ANDN U4341 ( .A(n4064), .B(n3867), .Z(n4063) );
  XOR U4342 ( .A(n4065), .B(n3882), .Z(o[1478]) );
  ANDN U4343 ( .A(n4066), .B(n3881), .Z(n4065) );
  XOR U4344 ( .A(n4067), .B(n3886), .Z(o[1477]) );
  ANDN U4345 ( .A(n4068), .B(n3885), .Z(n4067) );
  XOR U4346 ( .A(n4069), .B(n3890), .Z(o[1476]) );
  ANDN U4347 ( .A(n4070), .B(n3889), .Z(n4069) );
  XOR U4348 ( .A(n4071), .B(n3897), .Z(o[1475]) );
  ANDN U4349 ( .A(n4072), .B(n3896), .Z(n4071) );
  XOR U4350 ( .A(n4073), .B(n3912), .Z(o[1474]) );
  ANDN U4351 ( .A(n4074), .B(n3911), .Z(n4073) );
  XOR U4352 ( .A(n4075), .B(n3918), .Z(o[1473]) );
  ANDN U4353 ( .A(n4076), .B(n3917), .Z(n4075) );
  XOR U4354 ( .A(n4077), .B(n3931), .Z(o[1472]) );
  ANDN U4355 ( .A(n4078), .B(n3930), .Z(n4077) );
  XOR U4356 ( .A(n4079), .B(n3602), .Z(o[1471]) );
  XOR U4357 ( .A(n2280), .B(round_reg[788]), .Z(n3602) );
  ANDN U4358 ( .A(n4080), .B(n3939), .Z(n4079) );
  XOR U4359 ( .A(n4081), .B(n3615), .Z(o[1470]) );
  XOR U4360 ( .A(n2284), .B(round_reg[787]), .Z(n3615) );
  ANDN U4361 ( .A(n4082), .B(n3941), .Z(n4081) );
  XOR U4362 ( .A(n4083), .B(n3401), .Z(o[146]) );
  IV U4363 ( .A(n3536), .Z(n3401) );
  XNOR U4364 ( .A(n1971), .B(round_reg[683]), .Z(n3536) );
  ANDN U4365 ( .A(n1716), .B(n1717), .Z(n4083) );
  XNOR U4366 ( .A(n2321), .B(round_reg[208]), .Z(n1717) );
  XNOR U4367 ( .A(n2135), .B(round_reg[617]), .Z(n1716) );
  XOR U4368 ( .A(n4084), .B(n3619), .Z(o[1469]) );
  XOR U4369 ( .A(n2288), .B(round_reg[786]), .Z(n3619) );
  ANDN U4370 ( .A(n4085), .B(n3943), .Z(n4084) );
  XOR U4371 ( .A(n4086), .B(n3623), .Z(o[1468]) );
  XOR U4372 ( .A(n2292), .B(round_reg[785]), .Z(n3623) );
  ANDN U4373 ( .A(n4087), .B(n3945), .Z(n4086) );
  XOR U4374 ( .A(n4088), .B(n3627), .Z(o[1467]) );
  XOR U4375 ( .A(n2296), .B(round_reg[784]), .Z(n3627) );
  ANDN U4376 ( .A(n4089), .B(n3947), .Z(n4088) );
  XOR U4377 ( .A(n4090), .B(n3631), .Z(o[1466]) );
  XOR U4378 ( .A(n2300), .B(round_reg[783]), .Z(n3631) );
  ANDN U4379 ( .A(n4091), .B(n3949), .Z(n4090) );
  XOR U4380 ( .A(n4092), .B(n3635), .Z(o[1465]) );
  XOR U4381 ( .A(n2304), .B(round_reg[782]), .Z(n3635) );
  ANDN U4382 ( .A(n4093), .B(n3952), .Z(n4092) );
  XOR U4383 ( .A(n4094), .B(n3639), .Z(o[1464]) );
  XOR U4384 ( .A(n2312), .B(round_reg[781]), .Z(n3639) );
  ANDN U4385 ( .A(n4095), .B(n3954), .Z(n4094) );
  XOR U4386 ( .A(n4096), .B(n3643), .Z(o[1463]) );
  XOR U4387 ( .A(n2316), .B(round_reg[780]), .Z(n3643) );
  ANDN U4388 ( .A(n4097), .B(n3956), .Z(n4096) );
  XOR U4389 ( .A(n4098), .B(n3647), .Z(o[1462]) );
  XOR U4390 ( .A(n2320), .B(round_reg[779]), .Z(n3647) );
  ANDN U4391 ( .A(n4099), .B(n3958), .Z(n4098) );
  XOR U4392 ( .A(n4100), .B(n3652), .Z(o[1461]) );
  XOR U4393 ( .A(n2324), .B(round_reg[778]), .Z(n3652) );
  ANDN U4394 ( .A(n4101), .B(n3960), .Z(n4100) );
  XOR U4395 ( .A(n4102), .B(n3656), .Z(o[1460]) );
  XOR U4396 ( .A(n2328), .B(round_reg[777]), .Z(n3656) );
  ANDN U4397 ( .A(n4103), .B(n3962), .Z(n4102) );
  XOR U4398 ( .A(n4104), .B(n3405), .Z(o[145]) );
  IV U4399 ( .A(n3539), .Z(n3405) );
  XNOR U4400 ( .A(n1974), .B(round_reg[682]), .Z(n3539) );
  ANDN U4401 ( .A(n1750), .B(n1751), .Z(n4104) );
  XNOR U4402 ( .A(n2325), .B(round_reg[207]), .Z(n1751) );
  XNOR U4403 ( .A(n2139), .B(round_reg[616]), .Z(n1750) );
  XOR U4404 ( .A(n4105), .B(n3660), .Z(o[1459]) );
  XOR U4405 ( .A(n2332), .B(round_reg[776]), .Z(n3660) );
  ANDN U4406 ( .A(n4106), .B(n3964), .Z(n4105) );
  XOR U4407 ( .A(n4107), .B(n3664), .Z(o[1458]) );
  XOR U4408 ( .A(n2336), .B(round_reg[775]), .Z(n3664) );
  ANDN U4409 ( .A(n4108), .B(n3966), .Z(n4107) );
  XOR U4410 ( .A(n4109), .B(n3668), .Z(o[1457]) );
  XOR U4411 ( .A(n2340), .B(round_reg[774]), .Z(n3668) );
  ANDN U4412 ( .A(n4110), .B(n3968), .Z(n4109) );
  XOR U4413 ( .A(n4111), .B(n3672), .Z(o[1456]) );
  XOR U4414 ( .A(n2344), .B(round_reg[773]), .Z(n3672) );
  ANDN U4415 ( .A(n4112), .B(n3970), .Z(n4111) );
  XOR U4416 ( .A(n4113), .B(n3676), .Z(o[1455]) );
  XOR U4417 ( .A(n2348), .B(round_reg[772]), .Z(n3676) );
  ANDN U4418 ( .A(n4114), .B(n3973), .Z(n4113) );
  XOR U4419 ( .A(n4115), .B(n3680), .Z(o[1454]) );
  XOR U4420 ( .A(n2356), .B(round_reg[771]), .Z(n3680) );
  ANDN U4421 ( .A(n4116), .B(n3975), .Z(n4115) );
  XOR U4422 ( .A(n4117), .B(n3684), .Z(o[1453]) );
  XOR U4423 ( .A(n2360), .B(round_reg[770]), .Z(n3684) );
  ANDN U4424 ( .A(n4118), .B(n3977), .Z(n4117) );
  XOR U4425 ( .A(n4119), .B(n3688), .Z(o[1452]) );
  XOR U4426 ( .A(n2364), .B(round_reg[769]), .Z(n3688) );
  ANDN U4427 ( .A(n4120), .B(n3979), .Z(n4119) );
  XOR U4428 ( .A(n4121), .B(n3693), .Z(o[1451]) );
  XOR U4429 ( .A(n2368), .B(round_reg[768]), .Z(n3693) );
  ANDN U4430 ( .A(n4122), .B(n3981), .Z(n4121) );
  XOR U4431 ( .A(n4123), .B(n3697), .Z(o[1450]) );
  XOR U4432 ( .A(n2372), .B(round_reg[831]), .Z(n3697) );
  ANDN U4433 ( .A(n4124), .B(n3983), .Z(n4123) );
  XOR U4434 ( .A(n4125), .B(n3409), .Z(o[144]) );
  XOR U4435 ( .A(n1977), .B(round_reg[681]), .Z(n3409) );
  ANDN U4436 ( .A(n1784), .B(n1785), .Z(n4125) );
  XNOR U4437 ( .A(n2329), .B(round_reg[206]), .Z(n1785) );
  XNOR U4438 ( .A(n2143), .B(round_reg[615]), .Z(n1784) );
  XOR U4439 ( .A(n4126), .B(n3701), .Z(o[1449]) );
  XOR U4440 ( .A(n2376), .B(round_reg[830]), .Z(n3701) );
  ANDN U4441 ( .A(n4127), .B(n3985), .Z(n4126) );
  XOR U4442 ( .A(n4128), .B(n3705), .Z(o[1448]) );
  XOR U4443 ( .A(n2380), .B(round_reg[829]), .Z(n3705) );
  ANDN U4444 ( .A(n4129), .B(n3987), .Z(n4128) );
  XOR U4445 ( .A(n4130), .B(n3709), .Z(o[1447]) );
  XOR U4446 ( .A(n2384), .B(round_reg[828]), .Z(n3709) );
  ANDN U4447 ( .A(n4131), .B(n3989), .Z(n4130) );
  XOR U4448 ( .A(n4132), .B(n3713), .Z(o[1446]) );
  XOR U4449 ( .A(n2388), .B(round_reg[827]), .Z(n3713) );
  XOR U4450 ( .A(n4134), .B(n3717), .Z(o[1445]) );
  XOR U4451 ( .A(n2392), .B(round_reg[826]), .Z(n3717) );
  AND U4452 ( .A(n4135), .B(n4136), .Z(n4134) );
  IV U4453 ( .A(n3995), .Z(n4136) );
  XOR U4454 ( .A(n4137), .B(n3721), .Z(o[1444]) );
  XOR U4455 ( .A(n2114), .B(round_reg[825]), .Z(n3721) );
  AND U4456 ( .A(n4138), .B(n4139), .Z(n4137) );
  IV U4457 ( .A(n3997), .Z(n4139) );
  XOR U4458 ( .A(n4140), .B(n3725), .Z(o[1443]) );
  XOR U4459 ( .A(n2118), .B(round_reg[824]), .Z(n3725) );
  AND U4460 ( .A(n4141), .B(n4142), .Z(n4140) );
  IV U4461 ( .A(n4000), .Z(n4142) );
  XOR U4462 ( .A(n4143), .B(n3729), .Z(o[1442]) );
  XOR U4463 ( .A(n2122), .B(round_reg[823]), .Z(n3729) );
  AND U4464 ( .A(n4144), .B(n4145), .Z(n4143) );
  IV U4465 ( .A(n4003), .Z(n4145) );
  XOR U4466 ( .A(n4146), .B(n3734), .Z(o[1441]) );
  XOR U4467 ( .A(n2126), .B(round_reg[822]), .Z(n3734) );
  AND U4468 ( .A(n4147), .B(n4148), .Z(n4146) );
  IV U4469 ( .A(n4006), .Z(n4148) );
  XOR U4470 ( .A(n4149), .B(n3738), .Z(o[1440]) );
  XOR U4471 ( .A(n2137), .B(round_reg[821]), .Z(n3738) );
  ANDN U4472 ( .A(n4150), .B(n4009), .Z(n4149) );
  XOR U4473 ( .A(n4151), .B(n3413), .Z(o[143]) );
  XOR U4474 ( .A(n1979), .B(round_reg[680]), .Z(n3413) );
  ANDN U4475 ( .A(n1822), .B(n1823), .Z(n4151) );
  XNOR U4476 ( .A(n2333), .B(round_reg[205]), .Z(n1823) );
  XNOR U4477 ( .A(n2147), .B(round_reg[614]), .Z(n1822) );
  XOR U4478 ( .A(n4152), .B(n3744), .Z(o[1439]) );
  XOR U4479 ( .A(n2140), .B(round_reg[820]), .Z(n3744) );
  ANDN U4480 ( .A(n4153), .B(n4011), .Z(n4152) );
  XOR U4481 ( .A(n4154), .B(n3757), .Z(o[1438]) );
  XOR U4482 ( .A(n2144), .B(round_reg[819]), .Z(n3757) );
  ANDN U4483 ( .A(n4155), .B(n4013), .Z(n4154) );
  XOR U4484 ( .A(n4156), .B(n3761), .Z(o[1437]) );
  XOR U4485 ( .A(n2148), .B(round_reg[818]), .Z(n3761) );
  ANDN U4486 ( .A(n4157), .B(n4015), .Z(n4156) );
  XOR U4487 ( .A(n4158), .B(n3765), .Z(o[1436]) );
  XOR U4488 ( .A(n2152), .B(round_reg[817]), .Z(n3765) );
  ANDN U4489 ( .A(n4159), .B(n4017), .Z(n4158) );
  XOR U4490 ( .A(n4160), .B(n3769), .Z(o[1435]) );
  XOR U4491 ( .A(n2156), .B(round_reg[816]), .Z(n3769) );
  ANDN U4492 ( .A(n4161), .B(n4022), .Z(n4160) );
  XOR U4493 ( .A(n4162), .B(n3773), .Z(o[1434]) );
  XOR U4494 ( .A(n2160), .B(round_reg[815]), .Z(n3773) );
  ANDN U4495 ( .A(n4163), .B(n4024), .Z(n4162) );
  XOR U4496 ( .A(n4164), .B(n3777), .Z(o[1433]) );
  XOR U4497 ( .A(n2164), .B(round_reg[814]), .Z(n3777) );
  ANDN U4498 ( .A(n4165), .B(n4026), .Z(n4164) );
  XOR U4499 ( .A(n4166), .B(n3781), .Z(o[1432]) );
  XOR U4500 ( .A(n2168), .B(round_reg[813]), .Z(n3781) );
  ANDN U4501 ( .A(n4167), .B(n4028), .Z(n4166) );
  XOR U4502 ( .A(n4168), .B(n3786), .Z(o[1431]) );
  XNOR U4503 ( .A(n2172), .B(round_reg[812]), .Z(n3786) );
  ANDN U4504 ( .A(n4169), .B(n4030), .Z(n4168) );
  XOR U4505 ( .A(n4170), .B(n3790), .Z(o[1430]) );
  XNOR U4506 ( .A(n2180), .B(round_reg[811]), .Z(n3790) );
  ANDN U4507 ( .A(n4171), .B(n4032), .Z(n4170) );
  XOR U4508 ( .A(n4172), .B(n3417), .Z(o[142]) );
  XOR U4509 ( .A(n1981), .B(round_reg[679]), .Z(n3417) );
  ANDN U4510 ( .A(n1856), .B(n1857), .Z(n4172) );
  XNOR U4511 ( .A(n2337), .B(round_reg[204]), .Z(n1857) );
  XNOR U4512 ( .A(n2151), .B(round_reg[613]), .Z(n1856) );
  XOR U4513 ( .A(n4173), .B(n3794), .Z(o[1429]) );
  XOR U4514 ( .A(n2184), .B(round_reg[810]), .Z(n3794) );
  ANDN U4515 ( .A(n4174), .B(n4034), .Z(n4173) );
  XOR U4516 ( .A(n4175), .B(n3798), .Z(o[1428]) );
  XOR U4517 ( .A(n2188), .B(round_reg[809]), .Z(n3798) );
  ANDN U4518 ( .A(n4176), .B(n4036), .Z(n4175) );
  XOR U4519 ( .A(n4177), .B(n3802), .Z(o[1427]) );
  XOR U4520 ( .A(n2192), .B(round_reg[808]), .Z(n3802) );
  ANDN U4521 ( .A(n4178), .B(n4038), .Z(n4177) );
  XOR U4522 ( .A(n4179), .B(n3806), .Z(o[1426]) );
  XOR U4523 ( .A(n2196), .B(round_reg[807]), .Z(n3806) );
  ANDN U4524 ( .A(n4180), .B(n4040), .Z(n4179) );
  XOR U4525 ( .A(n4181), .B(n3810), .Z(o[1425]) );
  XOR U4526 ( .A(n2200), .B(round_reg[806]), .Z(n3810) );
  ANDN U4527 ( .A(n4182), .B(n4043), .Z(n4181) );
  XOR U4528 ( .A(n4183), .B(n3814), .Z(o[1424]) );
  XOR U4529 ( .A(n2204), .B(round_reg[805]), .Z(n3814) );
  ANDN U4530 ( .A(n4184), .B(n4045), .Z(n4183) );
  XOR U4531 ( .A(n4185), .B(n3820), .Z(o[1423]) );
  XOR U4532 ( .A(n2208), .B(round_reg[804]), .Z(n3820) );
  ANDN U4533 ( .A(n4186), .B(n4047), .Z(n4185) );
  XOR U4534 ( .A(n4187), .B(n3835), .Z(o[1422]) );
  XNOR U4535 ( .A(n2212), .B(round_reg[803]), .Z(n3835) );
  ANDN U4536 ( .A(n4188), .B(n4049), .Z(n4187) );
  XOR U4537 ( .A(n4189), .B(n3840), .Z(o[1421]) );
  XOR U4538 ( .A(n2216), .B(round_reg[802]), .Z(n3840) );
  ANDN U4539 ( .A(n4190), .B(n4051), .Z(n4189) );
  XOR U4540 ( .A(n4191), .B(n3844), .Z(o[1420]) );
  XOR U4541 ( .A(n2224), .B(round_reg[801]), .Z(n3844) );
  ANDN U4542 ( .A(n4192), .B(n4053), .Z(n4191) );
  XOR U4543 ( .A(n4193), .B(n3421), .Z(o[141]) );
  XOR U4544 ( .A(n1983), .B(round_reg[678]), .Z(n3421) );
  AND U4545 ( .A(n1892), .B(n1890), .Z(n4193) );
  XNOR U4546 ( .A(n2155), .B(round_reg[612]), .Z(n1890) );
  XOR U4547 ( .A(n4194), .B(n3849), .Z(o[1419]) );
  XOR U4548 ( .A(n2228), .B(round_reg[800]), .Z(n3849) );
  ANDN U4549 ( .A(n4195), .B(n4055), .Z(n4194) );
  XOR U4550 ( .A(n4196), .B(n3853), .Z(o[1418]) );
  XOR U4551 ( .A(n2232), .B(round_reg[799]), .Z(n3853) );
  ANDN U4552 ( .A(n4197), .B(n4057), .Z(n4196) );
  XOR U4553 ( .A(n4198), .B(n3857), .Z(o[1417]) );
  XOR U4554 ( .A(n2236), .B(round_reg[798]), .Z(n3857) );
  ANDN U4555 ( .A(n4199), .B(n4059), .Z(n4198) );
  XOR U4556 ( .A(n4200), .B(n3861), .Z(o[1416]) );
  XOR U4557 ( .A(n2240), .B(round_reg[797]), .Z(n3861) );
  ANDN U4558 ( .A(n4201), .B(n4061), .Z(n4200) );
  XOR U4559 ( .A(n4202), .B(n3867), .Z(o[1415]) );
  XOR U4560 ( .A(n2244), .B(round_reg[796]), .Z(n3867) );
  ANDN U4561 ( .A(n4203), .B(n4064), .Z(n4202) );
  XOR U4562 ( .A(n4204), .B(n3881), .Z(o[1414]) );
  XOR U4563 ( .A(n2248), .B(round_reg[795]), .Z(n3881) );
  ANDN U4564 ( .A(n4205), .B(n4066), .Z(n4204) );
  XOR U4565 ( .A(n4206), .B(n3885), .Z(o[1413]) );
  XOR U4566 ( .A(n2252), .B(round_reg[794]), .Z(n3885) );
  ANDN U4567 ( .A(n4207), .B(n4068), .Z(n4206) );
  XOR U4568 ( .A(n4208), .B(n3889), .Z(o[1412]) );
  XOR U4569 ( .A(n2256), .B(round_reg[793]), .Z(n3889) );
  ANDN U4570 ( .A(n4209), .B(n4070), .Z(n4208) );
  XOR U4571 ( .A(n4210), .B(n3896), .Z(o[1411]) );
  XOR U4572 ( .A(n2260), .B(round_reg[792]), .Z(n3896) );
  ANDN U4573 ( .A(n4211), .B(n4072), .Z(n4210) );
  XOR U4574 ( .A(n4212), .B(n3911), .Z(o[1410]) );
  XOR U4575 ( .A(n2268), .B(round_reg[791]), .Z(n3911) );
  ANDN U4576 ( .A(n4213), .B(n4074), .Z(n4212) );
  XOR U4577 ( .A(n4214), .B(n3424), .Z(o[140]) );
  XOR U4578 ( .A(n1989), .B(round_reg[677]), .Z(n3424) );
  AND U4579 ( .A(n1926), .B(n1924), .Z(n4214) );
  XNOR U4580 ( .A(n2159), .B(round_reg[611]), .Z(n1924) );
  XOR U4581 ( .A(n4215), .B(n3917), .Z(o[1409]) );
  XOR U4582 ( .A(n2272), .B(round_reg[790]), .Z(n3917) );
  ANDN U4583 ( .A(n4216), .B(n4076), .Z(n4215) );
  XOR U4584 ( .A(n4217), .B(n3930), .Z(o[1408]) );
  XOR U4585 ( .A(n2276), .B(round_reg[789]), .Z(n3930) );
  ANDN U4586 ( .A(n4218), .B(n4078), .Z(n4217) );
  XOR U4587 ( .A(n4219), .B(n3939), .Z(o[1407]) );
  XNOR U4588 ( .A(n1918), .B(round_reg[426]), .Z(n3939) );
  NOR U4589 ( .A(n4080), .B(n3599), .Z(n4219) );
  XOR U4590 ( .A(n4220), .B(n3941), .Z(o[1406]) );
  XNOR U4591 ( .A(n1921), .B(round_reg[425]), .Z(n3941) );
  NOR U4592 ( .A(n4082), .B(n3614), .Z(n4220) );
  XOR U4593 ( .A(n4221), .B(n3943), .Z(o[1405]) );
  XNOR U4594 ( .A(n1928), .B(round_reg[424]), .Z(n3943) );
  NOR U4595 ( .A(n4085), .B(n3618), .Z(n4221) );
  XOR U4596 ( .A(n4222), .B(n3945), .Z(o[1404]) );
  XNOR U4597 ( .A(n1931), .B(round_reg[423]), .Z(n3945) );
  NOR U4598 ( .A(n4087), .B(n3622), .Z(n4222) );
  XOR U4599 ( .A(n4223), .B(n3947), .Z(o[1403]) );
  XNOR U4600 ( .A(n1710), .B(round_reg[422]), .Z(n3947) );
  NOR U4601 ( .A(n4089), .B(n3626), .Z(n4223) );
  XOR U4602 ( .A(n4224), .B(n3949), .Z(o[1402]) );
  XNOR U4603 ( .A(n1713), .B(round_reg[421]), .Z(n3949) );
  ANDN U4604 ( .A(n3630), .B(n4091), .Z(n4224) );
  XOR U4605 ( .A(n4225), .B(n3952), .Z(o[1401]) );
  XNOR U4606 ( .A(n1720), .B(round_reg[420]), .Z(n3952) );
  ANDN U4607 ( .A(n3634), .B(n4093), .Z(n4225) );
  XOR U4608 ( .A(n4226), .B(n3954), .Z(o[1400]) );
  XNOR U4609 ( .A(n1723), .B(round_reg[419]), .Z(n3954) );
  NOR U4610 ( .A(n4095), .B(n3638), .Z(n4226) );
  XOR U4611 ( .A(n4227), .B(n1892), .Z(o[13]) );
  XOR U4612 ( .A(n2341), .B(round_reg[203]), .Z(n1892) );
  ANDN U4613 ( .A(n1891), .B(n3420), .Z(n4227) );
  XOR U4614 ( .A(n1766), .B(round_reg[1046]), .Z(n3420) );
  XNOR U4615 ( .A(n2300), .B(round_reg[1423]), .Z(n1891) );
  XOR U4616 ( .A(n4228), .B(n3427), .Z(o[139]) );
  XOR U4617 ( .A(n1991), .B(round_reg[676]), .Z(n3427) );
  AND U4618 ( .A(n1957), .B(n1955), .Z(n4228) );
  XNOR U4619 ( .A(n2163), .B(round_reg[610]), .Z(n1955) );
  XOR U4620 ( .A(n4229), .B(n3956), .Z(o[1399]) );
  XNOR U4621 ( .A(n1726), .B(round_reg[418]), .Z(n3956) );
  XOR U4622 ( .A(n4230), .B(n3958), .Z(o[1398]) );
  XNOR U4623 ( .A(n1729), .B(round_reg[417]), .Z(n3958) );
  XOR U4624 ( .A(n4231), .B(n3960), .Z(o[1397]) );
  XOR U4625 ( .A(n1732), .B(round_reg[416]), .Z(n3960) );
  XOR U4626 ( .A(n4232), .B(n3962), .Z(o[1396]) );
  XOR U4627 ( .A(n1735), .B(round_reg[415]), .Z(n3962) );
  XOR U4628 ( .A(n4233), .B(n3964), .Z(o[1395]) );
  XOR U4629 ( .A(n1738), .B(round_reg[414]), .Z(n3964) );
  XOR U4630 ( .A(n4234), .B(n3966), .Z(o[1394]) );
  XOR U4631 ( .A(n1741), .B(round_reg[413]), .Z(n3966) );
  XOR U4632 ( .A(n4235), .B(n3968), .Z(o[1393]) );
  XOR U4633 ( .A(n1744), .B(round_reg[412]), .Z(n3968) );
  XOR U4634 ( .A(n4236), .B(n3970), .Z(o[1392]) );
  XOR U4635 ( .A(n1747), .B(round_reg[411]), .Z(n3970) );
  XOR U4636 ( .A(n4237), .B(n3973), .Z(o[1391]) );
  XNOR U4637 ( .A(n1754), .B(round_reg[410]), .Z(n3973) );
  NOR U4638 ( .A(n4114), .B(n3675), .Z(n4237) );
  XOR U4639 ( .A(n4238), .B(n3975), .Z(o[1390]) );
  XNOR U4640 ( .A(n1757), .B(round_reg[409]), .Z(n3975) );
  NOR U4641 ( .A(n4116), .B(n3679), .Z(n4238) );
  XOR U4642 ( .A(n4239), .B(n3430), .Z(o[138]) );
  XOR U4643 ( .A(n1993), .B(round_reg[675]), .Z(n3430) );
  AND U4644 ( .A(n1987), .B(n1985), .Z(n4239) );
  XNOR U4645 ( .A(n2167), .B(round_reg[609]), .Z(n1985) );
  XOR U4646 ( .A(n4240), .B(n3977), .Z(o[1389]) );
  XNOR U4647 ( .A(n1760), .B(round_reg[408]), .Z(n3977) );
  ANDN U4648 ( .A(n3683), .B(n4118), .Z(n4240) );
  XOR U4649 ( .A(n4241), .B(n3979), .Z(o[1388]) );
  XNOR U4650 ( .A(n1763), .B(round_reg[407]), .Z(n3979) );
  ANDN U4651 ( .A(n3687), .B(n4120), .Z(n4241) );
  XOR U4652 ( .A(n4242), .B(n3981), .Z(o[1387]) );
  XNOR U4653 ( .A(n1766), .B(round_reg[406]), .Z(n3981) );
  NOR U4654 ( .A(n4122), .B(n3692), .Z(n4242) );
  XOR U4655 ( .A(n4243), .B(n3983), .Z(o[1386]) );
  XNOR U4656 ( .A(n1769), .B(round_reg[405]), .Z(n3983) );
  XOR U4657 ( .A(n4244), .B(n3985), .Z(o[1385]) );
  XNOR U4658 ( .A(n1772), .B(round_reg[404]), .Z(n3985) );
  XOR U4659 ( .A(n4245), .B(n3987), .Z(o[1384]) );
  XNOR U4660 ( .A(n1775), .B(round_reg[403]), .Z(n3987) );
  XOR U4661 ( .A(n4246), .B(n3989), .Z(o[1383]) );
  XOR U4662 ( .A(n1778), .B(round_reg[402]), .Z(n3989) );
  XOR U4663 ( .A(n4247), .B(n3991), .Z(o[1382]) );
  XOR U4664 ( .A(n1781), .B(round_reg[401]), .Z(n3991) );
  IV U4665 ( .A(n4248), .Z(n1781) );
  XOR U4666 ( .A(n4249), .B(n3995), .Z(o[1381]) );
  XOR U4667 ( .A(n1788), .B(round_reg[400]), .Z(n3995) );
  IV U4668 ( .A(n4250), .Z(n1788) );
  XOR U4669 ( .A(n4251), .B(n3997), .Z(o[1380]) );
  XOR U4670 ( .A(n1791), .B(round_reg[399]), .Z(n3997) );
  IV U4671 ( .A(n4252), .Z(n1791) );
  ANDN U4672 ( .A(n4253), .B(n3720), .Z(n4251) );
  IV U4673 ( .A(n4138), .Z(n4253) );
  XOR U4674 ( .A(n4254), .B(n3548), .Z(o[137]) );
  XOR U4675 ( .A(n1995), .B(round_reg[674]), .Z(n3548) );
  AND U4676 ( .A(n2009), .B(n1052), .Z(n4254) );
  IV U4677 ( .A(n2010), .Z(n1052) );
  XNOR U4678 ( .A(n2361), .B(round_reg[199]), .Z(n2010) );
  XNOR U4679 ( .A(n2171), .B(round_reg[608]), .Z(n2009) );
  XOR U4680 ( .A(n4255), .B(n4000), .Z(o[1379]) );
  XOR U4681 ( .A(n1794), .B(round_reg[398]), .Z(n4000) );
  IV U4682 ( .A(n4256), .Z(n1794) );
  ANDN U4683 ( .A(n4257), .B(n3724), .Z(n4255) );
  IV U4684 ( .A(n4141), .Z(n4257) );
  XOR U4685 ( .A(n4258), .B(n4003), .Z(o[1378]) );
  XOR U4686 ( .A(n1797), .B(round_reg[397]), .Z(n4003) );
  IV U4687 ( .A(n4259), .Z(n1797) );
  ANDN U4688 ( .A(n4260), .B(n3728), .Z(n4258) );
  IV U4689 ( .A(n4144), .Z(n4260) );
  XOR U4690 ( .A(n4261), .B(n4006), .Z(o[1377]) );
  XOR U4691 ( .A(n1800), .B(round_reg[396]), .Z(n4006) );
  IV U4692 ( .A(n4262), .Z(n1800) );
  NOR U4693 ( .A(n4147), .B(n3733), .Z(n4261) );
  XOR U4694 ( .A(n4263), .B(n4009), .Z(o[1376]) );
  XOR U4695 ( .A(n1803), .B(round_reg[395]), .Z(n4009) );
  NOR U4696 ( .A(n3737), .B(n4150), .Z(n4263) );
  XOR U4697 ( .A(n4264), .B(n4011), .Z(o[1375]) );
  XOR U4698 ( .A(n1806), .B(round_reg[394]), .Z(n4011) );
  ANDN U4699 ( .A(n3741), .B(n4153), .Z(n4264) );
  XOR U4700 ( .A(n4265), .B(n4013), .Z(o[1374]) );
  XOR U4701 ( .A(n1809), .B(round_reg[393]), .Z(n4013) );
  ANDN U4702 ( .A(n3756), .B(n4155), .Z(n4265) );
  XOR U4703 ( .A(n4266), .B(n4015), .Z(o[1373]) );
  XOR U4704 ( .A(n1812), .B(round_reg[392]), .Z(n4015) );
  ANDN U4705 ( .A(n3760), .B(n4157), .Z(n4266) );
  XOR U4706 ( .A(n4267), .B(n4017), .Z(o[1372]) );
  XOR U4707 ( .A(n1815), .B(round_reg[391]), .Z(n4017) );
  ANDN U4708 ( .A(n3764), .B(n4159), .Z(n4267) );
  XOR U4709 ( .A(n4268), .B(n4022), .Z(o[1371]) );
  XOR U4710 ( .A(n1826), .B(round_reg[390]), .Z(n4022) );
  ANDN U4711 ( .A(n3768), .B(n4161), .Z(n4268) );
  XOR U4712 ( .A(n4269), .B(n4024), .Z(o[1370]) );
  XOR U4713 ( .A(n1829), .B(round_reg[389]), .Z(n4024) );
  ANDN U4714 ( .A(n3772), .B(n4163), .Z(n4269) );
  XOR U4715 ( .A(n4270), .B(n3434), .Z(o[136]) );
  XOR U4716 ( .A(n1997), .B(round_reg[673]), .Z(n3434) );
  IV U4717 ( .A(n4271), .Z(n1997) );
  ANDN U4718 ( .A(n2034), .B(n1496), .Z(n4270) );
  XNOR U4719 ( .A(n2365), .B(round_reg[198]), .Z(n1496) );
  XNOR U4720 ( .A(n2179), .B(round_reg[607]), .Z(n2034) );
  XOR U4721 ( .A(n4272), .B(n4026), .Z(o[1369]) );
  XOR U4722 ( .A(n1832), .B(round_reg[388]), .Z(n4026) );
  NOR U4723 ( .A(n4165), .B(n3776), .Z(n4272) );
  XOR U4724 ( .A(n4273), .B(n4028), .Z(o[1368]) );
  XOR U4725 ( .A(n1835), .B(round_reg[387]), .Z(n4028) );
  NOR U4726 ( .A(n4167), .B(n3780), .Z(n4273) );
  XOR U4727 ( .A(n4274), .B(n4030), .Z(o[1367]) );
  XOR U4728 ( .A(n1838), .B(round_reg[386]), .Z(n4030) );
  NOR U4729 ( .A(n4169), .B(n3785), .Z(n4274) );
  XOR U4730 ( .A(n4275), .B(n4032), .Z(o[1366]) );
  XOR U4731 ( .A(n1841), .B(round_reg[385]), .Z(n4032) );
  NOR U4732 ( .A(n4171), .B(n3789), .Z(n4275) );
  XOR U4733 ( .A(n4276), .B(n4034), .Z(o[1365]) );
  XOR U4734 ( .A(n1844), .B(round_reg[384]), .Z(n4034) );
  NOR U4735 ( .A(n4174), .B(n3793), .Z(n4276) );
  XOR U4736 ( .A(n4277), .B(n4036), .Z(o[1364]) );
  XOR U4737 ( .A(n1847), .B(round_reg[447]), .Z(n4036) );
  NOR U4738 ( .A(n4176), .B(n3797), .Z(n4277) );
  XOR U4739 ( .A(n4278), .B(n4038), .Z(o[1363]) );
  XOR U4740 ( .A(n1850), .B(round_reg[446]), .Z(n4038) );
  NOR U4741 ( .A(n4178), .B(n3801), .Z(n4278) );
  XOR U4742 ( .A(n4279), .B(n4040), .Z(o[1362]) );
  XOR U4743 ( .A(n1853), .B(round_reg[445]), .Z(n4040) );
  NOR U4744 ( .A(n4180), .B(n3805), .Z(n4279) );
  XOR U4745 ( .A(n4280), .B(n4043), .Z(o[1361]) );
  XOR U4746 ( .A(n1860), .B(round_reg[444]), .Z(n4043) );
  NOR U4747 ( .A(n4182), .B(n3809), .Z(n4280) );
  XOR U4748 ( .A(n4281), .B(n4045), .Z(o[1360]) );
  XOR U4749 ( .A(n1863), .B(round_reg[443]), .Z(n4045) );
  NOR U4750 ( .A(n4184), .B(n3813), .Z(n4281) );
  XOR U4751 ( .A(n4282), .B(n3437), .Z(o[135]) );
  XOR U4752 ( .A(n1999), .B(round_reg[672]), .Z(n3437) );
  IV U4753 ( .A(n4283), .Z(n1999) );
  ANDN U4754 ( .A(n2065), .B(n1818), .Z(n4282) );
  XNOR U4755 ( .A(n2369), .B(round_reg[197]), .Z(n1818) );
  XNOR U4756 ( .A(n2183), .B(round_reg[606]), .Z(n2065) );
  XOR U4757 ( .A(n4284), .B(n4047), .Z(o[1359]) );
  XOR U4758 ( .A(n1866), .B(round_reg[442]), .Z(n4047) );
  NOR U4759 ( .A(n4186), .B(n3817), .Z(n4284) );
  XOR U4760 ( .A(n4285), .B(n4049), .Z(o[1358]) );
  XOR U4761 ( .A(n1869), .B(round_reg[441]), .Z(n4049) );
  NOR U4762 ( .A(n4188), .B(n3834), .Z(n4285) );
  XOR U4763 ( .A(n4286), .B(n4051), .Z(o[1357]) );
  XOR U4764 ( .A(n1872), .B(round_reg[440]), .Z(n4051) );
  NOR U4765 ( .A(n4190), .B(n3839), .Z(n4286) );
  XOR U4766 ( .A(n4287), .B(n4053), .Z(o[1356]) );
  XOR U4767 ( .A(n1875), .B(round_reg[439]), .Z(n4053) );
  NOR U4768 ( .A(n4192), .B(n3843), .Z(n4287) );
  XOR U4769 ( .A(n4288), .B(n4055), .Z(o[1355]) );
  XOR U4770 ( .A(n1878), .B(round_reg[438]), .Z(n4055) );
  NOR U4771 ( .A(n4195), .B(n3848), .Z(n4288) );
  XOR U4772 ( .A(n4289), .B(n4057), .Z(o[1354]) );
  XOR U4773 ( .A(n1881), .B(round_reg[437]), .Z(n4057) );
  NOR U4774 ( .A(n4197), .B(n3852), .Z(n4289) );
  XOR U4775 ( .A(n4290), .B(n4059), .Z(o[1353]) );
  XOR U4776 ( .A(n1884), .B(round_reg[436]), .Z(n4059) );
  NOR U4777 ( .A(n4199), .B(n3856), .Z(n4290) );
  XOR U4778 ( .A(n4291), .B(n4061), .Z(o[1352]) );
  XOR U4779 ( .A(n1887), .B(round_reg[435]), .Z(n4061) );
  NOR U4780 ( .A(n4201), .B(n3860), .Z(n4291) );
  XOR U4781 ( .A(n4292), .B(n4064), .Z(o[1351]) );
  XOR U4782 ( .A(n1894), .B(round_reg[434]), .Z(n4064) );
  NOR U4783 ( .A(n4203), .B(n3864), .Z(n4292) );
  XOR U4784 ( .A(n4293), .B(n4066), .Z(o[1350]) );
  XOR U4785 ( .A(n1897), .B(round_reg[433]), .Z(n4066) );
  NOR U4786 ( .A(n4205), .B(n3880), .Z(n4293) );
  XOR U4787 ( .A(n4294), .B(n3440), .Z(o[134]) );
  XOR U4788 ( .A(n2001), .B(round_reg[671]), .Z(n3440) );
  IV U4789 ( .A(n4295), .Z(n2001) );
  ANDN U4790 ( .A(n2091), .B(n2092), .Z(n4294) );
  XNOR U4791 ( .A(n2373), .B(round_reg[196]), .Z(n2092) );
  XNOR U4792 ( .A(n2187), .B(round_reg[605]), .Z(n2091) );
  XOR U4793 ( .A(n4296), .B(n4068), .Z(o[1349]) );
  XOR U4794 ( .A(n1900), .B(round_reg[432]), .Z(n4068) );
  ANDN U4795 ( .A(n3884), .B(n4207), .Z(n4296) );
  XOR U4796 ( .A(n4297), .B(n4070), .Z(o[1348]) );
  XOR U4797 ( .A(n1903), .B(round_reg[431]), .Z(n4070) );
  NOR U4798 ( .A(n4209), .B(n3888), .Z(n4297) );
  XOR U4799 ( .A(n4298), .B(n4072), .Z(o[1347]) );
  XOR U4800 ( .A(n1906), .B(round_reg[430]), .Z(n4072) );
  NOR U4801 ( .A(n4211), .B(n3893), .Z(n4298) );
  XOR U4802 ( .A(n4299), .B(n4074), .Z(o[1346]) );
  XOR U4803 ( .A(n1909), .B(round_reg[429]), .Z(n4074) );
  NOR U4804 ( .A(n4213), .B(n3910), .Z(n4299) );
  XOR U4805 ( .A(n4300), .B(n4076), .Z(o[1345]) );
  XNOR U4806 ( .A(n1912), .B(round_reg[428]), .Z(n4076) );
  NOR U4807 ( .A(n4216), .B(n3914), .Z(n4300) );
  XOR U4808 ( .A(n4301), .B(n4078), .Z(o[1344]) );
  XNOR U4809 ( .A(n1915), .B(round_reg[427]), .Z(n4078) );
  NOR U4810 ( .A(n4218), .B(n3927), .Z(n4301) );
  XOR U4811 ( .A(n4302), .B(n4080), .Z(o[1343]) );
  XOR U4812 ( .A(n1949), .B(round_reg[49]), .Z(n4080) );
  AND U4813 ( .A(n3599), .B(n3603), .Z(n4302) );
  XOR U4814 ( .A(n2305), .B(round_reg[1171]), .Z(n3603) );
  XNOR U4815 ( .A(n2319), .B(round_reg[1599]), .Z(n3599) );
  XOR U4816 ( .A(n4303), .B(n4082), .Z(o[1342]) );
  XOR U4817 ( .A(n1952), .B(round_reg[48]), .Z(n4082) );
  AND U4818 ( .A(n3614), .B(n3616), .Z(n4303) );
  XOR U4819 ( .A(n2313), .B(round_reg[1170]), .Z(n3616) );
  XNOR U4820 ( .A(n2323), .B(round_reg[1598]), .Z(n3614) );
  XOR U4821 ( .A(n4304), .B(n4085), .Z(o[1341]) );
  XOR U4822 ( .A(n1959), .B(round_reg[47]), .Z(n4085) );
  AND U4823 ( .A(n3618), .B(n3620), .Z(n4304) );
  XOR U4824 ( .A(n2317), .B(round_reg[1169]), .Z(n3620) );
  XNOR U4825 ( .A(n2327), .B(round_reg[1597]), .Z(n3618) );
  XOR U4826 ( .A(n4305), .B(n4087), .Z(o[1340]) );
  XOR U4827 ( .A(n1962), .B(round_reg[46]), .Z(n4087) );
  AND U4828 ( .A(n3622), .B(n3624), .Z(n4305) );
  XOR U4829 ( .A(n2321), .B(round_reg[1168]), .Z(n3624) );
  XNOR U4830 ( .A(n2331), .B(round_reg[1596]), .Z(n3622) );
  XOR U4831 ( .A(n4306), .B(n3442), .Z(o[133]) );
  XOR U4832 ( .A(n2003), .B(round_reg[670]), .Z(n3442) );
  IV U4833 ( .A(n4307), .Z(n2003) );
  ANDN U4834 ( .A(n2131), .B(n2132), .Z(n4306) );
  XNOR U4835 ( .A(n2377), .B(round_reg[195]), .Z(n2132) );
  XNOR U4836 ( .A(n2191), .B(round_reg[604]), .Z(n2131) );
  XOR U4837 ( .A(n4308), .B(n4089), .Z(o[1339]) );
  XOR U4838 ( .A(n1965), .B(round_reg[45]), .Z(n4089) );
  AND U4839 ( .A(n3626), .B(n3628), .Z(n4308) );
  XOR U4840 ( .A(n2325), .B(round_reg[1167]), .Z(n3628) );
  XNOR U4841 ( .A(n2335), .B(round_reg[1595]), .Z(n3626) );
  XOR U4842 ( .A(n4309), .B(n4091), .Z(o[1338]) );
  XOR U4843 ( .A(n1968), .B(round_reg[44]), .Z(n4091) );
  ANDN U4844 ( .A(n3632), .B(n3630), .Z(n4309) );
  XOR U4845 ( .A(n2339), .B(round_reg[1594]), .Z(n3630) );
  XOR U4846 ( .A(n2329), .B(round_reg[1166]), .Z(n3632) );
  XOR U4847 ( .A(n4310), .B(n4093), .Z(o[1337]) );
  XOR U4848 ( .A(n1971), .B(round_reg[43]), .Z(n4093) );
  ANDN U4849 ( .A(n3636), .B(n3634), .Z(n4310) );
  XOR U4850 ( .A(n2343), .B(round_reg[1593]), .Z(n3634) );
  XOR U4851 ( .A(n2333), .B(round_reg[1165]), .Z(n3636) );
  XOR U4852 ( .A(n4311), .B(n4095), .Z(o[1336]) );
  XOR U4853 ( .A(n1974), .B(round_reg[42]), .Z(n4095) );
  AND U4854 ( .A(n3638), .B(n3640), .Z(n4311) );
  XOR U4855 ( .A(n2337), .B(round_reg[1164]), .Z(n3640) );
  XNOR U4856 ( .A(n2347), .B(round_reg[1592]), .Z(n3638) );
  XOR U4857 ( .A(n4312), .B(n4097), .Z(o[1335]) );
  XOR U4858 ( .A(n1977), .B(round_reg[41]), .Z(n4097) );
  IV U4859 ( .A(n4313), .Z(n1977) );
  AND U4860 ( .A(n3642), .B(n3644), .Z(n4312) );
  XOR U4861 ( .A(n2341), .B(round_reg[1163]), .Z(n3644) );
  XNOR U4862 ( .A(n2355), .B(round_reg[1591]), .Z(n3642) );
  XOR U4863 ( .A(n4314), .B(n4099), .Z(o[1334]) );
  XOR U4864 ( .A(n1979), .B(round_reg[40]), .Z(n4099) );
  IV U4865 ( .A(n4315), .Z(n1979) );
  ANDN U4866 ( .A(n3648), .B(n3646), .Z(n4314) );
  XOR U4867 ( .A(n2359), .B(round_reg[1590]), .Z(n3646) );
  XOR U4868 ( .A(n2345), .B(round_reg[1162]), .Z(n3648) );
  XOR U4869 ( .A(n4316), .B(n4101), .Z(o[1333]) );
  XOR U4870 ( .A(n1981), .B(round_reg[39]), .Z(n4101) );
  IV U4871 ( .A(n4317), .Z(n1981) );
  AND U4872 ( .A(n3651), .B(n3653), .Z(n4316) );
  XOR U4873 ( .A(n2349), .B(round_reg[1161]), .Z(n3653) );
  XNOR U4874 ( .A(n2363), .B(round_reg[1589]), .Z(n3651) );
  IV U4875 ( .A(n4318), .Z(n2363) );
  XOR U4876 ( .A(n4319), .B(n4103), .Z(o[1332]) );
  XOR U4877 ( .A(n1983), .B(round_reg[38]), .Z(n4103) );
  IV U4878 ( .A(n4320), .Z(n1983) );
  AND U4879 ( .A(n3655), .B(n3657), .Z(n4319) );
  XOR U4880 ( .A(n2357), .B(round_reg[1160]), .Z(n3657) );
  XNOR U4881 ( .A(n2367), .B(round_reg[1588]), .Z(n3655) );
  IV U4882 ( .A(n4321), .Z(n2367) );
  XOR U4883 ( .A(n4322), .B(n4106), .Z(o[1331]) );
  XOR U4884 ( .A(n1989), .B(round_reg[37]), .Z(n4106) );
  IV U4885 ( .A(n4323), .Z(n1989) );
  AND U4886 ( .A(n3659), .B(n3661), .Z(n4322) );
  XOR U4887 ( .A(n2361), .B(round_reg[1159]), .Z(n3661) );
  XNOR U4888 ( .A(n2371), .B(round_reg[1587]), .Z(n3659) );
  IV U4889 ( .A(n4324), .Z(n2371) );
  XOR U4890 ( .A(n4325), .B(n4108), .Z(o[1330]) );
  XOR U4891 ( .A(n1991), .B(round_reg[36]), .Z(n4108) );
  IV U4892 ( .A(n4326), .Z(n1991) );
  AND U4893 ( .A(n3663), .B(n3665), .Z(n4325) );
  XOR U4894 ( .A(n2365), .B(round_reg[1158]), .Z(n3665) );
  XNOR U4895 ( .A(n2375), .B(round_reg[1586]), .Z(n3663) );
  IV U4896 ( .A(n4327), .Z(n2375) );
  XOR U4897 ( .A(n4328), .B(n3444), .Z(o[132]) );
  XOR U4898 ( .A(n2005), .B(round_reg[669]), .Z(n3444) );
  IV U4899 ( .A(n4329), .Z(n2005) );
  ANDN U4900 ( .A(n2175), .B(n2176), .Z(n4328) );
  XNOR U4901 ( .A(n2381), .B(round_reg[194]), .Z(n2176) );
  XNOR U4902 ( .A(n2195), .B(round_reg[603]), .Z(n2175) );
  XOR U4903 ( .A(n4330), .B(n4110), .Z(o[1329]) );
  XOR U4904 ( .A(n1993), .B(round_reg[35]), .Z(n4110) );
  IV U4905 ( .A(n4331), .Z(n1993) );
  AND U4906 ( .A(n3667), .B(n3669), .Z(n4330) );
  XOR U4907 ( .A(n2369), .B(round_reg[1157]), .Z(n3669) );
  XNOR U4908 ( .A(n2379), .B(round_reg[1585]), .Z(n3667) );
  IV U4909 ( .A(n4332), .Z(n2379) );
  XOR U4910 ( .A(n4333), .B(n4112), .Z(o[1328]) );
  XOR U4911 ( .A(n1995), .B(round_reg[34]), .Z(n4112) );
  IV U4912 ( .A(n4334), .Z(n1995) );
  AND U4913 ( .A(n3671), .B(n3673), .Z(n4333) );
  XOR U4914 ( .A(n2373), .B(round_reg[1156]), .Z(n3673) );
  XNOR U4915 ( .A(n2383), .B(round_reg[1584]), .Z(n3671) );
  IV U4916 ( .A(n4335), .Z(n2383) );
  XOR U4917 ( .A(n4336), .B(n4114), .Z(o[1327]) );
  XNOR U4918 ( .A(n4271), .B(round_reg[33]), .Z(n4114) );
  AND U4919 ( .A(n3675), .B(n3677), .Z(n4336) );
  XOR U4920 ( .A(n2377), .B(round_reg[1155]), .Z(n3677) );
  XNOR U4921 ( .A(n2387), .B(round_reg[1583]), .Z(n3675) );
  IV U4922 ( .A(n4337), .Z(n2387) );
  XOR U4923 ( .A(n4338), .B(n4116), .Z(o[1326]) );
  XNOR U4924 ( .A(n4283), .B(round_reg[32]), .Z(n4116) );
  AND U4925 ( .A(n3679), .B(n3681), .Z(n4338) );
  XOR U4926 ( .A(n2381), .B(round_reg[1154]), .Z(n3681) );
  XNOR U4927 ( .A(n2391), .B(round_reg[1582]), .Z(n3679) );
  IV U4928 ( .A(n4339), .Z(n2391) );
  XOR U4929 ( .A(n4340), .B(n4118), .Z(o[1325]) );
  XNOR U4930 ( .A(n4295), .B(round_reg[31]), .Z(n4118) );
  ANDN U4931 ( .A(n3685), .B(n3683), .Z(n4340) );
  XNOR U4932 ( .A(n3993), .B(round_reg[1581]), .Z(n3683) );
  XOR U4933 ( .A(n2385), .B(round_reg[1153]), .Z(n3685) );
  XOR U4934 ( .A(n4341), .B(n4120), .Z(o[1324]) );
  XNOR U4935 ( .A(n4307), .B(round_reg[30]), .Z(n4120) );
  ANDN U4936 ( .A(n3689), .B(n3687), .Z(n4341) );
  XNOR U4937 ( .A(n4020), .B(round_reg[1580]), .Z(n3687) );
  XOR U4938 ( .A(n2389), .B(round_reg[1152]), .Z(n3689) );
  XOR U4939 ( .A(n4342), .B(n4122), .Z(o[1323]) );
  XNOR U4940 ( .A(n4329), .B(round_reg[29]), .Z(n4122) );
  AND U4941 ( .A(n3692), .B(n3694), .Z(n4342) );
  XOR U4942 ( .A(n2393), .B(round_reg[1215]), .Z(n3694) );
  XNOR U4943 ( .A(n2120), .B(round_reg[1579]), .Z(n3692) );
  IV U4944 ( .A(n4343), .Z(n2120) );
  XOR U4945 ( .A(n4344), .B(n4124), .Z(o[1322]) );
  XOR U4946 ( .A(n2007), .B(round_reg[28]), .Z(n4124) );
  ANDN U4947 ( .A(n3696), .B(n3698), .Z(n4344) );
  XNOR U4948 ( .A(n3029), .B(round_reg[1214]), .Z(n3698) );
  XNOR U4949 ( .A(n2124), .B(round_reg[1578]), .Z(n3696) );
  IV U4950 ( .A(n4345), .Z(n2124) );
  XOR U4951 ( .A(n4346), .B(n4127), .Z(o[1321]) );
  XOR U4952 ( .A(n2012), .B(round_reg[27]), .Z(n4127) );
  AND U4953 ( .A(n3700), .B(n3702), .Z(n4346) );
  XOR U4954 ( .A(n2117), .B(round_reg[1213]), .Z(n3702) );
  XNOR U4955 ( .A(n2135), .B(round_reg[1577]), .Z(n3700) );
  IV U4956 ( .A(n4347), .Z(n2135) );
  XOR U4957 ( .A(n4348), .B(n4129), .Z(o[1320]) );
  XOR U4958 ( .A(n2014), .B(round_reg[26]), .Z(n4129) );
  AND U4959 ( .A(n3704), .B(n3706), .Z(n4348) );
  XOR U4960 ( .A(n2121), .B(round_reg[1212]), .Z(n3706) );
  XNOR U4961 ( .A(n2139), .B(round_reg[1576]), .Z(n3704) );
  IV U4962 ( .A(n4349), .Z(n2139) );
  XOR U4963 ( .A(n4350), .B(n3447), .Z(o[131]) );
  XOR U4964 ( .A(n2007), .B(round_reg[668]), .Z(n3447) );
  IV U4965 ( .A(n4351), .Z(n2007) );
  ANDN U4966 ( .A(n2219), .B(n2220), .Z(n4350) );
  XNOR U4967 ( .A(n2385), .B(round_reg[193]), .Z(n2220) );
  XNOR U4968 ( .A(n2199), .B(round_reg[602]), .Z(n2219) );
  XOR U4969 ( .A(n4352), .B(n4131), .Z(o[1319]) );
  XOR U4970 ( .A(n2016), .B(round_reg[25]), .Z(n4131) );
  AND U4971 ( .A(n3708), .B(n3710), .Z(n4352) );
  XOR U4972 ( .A(n2125), .B(round_reg[1211]), .Z(n3710) );
  XNOR U4973 ( .A(n2143), .B(round_reg[1575]), .Z(n3708) );
  IV U4974 ( .A(n4353), .Z(n2143) );
  XOR U4975 ( .A(n4354), .B(n4133), .Z(o[1318]) );
  XOR U4976 ( .A(n2018), .B(round_reg[24]), .Z(n4133) );
  IV U4977 ( .A(n4355), .Z(n2018) );
  AND U4978 ( .A(n3712), .B(n3714), .Z(n4354) );
  XOR U4979 ( .A(n2136), .B(round_reg[1210]), .Z(n3714) );
  XNOR U4980 ( .A(n2147), .B(round_reg[1574]), .Z(n3712) );
  IV U4981 ( .A(n4356), .Z(n2147) );
  XOR U4982 ( .A(n4357), .B(n4135), .Z(o[1317]) );
  XOR U4983 ( .A(n2020), .B(round_reg[23]), .Z(n4135) );
  IV U4984 ( .A(n4358), .Z(n2020) );
  AND U4985 ( .A(n3716), .B(n3718), .Z(n4357) );
  XOR U4986 ( .A(n2141), .B(round_reg[1209]), .Z(n3718) );
  XNOR U4987 ( .A(n2151), .B(round_reg[1573]), .Z(n3716) );
  IV U4988 ( .A(n4359), .Z(n2151) );
  XOR U4989 ( .A(n4360), .B(n4138), .Z(o[1316]) );
  XOR U4990 ( .A(n2022), .B(round_reg[22]), .Z(n4138) );
  IV U4991 ( .A(n4361), .Z(n2022) );
  AND U4992 ( .A(n3720), .B(n3722), .Z(n4360) );
  XOR U4993 ( .A(n2145), .B(round_reg[1208]), .Z(n3722) );
  XNOR U4994 ( .A(n2155), .B(round_reg[1572]), .Z(n3720) );
  IV U4995 ( .A(n4362), .Z(n2155) );
  XOR U4996 ( .A(n4363), .B(n4141), .Z(o[1315]) );
  XOR U4997 ( .A(n2024), .B(round_reg[21]), .Z(n4141) );
  IV U4998 ( .A(n4364), .Z(n2024) );
  AND U4999 ( .A(n3724), .B(n3726), .Z(n4363) );
  XOR U5000 ( .A(n2149), .B(round_reg[1207]), .Z(n3726) );
  XNOR U5001 ( .A(n2159), .B(round_reg[1571]), .Z(n3724) );
  IV U5002 ( .A(n4365), .Z(n2159) );
  XOR U5003 ( .A(n4366), .B(n4144), .Z(o[1314]) );
  XOR U5004 ( .A(n2026), .B(round_reg[20]), .Z(n4144) );
  IV U5005 ( .A(n4367), .Z(n2026) );
  AND U5006 ( .A(n3728), .B(n3730), .Z(n4366) );
  XOR U5007 ( .A(n2153), .B(round_reg[1206]), .Z(n3730) );
  XNOR U5008 ( .A(n2163), .B(round_reg[1570]), .Z(n3728) );
  IV U5009 ( .A(n4368), .Z(n2163) );
  XOR U5010 ( .A(n4369), .B(n4147), .Z(o[1313]) );
  XOR U5011 ( .A(n2028), .B(round_reg[19]), .Z(n4147) );
  AND U5012 ( .A(n3733), .B(n3735), .Z(n4369) );
  XOR U5013 ( .A(n2157), .B(round_reg[1205]), .Z(n3735) );
  XNOR U5014 ( .A(n2167), .B(round_reg[1569]), .Z(n3733) );
  IV U5015 ( .A(n4370), .Z(n2167) );
  XOR U5016 ( .A(n4371), .B(n4150), .Z(o[1312]) );
  XOR U5017 ( .A(n2031), .B(round_reg[18]), .Z(n4150) );
  AND U5018 ( .A(n3737), .B(n3739), .Z(n4371) );
  XOR U5019 ( .A(n2161), .B(round_reg[1204]), .Z(n3739) );
  XNOR U5020 ( .A(n2171), .B(round_reg[1568]), .Z(n3737) );
  IV U5021 ( .A(n4372), .Z(n2171) );
  XOR U5022 ( .A(n4373), .B(n4153), .Z(o[1311]) );
  XOR U5023 ( .A(n2036), .B(round_reg[17]), .Z(n4153) );
  ANDN U5024 ( .A(n3745), .B(n3741), .Z(n4373) );
  XOR U5025 ( .A(n2179), .B(round_reg[1567]), .Z(n3741) );
  XOR U5026 ( .A(n2165), .B(round_reg[1203]), .Z(n3745) );
  XOR U5027 ( .A(n4374), .B(n4155), .Z(o[1310]) );
  XOR U5028 ( .A(n2039), .B(round_reg[16]), .Z(n4155) );
  ANDN U5029 ( .A(n3758), .B(n3756), .Z(n4374) );
  XOR U5030 ( .A(n2183), .B(round_reg[1566]), .Z(n3756) );
  XOR U5031 ( .A(n2169), .B(round_reg[1202]), .Z(n3758) );
  XOR U5032 ( .A(n4375), .B(n3449), .Z(o[130]) );
  XOR U5033 ( .A(n2012), .B(round_reg[667]), .Z(n3449) );
  IV U5034 ( .A(n4376), .Z(n2012) );
  ANDN U5035 ( .A(n2263), .B(n2264), .Z(n4375) );
  XNOR U5036 ( .A(n2389), .B(round_reg[192]), .Z(n2264) );
  XNOR U5037 ( .A(n2203), .B(round_reg[601]), .Z(n2263) );
  XOR U5038 ( .A(n4377), .B(n4157), .Z(o[1309]) );
  XOR U5039 ( .A(n2042), .B(round_reg[15]), .Z(n4157) );
  ANDN U5040 ( .A(n3762), .B(n3760), .Z(n4377) );
  XOR U5041 ( .A(n2187), .B(round_reg[1565]), .Z(n3760) );
  XOR U5042 ( .A(n2173), .B(round_reg[1201]), .Z(n3762) );
  XOR U5043 ( .A(n4378), .B(n4159), .Z(o[1308]) );
  XOR U5044 ( .A(n2044), .B(round_reg[14]), .Z(n4159) );
  ANDN U5045 ( .A(n3766), .B(n3764), .Z(n4378) );
  XOR U5046 ( .A(n2191), .B(round_reg[1564]), .Z(n3764) );
  XOR U5047 ( .A(n2181), .B(round_reg[1200]), .Z(n3766) );
  XOR U5048 ( .A(n4379), .B(n4161), .Z(o[1307]) );
  XOR U5049 ( .A(n2047), .B(round_reg[13]), .Z(n4161) );
  ANDN U5050 ( .A(n3770), .B(n3768), .Z(n4379) );
  XOR U5051 ( .A(n2195), .B(round_reg[1563]), .Z(n3768) );
  XOR U5052 ( .A(n2185), .B(round_reg[1199]), .Z(n3770) );
  XOR U5053 ( .A(n4380), .B(n4163), .Z(o[1306]) );
  XOR U5054 ( .A(n2050), .B(round_reg[12]), .Z(n4163) );
  ANDN U5055 ( .A(n3774), .B(n3772), .Z(n4380) );
  XOR U5056 ( .A(n2199), .B(round_reg[1562]), .Z(n3772) );
  XOR U5057 ( .A(n2189), .B(round_reg[1198]), .Z(n3774) );
  XOR U5058 ( .A(n4381), .B(n4165), .Z(o[1305]) );
  XOR U5059 ( .A(n2053), .B(round_reg[11]), .Z(n4165) );
  AND U5060 ( .A(n3776), .B(n3778), .Z(n4381) );
  XOR U5061 ( .A(n2193), .B(round_reg[1197]), .Z(n3778) );
  XNOR U5062 ( .A(n2203), .B(round_reg[1561]), .Z(n3776) );
  IV U5063 ( .A(n4382), .Z(n2203) );
  XOR U5064 ( .A(n4383), .B(n4167), .Z(o[1304]) );
  XOR U5065 ( .A(n2056), .B(round_reg[10]), .Z(n4167) );
  AND U5066 ( .A(n3780), .B(n3782), .Z(n4383) );
  XOR U5067 ( .A(n2197), .B(round_reg[1196]), .Z(n3782) );
  XNOR U5068 ( .A(n2207), .B(round_reg[1560]), .Z(n3780) );
  XOR U5069 ( .A(n4384), .B(n4169), .Z(o[1303]) );
  XOR U5070 ( .A(n2059), .B(round_reg[9]), .Z(n4169) );
  AND U5071 ( .A(n3785), .B(n3787), .Z(n4384) );
  XOR U5072 ( .A(n2201), .B(round_reg[1195]), .Z(n3787) );
  XNOR U5073 ( .A(n2211), .B(round_reg[1559]), .Z(n3785) );
  XOR U5074 ( .A(n4385), .B(n4171), .Z(o[1302]) );
  XOR U5075 ( .A(n2062), .B(round_reg[8]), .Z(n4171) );
  AND U5076 ( .A(n3789), .B(n3791), .Z(n4385) );
  XOR U5077 ( .A(n2205), .B(round_reg[1194]), .Z(n3791) );
  XNOR U5078 ( .A(n2215), .B(round_reg[1558]), .Z(n3789) );
  XOR U5079 ( .A(n4386), .B(n4174), .Z(o[1301]) );
  XOR U5080 ( .A(n2067), .B(round_reg[7]), .Z(n4174) );
  AND U5081 ( .A(n3793), .B(n3795), .Z(n4386) );
  XOR U5082 ( .A(n2209), .B(round_reg[1193]), .Z(n3795) );
  XNOR U5083 ( .A(n2223), .B(round_reg[1557]), .Z(n3793) );
  XOR U5084 ( .A(n4387), .B(n4176), .Z(o[1300]) );
  XOR U5085 ( .A(n2070), .B(round_reg[6]), .Z(n4176) );
  AND U5086 ( .A(n3797), .B(n3799), .Z(n4387) );
  XOR U5087 ( .A(n2213), .B(round_reg[1192]), .Z(n3799) );
  XNOR U5088 ( .A(n2227), .B(round_reg[1556]), .Z(n3797) );
  XOR U5089 ( .A(n4388), .B(n1926), .Z(o[12]) );
  XOR U5090 ( .A(n2345), .B(round_reg[202]), .Z(n1926) );
  ANDN U5091 ( .A(n1925), .B(n3423), .Z(n4388) );
  XOR U5092 ( .A(n1769), .B(round_reg[1045]), .Z(n3423) );
  XNOR U5093 ( .A(n2304), .B(round_reg[1422]), .Z(n1925) );
  XOR U5094 ( .A(n4389), .B(n3452), .Z(o[129]) );
  XOR U5095 ( .A(n2014), .B(round_reg[666]), .Z(n3452) );
  IV U5096 ( .A(n4390), .Z(n2014) );
  ANDN U5097 ( .A(n2307), .B(n2308), .Z(n4389) );
  XNOR U5098 ( .A(n2393), .B(round_reg[255]), .Z(n2308) );
  XNOR U5099 ( .A(n2207), .B(round_reg[600]), .Z(n2307) );
  IV U5100 ( .A(n4391), .Z(n2207) );
  XOR U5101 ( .A(n4392), .B(n4178), .Z(o[1299]) );
  XOR U5102 ( .A(n2073), .B(round_reg[5]), .Z(n4178) );
  AND U5103 ( .A(n3801), .B(n3803), .Z(n4392) );
  XOR U5104 ( .A(n2217), .B(round_reg[1191]), .Z(n3803) );
  XNOR U5105 ( .A(n2231), .B(round_reg[1555]), .Z(n3801) );
  XOR U5106 ( .A(n4393), .B(n4180), .Z(o[1298]) );
  XOR U5107 ( .A(n2076), .B(round_reg[4]), .Z(n4180) );
  AND U5108 ( .A(n3805), .B(n3807), .Z(n4393) );
  XOR U5109 ( .A(n2225), .B(round_reg[1190]), .Z(n3807) );
  XNOR U5110 ( .A(n2235), .B(round_reg[1554]), .Z(n3805) );
  XOR U5111 ( .A(n4394), .B(n4182), .Z(o[1297]) );
  XOR U5112 ( .A(n2078), .B(round_reg[3]), .Z(n4182) );
  AND U5113 ( .A(n3809), .B(n3811), .Z(n4394) );
  XOR U5114 ( .A(n2229), .B(round_reg[1189]), .Z(n3811) );
  XNOR U5115 ( .A(n2239), .B(round_reg[1553]), .Z(n3809) );
  XOR U5116 ( .A(n4395), .B(n4184), .Z(o[1296]) );
  XOR U5117 ( .A(n2080), .B(round_reg[2]), .Z(n4184) );
  AND U5118 ( .A(n3813), .B(n3815), .Z(n4395) );
  XOR U5119 ( .A(n2233), .B(round_reg[1188]), .Z(n3815) );
  XNOR U5120 ( .A(n2243), .B(round_reg[1552]), .Z(n3813) );
  XOR U5121 ( .A(n4396), .B(n4186), .Z(o[1295]) );
  XOR U5122 ( .A(n2082), .B(round_reg[1]), .Z(n4186) );
  AND U5123 ( .A(n3817), .B(n3821), .Z(n4396) );
  XOR U5124 ( .A(n2237), .B(round_reg[1187]), .Z(n3821) );
  XNOR U5125 ( .A(n2247), .B(round_reg[1551]), .Z(n3817) );
  XOR U5126 ( .A(n4397), .B(n4188), .Z(o[1294]) );
  XOR U5127 ( .A(n2084), .B(round_reg[0]), .Z(n4188) );
  AND U5128 ( .A(n3834), .B(n3836), .Z(n4397) );
  XOR U5129 ( .A(n2241), .B(round_reg[1186]), .Z(n3836) );
  XNOR U5130 ( .A(n2251), .B(round_reg[1550]), .Z(n3834) );
  XOR U5131 ( .A(n4398), .B(n4190), .Z(o[1293]) );
  XNOR U5132 ( .A(n2086), .B(round_reg[63]), .Z(n4190) );
  AND U5133 ( .A(n3839), .B(n3841), .Z(n4398) );
  XOR U5134 ( .A(n2245), .B(round_reg[1185]), .Z(n3841) );
  XNOR U5135 ( .A(n2255), .B(round_reg[1549]), .Z(n3839) );
  XOR U5136 ( .A(n4399), .B(n4192), .Z(o[1292]) );
  XOR U5137 ( .A(n2088), .B(round_reg[62]), .Z(n4192) );
  AND U5138 ( .A(n3843), .B(n3846), .Z(n4399) );
  XNOR U5139 ( .A(n2249), .B(round_reg[1184]), .Z(n3846) );
  XNOR U5140 ( .A(n2259), .B(round_reg[1548]), .Z(n3843) );
  XOR U5141 ( .A(n4400), .B(n4195), .Z(o[1291]) );
  XOR U5142 ( .A(n2095), .B(round_reg[61]), .Z(n4195) );
  AND U5143 ( .A(n3848), .B(n3850), .Z(n4400) );
  XNOR U5144 ( .A(n2253), .B(round_reg[1183]), .Z(n3850) );
  XNOR U5145 ( .A(n2267), .B(round_reg[1547]), .Z(n3848) );
  XOR U5146 ( .A(n4401), .B(n4197), .Z(o[1290]) );
  XOR U5147 ( .A(n2098), .B(round_reg[60]), .Z(n4197) );
  AND U5148 ( .A(n3852), .B(n3854), .Z(n4401) );
  XNOR U5149 ( .A(n2257), .B(round_reg[1182]), .Z(n3854) );
  XNOR U5150 ( .A(n2271), .B(round_reg[1546]), .Z(n3852) );
  XOR U5151 ( .A(n4402), .B(n3456), .Z(o[128]) );
  XOR U5152 ( .A(n2016), .B(round_reg[665]), .Z(n3456) );
  IV U5153 ( .A(n4403), .Z(n2016) );
  AND U5154 ( .A(n2351), .B(n2353), .Z(n4402) );
  XNOR U5155 ( .A(n2211), .B(round_reg[599]), .Z(n2351) );
  IV U5156 ( .A(n4404), .Z(n2211) );
  XOR U5157 ( .A(n4405), .B(n4199), .Z(o[1289]) );
  XOR U5158 ( .A(n2101), .B(round_reg[59]), .Z(n4199) );
  AND U5159 ( .A(n3856), .B(n3858), .Z(n4405) );
  XNOR U5160 ( .A(n2261), .B(round_reg[1181]), .Z(n3858) );
  XNOR U5161 ( .A(n2275), .B(round_reg[1545]), .Z(n3856) );
  XOR U5162 ( .A(n4406), .B(n4201), .Z(o[1288]) );
  XOR U5163 ( .A(n2104), .B(round_reg[58]), .Z(n4201) );
  AND U5164 ( .A(n3860), .B(n3862), .Z(n4406) );
  XNOR U5165 ( .A(n2269), .B(round_reg[1180]), .Z(n3862) );
  XNOR U5166 ( .A(n2279), .B(round_reg[1544]), .Z(n3860) );
  XOR U5167 ( .A(n4407), .B(n4203), .Z(o[1287]) );
  XOR U5168 ( .A(n2107), .B(round_reg[57]), .Z(n4203) );
  AND U5169 ( .A(n3864), .B(n3868), .Z(n4407) );
  XOR U5170 ( .A(n2273), .B(round_reg[1179]), .Z(n3868) );
  XNOR U5171 ( .A(n2283), .B(round_reg[1543]), .Z(n3864) );
  XOR U5172 ( .A(n4408), .B(n4205), .Z(o[1286]) );
  XNOR U5173 ( .A(n4409), .B(round_reg[56]), .Z(n4205) );
  AND U5174 ( .A(n3880), .B(n3882), .Z(n4408) );
  XOR U5175 ( .A(n2277), .B(round_reg[1178]), .Z(n3882) );
  XNOR U5176 ( .A(n2287), .B(round_reg[1542]), .Z(n3880) );
  XOR U5177 ( .A(n4410), .B(n4207), .Z(o[1285]) );
  XNOR U5178 ( .A(n4411), .B(round_reg[55]), .Z(n4207) );
  ANDN U5179 ( .A(n3886), .B(n3884), .Z(n4410) );
  XOR U5180 ( .A(n2291), .B(round_reg[1541]), .Z(n3884) );
  XOR U5181 ( .A(n2281), .B(round_reg[1177]), .Z(n3886) );
  XOR U5182 ( .A(n4412), .B(n4209), .Z(o[1284]) );
  XNOR U5183 ( .A(n4413), .B(round_reg[54]), .Z(n4209) );
  AND U5184 ( .A(n3888), .B(n3890), .Z(n4412) );
  XOR U5185 ( .A(n2285), .B(round_reg[1176]), .Z(n3890) );
  XNOR U5186 ( .A(n2295), .B(round_reg[1540]), .Z(n3888) );
  XOR U5187 ( .A(n4414), .B(n4211), .Z(o[1283]) );
  XNOR U5188 ( .A(n4415), .B(round_reg[53]), .Z(n4211) );
  AND U5189 ( .A(n3893), .B(n3897), .Z(n4414) );
  XOR U5190 ( .A(n2289), .B(round_reg[1175]), .Z(n3897) );
  XNOR U5191 ( .A(n2299), .B(round_reg[1539]), .Z(n3893) );
  XOR U5192 ( .A(n4416), .B(n4213), .Z(o[1282]) );
  XOR U5193 ( .A(n1940), .B(round_reg[52]), .Z(n4213) );
  AND U5194 ( .A(n3910), .B(n3912), .Z(n4416) );
  XOR U5195 ( .A(n2293), .B(round_reg[1174]), .Z(n3912) );
  XNOR U5196 ( .A(n2303), .B(round_reg[1538]), .Z(n3910) );
  XOR U5197 ( .A(n4417), .B(n4216), .Z(o[1281]) );
  XOR U5198 ( .A(n1943), .B(round_reg[51]), .Z(n4216) );
  AND U5199 ( .A(n3914), .B(n3918), .Z(n4417) );
  XOR U5200 ( .A(n2297), .B(round_reg[1173]), .Z(n3918) );
  XNOR U5201 ( .A(n2311), .B(round_reg[1537]), .Z(n3914) );
  XOR U5202 ( .A(n4418), .B(n4218), .Z(o[1280]) );
  XOR U5203 ( .A(n1946), .B(round_reg[50]), .Z(n4218) );
  AND U5204 ( .A(n3927), .B(n3931), .Z(n4418) );
  XOR U5205 ( .A(n2301), .B(round_reg[1172]), .Z(n3931) );
  XNOR U5206 ( .A(n2315), .B(round_reg[1536]), .Z(n3927) );
  XOR U5207 ( .A(n4419), .B(n3459), .Z(o[127]) );
  XOR U5208 ( .A(n2215), .B(round_reg[598]), .Z(n3459) );
  IV U5209 ( .A(n4420), .Z(n2215) );
  ANDN U5210 ( .A(n2395), .B(n2396), .Z(n4419) );
  XNOR U5211 ( .A(n2364), .B(round_reg[1409]), .Z(n2396) );
  XNOR U5212 ( .A(n2117), .B(round_reg[253]), .Z(n2395) );
  XOR U5213 ( .A(n4421), .B(n4422), .Z(o[1279]) );
  XOR U5214 ( .A(n4425), .B(n4426), .Z(o[1278]) );
  XOR U5215 ( .A(n4429), .B(n4430), .Z(o[1277]) );
  ANDN U5216 ( .A(n4431), .B(n4432), .Z(n4429) );
  XOR U5217 ( .A(n4433), .B(n4434), .Z(o[1276]) );
  ANDN U5218 ( .A(n4435), .B(n4436), .Z(n4433) );
  XOR U5219 ( .A(n4437), .B(n4438), .Z(o[1275]) );
  ANDN U5220 ( .A(n4439), .B(n4440), .Z(n4437) );
  XOR U5221 ( .A(n4441), .B(n4442), .Z(o[1274]) );
  ANDN U5222 ( .A(n4443), .B(n4444), .Z(n4441) );
  XOR U5223 ( .A(n4445), .B(n4446), .Z(o[1273]) );
  ANDN U5224 ( .A(n4447), .B(n4448), .Z(n4445) );
  XOR U5225 ( .A(n4449), .B(n4450), .Z(o[1272]) );
  ANDN U5226 ( .A(n4451), .B(n4452), .Z(n4449) );
  XOR U5227 ( .A(n4453), .B(n4454), .Z(o[1271]) );
  ANDN U5228 ( .A(n4455), .B(n4456), .Z(n4453) );
  XOR U5229 ( .A(n4457), .B(n4458), .Z(o[1270]) );
  ANDN U5230 ( .A(n4459), .B(n4460), .Z(n4457) );
  XOR U5231 ( .A(n4461), .B(n3461), .Z(o[126]) );
  XOR U5232 ( .A(n2223), .B(round_reg[597]), .Z(n3461) );
  IV U5233 ( .A(n4462), .Z(n2223) );
  ANDN U5234 ( .A(n2439), .B(n2440), .Z(n4461) );
  XNOR U5235 ( .A(n2368), .B(round_reg[1408]), .Z(n2440) );
  XNOR U5236 ( .A(n2121), .B(round_reg[252]), .Z(n2439) );
  XOR U5237 ( .A(n4463), .B(n4464), .Z(o[1269]) );
  ANDN U5238 ( .A(n4465), .B(n4466), .Z(n4463) );
  XOR U5239 ( .A(n4467), .B(n4468), .Z(o[1268]) );
  ANDN U5240 ( .A(n4469), .B(n4470), .Z(n4467) );
  XOR U5241 ( .A(n4471), .B(n4472), .Z(o[1267]) );
  ANDN U5242 ( .A(n4473), .B(n4474), .Z(n4471) );
  XOR U5243 ( .A(n4475), .B(n4476), .Z(o[1266]) );
  ANDN U5244 ( .A(n4477), .B(n4478), .Z(n4475) );
  XOR U5245 ( .A(n4479), .B(n4480), .Z(o[1265]) );
  ANDN U5246 ( .A(n4481), .B(n4482), .Z(n4479) );
  XOR U5247 ( .A(n4483), .B(n4484), .Z(o[1264]) );
  ANDN U5248 ( .A(n4485), .B(n4486), .Z(n4483) );
  XOR U5249 ( .A(n4487), .B(n4488), .Z(o[1263]) );
  ANDN U5250 ( .A(n4489), .B(n4490), .Z(n4487) );
  XOR U5251 ( .A(n4491), .B(n4492), .Z(o[1262]) );
  ANDN U5252 ( .A(n4493), .B(n4494), .Z(n4491) );
  XOR U5253 ( .A(n4495), .B(n4496), .Z(o[1261]) );
  ANDN U5254 ( .A(n4497), .B(n4498), .Z(n4495) );
  XOR U5255 ( .A(n4499), .B(n4500), .Z(o[1260]) );
  ANDN U5256 ( .A(n4501), .B(n4502), .Z(n4499) );
  XOR U5257 ( .A(n4503), .B(n3463), .Z(o[125]) );
  XOR U5258 ( .A(n2227), .B(round_reg[596]), .Z(n3463) );
  IV U5259 ( .A(n4504), .Z(n2227) );
  ANDN U5260 ( .A(n2483), .B(n2484), .Z(n4503) );
  XNOR U5261 ( .A(n2372), .B(round_reg[1471]), .Z(n2484) );
  XNOR U5262 ( .A(n2125), .B(round_reg[251]), .Z(n2483) );
  XOR U5263 ( .A(n4505), .B(n4506), .Z(o[1259]) );
  ANDN U5264 ( .A(n4507), .B(n4508), .Z(n4505) );
  XOR U5265 ( .A(n4509), .B(n4510), .Z(o[1258]) );
  ANDN U5266 ( .A(n4511), .B(n4512), .Z(n4509) );
  XOR U5267 ( .A(n4513), .B(n4514), .Z(o[1257]) );
  ANDN U5268 ( .A(n4515), .B(n4516), .Z(n4513) );
  XOR U5269 ( .A(n4517), .B(n4518), .Z(o[1256]) );
  ANDN U5270 ( .A(n4519), .B(n4520), .Z(n4517) );
  XOR U5271 ( .A(n4521), .B(n1062), .Z(o[1255]) );
  ANDN U5272 ( .A(n4522), .B(n1061), .Z(n4521) );
  XNOR U5273 ( .A(n4523), .B(n1066), .Z(o[1254]) );
  ANDN U5274 ( .A(n4524), .B(n1065), .Z(n4523) );
  XOR U5275 ( .A(n4525), .B(n1070), .Z(o[1253]) );
  ANDN U5276 ( .A(n4526), .B(n1069), .Z(n4525) );
  XOR U5277 ( .A(n4527), .B(n1074), .Z(o[1252]) );
  ANDN U5278 ( .A(n4528), .B(n1073), .Z(n4527) );
  XOR U5279 ( .A(n4529), .B(n1078), .Z(o[1251]) );
  ANDN U5280 ( .A(n4530), .B(n1077), .Z(n4529) );
  XOR U5281 ( .A(n4531), .B(n1082), .Z(o[1250]) );
  ANDN U5282 ( .A(n4532), .B(n1081), .Z(n4531) );
  XOR U5283 ( .A(n4533), .B(n3465), .Z(o[124]) );
  XOR U5284 ( .A(n2231), .B(round_reg[595]), .Z(n3465) );
  IV U5285 ( .A(n4534), .Z(n2231) );
  ANDN U5286 ( .A(n2527), .B(n2528), .Z(n4533) );
  XNOR U5287 ( .A(n2376), .B(round_reg[1470]), .Z(n2528) );
  XNOR U5288 ( .A(n2136), .B(round_reg[250]), .Z(n2527) );
  XOR U5289 ( .A(n4535), .B(n1086), .Z(o[1249]) );
  ANDN U5290 ( .A(n4536), .B(n1085), .Z(n4535) );
  XOR U5291 ( .A(n4537), .B(n1090), .Z(o[1248]) );
  ANDN U5292 ( .A(n4538), .B(n1089), .Z(n4537) );
  XOR U5293 ( .A(n4539), .B(n1094), .Z(o[1247]) );
  ANDN U5294 ( .A(n4540), .B(n1093), .Z(n4539) );
  XOR U5295 ( .A(n4541), .B(n1098), .Z(o[1246]) );
  ANDN U5296 ( .A(n4542), .B(n1097), .Z(n4541) );
  XOR U5297 ( .A(n4543), .B(n1106), .Z(o[1245]) );
  ANDN U5298 ( .A(n4544), .B(n1105), .Z(n4543) );
  XOR U5299 ( .A(n4545), .B(n1110), .Z(o[1244]) );
  ANDN U5300 ( .A(n4546), .B(n1109), .Z(n4545) );
  XOR U5301 ( .A(n4547), .B(n1114), .Z(o[1243]) );
  ANDN U5302 ( .A(n4548), .B(n1113), .Z(n4547) );
  XOR U5303 ( .A(n4549), .B(n1118), .Z(o[1242]) );
  ANDN U5304 ( .A(n4550), .B(n1117), .Z(n4549) );
  XOR U5305 ( .A(n4551), .B(n1122), .Z(o[1241]) );
  ANDN U5306 ( .A(n4552), .B(n1121), .Z(n4551) );
  XOR U5307 ( .A(n4553), .B(n1126), .Z(o[1240]) );
  ANDN U5308 ( .A(n4554), .B(n1125), .Z(n4553) );
  XOR U5309 ( .A(n4555), .B(n3467), .Z(o[123]) );
  XOR U5310 ( .A(n2235), .B(round_reg[594]), .Z(n3467) );
  IV U5311 ( .A(n4556), .Z(n2235) );
  ANDN U5312 ( .A(n2574), .B(n2575), .Z(n4555) );
  XNOR U5313 ( .A(n2380), .B(round_reg[1469]), .Z(n2575) );
  XNOR U5314 ( .A(n2141), .B(round_reg[249]), .Z(n2574) );
  XOR U5315 ( .A(n4557), .B(n1130), .Z(o[1239]) );
  ANDN U5316 ( .A(n4558), .B(n1129), .Z(n4557) );
  XOR U5317 ( .A(n4559), .B(n1134), .Z(o[1238]) );
  ANDN U5318 ( .A(n4560), .B(n1133), .Z(n4559) );
  XOR U5319 ( .A(n4561), .B(n1138), .Z(o[1237]) );
  ANDN U5320 ( .A(n4562), .B(n1137), .Z(n4561) );
  XOR U5321 ( .A(n4563), .B(n1142), .Z(o[1236]) );
  ANDN U5322 ( .A(n4564), .B(n1141), .Z(n4563) );
  XOR U5323 ( .A(n4565), .B(n1150), .Z(o[1235]) );
  AND U5324 ( .A(n4566), .B(n1149), .Z(n4565) );
  IV U5325 ( .A(n4567), .Z(n1149) );
  XOR U5326 ( .A(n4568), .B(n1154), .Z(o[1234]) );
  ANDN U5327 ( .A(n4569), .B(n1153), .Z(n4568) );
  XOR U5328 ( .A(n4570), .B(n1158), .Z(o[1233]) );
  ANDN U5329 ( .A(n4571), .B(n1157), .Z(n4570) );
  XOR U5330 ( .A(n4572), .B(n1162), .Z(o[1232]) );
  ANDN U5331 ( .A(n4573), .B(n1161), .Z(n4572) );
  XOR U5332 ( .A(n4574), .B(n1166), .Z(o[1231]) );
  ANDN U5333 ( .A(n4575), .B(n1165), .Z(n4574) );
  XOR U5334 ( .A(n4576), .B(n1170), .Z(o[1230]) );
  ANDN U5335 ( .A(n4577), .B(n1169), .Z(n4576) );
  XOR U5336 ( .A(n4578), .B(n3469), .Z(o[122]) );
  XOR U5337 ( .A(n2239), .B(round_reg[593]), .Z(n3469) );
  IV U5338 ( .A(n4579), .Z(n2239) );
  ANDN U5339 ( .A(n2618), .B(n2619), .Z(n4578) );
  XNOR U5340 ( .A(n2384), .B(round_reg[1468]), .Z(n2619) );
  XNOR U5341 ( .A(n2145), .B(round_reg[248]), .Z(n2618) );
  XOR U5342 ( .A(n4580), .B(n1174), .Z(o[1229]) );
  ANDN U5343 ( .A(n4581), .B(n1173), .Z(n4580) );
  XOR U5344 ( .A(n4582), .B(n1178), .Z(o[1228]) );
  AND U5345 ( .A(n4583), .B(n1177), .Z(n4582) );
  IV U5346 ( .A(n4584), .Z(n1177) );
  XOR U5347 ( .A(n4585), .B(n1182), .Z(o[1227]) );
  AND U5348 ( .A(n4586), .B(n1181), .Z(n4585) );
  IV U5349 ( .A(n4587), .Z(n1181) );
  XOR U5350 ( .A(n4588), .B(n1186), .Z(o[1226]) );
  AND U5351 ( .A(n4589), .B(n1185), .Z(n4588) );
  IV U5352 ( .A(n4590), .Z(n1185) );
  XOR U5353 ( .A(n4591), .B(n1194), .Z(o[1225]) );
  AND U5354 ( .A(n4592), .B(n1193), .Z(n4591) );
  IV U5355 ( .A(n4593), .Z(n1193) );
  XOR U5356 ( .A(n4594), .B(n1198), .Z(o[1224]) );
  ANDN U5357 ( .A(n4595), .B(n1197), .Z(n4594) );
  XOR U5358 ( .A(n4596), .B(n1202), .Z(o[1223]) );
  ANDN U5359 ( .A(n4597), .B(n1201), .Z(n4596) );
  XOR U5360 ( .A(n4598), .B(n1206), .Z(o[1222]) );
  ANDN U5361 ( .A(n4599), .B(n1205), .Z(n4598) );
  XNOR U5362 ( .A(n4600), .B(n1209), .Z(o[1221]) );
  AND U5363 ( .A(n4601), .B(n4602), .Z(n4600) );
  XNOR U5364 ( .A(n4603), .B(n1213), .Z(o[1220]) );
  AND U5365 ( .A(n4604), .B(n4605), .Z(n4603) );
  XOR U5366 ( .A(n4606), .B(n3472), .Z(o[121]) );
  XOR U5367 ( .A(n2243), .B(round_reg[592]), .Z(n3472) );
  IV U5368 ( .A(n4607), .Z(n2243) );
  ANDN U5369 ( .A(n2662), .B(n2663), .Z(n4606) );
  XNOR U5370 ( .A(n2388), .B(round_reg[1467]), .Z(n2663) );
  XNOR U5371 ( .A(n2149), .B(round_reg[247]), .Z(n2662) );
  XNOR U5372 ( .A(n4608), .B(n1217), .Z(o[1219]) );
  AND U5373 ( .A(n4609), .B(n4610), .Z(n4608) );
  XNOR U5374 ( .A(n4611), .B(n1221), .Z(o[1218]) );
  AND U5375 ( .A(n4612), .B(n4613), .Z(n4611) );
  XNOR U5376 ( .A(n4614), .B(n1225), .Z(o[1217]) );
  AND U5377 ( .A(n4615), .B(n4616), .Z(n4614) );
  XNOR U5378 ( .A(n4617), .B(n1229), .Z(o[1216]) );
  AND U5379 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U5380 ( .A(n4620), .B(n4424), .Z(o[1215]) );
  ANDN U5381 ( .A(n4621), .B(n4423), .Z(n4620) );
  XOR U5382 ( .A(n4622), .B(n4428), .Z(o[1214]) );
  ANDN U5383 ( .A(n4623), .B(n4427), .Z(n4622) );
  XOR U5384 ( .A(n4624), .B(n4432), .Z(o[1213]) );
  ANDN U5385 ( .A(n4625), .B(n4431), .Z(n4624) );
  XOR U5386 ( .A(n4626), .B(n4436), .Z(o[1212]) );
  ANDN U5387 ( .A(n4627), .B(n4435), .Z(n4626) );
  XOR U5388 ( .A(n4628), .B(n4440), .Z(o[1211]) );
  ANDN U5389 ( .A(n4629), .B(n4439), .Z(n4628) );
  XOR U5390 ( .A(n4630), .B(n4444), .Z(o[1210]) );
  ANDN U5391 ( .A(n4631), .B(n4443), .Z(n4630) );
  XOR U5392 ( .A(n4632), .B(n3474), .Z(o[120]) );
  XOR U5393 ( .A(n2247), .B(round_reg[591]), .Z(n3474) );
  IV U5394 ( .A(n4633), .Z(n2247) );
  ANDN U5395 ( .A(n2700), .B(n2701), .Z(n4632) );
  XNOR U5396 ( .A(n2392), .B(round_reg[1466]), .Z(n2701) );
  XNOR U5397 ( .A(n2153), .B(round_reg[246]), .Z(n2700) );
  XOR U5398 ( .A(n4634), .B(n4448), .Z(o[1209]) );
  ANDN U5399 ( .A(n4635), .B(n4447), .Z(n4634) );
  XOR U5400 ( .A(n4636), .B(n4452), .Z(o[1208]) );
  ANDN U5401 ( .A(n4637), .B(n4451), .Z(n4636) );
  XOR U5402 ( .A(n4638), .B(n4456), .Z(o[1207]) );
  ANDN U5403 ( .A(n4639), .B(n4455), .Z(n4638) );
  XOR U5404 ( .A(n4640), .B(n4460), .Z(o[1206]) );
  ANDN U5405 ( .A(n4641), .B(n4459), .Z(n4640) );
  XOR U5406 ( .A(n4642), .B(n4466), .Z(o[1205]) );
  ANDN U5407 ( .A(n4643), .B(n4465), .Z(n4642) );
  XOR U5408 ( .A(n4644), .B(n4470), .Z(o[1204]) );
  ANDN U5409 ( .A(n4645), .B(n4469), .Z(n4644) );
  XOR U5410 ( .A(n4646), .B(n4474), .Z(o[1203]) );
  ANDN U5411 ( .A(n4647), .B(n4473), .Z(n4646) );
  XOR U5412 ( .A(n4648), .B(n4478), .Z(o[1202]) );
  ANDN U5413 ( .A(n4649), .B(n4477), .Z(n4648) );
  XOR U5414 ( .A(n4650), .B(n4482), .Z(o[1201]) );
  ANDN U5415 ( .A(n4651), .B(n4481), .Z(n4650) );
  XOR U5416 ( .A(n4652), .B(n4486), .Z(o[1200]) );
  ANDN U5417 ( .A(n4653), .B(n4485), .Z(n4652) );
  XOR U5418 ( .A(n4654), .B(n1957), .Z(o[11]) );
  XOR U5419 ( .A(n2349), .B(round_reg[201]), .Z(n1957) );
  ANDN U5420 ( .A(n1956), .B(n3426), .Z(n4654) );
  XOR U5421 ( .A(n1772), .B(round_reg[1044]), .Z(n3426) );
  XNOR U5422 ( .A(n2312), .B(round_reg[1421]), .Z(n1956) );
  XOR U5423 ( .A(n4655), .B(n3476), .Z(o[119]) );
  XOR U5424 ( .A(n2251), .B(round_reg[590]), .Z(n3476) );
  IV U5425 ( .A(n4656), .Z(n2251) );
  ANDN U5426 ( .A(n2734), .B(n2735), .Z(n4655) );
  XNOR U5427 ( .A(n2114), .B(round_reg[1465]), .Z(n2735) );
  IV U5428 ( .A(n4657), .Z(n2114) );
  XNOR U5429 ( .A(n2157), .B(round_reg[245]), .Z(n2734) );
  XOR U5430 ( .A(n4658), .B(n4490), .Z(o[1199]) );
  ANDN U5431 ( .A(n4659), .B(n4489), .Z(n4658) );
  XOR U5432 ( .A(n4660), .B(n4494), .Z(o[1198]) );
  ANDN U5433 ( .A(n4661), .B(n4493), .Z(n4660) );
  XOR U5434 ( .A(n4662), .B(n4498), .Z(o[1197]) );
  ANDN U5435 ( .A(n4663), .B(n4497), .Z(n4662) );
  XOR U5436 ( .A(n4664), .B(n4502), .Z(o[1196]) );
  ANDN U5437 ( .A(n4665), .B(n4501), .Z(n4664) );
  XOR U5438 ( .A(n4666), .B(n4508), .Z(o[1195]) );
  ANDN U5439 ( .A(n4667), .B(n4507), .Z(n4666) );
  XOR U5440 ( .A(n4668), .B(n4512), .Z(o[1194]) );
  ANDN U5441 ( .A(n4669), .B(n4511), .Z(n4668) );
  XOR U5442 ( .A(n4670), .B(n4516), .Z(o[1193]) );
  ANDN U5443 ( .A(n4671), .B(n4515), .Z(n4670) );
  XOR U5444 ( .A(n4672), .B(n4520), .Z(o[1192]) );
  ANDN U5445 ( .A(n4673), .B(n4519), .Z(n4672) );
  XOR U5446 ( .A(n4674), .B(n1061), .Z(o[1191]) );
  XOR U5447 ( .A(n2028), .B(round_reg[979]), .Z(n1061) );
  XOR U5448 ( .A(n4675), .B(n4676), .Z(n2028) );
  ANDN U5449 ( .A(n4677), .B(n4522), .Z(n4674) );
  XOR U5450 ( .A(n4678), .B(n1065), .Z(o[1190]) );
  XOR U5451 ( .A(n2031), .B(round_reg[978]), .Z(n1065) );
  XOR U5452 ( .A(n4679), .B(n4680), .Z(n2031) );
  ANDN U5453 ( .A(n4681), .B(n4524), .Z(n4678) );
  XOR U5454 ( .A(n4682), .B(n3478), .Z(o[118]) );
  XOR U5455 ( .A(n2255), .B(round_reg[589]), .Z(n3478) );
  IV U5456 ( .A(n4683), .Z(n2255) );
  ANDN U5457 ( .A(n2763), .B(n2764), .Z(n4682) );
  XNOR U5458 ( .A(n2118), .B(round_reg[1464]), .Z(n2764) );
  IV U5459 ( .A(n4684), .Z(n2118) );
  XNOR U5460 ( .A(n2161), .B(round_reg[244]), .Z(n2763) );
  XOR U5461 ( .A(n4685), .B(n1069), .Z(o[1189]) );
  XOR U5462 ( .A(n2036), .B(round_reg[977]), .Z(n1069) );
  XOR U5463 ( .A(n4686), .B(n4687), .Z(n2036) );
  ANDN U5464 ( .A(n4688), .B(n4526), .Z(n4685) );
  XOR U5465 ( .A(n4689), .B(n1073), .Z(o[1188]) );
  XOR U5466 ( .A(n2039), .B(round_reg[976]), .Z(n1073) );
  XOR U5467 ( .A(n4690), .B(n4691), .Z(n2039) );
  ANDN U5468 ( .A(n4692), .B(n4528), .Z(n4689) );
  XOR U5469 ( .A(n4693), .B(n1077), .Z(o[1187]) );
  XOR U5470 ( .A(n2042), .B(round_reg[975]), .Z(n1077) );
  XOR U5471 ( .A(n4694), .B(n4695), .Z(n2042) );
  ANDN U5472 ( .A(n4696), .B(n4530), .Z(n4693) );
  XOR U5473 ( .A(n4697), .B(n1081), .Z(o[1186]) );
  XOR U5474 ( .A(n2044), .B(round_reg[974]), .Z(n1081) );
  XOR U5475 ( .A(n4698), .B(n4699), .Z(n2044) );
  ANDN U5476 ( .A(n4700), .B(n4532), .Z(n4697) );
  XOR U5477 ( .A(n4701), .B(n1085), .Z(o[1185]) );
  XOR U5478 ( .A(n2047), .B(round_reg[973]), .Z(n1085) );
  XNOR U5479 ( .A(n4702), .B(n4703), .Z(n2047) );
  ANDN U5480 ( .A(n4704), .B(n4536), .Z(n4701) );
  XOR U5481 ( .A(n4705), .B(n1089), .Z(o[1184]) );
  XOR U5482 ( .A(n2050), .B(round_reg[972]), .Z(n1089) );
  XNOR U5483 ( .A(n4706), .B(n4707), .Z(n2050) );
  ANDN U5484 ( .A(n4708), .B(n4538), .Z(n4705) );
  XOR U5485 ( .A(n4709), .B(n1093), .Z(o[1183]) );
  XOR U5486 ( .A(n2053), .B(round_reg[971]), .Z(n1093) );
  XNOR U5487 ( .A(n4710), .B(n4711), .Z(n2053) );
  ANDN U5488 ( .A(n4712), .B(n4540), .Z(n4709) );
  XOR U5489 ( .A(n4713), .B(n1097), .Z(o[1182]) );
  XOR U5490 ( .A(n2056), .B(round_reg[970]), .Z(n1097) );
  XNOR U5491 ( .A(n4714), .B(n4715), .Z(n2056) );
  ANDN U5492 ( .A(n4716), .B(n4542), .Z(n4713) );
  XOR U5493 ( .A(n4717), .B(n1105), .Z(o[1181]) );
  XOR U5494 ( .A(n2059), .B(round_reg[969]), .Z(n1105) );
  XNOR U5495 ( .A(n4718), .B(n4719), .Z(n2059) );
  ANDN U5496 ( .A(n4720), .B(n4544), .Z(n4717) );
  XOR U5497 ( .A(n4721), .B(n1109), .Z(o[1180]) );
  XOR U5498 ( .A(n2062), .B(round_reg[968]), .Z(n1109) );
  XOR U5499 ( .A(n4722), .B(n4723), .Z(n2062) );
  ANDN U5500 ( .A(n4724), .B(n4546), .Z(n4721) );
  XOR U5501 ( .A(n4725), .B(n3480), .Z(o[117]) );
  XOR U5502 ( .A(n2259), .B(round_reg[588]), .Z(n3480) );
  IV U5503 ( .A(n4726), .Z(n2259) );
  ANDN U5504 ( .A(n2797), .B(n2798), .Z(n4725) );
  XNOR U5505 ( .A(n2122), .B(round_reg[1463]), .Z(n2798) );
  IV U5506 ( .A(n4727), .Z(n2122) );
  XNOR U5507 ( .A(n2165), .B(round_reg[243]), .Z(n2797) );
  XOR U5508 ( .A(n4728), .B(n1113), .Z(o[1179]) );
  XOR U5509 ( .A(n2067), .B(round_reg[967]), .Z(n1113) );
  XNOR U5510 ( .A(n4729), .B(n4730), .Z(n2067) );
  ANDN U5511 ( .A(n4731), .B(n4548), .Z(n4728) );
  XOR U5512 ( .A(n4732), .B(n1117), .Z(o[1178]) );
  XOR U5513 ( .A(n2070), .B(round_reg[966]), .Z(n1117) );
  XNOR U5514 ( .A(n4733), .B(n4734), .Z(n2070) );
  ANDN U5515 ( .A(n4735), .B(n4550), .Z(n4732) );
  XOR U5516 ( .A(n4736), .B(n1121), .Z(o[1177]) );
  XOR U5517 ( .A(n2073), .B(round_reg[965]), .Z(n1121) );
  XNOR U5518 ( .A(n4737), .B(n4738), .Z(n2073) );
  ANDN U5519 ( .A(n4739), .B(n4552), .Z(n4736) );
  XOR U5520 ( .A(n4740), .B(n1125), .Z(o[1176]) );
  XOR U5521 ( .A(n2076), .B(round_reg[964]), .Z(n1125) );
  XNOR U5522 ( .A(n4741), .B(n4742), .Z(n2076) );
  ANDN U5523 ( .A(n4743), .B(n4554), .Z(n4740) );
  XOR U5524 ( .A(n4744), .B(n1129), .Z(o[1175]) );
  XOR U5525 ( .A(n2078), .B(round_reg[963]), .Z(n1129) );
  XNOR U5526 ( .A(n4745), .B(n4746), .Z(n2078) );
  ANDN U5527 ( .A(n4747), .B(n4558), .Z(n4744) );
  XOR U5528 ( .A(n4748), .B(n1133), .Z(o[1174]) );
  XOR U5529 ( .A(n2080), .B(round_reg[962]), .Z(n1133) );
  XNOR U5530 ( .A(n4749), .B(n4750), .Z(n2080) );
  ANDN U5531 ( .A(n4751), .B(n4560), .Z(n4748) );
  XOR U5532 ( .A(n4752), .B(n1137), .Z(o[1173]) );
  XOR U5533 ( .A(n2082), .B(round_reg[961]), .Z(n1137) );
  XNOR U5534 ( .A(n4753), .B(n4754), .Z(n2082) );
  ANDN U5535 ( .A(n4755), .B(n4562), .Z(n4752) );
  XOR U5536 ( .A(n4756), .B(n1141), .Z(o[1172]) );
  XOR U5537 ( .A(n2084), .B(round_reg[960]), .Z(n1141) );
  XNOR U5538 ( .A(n4757), .B(n4758), .Z(n2084) );
  ANDN U5539 ( .A(n4759), .B(n4564), .Z(n4756) );
  XOR U5540 ( .A(n4760), .B(n4567), .Z(o[1171]) );
  XNOR U5541 ( .A(n2086), .B(round_reg[1023]), .Z(n4567) );
  ANDN U5542 ( .A(n4763), .B(n4566), .Z(n4760) );
  XOR U5543 ( .A(n4764), .B(n1153), .Z(o[1170]) );
  XOR U5544 ( .A(n2088), .B(round_reg[1022]), .Z(n1153) );
  XNOR U5545 ( .A(n4765), .B(n4766), .Z(n2088) );
  ANDN U5546 ( .A(n4767), .B(n4569), .Z(n4764) );
  XOR U5547 ( .A(n4768), .B(n3482), .Z(o[116]) );
  XOR U5548 ( .A(n2267), .B(round_reg[587]), .Z(n3482) );
  IV U5549 ( .A(n4769), .Z(n2267) );
  ANDN U5550 ( .A(n2831), .B(n2832), .Z(n4768) );
  XNOR U5551 ( .A(n2126), .B(round_reg[1462]), .Z(n2832) );
  IV U5552 ( .A(n4770), .Z(n2126) );
  XNOR U5553 ( .A(n2169), .B(round_reg[242]), .Z(n2831) );
  XOR U5554 ( .A(n4771), .B(n1157), .Z(o[1169]) );
  XOR U5555 ( .A(n2095), .B(round_reg[1021]), .Z(n1157) );
  XNOR U5556 ( .A(n4772), .B(n4773), .Z(n2095) );
  ANDN U5557 ( .A(n4774), .B(n4571), .Z(n4771) );
  XOR U5558 ( .A(n4775), .B(n1161), .Z(o[1168]) );
  XOR U5559 ( .A(n2098), .B(round_reg[1020]), .Z(n1161) );
  XNOR U5560 ( .A(n4776), .B(n4777), .Z(n2098) );
  ANDN U5561 ( .A(n4778), .B(n4573), .Z(n4775) );
  XOR U5562 ( .A(n4779), .B(n1165), .Z(o[1167]) );
  XOR U5563 ( .A(n2101), .B(round_reg[1019]), .Z(n1165) );
  XNOR U5564 ( .A(n4780), .B(n4781), .Z(n2101) );
  ANDN U5565 ( .A(n4782), .B(n4575), .Z(n4779) );
  XOR U5566 ( .A(n4783), .B(n1169), .Z(o[1166]) );
  XOR U5567 ( .A(n2104), .B(round_reg[1018]), .Z(n1169) );
  XNOR U5568 ( .A(n4784), .B(n4785), .Z(n2104) );
  ANDN U5569 ( .A(n4786), .B(n4577), .Z(n4783) );
  XOR U5570 ( .A(n4787), .B(n1173), .Z(o[1165]) );
  XOR U5571 ( .A(n2107), .B(round_reg[1017]), .Z(n1173) );
  XNOR U5572 ( .A(n4788), .B(n4789), .Z(n2107) );
  ANDN U5573 ( .A(n4790), .B(n4581), .Z(n4787) );
  XOR U5574 ( .A(n4791), .B(n4584), .Z(o[1164]) );
  XOR U5575 ( .A(n2110), .B(round_reg[1016]), .Z(n4584) );
  IV U5576 ( .A(n4409), .Z(n2110) );
  ANDN U5577 ( .A(n4794), .B(n4583), .Z(n4791) );
  XOR U5578 ( .A(n4795), .B(n4587), .Z(o[1163]) );
  XOR U5579 ( .A(n1934), .B(round_reg[1015]), .Z(n4587) );
  IV U5580 ( .A(n4411), .Z(n1934) );
  ANDN U5581 ( .A(n4798), .B(n4586), .Z(n4795) );
  XOR U5582 ( .A(n4799), .B(n4590), .Z(o[1162]) );
  XOR U5583 ( .A(n1936), .B(round_reg[1014]), .Z(n4590) );
  IV U5584 ( .A(n4413), .Z(n1936) );
  ANDN U5585 ( .A(n4802), .B(n4589), .Z(n4799) );
  XOR U5586 ( .A(n4803), .B(n4593), .Z(o[1161]) );
  XOR U5587 ( .A(n1938), .B(round_reg[1013]), .Z(n4593) );
  IV U5588 ( .A(n4415), .Z(n1938) );
  ANDN U5589 ( .A(n4806), .B(n4592), .Z(n4803) );
  XOR U5590 ( .A(n4807), .B(n1197), .Z(o[1160]) );
  XOR U5591 ( .A(n1940), .B(round_reg[1012]), .Z(n1197) );
  XNOR U5592 ( .A(n4808), .B(n4809), .Z(n1940) );
  ANDN U5593 ( .A(n4810), .B(n4595), .Z(n4807) );
  XOR U5594 ( .A(n4811), .B(n3484), .Z(o[115]) );
  XOR U5595 ( .A(n2271), .B(round_reg[586]), .Z(n3484) );
  IV U5596 ( .A(n4812), .Z(n2271) );
  ANDN U5597 ( .A(n2864), .B(n2865), .Z(n4811) );
  XNOR U5598 ( .A(n2137), .B(round_reg[1461]), .Z(n2865) );
  IV U5599 ( .A(n4813), .Z(n2137) );
  XNOR U5600 ( .A(n2173), .B(round_reg[241]), .Z(n2864) );
  XOR U5601 ( .A(n4814), .B(n1201), .Z(o[1159]) );
  XOR U5602 ( .A(n1943), .B(round_reg[1011]), .Z(n1201) );
  XNOR U5603 ( .A(n4815), .B(n4816), .Z(n1943) );
  ANDN U5604 ( .A(n4817), .B(n4597), .Z(n4814) );
  XOR U5605 ( .A(n4818), .B(n1205), .Z(o[1158]) );
  XOR U5606 ( .A(n1946), .B(round_reg[1010]), .Z(n1205) );
  XNOR U5607 ( .A(n4819), .B(n4820), .Z(n1946) );
  ANDN U5608 ( .A(n4821), .B(n4599), .Z(n4818) );
  XOR U5609 ( .A(n4822), .B(n1210), .Z(o[1157]) );
  IV U5610 ( .A(n4602), .Z(n1210) );
  XNOR U5611 ( .A(n1949), .B(round_reg[1009]), .Z(n4602) );
  XNOR U5612 ( .A(n4823), .B(n4824), .Z(n1949) );
  ANDN U5613 ( .A(n4825), .B(n4601), .Z(n4822) );
  XOR U5614 ( .A(n4826), .B(n1214), .Z(o[1156]) );
  IV U5615 ( .A(n4605), .Z(n1214) );
  XNOR U5616 ( .A(n1952), .B(round_reg[1008]), .Z(n4605) );
  XNOR U5617 ( .A(n4827), .B(n4828), .Z(n1952) );
  ANDN U5618 ( .A(n4829), .B(n4604), .Z(n4826) );
  XOR U5619 ( .A(n4830), .B(n1218), .Z(o[1155]) );
  IV U5620 ( .A(n4610), .Z(n1218) );
  XNOR U5621 ( .A(n1959), .B(round_reg[1007]), .Z(n4610) );
  XNOR U5622 ( .A(n4831), .B(n4832), .Z(n1959) );
  ANDN U5623 ( .A(n4833), .B(n4609), .Z(n4830) );
  XOR U5624 ( .A(n4834), .B(n1222), .Z(o[1154]) );
  IV U5625 ( .A(n4613), .Z(n1222) );
  XNOR U5626 ( .A(n1962), .B(round_reg[1006]), .Z(n4613) );
  XNOR U5627 ( .A(n4835), .B(n4836), .Z(n1962) );
  ANDN U5628 ( .A(n4837), .B(n4612), .Z(n4834) );
  XOR U5629 ( .A(n4838), .B(n1226), .Z(o[1153]) );
  IV U5630 ( .A(n4616), .Z(n1226) );
  XNOR U5631 ( .A(n1965), .B(round_reg[1005]), .Z(n4616) );
  XNOR U5632 ( .A(n4839), .B(n4840), .Z(n1965) );
  ANDN U5633 ( .A(n4841), .B(n4615), .Z(n4838) );
  XOR U5634 ( .A(n4842), .B(n1230), .Z(o[1152]) );
  IV U5635 ( .A(n4619), .Z(n1230) );
  XNOR U5636 ( .A(n1968), .B(round_reg[1004]), .Z(n4619) );
  XNOR U5637 ( .A(n4843), .B(n4844), .Z(n1968) );
  ANDN U5638 ( .A(n4845), .B(n4618), .Z(n4842) );
  XOR U5639 ( .A(n4846), .B(n4423), .Z(o[1151]) );
  XNOR U5640 ( .A(n4847), .B(round_reg[956]), .Z(n4423) );
  ANDN U5641 ( .A(n4848), .B(n4621), .Z(n4846) );
  XOR U5642 ( .A(n4849), .B(n4427), .Z(o[1150]) );
  XNOR U5643 ( .A(n4850), .B(round_reg[955]), .Z(n4427) );
  ANDN U5644 ( .A(n4851), .B(n4623), .Z(n4849) );
  XOR U5645 ( .A(n4852), .B(n3486), .Z(o[114]) );
  XOR U5646 ( .A(n2275), .B(round_reg[585]), .Z(n3486) );
  IV U5647 ( .A(n4853), .Z(n2275) );
  ANDN U5648 ( .A(n2896), .B(n2897), .Z(n4852) );
  XNOR U5649 ( .A(n2140), .B(round_reg[1460]), .Z(n2897) );
  XNOR U5650 ( .A(n2181), .B(round_reg[240]), .Z(n2896) );
  XOR U5651 ( .A(n4854), .B(n4431), .Z(o[1149]) );
  XOR U5652 ( .A(n2339), .B(round_reg[954]), .Z(n4431) );
  XOR U5653 ( .A(n4855), .B(n4856), .Z(n2339) );
  ANDN U5654 ( .A(n4857), .B(n4625), .Z(n4854) );
  XOR U5655 ( .A(n4858), .B(n4435), .Z(o[1148]) );
  XOR U5656 ( .A(n2343), .B(round_reg[953]), .Z(n4435) );
  XOR U5657 ( .A(n4859), .B(n4860), .Z(n2343) );
  ANDN U5658 ( .A(n4861), .B(n4627), .Z(n4858) );
  XOR U5659 ( .A(n4862), .B(n4439), .Z(o[1147]) );
  XOR U5660 ( .A(n2347), .B(round_reg[952]), .Z(n4439) );
  XOR U5661 ( .A(n4863), .B(n4864), .Z(n2347) );
  ANDN U5662 ( .A(n4865), .B(n4629), .Z(n4862) );
  XOR U5663 ( .A(n4866), .B(n4443), .Z(o[1146]) );
  XOR U5664 ( .A(n2355), .B(round_reg[951]), .Z(n4443) );
  XOR U5665 ( .A(n4867), .B(n4868), .Z(n2355) );
  ANDN U5666 ( .A(n4869), .B(n4631), .Z(n4866) );
  XOR U5667 ( .A(n4870), .B(n4447), .Z(o[1145]) );
  XOR U5668 ( .A(n2359), .B(round_reg[950]), .Z(n4447) );
  XNOR U5669 ( .A(n4871), .B(n4872), .Z(n2359) );
  ANDN U5670 ( .A(n4873), .B(n4635), .Z(n4870) );
  XOR U5671 ( .A(n4874), .B(n4451), .Z(o[1144]) );
  XNOR U5672 ( .A(n4318), .B(round_reg[949]), .Z(n4451) );
  XOR U5673 ( .A(n4875), .B(n4876), .Z(n4318) );
  ANDN U5674 ( .A(n4877), .B(n4637), .Z(n4874) );
  XOR U5675 ( .A(n4878), .B(n4455), .Z(o[1143]) );
  XNOR U5676 ( .A(n4321), .B(round_reg[948]), .Z(n4455) );
  XOR U5677 ( .A(n4879), .B(n4880), .Z(n4321) );
  ANDN U5678 ( .A(n4881), .B(n4639), .Z(n4878) );
  XOR U5679 ( .A(n4882), .B(n4459), .Z(o[1142]) );
  XNOR U5680 ( .A(n4324), .B(round_reg[947]), .Z(n4459) );
  XOR U5681 ( .A(n4883), .B(n4884), .Z(n4324) );
  ANDN U5682 ( .A(n4885), .B(n4641), .Z(n4882) );
  XOR U5683 ( .A(n4886), .B(n4465), .Z(o[1141]) );
  XNOR U5684 ( .A(n4327), .B(round_reg[946]), .Z(n4465) );
  XOR U5685 ( .A(n4887), .B(n4888), .Z(n4327) );
  ANDN U5686 ( .A(n4889), .B(n4643), .Z(n4886) );
  XOR U5687 ( .A(n4890), .B(n4469), .Z(o[1140]) );
  XNOR U5688 ( .A(n4332), .B(round_reg[945]), .Z(n4469) );
  XOR U5689 ( .A(n4891), .B(n4892), .Z(n4332) );
  ANDN U5690 ( .A(n4893), .B(n4645), .Z(n4890) );
  XOR U5691 ( .A(n4894), .B(n3488), .Z(o[113]) );
  XOR U5692 ( .A(n2279), .B(round_reg[584]), .Z(n3488) );
  IV U5693 ( .A(n4895), .Z(n2279) );
  ANDN U5694 ( .A(n2923), .B(n2924), .Z(n4894) );
  XNOR U5695 ( .A(n2144), .B(round_reg[1459]), .Z(n2924) );
  XNOR U5696 ( .A(n2185), .B(round_reg[239]), .Z(n2923) );
  XOR U5697 ( .A(n4896), .B(n4473), .Z(o[1139]) );
  XNOR U5698 ( .A(n4335), .B(round_reg[944]), .Z(n4473) );
  XOR U5699 ( .A(n4897), .B(n4898), .Z(n4335) );
  ANDN U5700 ( .A(n4899), .B(n4647), .Z(n4896) );
  XOR U5701 ( .A(n4900), .B(n4477), .Z(o[1138]) );
  XNOR U5702 ( .A(n4337), .B(round_reg[943]), .Z(n4477) );
  XOR U5703 ( .A(n4901), .B(n4902), .Z(n4337) );
  ANDN U5704 ( .A(n4903), .B(n4649), .Z(n4900) );
  XOR U5705 ( .A(n4904), .B(n4481), .Z(o[1137]) );
  XNOR U5706 ( .A(n4339), .B(round_reg[942]), .Z(n4481) );
  XOR U5707 ( .A(n4905), .B(n4906), .Z(n4339) );
  ANDN U5708 ( .A(n4907), .B(n4651), .Z(n4904) );
  XOR U5709 ( .A(n4908), .B(n4485), .Z(o[1136]) );
  XNOR U5710 ( .A(n3993), .B(round_reg[941]), .Z(n4485) );
  XOR U5711 ( .A(n4909), .B(n4910), .Z(n3993) );
  ANDN U5712 ( .A(n4911), .B(n4653), .Z(n4908) );
  XOR U5713 ( .A(n4912), .B(n4489), .Z(o[1135]) );
  XNOR U5714 ( .A(n4020), .B(round_reg[940]), .Z(n4489) );
  XOR U5715 ( .A(n4913), .B(n4914), .Z(n4020) );
  ANDN U5716 ( .A(n4915), .B(n4659), .Z(n4912) );
  XOR U5717 ( .A(n4916), .B(n4493), .Z(o[1134]) );
  XNOR U5718 ( .A(n4343), .B(round_reg[939]), .Z(n4493) );
  XOR U5719 ( .A(n4917), .B(n4918), .Z(n4343) );
  ANDN U5720 ( .A(n4919), .B(n4661), .Z(n4916) );
  XOR U5721 ( .A(n4920), .B(n4497), .Z(o[1133]) );
  XNOR U5722 ( .A(n4345), .B(round_reg[938]), .Z(n4497) );
  XOR U5723 ( .A(n4921), .B(n4922), .Z(n4345) );
  ANDN U5724 ( .A(n4923), .B(n4663), .Z(n4920) );
  XOR U5725 ( .A(n4924), .B(n4501), .Z(o[1132]) );
  XNOR U5726 ( .A(n4347), .B(round_reg[937]), .Z(n4501) );
  XOR U5727 ( .A(n4925), .B(n4926), .Z(n4347) );
  ANDN U5728 ( .A(n4927), .B(n4665), .Z(n4924) );
  XOR U5729 ( .A(n4928), .B(n4507), .Z(o[1131]) );
  XNOR U5730 ( .A(n4349), .B(round_reg[936]), .Z(n4507) );
  XOR U5731 ( .A(n4929), .B(n4930), .Z(n4349) );
  ANDN U5732 ( .A(n4931), .B(n4667), .Z(n4928) );
  XOR U5733 ( .A(n4932), .B(n4511), .Z(o[1130]) );
  XNOR U5734 ( .A(n4353), .B(round_reg[935]), .Z(n4511) );
  XOR U5735 ( .A(n4933), .B(n4934), .Z(n4353) );
  ANDN U5736 ( .A(n4935), .B(n4669), .Z(n4932) );
  XOR U5737 ( .A(n4936), .B(n3490), .Z(o[112]) );
  XOR U5738 ( .A(n2283), .B(round_reg[583]), .Z(n3490) );
  IV U5739 ( .A(n4937), .Z(n2283) );
  ANDN U5740 ( .A(n2947), .B(n2949), .Z(n4936) );
  XNOR U5741 ( .A(n2148), .B(round_reg[1458]), .Z(n2949) );
  XNOR U5742 ( .A(n2189), .B(round_reg[238]), .Z(n2947) );
  XOR U5743 ( .A(n4938), .B(n4515), .Z(o[1129]) );
  XNOR U5744 ( .A(n4356), .B(round_reg[934]), .Z(n4515) );
  XOR U5745 ( .A(n4939), .B(n4940), .Z(n4356) );
  ANDN U5746 ( .A(n4941), .B(n4671), .Z(n4938) );
  XOR U5747 ( .A(n4942), .B(n4519), .Z(o[1128]) );
  XNOR U5748 ( .A(n4359), .B(round_reg[933]), .Z(n4519) );
  XOR U5749 ( .A(n4943), .B(n4944), .Z(n4359) );
  ANDN U5750 ( .A(n4945), .B(n4673), .Z(n4942) );
  XOR U5751 ( .A(n4946), .B(n4522), .Z(o[1127]) );
  XNOR U5752 ( .A(n4362), .B(round_reg[932]), .Z(n4522) );
  XOR U5753 ( .A(n4947), .B(n4948), .Z(n4362) );
  ANDN U5754 ( .A(n1060), .B(n4677), .Z(n4946) );
  XOR U5755 ( .A(n4949), .B(n4524), .Z(o[1126]) );
  XNOR U5756 ( .A(n4365), .B(round_reg[931]), .Z(n4524) );
  XOR U5757 ( .A(n4950), .B(n4951), .Z(n4365) );
  ANDN U5758 ( .A(n1064), .B(n4681), .Z(n4949) );
  XOR U5759 ( .A(n4952), .B(n4526), .Z(o[1125]) );
  XNOR U5760 ( .A(n4368), .B(round_reg[930]), .Z(n4526) );
  XOR U5761 ( .A(n4953), .B(n4954), .Z(n4368) );
  ANDN U5762 ( .A(n1068), .B(n4688), .Z(n4952) );
  XOR U5763 ( .A(n4955), .B(n4528), .Z(o[1124]) );
  XNOR U5764 ( .A(n4370), .B(round_reg[929]), .Z(n4528) );
  XOR U5765 ( .A(n4956), .B(n4957), .Z(n4370) );
  ANDN U5766 ( .A(n1072), .B(n4692), .Z(n4955) );
  XOR U5767 ( .A(n4958), .B(n4530), .Z(o[1123]) );
  XNOR U5768 ( .A(n4372), .B(round_reg[928]), .Z(n4530) );
  XOR U5769 ( .A(n4959), .B(n4960), .Z(n4372) );
  ANDN U5770 ( .A(n1076), .B(n4696), .Z(n4958) );
  XOR U5771 ( .A(n4961), .B(n4532), .Z(o[1122]) );
  XOR U5772 ( .A(n2179), .B(round_reg[927]), .Z(n4532) );
  XNOR U5773 ( .A(n4962), .B(n4963), .Z(n2179) );
  ANDN U5774 ( .A(n1080), .B(n4700), .Z(n4961) );
  XOR U5775 ( .A(n4964), .B(n4536), .Z(o[1121]) );
  XOR U5776 ( .A(n2183), .B(round_reg[926]), .Z(n4536) );
  XNOR U5777 ( .A(n4965), .B(n4966), .Z(n2183) );
  ANDN U5778 ( .A(n1084), .B(n4704), .Z(n4964) );
  XOR U5779 ( .A(n4967), .B(n4538), .Z(o[1120]) );
  XOR U5780 ( .A(n2187), .B(round_reg[925]), .Z(n4538) );
  XNOR U5781 ( .A(n4968), .B(n4969), .Z(n2187) );
  ANDN U5782 ( .A(n1088), .B(n4708), .Z(n4967) );
  XOR U5783 ( .A(n4970), .B(n3493), .Z(o[111]) );
  XOR U5784 ( .A(n2287), .B(round_reg[582]), .Z(n3493) );
  IV U5785 ( .A(n4971), .Z(n2287) );
  ANDN U5786 ( .A(n2971), .B(n2973), .Z(n4970) );
  XNOR U5787 ( .A(n2152), .B(round_reg[1457]), .Z(n2973) );
  XNOR U5788 ( .A(n2193), .B(round_reg[237]), .Z(n2971) );
  XOR U5789 ( .A(n4972), .B(n4540), .Z(o[1119]) );
  XOR U5790 ( .A(n2191), .B(round_reg[924]), .Z(n4540) );
  XNOR U5791 ( .A(n4973), .B(n4974), .Z(n2191) );
  ANDN U5792 ( .A(n1092), .B(n4712), .Z(n4972) );
  XOR U5793 ( .A(n4975), .B(n4542), .Z(o[1118]) );
  XOR U5794 ( .A(n2195), .B(round_reg[923]), .Z(n4542) );
  XNOR U5795 ( .A(n4976), .B(n4977), .Z(n2195) );
  ANDN U5796 ( .A(n1096), .B(n4716), .Z(n4975) );
  XOR U5797 ( .A(n4978), .B(n4544), .Z(o[1117]) );
  XOR U5798 ( .A(n2199), .B(round_reg[922]), .Z(n4544) );
  XNOR U5799 ( .A(n4979), .B(n4980), .Z(n2199) );
  NOR U5800 ( .A(n1104), .B(n4720), .Z(n4978) );
  XOR U5801 ( .A(n4981), .B(n4546), .Z(o[1116]) );
  XNOR U5802 ( .A(n4382), .B(round_reg[921]), .Z(n4546) );
  XOR U5803 ( .A(n4982), .B(n4983), .Z(n4382) );
  NOR U5804 ( .A(n1108), .B(n4724), .Z(n4981) );
  XOR U5805 ( .A(n4984), .B(n4548), .Z(o[1115]) );
  XNOR U5806 ( .A(n4391), .B(round_reg[920]), .Z(n4548) );
  XOR U5807 ( .A(n4985), .B(n4986), .Z(n4391) );
  ANDN U5808 ( .A(n1112), .B(n4731), .Z(n4984) );
  XOR U5809 ( .A(n4987), .B(n4550), .Z(o[1114]) );
  XNOR U5810 ( .A(n4404), .B(round_reg[919]), .Z(n4550) );
  XOR U5811 ( .A(n4988), .B(n4989), .Z(n4404) );
  ANDN U5812 ( .A(n1116), .B(n4735), .Z(n4987) );
  XOR U5813 ( .A(n4990), .B(n4552), .Z(o[1113]) );
  XNOR U5814 ( .A(n4420), .B(round_reg[918]), .Z(n4552) );
  XOR U5815 ( .A(n4991), .B(n4992), .Z(n4420) );
  ANDN U5816 ( .A(n1120), .B(n4739), .Z(n4990) );
  XOR U5817 ( .A(n4993), .B(n4554), .Z(o[1112]) );
  XNOR U5818 ( .A(n4462), .B(round_reg[917]), .Z(n4554) );
  XOR U5819 ( .A(n4994), .B(n4995), .Z(n4462) );
  ANDN U5820 ( .A(n1124), .B(n4743), .Z(n4993) );
  XOR U5821 ( .A(n4996), .B(n4558), .Z(o[1111]) );
  XNOR U5822 ( .A(n4504), .B(round_reg[916]), .Z(n4558) );
  XOR U5823 ( .A(n4997), .B(n4998), .Z(n4504) );
  ANDN U5824 ( .A(n1128), .B(n4747), .Z(n4996) );
  XOR U5825 ( .A(n4999), .B(n4560), .Z(o[1110]) );
  XNOR U5826 ( .A(n4534), .B(round_reg[915]), .Z(n4560) );
  XOR U5827 ( .A(n5000), .B(n5001), .Z(n4534) );
  ANDN U5828 ( .A(n1132), .B(n4751), .Z(n4999) );
  XOR U5829 ( .A(n5002), .B(n3495), .Z(o[110]) );
  IV U5830 ( .A(n3580), .Z(n3495) );
  XNOR U5831 ( .A(n2291), .B(round_reg[581]), .Z(n3580) );
  ANDN U5832 ( .A(n2995), .B(n2997), .Z(n5002) );
  XNOR U5833 ( .A(n2156), .B(round_reg[1456]), .Z(n2997) );
  XNOR U5834 ( .A(n2197), .B(round_reg[236]), .Z(n2995) );
  XOR U5835 ( .A(n5003), .B(n4562), .Z(o[1109]) );
  XNOR U5836 ( .A(n4556), .B(round_reg[914]), .Z(n4562) );
  XOR U5837 ( .A(n5004), .B(n5005), .Z(n4556) );
  ANDN U5838 ( .A(n1136), .B(n4755), .Z(n5003) );
  XOR U5839 ( .A(n5006), .B(n4564), .Z(o[1108]) );
  XNOR U5840 ( .A(n4579), .B(round_reg[913]), .Z(n4564) );
  XOR U5841 ( .A(n5007), .B(n5008), .Z(n4579) );
  ANDN U5842 ( .A(n1140), .B(n4759), .Z(n5006) );
  XOR U5843 ( .A(n5009), .B(n4566), .Z(o[1107]) );
  XNOR U5844 ( .A(n4607), .B(round_reg[912]), .Z(n4566) );
  XOR U5845 ( .A(n5010), .B(n5011), .Z(n4607) );
  ANDN U5846 ( .A(n1148), .B(n4763), .Z(n5009) );
  XOR U5847 ( .A(n5012), .B(n4569), .Z(o[1106]) );
  XNOR U5848 ( .A(n4633), .B(round_reg[911]), .Z(n4569) );
  XOR U5849 ( .A(n5013), .B(n5014), .Z(n4633) );
  ANDN U5850 ( .A(n1152), .B(n4767), .Z(n5012) );
  XOR U5851 ( .A(n5015), .B(n4571), .Z(o[1105]) );
  XNOR U5852 ( .A(n4656), .B(round_reg[910]), .Z(n4571) );
  XOR U5853 ( .A(n5016), .B(n5017), .Z(n4656) );
  ANDN U5854 ( .A(n1156), .B(n4774), .Z(n5015) );
  XOR U5855 ( .A(n5018), .B(n4573), .Z(o[1104]) );
  XNOR U5856 ( .A(n4683), .B(round_reg[909]), .Z(n4573) );
  XOR U5857 ( .A(n5019), .B(n5020), .Z(n4683) );
  ANDN U5858 ( .A(n1160), .B(n4778), .Z(n5018) );
  XOR U5859 ( .A(n5021), .B(n4575), .Z(o[1103]) );
  XNOR U5860 ( .A(n4726), .B(round_reg[908]), .Z(n4575) );
  XOR U5861 ( .A(n5022), .B(n5023), .Z(n4726) );
  NOR U5862 ( .A(n1164), .B(n4782), .Z(n5021) );
  XOR U5863 ( .A(n5024), .B(n4577), .Z(o[1102]) );
  XNOR U5864 ( .A(n4769), .B(round_reg[907]), .Z(n4577) );
  XOR U5865 ( .A(n5025), .B(n5026), .Z(n4769) );
  ANDN U5866 ( .A(n1168), .B(n4786), .Z(n5024) );
  XOR U5867 ( .A(n5027), .B(n4581), .Z(o[1101]) );
  XNOR U5868 ( .A(n4812), .B(round_reg[906]), .Z(n4581) );
  XOR U5869 ( .A(n5028), .B(n5029), .Z(n4812) );
  ANDN U5870 ( .A(n1172), .B(n4790), .Z(n5027) );
  XOR U5871 ( .A(n5030), .B(n4583), .Z(o[1100]) );
  XNOR U5872 ( .A(n4853), .B(round_reg[905]), .Z(n4583) );
  XOR U5873 ( .A(n5031), .B(n5032), .Z(n4853) );
  ANDN U5874 ( .A(n1176), .B(n4794), .Z(n5030) );
  XOR U5875 ( .A(n5033), .B(n1987), .Z(o[10]) );
  XOR U5876 ( .A(n2357), .B(round_reg[200]), .Z(n1987) );
  ANDN U5877 ( .A(n1986), .B(n3429), .Z(n5033) );
  XOR U5878 ( .A(n1775), .B(round_reg[1043]), .Z(n3429) );
  XNOR U5879 ( .A(n2316), .B(round_reg[1420]), .Z(n1986) );
  XOR U5880 ( .A(n5034), .B(n3497), .Z(o[109]) );
  XOR U5881 ( .A(n2295), .B(round_reg[580]), .Z(n3497) );
  IV U5882 ( .A(n5035), .Z(n2295) );
  ANDN U5883 ( .A(n3019), .B(n3021), .Z(n5034) );
  XNOR U5884 ( .A(n2160), .B(round_reg[1455]), .Z(n3021) );
  XNOR U5885 ( .A(n2201), .B(round_reg[235]), .Z(n3019) );
  XOR U5886 ( .A(n5036), .B(n4586), .Z(o[1099]) );
  XNOR U5887 ( .A(n4895), .B(round_reg[904]), .Z(n4586) );
  XOR U5888 ( .A(n5037), .B(n5038), .Z(n4895) );
  ANDN U5889 ( .A(n1180), .B(n4798), .Z(n5036) );
  XOR U5890 ( .A(n5039), .B(n4589), .Z(o[1098]) );
  XNOR U5891 ( .A(n4937), .B(round_reg[903]), .Z(n4589) );
  XOR U5892 ( .A(n5040), .B(n5041), .Z(n4937) );
  ANDN U5893 ( .A(n1184), .B(n4802), .Z(n5039) );
  XOR U5894 ( .A(n5042), .B(n4592), .Z(o[1097]) );
  XNOR U5895 ( .A(n4971), .B(round_reg[902]), .Z(n4592) );
  XOR U5896 ( .A(n5043), .B(n5044), .Z(n4971) );
  ANDN U5897 ( .A(n1192), .B(n4806), .Z(n5042) );
  XOR U5898 ( .A(n5045), .B(n4595), .Z(o[1096]) );
  XOR U5899 ( .A(n2291), .B(round_reg[901]), .Z(n4595) );
  XNOR U5900 ( .A(n5046), .B(n5047), .Z(n2291) );
  NOR U5901 ( .A(n1196), .B(n4810), .Z(n5045) );
  XOR U5902 ( .A(n5048), .B(n4597), .Z(o[1095]) );
  XNOR U5903 ( .A(n5035), .B(round_reg[900]), .Z(n4597) );
  XOR U5904 ( .A(n5049), .B(n5050), .Z(n5035) );
  NOR U5905 ( .A(n1200), .B(n4817), .Z(n5048) );
  XOR U5906 ( .A(n5051), .B(n4599), .Z(o[1094]) );
  XNOR U5907 ( .A(n5052), .B(round_reg[899]), .Z(n4599) );
  NOR U5908 ( .A(n1204), .B(n4821), .Z(n5051) );
  XOR U5909 ( .A(n5053), .B(n4601), .Z(o[1093]) );
  XNOR U5910 ( .A(n5054), .B(round_reg[898]), .Z(n4601) );
  NOR U5911 ( .A(n1208), .B(n4825), .Z(n5053) );
  XOR U5912 ( .A(n5055), .B(n4604), .Z(o[1092]) );
  XNOR U5913 ( .A(n5056), .B(round_reg[897]), .Z(n4604) );
  NOR U5914 ( .A(n1212), .B(n4829), .Z(n5055) );
  XOR U5915 ( .A(n5057), .B(n4609), .Z(o[1091]) );
  XNOR U5916 ( .A(n5058), .B(round_reg[896]), .Z(n4609) );
  NOR U5917 ( .A(n1216), .B(n4833), .Z(n5057) );
  XOR U5918 ( .A(n5059), .B(n4612), .Z(o[1090]) );
  XNOR U5919 ( .A(n5060), .B(round_reg[959]), .Z(n4612) );
  NOR U5920 ( .A(n1220), .B(n4837), .Z(n5059) );
  XOR U5921 ( .A(n5061), .B(n3499), .Z(o[108]) );
  XOR U5922 ( .A(n2299), .B(round_reg[579]), .Z(n3499) );
  IV U5923 ( .A(n5052), .Z(n2299) );
  XOR U5924 ( .A(n5062), .B(n5063), .Z(n5052) );
  ANDN U5925 ( .A(n3044), .B(n3046), .Z(n5061) );
  XNOR U5926 ( .A(n2164), .B(round_reg[1454]), .Z(n3046) );
  XNOR U5927 ( .A(n2205), .B(round_reg[234]), .Z(n3044) );
  XOR U5928 ( .A(n5064), .B(n4615), .Z(o[1089]) );
  XNOR U5929 ( .A(n5065), .B(round_reg[958]), .Z(n4615) );
  NOR U5930 ( .A(n1224), .B(n4841), .Z(n5064) );
  XOR U5931 ( .A(n5066), .B(n4618), .Z(o[1088]) );
  XNOR U5932 ( .A(n5067), .B(round_reg[957]), .Z(n4618) );
  NOR U5933 ( .A(n1228), .B(n4845), .Z(n5066) );
  XOR U5934 ( .A(n5068), .B(n4621), .Z(o[1087]) );
  XOR U5935 ( .A(n2313), .B(round_reg[530]), .Z(n4621) );
  XNOR U5936 ( .A(n5069), .B(n4675), .Z(n2313) );
  XOR U5937 ( .A(n5070), .B(n5071), .Z(n4675) );
  XOR U5938 ( .A(round_reg[274]), .B(n5072), .Z(n5071) );
  XOR U5939 ( .A(round_reg[914]), .B(round_reg[594]), .Z(n5072) );
  XNOR U5940 ( .A(round_reg[1234]), .B(round_reg[1554]), .Z(n5070) );
  ANDN U5941 ( .A(n4422), .B(n4848), .Z(n5068) );
  XOR U5942 ( .A(n5073), .B(n4623), .Z(o[1086]) );
  XOR U5943 ( .A(n2317), .B(round_reg[529]), .Z(n4623) );
  XNOR U5944 ( .A(n5074), .B(n4679), .Z(n2317) );
  XOR U5945 ( .A(n5075), .B(n5076), .Z(n4679) );
  XOR U5946 ( .A(round_reg[273]), .B(n5077), .Z(n5076) );
  XOR U5947 ( .A(round_reg[913]), .B(round_reg[593]), .Z(n5077) );
  XNOR U5948 ( .A(round_reg[1233]), .B(round_reg[1553]), .Z(n5075) );
  ANDN U5949 ( .A(n4426), .B(n4851), .Z(n5073) );
  XOR U5950 ( .A(n5078), .B(n4625), .Z(o[1085]) );
  XOR U5951 ( .A(n2321), .B(round_reg[528]), .Z(n4625) );
  XNOR U5952 ( .A(n5079), .B(n4686), .Z(n2321) );
  XOR U5953 ( .A(n5080), .B(n5081), .Z(n4686) );
  XOR U5954 ( .A(round_reg[272]), .B(n5082), .Z(n5081) );
  XOR U5955 ( .A(round_reg[912]), .B(round_reg[592]), .Z(n5082) );
  XNOR U5956 ( .A(round_reg[1232]), .B(round_reg[1552]), .Z(n5080) );
  ANDN U5957 ( .A(n4430), .B(n4857), .Z(n5078) );
  XOR U5958 ( .A(n5083), .B(n4627), .Z(o[1084]) );
  XOR U5959 ( .A(n2325), .B(round_reg[527]), .Z(n4627) );
  XNOR U5960 ( .A(n5084), .B(n4690), .Z(n2325) );
  XOR U5961 ( .A(n5085), .B(n5086), .Z(n4690) );
  XOR U5962 ( .A(round_reg[271]), .B(n5087), .Z(n5086) );
  XOR U5963 ( .A(round_reg[911]), .B(round_reg[591]), .Z(n5087) );
  XNOR U5964 ( .A(round_reg[1231]), .B(round_reg[1551]), .Z(n5085) );
  ANDN U5965 ( .A(n4434), .B(n4861), .Z(n5083) );
  XOR U5966 ( .A(n5088), .B(n4629), .Z(o[1083]) );
  XOR U5967 ( .A(n2329), .B(round_reg[526]), .Z(n4629) );
  XNOR U5968 ( .A(n5089), .B(n4694), .Z(n2329) );
  XOR U5969 ( .A(n5090), .B(n5091), .Z(n4694) );
  XOR U5970 ( .A(round_reg[270]), .B(n5092), .Z(n5091) );
  XOR U5971 ( .A(round_reg[910]), .B(round_reg[590]), .Z(n5092) );
  XNOR U5972 ( .A(round_reg[1230]), .B(round_reg[1550]), .Z(n5090) );
  ANDN U5973 ( .A(n4438), .B(n4865), .Z(n5088) );
  XOR U5974 ( .A(n5093), .B(n4631), .Z(o[1082]) );
  XOR U5975 ( .A(n2333), .B(round_reg[525]), .Z(n4631) );
  XNOR U5976 ( .A(n5094), .B(n4698), .Z(n2333) );
  XOR U5977 ( .A(n5095), .B(n5096), .Z(n4698) );
  XOR U5978 ( .A(round_reg[269]), .B(n5097), .Z(n5096) );
  XOR U5979 ( .A(round_reg[909]), .B(round_reg[589]), .Z(n5097) );
  XNOR U5980 ( .A(round_reg[1229]), .B(round_reg[1549]), .Z(n5095) );
  ANDN U5981 ( .A(n4442), .B(n4869), .Z(n5093) );
  XOR U5982 ( .A(n5098), .B(n4635), .Z(o[1081]) );
  XOR U5983 ( .A(n2337), .B(round_reg[524]), .Z(n4635) );
  XNOR U5984 ( .A(n4702), .B(n5099), .Z(n2337) );
  XNOR U5985 ( .A(n5100), .B(n5101), .Z(n4702) );
  XOR U5986 ( .A(round_reg[268]), .B(n5102), .Z(n5101) );
  XOR U5987 ( .A(round_reg[908]), .B(round_reg[588]), .Z(n5102) );
  XNOR U5988 ( .A(round_reg[1228]), .B(round_reg[1548]), .Z(n5100) );
  ANDN U5989 ( .A(n4446), .B(n4873), .Z(n5098) );
  XOR U5990 ( .A(n5103), .B(n4637), .Z(o[1080]) );
  XOR U5991 ( .A(n2341), .B(round_reg[523]), .Z(n4637) );
  XNOR U5992 ( .A(n4706), .B(n5104), .Z(n2341) );
  XNOR U5993 ( .A(n5105), .B(n5106), .Z(n4706) );
  XOR U5994 ( .A(round_reg[267]), .B(n5107), .Z(n5106) );
  XOR U5995 ( .A(round_reg[907]), .B(round_reg[587]), .Z(n5107) );
  XNOR U5996 ( .A(round_reg[1227]), .B(round_reg[1547]), .Z(n5105) );
  ANDN U5997 ( .A(n4450), .B(n4877), .Z(n5103) );
  XOR U5998 ( .A(n5108), .B(n3501), .Z(o[107]) );
  XOR U5999 ( .A(n2303), .B(round_reg[578]), .Z(n3501) );
  IV U6000 ( .A(n5054), .Z(n2303) );
  XOR U6001 ( .A(n5109), .B(n5110), .Z(n5054) );
  ANDN U6002 ( .A(n3060), .B(n3062), .Z(n5108) );
  XNOR U6003 ( .A(n2168), .B(round_reg[1453]), .Z(n3062) );
  XNOR U6004 ( .A(n2209), .B(round_reg[233]), .Z(n3060) );
  XOR U6005 ( .A(n5111), .B(n4639), .Z(o[1079]) );
  XOR U6006 ( .A(n2345), .B(round_reg[522]), .Z(n4639) );
  XNOR U6007 ( .A(n4710), .B(n5112), .Z(n2345) );
  XNOR U6008 ( .A(n5113), .B(n5114), .Z(n4710) );
  XOR U6009 ( .A(round_reg[266]), .B(n5115), .Z(n5114) );
  XOR U6010 ( .A(round_reg[906]), .B(round_reg[586]), .Z(n5115) );
  XNOR U6011 ( .A(round_reg[1226]), .B(round_reg[1546]), .Z(n5113) );
  ANDN U6012 ( .A(n4454), .B(n4881), .Z(n5111) );
  XOR U6013 ( .A(n5116), .B(n4641), .Z(o[1078]) );
  XOR U6014 ( .A(n2349), .B(round_reg[521]), .Z(n4641) );
  XNOR U6015 ( .A(n4714), .B(n5117), .Z(n2349) );
  XNOR U6016 ( .A(n5118), .B(n5119), .Z(n4714) );
  XOR U6017 ( .A(round_reg[265]), .B(n5120), .Z(n5119) );
  XOR U6018 ( .A(round_reg[905]), .B(round_reg[585]), .Z(n5120) );
  XNOR U6019 ( .A(round_reg[1225]), .B(round_reg[1545]), .Z(n5118) );
  ANDN U6020 ( .A(n4458), .B(n4885), .Z(n5116) );
  XOR U6021 ( .A(n5121), .B(n4643), .Z(o[1077]) );
  XOR U6022 ( .A(n2357), .B(round_reg[520]), .Z(n4643) );
  XNOR U6023 ( .A(n4718), .B(n5122), .Z(n2357) );
  XNOR U6024 ( .A(n5123), .B(n5124), .Z(n4718) );
  XOR U6025 ( .A(round_reg[264]), .B(n5125), .Z(n5124) );
  XOR U6026 ( .A(round_reg[904]), .B(round_reg[584]), .Z(n5125) );
  XNOR U6027 ( .A(round_reg[1224]), .B(round_reg[1544]), .Z(n5123) );
  ANDN U6028 ( .A(n4464), .B(n4889), .Z(n5121) );
  XOR U6029 ( .A(n5126), .B(n4645), .Z(o[1076]) );
  XOR U6030 ( .A(n2361), .B(round_reg[519]), .Z(n4645) );
  XOR U6031 ( .A(n4723), .B(n5127), .Z(n2361) );
  XOR U6032 ( .A(n5128), .B(n5129), .Z(n4723) );
  XOR U6033 ( .A(round_reg[263]), .B(n5130), .Z(n5129) );
  XOR U6034 ( .A(round_reg[903]), .B(round_reg[583]), .Z(n5130) );
  XNOR U6035 ( .A(round_reg[1223]), .B(round_reg[1543]), .Z(n5128) );
  ANDN U6036 ( .A(n4468), .B(n4893), .Z(n5126) );
  XOR U6037 ( .A(n5131), .B(n4647), .Z(o[1075]) );
  XOR U6038 ( .A(n2365), .B(round_reg[518]), .Z(n4647) );
  XNOR U6039 ( .A(n4729), .B(n5132), .Z(n2365) );
  XNOR U6040 ( .A(n5133), .B(n5134), .Z(n4729) );
  XOR U6041 ( .A(round_reg[262]), .B(n5135), .Z(n5134) );
  XOR U6042 ( .A(round_reg[902]), .B(round_reg[582]), .Z(n5135) );
  XNOR U6043 ( .A(round_reg[1222]), .B(round_reg[1542]), .Z(n5133) );
  ANDN U6044 ( .A(n4472), .B(n4899), .Z(n5131) );
  XOR U6045 ( .A(n5136), .B(n4649), .Z(o[1074]) );
  XOR U6046 ( .A(n2369), .B(round_reg[517]), .Z(n4649) );
  XNOR U6047 ( .A(n4733), .B(n5137), .Z(n2369) );
  XNOR U6048 ( .A(n5138), .B(n5139), .Z(n4733) );
  XOR U6049 ( .A(round_reg[261]), .B(n5140), .Z(n5139) );
  XOR U6050 ( .A(round_reg[901]), .B(round_reg[581]), .Z(n5140) );
  XNOR U6051 ( .A(round_reg[1221]), .B(round_reg[1541]), .Z(n5138) );
  ANDN U6052 ( .A(n4476), .B(n4903), .Z(n5136) );
  XOR U6053 ( .A(n5141), .B(n4651), .Z(o[1073]) );
  XOR U6054 ( .A(n2373), .B(round_reg[516]), .Z(n4651) );
  XNOR U6055 ( .A(n4737), .B(n5142), .Z(n2373) );
  XNOR U6056 ( .A(n5143), .B(n5144), .Z(n4737) );
  XOR U6057 ( .A(round_reg[260]), .B(n5145), .Z(n5144) );
  XOR U6058 ( .A(round_reg[900]), .B(round_reg[580]), .Z(n5145) );
  XNOR U6059 ( .A(round_reg[1220]), .B(round_reg[1540]), .Z(n5143) );
  ANDN U6060 ( .A(n4480), .B(n4907), .Z(n5141) );
  XOR U6061 ( .A(n5146), .B(n4653), .Z(o[1072]) );
  XOR U6062 ( .A(n2377), .B(round_reg[515]), .Z(n4653) );
  XNOR U6063 ( .A(n4741), .B(n5147), .Z(n2377) );
  XNOR U6064 ( .A(n5148), .B(n5149), .Z(n4741) );
  XOR U6065 ( .A(round_reg[259]), .B(n5150), .Z(n5149) );
  XOR U6066 ( .A(round_reg[899]), .B(round_reg[579]), .Z(n5150) );
  XNOR U6067 ( .A(round_reg[1219]), .B(round_reg[1539]), .Z(n5148) );
  ANDN U6068 ( .A(n4484), .B(n4911), .Z(n5146) );
  XOR U6069 ( .A(n5151), .B(n4659), .Z(o[1071]) );
  XOR U6070 ( .A(n2381), .B(round_reg[514]), .Z(n4659) );
  XNOR U6071 ( .A(n4745), .B(n5152), .Z(n2381) );
  XNOR U6072 ( .A(n5153), .B(n5154), .Z(n4745) );
  XOR U6073 ( .A(round_reg[258]), .B(n5155), .Z(n5154) );
  XOR U6074 ( .A(round_reg[898]), .B(round_reg[578]), .Z(n5155) );
  XNOR U6075 ( .A(round_reg[1218]), .B(round_reg[1538]), .Z(n5153) );
  ANDN U6076 ( .A(n4488), .B(n4915), .Z(n5151) );
  XOR U6077 ( .A(n5156), .B(n4661), .Z(o[1070]) );
  XOR U6078 ( .A(n2385), .B(round_reg[513]), .Z(n4661) );
  XNOR U6079 ( .A(n4749), .B(n5157), .Z(n2385) );
  XNOR U6080 ( .A(n5158), .B(n5159), .Z(n4749) );
  XOR U6081 ( .A(round_reg[257]), .B(n5160), .Z(n5159) );
  XOR U6082 ( .A(round_reg[897]), .B(round_reg[577]), .Z(n5160) );
  XNOR U6083 ( .A(round_reg[1217]), .B(round_reg[1537]), .Z(n5158) );
  ANDN U6084 ( .A(n4492), .B(n4919), .Z(n5156) );
  XOR U6085 ( .A(n5161), .B(n3503), .Z(o[106]) );
  XOR U6086 ( .A(n2311), .B(round_reg[577]), .Z(n3503) );
  IV U6087 ( .A(n5056), .Z(n2311) );
  XOR U6088 ( .A(n5162), .B(n5163), .Z(n5056) );
  ANDN U6089 ( .A(n3080), .B(n3082), .Z(n5161) );
  XOR U6090 ( .A(n2172), .B(round_reg[1452]), .Z(n3082) );
  XNOR U6091 ( .A(n2213), .B(round_reg[232]), .Z(n3080) );
  XOR U6092 ( .A(n5164), .B(n4663), .Z(o[1069]) );
  XOR U6093 ( .A(n2389), .B(round_reg[512]), .Z(n4663) );
  XNOR U6094 ( .A(n4753), .B(n5165), .Z(n2389) );
  XNOR U6095 ( .A(n5166), .B(n5167), .Z(n4753) );
  XOR U6096 ( .A(round_reg[256]), .B(n5168), .Z(n5167) );
  XOR U6097 ( .A(round_reg[896]), .B(round_reg[576]), .Z(n5168) );
  XNOR U6098 ( .A(round_reg[1216]), .B(round_reg[1536]), .Z(n5166) );
  ANDN U6099 ( .A(n4496), .B(n4923), .Z(n5164) );
  XOR U6100 ( .A(n5169), .B(n4665), .Z(o[1068]) );
  XOR U6101 ( .A(n2393), .B(round_reg[575]), .Z(n4665) );
  XNOR U6102 ( .A(n4757), .B(n5170), .Z(n2393) );
  XNOR U6103 ( .A(n5171), .B(n5172), .Z(n4757) );
  XOR U6104 ( .A(round_reg[319]), .B(n5173), .Z(n5172) );
  XOR U6105 ( .A(round_reg[959]), .B(round_reg[639]), .Z(n5173) );
  XNOR U6106 ( .A(round_reg[1279]), .B(round_reg[1599]), .Z(n5171) );
  ANDN U6107 ( .A(n4500), .B(n4927), .Z(n5169) );
  XOR U6108 ( .A(n5174), .B(n4667), .Z(o[1067]) );
  XNOR U6109 ( .A(n2113), .B(round_reg[574]), .Z(n4667) );
  ANDN U6110 ( .A(n4506), .B(n4931), .Z(n5174) );
  XOR U6111 ( .A(n5175), .B(n4669), .Z(o[1066]) );
  XOR U6112 ( .A(n2117), .B(round_reg[573]), .Z(n4669) );
  XNOR U6113 ( .A(n4765), .B(n5176), .Z(n2117) );
  XNOR U6114 ( .A(n5177), .B(n5178), .Z(n4765) );
  XOR U6115 ( .A(round_reg[317]), .B(n5179), .Z(n5178) );
  XOR U6116 ( .A(round_reg[957]), .B(round_reg[637]), .Z(n5179) );
  XNOR U6117 ( .A(round_reg[1277]), .B(round_reg[1597]), .Z(n5177) );
  ANDN U6118 ( .A(n4510), .B(n4935), .Z(n5175) );
  XOR U6119 ( .A(n5180), .B(n4671), .Z(o[1065]) );
  XOR U6120 ( .A(n2121), .B(round_reg[572]), .Z(n4671) );
  XNOR U6121 ( .A(n4772), .B(n5181), .Z(n2121) );
  XNOR U6122 ( .A(n5182), .B(n5183), .Z(n4772) );
  XOR U6123 ( .A(round_reg[316]), .B(n5184), .Z(n5183) );
  XOR U6124 ( .A(round_reg[956]), .B(round_reg[636]), .Z(n5184) );
  XNOR U6125 ( .A(round_reg[1276]), .B(round_reg[1596]), .Z(n5182) );
  ANDN U6126 ( .A(n4514), .B(n4941), .Z(n5180) );
  XOR U6127 ( .A(n5185), .B(n4673), .Z(o[1064]) );
  XOR U6128 ( .A(n2125), .B(round_reg[571]), .Z(n4673) );
  XNOR U6129 ( .A(n4776), .B(n5186), .Z(n2125) );
  XNOR U6130 ( .A(n5187), .B(n5188), .Z(n4776) );
  XOR U6131 ( .A(round_reg[315]), .B(n5189), .Z(n5188) );
  XOR U6132 ( .A(round_reg[955]), .B(round_reg[635]), .Z(n5189) );
  XNOR U6133 ( .A(round_reg[1275]), .B(round_reg[1595]), .Z(n5187) );
  ANDN U6134 ( .A(n4518), .B(n4945), .Z(n5185) );
  XOR U6135 ( .A(n5190), .B(n4677), .Z(o[1063]) );
  XOR U6136 ( .A(n2136), .B(round_reg[570]), .Z(n4677) );
  XNOR U6137 ( .A(n4780), .B(n5191), .Z(n2136) );
  XNOR U6138 ( .A(n5192), .B(n5193), .Z(n4780) );
  XOR U6139 ( .A(round_reg[314]), .B(n5194), .Z(n5193) );
  XOR U6140 ( .A(round_reg[954]), .B(round_reg[634]), .Z(n5194) );
  XNOR U6141 ( .A(round_reg[1274]), .B(round_reg[1594]), .Z(n5192) );
  ANDN U6142 ( .A(n1062), .B(n1060), .Z(n5190) );
  XOR U6143 ( .A(n2184), .B(round_reg[170]), .Z(n1060) );
  XOR U6144 ( .A(n1803), .B(round_reg[1355]), .Z(n1062) );
  XOR U6145 ( .A(n5099), .B(n5029), .Z(n1803) );
  XOR U6146 ( .A(n5195), .B(n5196), .Z(n5029) );
  XOR U6147 ( .A(round_reg[330]), .B(n5197), .Z(n5196) );
  XOR U6148 ( .A(round_reg[970]), .B(round_reg[650]), .Z(n5197) );
  XNOR U6149 ( .A(round_reg[10]), .B(round_reg[1290]), .Z(n5195) );
  XOR U6150 ( .A(n5198), .B(n5199), .Z(n5099) );
  XOR U6151 ( .A(round_reg[1419]), .B(n5200), .Z(n5199) );
  XOR U6152 ( .A(round_reg[779]), .B(round_reg[459]), .Z(n5200) );
  XNOR U6153 ( .A(round_reg[1099]), .B(round_reg[139]), .Z(n5198) );
  XOR U6154 ( .A(n5201), .B(n4681), .Z(o[1062]) );
  XOR U6155 ( .A(n2141), .B(round_reg[569]), .Z(n4681) );
  XNOR U6156 ( .A(n4784), .B(n5202), .Z(n2141) );
  XNOR U6157 ( .A(n5203), .B(n5204), .Z(n4784) );
  XOR U6158 ( .A(round_reg[313]), .B(n5205), .Z(n5204) );
  XOR U6159 ( .A(round_reg[953]), .B(round_reg[633]), .Z(n5205) );
  XNOR U6160 ( .A(round_reg[1273]), .B(round_reg[1593]), .Z(n5203) );
  NOR U6161 ( .A(n1066), .B(n1064), .Z(n5201) );
  XOR U6162 ( .A(n2188), .B(round_reg[169]), .Z(n1064) );
  XNOR U6163 ( .A(n1806), .B(round_reg[1354]), .Z(n1066) );
  XOR U6164 ( .A(n5104), .B(n5032), .Z(n1806) );
  XOR U6165 ( .A(n5206), .B(n5207), .Z(n5032) );
  XOR U6166 ( .A(round_reg[649]), .B(n5208), .Z(n5207) );
  XOR U6167 ( .A(round_reg[9]), .B(round_reg[969]), .Z(n5208) );
  XNOR U6168 ( .A(round_reg[1289]), .B(round_reg[329]), .Z(n5206) );
  XOR U6169 ( .A(n5209), .B(n5210), .Z(n5104) );
  XOR U6170 ( .A(round_reg[1418]), .B(n5211), .Z(n5210) );
  XOR U6171 ( .A(round_reg[778]), .B(round_reg[458]), .Z(n5211) );
  XNOR U6172 ( .A(round_reg[1098]), .B(round_reg[138]), .Z(n5209) );
  XOR U6173 ( .A(n5212), .B(n4688), .Z(o[1061]) );
  XOR U6174 ( .A(n2145), .B(round_reg[568]), .Z(n4688) );
  XNOR U6175 ( .A(n4788), .B(n5213), .Z(n2145) );
  XNOR U6176 ( .A(n5214), .B(n5215), .Z(n4788) );
  XOR U6177 ( .A(round_reg[312]), .B(n5216), .Z(n5215) );
  XOR U6178 ( .A(round_reg[952]), .B(round_reg[632]), .Z(n5216) );
  XNOR U6179 ( .A(round_reg[1272]), .B(round_reg[1592]), .Z(n5214) );
  ANDN U6180 ( .A(n1070), .B(n1068), .Z(n5212) );
  XOR U6181 ( .A(n2192), .B(round_reg[168]), .Z(n1068) );
  XOR U6182 ( .A(n1809), .B(round_reg[1353]), .Z(n1070) );
  XOR U6183 ( .A(n5217), .B(n4692), .Z(o[1060]) );
  XOR U6184 ( .A(n2149), .B(round_reg[567]), .Z(n4692) );
  XNOR U6185 ( .A(n4792), .B(n5218), .Z(n2149) );
  XNOR U6186 ( .A(n5219), .B(n5220), .Z(n4792) );
  XOR U6187 ( .A(round_reg[311]), .B(n5221), .Z(n5220) );
  XOR U6188 ( .A(round_reg[951]), .B(round_reg[631]), .Z(n5221) );
  XNOR U6189 ( .A(round_reg[1271]), .B(round_reg[1591]), .Z(n5219) );
  ANDN U6190 ( .A(n1074), .B(n1072), .Z(n5217) );
  XOR U6191 ( .A(n2196), .B(round_reg[167]), .Z(n1072) );
  XOR U6192 ( .A(n1812), .B(round_reg[1352]), .Z(n1074) );
  XOR U6193 ( .A(n5117), .B(n5041), .Z(n1812) );
  XOR U6194 ( .A(n5222), .B(n5223), .Z(n5041) );
  XOR U6195 ( .A(round_reg[647]), .B(n5224), .Z(n5223) );
  XOR U6196 ( .A(round_reg[967]), .B(round_reg[7]), .Z(n5224) );
  XNOR U6197 ( .A(round_reg[1287]), .B(round_reg[327]), .Z(n5222) );
  XOR U6198 ( .A(n5225), .B(n5226), .Z(n5117) );
  XOR U6199 ( .A(round_reg[1416]), .B(n5227), .Z(n5226) );
  XOR U6200 ( .A(round_reg[776]), .B(round_reg[456]), .Z(n5227) );
  XNOR U6201 ( .A(round_reg[1096]), .B(round_reg[136]), .Z(n5225) );
  XOR U6202 ( .A(n5228), .B(n3505), .Z(o[105]) );
  XOR U6203 ( .A(n2315), .B(round_reg[576]), .Z(n3505) );
  IV U6204 ( .A(n5058), .Z(n2315) );
  XOR U6205 ( .A(n5229), .B(n5230), .Z(n5058) );
  ANDN U6206 ( .A(n3103), .B(n3105), .Z(n5228) );
  XOR U6207 ( .A(n2180), .B(round_reg[1451]), .Z(n3105) );
  XNOR U6208 ( .A(n2217), .B(round_reg[231]), .Z(n3103) );
  XOR U6209 ( .A(n5231), .B(n4696), .Z(o[1059]) );
  XOR U6210 ( .A(n2153), .B(round_reg[566]), .Z(n4696) );
  XNOR U6211 ( .A(n4796), .B(n5232), .Z(n2153) );
  XNOR U6212 ( .A(n5233), .B(n5234), .Z(n4796) );
  XOR U6213 ( .A(round_reg[310]), .B(n5235), .Z(n5234) );
  XOR U6214 ( .A(round_reg[950]), .B(round_reg[630]), .Z(n5235) );
  XNOR U6215 ( .A(round_reg[1270]), .B(round_reg[1590]), .Z(n5233) );
  ANDN U6216 ( .A(n1078), .B(n1076), .Z(n5231) );
  XOR U6217 ( .A(n2200), .B(round_reg[166]), .Z(n1076) );
  XOR U6218 ( .A(n1815), .B(round_reg[1351]), .Z(n1078) );
  XOR U6219 ( .A(n5122), .B(n5044), .Z(n1815) );
  XOR U6220 ( .A(n5236), .B(n5237), .Z(n5044) );
  XOR U6221 ( .A(round_reg[646]), .B(n5238), .Z(n5237) );
  XOR U6222 ( .A(round_reg[966]), .B(round_reg[6]), .Z(n5238) );
  XNOR U6223 ( .A(round_reg[1286]), .B(round_reg[326]), .Z(n5236) );
  XOR U6224 ( .A(n5239), .B(n5240), .Z(n5122) );
  XOR U6225 ( .A(round_reg[1415]), .B(n5241), .Z(n5240) );
  XOR U6226 ( .A(round_reg[775]), .B(round_reg[455]), .Z(n5241) );
  XNOR U6227 ( .A(round_reg[1095]), .B(round_reg[135]), .Z(n5239) );
  XOR U6228 ( .A(n5242), .B(n4700), .Z(o[1058]) );
  XOR U6229 ( .A(n2157), .B(round_reg[565]), .Z(n4700) );
  XNOR U6230 ( .A(n4800), .B(n5243), .Z(n2157) );
  XNOR U6231 ( .A(n5244), .B(n5245), .Z(n4800) );
  XOR U6232 ( .A(round_reg[309]), .B(n5246), .Z(n5245) );
  XOR U6233 ( .A(round_reg[949]), .B(round_reg[629]), .Z(n5246) );
  XNOR U6234 ( .A(round_reg[1269]), .B(round_reg[1589]), .Z(n5244) );
  ANDN U6235 ( .A(n1082), .B(n1080), .Z(n5242) );
  XOR U6236 ( .A(n2204), .B(round_reg[165]), .Z(n1080) );
  XOR U6237 ( .A(n4940), .B(n5247), .Z(n2204) );
  XOR U6238 ( .A(n5248), .B(n5249), .Z(n4940) );
  XOR U6239 ( .A(round_reg[229]), .B(n5250), .Z(n5249) );
  XOR U6240 ( .A(round_reg[869]), .B(round_reg[549]), .Z(n5250) );
  XNOR U6241 ( .A(round_reg[1189]), .B(round_reg[1509]), .Z(n5248) );
  XOR U6242 ( .A(n1826), .B(round_reg[1350]), .Z(n1082) );
  XOR U6243 ( .A(n5047), .B(n5127), .Z(n1826) );
  XOR U6244 ( .A(n5251), .B(n5252), .Z(n5127) );
  XOR U6245 ( .A(round_reg[1414]), .B(n5253), .Z(n5252) );
  XOR U6246 ( .A(round_reg[774]), .B(round_reg[454]), .Z(n5253) );
  XNOR U6247 ( .A(round_reg[1094]), .B(round_reg[134]), .Z(n5251) );
  XOR U6248 ( .A(n5254), .B(n5255), .Z(n5047) );
  XOR U6249 ( .A(round_reg[5]), .B(n5256), .Z(n5255) );
  XOR U6250 ( .A(round_reg[965]), .B(round_reg[645]), .Z(n5256) );
  XNOR U6251 ( .A(round_reg[1285]), .B(round_reg[325]), .Z(n5254) );
  XOR U6252 ( .A(n5257), .B(n4704), .Z(o[1057]) );
  XOR U6253 ( .A(n2161), .B(round_reg[564]), .Z(n4704) );
  XNOR U6254 ( .A(n4804), .B(n5258), .Z(n2161) );
  XNOR U6255 ( .A(n5259), .B(n5260), .Z(n4804) );
  XOR U6256 ( .A(round_reg[308]), .B(n5261), .Z(n5260) );
  XOR U6257 ( .A(round_reg[948]), .B(round_reg[628]), .Z(n5261) );
  XNOR U6258 ( .A(round_reg[1268]), .B(round_reg[1588]), .Z(n5259) );
  ANDN U6259 ( .A(n1086), .B(n1084), .Z(n5257) );
  XOR U6260 ( .A(n2208), .B(round_reg[164]), .Z(n1084) );
  XOR U6261 ( .A(n4944), .B(n5262), .Z(n2208) );
  XOR U6262 ( .A(n5263), .B(n5264), .Z(n4944) );
  XOR U6263 ( .A(round_reg[228]), .B(n5265), .Z(n5264) );
  XOR U6264 ( .A(round_reg[868]), .B(round_reg[548]), .Z(n5265) );
  XNOR U6265 ( .A(round_reg[1188]), .B(round_reg[1508]), .Z(n5263) );
  XOR U6266 ( .A(n1829), .B(round_reg[1349]), .Z(n1086) );
  XOR U6267 ( .A(n5132), .B(n5050), .Z(n1829) );
  XOR U6268 ( .A(n5266), .B(n5267), .Z(n5050) );
  XOR U6269 ( .A(round_reg[4]), .B(n5268), .Z(n5267) );
  XOR U6270 ( .A(round_reg[964]), .B(round_reg[644]), .Z(n5268) );
  XNOR U6271 ( .A(round_reg[1284]), .B(round_reg[324]), .Z(n5266) );
  XOR U6272 ( .A(n5269), .B(n5270), .Z(n5132) );
  XOR U6273 ( .A(round_reg[1413]), .B(n5271), .Z(n5270) );
  XOR U6274 ( .A(round_reg[773]), .B(round_reg[453]), .Z(n5271) );
  XNOR U6275 ( .A(round_reg[1093]), .B(round_reg[133]), .Z(n5269) );
  XOR U6276 ( .A(n5272), .B(n4708), .Z(o[1056]) );
  XOR U6277 ( .A(n2165), .B(round_reg[563]), .Z(n4708) );
  XNOR U6278 ( .A(n4808), .B(n5273), .Z(n2165) );
  XNOR U6279 ( .A(n5274), .B(n5275), .Z(n4808) );
  XOR U6280 ( .A(round_reg[307]), .B(n5276), .Z(n5275) );
  XOR U6281 ( .A(round_reg[947]), .B(round_reg[627]), .Z(n5276) );
  XNOR U6282 ( .A(round_reg[1267]), .B(round_reg[1587]), .Z(n5274) );
  ANDN U6283 ( .A(n1090), .B(n1088), .Z(n5272) );
  XNOR U6284 ( .A(n2212), .B(round_reg[163]), .Z(n1088) );
  XOR U6285 ( .A(n5278), .B(n5279), .Z(n4948) );
  XOR U6286 ( .A(round_reg[227]), .B(n5280), .Z(n5279) );
  XOR U6287 ( .A(round_reg[867]), .B(round_reg[547]), .Z(n5280) );
  XNOR U6288 ( .A(round_reg[1187]), .B(round_reg[1507]), .Z(n5278) );
  XOR U6289 ( .A(n1832), .B(round_reg[1348]), .Z(n1090) );
  XOR U6290 ( .A(n5137), .B(n5063), .Z(n1832) );
  XOR U6291 ( .A(n5281), .B(n5282), .Z(n5063) );
  XOR U6292 ( .A(round_reg[3]), .B(n5283), .Z(n5282) );
  XOR U6293 ( .A(round_reg[963]), .B(round_reg[643]), .Z(n5283) );
  XNOR U6294 ( .A(round_reg[1283]), .B(round_reg[323]), .Z(n5281) );
  XOR U6295 ( .A(n5284), .B(n5285), .Z(n5137) );
  XOR U6296 ( .A(round_reg[1412]), .B(n5286), .Z(n5285) );
  XOR U6297 ( .A(round_reg[772]), .B(round_reg[452]), .Z(n5286) );
  XNOR U6298 ( .A(round_reg[1092]), .B(round_reg[132]), .Z(n5284) );
  XOR U6299 ( .A(n5287), .B(n4712), .Z(o[1055]) );
  XOR U6300 ( .A(n2169), .B(round_reg[562]), .Z(n4712) );
  XNOR U6301 ( .A(n4815), .B(n5288), .Z(n2169) );
  XNOR U6302 ( .A(n5289), .B(n5290), .Z(n4815) );
  XOR U6303 ( .A(round_reg[306]), .B(n5291), .Z(n5290) );
  XOR U6304 ( .A(round_reg[946]), .B(round_reg[626]), .Z(n5291) );
  XNOR U6305 ( .A(round_reg[1266]), .B(round_reg[1586]), .Z(n5289) );
  ANDN U6306 ( .A(n1094), .B(n1092), .Z(n5287) );
  XOR U6307 ( .A(n2216), .B(round_reg[162]), .Z(n1092) );
  XOR U6308 ( .A(n4951), .B(n5292), .Z(n2216) );
  XOR U6309 ( .A(n5293), .B(n5294), .Z(n4951) );
  XOR U6310 ( .A(round_reg[226]), .B(n5295), .Z(n5294) );
  XOR U6311 ( .A(round_reg[866]), .B(round_reg[546]), .Z(n5295) );
  XNOR U6312 ( .A(round_reg[1186]), .B(round_reg[1506]), .Z(n5293) );
  XOR U6313 ( .A(n1835), .B(round_reg[1347]), .Z(n1094) );
  XOR U6314 ( .A(n5142), .B(n5110), .Z(n1835) );
  XOR U6315 ( .A(n5296), .B(n5297), .Z(n5110) );
  XOR U6316 ( .A(round_reg[322]), .B(n5298), .Z(n5297) );
  XOR U6317 ( .A(round_reg[962]), .B(round_reg[642]), .Z(n5298) );
  XNOR U6318 ( .A(round_reg[1282]), .B(round_reg[2]), .Z(n5296) );
  XOR U6319 ( .A(n5299), .B(n5300), .Z(n5142) );
  XOR U6320 ( .A(round_reg[1411]), .B(n5301), .Z(n5300) );
  XOR U6321 ( .A(round_reg[771]), .B(round_reg[451]), .Z(n5301) );
  XNOR U6322 ( .A(round_reg[1091]), .B(round_reg[131]), .Z(n5299) );
  XOR U6323 ( .A(n5302), .B(n4716), .Z(o[1054]) );
  XOR U6324 ( .A(n2173), .B(round_reg[561]), .Z(n4716) );
  XNOR U6325 ( .A(n4819), .B(n5303), .Z(n2173) );
  XNOR U6326 ( .A(n5304), .B(n5305), .Z(n4819) );
  XOR U6327 ( .A(round_reg[305]), .B(n5306), .Z(n5305) );
  XOR U6328 ( .A(round_reg[945]), .B(round_reg[625]), .Z(n5306) );
  XNOR U6329 ( .A(round_reg[1265]), .B(round_reg[1585]), .Z(n5304) );
  ANDN U6330 ( .A(n1098), .B(n1096), .Z(n5302) );
  XOR U6331 ( .A(n2224), .B(round_reg[161]), .Z(n1096) );
  XOR U6332 ( .A(n4954), .B(n5307), .Z(n2224) );
  XOR U6333 ( .A(n5308), .B(n5309), .Z(n4954) );
  XOR U6334 ( .A(round_reg[225]), .B(n5310), .Z(n5309) );
  XOR U6335 ( .A(round_reg[865]), .B(round_reg[545]), .Z(n5310) );
  XNOR U6336 ( .A(round_reg[1185]), .B(round_reg[1505]), .Z(n5308) );
  XOR U6337 ( .A(n1838), .B(round_reg[1346]), .Z(n1098) );
  XOR U6338 ( .A(n5147), .B(n5163), .Z(n1838) );
  XOR U6339 ( .A(n5311), .B(n5312), .Z(n5163) );
  XOR U6340 ( .A(round_reg[321]), .B(n5313), .Z(n5312) );
  XOR U6341 ( .A(round_reg[961]), .B(round_reg[641]), .Z(n5313) );
  XNOR U6342 ( .A(round_reg[1281]), .B(round_reg[1]), .Z(n5311) );
  XOR U6343 ( .A(n5314), .B(n5315), .Z(n5147) );
  XOR U6344 ( .A(round_reg[1410]), .B(n5316), .Z(n5315) );
  XOR U6345 ( .A(round_reg[770]), .B(round_reg[450]), .Z(n5316) );
  XNOR U6346 ( .A(round_reg[1090]), .B(round_reg[130]), .Z(n5314) );
  XOR U6347 ( .A(n5317), .B(n4720), .Z(o[1053]) );
  XOR U6348 ( .A(n2181), .B(round_reg[560]), .Z(n4720) );
  XNOR U6349 ( .A(n4823), .B(n5318), .Z(n2181) );
  XNOR U6350 ( .A(n5319), .B(n5320), .Z(n4823) );
  XOR U6351 ( .A(round_reg[304]), .B(n5321), .Z(n5320) );
  XOR U6352 ( .A(round_reg[944]), .B(round_reg[624]), .Z(n5321) );
  XNOR U6353 ( .A(round_reg[1264]), .B(round_reg[1584]), .Z(n5319) );
  AND U6354 ( .A(n1106), .B(n1104), .Z(n5317) );
  XNOR U6355 ( .A(n2228), .B(round_reg[160]), .Z(n1104) );
  XOR U6356 ( .A(n4957), .B(n5322), .Z(n2228) );
  XOR U6357 ( .A(n5323), .B(n5324), .Z(n4957) );
  XOR U6358 ( .A(round_reg[224]), .B(n5325), .Z(n5324) );
  XOR U6359 ( .A(round_reg[864]), .B(round_reg[544]), .Z(n5325) );
  XNOR U6360 ( .A(round_reg[1184]), .B(round_reg[1504]), .Z(n5323) );
  XOR U6361 ( .A(n1841), .B(round_reg[1345]), .Z(n1106) );
  XOR U6362 ( .A(n5152), .B(n5230), .Z(n1841) );
  XOR U6363 ( .A(n5326), .B(n5327), .Z(n5230) );
  XOR U6364 ( .A(round_reg[320]), .B(n5328), .Z(n5327) );
  XOR U6365 ( .A(round_reg[960]), .B(round_reg[640]), .Z(n5328) );
  XNOR U6366 ( .A(round_reg[0]), .B(round_reg[1280]), .Z(n5326) );
  XOR U6367 ( .A(n5329), .B(n5330), .Z(n5152) );
  XOR U6368 ( .A(round_reg[1409]), .B(n5331), .Z(n5330) );
  XOR U6369 ( .A(round_reg[769]), .B(round_reg[449]), .Z(n5331) );
  XNOR U6370 ( .A(round_reg[1089]), .B(round_reg[129]), .Z(n5329) );
  XOR U6371 ( .A(n5332), .B(n4724), .Z(o[1052]) );
  XOR U6372 ( .A(n2185), .B(round_reg[559]), .Z(n4724) );
  XNOR U6373 ( .A(n4827), .B(n5333), .Z(n2185) );
  XNOR U6374 ( .A(n5334), .B(n5335), .Z(n4827) );
  XOR U6375 ( .A(round_reg[303]), .B(n5336), .Z(n5335) );
  XOR U6376 ( .A(round_reg[943]), .B(round_reg[623]), .Z(n5336) );
  XNOR U6377 ( .A(round_reg[1263]), .B(round_reg[1583]), .Z(n5334) );
  AND U6378 ( .A(n1110), .B(n1108), .Z(n5332) );
  XNOR U6379 ( .A(n2232), .B(round_reg[159]), .Z(n1108) );
  XOR U6380 ( .A(n4960), .B(n5337), .Z(n2232) );
  XOR U6381 ( .A(n5338), .B(n5339), .Z(n4960) );
  XOR U6382 ( .A(round_reg[223]), .B(n5340), .Z(n5339) );
  XOR U6383 ( .A(round_reg[863]), .B(round_reg[543]), .Z(n5340) );
  XNOR U6384 ( .A(round_reg[1183]), .B(round_reg[1503]), .Z(n5338) );
  XOR U6385 ( .A(n1844), .B(round_reg[1344]), .Z(n1110) );
  XOR U6386 ( .A(n5157), .B(n5341), .Z(n1844) );
  XOR U6387 ( .A(n5342), .B(n5343), .Z(n5157) );
  XOR U6388 ( .A(round_reg[1408]), .B(n5344), .Z(n5343) );
  XOR U6389 ( .A(round_reg[768]), .B(round_reg[448]), .Z(n5344) );
  XNOR U6390 ( .A(round_reg[1088]), .B(round_reg[128]), .Z(n5342) );
  XOR U6391 ( .A(n5345), .B(n4731), .Z(o[1051]) );
  XOR U6392 ( .A(n2189), .B(round_reg[558]), .Z(n4731) );
  XNOR U6393 ( .A(n4831), .B(n5346), .Z(n2189) );
  XNOR U6394 ( .A(n5347), .B(n5348), .Z(n4831) );
  XOR U6395 ( .A(round_reg[302]), .B(n5349), .Z(n5348) );
  XOR U6396 ( .A(round_reg[942]), .B(round_reg[622]), .Z(n5349) );
  XNOR U6397 ( .A(round_reg[1262]), .B(round_reg[1582]), .Z(n5347) );
  ANDN U6398 ( .A(n1114), .B(n1112), .Z(n5345) );
  XOR U6399 ( .A(n2236), .B(round_reg[158]), .Z(n1112) );
  XOR U6400 ( .A(n4963), .B(n5350), .Z(n2236) );
  XOR U6401 ( .A(n5351), .B(n5352), .Z(n4963) );
  XOR U6402 ( .A(round_reg[222]), .B(n5353), .Z(n5352) );
  XOR U6403 ( .A(round_reg[862]), .B(round_reg[542]), .Z(n5353) );
  XNOR U6404 ( .A(round_reg[1182]), .B(round_reg[1502]), .Z(n5351) );
  XOR U6405 ( .A(n1847), .B(round_reg[1407]), .Z(n1114) );
  XOR U6406 ( .A(n5165), .B(n5354), .Z(n1847) );
  XOR U6407 ( .A(n5355), .B(n5356), .Z(n5165) );
  XOR U6408 ( .A(round_reg[191]), .B(n5357), .Z(n5356) );
  XOR U6409 ( .A(round_reg[831]), .B(round_reg[511]), .Z(n5357) );
  XNOR U6410 ( .A(round_reg[1151]), .B(round_reg[1471]), .Z(n5355) );
  XOR U6411 ( .A(n5358), .B(n4735), .Z(o[1050]) );
  XOR U6412 ( .A(n2193), .B(round_reg[557]), .Z(n4735) );
  XNOR U6413 ( .A(n4835), .B(n5359), .Z(n2193) );
  XNOR U6414 ( .A(n5360), .B(n5361), .Z(n4835) );
  XOR U6415 ( .A(round_reg[301]), .B(n5362), .Z(n5361) );
  XOR U6416 ( .A(round_reg[941]), .B(round_reg[621]), .Z(n5362) );
  XNOR U6417 ( .A(round_reg[1261]), .B(round_reg[1581]), .Z(n5360) );
  ANDN U6418 ( .A(n1118), .B(n1116), .Z(n5358) );
  XOR U6419 ( .A(n2240), .B(round_reg[157]), .Z(n1116) );
  XOR U6420 ( .A(n4966), .B(n5363), .Z(n2240) );
  XOR U6421 ( .A(n5364), .B(n5365), .Z(n4966) );
  XOR U6422 ( .A(round_reg[221]), .B(n5366), .Z(n5365) );
  XOR U6423 ( .A(round_reg[861]), .B(round_reg[541]), .Z(n5366) );
  XNOR U6424 ( .A(round_reg[1181]), .B(round_reg[1501]), .Z(n5364) );
  XOR U6425 ( .A(n1850), .B(round_reg[1406]), .Z(n1118) );
  XOR U6426 ( .A(n5170), .B(n5367), .Z(n1850) );
  XOR U6427 ( .A(n5368), .B(n5369), .Z(n5170) );
  XOR U6428 ( .A(round_reg[190]), .B(n5370), .Z(n5369) );
  XOR U6429 ( .A(round_reg[830]), .B(round_reg[510]), .Z(n5370) );
  XNOR U6430 ( .A(round_reg[1150]), .B(round_reg[1470]), .Z(n5368) );
  XOR U6431 ( .A(n5371), .B(n3507), .Z(o[104]) );
  XOR U6432 ( .A(n2319), .B(round_reg[639]), .Z(n3507) );
  IV U6433 ( .A(n5060), .Z(n2319) );
  XOR U6434 ( .A(n5372), .B(n5341), .Z(n5060) );
  XOR U6435 ( .A(n5373), .B(n5374), .Z(n5341) );
  XOR U6436 ( .A(round_reg[383]), .B(n5375), .Z(n5374) );
  XOR U6437 ( .A(round_reg[703]), .B(round_reg[63]), .Z(n5375) );
  XNOR U6438 ( .A(round_reg[1023]), .B(round_reg[1343]), .Z(n5373) );
  AND U6439 ( .A(n3125), .B(n3127), .Z(n5371) );
  XOR U6440 ( .A(n2184), .B(round_reg[1450]), .Z(n3127) );
  XOR U6441 ( .A(n4918), .B(n5376), .Z(n2184) );
  XOR U6442 ( .A(n5377), .B(n5378), .Z(n4918) );
  XOR U6443 ( .A(round_reg[234]), .B(n5379), .Z(n5378) );
  XOR U6444 ( .A(round_reg[874]), .B(round_reg[554]), .Z(n5379) );
  XNOR U6445 ( .A(round_reg[1194]), .B(round_reg[1514]), .Z(n5377) );
  XNOR U6446 ( .A(n2225), .B(round_reg[230]), .Z(n3125) );
  XOR U6447 ( .A(n5380), .B(n4739), .Z(o[1049]) );
  XOR U6448 ( .A(n2197), .B(round_reg[556]), .Z(n4739) );
  XNOR U6449 ( .A(n4839), .B(n5381), .Z(n2197) );
  XNOR U6450 ( .A(n5382), .B(n5383), .Z(n4839) );
  XOR U6451 ( .A(round_reg[300]), .B(n5384), .Z(n5383) );
  XOR U6452 ( .A(round_reg[940]), .B(round_reg[620]), .Z(n5384) );
  XNOR U6453 ( .A(round_reg[1260]), .B(round_reg[1580]), .Z(n5382) );
  ANDN U6454 ( .A(n1122), .B(n1120), .Z(n5380) );
  XOR U6455 ( .A(n2244), .B(round_reg[156]), .Z(n1120) );
  XOR U6456 ( .A(n4969), .B(n5385), .Z(n2244) );
  XOR U6457 ( .A(n5386), .B(n5387), .Z(n4969) );
  XOR U6458 ( .A(round_reg[220]), .B(n5388), .Z(n5387) );
  XOR U6459 ( .A(round_reg[860]), .B(round_reg[540]), .Z(n5388) );
  XNOR U6460 ( .A(round_reg[1180]), .B(round_reg[1500]), .Z(n5386) );
  XOR U6461 ( .A(n1853), .B(round_reg[1405]), .Z(n1122) );
  XOR U6462 ( .A(n5389), .B(n5390), .Z(n1853) );
  XOR U6463 ( .A(n5391), .B(n4743), .Z(o[1048]) );
  XOR U6464 ( .A(n2201), .B(round_reg[555]), .Z(n4743) );
  XNOR U6465 ( .A(n4843), .B(n5392), .Z(n2201) );
  XNOR U6466 ( .A(n5393), .B(n5394), .Z(n4843) );
  XOR U6467 ( .A(round_reg[299]), .B(n5395), .Z(n5394) );
  XOR U6468 ( .A(round_reg[939]), .B(round_reg[619]), .Z(n5395) );
  XNOR U6469 ( .A(round_reg[1259]), .B(round_reg[1579]), .Z(n5393) );
  ANDN U6470 ( .A(n1126), .B(n1124), .Z(n5391) );
  XOR U6471 ( .A(n2248), .B(round_reg[155]), .Z(n1124) );
  XOR U6472 ( .A(n4974), .B(n5396), .Z(n2248) );
  XOR U6473 ( .A(n5397), .B(n5398), .Z(n4974) );
  XOR U6474 ( .A(round_reg[219]), .B(n5399), .Z(n5398) );
  XOR U6475 ( .A(round_reg[859]), .B(round_reg[539]), .Z(n5399) );
  XNOR U6476 ( .A(round_reg[1179]), .B(round_reg[1499]), .Z(n5397) );
  XOR U6477 ( .A(n1860), .B(round_reg[1404]), .Z(n1126) );
  XOR U6478 ( .A(n5176), .B(n5400), .Z(n1860) );
  XOR U6479 ( .A(n5401), .B(n5402), .Z(n5176) );
  XOR U6480 ( .A(round_reg[188]), .B(n5403), .Z(n5402) );
  XOR U6481 ( .A(round_reg[828]), .B(round_reg[508]), .Z(n5403) );
  XNOR U6482 ( .A(round_reg[1148]), .B(round_reg[1468]), .Z(n5401) );
  XOR U6483 ( .A(n5404), .B(n4747), .Z(o[1047]) );
  XOR U6484 ( .A(n2205), .B(round_reg[554]), .Z(n4747) );
  XNOR U6485 ( .A(n5405), .B(n5406), .Z(n2205) );
  ANDN U6486 ( .A(n1130), .B(n1128), .Z(n5404) );
  XOR U6487 ( .A(n2252), .B(round_reg[154]), .Z(n1128) );
  XOR U6488 ( .A(n4977), .B(n5407), .Z(n2252) );
  XOR U6489 ( .A(n5408), .B(n5409), .Z(n4977) );
  XOR U6490 ( .A(round_reg[218]), .B(n5410), .Z(n5409) );
  XOR U6491 ( .A(round_reg[858]), .B(round_reg[538]), .Z(n5410) );
  XNOR U6492 ( .A(round_reg[1178]), .B(round_reg[1498]), .Z(n5408) );
  XOR U6493 ( .A(n1863), .B(round_reg[1403]), .Z(n1130) );
  XOR U6494 ( .A(n5181), .B(n4856), .Z(n1863) );
  XOR U6495 ( .A(n5411), .B(n5412), .Z(n4856) );
  XOR U6496 ( .A(round_reg[378]), .B(n5413), .Z(n5412) );
  XOR U6497 ( .A(round_reg[698]), .B(round_reg[58]), .Z(n5413) );
  XNOR U6498 ( .A(round_reg[1018]), .B(round_reg[1338]), .Z(n5411) );
  XOR U6499 ( .A(n5414), .B(n5415), .Z(n5181) );
  XOR U6500 ( .A(round_reg[187]), .B(n5416), .Z(n5415) );
  XOR U6501 ( .A(round_reg[827]), .B(round_reg[507]), .Z(n5416) );
  XNOR U6502 ( .A(round_reg[1147]), .B(round_reg[1467]), .Z(n5414) );
  XOR U6503 ( .A(n5417), .B(n4751), .Z(o[1046]) );
  XOR U6504 ( .A(n2209), .B(round_reg[553]), .Z(n4751) );
  XNOR U6505 ( .A(n5418), .B(n5419), .Z(n2209) );
  ANDN U6506 ( .A(n1134), .B(n1132), .Z(n5417) );
  XOR U6507 ( .A(n2256), .B(round_reg[153]), .Z(n1132) );
  XOR U6508 ( .A(n4980), .B(n5420), .Z(n2256) );
  XOR U6509 ( .A(n5421), .B(n5422), .Z(n4980) );
  XOR U6510 ( .A(round_reg[217]), .B(n5423), .Z(n5422) );
  XOR U6511 ( .A(round_reg[857]), .B(round_reg[537]), .Z(n5423) );
  XNOR U6512 ( .A(round_reg[1177]), .B(round_reg[1497]), .Z(n5421) );
  XOR U6513 ( .A(n1866), .B(round_reg[1402]), .Z(n1134) );
  XOR U6514 ( .A(n5186), .B(n4860), .Z(n1866) );
  XOR U6515 ( .A(n5424), .B(n5425), .Z(n4860) );
  XOR U6516 ( .A(round_reg[377]), .B(n5426), .Z(n5425) );
  XOR U6517 ( .A(round_reg[697]), .B(round_reg[57]), .Z(n5426) );
  XNOR U6518 ( .A(round_reg[1017]), .B(round_reg[1337]), .Z(n5424) );
  XOR U6519 ( .A(n5427), .B(n5428), .Z(n5186) );
  XOR U6520 ( .A(round_reg[186]), .B(n5429), .Z(n5428) );
  XOR U6521 ( .A(round_reg[826]), .B(round_reg[506]), .Z(n5429) );
  XNOR U6522 ( .A(round_reg[1146]), .B(round_reg[1466]), .Z(n5427) );
  XOR U6523 ( .A(n5430), .B(n4755), .Z(o[1045]) );
  XOR U6524 ( .A(n2213), .B(round_reg[552]), .Z(n4755) );
  XNOR U6525 ( .A(n5431), .B(n5432), .Z(n2213) );
  ANDN U6526 ( .A(n1138), .B(n1136), .Z(n5430) );
  XOR U6527 ( .A(n2260), .B(round_reg[152]), .Z(n1136) );
  XOR U6528 ( .A(n4983), .B(n5433), .Z(n2260) );
  XOR U6529 ( .A(n5434), .B(n5435), .Z(n4983) );
  XOR U6530 ( .A(round_reg[216]), .B(n5436), .Z(n5435) );
  XOR U6531 ( .A(round_reg[856]), .B(round_reg[536]), .Z(n5436) );
  XNOR U6532 ( .A(round_reg[1176]), .B(round_reg[1496]), .Z(n5434) );
  XOR U6533 ( .A(n1869), .B(round_reg[1401]), .Z(n1138) );
  XOR U6534 ( .A(n5191), .B(n4864), .Z(n1869) );
  XOR U6535 ( .A(n5437), .B(n5438), .Z(n4864) );
  XOR U6536 ( .A(round_reg[376]), .B(n5439), .Z(n5438) );
  XOR U6537 ( .A(round_reg[696]), .B(round_reg[56]), .Z(n5439) );
  XNOR U6538 ( .A(round_reg[1016]), .B(round_reg[1336]), .Z(n5437) );
  XOR U6539 ( .A(n5440), .B(n5441), .Z(n5191) );
  XOR U6540 ( .A(round_reg[185]), .B(n5442), .Z(n5441) );
  XOR U6541 ( .A(round_reg[825]), .B(round_reg[505]), .Z(n5442) );
  XNOR U6542 ( .A(round_reg[1145]), .B(round_reg[1465]), .Z(n5440) );
  XOR U6543 ( .A(n5443), .B(n4759), .Z(o[1044]) );
  XOR U6544 ( .A(n2217), .B(round_reg[551]), .Z(n4759) );
  XNOR U6545 ( .A(n5444), .B(n5445), .Z(n2217) );
  ANDN U6546 ( .A(n1142), .B(n1140), .Z(n5443) );
  XOR U6547 ( .A(n2268), .B(round_reg[151]), .Z(n1140) );
  XOR U6548 ( .A(n4986), .B(n5446), .Z(n2268) );
  XOR U6549 ( .A(n5447), .B(n5448), .Z(n4986) );
  XOR U6550 ( .A(round_reg[215]), .B(n5449), .Z(n5448) );
  XOR U6551 ( .A(round_reg[855]), .B(round_reg[535]), .Z(n5449) );
  XNOR U6552 ( .A(round_reg[1175]), .B(round_reg[1495]), .Z(n5447) );
  XOR U6553 ( .A(n1872), .B(round_reg[1400]), .Z(n1142) );
  XOR U6554 ( .A(n5202), .B(n4868), .Z(n1872) );
  XOR U6555 ( .A(n5450), .B(n5451), .Z(n4868) );
  XOR U6556 ( .A(round_reg[375]), .B(n5452), .Z(n5451) );
  XOR U6557 ( .A(round_reg[695]), .B(round_reg[55]), .Z(n5452) );
  XNOR U6558 ( .A(round_reg[1015]), .B(round_reg[1335]), .Z(n5450) );
  XOR U6559 ( .A(n5453), .B(n5454), .Z(n5202) );
  XOR U6560 ( .A(round_reg[184]), .B(n5455), .Z(n5454) );
  XOR U6561 ( .A(round_reg[824]), .B(round_reg[504]), .Z(n5455) );
  XNOR U6562 ( .A(round_reg[1144]), .B(round_reg[1464]), .Z(n5453) );
  XOR U6563 ( .A(n5456), .B(n4763), .Z(o[1043]) );
  XOR U6564 ( .A(n2225), .B(round_reg[550]), .Z(n4763) );
  XNOR U6565 ( .A(n5457), .B(n5458), .Z(n2225) );
  ANDN U6566 ( .A(n1150), .B(n1148), .Z(n5456) );
  XOR U6567 ( .A(n2272), .B(round_reg[150]), .Z(n1148) );
  XOR U6568 ( .A(n4989), .B(n5459), .Z(n2272) );
  XOR U6569 ( .A(n5460), .B(n5461), .Z(n4989) );
  XOR U6570 ( .A(round_reg[214]), .B(n5462), .Z(n5461) );
  XOR U6571 ( .A(round_reg[854]), .B(round_reg[534]), .Z(n5462) );
  XNOR U6572 ( .A(round_reg[1174]), .B(round_reg[1494]), .Z(n5460) );
  XOR U6573 ( .A(n1875), .B(round_reg[1399]), .Z(n1150) );
  XOR U6574 ( .A(n5213), .B(n4872), .Z(n1875) );
  XOR U6575 ( .A(n5463), .B(n5464), .Z(n4872) );
  XOR U6576 ( .A(round_reg[374]), .B(n5465), .Z(n5464) );
  XOR U6577 ( .A(round_reg[694]), .B(round_reg[54]), .Z(n5465) );
  XNOR U6578 ( .A(round_reg[1014]), .B(round_reg[1334]), .Z(n5463) );
  XOR U6579 ( .A(n5466), .B(n5467), .Z(n5213) );
  XOR U6580 ( .A(round_reg[183]), .B(n5468), .Z(n5467) );
  XOR U6581 ( .A(round_reg[823]), .B(round_reg[503]), .Z(n5468) );
  XNOR U6582 ( .A(round_reg[1143]), .B(round_reg[1463]), .Z(n5466) );
  XOR U6583 ( .A(n5469), .B(n4767), .Z(o[1042]) );
  XOR U6584 ( .A(n2229), .B(round_reg[549]), .Z(n4767) );
  ANDN U6585 ( .A(n1154), .B(n1152), .Z(n5469) );
  XOR U6586 ( .A(n2276), .B(round_reg[149]), .Z(n1152) );
  XOR U6587 ( .A(n4992), .B(n5470), .Z(n2276) );
  XOR U6588 ( .A(n5471), .B(n5472), .Z(n4992) );
  XOR U6589 ( .A(round_reg[213]), .B(n5473), .Z(n5472) );
  XOR U6590 ( .A(round_reg[853]), .B(round_reg[533]), .Z(n5473) );
  XNOR U6591 ( .A(round_reg[1173]), .B(round_reg[1493]), .Z(n5471) );
  XOR U6592 ( .A(n1878), .B(round_reg[1398]), .Z(n1154) );
  XOR U6593 ( .A(n5218), .B(n4876), .Z(n1878) );
  XOR U6594 ( .A(n5474), .B(n5475), .Z(n4876) );
  XOR U6595 ( .A(round_reg[373]), .B(n5476), .Z(n5475) );
  XOR U6596 ( .A(round_reg[693]), .B(round_reg[53]), .Z(n5476) );
  XNOR U6597 ( .A(round_reg[1013]), .B(round_reg[1333]), .Z(n5474) );
  XOR U6598 ( .A(n5477), .B(n5478), .Z(n5218) );
  XOR U6599 ( .A(round_reg[182]), .B(n5479), .Z(n5478) );
  XOR U6600 ( .A(round_reg[822]), .B(round_reg[502]), .Z(n5479) );
  XNOR U6601 ( .A(round_reg[1142]), .B(round_reg[1462]), .Z(n5477) );
  XOR U6602 ( .A(n5480), .B(n4774), .Z(o[1041]) );
  XOR U6603 ( .A(n2233), .B(round_reg[548]), .Z(n4774) );
  ANDN U6604 ( .A(n1158), .B(n1156), .Z(n5480) );
  XOR U6605 ( .A(n2280), .B(round_reg[148]), .Z(n1156) );
  XOR U6606 ( .A(n4995), .B(n4676), .Z(n2280) );
  XOR U6607 ( .A(n5481), .B(n5482), .Z(n4676) );
  XOR U6608 ( .A(round_reg[403]), .B(n5483), .Z(n5482) );
  XOR U6609 ( .A(round_reg[83]), .B(round_reg[723]), .Z(n5483) );
  XNOR U6610 ( .A(round_reg[1043]), .B(round_reg[1363]), .Z(n5481) );
  XOR U6611 ( .A(n5484), .B(n5485), .Z(n4995) );
  XOR U6612 ( .A(round_reg[212]), .B(n5486), .Z(n5485) );
  XOR U6613 ( .A(round_reg[852]), .B(round_reg[532]), .Z(n5486) );
  XNOR U6614 ( .A(round_reg[1172]), .B(round_reg[1492]), .Z(n5484) );
  XOR U6615 ( .A(n1881), .B(round_reg[1397]), .Z(n1158) );
  XOR U6616 ( .A(n5232), .B(n4880), .Z(n1881) );
  XOR U6617 ( .A(n5487), .B(n5488), .Z(n4880) );
  XOR U6618 ( .A(round_reg[372]), .B(n5489), .Z(n5488) );
  XOR U6619 ( .A(round_reg[692]), .B(round_reg[52]), .Z(n5489) );
  XNOR U6620 ( .A(round_reg[1012]), .B(round_reg[1332]), .Z(n5487) );
  XOR U6621 ( .A(n5490), .B(n5491), .Z(n5232) );
  XOR U6622 ( .A(round_reg[181]), .B(n5492), .Z(n5491) );
  XOR U6623 ( .A(round_reg[821]), .B(round_reg[501]), .Z(n5492) );
  XNOR U6624 ( .A(round_reg[1141]), .B(round_reg[1461]), .Z(n5490) );
  XOR U6625 ( .A(n5493), .B(n4778), .Z(o[1040]) );
  XOR U6626 ( .A(n2237), .B(round_reg[547]), .Z(n4778) );
  ANDN U6627 ( .A(n1162), .B(n1160), .Z(n5493) );
  XOR U6628 ( .A(n2284), .B(round_reg[147]), .Z(n1160) );
  XOR U6629 ( .A(n4998), .B(n4680), .Z(n2284) );
  XOR U6630 ( .A(n5494), .B(n5495), .Z(n4680) );
  XOR U6631 ( .A(round_reg[402]), .B(n5496), .Z(n5495) );
  XOR U6632 ( .A(round_reg[82]), .B(round_reg[722]), .Z(n5496) );
  XNOR U6633 ( .A(round_reg[1042]), .B(round_reg[1362]), .Z(n5494) );
  XOR U6634 ( .A(n5497), .B(n5498), .Z(n4998) );
  XOR U6635 ( .A(round_reg[211]), .B(n5499), .Z(n5498) );
  XOR U6636 ( .A(round_reg[851]), .B(round_reg[531]), .Z(n5499) );
  XNOR U6637 ( .A(round_reg[1171]), .B(round_reg[1491]), .Z(n5497) );
  XOR U6638 ( .A(n1884), .B(round_reg[1396]), .Z(n1162) );
  XOR U6639 ( .A(n5243), .B(n4884), .Z(n1884) );
  XOR U6640 ( .A(n5500), .B(n5501), .Z(n4884) );
  XOR U6641 ( .A(round_reg[371]), .B(n5502), .Z(n5501) );
  XOR U6642 ( .A(round_reg[691]), .B(round_reg[51]), .Z(n5502) );
  XNOR U6643 ( .A(round_reg[1011]), .B(round_reg[1331]), .Z(n5500) );
  XOR U6644 ( .A(n5503), .B(n5504), .Z(n5243) );
  XOR U6645 ( .A(round_reg[180]), .B(n5505), .Z(n5504) );
  XOR U6646 ( .A(round_reg[820]), .B(round_reg[500]), .Z(n5505) );
  XNOR U6647 ( .A(round_reg[1140]), .B(round_reg[1460]), .Z(n5503) );
  XOR U6648 ( .A(n5506), .B(n3509), .Z(o[103]) );
  XOR U6649 ( .A(n2323), .B(round_reg[638]), .Z(n3509) );
  IV U6650 ( .A(n5065), .Z(n2323) );
  XOR U6651 ( .A(n5507), .B(n5354), .Z(n5065) );
  XOR U6652 ( .A(n5508), .B(n5509), .Z(n5354) );
  XOR U6653 ( .A(round_reg[382]), .B(n5510), .Z(n5509) );
  XOR U6654 ( .A(round_reg[702]), .B(round_reg[62]), .Z(n5510) );
  XNOR U6655 ( .A(round_reg[1022]), .B(round_reg[1342]), .Z(n5508) );
  AND U6656 ( .A(n3151), .B(n3153), .Z(n5506) );
  XOR U6657 ( .A(n2188), .B(round_reg[1449]), .Z(n3153) );
  XOR U6658 ( .A(n4922), .B(n5511), .Z(n2188) );
  XOR U6659 ( .A(n5512), .B(n5513), .Z(n4922) );
  XOR U6660 ( .A(round_reg[233]), .B(n5514), .Z(n5513) );
  XOR U6661 ( .A(round_reg[873]), .B(round_reg[553]), .Z(n5514) );
  XNOR U6662 ( .A(round_reg[1193]), .B(round_reg[1513]), .Z(n5512) );
  XNOR U6663 ( .A(n2229), .B(round_reg[229]), .Z(n3151) );
  XNOR U6664 ( .A(n5515), .B(n5516), .Z(n2229) );
  XOR U6665 ( .A(n5517), .B(n4782), .Z(o[1039]) );
  XOR U6666 ( .A(n2241), .B(round_reg[546]), .Z(n4782) );
  AND U6667 ( .A(n1166), .B(n1164), .Z(n5517) );
  XNOR U6668 ( .A(n2288), .B(round_reg[146]), .Z(n1164) );
  XOR U6669 ( .A(n5001), .B(n4687), .Z(n2288) );
  XOR U6670 ( .A(n5518), .B(n5519), .Z(n4687) );
  XOR U6671 ( .A(round_reg[401]), .B(n5520), .Z(n5519) );
  XOR U6672 ( .A(round_reg[81]), .B(round_reg[721]), .Z(n5520) );
  XNOR U6673 ( .A(round_reg[1041]), .B(round_reg[1361]), .Z(n5518) );
  XOR U6674 ( .A(n5521), .B(n5522), .Z(n5001) );
  XOR U6675 ( .A(round_reg[210]), .B(n5523), .Z(n5522) );
  XOR U6676 ( .A(round_reg[850]), .B(round_reg[530]), .Z(n5523) );
  XNOR U6677 ( .A(round_reg[1170]), .B(round_reg[1490]), .Z(n5521) );
  XOR U6678 ( .A(n1887), .B(round_reg[1395]), .Z(n1166) );
  XOR U6679 ( .A(n5258), .B(n4888), .Z(n1887) );
  XOR U6680 ( .A(n5524), .B(n5525), .Z(n4888) );
  XOR U6681 ( .A(round_reg[370]), .B(n5526), .Z(n5525) );
  XOR U6682 ( .A(round_reg[690]), .B(round_reg[50]), .Z(n5526) );
  XNOR U6683 ( .A(round_reg[1010]), .B(round_reg[1330]), .Z(n5524) );
  XOR U6684 ( .A(n5527), .B(n5528), .Z(n5258) );
  XOR U6685 ( .A(round_reg[179]), .B(n5529), .Z(n5528) );
  XOR U6686 ( .A(round_reg[819]), .B(round_reg[499]), .Z(n5529) );
  XNOR U6687 ( .A(round_reg[1139]), .B(round_reg[1459]), .Z(n5527) );
  XOR U6688 ( .A(n5530), .B(n4786), .Z(o[1038]) );
  XOR U6689 ( .A(n2245), .B(round_reg[545]), .Z(n4786) );
  XOR U6690 ( .A(n5531), .B(n5532), .Z(n2245) );
  ANDN U6691 ( .A(n1170), .B(n1168), .Z(n5530) );
  XOR U6692 ( .A(n2292), .B(round_reg[145]), .Z(n1168) );
  XOR U6693 ( .A(n5005), .B(n4691), .Z(n2292) );
  XOR U6694 ( .A(n5533), .B(n5534), .Z(n4691) );
  XOR U6695 ( .A(round_reg[400]), .B(n5535), .Z(n5534) );
  XOR U6696 ( .A(round_reg[80]), .B(round_reg[720]), .Z(n5535) );
  XNOR U6697 ( .A(round_reg[1040]), .B(round_reg[1360]), .Z(n5533) );
  XOR U6698 ( .A(n5536), .B(n5537), .Z(n5005) );
  XOR U6699 ( .A(round_reg[209]), .B(n5538), .Z(n5537) );
  XOR U6700 ( .A(round_reg[849]), .B(round_reg[529]), .Z(n5538) );
  XNOR U6701 ( .A(round_reg[1169]), .B(round_reg[1489]), .Z(n5536) );
  XOR U6702 ( .A(n1894), .B(round_reg[1394]), .Z(n1170) );
  XOR U6703 ( .A(n5273), .B(n4892), .Z(n1894) );
  XOR U6704 ( .A(n5539), .B(n5540), .Z(n4892) );
  XOR U6705 ( .A(round_reg[369]), .B(n5541), .Z(n5540) );
  XOR U6706 ( .A(round_reg[689]), .B(round_reg[49]), .Z(n5541) );
  XNOR U6707 ( .A(round_reg[1009]), .B(round_reg[1329]), .Z(n5539) );
  XOR U6708 ( .A(n5542), .B(n5543), .Z(n5273) );
  XOR U6709 ( .A(round_reg[178]), .B(n5544), .Z(n5543) );
  XOR U6710 ( .A(round_reg[818]), .B(round_reg[498]), .Z(n5544) );
  XNOR U6711 ( .A(round_reg[1138]), .B(round_reg[1458]), .Z(n5542) );
  XOR U6712 ( .A(n5545), .B(n4790), .Z(o[1037]) );
  XNOR U6713 ( .A(n2249), .B(round_reg[544]), .Z(n4790) );
  ANDN U6714 ( .A(n1174), .B(n1172), .Z(n5545) );
  XOR U6715 ( .A(n2296), .B(round_reg[144]), .Z(n1172) );
  XNOR U6716 ( .A(n5007), .B(n4695), .Z(n2296) );
  XOR U6717 ( .A(n5548), .B(n5549), .Z(n4695) );
  XOR U6718 ( .A(round_reg[399]), .B(n5550), .Z(n5549) );
  XOR U6719 ( .A(round_reg[79]), .B(round_reg[719]), .Z(n5550) );
  XNOR U6720 ( .A(round_reg[1039]), .B(round_reg[1359]), .Z(n5548) );
  XNOR U6721 ( .A(n5551), .B(n5552), .Z(n5007) );
  XOR U6722 ( .A(round_reg[208]), .B(n5553), .Z(n5552) );
  XOR U6723 ( .A(round_reg[848]), .B(round_reg[528]), .Z(n5553) );
  XNOR U6724 ( .A(round_reg[1168]), .B(round_reg[1488]), .Z(n5551) );
  XOR U6725 ( .A(n1897), .B(round_reg[1393]), .Z(n1174) );
  XOR U6726 ( .A(n5288), .B(n4898), .Z(n1897) );
  XOR U6727 ( .A(n5554), .B(n5555), .Z(n4898) );
  XOR U6728 ( .A(round_reg[368]), .B(n5556), .Z(n5555) );
  XOR U6729 ( .A(round_reg[688]), .B(round_reg[48]), .Z(n5556) );
  XNOR U6730 ( .A(round_reg[1008]), .B(round_reg[1328]), .Z(n5554) );
  XOR U6731 ( .A(n5557), .B(n5558), .Z(n5288) );
  XOR U6732 ( .A(round_reg[177]), .B(n5559), .Z(n5558) );
  XOR U6733 ( .A(round_reg[817]), .B(round_reg[497]), .Z(n5559) );
  XNOR U6734 ( .A(round_reg[1137]), .B(round_reg[1457]), .Z(n5557) );
  XOR U6735 ( .A(n5560), .B(n4794), .Z(o[1036]) );
  XNOR U6736 ( .A(n2253), .B(round_reg[543]), .Z(n4794) );
  ANDN U6737 ( .A(n1178), .B(n1176), .Z(n5560) );
  XOR U6738 ( .A(n2300), .B(round_reg[143]), .Z(n1176) );
  XOR U6739 ( .A(n5011), .B(n4699), .Z(n2300) );
  XOR U6740 ( .A(n5563), .B(n5564), .Z(n4699) );
  XOR U6741 ( .A(round_reg[398]), .B(n5565), .Z(n5564) );
  XOR U6742 ( .A(round_reg[78]), .B(round_reg[718]), .Z(n5565) );
  XNOR U6743 ( .A(round_reg[1038]), .B(round_reg[1358]), .Z(n5563) );
  XOR U6744 ( .A(n5566), .B(n5567), .Z(n5011) );
  XOR U6745 ( .A(round_reg[207]), .B(n5568), .Z(n5567) );
  XOR U6746 ( .A(round_reg[847]), .B(round_reg[527]), .Z(n5568) );
  XNOR U6747 ( .A(round_reg[1167]), .B(round_reg[1487]), .Z(n5566) );
  XOR U6748 ( .A(n1900), .B(round_reg[1392]), .Z(n1178) );
  XOR U6749 ( .A(n5303), .B(n4902), .Z(n1900) );
  XOR U6750 ( .A(n5569), .B(n5570), .Z(n4902) );
  XOR U6751 ( .A(round_reg[367]), .B(n5571), .Z(n5570) );
  XOR U6752 ( .A(round_reg[687]), .B(round_reg[47]), .Z(n5571) );
  XNOR U6753 ( .A(round_reg[1007]), .B(round_reg[1327]), .Z(n5569) );
  XOR U6754 ( .A(n5572), .B(n5573), .Z(n5303) );
  XOR U6755 ( .A(round_reg[176]), .B(n5574), .Z(n5573) );
  XOR U6756 ( .A(round_reg[816]), .B(round_reg[496]), .Z(n5574) );
  XNOR U6757 ( .A(round_reg[1136]), .B(round_reg[1456]), .Z(n5572) );
  XOR U6758 ( .A(n5575), .B(n4798), .Z(o[1035]) );
  XNOR U6759 ( .A(n2257), .B(round_reg[542]), .Z(n4798) );
  ANDN U6760 ( .A(n1182), .B(n1180), .Z(n5575) );
  XOR U6761 ( .A(n2304), .B(round_reg[142]), .Z(n1180) );
  XOR U6762 ( .A(n5014), .B(n4703), .Z(n2304) );
  XOR U6763 ( .A(n5578), .B(n5579), .Z(n4703) );
  XOR U6764 ( .A(round_reg[397]), .B(n5580), .Z(n5579) );
  XOR U6765 ( .A(round_reg[77]), .B(round_reg[717]), .Z(n5580) );
  XNOR U6766 ( .A(round_reg[1037]), .B(round_reg[1357]), .Z(n5578) );
  XOR U6767 ( .A(n5581), .B(n5582), .Z(n5014) );
  XOR U6768 ( .A(round_reg[206]), .B(n5583), .Z(n5582) );
  XOR U6769 ( .A(round_reg[846]), .B(round_reg[526]), .Z(n5583) );
  XNOR U6770 ( .A(round_reg[1166]), .B(round_reg[1486]), .Z(n5581) );
  XOR U6771 ( .A(n1903), .B(round_reg[1391]), .Z(n1182) );
  XOR U6772 ( .A(n5318), .B(n4906), .Z(n1903) );
  XOR U6773 ( .A(n5584), .B(n5585), .Z(n4906) );
  XOR U6774 ( .A(round_reg[366]), .B(n5586), .Z(n5585) );
  XOR U6775 ( .A(round_reg[686]), .B(round_reg[46]), .Z(n5586) );
  XNOR U6776 ( .A(round_reg[1006]), .B(round_reg[1326]), .Z(n5584) );
  XOR U6777 ( .A(n5587), .B(n5588), .Z(n5318) );
  XOR U6778 ( .A(round_reg[175]), .B(n5589), .Z(n5588) );
  XOR U6779 ( .A(round_reg[815]), .B(round_reg[495]), .Z(n5589) );
  XNOR U6780 ( .A(round_reg[1135]), .B(round_reg[1455]), .Z(n5587) );
  XOR U6781 ( .A(n5590), .B(n4802), .Z(o[1034]) );
  XNOR U6782 ( .A(n2261), .B(round_reg[541]), .Z(n4802) );
  ANDN U6783 ( .A(n1186), .B(n1184), .Z(n5590) );
  XOR U6784 ( .A(n2312), .B(round_reg[141]), .Z(n1184) );
  XOR U6785 ( .A(n5017), .B(n4707), .Z(n2312) );
  XOR U6786 ( .A(n5593), .B(n5594), .Z(n4707) );
  XOR U6787 ( .A(round_reg[396]), .B(n5595), .Z(n5594) );
  XOR U6788 ( .A(round_reg[76]), .B(round_reg[716]), .Z(n5595) );
  XNOR U6789 ( .A(round_reg[1036]), .B(round_reg[1356]), .Z(n5593) );
  XOR U6790 ( .A(n5596), .B(n5597), .Z(n5017) );
  XOR U6791 ( .A(round_reg[205]), .B(n5598), .Z(n5597) );
  XOR U6792 ( .A(round_reg[845]), .B(round_reg[525]), .Z(n5598) );
  XNOR U6793 ( .A(round_reg[1165]), .B(round_reg[1485]), .Z(n5596) );
  XOR U6794 ( .A(n1906), .B(round_reg[1390]), .Z(n1186) );
  XOR U6795 ( .A(n5333), .B(n4910), .Z(n1906) );
  XOR U6796 ( .A(n5599), .B(n5600), .Z(n4910) );
  XOR U6797 ( .A(round_reg[365]), .B(n5601), .Z(n5600) );
  XOR U6798 ( .A(round_reg[685]), .B(round_reg[45]), .Z(n5601) );
  XNOR U6799 ( .A(round_reg[1005]), .B(round_reg[1325]), .Z(n5599) );
  XOR U6800 ( .A(n5602), .B(n5603), .Z(n5333) );
  XOR U6801 ( .A(round_reg[174]), .B(n5604), .Z(n5603) );
  XOR U6802 ( .A(round_reg[814]), .B(round_reg[494]), .Z(n5604) );
  XNOR U6803 ( .A(round_reg[1134]), .B(round_reg[1454]), .Z(n5602) );
  XOR U6804 ( .A(n5605), .B(n4806), .Z(o[1033]) );
  XNOR U6805 ( .A(n2269), .B(round_reg[540]), .Z(n4806) );
  ANDN U6806 ( .A(n1194), .B(n1192), .Z(n5605) );
  XOR U6807 ( .A(n2316), .B(round_reg[140]), .Z(n1192) );
  XOR U6808 ( .A(n5020), .B(n4711), .Z(n2316) );
  XOR U6809 ( .A(n5608), .B(n5609), .Z(n4711) );
  XOR U6810 ( .A(round_reg[395]), .B(n5610), .Z(n5609) );
  XOR U6811 ( .A(round_reg[75]), .B(round_reg[715]), .Z(n5610) );
  XNOR U6812 ( .A(round_reg[1035]), .B(round_reg[1355]), .Z(n5608) );
  XOR U6813 ( .A(n5611), .B(n5612), .Z(n5020) );
  XOR U6814 ( .A(round_reg[204]), .B(n5613), .Z(n5612) );
  XOR U6815 ( .A(round_reg[844]), .B(round_reg[524]), .Z(n5613) );
  XNOR U6816 ( .A(round_reg[1164]), .B(round_reg[1484]), .Z(n5611) );
  XOR U6817 ( .A(n1909), .B(round_reg[1389]), .Z(n1194) );
  XOR U6818 ( .A(n5346), .B(n4914), .Z(n1909) );
  XOR U6819 ( .A(n5614), .B(n5615), .Z(n4914) );
  XOR U6820 ( .A(round_reg[364]), .B(n5616), .Z(n5615) );
  XOR U6821 ( .A(round_reg[684]), .B(round_reg[44]), .Z(n5616) );
  XNOR U6822 ( .A(round_reg[1004]), .B(round_reg[1324]), .Z(n5614) );
  XOR U6823 ( .A(n5617), .B(n5618), .Z(n5346) );
  XOR U6824 ( .A(round_reg[173]), .B(n5619), .Z(n5618) );
  XOR U6825 ( .A(round_reg[813]), .B(round_reg[493]), .Z(n5619) );
  XNOR U6826 ( .A(round_reg[1133]), .B(round_reg[1453]), .Z(n5617) );
  XOR U6827 ( .A(n5620), .B(n4810), .Z(o[1032]) );
  XOR U6828 ( .A(n2273), .B(round_reg[539]), .Z(n4810) );
  XNOR U6829 ( .A(n5621), .B(n5622), .Z(n2273) );
  AND U6830 ( .A(n1198), .B(n1196), .Z(n5620) );
  XNOR U6831 ( .A(n2320), .B(round_reg[139]), .Z(n1196) );
  XOR U6832 ( .A(n5023), .B(n4715), .Z(n2320) );
  XOR U6833 ( .A(n5623), .B(n5624), .Z(n4715) );
  XOR U6834 ( .A(round_reg[394]), .B(n5625), .Z(n5624) );
  XOR U6835 ( .A(round_reg[74]), .B(round_reg[714]), .Z(n5625) );
  XNOR U6836 ( .A(round_reg[1034]), .B(round_reg[1354]), .Z(n5623) );
  XOR U6837 ( .A(n5626), .B(n5627), .Z(n5023) );
  XOR U6838 ( .A(round_reg[203]), .B(n5628), .Z(n5627) );
  XOR U6839 ( .A(round_reg[843]), .B(round_reg[523]), .Z(n5628) );
  XNOR U6840 ( .A(round_reg[1163]), .B(round_reg[1483]), .Z(n5626) );
  XNOR U6841 ( .A(n1912), .B(round_reg[1388]), .Z(n1198) );
  XNOR U6842 ( .A(n5629), .B(n5630), .Z(n4917) );
  XOR U6843 ( .A(round_reg[363]), .B(n5631), .Z(n5630) );
  XOR U6844 ( .A(round_reg[683]), .B(round_reg[43]), .Z(n5631) );
  XNOR U6845 ( .A(round_reg[1003]), .B(round_reg[1323]), .Z(n5629) );
  XOR U6846 ( .A(n5632), .B(n5633), .Z(n5359) );
  XOR U6847 ( .A(round_reg[172]), .B(n5634), .Z(n5633) );
  XOR U6848 ( .A(round_reg[812]), .B(round_reg[492]), .Z(n5634) );
  XNOR U6849 ( .A(round_reg[1132]), .B(round_reg[1452]), .Z(n5632) );
  XOR U6850 ( .A(n5635), .B(n4817), .Z(o[1031]) );
  XOR U6851 ( .A(n2277), .B(round_reg[538]), .Z(n4817) );
  XNOR U6852 ( .A(n5636), .B(n5637), .Z(n2277) );
  AND U6853 ( .A(n1202), .B(n1200), .Z(n5635) );
  XNOR U6854 ( .A(n2324), .B(round_reg[138]), .Z(n1200) );
  XOR U6855 ( .A(n5026), .B(n4719), .Z(n2324) );
  XOR U6856 ( .A(n5638), .B(n5639), .Z(n4719) );
  XOR U6857 ( .A(round_reg[393]), .B(n5640), .Z(n5639) );
  XOR U6858 ( .A(round_reg[73]), .B(round_reg[713]), .Z(n5640) );
  XNOR U6859 ( .A(round_reg[1033]), .B(round_reg[1353]), .Z(n5638) );
  XOR U6860 ( .A(n5641), .B(n5642), .Z(n5026) );
  XOR U6861 ( .A(round_reg[202]), .B(n5643), .Z(n5642) );
  XOR U6862 ( .A(round_reg[842]), .B(round_reg[522]), .Z(n5643) );
  XNOR U6863 ( .A(round_reg[1162]), .B(round_reg[1482]), .Z(n5641) );
  XNOR U6864 ( .A(n1915), .B(round_reg[1387]), .Z(n1202) );
  XNOR U6865 ( .A(n5644), .B(n5645), .Z(n4921) );
  XOR U6866 ( .A(round_reg[362]), .B(n5646), .Z(n5645) );
  XOR U6867 ( .A(round_reg[682]), .B(round_reg[42]), .Z(n5646) );
  XNOR U6868 ( .A(round_reg[1002]), .B(round_reg[1322]), .Z(n5644) );
  XOR U6869 ( .A(n5647), .B(n5648), .Z(n5381) );
  XOR U6870 ( .A(round_reg[171]), .B(n5649), .Z(n5648) );
  XOR U6871 ( .A(round_reg[811]), .B(round_reg[491]), .Z(n5649) );
  XNOR U6872 ( .A(round_reg[1131]), .B(round_reg[1451]), .Z(n5647) );
  XOR U6873 ( .A(n5650), .B(n4821), .Z(o[1030]) );
  XOR U6874 ( .A(n2281), .B(round_reg[537]), .Z(n4821) );
  XNOR U6875 ( .A(n5651), .B(n5652), .Z(n2281) );
  AND U6876 ( .A(n1206), .B(n1204), .Z(n5650) );
  XNOR U6877 ( .A(n2328), .B(round_reg[137]), .Z(n1204) );
  XNOR U6878 ( .A(n5028), .B(n4722), .Z(n2328) );
  XOR U6879 ( .A(n5653), .B(n5654), .Z(n4722) );
  XOR U6880 ( .A(round_reg[392]), .B(n5655), .Z(n5654) );
  XOR U6881 ( .A(round_reg[72]), .B(round_reg[712]), .Z(n5655) );
  XNOR U6882 ( .A(round_reg[1032]), .B(round_reg[1352]), .Z(n5653) );
  XNOR U6883 ( .A(n5656), .B(n5657), .Z(n5028) );
  XOR U6884 ( .A(round_reg[201]), .B(n5658), .Z(n5657) );
  XOR U6885 ( .A(round_reg[841]), .B(round_reg[521]), .Z(n5658) );
  XNOR U6886 ( .A(round_reg[1161]), .B(round_reg[1481]), .Z(n5656) );
  XNOR U6887 ( .A(n1918), .B(round_reg[1386]), .Z(n1206) );
  XNOR U6888 ( .A(n5659), .B(n5660), .Z(n4925) );
  XOR U6889 ( .A(round_reg[361]), .B(n5661), .Z(n5660) );
  XOR U6890 ( .A(round_reg[681]), .B(round_reg[41]), .Z(n5661) );
  XNOR U6891 ( .A(round_reg[1001]), .B(round_reg[1321]), .Z(n5659) );
  XOR U6892 ( .A(n5662), .B(n5663), .Z(n5392) );
  XOR U6893 ( .A(round_reg[170]), .B(n5664), .Z(n5663) );
  XOR U6894 ( .A(round_reg[810]), .B(round_reg[490]), .Z(n5664) );
  XNOR U6895 ( .A(round_reg[1130]), .B(round_reg[1450]), .Z(n5662) );
  XOR U6896 ( .A(n5665), .B(n3511), .Z(o[102]) );
  XOR U6897 ( .A(n2327), .B(round_reg[637]), .Z(n3511) );
  IV U6898 ( .A(n5067), .Z(n2327) );
  XOR U6899 ( .A(n5666), .B(n5367), .Z(n5067) );
  XOR U6900 ( .A(n5667), .B(n5668), .Z(n5367) );
  XOR U6901 ( .A(round_reg[381]), .B(n5669), .Z(n5668) );
  XOR U6902 ( .A(round_reg[701]), .B(round_reg[61]), .Z(n5669) );
  XNOR U6903 ( .A(round_reg[1021]), .B(round_reg[1341]), .Z(n5667) );
  AND U6904 ( .A(n3171), .B(n3173), .Z(n5665) );
  XOR U6905 ( .A(n2192), .B(round_reg[1448]), .Z(n3173) );
  XOR U6906 ( .A(n4926), .B(n5670), .Z(n2192) );
  XOR U6907 ( .A(n5671), .B(n5672), .Z(n4926) );
  XOR U6908 ( .A(round_reg[232]), .B(n5673), .Z(n5672) );
  XOR U6909 ( .A(round_reg[872]), .B(round_reg[552]), .Z(n5673) );
  XNOR U6910 ( .A(round_reg[1192]), .B(round_reg[1512]), .Z(n5671) );
  XNOR U6911 ( .A(n2233), .B(round_reg[228]), .Z(n3171) );
  XNOR U6912 ( .A(n5674), .B(n5675), .Z(n2233) );
  XOR U6913 ( .A(n5676), .B(n4825), .Z(o[1029]) );
  XOR U6914 ( .A(n2285), .B(round_reg[536]), .Z(n4825) );
  XNOR U6915 ( .A(n5677), .B(n5678), .Z(n2285) );
  ANDN U6916 ( .A(n1208), .B(n1209), .Z(n5676) );
  XOR U6917 ( .A(n1921), .B(round_reg[1385]), .Z(n1209) );
  XNOR U6918 ( .A(n5679), .B(n5680), .Z(n4929) );
  XOR U6919 ( .A(round_reg[360]), .B(n5681), .Z(n5680) );
  XOR U6920 ( .A(round_reg[680]), .B(round_reg[40]), .Z(n5681) );
  XNOR U6921 ( .A(round_reg[1000]), .B(round_reg[1320]), .Z(n5679) );
  XOR U6922 ( .A(n5682), .B(n5683), .Z(n5406) );
  XOR U6923 ( .A(round_reg[169]), .B(n5684), .Z(n5683) );
  XOR U6924 ( .A(round_reg[809]), .B(round_reg[489]), .Z(n5684) );
  XNOR U6925 ( .A(round_reg[1129]), .B(round_reg[1449]), .Z(n5682) );
  XNOR U6926 ( .A(n2332), .B(round_reg[136]), .Z(n1208) );
  XNOR U6927 ( .A(n5031), .B(n4730), .Z(n2332) );
  XOR U6928 ( .A(n5685), .B(n5686), .Z(n4730) );
  XOR U6929 ( .A(round_reg[391]), .B(n5687), .Z(n5686) );
  XOR U6930 ( .A(round_reg[71]), .B(round_reg[711]), .Z(n5687) );
  XNOR U6931 ( .A(round_reg[1031]), .B(round_reg[1351]), .Z(n5685) );
  XNOR U6932 ( .A(n5688), .B(n5689), .Z(n5031) );
  XOR U6933 ( .A(round_reg[200]), .B(n5690), .Z(n5689) );
  XOR U6934 ( .A(round_reg[840]), .B(round_reg[520]), .Z(n5690) );
  XNOR U6935 ( .A(round_reg[1160]), .B(round_reg[1480]), .Z(n5688) );
  XOR U6936 ( .A(n5691), .B(n4829), .Z(o[1028]) );
  XOR U6937 ( .A(n2289), .B(round_reg[535]), .Z(n4829) );
  XNOR U6938 ( .A(n5692), .B(n5693), .Z(n2289) );
  ANDN U6939 ( .A(n1212), .B(n1213), .Z(n5691) );
  XOR U6940 ( .A(n1928), .B(round_reg[1384]), .Z(n1213) );
  XNOR U6941 ( .A(n5694), .B(n5695), .Z(n4933) );
  XOR U6942 ( .A(round_reg[39]), .B(n5696), .Z(n5695) );
  XOR U6943 ( .A(round_reg[999]), .B(round_reg[679]), .Z(n5696) );
  XNOR U6944 ( .A(round_reg[1319]), .B(round_reg[359]), .Z(n5694) );
  XOR U6945 ( .A(n5697), .B(n5698), .Z(n5419) );
  XOR U6946 ( .A(round_reg[168]), .B(n5699), .Z(n5698) );
  XOR U6947 ( .A(round_reg[808]), .B(round_reg[488]), .Z(n5699) );
  XNOR U6948 ( .A(round_reg[1128]), .B(round_reg[1448]), .Z(n5697) );
  XNOR U6949 ( .A(n2336), .B(round_reg[135]), .Z(n1212) );
  XNOR U6950 ( .A(n5037), .B(n4734), .Z(n2336) );
  XOR U6951 ( .A(n5700), .B(n5701), .Z(n4734) );
  XOR U6952 ( .A(round_reg[390]), .B(n5702), .Z(n5701) );
  XOR U6953 ( .A(round_reg[710]), .B(round_reg[70]), .Z(n5702) );
  XNOR U6954 ( .A(round_reg[1030]), .B(round_reg[1350]), .Z(n5700) );
  XNOR U6955 ( .A(n5703), .B(n5704), .Z(n5037) );
  XOR U6956 ( .A(round_reg[199]), .B(n5705), .Z(n5704) );
  XOR U6957 ( .A(round_reg[839]), .B(round_reg[519]), .Z(n5705) );
  XNOR U6958 ( .A(round_reg[1159]), .B(round_reg[1479]), .Z(n5703) );
  XOR U6959 ( .A(n5706), .B(n4833), .Z(o[1027]) );
  XOR U6960 ( .A(n2293), .B(round_reg[534]), .Z(n4833) );
  XNOR U6961 ( .A(n5707), .B(n5708), .Z(n2293) );
  ANDN U6962 ( .A(n1216), .B(n1217), .Z(n5706) );
  XOR U6963 ( .A(n1931), .B(round_reg[1383]), .Z(n1217) );
  XNOR U6964 ( .A(n5709), .B(n5710), .Z(n4939) );
  XOR U6965 ( .A(round_reg[38]), .B(n5711), .Z(n5710) );
  XOR U6966 ( .A(round_reg[998]), .B(round_reg[678]), .Z(n5711) );
  XNOR U6967 ( .A(round_reg[1318]), .B(round_reg[358]), .Z(n5709) );
  XOR U6968 ( .A(n5712), .B(n5713), .Z(n5432) );
  XOR U6969 ( .A(round_reg[167]), .B(n5714), .Z(n5713) );
  XOR U6970 ( .A(round_reg[807]), .B(round_reg[487]), .Z(n5714) );
  XNOR U6971 ( .A(round_reg[1127]), .B(round_reg[1447]), .Z(n5712) );
  XNOR U6972 ( .A(n2340), .B(round_reg[134]), .Z(n1216) );
  XNOR U6973 ( .A(n5040), .B(n4738), .Z(n2340) );
  XOR U6974 ( .A(n5715), .B(n5716), .Z(n4738) );
  XOR U6975 ( .A(round_reg[389]), .B(n5717), .Z(n5716) );
  XOR U6976 ( .A(round_reg[709]), .B(round_reg[69]), .Z(n5717) );
  XNOR U6977 ( .A(round_reg[1029]), .B(round_reg[1349]), .Z(n5715) );
  XNOR U6978 ( .A(n5718), .B(n5719), .Z(n5040) );
  XOR U6979 ( .A(round_reg[198]), .B(n5720), .Z(n5719) );
  XOR U6980 ( .A(round_reg[838]), .B(round_reg[518]), .Z(n5720) );
  XNOR U6981 ( .A(round_reg[1158]), .B(round_reg[1478]), .Z(n5718) );
  XOR U6982 ( .A(n5721), .B(n4837), .Z(o[1026]) );
  XOR U6983 ( .A(n2297), .B(round_reg[533]), .Z(n4837) );
  XNOR U6984 ( .A(n5722), .B(n5723), .Z(n2297) );
  ANDN U6985 ( .A(n1220), .B(n1221), .Z(n5721) );
  XOR U6986 ( .A(n1710), .B(round_reg[1382]), .Z(n1221) );
  XNOR U6987 ( .A(n5724), .B(n5725), .Z(n4943) );
  XOR U6988 ( .A(round_reg[37]), .B(n5726), .Z(n5725) );
  XOR U6989 ( .A(round_reg[997]), .B(round_reg[677]), .Z(n5726) );
  XNOR U6990 ( .A(round_reg[1317]), .B(round_reg[357]), .Z(n5724) );
  XOR U6991 ( .A(n5727), .B(n5728), .Z(n5445) );
  XOR U6992 ( .A(round_reg[166]), .B(n5729), .Z(n5728) );
  XOR U6993 ( .A(round_reg[806]), .B(round_reg[486]), .Z(n5729) );
  XNOR U6994 ( .A(round_reg[1126]), .B(round_reg[1446]), .Z(n5727) );
  XNOR U6995 ( .A(n2344), .B(round_reg[133]), .Z(n1220) );
  XNOR U6996 ( .A(n5043), .B(n4742), .Z(n2344) );
  XOR U6997 ( .A(n5730), .B(n5731), .Z(n4742) );
  XOR U6998 ( .A(round_reg[388]), .B(n5732), .Z(n5731) );
  XOR U6999 ( .A(round_reg[708]), .B(round_reg[68]), .Z(n5732) );
  XNOR U7000 ( .A(round_reg[1028]), .B(round_reg[1348]), .Z(n5730) );
  XNOR U7001 ( .A(n5733), .B(n5734), .Z(n5043) );
  XOR U7002 ( .A(round_reg[197]), .B(n5735), .Z(n5734) );
  XOR U7003 ( .A(round_reg[837]), .B(round_reg[517]), .Z(n5735) );
  XNOR U7004 ( .A(round_reg[1157]), .B(round_reg[1477]), .Z(n5733) );
  XOR U7005 ( .A(n5736), .B(n4841), .Z(o[1025]) );
  XOR U7006 ( .A(n2301), .B(round_reg[532]), .Z(n4841) );
  XNOR U7007 ( .A(n5737), .B(n5738), .Z(n2301) );
  ANDN U7008 ( .A(n1224), .B(n1225), .Z(n5736) );
  XOR U7009 ( .A(n1713), .B(round_reg[1381]), .Z(n1225) );
  XNOR U7010 ( .A(n5739), .B(n5740), .Z(n4947) );
  XOR U7011 ( .A(round_reg[36]), .B(n5741), .Z(n5740) );
  XOR U7012 ( .A(round_reg[996]), .B(round_reg[676]), .Z(n5741) );
  XNOR U7013 ( .A(round_reg[1316]), .B(round_reg[356]), .Z(n5739) );
  XOR U7014 ( .A(n5742), .B(n5743), .Z(n5458) );
  XOR U7015 ( .A(round_reg[165]), .B(n5744), .Z(n5743) );
  XOR U7016 ( .A(round_reg[805]), .B(round_reg[485]), .Z(n5744) );
  XNOR U7017 ( .A(round_reg[1125]), .B(round_reg[1445]), .Z(n5742) );
  XNOR U7018 ( .A(n2348), .B(round_reg[132]), .Z(n1224) );
  XNOR U7019 ( .A(n5046), .B(n4746), .Z(n2348) );
  XOR U7020 ( .A(n5745), .B(n5746), .Z(n4746) );
  XOR U7021 ( .A(round_reg[387]), .B(n5747), .Z(n5746) );
  XOR U7022 ( .A(round_reg[707]), .B(round_reg[67]), .Z(n5747) );
  XNOR U7023 ( .A(round_reg[1027]), .B(round_reg[1347]), .Z(n5745) );
  XNOR U7024 ( .A(n5748), .B(n5749), .Z(n5046) );
  XOR U7025 ( .A(round_reg[196]), .B(n5750), .Z(n5749) );
  XOR U7026 ( .A(round_reg[836]), .B(round_reg[516]), .Z(n5750) );
  XNOR U7027 ( .A(round_reg[1156]), .B(round_reg[1476]), .Z(n5748) );
  XOR U7028 ( .A(n5751), .B(n4845), .Z(o[1024]) );
  XOR U7029 ( .A(n2305), .B(round_reg[531]), .Z(n4845) );
  XNOR U7030 ( .A(n5752), .B(n5753), .Z(n2305) );
  ANDN U7031 ( .A(n1228), .B(n1229), .Z(n5751) );
  XOR U7032 ( .A(n1720), .B(round_reg[1380]), .Z(n1229) );
  XNOR U7033 ( .A(n5754), .B(n5755), .Z(n4950) );
  XOR U7034 ( .A(round_reg[35]), .B(n5756), .Z(n5755) );
  XOR U7035 ( .A(round_reg[995]), .B(round_reg[675]), .Z(n5756) );
  XNOR U7036 ( .A(round_reg[1315]), .B(round_reg[355]), .Z(n5754) );
  XOR U7037 ( .A(n5757), .B(n5758), .Z(n5516) );
  XOR U7038 ( .A(round_reg[164]), .B(n5759), .Z(n5758) );
  XOR U7039 ( .A(round_reg[804]), .B(round_reg[484]), .Z(n5759) );
  XNOR U7040 ( .A(round_reg[1124]), .B(round_reg[1444]), .Z(n5757) );
  XNOR U7041 ( .A(n2356), .B(round_reg[131]), .Z(n1228) );
  XNOR U7042 ( .A(n5049), .B(n4750), .Z(n2356) );
  XOR U7043 ( .A(n5760), .B(n5761), .Z(n4750) );
  XOR U7044 ( .A(round_reg[386]), .B(n5762), .Z(n5761) );
  XOR U7045 ( .A(round_reg[706]), .B(round_reg[66]), .Z(n5762) );
  XNOR U7046 ( .A(round_reg[1026]), .B(round_reg[1346]), .Z(n5760) );
  XNOR U7047 ( .A(n5763), .B(n5764), .Z(n5049) );
  XOR U7048 ( .A(round_reg[195]), .B(n5765), .Z(n5764) );
  XOR U7049 ( .A(round_reg[835]), .B(round_reg[515]), .Z(n5765) );
  XNOR U7050 ( .A(round_reg[1155]), .B(round_reg[1475]), .Z(n5763) );
  XOR U7051 ( .A(n5766), .B(n4848), .Z(o[1023]) );
  XOR U7052 ( .A(n2360), .B(round_reg[130]), .Z(n4848) );
  ANDN U7053 ( .A(n4424), .B(n4422), .Z(n5766) );
  XNOR U7054 ( .A(n1723), .B(round_reg[1379]), .Z(n4422) );
  XNOR U7055 ( .A(n5767), .B(n5768), .Z(n4953) );
  XOR U7056 ( .A(round_reg[354]), .B(n5769), .Z(n5768) );
  XOR U7057 ( .A(round_reg[994]), .B(round_reg[674]), .Z(n5769) );
  XNOR U7058 ( .A(round_reg[1314]), .B(round_reg[34]), .Z(n5767) );
  XOR U7059 ( .A(n5770), .B(n5771), .Z(n5675) );
  XOR U7060 ( .A(round_reg[163]), .B(n5772), .Z(n5771) );
  XOR U7061 ( .A(round_reg[803]), .B(round_reg[483]), .Z(n5772) );
  XNOR U7062 ( .A(round_reg[1123]), .B(round_reg[1443]), .Z(n5770) );
  XOR U7063 ( .A(n1971), .B(round_reg[1003]), .Z(n4424) );
  XNOR U7064 ( .A(n5405), .B(n5773), .Z(n1971) );
  XNOR U7065 ( .A(n5774), .B(n5775), .Z(n5405) );
  XOR U7066 ( .A(round_reg[298]), .B(n5776), .Z(n5775) );
  XOR U7067 ( .A(round_reg[938]), .B(round_reg[618]), .Z(n5776) );
  XNOR U7068 ( .A(round_reg[1258]), .B(round_reg[1578]), .Z(n5774) );
  XOR U7069 ( .A(n5777), .B(n4851), .Z(o[1022]) );
  XOR U7070 ( .A(n2364), .B(round_reg[129]), .Z(n4851) );
  XNOR U7071 ( .A(n5109), .B(n4758), .Z(n2364) );
  XOR U7072 ( .A(n5778), .B(n5779), .Z(n4758) );
  XOR U7073 ( .A(round_reg[384]), .B(n5780), .Z(n5779) );
  XOR U7074 ( .A(round_reg[704]), .B(round_reg[64]), .Z(n5780) );
  XNOR U7075 ( .A(round_reg[1024]), .B(round_reg[1344]), .Z(n5778) );
  XNOR U7076 ( .A(n5781), .B(n5782), .Z(n5109) );
  XOR U7077 ( .A(round_reg[193]), .B(n5783), .Z(n5782) );
  XOR U7078 ( .A(round_reg[833]), .B(round_reg[513]), .Z(n5783) );
  XNOR U7079 ( .A(round_reg[1153]), .B(round_reg[1473]), .Z(n5781) );
  ANDN U7080 ( .A(n4428), .B(n4426), .Z(n5777) );
  XNOR U7081 ( .A(n1726), .B(round_reg[1378]), .Z(n4426) );
  XNOR U7082 ( .A(n5785), .B(n5786), .Z(n4956) );
  XOR U7083 ( .A(round_reg[353]), .B(n5787), .Z(n5786) );
  XOR U7084 ( .A(round_reg[993]), .B(round_reg[673]), .Z(n5787) );
  XNOR U7085 ( .A(round_reg[1313]), .B(round_reg[33]), .Z(n5785) );
  XOR U7086 ( .A(n1974), .B(round_reg[1002]), .Z(n4428) );
  XNOR U7087 ( .A(n5418), .B(n5788), .Z(n1974) );
  XNOR U7088 ( .A(n5789), .B(n5790), .Z(n5418) );
  XOR U7089 ( .A(round_reg[297]), .B(n5791), .Z(n5790) );
  XOR U7090 ( .A(round_reg[937]), .B(round_reg[617]), .Z(n5791) );
  XNOR U7091 ( .A(round_reg[1257]), .B(round_reg[1577]), .Z(n5789) );
  XOR U7092 ( .A(n5792), .B(n4857), .Z(o[1021]) );
  XOR U7093 ( .A(n2368), .B(round_reg[128]), .Z(n4857) );
  XNOR U7094 ( .A(n5162), .B(n4761), .Z(n2368) );
  XOR U7095 ( .A(n5793), .B(n5794), .Z(n4761) );
  XOR U7096 ( .A(round_reg[1407]), .B(n5795), .Z(n5794) );
  XOR U7097 ( .A(round_reg[767]), .B(round_reg[447]), .Z(n5795) );
  XNOR U7098 ( .A(round_reg[1087]), .B(round_reg[127]), .Z(n5793) );
  XNOR U7099 ( .A(n5796), .B(n5797), .Z(n5162) );
  XOR U7100 ( .A(round_reg[192]), .B(n5798), .Z(n5797) );
  XOR U7101 ( .A(round_reg[832]), .B(round_reg[512]), .Z(n5798) );
  XNOR U7102 ( .A(round_reg[1152]), .B(round_reg[1472]), .Z(n5796) );
  ANDN U7103 ( .A(n4432), .B(n4430), .Z(n5792) );
  XNOR U7104 ( .A(n1729), .B(round_reg[1377]), .Z(n4430) );
  XNOR U7105 ( .A(n5800), .B(n5801), .Z(n4959) );
  XOR U7106 ( .A(round_reg[352]), .B(n5802), .Z(n5801) );
  XOR U7107 ( .A(round_reg[992]), .B(round_reg[672]), .Z(n5802) );
  XNOR U7108 ( .A(round_reg[1312]), .B(round_reg[32]), .Z(n5800) );
  XNOR U7109 ( .A(n4313), .B(round_reg[1001]), .Z(n4432) );
  XOR U7110 ( .A(n5431), .B(n5376), .Z(n4313) );
  XOR U7111 ( .A(n5803), .B(n5804), .Z(n5376) );
  XOR U7112 ( .A(round_reg[1385]), .B(n5805), .Z(n5804) );
  XOR U7113 ( .A(round_reg[745]), .B(round_reg[425]), .Z(n5805) );
  XNOR U7114 ( .A(round_reg[105]), .B(round_reg[1065]), .Z(n5803) );
  XNOR U7115 ( .A(n5806), .B(n5807), .Z(n5431) );
  XOR U7116 ( .A(round_reg[296]), .B(n5808), .Z(n5807) );
  XOR U7117 ( .A(round_reg[936]), .B(round_reg[616]), .Z(n5808) );
  XNOR U7118 ( .A(round_reg[1256]), .B(round_reg[1576]), .Z(n5806) );
  XOR U7119 ( .A(n5809), .B(n4861), .Z(o[1020]) );
  XOR U7120 ( .A(n2372), .B(round_reg[191]), .Z(n4861) );
  XNOR U7121 ( .A(n5229), .B(n4766), .Z(n2372) );
  XOR U7122 ( .A(n5810), .B(n5811), .Z(n4766) );
  XOR U7123 ( .A(round_reg[1406]), .B(n5812), .Z(n5811) );
  XOR U7124 ( .A(round_reg[766]), .B(round_reg[446]), .Z(n5812) );
  XNOR U7125 ( .A(round_reg[1086]), .B(round_reg[126]), .Z(n5810) );
  XNOR U7126 ( .A(n5813), .B(n5814), .Z(n5229) );
  XOR U7127 ( .A(round_reg[255]), .B(n5815), .Z(n5814) );
  XOR U7128 ( .A(round_reg[895]), .B(round_reg[575]), .Z(n5815) );
  XNOR U7129 ( .A(round_reg[1215]), .B(round_reg[1535]), .Z(n5813) );
  ANDN U7130 ( .A(n4436), .B(n4434), .Z(n5809) );
  XOR U7131 ( .A(n1732), .B(round_reg[1376]), .Z(n4434) );
  XNOR U7132 ( .A(n4962), .B(n5532), .Z(n1732) );
  XOR U7133 ( .A(n5816), .B(n5817), .Z(n5532) );
  XOR U7134 ( .A(round_reg[160]), .B(n5818), .Z(n5817) );
  XOR U7135 ( .A(round_reg[800]), .B(round_reg[480]), .Z(n5818) );
  XNOR U7136 ( .A(round_reg[1120]), .B(round_reg[1440]), .Z(n5816) );
  XNOR U7137 ( .A(n5819), .B(n5820), .Z(n4962) );
  XOR U7138 ( .A(round_reg[351]), .B(n5821), .Z(n5820) );
  XOR U7139 ( .A(round_reg[991]), .B(round_reg[671]), .Z(n5821) );
  XNOR U7140 ( .A(round_reg[1311]), .B(round_reg[31]), .Z(n5819) );
  XNOR U7141 ( .A(n4315), .B(round_reg[1000]), .Z(n4436) );
  XOR U7142 ( .A(n5444), .B(n5511), .Z(n4315) );
  XOR U7143 ( .A(n5822), .B(n5823), .Z(n5511) );
  XOR U7144 ( .A(round_reg[1384]), .B(n5824), .Z(n5823) );
  XOR U7145 ( .A(round_reg[744]), .B(round_reg[424]), .Z(n5824) );
  XNOR U7146 ( .A(round_reg[104]), .B(round_reg[1064]), .Z(n5822) );
  XNOR U7147 ( .A(n5825), .B(n5826), .Z(n5444) );
  XOR U7148 ( .A(round_reg[295]), .B(n5827), .Z(n5826) );
  XOR U7149 ( .A(round_reg[935]), .B(round_reg[615]), .Z(n5827) );
  XNOR U7150 ( .A(round_reg[1255]), .B(round_reg[1575]), .Z(n5825) );
  XOR U7151 ( .A(n5828), .B(n3514), .Z(o[101]) );
  XOR U7152 ( .A(n2331), .B(round_reg[636]), .Z(n3514) );
  IV U7153 ( .A(n4847), .Z(n2331) );
  XOR U7154 ( .A(n5829), .B(n5390), .Z(n4847) );
  XOR U7155 ( .A(n5830), .B(n5831), .Z(n5390) );
  XOR U7156 ( .A(round_reg[380]), .B(n5832), .Z(n5831) );
  XOR U7157 ( .A(round_reg[700]), .B(round_reg[60]), .Z(n5832) );
  XNOR U7158 ( .A(round_reg[1020]), .B(round_reg[1340]), .Z(n5830) );
  AND U7159 ( .A(n3185), .B(n3187), .Z(n5828) );
  XOR U7160 ( .A(n2196), .B(round_reg[1447]), .Z(n3187) );
  XOR U7161 ( .A(n4930), .B(n5833), .Z(n2196) );
  XOR U7162 ( .A(n5834), .B(n5835), .Z(n4930) );
  XOR U7163 ( .A(round_reg[231]), .B(n5836), .Z(n5835) );
  XOR U7164 ( .A(round_reg[871]), .B(round_reg[551]), .Z(n5836) );
  XNOR U7165 ( .A(round_reg[1191]), .B(round_reg[1511]), .Z(n5834) );
  XNOR U7166 ( .A(n2237), .B(round_reg[227]), .Z(n3185) );
  XNOR U7167 ( .A(n5837), .B(n5784), .Z(n2237) );
  XOR U7168 ( .A(n5838), .B(n5839), .Z(n5784) );
  XOR U7169 ( .A(round_reg[162]), .B(n5840), .Z(n5839) );
  XOR U7170 ( .A(round_reg[802]), .B(round_reg[482]), .Z(n5840) );
  XNOR U7171 ( .A(round_reg[1122]), .B(round_reg[1442]), .Z(n5838) );
  XOR U7172 ( .A(n5841), .B(n4865), .Z(o[1019]) );
  XOR U7173 ( .A(n2376), .B(round_reg[190]), .Z(n4865) );
  XNOR U7174 ( .A(n5372), .B(n4773), .Z(n2376) );
  XOR U7175 ( .A(n5842), .B(n5843), .Z(n4773) );
  XOR U7176 ( .A(round_reg[1405]), .B(n5844), .Z(n5843) );
  XOR U7177 ( .A(round_reg[765]), .B(round_reg[445]), .Z(n5844) );
  XNOR U7178 ( .A(round_reg[1085]), .B(round_reg[125]), .Z(n5842) );
  XNOR U7179 ( .A(n5845), .B(n5846), .Z(n5372) );
  XOR U7180 ( .A(round_reg[254]), .B(n5847), .Z(n5846) );
  XOR U7181 ( .A(round_reg[894]), .B(round_reg[574]), .Z(n5847) );
  XNOR U7182 ( .A(round_reg[1214]), .B(round_reg[1534]), .Z(n5845) );
  ANDN U7183 ( .A(n4440), .B(n4438), .Z(n5841) );
  XOR U7184 ( .A(n1735), .B(round_reg[1375]), .Z(n4438) );
  XNOR U7185 ( .A(n4965), .B(n5546), .Z(n1735) );
  XOR U7186 ( .A(n5848), .B(n5849), .Z(n5546) );
  XOR U7187 ( .A(round_reg[159]), .B(n5850), .Z(n5849) );
  XOR U7188 ( .A(round_reg[799]), .B(round_reg[479]), .Z(n5850) );
  XNOR U7189 ( .A(round_reg[1119]), .B(round_reg[1439]), .Z(n5848) );
  XNOR U7190 ( .A(n5851), .B(n5852), .Z(n4965) );
  XOR U7191 ( .A(round_reg[350]), .B(n5853), .Z(n5852) );
  XOR U7192 ( .A(round_reg[990]), .B(round_reg[670]), .Z(n5853) );
  XNOR U7193 ( .A(round_reg[1310]), .B(round_reg[30]), .Z(n5851) );
  XNOR U7194 ( .A(n4317), .B(round_reg[999]), .Z(n4440) );
  XOR U7195 ( .A(n5457), .B(n5670), .Z(n4317) );
  XOR U7196 ( .A(n5854), .B(n5855), .Z(n5670) );
  XOR U7197 ( .A(round_reg[1383]), .B(n5856), .Z(n5855) );
  XOR U7198 ( .A(round_reg[743]), .B(round_reg[423]), .Z(n5856) );
  XNOR U7199 ( .A(round_reg[103]), .B(round_reg[1063]), .Z(n5854) );
  XNOR U7200 ( .A(n5857), .B(n5858), .Z(n5457) );
  XOR U7201 ( .A(round_reg[294]), .B(n5859), .Z(n5858) );
  XOR U7202 ( .A(round_reg[934]), .B(round_reg[614]), .Z(n5859) );
  XNOR U7203 ( .A(round_reg[1254]), .B(round_reg[1574]), .Z(n5857) );
  XOR U7204 ( .A(n5860), .B(n4869), .Z(o[1018]) );
  XOR U7205 ( .A(n2380), .B(round_reg[189]), .Z(n4869) );
  XNOR U7206 ( .A(n5507), .B(n4777), .Z(n2380) );
  XOR U7207 ( .A(n5861), .B(n5862), .Z(n4777) );
  XOR U7208 ( .A(round_reg[1404]), .B(n5863), .Z(n5862) );
  XOR U7209 ( .A(round_reg[764]), .B(round_reg[444]), .Z(n5863) );
  XNOR U7210 ( .A(round_reg[1084]), .B(round_reg[124]), .Z(n5861) );
  XNOR U7211 ( .A(n5864), .B(n5865), .Z(n5507) );
  XOR U7212 ( .A(round_reg[253]), .B(n5866), .Z(n5865) );
  XOR U7213 ( .A(round_reg[893]), .B(round_reg[573]), .Z(n5866) );
  XNOR U7214 ( .A(round_reg[1213]), .B(round_reg[1533]), .Z(n5864) );
  ANDN U7215 ( .A(n4444), .B(n4442), .Z(n5860) );
  XOR U7216 ( .A(n1738), .B(round_reg[1374]), .Z(n4442) );
  XNOR U7217 ( .A(n4968), .B(n5561), .Z(n1738) );
  XOR U7218 ( .A(n5867), .B(n5868), .Z(n5561) );
  XOR U7219 ( .A(round_reg[158]), .B(n5869), .Z(n5868) );
  XOR U7220 ( .A(round_reg[798]), .B(round_reg[478]), .Z(n5869) );
  XNOR U7221 ( .A(round_reg[1118]), .B(round_reg[1438]), .Z(n5867) );
  XNOR U7222 ( .A(n5870), .B(n5871), .Z(n4968) );
  XOR U7223 ( .A(round_reg[349]), .B(n5872), .Z(n5871) );
  XOR U7224 ( .A(round_reg[989]), .B(round_reg[669]), .Z(n5872) );
  XNOR U7225 ( .A(round_reg[1309]), .B(round_reg[29]), .Z(n5870) );
  XNOR U7226 ( .A(n4320), .B(round_reg[998]), .Z(n4444) );
  XOR U7227 ( .A(n5515), .B(n5833), .Z(n4320) );
  XOR U7228 ( .A(n5873), .B(n5874), .Z(n5833) );
  XOR U7229 ( .A(round_reg[1382]), .B(n5875), .Z(n5874) );
  XOR U7230 ( .A(round_reg[742]), .B(round_reg[422]), .Z(n5875) );
  XNOR U7231 ( .A(round_reg[102]), .B(round_reg[1062]), .Z(n5873) );
  XNOR U7232 ( .A(n5876), .B(n5877), .Z(n5515) );
  XOR U7233 ( .A(round_reg[293]), .B(n5878), .Z(n5877) );
  XOR U7234 ( .A(round_reg[933]), .B(round_reg[613]), .Z(n5878) );
  XNOR U7235 ( .A(round_reg[1253]), .B(round_reg[1573]), .Z(n5876) );
  XOR U7236 ( .A(n5879), .B(n4873), .Z(o[1017]) );
  XOR U7237 ( .A(n2384), .B(round_reg[188]), .Z(n4873) );
  XNOR U7238 ( .A(n5666), .B(n4781), .Z(n2384) );
  XOR U7239 ( .A(n5880), .B(n5881), .Z(n4781) );
  XOR U7240 ( .A(round_reg[1403]), .B(n5882), .Z(n5881) );
  XOR U7241 ( .A(round_reg[763]), .B(round_reg[443]), .Z(n5882) );
  XNOR U7242 ( .A(round_reg[1083]), .B(round_reg[123]), .Z(n5880) );
  XNOR U7243 ( .A(n5883), .B(n5884), .Z(n5666) );
  XOR U7244 ( .A(round_reg[252]), .B(n5885), .Z(n5884) );
  XOR U7245 ( .A(round_reg[892]), .B(round_reg[572]), .Z(n5885) );
  XNOR U7246 ( .A(round_reg[1212]), .B(round_reg[1532]), .Z(n5883) );
  ANDN U7247 ( .A(n4448), .B(n4446), .Z(n5879) );
  XOR U7248 ( .A(n1741), .B(round_reg[1373]), .Z(n4446) );
  XNOR U7249 ( .A(n4973), .B(n5576), .Z(n1741) );
  XOR U7250 ( .A(n5886), .B(n5887), .Z(n5576) );
  XOR U7251 ( .A(round_reg[157]), .B(n5888), .Z(n5887) );
  XOR U7252 ( .A(round_reg[797]), .B(round_reg[477]), .Z(n5888) );
  XNOR U7253 ( .A(round_reg[1117]), .B(round_reg[1437]), .Z(n5886) );
  XNOR U7254 ( .A(n5889), .B(n5890), .Z(n4973) );
  XOR U7255 ( .A(round_reg[348]), .B(n5891), .Z(n5890) );
  XOR U7256 ( .A(round_reg[988]), .B(round_reg[668]), .Z(n5891) );
  XNOR U7257 ( .A(round_reg[1308]), .B(round_reg[28]), .Z(n5889) );
  XNOR U7258 ( .A(n4323), .B(round_reg[997]), .Z(n4448) );
  XOR U7259 ( .A(n5674), .B(n5892), .Z(n4323) );
  XNOR U7260 ( .A(n5893), .B(n5894), .Z(n5674) );
  XOR U7261 ( .A(round_reg[292]), .B(n5895), .Z(n5894) );
  XOR U7262 ( .A(round_reg[932]), .B(round_reg[612]), .Z(n5895) );
  XNOR U7263 ( .A(round_reg[1252]), .B(round_reg[1572]), .Z(n5893) );
  XOR U7264 ( .A(n5896), .B(n4877), .Z(o[1016]) );
  XOR U7265 ( .A(n2388), .B(round_reg[187]), .Z(n4877) );
  XNOR U7266 ( .A(n5829), .B(n4785), .Z(n2388) );
  XOR U7267 ( .A(n5897), .B(n5898), .Z(n4785) );
  XOR U7268 ( .A(round_reg[1402]), .B(n5899), .Z(n5898) );
  XOR U7269 ( .A(round_reg[762]), .B(round_reg[442]), .Z(n5899) );
  XNOR U7270 ( .A(round_reg[1082]), .B(round_reg[122]), .Z(n5897) );
  XNOR U7271 ( .A(n5900), .B(n5901), .Z(n5829) );
  XOR U7272 ( .A(round_reg[251]), .B(n5902), .Z(n5901) );
  XOR U7273 ( .A(round_reg[891]), .B(round_reg[571]), .Z(n5902) );
  XNOR U7274 ( .A(round_reg[1211]), .B(round_reg[1531]), .Z(n5900) );
  ANDN U7275 ( .A(n4452), .B(n4450), .Z(n5896) );
  XOR U7276 ( .A(n1744), .B(round_reg[1372]), .Z(n4450) );
  XNOR U7277 ( .A(n4976), .B(n5591), .Z(n1744) );
  XOR U7278 ( .A(n5903), .B(n5904), .Z(n5591) );
  XOR U7279 ( .A(round_reg[156]), .B(n5905), .Z(n5904) );
  XOR U7280 ( .A(round_reg[796]), .B(round_reg[476]), .Z(n5905) );
  XNOR U7281 ( .A(round_reg[1116]), .B(round_reg[1436]), .Z(n5903) );
  XNOR U7282 ( .A(n5906), .B(n5907), .Z(n4976) );
  XOR U7283 ( .A(round_reg[347]), .B(n5908), .Z(n5907) );
  XOR U7284 ( .A(round_reg[987]), .B(round_reg[667]), .Z(n5908) );
  XNOR U7285 ( .A(round_reg[1307]), .B(round_reg[27]), .Z(n5906) );
  XNOR U7286 ( .A(n4326), .B(round_reg[996]), .Z(n4452) );
  XOR U7287 ( .A(n5837), .B(n5247), .Z(n4326) );
  XOR U7288 ( .A(n5909), .B(n5910), .Z(n5247) );
  XOR U7289 ( .A(round_reg[1380]), .B(n5911), .Z(n5910) );
  XOR U7290 ( .A(round_reg[740]), .B(round_reg[420]), .Z(n5911) );
  XNOR U7291 ( .A(round_reg[100]), .B(round_reg[1060]), .Z(n5909) );
  XNOR U7292 ( .A(n5912), .B(n5913), .Z(n5837) );
  XOR U7293 ( .A(round_reg[291]), .B(n5914), .Z(n5913) );
  XOR U7294 ( .A(round_reg[931]), .B(round_reg[611]), .Z(n5914) );
  XNOR U7295 ( .A(round_reg[1251]), .B(round_reg[1571]), .Z(n5912) );
  XOR U7296 ( .A(n5915), .B(n4881), .Z(o[1015]) );
  XOR U7297 ( .A(n2392), .B(round_reg[186]), .Z(n4881) );
  XNOR U7298 ( .A(n5916), .B(n4789), .Z(n2392) );
  XOR U7299 ( .A(n5917), .B(n5918), .Z(n4789) );
  XOR U7300 ( .A(round_reg[1401]), .B(n5919), .Z(n5918) );
  XOR U7301 ( .A(round_reg[761]), .B(round_reg[441]), .Z(n5919) );
  XNOR U7302 ( .A(round_reg[1081]), .B(round_reg[121]), .Z(n5917) );
  ANDN U7303 ( .A(n4456), .B(n4454), .Z(n5915) );
  XOR U7304 ( .A(n1747), .B(round_reg[1371]), .Z(n4454) );
  XNOR U7305 ( .A(n4979), .B(n5606), .Z(n1747) );
  XOR U7306 ( .A(n5920), .B(n5921), .Z(n5606) );
  XOR U7307 ( .A(round_reg[155]), .B(n5922), .Z(n5921) );
  XOR U7308 ( .A(round_reg[795]), .B(round_reg[475]), .Z(n5922) );
  XNOR U7309 ( .A(round_reg[1115]), .B(round_reg[1435]), .Z(n5920) );
  XNOR U7310 ( .A(n5923), .B(n5924), .Z(n4979) );
  XOR U7311 ( .A(round_reg[346]), .B(n5925), .Z(n5924) );
  XOR U7312 ( .A(round_reg[986]), .B(round_reg[666]), .Z(n5925) );
  XNOR U7313 ( .A(round_reg[1306]), .B(round_reg[26]), .Z(n5923) );
  XNOR U7314 ( .A(n4331), .B(round_reg[995]), .Z(n4456) );
  XOR U7315 ( .A(n5926), .B(n5262), .Z(n4331) );
  XOR U7316 ( .A(n5927), .B(n5928), .Z(n5262) );
  XOR U7317 ( .A(round_reg[419]), .B(n5929), .Z(n5928) );
  XOR U7318 ( .A(round_reg[99]), .B(round_reg[739]), .Z(n5929) );
  XNOR U7319 ( .A(round_reg[1059]), .B(round_reg[1379]), .Z(n5927) );
  XOR U7320 ( .A(n5930), .B(n4885), .Z(o[1014]) );
  XNOR U7321 ( .A(n4657), .B(round_reg[185]), .Z(n4885) );
  XOR U7322 ( .A(n4793), .B(n4855), .Z(n4657) );
  XOR U7323 ( .A(n5931), .B(n5932), .Z(n4855) );
  XOR U7324 ( .A(round_reg[249]), .B(n5933), .Z(n5932) );
  XOR U7325 ( .A(round_reg[889]), .B(round_reg[569]), .Z(n5933) );
  XNOR U7326 ( .A(round_reg[1209]), .B(round_reg[1529]), .Z(n5931) );
  XNOR U7327 ( .A(n5934), .B(n5935), .Z(n4793) );
  XOR U7328 ( .A(round_reg[1400]), .B(n5936), .Z(n5935) );
  XOR U7329 ( .A(round_reg[760]), .B(round_reg[440]), .Z(n5936) );
  XNOR U7330 ( .A(round_reg[1080]), .B(round_reg[120]), .Z(n5934) );
  ANDN U7331 ( .A(n4460), .B(n4458), .Z(n5930) );
  XNOR U7332 ( .A(n1754), .B(round_reg[1370]), .Z(n4458) );
  XNOR U7333 ( .A(n5937), .B(n5938), .Z(n4982) );
  XOR U7334 ( .A(round_reg[345]), .B(n5939), .Z(n5938) );
  XOR U7335 ( .A(round_reg[985]), .B(round_reg[665]), .Z(n5939) );
  XNOR U7336 ( .A(round_reg[1305]), .B(round_reg[25]), .Z(n5937) );
  XOR U7337 ( .A(n5940), .B(n5941), .Z(n5622) );
  XOR U7338 ( .A(round_reg[154]), .B(n5942), .Z(n5941) );
  XOR U7339 ( .A(round_reg[794]), .B(round_reg[474]), .Z(n5942) );
  XNOR U7340 ( .A(round_reg[1114]), .B(round_reg[1434]), .Z(n5940) );
  XNOR U7341 ( .A(n4334), .B(round_reg[994]), .Z(n4460) );
  XOR U7342 ( .A(n5277), .B(n5531), .Z(n4334) );
  XOR U7343 ( .A(n5943), .B(n5944), .Z(n5531) );
  XOR U7344 ( .A(round_reg[289]), .B(n5945), .Z(n5944) );
  XOR U7345 ( .A(round_reg[929]), .B(round_reg[609]), .Z(n5945) );
  XNOR U7346 ( .A(round_reg[1249]), .B(round_reg[1569]), .Z(n5943) );
  XNOR U7347 ( .A(n5946), .B(n5947), .Z(n5277) );
  XOR U7348 ( .A(round_reg[418]), .B(n5948), .Z(n5947) );
  XOR U7349 ( .A(round_reg[98]), .B(round_reg[738]), .Z(n5948) );
  XNOR U7350 ( .A(round_reg[1058]), .B(round_reg[1378]), .Z(n5946) );
  XOR U7351 ( .A(n5949), .B(n4889), .Z(o[1013]) );
  XNOR U7352 ( .A(n4684), .B(round_reg[184]), .Z(n4889) );
  XOR U7353 ( .A(n4797), .B(n4859), .Z(n4684) );
  XOR U7354 ( .A(n5950), .B(n5951), .Z(n4859) );
  XOR U7355 ( .A(round_reg[248]), .B(n5952), .Z(n5951) );
  XOR U7356 ( .A(round_reg[888]), .B(round_reg[568]), .Z(n5952) );
  XNOR U7357 ( .A(round_reg[1208]), .B(round_reg[1528]), .Z(n5950) );
  XNOR U7358 ( .A(n5953), .B(n5954), .Z(n4797) );
  XOR U7359 ( .A(round_reg[1399]), .B(n5955), .Z(n5954) );
  XOR U7360 ( .A(round_reg[759]), .B(round_reg[439]), .Z(n5955) );
  XNOR U7361 ( .A(round_reg[1079]), .B(round_reg[119]), .Z(n5953) );
  ANDN U7362 ( .A(n4466), .B(n4464), .Z(n5949) );
  XNOR U7363 ( .A(n1757), .B(round_reg[1369]), .Z(n4464) );
  XNOR U7364 ( .A(n5956), .B(n5957), .Z(n4985) );
  XOR U7365 ( .A(round_reg[344]), .B(n5958), .Z(n5957) );
  XOR U7366 ( .A(round_reg[984]), .B(round_reg[664]), .Z(n5958) );
  XNOR U7367 ( .A(round_reg[1304]), .B(round_reg[24]), .Z(n5956) );
  XOR U7368 ( .A(n5959), .B(n5960), .Z(n5637) );
  XOR U7369 ( .A(round_reg[153]), .B(n5961), .Z(n5960) );
  XOR U7370 ( .A(round_reg[793]), .B(round_reg[473]), .Z(n5961) );
  XNOR U7371 ( .A(round_reg[1113]), .B(round_reg[1433]), .Z(n5959) );
  XNOR U7372 ( .A(n4271), .B(round_reg[993]), .Z(n4466) );
  XOR U7373 ( .A(n5547), .B(n5292), .Z(n4271) );
  XOR U7374 ( .A(n5962), .B(n5963), .Z(n5292) );
  XOR U7375 ( .A(round_reg[417]), .B(n5964), .Z(n5963) );
  XOR U7376 ( .A(round_reg[97]), .B(round_reg[737]), .Z(n5964) );
  XNOR U7377 ( .A(round_reg[1057]), .B(round_reg[1377]), .Z(n5962) );
  XNOR U7378 ( .A(n5965), .B(n5966), .Z(n5547) );
  XOR U7379 ( .A(round_reg[288]), .B(n5967), .Z(n5966) );
  XOR U7380 ( .A(round_reg[928]), .B(round_reg[608]), .Z(n5967) );
  XNOR U7381 ( .A(round_reg[1248]), .B(round_reg[1568]), .Z(n5965) );
  XOR U7382 ( .A(n5968), .B(n4893), .Z(o[1012]) );
  XNOR U7383 ( .A(n4727), .B(round_reg[183]), .Z(n4893) );
  XOR U7384 ( .A(n4801), .B(n4863), .Z(n4727) );
  XOR U7385 ( .A(n5969), .B(n5970), .Z(n4863) );
  XOR U7386 ( .A(round_reg[247]), .B(n5971), .Z(n5970) );
  XOR U7387 ( .A(round_reg[887]), .B(round_reg[567]), .Z(n5971) );
  XNOR U7388 ( .A(round_reg[1207]), .B(round_reg[1527]), .Z(n5969) );
  XNOR U7389 ( .A(n5972), .B(n5973), .Z(n4801) );
  XOR U7390 ( .A(round_reg[1398]), .B(n5974), .Z(n5973) );
  XOR U7391 ( .A(round_reg[758]), .B(round_reg[438]), .Z(n5974) );
  XNOR U7392 ( .A(round_reg[1078]), .B(round_reg[118]), .Z(n5972) );
  ANDN U7393 ( .A(n4470), .B(n4468), .Z(n5968) );
  XNOR U7394 ( .A(n1760), .B(round_reg[1368]), .Z(n4468) );
  XNOR U7395 ( .A(n5975), .B(n5976), .Z(n4988) );
  XOR U7396 ( .A(round_reg[343]), .B(n5977), .Z(n5976) );
  XOR U7397 ( .A(round_reg[983]), .B(round_reg[663]), .Z(n5977) );
  XNOR U7398 ( .A(round_reg[1303]), .B(round_reg[23]), .Z(n5975) );
  XOR U7399 ( .A(n5978), .B(n5979), .Z(n5652) );
  XOR U7400 ( .A(round_reg[152]), .B(n5980), .Z(n5979) );
  XOR U7401 ( .A(round_reg[792]), .B(round_reg[472]), .Z(n5980) );
  XNOR U7402 ( .A(round_reg[1112]), .B(round_reg[1432]), .Z(n5978) );
  XNOR U7403 ( .A(n4283), .B(round_reg[992]), .Z(n4470) );
  XOR U7404 ( .A(n5562), .B(n5307), .Z(n4283) );
  XOR U7405 ( .A(n5981), .B(n5982), .Z(n5307) );
  XOR U7406 ( .A(round_reg[416]), .B(n5983), .Z(n5982) );
  XOR U7407 ( .A(round_reg[96]), .B(round_reg[736]), .Z(n5983) );
  XNOR U7408 ( .A(round_reg[1056]), .B(round_reg[1376]), .Z(n5981) );
  XNOR U7409 ( .A(n5984), .B(n5985), .Z(n5562) );
  XOR U7410 ( .A(round_reg[287]), .B(n5986), .Z(n5985) );
  XOR U7411 ( .A(round_reg[927]), .B(round_reg[607]), .Z(n5986) );
  XNOR U7412 ( .A(round_reg[1247]), .B(round_reg[1567]), .Z(n5984) );
  XOR U7413 ( .A(n5987), .B(n4899), .Z(o[1011]) );
  XNOR U7414 ( .A(n4770), .B(round_reg[182]), .Z(n4899) );
  XOR U7415 ( .A(n4805), .B(n4867), .Z(n4770) );
  XOR U7416 ( .A(n5988), .B(n5989), .Z(n4867) );
  XOR U7417 ( .A(round_reg[246]), .B(n5990), .Z(n5989) );
  XOR U7418 ( .A(round_reg[886]), .B(round_reg[566]), .Z(n5990) );
  XNOR U7419 ( .A(round_reg[1206]), .B(round_reg[1526]), .Z(n5988) );
  XNOR U7420 ( .A(n5991), .B(n5992), .Z(n4805) );
  XOR U7421 ( .A(round_reg[1397]), .B(n5993), .Z(n5992) );
  XOR U7422 ( .A(round_reg[757]), .B(round_reg[437]), .Z(n5993) );
  XNOR U7423 ( .A(round_reg[1077]), .B(round_reg[117]), .Z(n5991) );
  ANDN U7424 ( .A(n4474), .B(n4472), .Z(n5987) );
  XNOR U7425 ( .A(n1763), .B(round_reg[1367]), .Z(n4472) );
  XNOR U7426 ( .A(n5994), .B(n5995), .Z(n4991) );
  XOR U7427 ( .A(round_reg[342]), .B(n5996), .Z(n5995) );
  XOR U7428 ( .A(round_reg[982]), .B(round_reg[662]), .Z(n5996) );
  XNOR U7429 ( .A(round_reg[1302]), .B(round_reg[22]), .Z(n5994) );
  XOR U7430 ( .A(n5997), .B(n5998), .Z(n5678) );
  XOR U7431 ( .A(round_reg[151]), .B(n5999), .Z(n5998) );
  XOR U7432 ( .A(round_reg[791]), .B(round_reg[471]), .Z(n5999) );
  XNOR U7433 ( .A(round_reg[1111]), .B(round_reg[1431]), .Z(n5997) );
  XNOR U7434 ( .A(n4295), .B(round_reg[991]), .Z(n4474) );
  XOR U7435 ( .A(n5577), .B(n5322), .Z(n4295) );
  XOR U7436 ( .A(n6000), .B(n6001), .Z(n5322) );
  XOR U7437 ( .A(round_reg[415]), .B(n6002), .Z(n6001) );
  XOR U7438 ( .A(round_reg[95]), .B(round_reg[735]), .Z(n6002) );
  XNOR U7439 ( .A(round_reg[1055]), .B(round_reg[1375]), .Z(n6000) );
  XNOR U7440 ( .A(n6003), .B(n6004), .Z(n5577) );
  XOR U7441 ( .A(round_reg[286]), .B(n6005), .Z(n6004) );
  XOR U7442 ( .A(round_reg[926]), .B(round_reg[606]), .Z(n6005) );
  XNOR U7443 ( .A(round_reg[1246]), .B(round_reg[1566]), .Z(n6003) );
  XOR U7444 ( .A(n6006), .B(n4903), .Z(o[1010]) );
  XNOR U7445 ( .A(n4813), .B(round_reg[181]), .Z(n4903) );
  XOR U7446 ( .A(n4871), .B(n4809), .Z(n4813) );
  XOR U7447 ( .A(n6007), .B(n6008), .Z(n4809) );
  XOR U7448 ( .A(round_reg[1396]), .B(n6009), .Z(n6008) );
  XOR U7449 ( .A(round_reg[756]), .B(round_reg[436]), .Z(n6009) );
  XNOR U7450 ( .A(round_reg[1076]), .B(round_reg[116]), .Z(n6007) );
  XNOR U7451 ( .A(n6010), .B(n6011), .Z(n4871) );
  XOR U7452 ( .A(round_reg[245]), .B(n6012), .Z(n6011) );
  XOR U7453 ( .A(round_reg[885]), .B(round_reg[565]), .Z(n6012) );
  XNOR U7454 ( .A(round_reg[1205]), .B(round_reg[1525]), .Z(n6010) );
  ANDN U7455 ( .A(n4478), .B(n4476), .Z(n6006) );
  XNOR U7456 ( .A(n1766), .B(round_reg[1366]), .Z(n4476) );
  XNOR U7457 ( .A(n6013), .B(n6014), .Z(n4994) );
  XOR U7458 ( .A(round_reg[341]), .B(n6015), .Z(n6014) );
  XOR U7459 ( .A(round_reg[981]), .B(round_reg[661]), .Z(n6015) );
  XNOR U7460 ( .A(round_reg[1301]), .B(round_reg[21]), .Z(n6013) );
  XOR U7461 ( .A(n6016), .B(n6017), .Z(n5693) );
  XOR U7462 ( .A(round_reg[150]), .B(n6018), .Z(n6017) );
  XOR U7463 ( .A(round_reg[790]), .B(round_reg[470]), .Z(n6018) );
  XNOR U7464 ( .A(round_reg[1110]), .B(round_reg[1430]), .Z(n6016) );
  XNOR U7465 ( .A(n4307), .B(round_reg[990]), .Z(n4478) );
  XOR U7466 ( .A(n5592), .B(n5337), .Z(n4307) );
  XOR U7467 ( .A(n6019), .B(n6020), .Z(n5337) );
  XOR U7468 ( .A(round_reg[414]), .B(n6021), .Z(n6020) );
  XOR U7469 ( .A(round_reg[94]), .B(round_reg[734]), .Z(n6021) );
  XNOR U7470 ( .A(round_reg[1054]), .B(round_reg[1374]), .Z(n6019) );
  XNOR U7471 ( .A(n6022), .B(n6023), .Z(n5592) );
  XOR U7472 ( .A(round_reg[285]), .B(n6024), .Z(n6023) );
  XOR U7473 ( .A(round_reg[925]), .B(round_reg[605]), .Z(n6024) );
  XNOR U7474 ( .A(round_reg[1245]), .B(round_reg[1565]), .Z(n6022) );
  XOR U7475 ( .A(n6025), .B(n3516), .Z(o[100]) );
  XOR U7476 ( .A(n2335), .B(round_reg[635]), .Z(n3516) );
  IV U7477 ( .A(n4850), .Z(n2335) );
  XOR U7478 ( .A(n5916), .B(n5400), .Z(n4850) );
  XOR U7479 ( .A(n6026), .B(n6027), .Z(n5400) );
  XOR U7480 ( .A(round_reg[379]), .B(n6028), .Z(n6027) );
  XOR U7481 ( .A(round_reg[699]), .B(round_reg[59]), .Z(n6028) );
  XNOR U7482 ( .A(round_reg[1019]), .B(round_reg[1339]), .Z(n6026) );
  XNOR U7483 ( .A(n6029), .B(n6030), .Z(n5916) );
  XOR U7484 ( .A(round_reg[250]), .B(n6031), .Z(n6030) );
  XOR U7485 ( .A(round_reg[890]), .B(round_reg[570]), .Z(n6031) );
  XNOR U7486 ( .A(round_reg[1210]), .B(round_reg[1530]), .Z(n6029) );
  AND U7487 ( .A(n3199), .B(n3201), .Z(n6025) );
  XOR U7488 ( .A(n2200), .B(round_reg[1446]), .Z(n3201) );
  XOR U7489 ( .A(n4934), .B(n5892), .Z(n2200) );
  XOR U7490 ( .A(n6032), .B(n6033), .Z(n5892) );
  XOR U7491 ( .A(round_reg[1381]), .B(n6034), .Z(n6033) );
  XOR U7492 ( .A(round_reg[741]), .B(round_reg[421]), .Z(n6034) );
  XNOR U7493 ( .A(round_reg[101]), .B(round_reg[1061]), .Z(n6032) );
  XOR U7494 ( .A(n6035), .B(n6036), .Z(n4934) );
  XOR U7495 ( .A(round_reg[230]), .B(n6037), .Z(n6036) );
  XOR U7496 ( .A(round_reg[870]), .B(round_reg[550]), .Z(n6037) );
  XNOR U7497 ( .A(round_reg[1190]), .B(round_reg[1510]), .Z(n6035) );
  XNOR U7498 ( .A(n2241), .B(round_reg[226]), .Z(n3199) );
  XNOR U7499 ( .A(n5926), .B(n5799), .Z(n2241) );
  XOR U7500 ( .A(n6038), .B(n6039), .Z(n5799) );
  XOR U7501 ( .A(round_reg[161]), .B(n6040), .Z(n6039) );
  XOR U7502 ( .A(round_reg[801]), .B(round_reg[481]), .Z(n6040) );
  XNOR U7503 ( .A(round_reg[1121]), .B(round_reg[1441]), .Z(n6038) );
  XNOR U7504 ( .A(n6041), .B(n6042), .Z(n5926) );
  XOR U7505 ( .A(round_reg[290]), .B(n6043), .Z(n6042) );
  XOR U7506 ( .A(round_reg[930]), .B(round_reg[610]), .Z(n6043) );
  XNOR U7507 ( .A(round_reg[1250]), .B(round_reg[1570]), .Z(n6041) );
  XOR U7508 ( .A(n6044), .B(n4907), .Z(o[1009]) );
  XOR U7509 ( .A(n2140), .B(round_reg[180]), .Z(n4907) );
  XNOR U7510 ( .A(n4875), .B(n4816), .Z(n2140) );
  XOR U7511 ( .A(n6045), .B(n6046), .Z(n4816) );
  XOR U7512 ( .A(round_reg[1395]), .B(n6047), .Z(n6046) );
  XOR U7513 ( .A(round_reg[755]), .B(round_reg[435]), .Z(n6047) );
  XNOR U7514 ( .A(round_reg[1075]), .B(round_reg[115]), .Z(n6045) );
  XNOR U7515 ( .A(n6048), .B(n6049), .Z(n4875) );
  XOR U7516 ( .A(round_reg[244]), .B(n6050), .Z(n6049) );
  XOR U7517 ( .A(round_reg[884]), .B(round_reg[564]), .Z(n6050) );
  XNOR U7518 ( .A(round_reg[1204]), .B(round_reg[1524]), .Z(n6048) );
  ANDN U7519 ( .A(n4482), .B(n4480), .Z(n6044) );
  XNOR U7520 ( .A(n1769), .B(round_reg[1365]), .Z(n4480) );
  XNOR U7521 ( .A(n6051), .B(n6052), .Z(n4997) );
  XOR U7522 ( .A(round_reg[340]), .B(n6053), .Z(n6052) );
  XOR U7523 ( .A(round_reg[980]), .B(round_reg[660]), .Z(n6053) );
  XNOR U7524 ( .A(round_reg[1300]), .B(round_reg[20]), .Z(n6051) );
  XOR U7525 ( .A(n6054), .B(n6055), .Z(n5708) );
  XOR U7526 ( .A(round_reg[149]), .B(n6056), .Z(n6055) );
  XOR U7527 ( .A(round_reg[789]), .B(round_reg[469]), .Z(n6056) );
  XNOR U7528 ( .A(round_reg[1109]), .B(round_reg[1429]), .Z(n6054) );
  XNOR U7529 ( .A(n4329), .B(round_reg[989]), .Z(n4482) );
  XOR U7530 ( .A(n5607), .B(n5350), .Z(n4329) );
  XOR U7531 ( .A(n6057), .B(n6058), .Z(n5350) );
  XOR U7532 ( .A(round_reg[413]), .B(n6059), .Z(n6058) );
  XOR U7533 ( .A(round_reg[93]), .B(round_reg[733]), .Z(n6059) );
  XNOR U7534 ( .A(round_reg[1053]), .B(round_reg[1373]), .Z(n6057) );
  XNOR U7535 ( .A(n6060), .B(n6061), .Z(n5607) );
  XOR U7536 ( .A(round_reg[284]), .B(n6062), .Z(n6061) );
  XOR U7537 ( .A(round_reg[924]), .B(round_reg[604]), .Z(n6062) );
  XNOR U7538 ( .A(round_reg[1244]), .B(round_reg[1564]), .Z(n6060) );
  XOR U7539 ( .A(n6063), .B(n4911), .Z(o[1008]) );
  XOR U7540 ( .A(n2144), .B(round_reg[179]), .Z(n4911) );
  XNOR U7541 ( .A(n4879), .B(n4820), .Z(n2144) );
  XOR U7542 ( .A(n6064), .B(n6065), .Z(n4820) );
  XOR U7543 ( .A(round_reg[1394]), .B(n6066), .Z(n6065) );
  XOR U7544 ( .A(round_reg[754]), .B(round_reg[434]), .Z(n6066) );
  XNOR U7545 ( .A(round_reg[1074]), .B(round_reg[114]), .Z(n6064) );
  XNOR U7546 ( .A(n6067), .B(n6068), .Z(n4879) );
  XOR U7547 ( .A(round_reg[243]), .B(n6069), .Z(n6068) );
  XOR U7548 ( .A(round_reg[883]), .B(round_reg[563]), .Z(n6069) );
  XNOR U7549 ( .A(round_reg[1203]), .B(round_reg[1523]), .Z(n6067) );
  ANDN U7550 ( .A(n4486), .B(n4484), .Z(n6063) );
  XNOR U7551 ( .A(n1772), .B(round_reg[1364]), .Z(n4484) );
  XNOR U7552 ( .A(n6070), .B(n6071), .Z(n5000) );
  XOR U7553 ( .A(round_reg[339]), .B(n6072), .Z(n6071) );
  XOR U7554 ( .A(round_reg[979]), .B(round_reg[659]), .Z(n6072) );
  XNOR U7555 ( .A(round_reg[1299]), .B(round_reg[19]), .Z(n6070) );
  XOR U7556 ( .A(n6073), .B(n6074), .Z(n5723) );
  XOR U7557 ( .A(round_reg[148]), .B(n6075), .Z(n6074) );
  XOR U7558 ( .A(round_reg[788]), .B(round_reg[468]), .Z(n6075) );
  XNOR U7559 ( .A(round_reg[1108]), .B(round_reg[1428]), .Z(n6073) );
  XNOR U7560 ( .A(n4351), .B(round_reg[988]), .Z(n4486) );
  XOR U7561 ( .A(n5621), .B(n5363), .Z(n4351) );
  XOR U7562 ( .A(n6076), .B(n6077), .Z(n5363) );
  XOR U7563 ( .A(round_reg[412]), .B(n6078), .Z(n6077) );
  XOR U7564 ( .A(round_reg[92]), .B(round_reg[732]), .Z(n6078) );
  XNOR U7565 ( .A(round_reg[1052]), .B(round_reg[1372]), .Z(n6076) );
  XNOR U7566 ( .A(n6079), .B(n6080), .Z(n5621) );
  XOR U7567 ( .A(round_reg[283]), .B(n6081), .Z(n6080) );
  XOR U7568 ( .A(round_reg[923]), .B(round_reg[603]), .Z(n6081) );
  XNOR U7569 ( .A(round_reg[1243]), .B(round_reg[1563]), .Z(n6079) );
  XOR U7570 ( .A(n6082), .B(n4915), .Z(o[1007]) );
  XOR U7571 ( .A(n2148), .B(round_reg[178]), .Z(n4915) );
  XNOR U7572 ( .A(n4883), .B(n4824), .Z(n2148) );
  XOR U7573 ( .A(n6083), .B(n6084), .Z(n4824) );
  XOR U7574 ( .A(round_reg[1393]), .B(n6085), .Z(n6084) );
  XOR U7575 ( .A(round_reg[753]), .B(round_reg[433]), .Z(n6085) );
  XNOR U7576 ( .A(round_reg[1073]), .B(round_reg[113]), .Z(n6083) );
  XNOR U7577 ( .A(n6086), .B(n6087), .Z(n4883) );
  XOR U7578 ( .A(round_reg[242]), .B(n6088), .Z(n6087) );
  XOR U7579 ( .A(round_reg[882]), .B(round_reg[562]), .Z(n6088) );
  XNOR U7580 ( .A(round_reg[1202]), .B(round_reg[1522]), .Z(n6086) );
  ANDN U7581 ( .A(n4490), .B(n4488), .Z(n6082) );
  XNOR U7582 ( .A(n1775), .B(round_reg[1363]), .Z(n4488) );
  XNOR U7583 ( .A(n6089), .B(n6090), .Z(n5004) );
  XOR U7584 ( .A(round_reg[338]), .B(n6091), .Z(n6090) );
  XOR U7585 ( .A(round_reg[978]), .B(round_reg[658]), .Z(n6091) );
  XNOR U7586 ( .A(round_reg[1298]), .B(round_reg[18]), .Z(n6089) );
  XOR U7587 ( .A(n6092), .B(n6093), .Z(n5738) );
  XOR U7588 ( .A(round_reg[147]), .B(n6094), .Z(n6093) );
  XOR U7589 ( .A(round_reg[787]), .B(round_reg[467]), .Z(n6094) );
  XNOR U7590 ( .A(round_reg[1107]), .B(round_reg[1427]), .Z(n6092) );
  XNOR U7591 ( .A(n4376), .B(round_reg[987]), .Z(n4490) );
  XOR U7592 ( .A(n5636), .B(n5385), .Z(n4376) );
  XOR U7593 ( .A(n6095), .B(n6096), .Z(n5385) );
  XOR U7594 ( .A(round_reg[411]), .B(n6097), .Z(n6096) );
  XOR U7595 ( .A(round_reg[91]), .B(round_reg[731]), .Z(n6097) );
  XNOR U7596 ( .A(round_reg[1051]), .B(round_reg[1371]), .Z(n6095) );
  XNOR U7597 ( .A(n6098), .B(n6099), .Z(n5636) );
  XOR U7598 ( .A(round_reg[282]), .B(n6100), .Z(n6099) );
  XOR U7599 ( .A(round_reg[922]), .B(round_reg[602]), .Z(n6100) );
  XNOR U7600 ( .A(round_reg[1242]), .B(round_reg[1562]), .Z(n6098) );
  XOR U7601 ( .A(n6101), .B(n4919), .Z(o[1006]) );
  XOR U7602 ( .A(n2152), .B(round_reg[177]), .Z(n4919) );
  XNOR U7603 ( .A(n4887), .B(n4828), .Z(n2152) );
  XOR U7604 ( .A(n6102), .B(n6103), .Z(n4828) );
  XOR U7605 ( .A(round_reg[1392]), .B(n6104), .Z(n6103) );
  XOR U7606 ( .A(round_reg[752]), .B(round_reg[432]), .Z(n6104) );
  XNOR U7607 ( .A(round_reg[1072]), .B(round_reg[112]), .Z(n6102) );
  XNOR U7608 ( .A(n6105), .B(n6106), .Z(n4887) );
  XOR U7609 ( .A(round_reg[241]), .B(n6107), .Z(n6106) );
  XOR U7610 ( .A(round_reg[881]), .B(round_reg[561]), .Z(n6107) );
  XNOR U7611 ( .A(round_reg[1201]), .B(round_reg[1521]), .Z(n6105) );
  ANDN U7612 ( .A(n4494), .B(n4492), .Z(n6101) );
  XOR U7613 ( .A(n1778), .B(round_reg[1362]), .Z(n4492) );
  XOR U7614 ( .A(n5753), .B(n5008), .Z(n1778) );
  XOR U7615 ( .A(n6108), .B(n6109), .Z(n5008) );
  XOR U7616 ( .A(round_reg[337]), .B(n6110), .Z(n6109) );
  XOR U7617 ( .A(round_reg[977]), .B(round_reg[657]), .Z(n6110) );
  XNOR U7618 ( .A(round_reg[1297]), .B(round_reg[17]), .Z(n6108) );
  XOR U7619 ( .A(n6111), .B(n6112), .Z(n5753) );
  XOR U7620 ( .A(round_reg[146]), .B(n6113), .Z(n6112) );
  XOR U7621 ( .A(round_reg[786]), .B(round_reg[466]), .Z(n6113) );
  XNOR U7622 ( .A(round_reg[1106]), .B(round_reg[1426]), .Z(n6111) );
  XNOR U7623 ( .A(n4390), .B(round_reg[986]), .Z(n4494) );
  XOR U7624 ( .A(n5651), .B(n5396), .Z(n4390) );
  XOR U7625 ( .A(n6114), .B(n6115), .Z(n5396) );
  XOR U7626 ( .A(round_reg[410]), .B(n6116), .Z(n6115) );
  XOR U7627 ( .A(round_reg[90]), .B(round_reg[730]), .Z(n6116) );
  XNOR U7628 ( .A(round_reg[1050]), .B(round_reg[1370]), .Z(n6114) );
  XNOR U7629 ( .A(n6117), .B(n6118), .Z(n5651) );
  XOR U7630 ( .A(round_reg[281]), .B(n6119), .Z(n6118) );
  XOR U7631 ( .A(round_reg[921]), .B(round_reg[601]), .Z(n6119) );
  XNOR U7632 ( .A(round_reg[1241]), .B(round_reg[1561]), .Z(n6117) );
  XOR U7633 ( .A(n6120), .B(n4923), .Z(o[1005]) );
  XOR U7634 ( .A(n2156), .B(round_reg[176]), .Z(n4923) );
  XNOR U7635 ( .A(n4891), .B(n4832), .Z(n2156) );
  XOR U7636 ( .A(n6121), .B(n6122), .Z(n4832) );
  XOR U7637 ( .A(round_reg[1391]), .B(n6123), .Z(n6122) );
  XOR U7638 ( .A(round_reg[751]), .B(round_reg[431]), .Z(n6123) );
  XNOR U7639 ( .A(round_reg[1071]), .B(round_reg[111]), .Z(n6121) );
  XNOR U7640 ( .A(n6124), .B(n6125), .Z(n4891) );
  XOR U7641 ( .A(round_reg[240]), .B(n6126), .Z(n6125) );
  XOR U7642 ( .A(round_reg[880]), .B(round_reg[560]), .Z(n6126) );
  XNOR U7643 ( .A(round_reg[1200]), .B(round_reg[1520]), .Z(n6124) );
  ANDN U7644 ( .A(n4498), .B(n4496), .Z(n6120) );
  XNOR U7645 ( .A(n4248), .B(round_reg[1361]), .Z(n4496) );
  XNOR U7646 ( .A(n6127), .B(n6128), .Z(n5010) );
  XOR U7647 ( .A(round_reg[336]), .B(n6129), .Z(n6128) );
  XOR U7648 ( .A(round_reg[976]), .B(round_reg[656]), .Z(n6129) );
  XNOR U7649 ( .A(round_reg[1296]), .B(round_reg[16]), .Z(n6127) );
  XNOR U7650 ( .A(n6130), .B(n6131), .Z(n5069) );
  XOR U7651 ( .A(round_reg[145]), .B(n6132), .Z(n6131) );
  XOR U7652 ( .A(round_reg[785]), .B(round_reg[465]), .Z(n6132) );
  XNOR U7653 ( .A(round_reg[1105]), .B(round_reg[1425]), .Z(n6130) );
  XNOR U7654 ( .A(n4403), .B(round_reg[985]), .Z(n4498) );
  XOR U7655 ( .A(n5677), .B(n5407), .Z(n4403) );
  XOR U7656 ( .A(n6133), .B(n6134), .Z(n5407) );
  XOR U7657 ( .A(round_reg[409]), .B(n6135), .Z(n6134) );
  XOR U7658 ( .A(round_reg[89]), .B(round_reg[729]), .Z(n6135) );
  XNOR U7659 ( .A(round_reg[1049]), .B(round_reg[1369]), .Z(n6133) );
  XNOR U7660 ( .A(n6136), .B(n6137), .Z(n5677) );
  XOR U7661 ( .A(round_reg[280]), .B(n6138), .Z(n6137) );
  XOR U7662 ( .A(round_reg[920]), .B(round_reg[600]), .Z(n6138) );
  XNOR U7663 ( .A(round_reg[1240]), .B(round_reg[1560]), .Z(n6136) );
  XOR U7664 ( .A(n6139), .B(n4927), .Z(o[1004]) );
  XOR U7665 ( .A(n2160), .B(round_reg[175]), .Z(n4927) );
  XNOR U7666 ( .A(n4897), .B(n4836), .Z(n2160) );
  XOR U7667 ( .A(n6140), .B(n6141), .Z(n4836) );
  XOR U7668 ( .A(round_reg[1390]), .B(n6142), .Z(n6141) );
  XOR U7669 ( .A(round_reg[750]), .B(round_reg[430]), .Z(n6142) );
  XNOR U7670 ( .A(round_reg[1070]), .B(round_reg[110]), .Z(n6140) );
  XNOR U7671 ( .A(n6143), .B(n6144), .Z(n4897) );
  XOR U7672 ( .A(round_reg[239]), .B(n6145), .Z(n6144) );
  XOR U7673 ( .A(round_reg[879]), .B(round_reg[559]), .Z(n6145) );
  XNOR U7674 ( .A(round_reg[1199]), .B(round_reg[1519]), .Z(n6143) );
  ANDN U7675 ( .A(n4502), .B(n4500), .Z(n6139) );
  XNOR U7676 ( .A(n4250), .B(round_reg[1360]), .Z(n4500) );
  XOR U7677 ( .A(n5074), .B(n6146), .Z(n4250) );
  IV U7678 ( .A(n5013), .Z(n6146) );
  XNOR U7679 ( .A(n6147), .B(n6148), .Z(n5013) );
  XOR U7680 ( .A(round_reg[335]), .B(n6149), .Z(n6148) );
  XOR U7681 ( .A(round_reg[975]), .B(round_reg[655]), .Z(n6149) );
  XNOR U7682 ( .A(round_reg[1295]), .B(round_reg[15]), .Z(n6147) );
  XNOR U7683 ( .A(n6150), .B(n6151), .Z(n5074) );
  XOR U7684 ( .A(round_reg[144]), .B(n6152), .Z(n6151) );
  XOR U7685 ( .A(round_reg[784]), .B(round_reg[464]), .Z(n6152) );
  XNOR U7686 ( .A(round_reg[1104]), .B(round_reg[1424]), .Z(n6150) );
  XNOR U7687 ( .A(n4355), .B(round_reg[984]), .Z(n4502) );
  XOR U7688 ( .A(n5692), .B(n5420), .Z(n4355) );
  XOR U7689 ( .A(n6153), .B(n6154), .Z(n5420) );
  XOR U7690 ( .A(round_reg[408]), .B(n6155), .Z(n6154) );
  XOR U7691 ( .A(round_reg[88]), .B(round_reg[728]), .Z(n6155) );
  XNOR U7692 ( .A(round_reg[1048]), .B(round_reg[1368]), .Z(n6153) );
  XNOR U7693 ( .A(n6156), .B(n6157), .Z(n5692) );
  XOR U7694 ( .A(round_reg[279]), .B(n6158), .Z(n6157) );
  XOR U7695 ( .A(round_reg[919]), .B(round_reg[599]), .Z(n6158) );
  XNOR U7696 ( .A(round_reg[1239]), .B(round_reg[1559]), .Z(n6156) );
  XOR U7697 ( .A(n6159), .B(n4931), .Z(o[1003]) );
  XOR U7698 ( .A(n2164), .B(round_reg[174]), .Z(n4931) );
  XNOR U7699 ( .A(n4901), .B(n4840), .Z(n2164) );
  XOR U7700 ( .A(n6160), .B(n6161), .Z(n4840) );
  XOR U7701 ( .A(round_reg[1389]), .B(n6162), .Z(n6161) );
  XOR U7702 ( .A(round_reg[749]), .B(round_reg[429]), .Z(n6162) );
  XNOR U7703 ( .A(round_reg[1069]), .B(round_reg[109]), .Z(n6160) );
  XNOR U7704 ( .A(n6163), .B(n6164), .Z(n4901) );
  XOR U7705 ( .A(round_reg[238]), .B(n6165), .Z(n6164) );
  XOR U7706 ( .A(round_reg[878]), .B(round_reg[558]), .Z(n6165) );
  XNOR U7707 ( .A(round_reg[1198]), .B(round_reg[1518]), .Z(n6163) );
  ANDN U7708 ( .A(n4508), .B(n4506), .Z(n6159) );
  XNOR U7709 ( .A(n4252), .B(round_reg[1359]), .Z(n4506) );
  XOR U7710 ( .A(n5079), .B(n6166), .Z(n4252) );
  IV U7711 ( .A(n5016), .Z(n6166) );
  XNOR U7712 ( .A(n6167), .B(n6168), .Z(n5016) );
  XOR U7713 ( .A(round_reg[334]), .B(n6169), .Z(n6168) );
  XOR U7714 ( .A(round_reg[974]), .B(round_reg[654]), .Z(n6169) );
  XNOR U7715 ( .A(round_reg[1294]), .B(round_reg[14]), .Z(n6167) );
  XNOR U7716 ( .A(n6170), .B(n6171), .Z(n5079) );
  XOR U7717 ( .A(round_reg[143]), .B(n6172), .Z(n6171) );
  XOR U7718 ( .A(round_reg[783]), .B(round_reg[463]), .Z(n6172) );
  XNOR U7719 ( .A(round_reg[1103]), .B(round_reg[1423]), .Z(n6170) );
  XNOR U7720 ( .A(n4358), .B(round_reg[983]), .Z(n4508) );
  XOR U7721 ( .A(n5707), .B(n5433), .Z(n4358) );
  XOR U7722 ( .A(n6173), .B(n6174), .Z(n5433) );
  XOR U7723 ( .A(round_reg[407]), .B(n6175), .Z(n6174) );
  XOR U7724 ( .A(round_reg[87]), .B(round_reg[727]), .Z(n6175) );
  XNOR U7725 ( .A(round_reg[1047]), .B(round_reg[1367]), .Z(n6173) );
  XNOR U7726 ( .A(n6176), .B(n6177), .Z(n5707) );
  XOR U7727 ( .A(round_reg[278]), .B(n6178), .Z(n6177) );
  XOR U7728 ( .A(round_reg[918]), .B(round_reg[598]), .Z(n6178) );
  XNOR U7729 ( .A(round_reg[1238]), .B(round_reg[1558]), .Z(n6176) );
  XOR U7730 ( .A(n6179), .B(n4935), .Z(o[1002]) );
  XOR U7731 ( .A(n2168), .B(round_reg[173]), .Z(n4935) );
  XNOR U7732 ( .A(n4905), .B(n4844), .Z(n2168) );
  XOR U7733 ( .A(n6180), .B(n6181), .Z(n4844) );
  XOR U7734 ( .A(round_reg[1388]), .B(n6182), .Z(n6181) );
  XOR U7735 ( .A(round_reg[748]), .B(round_reg[428]), .Z(n6182) );
  XNOR U7736 ( .A(round_reg[1068]), .B(round_reg[108]), .Z(n6180) );
  XNOR U7737 ( .A(n6183), .B(n6184), .Z(n4905) );
  XOR U7738 ( .A(round_reg[237]), .B(n6185), .Z(n6184) );
  XOR U7739 ( .A(round_reg[877]), .B(round_reg[557]), .Z(n6185) );
  XNOR U7740 ( .A(round_reg[1197]), .B(round_reg[1517]), .Z(n6183) );
  ANDN U7741 ( .A(n4512), .B(n4510), .Z(n6179) );
  XNOR U7742 ( .A(n4256), .B(round_reg[1358]), .Z(n4510) );
  XOR U7743 ( .A(n5084), .B(n6186), .Z(n4256) );
  IV U7744 ( .A(n5019), .Z(n6186) );
  XNOR U7745 ( .A(n6187), .B(n6188), .Z(n5019) );
  XOR U7746 ( .A(round_reg[333]), .B(n6189), .Z(n6188) );
  XOR U7747 ( .A(round_reg[973]), .B(round_reg[653]), .Z(n6189) );
  XNOR U7748 ( .A(round_reg[1293]), .B(round_reg[13]), .Z(n6187) );
  XNOR U7749 ( .A(n6190), .B(n6191), .Z(n5084) );
  XOR U7750 ( .A(round_reg[142]), .B(n6192), .Z(n6191) );
  XOR U7751 ( .A(round_reg[782]), .B(round_reg[462]), .Z(n6192) );
  XNOR U7752 ( .A(round_reg[1102]), .B(round_reg[1422]), .Z(n6190) );
  XNOR U7753 ( .A(n4361), .B(round_reg[982]), .Z(n4512) );
  XOR U7754 ( .A(n5722), .B(n5446), .Z(n4361) );
  XOR U7755 ( .A(n6193), .B(n6194), .Z(n5446) );
  XOR U7756 ( .A(round_reg[406]), .B(n6195), .Z(n6194) );
  XOR U7757 ( .A(round_reg[86]), .B(round_reg[726]), .Z(n6195) );
  XNOR U7758 ( .A(round_reg[1046]), .B(round_reg[1366]), .Z(n6193) );
  XNOR U7759 ( .A(n6196), .B(n6197), .Z(n5722) );
  XOR U7760 ( .A(round_reg[277]), .B(n6198), .Z(n6197) );
  XOR U7761 ( .A(round_reg[917]), .B(round_reg[597]), .Z(n6198) );
  XNOR U7762 ( .A(round_reg[1237]), .B(round_reg[1557]), .Z(n6196) );
  XOR U7763 ( .A(n6199), .B(n4941), .Z(o[1001]) );
  XNOR U7764 ( .A(n2172), .B(round_reg[172]), .Z(n4941) );
  XNOR U7765 ( .A(n6200), .B(n6201), .Z(n4909) );
  XOR U7766 ( .A(round_reg[236]), .B(n6202), .Z(n6201) );
  XOR U7767 ( .A(round_reg[876]), .B(round_reg[556]), .Z(n6202) );
  XNOR U7768 ( .A(round_reg[1196]), .B(round_reg[1516]), .Z(n6200) );
  XOR U7769 ( .A(n6203), .B(n6204), .Z(n5773) );
  XOR U7770 ( .A(round_reg[1387]), .B(n6205), .Z(n6204) );
  XOR U7771 ( .A(round_reg[747]), .B(round_reg[427]), .Z(n6205) );
  XNOR U7772 ( .A(round_reg[1067]), .B(round_reg[107]), .Z(n6203) );
  ANDN U7773 ( .A(n4516), .B(n4514), .Z(n6199) );
  XNOR U7774 ( .A(n4259), .B(round_reg[1357]), .Z(n4514) );
  XOR U7775 ( .A(n5089), .B(n6206), .Z(n4259) );
  IV U7776 ( .A(n5022), .Z(n6206) );
  XNOR U7777 ( .A(n6207), .B(n6208), .Z(n5022) );
  XOR U7778 ( .A(round_reg[332]), .B(n6209), .Z(n6208) );
  XOR U7779 ( .A(round_reg[972]), .B(round_reg[652]), .Z(n6209) );
  XNOR U7780 ( .A(round_reg[1292]), .B(round_reg[12]), .Z(n6207) );
  XNOR U7781 ( .A(n6210), .B(n6211), .Z(n5089) );
  XOR U7782 ( .A(round_reg[1421]), .B(n6212), .Z(n6211) );
  XOR U7783 ( .A(round_reg[781]), .B(round_reg[461]), .Z(n6212) );
  XNOR U7784 ( .A(round_reg[1101]), .B(round_reg[141]), .Z(n6210) );
  XNOR U7785 ( .A(n4364), .B(round_reg[981]), .Z(n4516) );
  XOR U7786 ( .A(n5737), .B(n5459), .Z(n4364) );
  XOR U7787 ( .A(n6213), .B(n6214), .Z(n5459) );
  XOR U7788 ( .A(round_reg[405]), .B(n6215), .Z(n6214) );
  XOR U7789 ( .A(round_reg[85]), .B(round_reg[725]), .Z(n6215) );
  XNOR U7790 ( .A(round_reg[1045]), .B(round_reg[1365]), .Z(n6213) );
  XNOR U7791 ( .A(n6216), .B(n6217), .Z(n5737) );
  XOR U7792 ( .A(round_reg[276]), .B(n6218), .Z(n6217) );
  XOR U7793 ( .A(round_reg[916]), .B(round_reg[596]), .Z(n6218) );
  XNOR U7794 ( .A(round_reg[1236]), .B(round_reg[1556]), .Z(n6216) );
  XOR U7795 ( .A(n6219), .B(n4945), .Z(o[1000]) );
  XNOR U7796 ( .A(n2180), .B(round_reg[171]), .Z(n4945) );
  XNOR U7797 ( .A(n6220), .B(n6221), .Z(n4913) );
  XOR U7798 ( .A(round_reg[235]), .B(n6222), .Z(n6221) );
  XOR U7799 ( .A(round_reg[875]), .B(round_reg[555]), .Z(n6222) );
  XNOR U7800 ( .A(round_reg[1195]), .B(round_reg[1515]), .Z(n6220) );
  XOR U7801 ( .A(n6223), .B(n6224), .Z(n5788) );
  XOR U7802 ( .A(round_reg[1386]), .B(n6225), .Z(n6224) );
  XOR U7803 ( .A(round_reg[746]), .B(round_reg[426]), .Z(n6225) );
  XNOR U7804 ( .A(round_reg[1066]), .B(round_reg[106]), .Z(n6223) );
  ANDN U7805 ( .A(n4520), .B(n4518), .Z(n6219) );
  XNOR U7806 ( .A(n4262), .B(round_reg[1356]), .Z(n4518) );
  XOR U7807 ( .A(n5094), .B(n6226), .Z(n4262) );
  IV U7808 ( .A(n5025), .Z(n6226) );
  XNOR U7809 ( .A(n6227), .B(n6228), .Z(n5025) );
  XOR U7810 ( .A(round_reg[331]), .B(n6229), .Z(n6228) );
  XOR U7811 ( .A(round_reg[971]), .B(round_reg[651]), .Z(n6229) );
  XNOR U7812 ( .A(round_reg[11]), .B(round_reg[1291]), .Z(n6227) );
  XNOR U7813 ( .A(n6230), .B(n6231), .Z(n5094) );
  XOR U7814 ( .A(round_reg[1420]), .B(n6232), .Z(n6231) );
  XOR U7815 ( .A(round_reg[780]), .B(round_reg[460]), .Z(n6232) );
  XNOR U7816 ( .A(round_reg[1100]), .B(round_reg[140]), .Z(n6230) );
  XNOR U7817 ( .A(n4367), .B(round_reg[980]), .Z(n4520) );
  XOR U7818 ( .A(n5752), .B(n5470), .Z(n4367) );
  XOR U7819 ( .A(n6233), .B(n6234), .Z(n5470) );
  XOR U7820 ( .A(round_reg[404]), .B(n6235), .Z(n6234) );
  XOR U7821 ( .A(round_reg[84]), .B(round_reg[724]), .Z(n6235) );
  XNOR U7822 ( .A(round_reg[1044]), .B(round_reg[1364]), .Z(n6233) );
  XNOR U7823 ( .A(n6236), .B(n6237), .Z(n5752) );
  XOR U7824 ( .A(round_reg[275]), .B(n6238), .Z(n6237) );
  XOR U7825 ( .A(round_reg[915]), .B(round_reg[595]), .Z(n6238) );
  XNOR U7826 ( .A(round_reg[1235]), .B(round_reg[1555]), .Z(n6236) );
  XOR U7827 ( .A(n6239), .B(n2353), .Z(o[0]) );
  XOR U7828 ( .A(n3029), .B(round_reg[254]), .Z(n2353) );
  IV U7829 ( .A(n2113), .Z(n3029) );
  XOR U7830 ( .A(n4762), .B(n5389), .Z(n2113) );
  XOR U7831 ( .A(n6240), .B(n6241), .Z(n5389) );
  XOR U7832 ( .A(round_reg[189]), .B(n6242), .Z(n6241) );
  XOR U7833 ( .A(round_reg[829]), .B(round_reg[509]), .Z(n6242) );
  XNOR U7834 ( .A(round_reg[1149]), .B(round_reg[1469]), .Z(n6240) );
  XNOR U7835 ( .A(n6243), .B(n6244), .Z(n4762) );
  XOR U7836 ( .A(round_reg[318]), .B(n6245), .Z(n6244) );
  XOR U7837 ( .A(round_reg[958]), .B(round_reg[638]), .Z(n6245) );
  XNOR U7838 ( .A(round_reg[1278]), .B(round_reg[1598]), .Z(n6243) );
  AND U7839 ( .A(n3457), .B(n3455), .Z(n6239) );
  XNOR U7840 ( .A(n2360), .B(round_reg[1410]), .Z(n3455) );
  XNOR U7841 ( .A(n5062), .B(n4754), .Z(n2360) );
  XOR U7842 ( .A(n6246), .B(n6247), .Z(n4754) );
  XOR U7843 ( .A(round_reg[385]), .B(n6248), .Z(n6247) );
  XOR U7844 ( .A(round_reg[705]), .B(round_reg[65]), .Z(n6248) );
  XNOR U7845 ( .A(round_reg[1025]), .B(round_reg[1345]), .Z(n6246) );
  XNOR U7846 ( .A(n6249), .B(n6250), .Z(n5062) );
  XOR U7847 ( .A(round_reg[194]), .B(n6251), .Z(n6250) );
  XOR U7848 ( .A(round_reg[834]), .B(round_reg[514]), .Z(n6251) );
  XNOR U7849 ( .A(round_reg[1154]), .B(round_reg[1474]), .Z(n6249) );
  XOR U7850 ( .A(n1809), .B(round_reg[1033]), .Z(n3457) );
  XOR U7851 ( .A(n5112), .B(n5038), .Z(n1809) );
  XOR U7852 ( .A(n6252), .B(n6253), .Z(n5038) );
  XOR U7853 ( .A(round_reg[648]), .B(n6254), .Z(n6253) );
  XOR U7854 ( .A(round_reg[968]), .B(round_reg[8]), .Z(n6254) );
  XNOR U7855 ( .A(round_reg[1288]), .B(round_reg[328]), .Z(n6252) );
  XOR U7856 ( .A(n6255), .B(n6256), .Z(n5112) );
  XOR U7857 ( .A(round_reg[1417]), .B(n6257), .Z(n6256) );
  XOR U7858 ( .A(round_reg[777]), .B(round_reg[457]), .Z(n6257) );
  XNOR U7859 ( .A(round_reg[1097]), .B(round_reg[137]), .Z(n6255) );
  IV U7860 ( .A(init), .Z(n1050) );
endmodule

