
module mult_N64_CC1 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341;

  XNOR U2 ( .A(n304), .B(n305), .Z(n306) );
  XOR U3 ( .A(n970), .B(n971), .Z(n973) );
  XOR U4 ( .A(n7701), .B(n7702), .Z(n8083) );
  XNOR U5 ( .A(n18982), .B(n18983), .Z(n19361) );
  XNOR U6 ( .A(n7891), .B(n7892), .Z(n8274) );
  XNOR U7 ( .A(n624), .B(n625), .Z(n626) );
  XNOR U8 ( .A(n306), .B(n307), .Z(n384) );
  XNOR U9 ( .A(n436), .B(n437), .Z(n438) );
  XNOR U10 ( .A(n1360), .B(n1361), .Z(n1562) );
  XNOR U11 ( .A(n1202), .B(n1203), .Z(n1282) );
  XNOR U12 ( .A(n2722), .B(n2723), .Z(n3036) );
  XOR U13 ( .A(n2434), .B(n2435), .Z(n2637) );
  XNOR U14 ( .A(n826), .B(n827), .Z(n967) );
  XNOR U15 ( .A(n3052), .B(n3053), .Z(n3182) );
  XNOR U16 ( .A(n4680), .B(n4681), .Z(n5103) );
  XNOR U17 ( .A(n5418), .B(n5419), .Z(n5850) );
  XOR U18 ( .A(n4284), .B(n4285), .Z(n4286) );
  XNOR U19 ( .A(n3082), .B(n3083), .Z(n3172) );
  XNOR U20 ( .A(n7248), .B(n7249), .Z(n7701) );
  XNOR U21 ( .A(n7699), .B(n7700), .Z(n8082) );
  XNOR U22 ( .A(n5444), .B(n5445), .Z(n5836) );
  XOR U23 ( .A(n7713), .B(n7714), .Z(n8095) );
  XOR U24 ( .A(n9228), .B(n9229), .Z(n9610) );
  XNOR U25 ( .A(n3112), .B(n3113), .Z(n3114) );
  XOR U26 ( .A(n7725), .B(n7726), .Z(n8107) );
  XNOR U27 ( .A(n6488), .B(n6489), .Z(n7074) );
  XOR U28 ( .A(n7737), .B(n7738), .Z(n8119) );
  XOR U29 ( .A(n10766), .B(n10767), .Z(n11148) );
  XOR U30 ( .A(n7749), .B(n7750), .Z(n8131) );
  XOR U31 ( .A(n7761), .B(n7762), .Z(n8143) );
  XOR U32 ( .A(n12300), .B(n12301), .Z(n12684) );
  XOR U33 ( .A(n7773), .B(n7774), .Z(n8155) );
  XOR U34 ( .A(n15928), .B(n15929), .Z(n15930) );
  XOR U35 ( .A(n7785), .B(n7786), .Z(n8167) );
  XNOR U36 ( .A(n3942), .B(n3943), .Z(n4216) );
  XNOR U37 ( .A(n3496), .B(n3497), .Z(n3946) );
  XOR U38 ( .A(n13844), .B(n13845), .Z(n14226) );
  XOR U39 ( .A(n7797), .B(n7798), .Z(n8179) );
  XNOR U40 ( .A(n5202), .B(n5203), .Z(n5508) );
  XOR U41 ( .A(n7809), .B(n7810), .Z(n8191) );
  XOR U42 ( .A(n15380), .B(n15381), .Z(n15762) );
  XNOR U43 ( .A(n4923), .B(n4922), .Z(n4812) );
  XNOR U44 ( .A(n4802), .B(n4803), .Z(n4804) );
  XOR U45 ( .A(n7833), .B(n7834), .Z(n8215) );
  XNOR U46 ( .A(n5532), .B(n5533), .Z(n6110) );
  XOR U47 ( .A(n7845), .B(n7846), .Z(n8227) );
  XNOR U48 ( .A(n18577), .B(n18578), .Z(n18966) );
  XOR U49 ( .A(n18984), .B(n18985), .Z(n19362) );
  XOR U50 ( .A(n7857), .B(n7858), .Z(n8239) );
  XNOR U51 ( .A(n19359), .B(n19360), .Z(n19752) );
  XOR U52 ( .A(n18833), .B(n18834), .Z(n19221) );
  XOR U53 ( .A(n7869), .B(n7870), .Z(n8251) );
  XNOR U54 ( .A(n19740), .B(n19741), .Z(n20127) );
  XOR U55 ( .A(n19748), .B(n19749), .Z(n20132) );
  XOR U56 ( .A(n7881), .B(n7882), .Z(n8263) );
  XOR U57 ( .A(n20377), .B(n20378), .Z(n20751) );
  XOR U58 ( .A(n7893), .B(n7894), .Z(n8275) );
  ANDN U59 ( .B(n15102), .A(n15101), .Z(n24155) );
  XNOR U60 ( .A(n626), .B(n627), .Z(n768) );
  XNOR U61 ( .A(n312), .B(n313), .Z(n382) );
  XNOR U62 ( .A(n532), .B(n533), .Z(n534) );
  XNOR U63 ( .A(n438), .B(n439), .Z(n538) );
  XNOR U64 ( .A(n1630), .B(n1631), .Z(n1804) );
  XNOR U65 ( .A(n5944), .B(n5945), .Z(n5947) );
  XNOR U66 ( .A(n2200), .B(n2201), .Z(n2434) );
  XOR U67 ( .A(n1562), .B(n1563), .Z(n1645) );
  XNOR U68 ( .A(n1206), .B(n1207), .Z(n1278) );
  XNOR U69 ( .A(n556), .B(n557), .Z(n674) );
  XNOR U70 ( .A(n342), .B(n343), .Z(n344) );
  XNOR U71 ( .A(n5372), .B(n5373), .Z(n5958) );
  XNOR U72 ( .A(n4382), .B(n4383), .Z(n4648) );
  XNOR U73 ( .A(n3814), .B(n3815), .Z(n4080) );
  XNOR U74 ( .A(n3032), .B(n3033), .Z(n3273) );
  XNOR U75 ( .A(n2432), .B(n2433), .Z(n2636) );
  NAND U76 ( .A(n2211), .B(n2209), .Z(n2) );
  XOR U77 ( .A(n2209), .B(n2211), .Z(n3) );
  NAND U78 ( .A(n3), .B(n2208), .Z(n4) );
  NAND U79 ( .A(n2), .B(n4), .Z(n1884) );
  XNOR U80 ( .A(n1058), .B(n1059), .Z(n1120) );
  XNOR U81 ( .A(n3036), .B(n3037), .Z(n3038) );
  XNOR U82 ( .A(n832), .B(n833), .Z(n964) );
  XNOR U83 ( .A(n684), .B(n685), .Z(n687) );
  XNOR U84 ( .A(n3048), .B(n3049), .Z(n3184) );
  XNOR U85 ( .A(n2736), .B(n2737), .Z(n2944) );
  XNOR U86 ( .A(n2232), .B(n2233), .Z(n2338) );
  XNOR U87 ( .A(n1388), .B(n1389), .Z(n1551) );
  XNOR U88 ( .A(n1228), .B(n1229), .Z(n1393) );
  XNOR U89 ( .A(n4664), .B(n4665), .Z(n4968) );
  XOR U90 ( .A(n3724), .B(n3725), .Z(n3727) );
  XNOR U91 ( .A(n1398), .B(n1399), .Z(n1544) );
  XNOR U92 ( .A(n1238), .B(n1239), .Z(n1272) );
  XNOR U93 ( .A(n10953), .B(n10954), .Z(n11332) );
  XNOR U94 ( .A(n11328), .B(n11329), .Z(n11703) );
  XOR U95 ( .A(n5420), .B(n5421), .Z(n5851) );
  XOR U96 ( .A(n3316), .B(n3317), .Z(n3717) );
  XNOR U97 ( .A(n1924), .B(n1925), .Z(n2261) );
  XNOR U98 ( .A(n7244), .B(n7245), .Z(n7695) );
  XOR U99 ( .A(n4962), .B(n4963), .Z(n4964) );
  XOR U100 ( .A(n12515), .B(n12516), .Z(n12517) );
  XOR U101 ( .A(n3714), .B(n3715), .Z(n3874) );
  XNOR U102 ( .A(n2782), .B(n2783), .Z(n2926) );
  XOR U103 ( .A(n8082), .B(n8083), .Z(n8465) );
  XNOR U104 ( .A(n5128), .B(n5129), .Z(n5269) );
  XNOR U105 ( .A(n7256), .B(n7257), .Z(n7713) );
  XNOR U106 ( .A(n1710), .B(n1711), .Z(n1712) );
  XNOR U107 ( .A(n7711), .B(n7712), .Z(n8094) );
  XNOR U108 ( .A(n5448), .B(n5449), .Z(n6024) );
  XNOR U109 ( .A(n7264), .B(n7265), .Z(n7725) );
  XOR U110 ( .A(n4270), .B(n4271), .Z(n4729) );
  XNOR U111 ( .A(n3894), .B(n3895), .Z(n3964) );
  XNOR U112 ( .A(n3114), .B(n3115), .Z(n3164) );
  XOR U113 ( .A(n2610), .B(n2611), .Z(n2800) );
  XNOR U114 ( .A(n2500), .B(n2501), .Z(n2804) );
  XNOR U115 ( .A(n3644), .B(n3645), .Z(n3624) );
  XOR U116 ( .A(n9609), .B(n9610), .Z(n9997) );
  XNOR U117 ( .A(n7723), .B(n7724), .Z(n8106) );
  XNOR U118 ( .A(n4156), .B(n4157), .Z(n4264) );
  XOR U119 ( .A(n13972), .B(n13973), .Z(n14038) );
  XNOR U120 ( .A(n7272), .B(n7273), .Z(n7737) );
  XNOR U121 ( .A(n2034), .B(n2035), .Z(n2300) );
  XNOR U122 ( .A(n5616), .B(n5617), .Z(n5596) );
  XNOR U123 ( .A(n7735), .B(n7736), .Z(n8118) );
  XNOR U124 ( .A(n4738), .B(n4739), .Z(n4952) );
  XOR U125 ( .A(n14347), .B(n14348), .Z(n14389) );
  XNOR U126 ( .A(n7280), .B(n7281), .Z(n7749) );
  XNOR U127 ( .A(n5468), .B(n5469), .Z(n6045) );
  XOR U128 ( .A(n14726), .B(n14727), .Z(n14816) );
  XOR U129 ( .A(n11147), .B(n11148), .Z(n11531) );
  XNOR U130 ( .A(n7747), .B(n7748), .Z(n8130) );
  XNOR U131 ( .A(n6498), .B(n6499), .Z(n7067) );
  XNOR U132 ( .A(n7288), .B(n7289), .Z(n7761) );
  XNOR U133 ( .A(n6816), .B(n6817), .Z(n6796) );
  XNOR U134 ( .A(n7759), .B(n7760), .Z(n8142) );
  XNOR U135 ( .A(n6508), .B(n6509), .Z(n7063) );
  XOR U136 ( .A(n15482), .B(n15483), .Z(n15596) );
  XNOR U137 ( .A(n7296), .B(n7297), .Z(n7773) );
  XOR U138 ( .A(n12683), .B(n12684), .Z(n13073) );
  XNOR U139 ( .A(n7771), .B(n7772), .Z(n8154) );
  XOR U140 ( .A(n6274), .B(n6275), .Z(n6518) );
  XOR U141 ( .A(n4202), .B(n4203), .Z(n4241) );
  XNOR U142 ( .A(n7304), .B(n7305), .Z(n7785) );
  XNOR U143 ( .A(n3674), .B(n3675), .Z(n3594) );
  XOR U144 ( .A(n16238), .B(n16239), .Z(n16316) );
  XOR U145 ( .A(n16369), .B(n16370), .Z(n16372) );
  XNOR U146 ( .A(n7783), .B(n7784), .Z(n8166) );
  XNOR U147 ( .A(n16305), .B(n16306), .Z(n16700) );
  XNOR U148 ( .A(n7312), .B(n7313), .Z(n7797) );
  XNOR U149 ( .A(n5194), .B(n5195), .Z(n5236) );
  XNOR U150 ( .A(n4782), .B(n4783), .Z(n4936) );
  XOR U151 ( .A(n16722), .B(n16723), .Z(n17084) );
  XOR U152 ( .A(n16625), .B(n16626), .Z(n16751) );
  XOR U153 ( .A(n14225), .B(n14226), .Z(n14609) );
  XNOR U154 ( .A(n7795), .B(n7796), .Z(n8178) );
  XNOR U155 ( .A(n6540), .B(n6541), .Z(n7051) );
  XNOR U156 ( .A(n4222), .B(n4223), .Z(n4225) );
  XNOR U157 ( .A(n4910), .B(n4911), .Z(n4818) );
  XNOR U158 ( .A(n16287), .B(n16288), .Z(n16684) );
  NAND U159 ( .A(b[12]), .B(a[17]), .Z(n17080) );
  XNOR U160 ( .A(n7320), .B(n7321), .Z(n7809) );
  XNOR U161 ( .A(n16690), .B(n16691), .Z(n17051) );
  XNOR U162 ( .A(n7807), .B(n7808), .Z(n8190) );
  XOR U163 ( .A(n5234), .B(n5235), .Z(n5515) );
  XNOR U164 ( .A(n6920), .B(n6921), .Z(n6922) );
  XOR U165 ( .A(n15761), .B(n15762), .Z(n16147) );
  XNOR U166 ( .A(n7819), .B(n7820), .Z(n8202) );
  XOR U167 ( .A(n6268), .B(n6269), .Z(n6270) );
  XNOR U168 ( .A(n4804), .B(n4805), .Z(n4927) );
  XNOR U169 ( .A(n7336), .B(n7337), .Z(n7833) );
  XNOR U170 ( .A(n5548), .B(n5549), .Z(n5550) );
  XNOR U171 ( .A(n7831), .B(n7832), .Z(n8214) );
  XNOR U172 ( .A(n5530), .B(n5531), .Z(n5532) );
  XNOR U173 ( .A(n7344), .B(n7345), .Z(n7845) );
  XNOR U174 ( .A(n5545), .B(n5544), .Z(n5536) );
  XOR U175 ( .A(n16932), .B(n16933), .Z(n17302) );
  XNOR U176 ( .A(n7843), .B(n7844), .Z(n8226) );
  XNOR U177 ( .A(n6578), .B(n6579), .Z(n7034) );
  XNOR U178 ( .A(n7352), .B(n7353), .Z(n7857) );
  XOR U179 ( .A(n18966), .B(n18967), .Z(n19342) );
  XNOR U180 ( .A(n7855), .B(n7856), .Z(n8238) );
  XNOR U181 ( .A(n6600), .B(n6601), .Z(n6602) );
  XOR U182 ( .A(n19361), .B(n19362), .Z(n19753) );
  XNOR U183 ( .A(n7360), .B(n7361), .Z(n7869) );
  XNOR U184 ( .A(n19353), .B(n19354), .Z(n19748) );
  XOR U185 ( .A(n16952), .B(n16953), .Z(n17326) );
  XNOR U186 ( .A(n7867), .B(n7868), .Z(n8250) );
  XNOR U187 ( .A(n19746), .B(n19747), .Z(n20131) );
  XOR U188 ( .A(n19220), .B(n19221), .Z(n19602) );
  XNOR U189 ( .A(n7368), .B(n7369), .Z(n7881) );
  XOR U190 ( .A(n20127), .B(n20128), .Z(n20505) );
  XNOR U191 ( .A(n20161), .B(n20162), .Z(n20538) );
  XNOR U192 ( .A(n7879), .B(n7880), .Z(n8262) );
  XNOR U193 ( .A(n7376), .B(n7377), .Z(n7893) );
  XNOR U194 ( .A(n20474), .B(n20475), .Z(n20852) );
  XOR U195 ( .A(n20769), .B(n20770), .Z(n20929) );
  XOR U196 ( .A(n20750), .B(n20751), .Z(n21133) );
  XOR U197 ( .A(n8280), .B(n8281), .Z(n8286) );
  XNOR U198 ( .A(n18115), .B(n18116), .Z(n18495) );
  OR U199 ( .A(n23950), .B(n23951), .Z(n5) );
  NANDN U200 ( .A(n23953), .B(n23952), .Z(n6) );
  AND U201 ( .A(n5), .B(n6), .Z(n23959) );
  ANDN U202 ( .B(n15858), .A(n15857), .Z(n21963) );
  XOR U203 ( .A(n24157), .B(n24155), .Z(n7) );
  NAND U204 ( .A(n7), .B(n24154), .Z(n8) );
  NAND U205 ( .A(n24157), .B(n24155), .Z(n9) );
  AND U206 ( .A(n8), .B(n9), .Z(n24159) );
  OR U207 ( .A(n22441), .B(n22442), .Z(n10) );
  NANDN U208 ( .A(n22444), .B(n22443), .Z(n11) );
  AND U209 ( .A(n10), .B(n11), .Z(n22580) );
  OR U210 ( .A(n23374), .B(n23375), .Z(n12) );
  NANDN U211 ( .A(n23377), .B(n23376), .Z(n13) );
  AND U212 ( .A(n12), .B(n13), .Z(n23463) );
  OR U213 ( .A(n23618), .B(n23619), .Z(n14) );
  NANDN U214 ( .A(n23621), .B(n23620), .Z(n15) );
  AND U215 ( .A(n14), .B(n15), .Z(n23693) );
  OR U216 ( .A(n23814), .B(n23815), .Z(n16) );
  NANDN U217 ( .A(n23817), .B(n23816), .Z(n17) );
  AND U218 ( .A(n16), .B(n17), .Z(n23869) );
  OR U219 ( .A(n23954), .B(n23955), .Z(n18) );
  NANDN U220 ( .A(n23957), .B(n23956), .Z(n19) );
  AND U221 ( .A(n18), .B(n19), .Z(n23993) );
  OR U222 ( .A(n24044), .B(n24045), .Z(n20) );
  NANDN U223 ( .A(n24047), .B(n24046), .Z(n21) );
  AND U224 ( .A(n20), .B(n21), .Z(n24065) );
  XNOR U225 ( .A(n768), .B(n769), .Z(n771) );
  XNOR U226 ( .A(n520), .B(n521), .Z(n594) );
  XNOR U227 ( .A(n382), .B(n383), .Z(n422) );
  XNOR U228 ( .A(n1186), .B(n1187), .Z(n1290) );
  XNOR U229 ( .A(n1034), .B(n1035), .Z(n1132) );
  XNOR U230 ( .A(n7563), .B(n7564), .Z(n7944) );
  XNOR U231 ( .A(n7587), .B(n7588), .Z(n7966) );
  XNOR U232 ( .A(n792), .B(n793), .Z(n976) );
  XNOR U233 ( .A(n1352), .B(n1353), .Z(n1564) );
  XNOR U234 ( .A(n1194), .B(n1195), .Z(n1286) );
  XNOR U235 ( .A(n592), .B(n593), .Z(n656) );
  XOR U236 ( .A(n538), .B(n539), .Z(n541) );
  XNOR U237 ( .A(n442), .B(n443), .Z(n544) );
  XOR U238 ( .A(n8338), .B(n8339), .Z(n8341) );
  XNOR U239 ( .A(n1874), .B(n1875), .Z(n2125) );
  XNOR U240 ( .A(n5052), .B(n5053), .Z(n5364) );
  XNOR U241 ( .A(n3256), .B(n3257), .Z(n3806) );
  XNOR U242 ( .A(n1050), .B(n1051), .Z(n1124) );
  XOR U243 ( .A(n8362), .B(n8363), .Z(n8365) );
  XNOR U244 ( .A(n344), .B(n345), .Z(n370) );
  XNOR U245 ( .A(n5952), .B(n5953), .Z(n6402) );
  XNOR U246 ( .A(n7992), .B(n7993), .Z(n8375) );
  XNOR U247 ( .A(n5062), .B(n5063), .Z(n5377) );
  XOR U248 ( .A(n1884), .B(n1885), .Z(n2219) );
  XOR U249 ( .A(n1560), .B(n1561), .Z(n1649) );
  XNOR U250 ( .A(n820), .B(n821), .Z(n968) );
  XNOR U251 ( .A(n674), .B(n675), .Z(n677) );
  XNOR U252 ( .A(n5958), .B(n5959), .Z(n6310) );
  XNOR U253 ( .A(n7623), .B(n7624), .Z(n8002) );
  XNOR U254 ( .A(n4648), .B(n4649), .Z(n4976) );
  XNOR U255 ( .A(n4080), .B(n4081), .Z(n4296) );
  XNOR U256 ( .A(n3038), .B(n3039), .Z(n3278) );
  XOR U257 ( .A(n2636), .B(n2637), .Z(n2639) );
  XNOR U258 ( .A(n2216), .B(n2217), .Z(n2346) );
  XOR U259 ( .A(n1370), .B(n1371), .Z(n1372) );
  XOR U260 ( .A(n1214), .B(n1215), .Z(n1376) );
  XNOR U261 ( .A(n9142), .B(n9143), .Z(n9526) );
  XNOR U262 ( .A(n1066), .B(n1067), .Z(n1222) );
  XNOR U263 ( .A(n9816), .B(n9817), .Z(n10195) );
  XNOR U264 ( .A(n2228), .B(n2229), .Z(n2340) );
  XOR U265 ( .A(n1898), .B(n1899), .Z(n1901) );
  XNOR U266 ( .A(n8014), .B(n8015), .Z(n8399) );
  XNOR U267 ( .A(n3290), .B(n3291), .Z(n3838) );
  XNOR U268 ( .A(n1074), .B(n1075), .Z(n1076) );
  XNOR U269 ( .A(n10191), .B(n10192), .Z(n10578) );
  XNOR U270 ( .A(n10261), .B(n10262), .Z(n10651) );
  XNOR U271 ( .A(n8779), .B(n8780), .Z(n8781) );
  XNOR U272 ( .A(n7647), .B(n7648), .Z(n8026) );
  XNOR U273 ( .A(n3056), .B(n3057), .Z(n3298) );
  XNOR U274 ( .A(n2746), .B(n2747), .Z(n2940) );
  XNOR U275 ( .A(n2456), .B(n2457), .Z(n2627) );
  XNOR U276 ( .A(n1668), .B(n1669), .Z(n1789) );
  XNOR U277 ( .A(n10574), .B(n10575), .Z(n10957) );
  XNOR U278 ( .A(n4968), .B(n4969), .Z(n5086) );
  XNOR U279 ( .A(n3060), .B(n3061), .Z(n3180) );
  XOR U280 ( .A(n1546), .B(n1547), .Z(n1549) );
  XOR U281 ( .A(n4104), .B(n4105), .Z(n4289) );
  XNOR U282 ( .A(n5988), .B(n5989), .Z(n6434) );
  XNOR U283 ( .A(n1402), .B(n1403), .Z(n1540) );
  XNOR U284 ( .A(n10969), .B(n10970), .Z(n11350) );
  XOR U285 ( .A(n9557), .B(n9558), .Z(n9940) );
  XOR U286 ( .A(n2332), .B(n2333), .Z(n2762) );
  XNOR U287 ( .A(n894), .B(n895), .Z(n889) );
  XNOR U288 ( .A(n1466), .B(n1467), .Z(n1446) );
  XNOR U289 ( .A(n11378), .B(n11379), .Z(n11381) );
  XNOR U290 ( .A(n4114), .B(n4115), .Z(n4284) );
  XNOR U291 ( .A(n3074), .B(n3075), .Z(n3316) );
  XNOR U292 ( .A(n3856), .B(n3857), .Z(n3976) );
  XNOR U293 ( .A(n1252), .B(n1253), .Z(n1416) );
  XNOR U294 ( .A(n11334), .B(n11335), .Z(n11710) );
  XNOR U295 ( .A(n11344), .B(n11345), .Z(n11721) );
  XNOR U296 ( .A(n8428), .B(n8429), .Z(n8816) );
  XNOR U297 ( .A(n9190), .B(n9191), .Z(n9574) );
  XNOR U298 ( .A(n10704), .B(n10705), .Z(n11088) );
  XNOR U299 ( .A(n4690), .B(n4691), .Z(n5112) );
  XNOR U300 ( .A(n3314), .B(n3315), .Z(n3716) );
  XOR U301 ( .A(n5850), .B(n5851), .Z(n5853) );
  XNOR U302 ( .A(n2256), .B(n2257), .Z(n2323) );
  XNOR U303 ( .A(n11699), .B(n11700), .Z(n12090) );
  XNOR U304 ( .A(n11715), .B(n11716), .Z(n12108) );
  XNOR U305 ( .A(n4430), .B(n4431), .Z(n4698) );
  XNOR U306 ( .A(n4122), .B(n4123), .Z(n4280) );
  XNOR U307 ( .A(n3086), .B(n3087), .Z(n3170) );
  XOR U308 ( .A(n2772), .B(n2773), .Z(n2774) );
  XNOR U309 ( .A(n1930), .B(n1931), .Z(n2266) );
  XNOR U310 ( .A(n12086), .B(n12087), .Z(n12469) );
  XOR U311 ( .A(n12156), .B(n12157), .Z(n12539) );
  XNOR U312 ( .A(n12160), .B(n12161), .Z(n12163) );
  XNOR U313 ( .A(n6006), .B(n6007), .Z(n6460) );
  XNOR U314 ( .A(n5430), .B(n5431), .Z(n5845) );
  XNOR U315 ( .A(n12138), .B(n12139), .Z(n12524) );
  XOR U316 ( .A(n7695), .B(n7696), .Z(n8075) );
  XNOR U317 ( .A(n4132), .B(n4133), .Z(n4274) );
  XNOR U318 ( .A(n12465), .B(n12466), .Z(n12852) );
  XNOR U319 ( .A(n12481), .B(n12482), .Z(n12870) );
  XOR U320 ( .A(n12521), .B(n12522), .Z(n12911) );
  XNOR U321 ( .A(n11480), .B(n11481), .Z(n11858) );
  XNOR U322 ( .A(n7252), .B(n7253), .Z(n7705) );
  XNOR U323 ( .A(n8080), .B(n8081), .Z(n8464) );
  XNOR U324 ( .A(n6014), .B(n6015), .Z(n6472) );
  XOR U325 ( .A(n3342), .B(n3343), .Z(n3885) );
  XNOR U326 ( .A(n2488), .B(n2489), .Z(n2612) );
  XNOR U327 ( .A(n1942), .B(n1943), .Z(n2099) );
  XOR U328 ( .A(n12833), .B(n12834), .Z(n12923) );
  XOR U329 ( .A(n12944), .B(n12945), .Z(n12947) );
  XNOR U330 ( .A(n7707), .B(n7708), .Z(n8086) );
  XNOR U331 ( .A(n4142), .B(n4143), .Z(n4272) );
  XOR U332 ( .A(n5840), .B(n5841), .Z(n6019) );
  XOR U333 ( .A(n3102), .B(n3103), .Z(n3105) );
  XNOR U334 ( .A(n2492), .B(n2493), .Z(n2794) );
  XNOR U335 ( .A(n1712), .B(n1713), .Z(n1952) );
  XNOR U336 ( .A(n12848), .B(n12849), .Z(n13233) );
  XNOR U337 ( .A(n12864), .B(n12865), .Z(n13251) );
  XNOR U338 ( .A(n12876), .B(n12877), .Z(n13262) );
  XNOR U339 ( .A(n7260), .B(n7261), .Z(n7717) );
  XOR U340 ( .A(n8094), .B(n8095), .Z(n8477) );
  XNOR U341 ( .A(n5138), .B(n5139), .Z(n5264) );
  XNOR U342 ( .A(n4718), .B(n4719), .Z(n4959) );
  XOR U343 ( .A(n5836), .B(n5837), .Z(n5839) );
  XNOR U344 ( .A(n13245), .B(n13246), .Z(n13630) );
  XOR U345 ( .A(n13329), .B(n13330), .Z(n13717) );
  XNOR U346 ( .A(n7719), .B(n7720), .Z(n8098) );
  XNOR U347 ( .A(n3624), .B(n3625), .Z(n3626) );
  XNOR U348 ( .A(n13229), .B(n13230), .Z(n13612) );
  XNOR U349 ( .A(n13652), .B(n13653), .Z(n13972) );
  XOR U350 ( .A(n13593), .B(n13594), .Z(n13707) );
  XNOR U351 ( .A(n7268), .B(n7269), .Z(n7729) );
  XOR U352 ( .A(n8106), .B(n8107), .Z(n8489) );
  XOR U353 ( .A(n4728), .B(n4729), .Z(n4955) );
  XOR U354 ( .A(n5832), .B(n5833), .Z(n5834) );
  XNOR U355 ( .A(n5456), .B(n5457), .Z(n5830) );
  XNOR U356 ( .A(n3898), .B(n3899), .Z(n4164) );
  XNOR U357 ( .A(n3120), .B(n3121), .Z(n3364) );
  XNOR U358 ( .A(n2804), .B(n2805), .Z(n2806) );
  XOR U359 ( .A(n9996), .B(n9997), .Z(n10376) );
  XNOR U360 ( .A(n7731), .B(n7732), .Z(n8110) );
  XNOR U361 ( .A(n4460), .B(n4461), .Z(n4536) );
  XNOR U362 ( .A(n2608), .B(n2609), .Z(n2810) );
  XNOR U363 ( .A(n2296), .B(n2297), .Z(n2514) );
  XNOR U364 ( .A(n5596), .B(n5597), .Z(n5599) );
  XNOR U365 ( .A(n13608), .B(n13609), .Z(n13993) );
  XNOR U366 ( .A(n14009), .B(n14010), .Z(n14347) );
  XNOR U367 ( .A(n14027), .B(n14028), .Z(n14404) );
  XNOR U368 ( .A(n12653), .B(n12654), .Z(n13041) );
  XNOR U369 ( .A(n7276), .B(n7277), .Z(n7741) );
  XOR U370 ( .A(n8118), .B(n8119), .Z(n8501) );
  XNOR U371 ( .A(n6036), .B(n6037), .Z(n6280) );
  XNOR U372 ( .A(n2300), .B(n2301), .Z(n2303) );
  XNOR U373 ( .A(n2840), .B(n2841), .Z(n2842) );
  XOR U374 ( .A(n14345), .B(n14346), .Z(n14423) );
  XNOR U375 ( .A(n12280), .B(n12281), .Z(n12283) );
  XNOR U376 ( .A(n7743), .B(n7744), .Z(n8122) );
  XNOR U377 ( .A(n5160), .B(n5161), .Z(n5254) );
  XOR U378 ( .A(n3910), .B(n3911), .Z(n3913) );
  XNOR U379 ( .A(n3372), .B(n3373), .Z(n3375) );
  XNOR U380 ( .A(n13989), .B(n13990), .Z(n14366) );
  XOR U381 ( .A(n14779), .B(n14780), .Z(n14782) );
  XNOR U382 ( .A(n14412), .B(n14413), .Z(n14800) );
  XNOR U383 ( .A(n7284), .B(n7285), .Z(n7753) );
  XOR U384 ( .A(n8130), .B(n8131), .Z(n8513) );
  XNOR U385 ( .A(n4176), .B(n4177), .Z(n4250) );
  XNOR U386 ( .A(n6046), .B(n6047), .Z(n6276) );
  XNOR U387 ( .A(n14362), .B(n14363), .Z(n14745) );
  XOR U388 ( .A(n11530), .B(n11531), .Z(n11906) );
  XNOR U389 ( .A(n7755), .B(n7756), .Z(n8134) );
  XNOR U390 ( .A(n3158), .B(n3159), .Z(n3384) );
  XNOR U391 ( .A(n3142), .B(n3143), .Z(n3388) );
  XNOR U392 ( .A(n6796), .B(n6797), .Z(n6798) );
  XNOR U393 ( .A(n14741), .B(n14742), .Z(n15126) );
  XOR U394 ( .A(n15166), .B(n15167), .Z(n15552) );
  XOR U395 ( .A(n15105), .B(n15106), .Z(n15207) );
  XNOR U396 ( .A(n11917), .B(n11918), .Z(n12310) );
  XNOR U397 ( .A(n7292), .B(n7293), .Z(n7765) );
  XOR U398 ( .A(n8142), .B(n8143), .Z(n8525) );
  XOR U399 ( .A(n6056), .B(n6057), .Z(n6512) );
  XNOR U400 ( .A(n5482), .B(n5483), .Z(n5822) );
  XNOR U401 ( .A(n15122), .B(n15123), .Z(n15505) );
  XOR U402 ( .A(n15486), .B(n15487), .Z(n15576) );
  XNOR U403 ( .A(n7767), .B(n7768), .Z(n8146) );
  XNOR U404 ( .A(n5176), .B(n5177), .Z(n5246) );
  XNOR U405 ( .A(n4762), .B(n4763), .Z(n4943) );
  XNOR U406 ( .A(n4190), .B(n4191), .Z(n4245) );
  XNOR U407 ( .A(n3668), .B(n3669), .Z(n3600) );
  XNOR U408 ( .A(n15501), .B(n15502), .Z(n15880) );
  XNOR U409 ( .A(n7300), .B(n7301), .Z(n7777) );
  XOR U410 ( .A(n8154), .B(n8155), .Z(n8537) );
  XNOR U411 ( .A(n15934), .B(n15935), .Z(n16238) );
  XOR U412 ( .A(n15859), .B(n15860), .Z(n15985) );
  XOR U413 ( .A(n13072), .B(n13073), .Z(n13456) );
  XNOR U414 ( .A(n7779), .B(n7780), .Z(n8158) );
  XNOR U415 ( .A(n4208), .B(n4209), .Z(n4494) );
  XNOR U416 ( .A(n3594), .B(n3595), .Z(n3596) );
  XNOR U417 ( .A(n15876), .B(n15877), .Z(n16255) );
  XOR U418 ( .A(n16236), .B(n16237), .Z(n16350) );
  XNOR U419 ( .A(n7308), .B(n7309), .Z(n7789) );
  XOR U420 ( .A(n8166), .B(n8167), .Z(n8549) );
  XNOR U421 ( .A(n5190), .B(n5191), .Z(n5238) );
  XNOR U422 ( .A(n16251), .B(n16252), .Z(n16648) );
  XNOR U423 ( .A(n16319), .B(n16320), .Z(n16627) );
  XNOR U424 ( .A(n7791), .B(n7792), .Z(n8170) );
  XOR U425 ( .A(n6534), .B(n6535), .Z(n6536) );
  XNOR U426 ( .A(n6078), .B(n6079), .Z(n6272) );
  XNOR U427 ( .A(n4216), .B(n4217), .Z(n4218) );
  XNOR U428 ( .A(n3946), .B(n3947), .Z(n3948) );
  XNOR U429 ( .A(n16297), .B(n16298), .Z(n16694) );
  XNOR U430 ( .A(n16726), .B(n16727), .Z(n16729) );
  XNOR U431 ( .A(n16738), .B(n16739), .Z(n16741) );
  XOR U432 ( .A(n16754), .B(n16755), .Z(n17120) );
  XOR U433 ( .A(n16766), .B(n16767), .Z(n17132) );
  XNOR U434 ( .A(n16770), .B(n16771), .Z(n16773) );
  XNOR U435 ( .A(n16782), .B(n16783), .Z(n16785) );
  XNOR U436 ( .A(n16794), .B(n16795), .Z(n16797) );
  XNOR U437 ( .A(n16806), .B(n16807), .Z(n16809) );
  XNOR U438 ( .A(n16818), .B(n16819), .Z(n16821) );
  XNOR U439 ( .A(n16830), .B(n16831), .Z(n16833) );
  XNOR U440 ( .A(n16842), .B(n16843), .Z(n16845) );
  XNOR U441 ( .A(n16854), .B(n16855), .Z(n16857) );
  XNOR U442 ( .A(n16866), .B(n16867), .Z(n16869) );
  XNOR U443 ( .A(n16878), .B(n16879), .Z(n16881) );
  XOR U444 ( .A(n8178), .B(n8179), .Z(n8561) );
  XNOR U445 ( .A(n5198), .B(n5199), .Z(n5502) );
  OR U446 ( .A(n22189), .B(n22190), .Z(n22) );
  NANDN U447 ( .A(n22192), .B(n22191), .Z(n23) );
  NAND U448 ( .A(n22), .B(n23), .Z(n22412) );
  XNOR U449 ( .A(n16644), .B(n16645), .Z(n17003) );
  XOR U450 ( .A(n14608), .B(n14609), .Z(n14994) );
  XNOR U451 ( .A(n16890), .B(n16891), .Z(n16893) );
  XNOR U452 ( .A(n4792), .B(n4793), .Z(n4932) );
  XOR U453 ( .A(n5508), .B(n5509), .Z(n5511) );
  XNOR U454 ( .A(n5560), .B(n5561), .Z(n5563) );
  XOR U455 ( .A(n17079), .B(n17080), .Z(n17471) );
  XOR U456 ( .A(n17089), .B(n17090), .Z(n17483) );
  XOR U457 ( .A(n17101), .B(n17102), .Z(n17495) );
  XOR U458 ( .A(n17113), .B(n17114), .Z(n17507) );
  XOR U459 ( .A(n17137), .B(n17138), .Z(n17531) );
  XOR U460 ( .A(n17149), .B(n17150), .Z(n17543) );
  XOR U461 ( .A(n17161), .B(n17162), .Z(n17555) );
  XOR U462 ( .A(n17173), .B(n17174), .Z(n17567) );
  XOR U463 ( .A(n17185), .B(n17186), .Z(n17579) );
  XOR U464 ( .A(n17197), .B(n17198), .Z(n17591) );
  XOR U465 ( .A(n17209), .B(n17210), .Z(n17603) );
  XOR U466 ( .A(n17221), .B(n17222), .Z(n17615) );
  XOR U467 ( .A(n17233), .B(n17234), .Z(n17627) );
  XOR U468 ( .A(n17245), .B(n17246), .Z(n17639) );
  XOR U469 ( .A(n17257), .B(n17258), .Z(n17651) );
  XNOR U470 ( .A(n7324), .B(n7325), .Z(n7813) );
  XOR U471 ( .A(n8190), .B(n8191), .Z(n8573) );
  XNOR U472 ( .A(n4512), .B(n4513), .Z(n4515) );
  XNOR U473 ( .A(n4920), .B(n4921), .Z(n4923) );
  XNOR U474 ( .A(n6624), .B(n6625), .Z(n6626) );
  XNOR U475 ( .A(n16999), .B(n17000), .Z(n17388) );
  XNOR U476 ( .A(n17454), .B(n17455), .Z(n17746) );
  XNOR U477 ( .A(n16902), .B(n16903), .Z(n16905) );
  XNOR U478 ( .A(n7815), .B(n7816), .Z(n8194) );
  XNOR U479 ( .A(n7502), .B(n7503), .Z(n7505) );
  XNOR U480 ( .A(n17384), .B(n17385), .Z(n17763) );
  XOR U481 ( .A(n17436), .B(n17437), .Z(n17439) );
  XOR U482 ( .A(n17442), .B(n17443), .Z(n17824) );
  XOR U483 ( .A(n17269), .B(n17270), .Z(n17663) );
  XNOR U484 ( .A(n7332), .B(n7333), .Z(n7825) );
  XOR U485 ( .A(n8202), .B(n8203), .Z(n8585) );
  XNOR U486 ( .A(n6098), .B(n6099), .Z(n6266) );
  XNOR U487 ( .A(n17759), .B(n17760), .Z(n18142) );
  XOR U488 ( .A(n16146), .B(n16147), .Z(n16526) );
  XNOR U489 ( .A(n7827), .B(n7828), .Z(n8206) );
  XNOR U490 ( .A(n18138), .B(n18139), .Z(n18525) );
  XNOR U491 ( .A(n7340), .B(n7341), .Z(n7837) );
  XOR U492 ( .A(n8214), .B(n8215), .Z(n8597) );
  XNOR U493 ( .A(n5222), .B(n5223), .Z(n5224) );
  XOR U494 ( .A(n5550), .B(n5551), .Z(n5662) );
  XNOR U495 ( .A(n5792), .B(n5793), .Z(n5684) );
  OR U496 ( .A(n23002), .B(n23003), .Z(n24) );
  NANDN U497 ( .A(n23005), .B(n23004), .Z(n25) );
  NAND U498 ( .A(n24), .B(n25), .Z(n23121) );
  XNOR U499 ( .A(n18224), .B(n18225), .Z(n18610) );
  XNOR U500 ( .A(n7839), .B(n7840), .Z(n8218) );
  XNOR U501 ( .A(n6110), .B(n6111), .Z(n6576) );
  XNOR U502 ( .A(n5536), .B(n5537), .Z(n6114) );
  XNOR U503 ( .A(n18055), .B(n18056), .Z(n18439) );
  XNOR U504 ( .A(n7348), .B(n7349), .Z(n7849) );
  XNOR U505 ( .A(n6614), .B(n6615), .Z(n6722) );
  XNOR U506 ( .A(n6904), .B(n6905), .Z(n7004) );
  XNOR U507 ( .A(n7420), .B(n7421), .Z(n7516) );
  XNOR U508 ( .A(n22109), .B(n22110), .Z(n22111) );
  XOR U509 ( .A(n19004), .B(n19005), .Z(n19384) );
  XOR U510 ( .A(n8226), .B(n8227), .Z(n8609) );
  XNOR U511 ( .A(n7851), .B(n7852), .Z(n8230) );
  XOR U512 ( .A(n18063), .B(n18064), .Z(n18445) );
  XOR U513 ( .A(n17694), .B(n17695), .Z(n18074) );
  XNOR U514 ( .A(n7356), .B(n7357), .Z(n7861) );
  XNOR U515 ( .A(n6728), .B(n6729), .Z(n6600) );
  OR U516 ( .A(n23410), .B(n23411), .Z(n26) );
  NANDN U517 ( .A(n23413), .B(n23412), .Z(n27) );
  NAND U518 ( .A(n26), .B(n27), .Z(n23509) );
  XNOR U519 ( .A(n19289), .B(n19290), .Z(n19679) );
  XOR U520 ( .A(n19341), .B(n19342), .Z(n19735) );
  XNOR U521 ( .A(n18071), .B(n18072), .Z(n18456) );
  XOR U522 ( .A(n8238), .B(n8239), .Z(n8621) );
  XNOR U523 ( .A(n7863), .B(n7864), .Z(n8242) );
  XOR U524 ( .A(n19684), .B(n19685), .Z(n20072) );
  XOR U525 ( .A(n19752), .B(n19753), .Z(n20138) );
  XOR U526 ( .A(n17704), .B(n17705), .Z(n17706) );
  XOR U527 ( .A(n17319), .B(n17320), .Z(n17713) );
  XNOR U528 ( .A(n7364), .B(n7365), .Z(n7873) );
  XOR U529 ( .A(n8250), .B(n8251), .Z(n8633) );
  XOR U530 ( .A(n6734), .B(n6735), .Z(n6259) );
  XNOR U531 ( .A(n19770), .B(n19771), .Z(n20156) );
  XNOR U532 ( .A(n7875), .B(n7876), .Z(n8254) );
  OR U533 ( .A(n20426), .B(n20427), .Z(n28) );
  NANDN U534 ( .A(n20802), .B(n20803), .Z(n29) );
  NAND U535 ( .A(n28), .B(n29), .Z(n20428) );
  XOR U536 ( .A(n20131), .B(n20132), .Z(n20511) );
  XOR U537 ( .A(n19601), .B(n19602), .Z(n19991) );
  XOR U538 ( .A(n17329), .B(n17330), .Z(n17723) );
  XOR U539 ( .A(n16962), .B(n16963), .Z(n17338) );
  XNOR U540 ( .A(n11668), .B(n11669), .Z(n12045) );
  XOR U541 ( .A(n8262), .B(n8263), .Z(n8645) );
  OR U542 ( .A(n23726), .B(n23727), .Z(n30) );
  NANDN U543 ( .A(n23729), .B(n23728), .Z(n31) );
  NAND U544 ( .A(n30), .B(n31), .Z(n23791) );
  XOR U545 ( .A(n20504), .B(n20505), .Z(n20883) );
  XOR U546 ( .A(n20395), .B(n20396), .Z(n20543) );
  XOR U547 ( .A(n12043), .B(n12044), .Z(n12437) );
  XNOR U548 ( .A(n20488), .B(n20489), .Z(n20864) );
  XOR U549 ( .A(n20399), .B(n20400), .Z(n20523) );
  XNOR U550 ( .A(n22141), .B(n22142), .Z(n22145) );
  XOR U551 ( .A(n20852), .B(n20853), .Z(n21241) );
  XOR U552 ( .A(n20910), .B(n20911), .Z(n21149) );
  XOR U553 ( .A(n21139), .B(n21137), .Z(n32) );
  NAND U554 ( .A(n32), .B(n21136), .Z(n33) );
  NAND U555 ( .A(n21139), .B(n21137), .Z(n34) );
  AND U556 ( .A(n33), .B(n34), .Z(n20763) );
  XOR U557 ( .A(n8656), .B(n8657), .Z(n9043) );
  XNOR U558 ( .A(n21262), .B(n21263), .Z(n21563) );
  XNOR U559 ( .A(n20900), .B(n20901), .Z(n21286) );
  XOR U560 ( .A(n21146), .B(n21147), .Z(n21321) );
  XOR U561 ( .A(n21132), .B(n21133), .Z(n21517) );
  NANDN U562 ( .A(n20761), .B(n20760), .Z(n35) );
  NANDN U563 ( .A(n20383), .B(n20384), .Z(n36) );
  NAND U564 ( .A(n35), .B(n36), .Z(n20389) );
  NANDN U565 ( .A(n17353), .B(n17354), .Z(n37) );
  NANDN U566 ( .A(n16978), .B(n16979), .Z(n38) );
  AND U567 ( .A(n37), .B(n38), .Z(n17362) );
  OR U568 ( .A(n16231), .B(n16230), .Z(n39) );
  NANDN U569 ( .A(n16610), .B(n16609), .Z(n40) );
  NAND U570 ( .A(n39), .B(n40), .Z(n16611) );
  XOR U571 ( .A(n8285), .B(n8286), .Z(n8667) );
  OR U572 ( .A(n23456), .B(n23457), .Z(n41) );
  NANDN U573 ( .A(n23459), .B(n23458), .Z(n42) );
  AND U574 ( .A(n41), .B(n42), .Z(n23465) );
  XNOR U575 ( .A(n21288), .B(n21289), .Z(n21707) );
  XNOR U576 ( .A(n21310), .B(n21311), .Z(n21731) );
  NOR U577 ( .A(n18497), .B(n18496), .Z(n24127) );
  XOR U578 ( .A(n24150), .B(n24151), .Z(n43) );
  NANDN U579 ( .A(n24153), .B(n43), .Z(n44) );
  NAND U580 ( .A(n24150), .B(n24151), .Z(n45) );
  AND U581 ( .A(n44), .B(n45), .Z(n24157) );
  XOR U582 ( .A(n24165), .B(n24162), .Z(n46) );
  NANDN U583 ( .A(n24163), .B(n46), .Z(n47) );
  NAND U584 ( .A(n24165), .B(n24162), .Z(n48) );
  AND U585 ( .A(n47), .B(n48), .Z(n24167) );
  OR U586 ( .A(n21971), .B(n21970), .Z(n49) );
  NANDN U587 ( .A(n24170), .B(n24171), .Z(n50) );
  AND U588 ( .A(n49), .B(n50), .Z(n24172) );
  OR U589 ( .A(n21993), .B(n21992), .Z(n51) );
  NANDN U590 ( .A(n24202), .B(n24203), .Z(n52) );
  NAND U591 ( .A(n51), .B(n52), .Z(n24204) );
  OR U592 ( .A(n22577), .B(n22578), .Z(n53) );
  NANDN U593 ( .A(n22580), .B(n22579), .Z(n54) );
  AND U594 ( .A(n53), .B(n54), .Z(n22584) );
  OR U595 ( .A(n23180), .B(n23181), .Z(n55) );
  NANDN U596 ( .A(n23183), .B(n23182), .Z(n56) );
  AND U597 ( .A(n55), .B(n56), .Z(n23281) );
  OR U598 ( .A(n23460), .B(n23461), .Z(n57) );
  NANDN U599 ( .A(n23463), .B(n23462), .Z(n58) );
  AND U600 ( .A(n57), .B(n58), .Z(n23547) );
  OR U601 ( .A(n23690), .B(n23691), .Z(n59) );
  NANDN U602 ( .A(n23693), .B(n23692), .Z(n60) );
  AND U603 ( .A(n59), .B(n60), .Z(n23757) );
  OR U604 ( .A(n23866), .B(n23867), .Z(n61) );
  NANDN U605 ( .A(n23869), .B(n23868), .Z(n62) );
  AND U606 ( .A(n61), .B(n62), .Z(n23917) );
  OR U607 ( .A(n23990), .B(n23991), .Z(n63) );
  NANDN U608 ( .A(n23993), .B(n23992), .Z(n64) );
  AND U609 ( .A(n63), .B(n64), .Z(n24023) );
  OR U610 ( .A(n24062), .B(n24063), .Z(n65) );
  NANDN U611 ( .A(n24065), .B(n24064), .Z(n66) );
  AND U612 ( .A(n65), .B(n66), .Z(n24078) );
  NAND U613 ( .A(b[54]), .B(a[0]), .Z(n1824) );
  NAND U614 ( .A(b[55]), .B(a[0]), .Z(n1584) );
  NAND U615 ( .A(b[56]), .B(a[0]), .Z(n1306) );
  NAND U616 ( .A(b[57]), .B(a[0]), .Z(n1148) );
  NAND U617 ( .A(b[58]), .B(a[0]), .Z(n994) );
  NAND U618 ( .A(b[59]), .B(a[0]), .Z(n742) );
  NAND U619 ( .A(b[60]), .B(a[0]), .Z(n604) );
  NAND U620 ( .A(b[44]), .B(a[0]), .Z(n5002) );
  NAND U621 ( .A(b[45]), .B(a[0]), .Z(n4580) );
  NAND U622 ( .A(b[46]), .B(a[0]), .Z(n4320) );
  NAND U623 ( .A(b[47]), .B(a[0]), .Z(n4012) );
  NAND U624 ( .A(b[48]), .B(a[0]), .Z(n3752) );
  NAND U625 ( .A(b[49]), .B(a[0]), .Z(n3206) );
  NAND U626 ( .A(b[50]), .B(a[0]), .Z(n2972) );
  NAND U627 ( .A(b[53]), .B(a[0]), .Z(n2146) );
  NAND U628 ( .A(b[52]), .B(a[0]), .Z(n2372) );
  NAND U629 ( .A(b[41]), .B(a[0]), .Z(n6336) );
  XNOR U630 ( .A(n508), .B(n509), .Z(n624) );
  XNOR U631 ( .A(n384), .B(n385), .Z(n387) );
  XOR U632 ( .A(n776), .B(n777), .Z(n1028) );
  XNOR U633 ( .A(n422), .B(n423), .Z(n478) );
  NAND U634 ( .A(b[39]), .B(a[0]), .Z(n7536) );
  XNOR U635 ( .A(n640), .B(n641), .Z(n734) );
  XNOR U636 ( .A(n7948), .B(n7949), .Z(n7950) );
  XNOR U637 ( .A(n1190), .B(n1191), .Z(n1288) );
  XNOR U638 ( .A(n1038), .B(n1039), .Z(n1130) );
  XNOR U639 ( .A(n7944), .B(n7945), .Z(n8327) );
  XNOR U640 ( .A(n7966), .B(n7967), .Z(n8351) );
  XOR U641 ( .A(n976), .B(n977), .Z(n979) );
  XNOR U642 ( .A(n656), .B(n657), .Z(n732) );
  XNOR U643 ( .A(n8344), .B(n8345), .Z(n8732) );
  XNOR U644 ( .A(n1634), .B(n1635), .Z(n1802) );
  XNOR U645 ( .A(n1356), .B(n1357), .Z(n1638) );
  XNOR U646 ( .A(n660), .B(n661), .Z(n663) );
  XNOR U647 ( .A(n544), .B(n545), .Z(n547) );
  XOR U648 ( .A(n6314), .B(n6315), .Z(n6385) );
  XNOR U649 ( .A(n5364), .B(n5365), .Z(n5367) );
  XNOR U650 ( .A(n8691), .B(n8692), .Z(n9077) );
  XNOR U651 ( .A(n8701), .B(n8702), .Z(n9089) );
  XNOR U652 ( .A(n8727), .B(n8728), .Z(n9113) );
  XNOR U653 ( .A(n6388), .B(n6389), .Z(n6391) );
  XNOR U654 ( .A(n7984), .B(n7985), .Z(n7986) );
  XNOR U655 ( .A(n7611), .B(n7612), .Z(n7992) );
  XNOR U656 ( .A(n5056), .B(n5057), .Z(n5059) );
  XNOR U657 ( .A(n4634), .B(n4635), .Z(n4637) );
  XNOR U658 ( .A(n4374), .B(n4375), .Z(n4377) );
  XNOR U659 ( .A(n4066), .B(n4067), .Z(n4069) );
  XNOR U660 ( .A(n3806), .B(n3807), .Z(n3809) );
  XNOR U661 ( .A(n3260), .B(n3261), .Z(n3263) );
  XNOR U662 ( .A(n3026), .B(n3027), .Z(n3029) );
  XOR U663 ( .A(n2204), .B(n2205), .Z(n2438) );
  XNOR U664 ( .A(n1364), .B(n1365), .Z(n1560) );
  XOR U665 ( .A(n370), .B(n371), .Z(n373) );
  XNOR U666 ( .A(n9072), .B(n9073), .Z(n9454) );
  XNOR U667 ( .A(n9106), .B(n9107), .Z(n9490) );
  XNOR U668 ( .A(n8749), .B(n8750), .Z(n9137) );
  XNOR U669 ( .A(n1210), .B(n1211), .Z(n1370) );
  XNOR U670 ( .A(n456), .B(n457), .Z(n459) );
  XNOR U671 ( .A(n9501), .B(n9502), .Z(n9504) );
  XNOR U672 ( .A(n6402), .B(n6403), .Z(n7111) );
  XOR U673 ( .A(n5286), .B(n5287), .Z(n5289) );
  XOR U674 ( .A(n1890), .B(n1891), .Z(n2223) );
  XNOR U675 ( .A(n1062), .B(n1063), .Z(n1118) );
  XNOR U676 ( .A(n824), .B(n825), .Z(n826) );
  XNOR U677 ( .A(n9449), .B(n9450), .Z(n9833) );
  XNOR U678 ( .A(n9483), .B(n9484), .Z(n9869) );
  XOR U679 ( .A(n6310), .B(n6311), .Z(n6313) );
  XNOR U680 ( .A(n8380), .B(n8381), .Z(n8768) );
  XNOR U681 ( .A(n8002), .B(n8003), .Z(n8387) );
  XOR U682 ( .A(n4976), .B(n4977), .Z(n4979) );
  XOR U683 ( .A(n4556), .B(n4557), .Z(n4559) );
  XOR U684 ( .A(n4296), .B(n4297), .Z(n4299) );
  XOR U685 ( .A(n3988), .B(n3989), .Z(n3991) );
  XNOR U686 ( .A(n3278), .B(n3279), .Z(n3281) );
  XOR U687 ( .A(n3042), .B(n3043), .Z(n3045) );
  XOR U688 ( .A(n2346), .B(n2347), .Z(n2348) );
  XNOR U689 ( .A(n1656), .B(n1657), .Z(n1898) );
  XNOR U690 ( .A(n9828), .B(n9829), .Z(n10208) );
  XNOR U691 ( .A(n9850), .B(n9851), .Z(n10232) );
  XNOR U692 ( .A(n9862), .B(n9863), .Z(n10244) );
  XNOR U693 ( .A(n9898), .B(n9899), .Z(n10280) );
  XNOR U694 ( .A(n8008), .B(n8009), .Z(n8010) );
  XNOR U695 ( .A(n7635), .B(n7636), .Z(n8014) );
  XNOR U696 ( .A(n2732), .B(n2733), .Z(n2947) );
  XNOR U697 ( .A(n5388), .B(n5389), .Z(n5863) );
  XNOR U698 ( .A(n1382), .B(n1383), .Z(n1552) );
  XOR U699 ( .A(n1222), .B(n1223), .Z(n1224) );
  XNOR U700 ( .A(n1070), .B(n1071), .Z(n1117) );
  XNOR U701 ( .A(n838), .B(n839), .Z(n1074) );
  XNOR U702 ( .A(n6412), .B(n6413), .Z(n7105) );
  XNOR U703 ( .A(n9531), .B(n9532), .Z(n9917) );
  XNOR U704 ( .A(n5078), .B(n5079), .Z(n5281) );
  XNOR U705 ( .A(n4658), .B(n4659), .Z(n4971) );
  XNOR U706 ( .A(n2452), .B(n2453), .Z(n2628) );
  XNOR U707 ( .A(n716), .B(n717), .Z(n720) );
  XNOR U708 ( .A(n10197), .B(n10198), .Z(n10585) );
  XNOR U709 ( .A(n10203), .B(n10204), .Z(n10591) );
  XNOR U710 ( .A(n10225), .B(n10226), .Z(n10615) );
  XNOR U711 ( .A(n4406), .B(n4407), .Z(n4669) );
  XOR U712 ( .A(n3838), .B(n3839), .Z(n3840) );
  XNOR U713 ( .A(n3294), .B(n3295), .Z(n3724) );
  XOR U714 ( .A(n2236), .B(n2237), .Z(n2460) );
  XNOR U715 ( .A(n1394), .B(n1395), .Z(n1546) );
  XNOR U716 ( .A(n1234), .B(n1235), .Z(n1274) );
  XNOR U717 ( .A(n10610), .B(n10611), .Z(n10992) );
  XNOR U718 ( .A(n10656), .B(n10657), .Z(n11040) );
  XNOR U719 ( .A(n8026), .B(n8027), .Z(n8411) );
  XNOR U720 ( .A(n8406), .B(n8407), .Z(n8792) );
  XNOR U721 ( .A(n5086), .B(n5087), .Z(n5279) );
  XOR U722 ( .A(n3298), .B(n3299), .Z(n3301) );
  XOR U723 ( .A(n2750), .B(n2751), .Z(n3068) );
  XNOR U724 ( .A(n10580), .B(n10581), .Z(n10964) );
  XNOR U725 ( .A(n9549), .B(n9550), .Z(n9551) );
  XNOR U726 ( .A(n9172), .B(n9173), .Z(n9175) );
  XOR U727 ( .A(n7659), .B(n7660), .Z(n8041) );
  XOR U728 ( .A(n4102), .B(n4103), .Z(n4288) );
  XNOR U729 ( .A(n3064), .B(n3065), .Z(n3179) );
  XOR U730 ( .A(n2112), .B(n2113), .Z(n2245) );
  XNOR U731 ( .A(n1912), .B(n1913), .Z(n2111) );
  XNOR U732 ( .A(n1674), .B(n1675), .Z(n1782) );
  XNOR U733 ( .A(n1242), .B(n1243), .Z(n1271) );
  XNOR U734 ( .A(n952), .B(n953), .Z(n932) );
  XNOR U735 ( .A(n10959), .B(n10960), .Z(n11339) );
  XNOR U736 ( .A(n10987), .B(n10988), .Z(n11367) );
  XNOR U737 ( .A(n6430), .B(n6431), .Z(n7097) );
  XNOR U738 ( .A(n6434), .B(n6435), .Z(n6437) );
  XOR U739 ( .A(n4108), .B(n4109), .Z(n4111) );
  XNOR U740 ( .A(n5414), .B(n5415), .Z(n5854) );
  XOR U741 ( .A(n1540), .B(n1541), .Z(n1543) );
  XNOR U742 ( .A(n11362), .B(n11363), .Z(n11738) );
  XOR U743 ( .A(n7671), .B(n7672), .Z(n8053) );
  XNOR U744 ( .A(n5100), .B(n5101), .Z(n5420) );
  XOR U745 ( .A(n4686), .B(n4687), .Z(n5106) );
  XNOR U746 ( .A(n11356), .B(n11357), .Z(n11734) );
  XNOR U747 ( .A(n11761), .B(n11762), .Z(n11764) );
  XNOR U748 ( .A(n9948), .B(n9949), .Z(n10328) );
  XNOR U749 ( .A(n6446), .B(n6447), .Z(n7090) );
  XOR U750 ( .A(n3078), .B(n3079), .Z(n3320) );
  XNOR U751 ( .A(n4118), .B(n4119), .Z(n4282) );
  XNOR U752 ( .A(n3860), .B(n3861), .Z(n3974) );
  XNOR U753 ( .A(n2768), .B(n2769), .Z(n2932) );
  XNOR U754 ( .A(n2474), .B(n2475), .Z(n2772) );
  XNOR U755 ( .A(n1686), .B(n1687), .Z(n1689) );
  XNOR U756 ( .A(n1416), .B(n1417), .Z(n1419) );
  XNOR U757 ( .A(n1258), .B(n1259), .Z(n1268) );
  XNOR U758 ( .A(n1102), .B(n1103), .Z(n1105) );
  XNOR U759 ( .A(n1524), .B(n1525), .Z(n1501) );
  XNOR U760 ( .A(n11705), .B(n11706), .Z(n12097) );
  XNOR U761 ( .A(n11727), .B(n11728), .Z(n12121) );
  XOR U762 ( .A(n11757), .B(n11758), .Z(n12148) );
  XOR U763 ( .A(n7683), .B(n7684), .Z(n8065) );
  XNOR U764 ( .A(n6450), .B(n6451), .Z(n7088) );
  XOR U765 ( .A(n5112), .B(n5113), .Z(n5114) );
  XNOR U766 ( .A(n4694), .B(n4695), .Z(n4962) );
  XOR U767 ( .A(n3716), .B(n3717), .Z(n3865) );
  XOR U768 ( .A(n6002), .B(n6003), .Z(n6454) );
  XNOR U769 ( .A(n2262), .B(n2263), .Z(n2320) );
  XNOR U770 ( .A(n8440), .B(n8441), .Z(n8828) );
  XOR U771 ( .A(n8823), .B(n8824), .Z(n9208) );
  XNOR U772 ( .A(n9579), .B(n9580), .Z(n9965) );
  XNOR U773 ( .A(n11093), .B(n11094), .Z(n11475) );
  XNOR U774 ( .A(n4434), .B(n4435), .Z(n4545) );
  XNOR U775 ( .A(n3326), .B(n3327), .Z(n3714) );
  XOR U776 ( .A(n2266), .B(n2267), .Z(n2268) );
  XNOR U777 ( .A(n1698), .B(n1699), .Z(n1774) );
  XNOR U778 ( .A(n2076), .B(n2077), .Z(n2056) );
  XNOR U779 ( .A(n12092), .B(n12093), .Z(n12476) );
  XNOR U780 ( .A(n12102), .B(n12103), .Z(n12487) );
  XNOR U781 ( .A(n12114), .B(n12115), .Z(n12500) );
  XNOR U782 ( .A(n12551), .B(n12552), .Z(n12554) );
  XOR U783 ( .A(n8074), .B(n8075), .Z(n8076) );
  XOR U784 ( .A(n6460), .B(n6461), .Z(n7085) );
  XNOR U785 ( .A(n5122), .B(n5123), .Z(n5434) );
  XOR U786 ( .A(n6010), .B(n6011), .Z(n6466) );
  XNOR U787 ( .A(n3336), .B(n3337), .Z(n3708) );
  XNOR U788 ( .A(n2572), .B(n2573), .Z(n2576) );
  XNOR U789 ( .A(n12471), .B(n12472), .Z(n12859) );
  XNOR U790 ( .A(n12493), .B(n12494), .Z(n12883) );
  XOR U791 ( .A(n12547), .B(n12548), .Z(n12932) );
  XOR U792 ( .A(n4138), .B(n4139), .Z(n4444) );
  XOR U793 ( .A(n5268), .B(n5269), .Z(n5441) );
  XNOR U794 ( .A(n2786), .B(n2787), .Z(n3102) );
  XNOR U795 ( .A(n1764), .B(n1765), .Z(n1720) );
  XOR U796 ( .A(n12910), .B(n12911), .Z(n12913) );
  XOR U797 ( .A(n12956), .B(n12957), .Z(n12959) );
  XOR U798 ( .A(n12968), .B(n12969), .Z(n12971) );
  XOR U799 ( .A(n12980), .B(n12981), .Z(n12983) );
  XOR U800 ( .A(n12992), .B(n12993), .Z(n12995) );
  XOR U801 ( .A(n13004), .B(n13005), .Z(n13007) );
  XOR U802 ( .A(n7705), .B(n7706), .Z(n8087) );
  XOR U803 ( .A(n8464), .B(n8465), .Z(n8466) );
  XOR U804 ( .A(n6472), .B(n6473), .Z(n6474) );
  XNOR U805 ( .A(n5134), .B(n5135), .Z(n5266) );
  XNOR U806 ( .A(n4714), .B(n4715), .Z(n4960) );
  XNOR U807 ( .A(n2612), .B(n2613), .Z(n2615) );
  XNOR U808 ( .A(n1948), .B(n1949), .Z(n2096) );
  XNOR U809 ( .A(n12854), .B(n12855), .Z(n13242) );
  XOR U810 ( .A(n13214), .B(n13215), .Z(n13292) );
  XOR U811 ( .A(n13212), .B(n13213), .Z(n13314) );
  XOR U812 ( .A(n8839), .B(n8840), .Z(n9229) );
  XNOR U813 ( .A(n9603), .B(n9604), .Z(n9989) );
  XNOR U814 ( .A(n11492), .B(n11493), .Z(n11870) );
  XNOR U815 ( .A(n11863), .B(n11864), .Z(n12257) );
  XNOR U816 ( .A(n10357), .B(n10358), .Z(n10747) );
  XNOR U817 ( .A(n4450), .B(n4451), .Z(n4538) );
  XNOR U818 ( .A(n3890), .B(n3891), .Z(n3966) );
  XNOR U819 ( .A(n3352), .B(n3353), .Z(n3704) );
  XNOR U820 ( .A(n2794), .B(n2795), .Z(n2797) );
  XNOR U821 ( .A(n1952), .B(n1953), .Z(n1955) );
  XNOR U822 ( .A(n2082), .B(n2083), .Z(n2038) );
  XNOR U823 ( .A(n13257), .B(n13258), .Z(n13643) );
  XOR U824 ( .A(n13016), .B(n13017), .Z(n13019) );
  XOR U825 ( .A(n7717), .B(n7718), .Z(n8099) );
  XOR U826 ( .A(n8476), .B(n8477), .Z(n8478) );
  XOR U827 ( .A(n6482), .B(n6483), .Z(n6485) );
  XOR U828 ( .A(n6024), .B(n6025), .Z(n6027) );
  XNOR U829 ( .A(n5452), .B(n5453), .Z(n5832) );
  XNOR U830 ( .A(n1970), .B(n1971), .Z(n1972) );
  XNOR U831 ( .A(n3532), .B(n3533), .Z(n3557) );
  XNOR U832 ( .A(n13235), .B(n13236), .Z(n13621) );
  XOR U833 ( .A(n13716), .B(n13717), .Z(n13719) );
  XNOR U834 ( .A(n5146), .B(n5147), .Z(n5260) );
  XOR U835 ( .A(n4456), .B(n4457), .Z(n4732) );
  XNOR U836 ( .A(n3164), .B(n3165), .Z(n3166) );
  XNOR U837 ( .A(n2806), .B(n2807), .Z(n2922) );
  XNOR U838 ( .A(n13638), .B(n13639), .Z(n14024) );
  XNOR U839 ( .A(n13648), .B(n13649), .Z(n14033) );
  XOR U840 ( .A(n13970), .B(n13971), .Z(n14096) );
  XNOR U841 ( .A(n11881), .B(n11882), .Z(n11884) );
  XOR U842 ( .A(n13028), .B(n13029), .Z(n13031) );
  XOR U843 ( .A(n7729), .B(n7730), .Z(n8111) );
  XOR U844 ( .A(n8488), .B(n8489), .Z(n8490) );
  XOR U845 ( .A(n4954), .B(n4955), .Z(n5150) );
  XNOR U846 ( .A(n4160), .B(n4161), .Z(n4262) );
  XNOR U847 ( .A(n6032), .B(n6033), .Z(n6285) );
  XOR U848 ( .A(n4164), .B(n4165), .Z(n4166) );
  XOR U849 ( .A(n3364), .B(n3365), .Z(n3366) );
  XNOR U850 ( .A(n2810), .B(n2811), .Z(n2921) );
  XNOR U851 ( .A(n2510), .B(n2511), .Z(n2606) );
  XNOR U852 ( .A(n3468), .B(n3469), .Z(n3424) );
  XNOR U853 ( .A(n4862), .B(n4863), .Z(n4887) );
  XNOR U854 ( .A(n13614), .B(n13615), .Z(n14002) );
  XNOR U855 ( .A(n14017), .B(n14018), .Z(n14395) );
  XNOR U856 ( .A(n14041), .B(n14042), .Z(n14345) );
  XOR U857 ( .A(n10375), .B(n10376), .Z(n10767) );
  XNOR U858 ( .A(n3162), .B(n3163), .Z(n3910) );
  XNOR U859 ( .A(n2514), .B(n2515), .Z(n2517) );
  XNOR U860 ( .A(n5599), .B(n5598), .Z(n5622) );
  XOR U861 ( .A(n14392), .B(n14393), .Z(n14780) );
  XNOR U862 ( .A(n14426), .B(n14427), .Z(n14726) );
  XOR U863 ( .A(n13040), .B(n13041), .Z(n13043) );
  XOR U864 ( .A(n7741), .B(n7742), .Z(n8123) );
  XOR U865 ( .A(n8500), .B(n8501), .Z(n8502) );
  XOR U866 ( .A(n6280), .B(n6281), .Z(n6283) );
  XNOR U867 ( .A(n4742), .B(n4743), .Z(n4950) );
  XOR U868 ( .A(n2306), .B(n2307), .Z(n2521) );
  XNOR U869 ( .A(n2596), .B(n2597), .Z(n2528) );
  XNOR U870 ( .A(n5756), .B(n5757), .Z(n5733) );
  XNOR U871 ( .A(n13995), .B(n13996), .Z(n14375) );
  XOR U872 ( .A(n14803), .B(n14804), .Z(n14805) );
  XNOR U873 ( .A(n4746), .B(n4747), .Z(n4748) );
  XNOR U874 ( .A(n5472), .B(n5473), .Z(n5824) );
  XNOR U875 ( .A(n3380), .B(n3381), .Z(n3694) );
  XNOR U876 ( .A(n3420), .B(n3421), .Z(n3481) );
  XNOR U877 ( .A(n14793), .B(n14794), .Z(n15181) );
  XNOR U878 ( .A(n14819), .B(n14820), .Z(n15105) );
  XNOR U879 ( .A(n12671), .B(n12672), .Z(n12674) );
  XOR U880 ( .A(n11911), .B(n11912), .Z(n11913) );
  XOR U881 ( .A(n7753), .B(n7754), .Z(n8135) );
  XOR U882 ( .A(n8512), .B(n8513), .Z(n8900) );
  XNOR U883 ( .A(n6502), .B(n6503), .Z(n7064) );
  XNOR U884 ( .A(n4180), .B(n4181), .Z(n4248) );
  XOR U885 ( .A(n4250), .B(n4251), .Z(n4253) );
  XNOR U886 ( .A(n3384), .B(n3385), .Z(n3693) );
  XNOR U887 ( .A(n3606), .B(n3607), .Z(n3608) );
  XNOR U888 ( .A(n6656), .B(n6657), .Z(n6681) );
  XNOR U889 ( .A(n14368), .B(n14369), .Z(n14754) );
  XOR U890 ( .A(n15160), .B(n15161), .Z(n15162) );
  XNOR U891 ( .A(n15210), .B(n15211), .Z(n15482) );
  XOR U892 ( .A(n11905), .B(n11906), .Z(n12301) );
  XNOR U893 ( .A(n5172), .B(n5173), .Z(n5250) );
  XNOR U894 ( .A(n3388), .B(n3389), .Z(n3391) );
  XNOR U895 ( .A(n3506), .B(n3507), .Z(n3508) );
  XNOR U896 ( .A(n14747), .B(n14748), .Z(n15135) );
  XOR U897 ( .A(n15551), .B(n15552), .Z(n15554) );
  XNOR U898 ( .A(n11548), .B(n11549), .Z(n11923) );
  XOR U899 ( .A(n12310), .B(n12311), .Z(n12312) );
  XOR U900 ( .A(n7765), .B(n7766), .Z(n8147) );
  XOR U901 ( .A(n8524), .B(n8525), .Z(n8911) );
  XOR U902 ( .A(n4478), .B(n4479), .Z(n4766) );
  XNOR U903 ( .A(n6060), .B(n6061), .Z(n6274) );
  XOR U904 ( .A(n5246), .B(n5247), .Z(n5248) );
  XNOR U905 ( .A(n3150), .B(n3151), .Z(n3155) );
  XNOR U906 ( .A(n6212), .B(n6213), .Z(n6168) );
  XNOR U907 ( .A(n6976), .B(n6977), .Z(n6953) );
  XNOR U908 ( .A(n15128), .B(n15129), .Z(n15514) );
  XNOR U909 ( .A(n15599), .B(n15600), .Z(n15859) );
  XNOR U910 ( .A(n13830), .B(n13831), .Z(n14214) );
  XNOR U911 ( .A(n5180), .B(n5181), .Z(n5244) );
  XNOR U912 ( .A(n4196), .B(n4197), .Z(n4242) );
  XNOR U913 ( .A(n15507), .B(n15508), .Z(n15889) );
  XOR U914 ( .A(n15863), .B(n15864), .Z(n15965) );
  XOR U915 ( .A(n15988), .B(n15989), .Z(n16370) );
  XNOR U916 ( .A(n11560), .B(n11561), .Z(n11935) );
  XOR U917 ( .A(n12322), .B(n12323), .Z(n12324) );
  XOR U918 ( .A(n7777), .B(n7778), .Z(n8159) );
  XOR U919 ( .A(n8536), .B(n8537), .Z(n8924) );
  XNOR U920 ( .A(n6524), .B(n6525), .Z(n7057) );
  XNOR U921 ( .A(n3936), .B(n3937), .Z(n3956) );
  XNOR U922 ( .A(n4904), .B(n4905), .Z(n4832) );
  XNOR U923 ( .A(n5640), .B(n5641), .Z(n5572) );
  XNOR U924 ( .A(n22039), .B(n22040), .Z(n22064) );
  XNOR U925 ( .A(n15882), .B(n15883), .Z(n16264) );
  XOR U926 ( .A(n13455), .B(n13456), .Z(n13845) );
  XNOR U927 ( .A(n6074), .B(n6075), .Z(n6534) );
  XNOR U928 ( .A(n5494), .B(n5495), .Z(n5816) );
  XOR U929 ( .A(n4494), .B(n4495), .Z(n4496) );
  XNOR U930 ( .A(n6636), .B(n6637), .Z(n6638) );
  XNOR U931 ( .A(n11572), .B(n11573), .Z(n11947) );
  XOR U932 ( .A(n12334), .B(n12335), .Z(n12336) );
  XOR U933 ( .A(n7789), .B(n7790), .Z(n8171) );
  XOR U934 ( .A(n8548), .B(n8549), .Z(n8937) );
  XOR U935 ( .A(n5236), .B(n5237), .Z(n5498) );
  XNOR U936 ( .A(n4218), .B(n4219), .Z(n4236) );
  XNOR U937 ( .A(n3948), .B(n3949), .Z(n4222) );
  XNOR U938 ( .A(n3680), .B(n3681), .Z(n3590) );
  XNOR U939 ( .A(n7456), .B(n7457), .Z(n7496) );
  XNOR U940 ( .A(n16257), .B(n16258), .Z(n16657) );
  XOR U941 ( .A(n16629), .B(n16630), .Z(n16707) );
  XOR U942 ( .A(n16710), .B(n16711), .Z(n16984) );
  XOR U943 ( .A(n16627), .B(n16628), .Z(n16717) );
  XOR U944 ( .A(n7316), .B(n7317), .Z(n7801) );
  XOR U945 ( .A(n5502), .B(n5503), .Z(n5505) );
  XNOR U946 ( .A(n5568), .B(n5569), .Z(n5652) );
  XNOR U947 ( .A(n22075), .B(n22076), .Z(n22031) );
  XNOR U948 ( .A(n16650), .B(n16651), .Z(n17012) );
  XOR U949 ( .A(n16694), .B(n16695), .Z(n16696) );
  XNOR U950 ( .A(n17083), .B(n17084), .Z(n17086) );
  XNOR U951 ( .A(n17095), .B(n17096), .Z(n17098) );
  XNOR U952 ( .A(n17107), .B(n17108), .Z(n17110) );
  XOR U953 ( .A(n17119), .B(n17120), .Z(n17122) );
  XNOR U954 ( .A(n17131), .B(n17132), .Z(n17134) );
  XNOR U955 ( .A(n17143), .B(n17144), .Z(n17146) );
  XNOR U956 ( .A(n17155), .B(n17156), .Z(n17158) );
  XNOR U957 ( .A(n17167), .B(n17168), .Z(n17170) );
  XNOR U958 ( .A(n17179), .B(n17180), .Z(n17182) );
  XNOR U959 ( .A(n17191), .B(n17192), .Z(n17194) );
  XNOR U960 ( .A(n17203), .B(n17204), .Z(n17206) );
  XNOR U961 ( .A(n17215), .B(n17216), .Z(n17218) );
  XNOR U962 ( .A(n17227), .B(n17228), .Z(n17230) );
  XNOR U963 ( .A(n17239), .B(n17240), .Z(n17242) );
  XNOR U964 ( .A(n17251), .B(n17252), .Z(n17254) );
  XNOR U965 ( .A(n11584), .B(n11585), .Z(n11959) );
  XOR U966 ( .A(n12346), .B(n12347), .Z(n12348) );
  XNOR U967 ( .A(n7803), .B(n7804), .Z(n8182) );
  XOR U968 ( .A(n8560), .B(n8561), .Z(n8948) );
  XNOR U969 ( .A(n6544), .B(n6545), .Z(n6547) );
  XNOR U970 ( .A(n4230), .B(n4231), .Z(n4512) );
  XNOR U971 ( .A(n6632), .B(n6633), .Z(n6704) );
  XOR U972 ( .A(n14993), .B(n14994), .Z(n15381) );
  XNOR U973 ( .A(n5206), .B(n5207), .Z(n5234) );
  XNOR U974 ( .A(n4916), .B(n4917), .Z(n4920) );
  XNOR U975 ( .A(n5563), .B(n5562), .Z(n5658) );
  OR U976 ( .A(n22477), .B(n22478), .Z(n67) );
  NANDN U977 ( .A(n22479), .B(n22480), .Z(n68) );
  NAND U978 ( .A(n67), .B(n68), .Z(n22636) );
  XNOR U979 ( .A(n17005), .B(n17006), .Z(n17397) );
  XOR U980 ( .A(n17043), .B(n17044), .Z(n17437) );
  XOR U981 ( .A(n17482), .B(n17483), .Z(n17485) );
  XOR U982 ( .A(n17494), .B(n17495), .Z(n17497) );
  XOR U983 ( .A(n17506), .B(n17507), .Z(n17509) );
  XOR U984 ( .A(n17530), .B(n17531), .Z(n17533) );
  XOR U985 ( .A(n17542), .B(n17543), .Z(n17545) );
  XOR U986 ( .A(n17554), .B(n17555), .Z(n17557) );
  XOR U987 ( .A(n17566), .B(n17567), .Z(n17569) );
  XOR U988 ( .A(n17578), .B(n17579), .Z(n17581) );
  XOR U989 ( .A(n17590), .B(n17591), .Z(n17593) );
  XOR U990 ( .A(n17602), .B(n17603), .Z(n17605) );
  XOR U991 ( .A(n17614), .B(n17615), .Z(n17617) );
  XOR U992 ( .A(n17626), .B(n17627), .Z(n17629) );
  XOR U993 ( .A(n17638), .B(n17639), .Z(n17641) );
  XNOR U994 ( .A(n17263), .B(n17264), .Z(n17266) );
  XOR U995 ( .A(n17650), .B(n17651), .Z(n17653) );
  XNOR U996 ( .A(n11596), .B(n11597), .Z(n11971) );
  XOR U997 ( .A(n12358), .B(n12359), .Z(n12360) );
  XOR U998 ( .A(n7813), .B(n7814), .Z(n8195) );
  XOR U999 ( .A(n8572), .B(n8573), .Z(n8960) );
  XNOR U1000 ( .A(n6094), .B(n6095), .Z(n6268) );
  XOR U1001 ( .A(n17746), .B(n17747), .Z(n17835) );
  XNOR U1002 ( .A(n17460), .B(n17461), .Z(n17839) );
  XNOR U1003 ( .A(n17472), .B(n17473), .Z(n17854) );
  XNOR U1004 ( .A(n17520), .B(n17521), .Z(n17902) );
  XNOR U1005 ( .A(n4812), .B(n4813), .Z(n4814) );
  XNOR U1006 ( .A(n6710), .B(n6711), .Z(n6618) );
  XNOR U1007 ( .A(n7505), .B(n7504), .Z(n7432) );
  XNOR U1008 ( .A(n22093), .B(n22094), .Z(n22025) );
  OR U1009 ( .A(n22211), .B(n22212), .Z(n69) );
  NANDN U1010 ( .A(n22214), .B(n22213), .Z(n70) );
  NAND U1011 ( .A(n69), .B(n70), .Z(n22364) );
  XNOR U1012 ( .A(n17390), .B(n17391), .Z(n17772) );
  XOR U1013 ( .A(n17823), .B(n17824), .Z(n17826) );
  XNOR U1014 ( .A(n17847), .B(n17848), .Z(n18231) );
  XOR U1015 ( .A(n17662), .B(n17663), .Z(n17665) );
  XNOR U1016 ( .A(n11608), .B(n11609), .Z(n11983) );
  XOR U1017 ( .A(n12370), .B(n12371), .Z(n12372) );
  XOR U1018 ( .A(n7825), .B(n7826), .Z(n8207) );
  XOR U1019 ( .A(n8584), .B(n8585), .Z(n8972) );
  XNOR U1020 ( .A(n6564), .B(n6565), .Z(n7041) );
  XOR U1021 ( .A(n6102), .B(n6103), .Z(n6568) );
  XNOR U1022 ( .A(n6242), .B(n6243), .Z(n6138) );
  XNOR U1023 ( .A(n6852), .B(n6853), .Z(n6760) );
  XNOR U1024 ( .A(n7000), .B(n7001), .Z(n6916) );
  XNOR U1025 ( .A(n17765), .B(n17766), .Z(n18151) );
  XOR U1026 ( .A(n16525), .B(n16526), .Z(n16923) );
  XNOR U1027 ( .A(n5224), .B(n5225), .Z(n5530) );
  XNOR U1028 ( .A(n18144), .B(n18145), .Z(n18534) );
  XNOR U1029 ( .A(n17676), .B(n17677), .Z(n18055) );
  XNOR U1030 ( .A(n11620), .B(n11621), .Z(n11995) );
  XOR U1031 ( .A(n12382), .B(n12383), .Z(n12384) );
  XOR U1032 ( .A(n7837), .B(n7838), .Z(n8219) );
  XOR U1033 ( .A(n8596), .B(n8597), .Z(n8985) );
  XNOR U1034 ( .A(n5664), .B(n5665), .Z(n5542) );
  XNOR U1035 ( .A(n5684), .B(n5685), .Z(n5676) );
  XNOR U1036 ( .A(n22021), .B(n22022), .Z(n22105) );
  XNOR U1037 ( .A(n18527), .B(n18528), .Z(n18915) );
  XOR U1038 ( .A(n17295), .B(n17296), .Z(n17686) );
  OR U1039 ( .A(n22772), .B(n22773), .Z(n71) );
  NANDN U1040 ( .A(n22775), .B(n22774), .Z(n72) );
  NAND U1041 ( .A(n71), .B(n72), .Z(n22873) );
  OR U1042 ( .A(n23216), .B(n23217), .Z(n73) );
  NANDN U1043 ( .A(n23219), .B(n23218), .Z(n74) );
  NAND U1044 ( .A(n73), .B(n74), .Z(n23339) );
  XNOR U1045 ( .A(n18593), .B(n18594), .Z(n18984) );
  XNOR U1046 ( .A(n11632), .B(n11633), .Z(n12007) );
  XOR U1047 ( .A(n12394), .B(n12395), .Z(n12396) );
  XOR U1048 ( .A(n7849), .B(n7850), .Z(n8231) );
  XNOR U1049 ( .A(n6582), .B(n6583), .Z(n6585) );
  XNOR U1050 ( .A(n7004), .B(n7005), .Z(n7006) );
  XNOR U1051 ( .A(n6606), .B(n6607), .Z(n6608) );
  XNOR U1052 ( .A(n6120), .B(n6121), .Z(n6261) );
  XNOR U1053 ( .A(n7516), .B(n7517), .Z(n7412) );
  XNOR U1054 ( .A(n19000), .B(n19001), .Z(n19377) );
  XOR U1055 ( .A(n19383), .B(n19384), .Z(n19386) );
  XOR U1056 ( .A(n17307), .B(n17308), .Z(n17701) );
  XOR U1057 ( .A(n16942), .B(n16943), .Z(n17314) );
  XOR U1058 ( .A(n8608), .B(n8609), .Z(n8996) );
  XOR U1059 ( .A(n6129), .B(n6128), .Z(n5797) );
  OR U1060 ( .A(n22245), .B(n22246), .Z(n75) );
  NANDN U1061 ( .A(n22248), .B(n22247), .Z(n76) );
  NAND U1062 ( .A(n75), .B(n76), .Z(n22328) );
  XOR U1063 ( .A(n18444), .B(n18445), .Z(n18834) );
  XNOR U1064 ( .A(n11644), .B(n11645), .Z(n12019) );
  XOR U1065 ( .A(n12406), .B(n12407), .Z(n12408) );
  XOR U1066 ( .A(n7861), .B(n7862), .Z(n8243) );
  XOR U1067 ( .A(n6602), .B(n6603), .Z(n6732) );
  XNOR U1068 ( .A(n6870), .B(n6871), .Z(n6742) );
  XNOR U1069 ( .A(n19674), .B(n19675), .Z(n20060) );
  XOR U1070 ( .A(n19734), .B(n19735), .Z(n19737) );
  XOR U1071 ( .A(n18456), .B(n18457), .Z(n18458) );
  XOR U1072 ( .A(n8620), .B(n8621), .Z(n9008) );
  XNOR U1073 ( .A(n6892), .B(n6893), .Z(n7013) );
  OR U1074 ( .A(n23238), .B(n23239), .Z(n77) );
  NANDN U1075 ( .A(n23241), .B(n23240), .Z(n78) );
  NAND U1076 ( .A(n77), .B(n78), .Z(n23303) );
  OR U1077 ( .A(n23580), .B(n23581), .Z(n79) );
  NANDN U1078 ( .A(n23583), .B(n23582), .Z(n80) );
  NAND U1079 ( .A(n79), .B(n80), .Z(n23655) );
  XOR U1080 ( .A(n20071), .B(n20072), .Z(n20074) );
  XOR U1081 ( .A(n20137), .B(n20138), .Z(n20140) );
  OR U1082 ( .A(n13929), .B(n13928), .Z(n81) );
  NANDN U1083 ( .A(n14310), .B(n14309), .Z(n82) );
  NAND U1084 ( .A(n81), .B(n82), .Z(n13933) );
  XNOR U1085 ( .A(n11656), .B(n11657), .Z(n12031) );
  XOR U1086 ( .A(n12418), .B(n12419), .Z(n12420) );
  XOR U1087 ( .A(n7873), .B(n7874), .Z(n8255) );
  XOR U1088 ( .A(n8632), .B(n8633), .Z(n9020) );
  XNOR U1089 ( .A(n20055), .B(n20056), .Z(n20435) );
  XNOR U1090 ( .A(n20165), .B(n20166), .Z(n20395) );
  XOR U1091 ( .A(n18468), .B(n18469), .Z(n18470) );
  XOR U1092 ( .A(n17716), .B(n17717), .Z(n17718) );
  OR U1093 ( .A(n10153), .B(n10152), .Z(n83) );
  NANDN U1094 ( .A(n10532), .B(n10531), .Z(n84) );
  NAND U1095 ( .A(n83), .B(n84), .Z(n10157) );
  XOR U1096 ( .A(n7372), .B(n7373), .Z(n7885) );
  XNOR U1097 ( .A(n6880), .B(n6881), .Z(n7022) );
  XNOR U1098 ( .A(n20430), .B(n20431), .Z(n20805) );
  XOR U1099 ( .A(n20510), .B(n20511), .Z(n20513) );
  XNOR U1100 ( .A(n20546), .B(n20547), .Z(n20769) );
  XOR U1101 ( .A(n19990), .B(n19991), .Z(n20378) );
  XOR U1102 ( .A(n12430), .B(n12431), .Z(n12432) );
  XNOR U1103 ( .A(n7887), .B(n7888), .Z(n8266) );
  XOR U1104 ( .A(n8644), .B(n8645), .Z(n9032) );
  OR U1105 ( .A(n21193), .B(n21192), .Z(n85) );
  NANDN U1106 ( .A(n20800), .B(n20801), .Z(n86) );
  AND U1107 ( .A(n85), .B(n86), .Z(n20807) );
  XNOR U1108 ( .A(n20470), .B(n20471), .Z(n20844) );
  XOR U1109 ( .A(n20882), .B(n20883), .Z(n20885) );
  XNOR U1110 ( .A(n20532), .B(n20533), .Z(n20910) );
  OR U1111 ( .A(n19247), .B(n19246), .Z(n87) );
  NANDN U1112 ( .A(n19624), .B(n19623), .Z(n88) );
  NAND U1113 ( .A(n87), .B(n88), .Z(n19251) );
  XOR U1114 ( .A(n17728), .B(n17729), .Z(n17730) );
  XOR U1115 ( .A(n17341), .B(n17342), .Z(n17735) );
  OR U1116 ( .A(n13193), .B(n13192), .Z(n89) );
  NANDN U1117 ( .A(n13576), .B(n13575), .Z(n90) );
  NAND U1118 ( .A(n89), .B(n90), .Z(n13197) );
  XOR U1119 ( .A(n12049), .B(n12050), .Z(n12072) );
  XOR U1120 ( .A(n12436), .B(n12437), .Z(n12822) );
  XOR U1121 ( .A(n8274), .B(n8275), .Z(n8657) );
  OR U1122 ( .A(n22279), .B(n22280), .Z(n91) );
  NANDN U1123 ( .A(n22282), .B(n22281), .Z(n92) );
  NAND U1124 ( .A(n91), .B(n92), .Z(n22430) );
  OR U1125 ( .A(n23060), .B(n23061), .Z(n93) );
  NANDN U1126 ( .A(n23063), .B(n23062), .Z(n94) );
  NAND U1127 ( .A(n93), .B(n94), .Z(n23169) );
  OR U1128 ( .A(n23602), .B(n23603), .Z(n95) );
  NANDN U1129 ( .A(n23605), .B(n23604), .Z(n96) );
  NAND U1130 ( .A(n95), .B(n96), .Z(n23679) );
  OR U1131 ( .A(n23850), .B(n23851), .Z(n97) );
  NANDN U1132 ( .A(n23853), .B(n23852), .Z(n98) );
  NAND U1133 ( .A(n97), .B(n98), .Z(n23903) );
  XNOR U1134 ( .A(n20824), .B(n20825), .Z(n21217) );
  XOR U1135 ( .A(n20856), .B(n20857), .Z(n21157) );
  XNOR U1136 ( .A(n20918), .B(n20919), .Z(n21303) );
  XNOR U1137 ( .A(n20932), .B(n20933), .Z(n21146) );
  XOR U1138 ( .A(n20759), .B(n20757), .Z(n99) );
  NANDN U1139 ( .A(n20756), .B(n99), .Z(n100) );
  NAND U1140 ( .A(n20759), .B(n20757), .Z(n101) );
  AND U1141 ( .A(n100), .B(n101), .Z(n20384) );
  NANDN U1142 ( .A(n14708), .B(n14709), .Z(n102) );
  NANDN U1143 ( .A(n14328), .B(n14327), .Z(n103) );
  NAND U1144 ( .A(n102), .B(n103), .Z(n14334) );
  AND U1145 ( .A(a[62]), .B(b[39]), .Z(n22148) );
  XOR U1146 ( .A(n21240), .B(n21241), .Z(n21567) );
  XNOR U1147 ( .A(n21252), .B(n21253), .Z(n21565) );
  XNOR U1148 ( .A(n21282), .B(n21283), .Z(n21559) );
  XNOR U1149 ( .A(n21304), .B(n21305), .Z(n21557) );
  XNOR U1150 ( .A(n21326), .B(n21327), .Z(n21555) );
  XOR U1151 ( .A(n17361), .B(n17362), .Z(n17364) );
  OR U1152 ( .A(n10175), .B(n10174), .Z(n104) );
  NANDN U1153 ( .A(n10179), .B(n10178), .Z(n105) );
  NAND U1154 ( .A(n104), .B(n105), .Z(n10555) );
  XNOR U1155 ( .A(n21634), .B(n21635), .Z(n21636) );
  XNOR U1156 ( .A(n21256), .B(n21257), .Z(n21673) );
  XOR U1157 ( .A(n21286), .B(n21287), .Z(n21706) );
  XOR U1158 ( .A(n21734), .B(n21735), .Z(n21736) );
  XOR U1159 ( .A(n21516), .B(n21517), .Z(n21912) );
  XOR U1160 ( .A(n21525), .B(n21523), .Z(n106) );
  NANDN U1161 ( .A(n21522), .B(n106), .Z(n107) );
  NAND U1162 ( .A(n21525), .B(n21523), .Z(n108) );
  AND U1163 ( .A(n107), .B(n108), .Z(n21145) );
  NAND U1164 ( .A(n17741), .B(n17740), .Z(n109) );
  NANDN U1165 ( .A(n17743), .B(n17742), .Z(n110) );
  AND U1166 ( .A(n109), .B(n110), .Z(n21942) );
  OR U1167 ( .A(n15477), .B(n15476), .Z(n111) );
  NANDN U1168 ( .A(n15481), .B(n15480), .Z(n112) );
  AND U1169 ( .A(n111), .B(n112), .Z(n15478) );
  OR U1170 ( .A(n22830), .B(n22831), .Z(n113) );
  NAND U1171 ( .A(n22833), .B(n22832), .Z(n114) );
  NAND U1172 ( .A(n113), .B(n114), .Z(n22951) );
  ANDN U1173 ( .B(n20394), .A(n20393), .Z(n24105) );
  NAND U1174 ( .A(n24117), .B(n24119), .Z(n24122) );
  NANDN U1175 ( .A(n24146), .B(n24147), .Z(n115) );
  NANDN U1176 ( .A(n21961), .B(n21960), .Z(n116) );
  NAND U1177 ( .A(n115), .B(n116), .Z(n24149) );
  XOR U1178 ( .A(n24159), .B(n24161), .Z(n117) );
  NANDN U1179 ( .A(n24158), .B(n117), .Z(n118) );
  NAND U1180 ( .A(n24159), .B(n24161), .Z(n119) );
  AND U1181 ( .A(n118), .B(n119), .Z(n24165) );
  OR U1182 ( .A(n21969), .B(n21968), .Z(n120) );
  NANDN U1183 ( .A(n24168), .B(n24169), .Z(n121) );
  AND U1184 ( .A(n120), .B(n121), .Z(n24170) );
  NAND U1185 ( .A(n24180), .B(n21975), .Z(n122) );
  ANDN U1186 ( .B(n122), .A(n24179), .Z(n123) );
  NAND U1187 ( .A(n21976), .B(n24175), .Z(n124) );
  NAND U1188 ( .A(n124), .B(n24176), .Z(n125) );
  AND U1189 ( .A(n123), .B(n125), .Z(n126) );
  ANDN U1190 ( .B(n24190), .A(n24187), .Z(n127) );
  NANDN U1191 ( .A(n24182), .B(n21977), .Z(n128) );
  NANDN U1192 ( .A(n126), .B(n127), .Z(n129) );
  NAND U1193 ( .A(n128), .B(n129), .Z(n130) );
  NANDN U1194 ( .A(n24193), .B(n24192), .Z(n131) );
  XNOR U1195 ( .A(n24193), .B(n24192), .Z(n132) );
  NAND U1196 ( .A(n132), .B(n130), .Z(n133) );
  NAND U1197 ( .A(n131), .B(n133), .Z(n24196) );
  OR U1198 ( .A(n21999), .B(n21998), .Z(n134) );
  NANDN U1199 ( .A(n24207), .B(n24206), .Z(n135) );
  AND U1200 ( .A(n134), .B(n135), .Z(n24208) );
  OR U1201 ( .A(n22581), .B(n22582), .Z(n136) );
  NANDN U1202 ( .A(n22584), .B(n22583), .Z(n137) );
  NAND U1203 ( .A(n136), .B(n137), .Z(n22952) );
  OR U1204 ( .A(n23278), .B(n23279), .Z(n138) );
  NANDN U1205 ( .A(n23281), .B(n23280), .Z(n139) );
  AND U1206 ( .A(n138), .B(n139), .Z(n23377) );
  OR U1207 ( .A(n23544), .B(n23545), .Z(n140) );
  NANDN U1208 ( .A(n23547), .B(n23546), .Z(n141) );
  AND U1209 ( .A(n140), .B(n141), .Z(n23621) );
  OR U1210 ( .A(n23754), .B(n23755), .Z(n142) );
  NANDN U1211 ( .A(n23757), .B(n23756), .Z(n143) );
  AND U1212 ( .A(n142), .B(n143), .Z(n23817) );
  OR U1213 ( .A(n23914), .B(n23915), .Z(n144) );
  NANDN U1214 ( .A(n23917), .B(n23916), .Z(n145) );
  AND U1215 ( .A(n144), .B(n145), .Z(n23957) );
  OR U1216 ( .A(n24020), .B(n24021), .Z(n146) );
  NANDN U1217 ( .A(n24023), .B(n24022), .Z(n147) );
  AND U1218 ( .A(n146), .B(n147), .Z(n24047) );
  OR U1219 ( .A(n24075), .B(n24076), .Z(n148) );
  NANDN U1220 ( .A(n24078), .B(n24077), .Z(n149) );
  AND U1221 ( .A(n148), .B(n149), .Z(n24080) );
  IV U1222 ( .A(b[1]), .Z(n150) );
  IV U1223 ( .A(b[2]), .Z(n151) );
  IV U1224 ( .A(b[3]), .Z(n152) );
  IV U1225 ( .A(b[13]), .Z(n153) );
  IV U1226 ( .A(b[40]), .Z(n154) );
  IV U1227 ( .A(b[42]), .Z(n155) );
  IV U1228 ( .A(b[43]), .Z(n156) );
  IV U1229 ( .A(b[51]), .Z(n157) );
  IV U1230 ( .A(b[61]), .Z(n158) );
  IV U1231 ( .A(b[62]), .Z(n159) );
  IV U1232 ( .A(b[63]), .Z(n160) );
  IV U1233 ( .A(a[0]), .Z(n161) );
  IV U1234 ( .A(a[2]), .Z(n162) );
  IV U1235 ( .A(a[4]), .Z(n163) );
  IV U1236 ( .A(a[5]), .Z(n164) );
  IV U1237 ( .A(a[6]), .Z(n165) );
  IV U1238 ( .A(a[7]), .Z(n166) );
  IV U1239 ( .A(a[8]), .Z(n167) );
  IV U1240 ( .A(a[10]), .Z(n168) );
  IV U1241 ( .A(a[12]), .Z(n169) );
  IV U1242 ( .A(a[13]), .Z(n170) );
  IV U1243 ( .A(a[14]), .Z(n171) );
  IV U1244 ( .A(a[15]), .Z(n172) );
  IV U1245 ( .A(a[16]), .Z(n173) );
  IV U1246 ( .A(a[17]), .Z(n174) );
  IV U1247 ( .A(a[18]), .Z(n175) );
  IV U1248 ( .A(a[20]), .Z(n176) );
  IV U1249 ( .A(a[22]), .Z(n177) );
  IV U1250 ( .A(a[24]), .Z(n178) );
  IV U1251 ( .A(a[26]), .Z(n179) );
  IV U1252 ( .A(a[28]), .Z(n180) );
  IV U1253 ( .A(a[30]), .Z(n181) );
  IV U1254 ( .A(a[32]), .Z(n182) );
  IV U1255 ( .A(a[34]), .Z(n183) );
  IV U1256 ( .A(a[35]), .Z(n184) );
  IV U1257 ( .A(a[36]), .Z(n185) );
  IV U1258 ( .A(a[38]), .Z(n186) );
  IV U1259 ( .A(a[39]), .Z(n187) );
  IV U1260 ( .A(a[40]), .Z(n188) );
  IV U1261 ( .A(a[41]), .Z(n189) );
  IV U1262 ( .A(a[42]), .Z(n190) );
  IV U1263 ( .A(a[43]), .Z(n191) );
  IV U1264 ( .A(a[44]), .Z(n192) );
  IV U1265 ( .A(a[45]), .Z(n193) );
  IV U1266 ( .A(a[46]), .Z(n194) );
  IV U1267 ( .A(a[47]), .Z(n195) );
  IV U1268 ( .A(a[48]), .Z(n196) );
  IV U1269 ( .A(a[49]), .Z(n197) );
  IV U1270 ( .A(a[50]), .Z(n198) );
  IV U1271 ( .A(a[51]), .Z(n199) );
  IV U1272 ( .A(a[52]), .Z(n200) );
  IV U1273 ( .A(a[53]), .Z(n201) );
  IV U1274 ( .A(a[54]), .Z(n202) );
  IV U1275 ( .A(a[55]), .Z(n203) );
  IV U1276 ( .A(a[56]), .Z(n204) );
  IV U1277 ( .A(a[57]), .Z(n205) );
  IV U1278 ( .A(a[58]), .Z(n206) );
  IV U1279 ( .A(a[59]), .Z(n207) );
  IV U1280 ( .A(a[60]), .Z(n208) );
  IV U1281 ( .A(a[61]), .Z(n209) );
  IV U1282 ( .A(a[63]), .Z(n210) );
  NAND U1283 ( .A(a[57]), .B(b[40]), .Z(n6735) );
  ANDN U1284 ( .B(b[40]), .A(n204), .Z(n5796) );
  NAND U1285 ( .A(a[54]), .B(b[41]), .Z(n5540) );
  NAND U1286 ( .A(a[53]), .B(b[41]), .Z(n5537) );
  NAND U1287 ( .A(b[42]), .B(a[52]), .Z(n5544) );
  NAND U1288 ( .A(a[51]), .B(b[43]), .Z(n5665) );
  NAND U1289 ( .A(b[45]), .B(a[48]), .Z(n4922) );
  ANDN U1290 ( .B(b[47]), .A(n194), .Z(n4820) );
  NAND U1291 ( .A(a[41]), .B(b[49]), .Z(n3409) );
  NAND U1292 ( .A(a[39]), .B(b[50]), .Z(n2907) );
  NAND U1293 ( .A(a[36]), .B(b[52]), .Z(n2595) );
  NAND U1294 ( .A(a[35]), .B(b[52]), .Z(n1969) );
  IV U1295 ( .A(a[33]), .Z(n21751) );
  ANDN U1296 ( .B(b[53]), .A(n21751), .Z(n1973) );
  IV U1297 ( .A(a[31]), .Z(n21740) );
  ANDN U1298 ( .B(b[54]), .A(n21740), .Z(n1768) );
  ANDN U1299 ( .B(b[55]), .A(n180), .Z(n1436) );
  NAND U1300 ( .A(a[26]), .B(b[57]), .Z(n1443) );
  ANDN U1301 ( .B(b[58]), .A(n177), .Z(n860) );
  ANDN U1302 ( .B(b[59]), .A(n176), .Z(n722) );
  ANDN U1303 ( .B(b[61]), .A(n175), .Z(n704) );
  ANDN U1304 ( .B(b[63]), .A(n172), .Z(n364) );
  ANDN U1305 ( .B(a[16]), .A(n159), .Z(n362) );
  NAND U1306 ( .A(b[62]), .B(a[12]), .Z(n252) );
  AND U1307 ( .A(b[63]), .B(a[11]), .Z(n251) );
  NANDN U1308 ( .A(n252), .B(n251), .Z(n254) );
  NAND U1309 ( .A(b[62]), .B(a[4]), .Z(n212) );
  NAND U1310 ( .A(a[3]), .B(b[63]), .Z(n211) );
  OR U1311 ( .A(n212), .B(n211), .Z(n222) );
  XNOR U1312 ( .A(n212), .B(n211), .Z(n298) );
  NAND U1313 ( .A(b[63]), .B(a[0]), .Z(n283) );
  ANDN U1314 ( .B(a[1]), .A(n159), .Z(n286) );
  NANDN U1315 ( .A(n283), .B(n286), .Z(n215) );
  NAND U1316 ( .A(b[62]), .B(a[2]), .Z(n282) );
  NANDN U1317 ( .A(n161), .B(b[62]), .Z(n398) );
  AND U1318 ( .A(a[1]), .B(n398), .Z(n213) );
  NAND U1319 ( .A(b[63]), .B(n213), .Z(n281) );
  OR U1320 ( .A(n282), .B(n281), .Z(n214) );
  NAND U1321 ( .A(n215), .B(n214), .Z(n216) );
  NAND U1322 ( .A(a[2]), .B(n216), .Z(n220) );
  NAND U1323 ( .A(b[62]), .B(a[3]), .Z(n280) );
  XOR U1324 ( .A(a[2]), .B(n216), .Z(n218) );
  NAND U1325 ( .A(a[2]), .B(n160), .Z(n217) );
  AND U1326 ( .A(n218), .B(n217), .Z(n279) );
  NANDN U1327 ( .A(n280), .B(n279), .Z(n219) );
  NAND U1328 ( .A(n220), .B(n219), .Z(n299) );
  NANDN U1329 ( .A(n298), .B(n299), .Z(n221) );
  NAND U1330 ( .A(n222), .B(n221), .Z(n223) );
  ANDN U1331 ( .B(a[4]), .A(n160), .Z(n224) );
  OR U1332 ( .A(n223), .B(n224), .Z(n226) );
  XOR U1333 ( .A(n224), .B(n223), .Z(n304) );
  NAND U1334 ( .A(a[5]), .B(b[62]), .Z(n305) );
  NAND U1335 ( .A(n304), .B(n305), .Z(n225) );
  AND U1336 ( .A(n226), .B(n225), .Z(n227) );
  ANDN U1337 ( .B(a[5]), .A(n160), .Z(n228) );
  OR U1338 ( .A(n227), .B(n228), .Z(n230) );
  XNOR U1339 ( .A(n228), .B(n227), .Z(n310) );
  ANDN U1340 ( .B(a[6]), .A(n159), .Z(n311) );
  OR U1341 ( .A(n310), .B(n311), .Z(n229) );
  AND U1342 ( .A(n230), .B(n229), .Z(n231) );
  ANDN U1343 ( .B(a[6]), .A(n160), .Z(n232) );
  OR U1344 ( .A(n231), .B(n232), .Z(n234) );
  XNOR U1345 ( .A(n232), .B(n231), .Z(n277) );
  ANDN U1346 ( .B(a[7]), .A(n159), .Z(n278) );
  OR U1347 ( .A(n277), .B(n278), .Z(n233) );
  AND U1348 ( .A(n234), .B(n233), .Z(n235) );
  ANDN U1349 ( .B(a[7]), .A(n160), .Z(n236) );
  OR U1350 ( .A(n235), .B(n236), .Z(n238) );
  XNOR U1351 ( .A(n236), .B(n235), .Z(n275) );
  ANDN U1352 ( .B(a[8]), .A(n159), .Z(n276) );
  OR U1353 ( .A(n275), .B(n276), .Z(n237) );
  AND U1354 ( .A(n238), .B(n237), .Z(n239) );
  ANDN U1355 ( .B(a[8]), .A(n160), .Z(n240) );
  OR U1356 ( .A(n239), .B(n240), .Z(n242) );
  XNOR U1357 ( .A(n240), .B(n239), .Z(n324) );
  ANDN U1358 ( .B(a[9]), .A(n159), .Z(n325) );
  OR U1359 ( .A(n324), .B(n325), .Z(n241) );
  AND U1360 ( .A(n242), .B(n241), .Z(n243) );
  ANDN U1361 ( .B(a[9]), .A(n160), .Z(n244) );
  OR U1362 ( .A(n243), .B(n244), .Z(n246) );
  XNOR U1363 ( .A(n244), .B(n243), .Z(n273) );
  ANDN U1364 ( .B(a[10]), .A(n159), .Z(n274) );
  OR U1365 ( .A(n273), .B(n274), .Z(n245) );
  AND U1366 ( .A(n246), .B(n245), .Z(n247) );
  ANDN U1367 ( .B(a[10]), .A(n160), .Z(n248) );
  OR U1368 ( .A(n247), .B(n248), .Z(n250) );
  XNOR U1369 ( .A(n248), .B(n247), .Z(n271) );
  ANDN U1370 ( .B(a[11]), .A(n159), .Z(n272) );
  OR U1371 ( .A(n271), .B(n272), .Z(n249) );
  NAND U1372 ( .A(n250), .B(n249), .Z(n270) );
  XNOR U1373 ( .A(n252), .B(n251), .Z(n269) );
  NANDN U1374 ( .A(n270), .B(n269), .Z(n253) );
  NAND U1375 ( .A(n254), .B(n253), .Z(n255) );
  ANDN U1376 ( .B(a[12]), .A(n160), .Z(n256) );
  OR U1377 ( .A(n255), .B(n256), .Z(n258) );
  XOR U1378 ( .A(n256), .B(n255), .Z(n342) );
  NAND U1379 ( .A(a[13]), .B(b[62]), .Z(n343) );
  NAND U1380 ( .A(n342), .B(n343), .Z(n257) );
  AND U1381 ( .A(n258), .B(n257), .Z(n259) );
  ANDN U1382 ( .B(b[63]), .A(n170), .Z(n260) );
  OR U1383 ( .A(n259), .B(n260), .Z(n262) );
  XNOR U1384 ( .A(n260), .B(n259), .Z(n348) );
  ANDN U1385 ( .B(a[14]), .A(n159), .Z(n349) );
  OR U1386 ( .A(n348), .B(n349), .Z(n261) );
  AND U1387 ( .A(n262), .B(n261), .Z(n263) );
  ANDN U1388 ( .B(a[15]), .A(n159), .Z(n264) );
  OR U1389 ( .A(n263), .B(n264), .Z(n266) );
  XNOR U1390 ( .A(n264), .B(n263), .Z(n267) );
  ANDN U1391 ( .B(a[14]), .A(n160), .Z(n268) );
  OR U1392 ( .A(n267), .B(n268), .Z(n265) );
  AND U1393 ( .A(n266), .B(n265), .Z(n363) );
  XNOR U1394 ( .A(n362), .B(n363), .Z(n365) );
  XNOR U1395 ( .A(n364), .B(n365), .Z(n358) );
  XNOR U1396 ( .A(n268), .B(n267), .Z(n354) );
  XNOR U1397 ( .A(n270), .B(n269), .Z(n338) );
  XNOR U1398 ( .A(n272), .B(n271), .Z(n335) );
  XNOR U1399 ( .A(n274), .B(n273), .Z(n330) );
  ANDN U1400 ( .B(b[61]), .A(n168), .Z(n326) );
  XNOR U1401 ( .A(n276), .B(n275), .Z(n321) );
  XNOR U1402 ( .A(n278), .B(n277), .Z(n317) );
  NAND U1403 ( .A(a[4]), .B(b[61]), .Z(n295) );
  XNOR U1404 ( .A(n280), .B(n279), .Z(n294) );
  NANDN U1405 ( .A(n295), .B(n294), .Z(n297) );
  XOR U1406 ( .A(n282), .B(n281), .Z(n290) );
  XOR U1407 ( .A(n286), .B(n283), .Z(n285) );
  NAND U1408 ( .A(b[61]), .B(n286), .Z(n284) );
  AND U1409 ( .A(n285), .B(n284), .Z(n289) );
  NANDN U1410 ( .A(n158), .B(a[0]), .Z(n492) );
  ANDN U1411 ( .B(n286), .A(n492), .Z(n401) );
  NAND U1412 ( .A(n160), .B(n401), .Z(n287) );
  NANDN U1413 ( .A(n289), .B(n287), .Z(n397) );
  ANDN U1414 ( .B(b[61]), .A(n162), .Z(n396) );
  OR U1415 ( .A(n397), .B(n396), .Z(n288) );
  NANDN U1416 ( .A(n289), .B(n288), .Z(n291) );
  NANDN U1417 ( .A(n290), .B(n291), .Z(n293) );
  XOR U1418 ( .A(n291), .B(n290), .Z(n394) );
  IV U1419 ( .A(a[3]), .Z(n21580) );
  ANDN U1420 ( .B(b[61]), .A(n21580), .Z(n395) );
  OR U1421 ( .A(n394), .B(n395), .Z(n292) );
  NAND U1422 ( .A(n293), .B(n292), .Z(n393) );
  XNOR U1423 ( .A(n295), .B(n294), .Z(n392) );
  NANDN U1424 ( .A(n393), .B(n392), .Z(n296) );
  NAND U1425 ( .A(n297), .B(n296), .Z(n300) );
  XOR U1426 ( .A(n299), .B(n298), .Z(n301) );
  NANDN U1427 ( .A(n300), .B(n301), .Z(n303) );
  XOR U1428 ( .A(n301), .B(n300), .Z(n389) );
  NANDN U1429 ( .A(n158), .B(a[5]), .Z(n388) );
  NANDN U1430 ( .A(n389), .B(n388), .Z(n302) );
  NAND U1431 ( .A(n303), .B(n302), .Z(n307) );
  NANDN U1432 ( .A(n307), .B(n306), .Z(n309) );
  NAND U1433 ( .A(a[6]), .B(b[61]), .Z(n385) );
  NANDN U1434 ( .A(n385), .B(n384), .Z(n308) );
  NAND U1435 ( .A(n309), .B(n308), .Z(n313) );
  XOR U1436 ( .A(n311), .B(n310), .Z(n312) );
  NANDN U1437 ( .A(n313), .B(n312), .Z(n315) );
  NAND U1438 ( .A(b[61]), .B(a[7]), .Z(n383) );
  NAND U1439 ( .A(n382), .B(n383), .Z(n314) );
  AND U1440 ( .A(n315), .B(n314), .Z(n316) );
  OR U1441 ( .A(n317), .B(n316), .Z(n319) );
  XNOR U1442 ( .A(n317), .B(n316), .Z(n380) );
  ANDN U1443 ( .B(b[61]), .A(n167), .Z(n381) );
  OR U1444 ( .A(n380), .B(n381), .Z(n318) );
  AND U1445 ( .A(n319), .B(n318), .Z(n320) );
  OR U1446 ( .A(n321), .B(n320), .Z(n323) );
  XNOR U1447 ( .A(n321), .B(n320), .Z(n431) );
  IV U1448 ( .A(a[9]), .Z(n21615) );
  ANDN U1449 ( .B(b[61]), .A(n21615), .Z(n430) );
  OR U1450 ( .A(n431), .B(n430), .Z(n322) );
  AND U1451 ( .A(n323), .B(n322), .Z(n327) );
  OR U1452 ( .A(n326), .B(n327), .Z(n329) );
  XNOR U1453 ( .A(n325), .B(n324), .Z(n437) );
  XOR U1454 ( .A(n327), .B(n326), .Z(n436) );
  NANDN U1455 ( .A(n437), .B(n436), .Z(n328) );
  AND U1456 ( .A(n329), .B(n328), .Z(n331) );
  OR U1457 ( .A(n330), .B(n331), .Z(n333) );
  XNOR U1458 ( .A(n331), .B(n330), .Z(n378) );
  NAND U1459 ( .A(b[61]), .B(a[11]), .Z(n379) );
  NANDN U1460 ( .A(n378), .B(n379), .Z(n332) );
  AND U1461 ( .A(n333), .B(n332), .Z(n334) );
  OR U1462 ( .A(n335), .B(n334), .Z(n337) );
  XNOR U1463 ( .A(n335), .B(n334), .Z(n377) );
  ANDN U1464 ( .B(b[61]), .A(n169), .Z(n376) );
  OR U1465 ( .A(n377), .B(n376), .Z(n336) );
  AND U1466 ( .A(n337), .B(n336), .Z(n339) );
  OR U1467 ( .A(n338), .B(n339), .Z(n341) );
  XNOR U1468 ( .A(n339), .B(n338), .Z(n374) );
  ANDN U1469 ( .B(b[61]), .A(n170), .Z(n375) );
  OR U1470 ( .A(n374), .B(n375), .Z(n340) );
  NAND U1471 ( .A(n341), .B(n340), .Z(n345) );
  NANDN U1472 ( .A(n345), .B(n344), .Z(n347) );
  NAND U1473 ( .A(a[14]), .B(b[61]), .Z(n371) );
  NANDN U1474 ( .A(n371), .B(n370), .Z(n346) );
  NAND U1475 ( .A(n347), .B(n346), .Z(n351) );
  ANDN U1476 ( .B(b[61]), .A(n172), .Z(n350) );
  OR U1477 ( .A(n351), .B(n350), .Z(n353) );
  XNOR U1478 ( .A(n349), .B(n348), .Z(n457) );
  XOR U1479 ( .A(n351), .B(n350), .Z(n456) );
  NANDN U1480 ( .A(n457), .B(n456), .Z(n352) );
  AND U1481 ( .A(n353), .B(n352), .Z(n355) );
  OR U1482 ( .A(n354), .B(n355), .Z(n357) );
  XNOR U1483 ( .A(n355), .B(n354), .Z(n463) );
  ANDN U1484 ( .B(b[61]), .A(n173), .Z(n462) );
  OR U1485 ( .A(n463), .B(n462), .Z(n356) );
  AND U1486 ( .A(n357), .B(n356), .Z(n359) );
  OR U1487 ( .A(n358), .B(n359), .Z(n361) );
  XNOR U1488 ( .A(n359), .B(n358), .Z(n368) );
  ANDN U1489 ( .B(b[61]), .A(n174), .Z(n369) );
  OR U1490 ( .A(n368), .B(n369), .Z(n360) );
  AND U1491 ( .A(n361), .B(n360), .Z(n702) );
  ANDN U1492 ( .B(b[63]), .A(n173), .Z(n710) );
  ANDN U1493 ( .B(a[17]), .A(n159), .Z(n708) );
  OR U1494 ( .A(n363), .B(n362), .Z(n367) );
  OR U1495 ( .A(n365), .B(n364), .Z(n366) );
  AND U1496 ( .A(n367), .B(n366), .Z(n709) );
  XNOR U1497 ( .A(n708), .B(n709), .Z(n711) );
  XNOR U1498 ( .A(n710), .B(n711), .Z(n703) );
  XNOR U1499 ( .A(n702), .B(n703), .Z(n705) );
  XNOR U1500 ( .A(n704), .B(n705), .Z(n717) );
  IV U1501 ( .A(a[19]), .Z(n21670) );
  ANDN U1502 ( .B(b[60]), .A(n21670), .Z(n714) );
  XNOR U1503 ( .A(n369), .B(n368), .Z(n469) );
  AND U1504 ( .A(a[15]), .B(b[60]), .Z(n372) );
  NANDN U1505 ( .A(n373), .B(n372), .Z(n455) );
  XOR U1506 ( .A(n373), .B(n372), .Z(n561) );
  XNOR U1507 ( .A(n375), .B(n374), .Z(n450) );
  XNOR U1508 ( .A(n377), .B(n376), .Z(n447) );
  NAND U1509 ( .A(a[12]), .B(b[60]), .Z(n443) );
  XOR U1510 ( .A(n379), .B(n378), .Z(n442) );
  NANDN U1511 ( .A(n443), .B(n442), .Z(n445) );
  XNOR U1512 ( .A(n381), .B(n380), .Z(n427) );
  NAND U1513 ( .A(a[8]), .B(b[60]), .Z(n423) );
  NANDN U1514 ( .A(n423), .B(n422), .Z(n425) );
  NAND U1515 ( .A(b[60]), .B(a[7]), .Z(n386) );
  NANDN U1516 ( .A(n386), .B(n387), .Z(n421) );
  XOR U1517 ( .A(n387), .B(n386), .Z(n480) );
  XNOR U1518 ( .A(n389), .B(n388), .Z(n391) );
  NAND U1519 ( .A(a[6]), .B(b[60]), .Z(n390) );
  OR U1520 ( .A(n391), .B(n390), .Z(n419) );
  XNOR U1521 ( .A(n391), .B(n390), .Z(n514) );
  XOR U1522 ( .A(n393), .B(n392), .Z(n415) );
  XNOR U1523 ( .A(n395), .B(n394), .Z(n410) );
  XNOR U1524 ( .A(n397), .B(n396), .Z(n406) );
  NAND U1525 ( .A(b[61]), .B(a[1]), .Z(n399) );
  NAND U1526 ( .A(n399), .B(n398), .Z(n402) );
  OR U1527 ( .A(n399), .B(n604), .Z(n495) );
  NAND U1528 ( .A(n495), .B(n401), .Z(n400) );
  AND U1529 ( .A(n402), .B(n400), .Z(n405) );
  XOR U1530 ( .A(n495), .B(n401), .Z(n403) );
  NAND U1531 ( .A(n403), .B(n402), .Z(n491) );
  ANDN U1532 ( .B(b[60]), .A(n162), .Z(n490) );
  OR U1533 ( .A(n491), .B(n490), .Z(n404) );
  AND U1534 ( .A(n405), .B(n404), .Z(n407) );
  OR U1535 ( .A(n406), .B(n407), .Z(n409) );
  XNOR U1536 ( .A(n407), .B(n406), .Z(n488) );
  ANDN U1537 ( .B(b[60]), .A(n21580), .Z(n489) );
  OR U1538 ( .A(n488), .B(n489), .Z(n408) );
  AND U1539 ( .A(n409), .B(n408), .Z(n411) );
  OR U1540 ( .A(n410), .B(n411), .Z(n413) );
  XNOR U1541 ( .A(n411), .B(n410), .Z(n486) );
  NAND U1542 ( .A(b[60]), .B(a[4]), .Z(n487) );
  NANDN U1543 ( .A(n486), .B(n487), .Z(n412) );
  NAND U1544 ( .A(n413), .B(n412), .Z(n414) );
  OR U1545 ( .A(n415), .B(n414), .Z(n417) );
  NAND U1546 ( .A(a[5]), .B(b[60]), .Z(n483) );
  XOR U1547 ( .A(n415), .B(n414), .Z(n482) );
  NANDN U1548 ( .A(n483), .B(n482), .Z(n416) );
  NAND U1549 ( .A(n417), .B(n416), .Z(n515) );
  NANDN U1550 ( .A(n514), .B(n515), .Z(n418) );
  NAND U1551 ( .A(n419), .B(n418), .Z(n481) );
  NANDN U1552 ( .A(n480), .B(n481), .Z(n420) );
  AND U1553 ( .A(n421), .B(n420), .Z(n479) );
  NANDN U1554 ( .A(n479), .B(n478), .Z(n424) );
  NAND U1555 ( .A(n425), .B(n424), .Z(n426) );
  OR U1556 ( .A(n427), .B(n426), .Z(n429) );
  XNOR U1557 ( .A(n427), .B(n426), .Z(n477) );
  ANDN U1558 ( .B(b[60]), .A(n21615), .Z(n476) );
  OR U1559 ( .A(n477), .B(n476), .Z(n428) );
  NAND U1560 ( .A(n429), .B(n428), .Z(n432) );
  XOR U1561 ( .A(n431), .B(n430), .Z(n433) );
  OR U1562 ( .A(n432), .B(n433), .Z(n435) );
  NAND U1563 ( .A(a[10]), .B(b[60]), .Z(n533) );
  XOR U1564 ( .A(n433), .B(n432), .Z(n532) );
  NANDN U1565 ( .A(n533), .B(n532), .Z(n434) );
  NAND U1566 ( .A(n435), .B(n434), .Z(n439) );
  NANDN U1567 ( .A(n439), .B(n438), .Z(n441) );
  IV U1568 ( .A(a[11]), .Z(n21164) );
  ANDN U1569 ( .B(b[60]), .A(n21164), .Z(n539) );
  NANDN U1570 ( .A(n539), .B(n538), .Z(n440) );
  NAND U1571 ( .A(n441), .B(n440), .Z(n545) );
  NANDN U1572 ( .A(n545), .B(n544), .Z(n444) );
  NAND U1573 ( .A(n445), .B(n444), .Z(n446) );
  OR U1574 ( .A(n447), .B(n446), .Z(n449) );
  XNOR U1575 ( .A(n447), .B(n446), .Z(n474) );
  ANDN U1576 ( .B(b[60]), .A(n170), .Z(n475) );
  OR U1577 ( .A(n474), .B(n475), .Z(n448) );
  AND U1578 ( .A(n449), .B(n448), .Z(n451) );
  OR U1579 ( .A(n450), .B(n451), .Z(n453) );
  XNOR U1580 ( .A(n451), .B(n450), .Z(n554) );
  NAND U1581 ( .A(b[60]), .B(a[14]), .Z(n555) );
  NANDN U1582 ( .A(n554), .B(n555), .Z(n452) );
  NAND U1583 ( .A(n453), .B(n452), .Z(n560) );
  OR U1584 ( .A(n561), .B(n560), .Z(n454) );
  NAND U1585 ( .A(n455), .B(n454), .Z(n458) );
  NANDN U1586 ( .A(n458), .B(n459), .Z(n461) );
  XOR U1587 ( .A(n459), .B(n458), .Z(n567) );
  ANDN U1588 ( .B(b[60]), .A(n173), .Z(n566) );
  OR U1589 ( .A(n567), .B(n566), .Z(n460) );
  NAND U1590 ( .A(n461), .B(n460), .Z(n465) );
  XOR U1591 ( .A(n463), .B(n462), .Z(n464) );
  OR U1592 ( .A(n465), .B(n464), .Z(n467) );
  XNOR U1593 ( .A(n465), .B(n464), .Z(n573) );
  AND U1594 ( .A(a[17]), .B(b[60]), .Z(n572) );
  NANDN U1595 ( .A(n573), .B(n572), .Z(n466) );
  NAND U1596 ( .A(n467), .B(n466), .Z(n468) );
  OR U1597 ( .A(n469), .B(n468), .Z(n471) );
  XNOR U1598 ( .A(n469), .B(n468), .Z(n472) );
  ANDN U1599 ( .B(b[60]), .A(n175), .Z(n473) );
  OR U1600 ( .A(n472), .B(n473), .Z(n470) );
  AND U1601 ( .A(n471), .B(n470), .Z(n715) );
  XOR U1602 ( .A(n714), .B(n715), .Z(n716) );
  XNOR U1603 ( .A(n473), .B(n472), .Z(n579) );
  NAND U1604 ( .A(a[18]), .B(b[59]), .Z(n574) );
  XNOR U1605 ( .A(n475), .B(n474), .Z(n551) );
  XOR U1606 ( .A(n477), .B(n476), .Z(n528) );
  NAND U1607 ( .A(a[9]), .B(b[59]), .Z(n525) );
  XOR U1608 ( .A(n479), .B(n478), .Z(n524) );
  OR U1609 ( .A(n525), .B(n524), .Z(n527) );
  XOR U1610 ( .A(n481), .B(n480), .Z(n521) );
  NAND U1611 ( .A(a[6]), .B(b[59]), .Z(n485) );
  XNOR U1612 ( .A(n483), .B(n482), .Z(n484) );
  NANDN U1613 ( .A(n485), .B(n484), .Z(n513) );
  XOR U1614 ( .A(n485), .B(n484), .Z(n597) );
  NAND U1615 ( .A(a[5]), .B(b[59]), .Z(n509) );
  XOR U1616 ( .A(n487), .B(n486), .Z(n508) );
  NANDN U1617 ( .A(n509), .B(n508), .Z(n511) );
  XNOR U1618 ( .A(n489), .B(n488), .Z(n504) );
  XNOR U1619 ( .A(n491), .B(n490), .Z(n500) );
  NAND U1620 ( .A(b[60]), .B(a[1]), .Z(n493) );
  NAND U1621 ( .A(n493), .B(n492), .Z(n496) );
  OR U1622 ( .A(n493), .B(n742), .Z(n607) );
  NANDN U1623 ( .A(n495), .B(n607), .Z(n494) );
  AND U1624 ( .A(n496), .B(n494), .Z(n499) );
  XNOR U1625 ( .A(n607), .B(n495), .Z(n497) );
  NAND U1626 ( .A(n497), .B(n496), .Z(n603) );
  ANDN U1627 ( .B(b[59]), .A(n162), .Z(n602) );
  OR U1628 ( .A(n603), .B(n602), .Z(n498) );
  AND U1629 ( .A(n499), .B(n498), .Z(n501) );
  OR U1630 ( .A(n500), .B(n501), .Z(n503) );
  XNOR U1631 ( .A(n501), .B(n500), .Z(n600) );
  ANDN U1632 ( .B(b[59]), .A(n21580), .Z(n601) );
  OR U1633 ( .A(n600), .B(n601), .Z(n502) );
  AND U1634 ( .A(n503), .B(n502), .Z(n505) );
  OR U1635 ( .A(n504), .B(n505), .Z(n507) );
  XNOR U1636 ( .A(n505), .B(n504), .Z(n598) );
  ANDN U1637 ( .B(b[59]), .A(n163), .Z(n599) );
  OR U1638 ( .A(n598), .B(n599), .Z(n506) );
  NAND U1639 ( .A(n507), .B(n506), .Z(n625) );
  NANDN U1640 ( .A(n625), .B(n624), .Z(n510) );
  NAND U1641 ( .A(n511), .B(n510), .Z(n596) );
  NANDN U1642 ( .A(n597), .B(n596), .Z(n512) );
  NAND U1643 ( .A(n513), .B(n512), .Z(n516) );
  XOR U1644 ( .A(n515), .B(n514), .Z(n517) );
  NANDN U1645 ( .A(n516), .B(n517), .Z(n519) );
  ANDN U1646 ( .B(b[59]), .A(n166), .Z(n635) );
  XOR U1647 ( .A(n517), .B(n516), .Z(n634) );
  OR U1648 ( .A(n635), .B(n634), .Z(n518) );
  AND U1649 ( .A(n519), .B(n518), .Z(n520) );
  NANDN U1650 ( .A(n521), .B(n520), .Z(n523) );
  NAND U1651 ( .A(a[8]), .B(b[59]), .Z(n595) );
  NANDN U1652 ( .A(n595), .B(n594), .Z(n522) );
  AND U1653 ( .A(n523), .B(n522), .Z(n644) );
  XNOR U1654 ( .A(n525), .B(n524), .Z(n645) );
  OR U1655 ( .A(n644), .B(n645), .Z(n526) );
  AND U1656 ( .A(n527), .B(n526), .Z(n529) );
  OR U1657 ( .A(n528), .B(n529), .Z(n531) );
  XNOR U1658 ( .A(n529), .B(n528), .Z(n651) );
  AND U1659 ( .A(a[10]), .B(b[59]), .Z(n650) );
  NANDN U1660 ( .A(n651), .B(n650), .Z(n530) );
  NAND U1661 ( .A(n531), .B(n530), .Z(n535) );
  OR U1662 ( .A(n535), .B(n534), .Z(n537) );
  XOR U1663 ( .A(n535), .B(n534), .Z(n592) );
  NAND U1664 ( .A(b[59]), .B(a[11]), .Z(n593) );
  NAND U1665 ( .A(n592), .B(n593), .Z(n536) );
  NAND U1666 ( .A(n537), .B(n536), .Z(n540) );
  NANDN U1667 ( .A(n540), .B(n541), .Z(n543) );
  NAND U1668 ( .A(a[12]), .B(b[59]), .Z(n661) );
  XNOR U1669 ( .A(n541), .B(n540), .Z(n660) );
  NANDN U1670 ( .A(n661), .B(n660), .Z(n542) );
  NAND U1671 ( .A(n543), .B(n542), .Z(n546) );
  OR U1672 ( .A(n546), .B(n547), .Z(n549) );
  ANDN U1673 ( .B(b[59]), .A(n170), .Z(n590) );
  XOR U1674 ( .A(n547), .B(n546), .Z(n591) );
  NANDN U1675 ( .A(n590), .B(n591), .Z(n548) );
  AND U1676 ( .A(n549), .B(n548), .Z(n550) );
  OR U1677 ( .A(n551), .B(n550), .Z(n553) );
  XNOR U1678 ( .A(n551), .B(n550), .Z(n588) );
  ANDN U1679 ( .B(b[59]), .A(n171), .Z(n589) );
  OR U1680 ( .A(n588), .B(n589), .Z(n552) );
  NAND U1681 ( .A(n553), .B(n552), .Z(n557) );
  XOR U1682 ( .A(n555), .B(n554), .Z(n556) );
  NANDN U1683 ( .A(n557), .B(n556), .Z(n559) );
  NAND U1684 ( .A(a[15]), .B(b[59]), .Z(n675) );
  NANDN U1685 ( .A(n675), .B(n674), .Z(n558) );
  NAND U1686 ( .A(n559), .B(n558), .Z(n562) );
  XOR U1687 ( .A(n561), .B(n560), .Z(n563) );
  OR U1688 ( .A(n562), .B(n563), .Z(n565) );
  ANDN U1689 ( .B(b[59]), .A(n173), .Z(n586) );
  XOR U1690 ( .A(n563), .B(n562), .Z(n587) );
  NANDN U1691 ( .A(n586), .B(n587), .Z(n564) );
  NAND U1692 ( .A(n565), .B(n564), .Z(n568) );
  XOR U1693 ( .A(n567), .B(n566), .Z(n569) );
  OR U1694 ( .A(n568), .B(n569), .Z(n571) );
  NAND U1695 ( .A(a[17]), .B(b[59]), .Z(n685) );
  XOR U1696 ( .A(n569), .B(n568), .Z(n684) );
  NANDN U1697 ( .A(n685), .B(n684), .Z(n570) );
  AND U1698 ( .A(n571), .B(n570), .Z(n575) );
  OR U1699 ( .A(n574), .B(n575), .Z(n577) );
  XOR U1700 ( .A(n573), .B(n572), .Z(n585) );
  XNOR U1701 ( .A(n575), .B(n574), .Z(n584) );
  OR U1702 ( .A(n585), .B(n584), .Z(n576) );
  NAND U1703 ( .A(n577), .B(n576), .Z(n578) );
  OR U1704 ( .A(n579), .B(n578), .Z(n581) );
  XNOR U1705 ( .A(n579), .B(n578), .Z(n583) );
  ANDN U1706 ( .B(b[59]), .A(n21670), .Z(n582) );
  OR U1707 ( .A(n583), .B(n582), .Z(n580) );
  AND U1708 ( .A(n581), .B(n580), .Z(n721) );
  XOR U1709 ( .A(n720), .B(n721), .Z(n723) );
  XNOR U1710 ( .A(n722), .B(n723), .Z(n699) );
  NAND U1711 ( .A(a[20]), .B(b[58]), .Z(n694) );
  XOR U1712 ( .A(n583), .B(n582), .Z(n695) );
  OR U1713 ( .A(n694), .B(n695), .Z(n697) );
  XOR U1714 ( .A(n585), .B(n584), .Z(n690) );
  XOR U1715 ( .A(n587), .B(n586), .Z(n680) );
  XNOR U1716 ( .A(n589), .B(n588), .Z(n670) );
  XOR U1717 ( .A(n591), .B(n590), .Z(n666) );
  NAND U1718 ( .A(a[12]), .B(b[58]), .Z(n657) );
  NANDN U1719 ( .A(n657), .B(n656), .Z(n659) );
  XNOR U1720 ( .A(n595), .B(n594), .Z(n641) );
  XOR U1721 ( .A(n597), .B(n596), .Z(n631) );
  NAND U1722 ( .A(b[58]), .B(a[7]), .Z(n630) );
  OR U1723 ( .A(n631), .B(n630), .Z(n633) );
  XNOR U1724 ( .A(n599), .B(n598), .Z(n620) );
  XNOR U1725 ( .A(n601), .B(n600), .Z(n616) );
  XNOR U1726 ( .A(n603), .B(n602), .Z(n612) );
  NAND U1727 ( .A(b[59]), .B(a[1]), .Z(n605) );
  NAND U1728 ( .A(n605), .B(n604), .Z(n608) );
  OR U1729 ( .A(n605), .B(n994), .Z(n745) );
  NANDN U1730 ( .A(n607), .B(n745), .Z(n606) );
  AND U1731 ( .A(n608), .B(n606), .Z(n611) );
  XNOR U1732 ( .A(n745), .B(n607), .Z(n609) );
  NAND U1733 ( .A(n609), .B(n608), .Z(n741) );
  ANDN U1734 ( .B(b[58]), .A(n162), .Z(n740) );
  OR U1735 ( .A(n741), .B(n740), .Z(n610) );
  AND U1736 ( .A(n611), .B(n610), .Z(n613) );
  OR U1737 ( .A(n612), .B(n613), .Z(n615) );
  XNOR U1738 ( .A(n613), .B(n612), .Z(n738) );
  ANDN U1739 ( .B(b[58]), .A(n21580), .Z(n739) );
  OR U1740 ( .A(n738), .B(n739), .Z(n614) );
  AND U1741 ( .A(n615), .B(n614), .Z(n617) );
  OR U1742 ( .A(n616), .B(n617), .Z(n619) );
  XNOR U1743 ( .A(n617), .B(n616), .Z(n736) );
  ANDN U1744 ( .B(b[58]), .A(n163), .Z(n737) );
  OR U1745 ( .A(n736), .B(n737), .Z(n618) );
  AND U1746 ( .A(n619), .B(n618), .Z(n621) );
  OR U1747 ( .A(n620), .B(n621), .Z(n623) );
  XNOR U1748 ( .A(n621), .B(n620), .Z(n764) );
  NAND U1749 ( .A(b[58]), .B(a[5]), .Z(n765) );
  NANDN U1750 ( .A(n764), .B(n765), .Z(n622) );
  NAND U1751 ( .A(n623), .B(n622), .Z(n627) );
  NANDN U1752 ( .A(n627), .B(n626), .Z(n629) );
  NAND U1753 ( .A(a[6]), .B(b[58]), .Z(n769) );
  NANDN U1754 ( .A(n769), .B(n768), .Z(n628) );
  AND U1755 ( .A(n629), .B(n628), .Z(n774) );
  XOR U1756 ( .A(n631), .B(n630), .Z(n775) );
  NANDN U1757 ( .A(n774), .B(n775), .Z(n632) );
  NAND U1758 ( .A(n633), .B(n632), .Z(n637) );
  XOR U1759 ( .A(n635), .B(n634), .Z(n636) );
  NANDN U1760 ( .A(n637), .B(n636), .Z(n639) );
  ANDN U1761 ( .B(b[58]), .A(n167), .Z(n781) );
  XOR U1762 ( .A(n637), .B(n636), .Z(n780) );
  OR U1763 ( .A(n781), .B(n780), .Z(n638) );
  NAND U1764 ( .A(n639), .B(n638), .Z(n640) );
  NANDN U1765 ( .A(n641), .B(n640), .Z(n643) );
  ANDN U1766 ( .B(b[58]), .A(n21615), .Z(n735) );
  NANDN U1767 ( .A(n735), .B(n734), .Z(n642) );
  NAND U1768 ( .A(n643), .B(n642), .Z(n647) );
  XOR U1769 ( .A(n645), .B(n644), .Z(n646) );
  NANDN U1770 ( .A(n647), .B(n646), .Z(n649) );
  NAND U1771 ( .A(a[10]), .B(b[58]), .Z(n790) );
  XNOR U1772 ( .A(n647), .B(n646), .Z(n791) );
  NANDN U1773 ( .A(n790), .B(n791), .Z(n648) );
  AND U1774 ( .A(n649), .B(n648), .Z(n652) );
  XOR U1775 ( .A(n651), .B(n650), .Z(n653) );
  OR U1776 ( .A(n652), .B(n653), .Z(n655) );
  NAND U1777 ( .A(a[11]), .B(b[58]), .Z(n797) );
  XOR U1778 ( .A(n653), .B(n652), .Z(n796) );
  NANDN U1779 ( .A(n797), .B(n796), .Z(n654) );
  AND U1780 ( .A(n655), .B(n654), .Z(n733) );
  NANDN U1781 ( .A(n733), .B(n732), .Z(n658) );
  NAND U1782 ( .A(n659), .B(n658), .Z(n662) );
  OR U1783 ( .A(n662), .B(n663), .Z(n665) );
  ANDN U1784 ( .B(b[58]), .A(n170), .Z(n807) );
  XOR U1785 ( .A(n663), .B(n662), .Z(n806) );
  NANDN U1786 ( .A(n807), .B(n806), .Z(n664) );
  AND U1787 ( .A(n665), .B(n664), .Z(n667) );
  OR U1788 ( .A(n666), .B(n667), .Z(n669) );
  XNOR U1789 ( .A(n667), .B(n666), .Z(n812) );
  NAND U1790 ( .A(b[58]), .B(a[14]), .Z(n813) );
  NANDN U1791 ( .A(n812), .B(n813), .Z(n668) );
  AND U1792 ( .A(n669), .B(n668), .Z(n671) );
  OR U1793 ( .A(n670), .B(n671), .Z(n673) );
  XNOR U1794 ( .A(n671), .B(n670), .Z(n818) );
  ANDN U1795 ( .B(b[58]), .A(n172), .Z(n819) );
  OR U1796 ( .A(n818), .B(n819), .Z(n672) );
  AND U1797 ( .A(n673), .B(n672), .Z(n676) );
  OR U1798 ( .A(n676), .B(n677), .Z(n679) );
  XOR U1799 ( .A(n677), .B(n676), .Z(n824) );
  NAND U1800 ( .A(b[58]), .B(a[16]), .Z(n825) );
  NAND U1801 ( .A(n824), .B(n825), .Z(n678) );
  AND U1802 ( .A(n679), .B(n678), .Z(n681) );
  OR U1803 ( .A(n680), .B(n681), .Z(n683) );
  XNOR U1804 ( .A(n681), .B(n680), .Z(n830) );
  NAND U1805 ( .A(b[58]), .B(a[17]), .Z(n831) );
  NANDN U1806 ( .A(n830), .B(n831), .Z(n682) );
  AND U1807 ( .A(n683), .B(n682), .Z(n686) );
  OR U1808 ( .A(n686), .B(n687), .Z(n689) );
  XOR U1809 ( .A(n687), .B(n686), .Z(n838) );
  NAND U1810 ( .A(b[58]), .B(a[18]), .Z(n839) );
  NAND U1811 ( .A(n838), .B(n839), .Z(n688) );
  AND U1812 ( .A(n689), .B(n688), .Z(n691) );
  OR U1813 ( .A(n690), .B(n691), .Z(n693) );
  XNOR U1814 ( .A(n691), .B(n690), .Z(n731) );
  ANDN U1815 ( .B(b[58]), .A(n21670), .Z(n730) );
  OR U1816 ( .A(n731), .B(n730), .Z(n692) );
  NAND U1817 ( .A(n693), .B(n692), .Z(n728) );
  XOR U1818 ( .A(n695), .B(n694), .Z(n729) );
  NANDN U1819 ( .A(n728), .B(n729), .Z(n696) );
  NAND U1820 ( .A(n697), .B(n696), .Z(n698) );
  OR U1821 ( .A(n699), .B(n698), .Z(n701) );
  XNOR U1822 ( .A(n699), .B(n698), .Z(n727) );
  IV U1823 ( .A(a[21]), .Z(n21681) );
  ANDN U1824 ( .B(b[58]), .A(n21681), .Z(n726) );
  OR U1825 ( .A(n727), .B(n726), .Z(n700) );
  AND U1826 ( .A(n701), .B(n700), .Z(n858) );
  NAND U1827 ( .A(b[61]), .B(a[19]), .Z(n866) );
  OR U1828 ( .A(n703), .B(n702), .Z(n707) );
  OR U1829 ( .A(n705), .B(n704), .Z(n706) );
  AND U1830 ( .A(n707), .B(n706), .Z(n864) );
  ANDN U1831 ( .B(b[63]), .A(n174), .Z(n872) );
  ANDN U1832 ( .B(a[18]), .A(n159), .Z(n870) );
  OR U1833 ( .A(n709), .B(n708), .Z(n713) );
  OR U1834 ( .A(n711), .B(n710), .Z(n712) );
  AND U1835 ( .A(n713), .B(n712), .Z(n871) );
  XNOR U1836 ( .A(n870), .B(n871), .Z(n873) );
  XNOR U1837 ( .A(n872), .B(n873), .Z(n865) );
  XNOR U1838 ( .A(n864), .B(n865), .Z(n867) );
  XOR U1839 ( .A(n866), .B(n867), .Z(n878) );
  NAND U1840 ( .A(a[20]), .B(b[60]), .Z(n877) );
  OR U1841 ( .A(n715), .B(n714), .Z(n719) );
  NANDN U1842 ( .A(n717), .B(n716), .Z(n718) );
  NAND U1843 ( .A(n719), .B(n718), .Z(n876) );
  XNOR U1844 ( .A(n877), .B(n876), .Z(n879) );
  XNOR U1845 ( .A(n878), .B(n879), .Z(n882) );
  NANDN U1846 ( .A(n721), .B(n720), .Z(n725) );
  OR U1847 ( .A(n723), .B(n722), .Z(n724) );
  AND U1848 ( .A(n725), .B(n724), .Z(n883) );
  XNOR U1849 ( .A(n882), .B(n883), .Z(n885) );
  ANDN U1850 ( .B(b[59]), .A(n21681), .Z(n884) );
  XNOR U1851 ( .A(n885), .B(n884), .Z(n859) );
  XNOR U1852 ( .A(n858), .B(n859), .Z(n861) );
  XNOR U1853 ( .A(n860), .B(n861), .Z(n855) );
  XNOR U1854 ( .A(n727), .B(n726), .Z(n851) );
  XNOR U1855 ( .A(n729), .B(n728), .Z(n846) );
  XNOR U1856 ( .A(n731), .B(n730), .Z(n843) );
  NAND U1857 ( .A(a[19]), .B(b[57]), .Z(n836) );
  XOR U1858 ( .A(n733), .B(n732), .Z(n803) );
  NAND U1859 ( .A(b[57]), .B(a[13]), .Z(n802) );
  OR U1860 ( .A(n803), .B(n802), .Z(n805) );
  ANDN U1861 ( .B(b[57]), .A(n168), .Z(n786) );
  XOR U1862 ( .A(n735), .B(n734), .Z(n787) );
  OR U1863 ( .A(n786), .B(n787), .Z(n789) );
  XNOR U1864 ( .A(n737), .B(n736), .Z(n759) );
  XNOR U1865 ( .A(n739), .B(n738), .Z(n754) );
  XNOR U1866 ( .A(n741), .B(n740), .Z(n750) );
  NAND U1867 ( .A(b[58]), .B(a[1]), .Z(n743) );
  NAND U1868 ( .A(n743), .B(n742), .Z(n746) );
  OR U1869 ( .A(n743), .B(n1148), .Z(n997) );
  NANDN U1870 ( .A(n745), .B(n997), .Z(n744) );
  AND U1871 ( .A(n746), .B(n744), .Z(n749) );
  XNOR U1872 ( .A(n997), .B(n745), .Z(n747) );
  NAND U1873 ( .A(n747), .B(n746), .Z(n993) );
  ANDN U1874 ( .B(b[57]), .A(n162), .Z(n992) );
  OR U1875 ( .A(n993), .B(n992), .Z(n748) );
  AND U1876 ( .A(n749), .B(n748), .Z(n751) );
  OR U1877 ( .A(n750), .B(n751), .Z(n753) );
  XNOR U1878 ( .A(n751), .B(n750), .Z(n990) );
  ANDN U1879 ( .B(b[57]), .A(n21580), .Z(n991) );
  OR U1880 ( .A(n990), .B(n991), .Z(n752) );
  AND U1881 ( .A(n753), .B(n752), .Z(n755) );
  OR U1882 ( .A(n754), .B(n755), .Z(n757) );
  XNOR U1883 ( .A(n755), .B(n754), .Z(n988) );
  ANDN U1884 ( .B(b[57]), .A(n163), .Z(n989) );
  OR U1885 ( .A(n988), .B(n989), .Z(n756) );
  AND U1886 ( .A(n757), .B(n756), .Z(n758) );
  OR U1887 ( .A(n759), .B(n758), .Z(n761) );
  XNOR U1888 ( .A(n759), .B(n758), .Z(n1016) );
  NAND U1889 ( .A(b[57]), .B(a[5]), .Z(n1017) );
  NANDN U1890 ( .A(n1016), .B(n1017), .Z(n760) );
  NAND U1891 ( .A(n761), .B(n760), .Z(n763) );
  AND U1892 ( .A(a[6]), .B(b[57]), .Z(n762) );
  NANDN U1893 ( .A(n763), .B(n762), .Z(n767) );
  XOR U1894 ( .A(n763), .B(n762), .Z(n984) );
  XOR U1895 ( .A(n765), .B(n764), .Z(n985) );
  NANDN U1896 ( .A(n984), .B(n985), .Z(n766) );
  AND U1897 ( .A(n767), .B(n766), .Z(n770) );
  NANDN U1898 ( .A(n770), .B(n771), .Z(n773) );
  XOR U1899 ( .A(n771), .B(n770), .Z(n1023) );
  AND U1900 ( .A(a[7]), .B(b[57]), .Z(n1022) );
  NANDN U1901 ( .A(n1023), .B(n1022), .Z(n772) );
  NAND U1902 ( .A(n773), .B(n772), .Z(n777) );
  XOR U1903 ( .A(n775), .B(n774), .Z(n776) );
  NANDN U1904 ( .A(n777), .B(n776), .Z(n779) );
  ANDN U1905 ( .B(b[57]), .A(n167), .Z(n1029) );
  OR U1906 ( .A(n1029), .B(n1028), .Z(n778) );
  NAND U1907 ( .A(n779), .B(n778), .Z(n782) );
  XNOR U1908 ( .A(n781), .B(n780), .Z(n783) );
  NANDN U1909 ( .A(n782), .B(n783), .Z(n785) );
  XOR U1910 ( .A(n783), .B(n782), .Z(n982) );
  NAND U1911 ( .A(a[9]), .B(b[57]), .Z(n983) );
  OR U1912 ( .A(n982), .B(n983), .Z(n784) );
  AND U1913 ( .A(n785), .B(n784), .Z(n980) );
  XOR U1914 ( .A(n787), .B(n786), .Z(n981) );
  NAND U1915 ( .A(n980), .B(n981), .Z(n788) );
  AND U1916 ( .A(n789), .B(n788), .Z(n793) );
  XOR U1917 ( .A(n791), .B(n790), .Z(n792) );
  NANDN U1918 ( .A(n793), .B(n792), .Z(n795) );
  ANDN U1919 ( .B(b[57]), .A(n21164), .Z(n977) );
  NANDN U1920 ( .A(n977), .B(n976), .Z(n794) );
  NAND U1921 ( .A(n795), .B(n794), .Z(n799) );
  XNOR U1922 ( .A(n797), .B(n796), .Z(n798) );
  NANDN U1923 ( .A(n799), .B(n798), .Z(n801) );
  NAND U1924 ( .A(a[12]), .B(b[57]), .Z(n975) );
  XNOR U1925 ( .A(n799), .B(n798), .Z(n974) );
  NANDN U1926 ( .A(n975), .B(n974), .Z(n800) );
  AND U1927 ( .A(n801), .B(n800), .Z(n1048) );
  XOR U1928 ( .A(n803), .B(n802), .Z(n1049) );
  NANDN U1929 ( .A(n1048), .B(n1049), .Z(n804) );
  NAND U1930 ( .A(n805), .B(n804), .Z(n809) );
  XOR U1931 ( .A(n807), .B(n806), .Z(n808) );
  OR U1932 ( .A(n809), .B(n808), .Z(n811) );
  ANDN U1933 ( .B(b[57]), .A(n171), .Z(n971) );
  XOR U1934 ( .A(n809), .B(n808), .Z(n970) );
  NANDN U1935 ( .A(n971), .B(n970), .Z(n810) );
  NAND U1936 ( .A(n811), .B(n810), .Z(n815) );
  XOR U1937 ( .A(n813), .B(n812), .Z(n814) );
  NANDN U1938 ( .A(n815), .B(n814), .Z(n817) );
  NAND U1939 ( .A(a[15]), .B(b[57]), .Z(n1056) );
  XNOR U1940 ( .A(n815), .B(n814), .Z(n1057) );
  NANDN U1941 ( .A(n1056), .B(n1057), .Z(n816) );
  NAND U1942 ( .A(n817), .B(n816), .Z(n821) );
  XOR U1943 ( .A(n819), .B(n818), .Z(n820) );
  NANDN U1944 ( .A(n821), .B(n820), .Z(n823) );
  ANDN U1945 ( .B(b[57]), .A(n173), .Z(n969) );
  NANDN U1946 ( .A(n969), .B(n968), .Z(n822) );
  NAND U1947 ( .A(n823), .B(n822), .Z(n827) );
  NANDN U1948 ( .A(n827), .B(n826), .Z(n829) );
  NAND U1949 ( .A(a[17]), .B(b[57]), .Z(n966) );
  NANDN U1950 ( .A(n966), .B(n967), .Z(n828) );
  AND U1951 ( .A(n829), .B(n828), .Z(n833) );
  XOR U1952 ( .A(n831), .B(n830), .Z(n832) );
  NANDN U1953 ( .A(n833), .B(n832), .Z(n835) );
  NAND U1954 ( .A(a[18]), .B(b[57]), .Z(n965) );
  NANDN U1955 ( .A(n965), .B(n964), .Z(n834) );
  AND U1956 ( .A(n835), .B(n834), .Z(n837) );
  OR U1957 ( .A(n836), .B(n837), .Z(n841) );
  XNOR U1958 ( .A(n837), .B(n836), .Z(n1075) );
  NANDN U1959 ( .A(n1075), .B(n1074), .Z(n840) );
  NAND U1960 ( .A(n841), .B(n840), .Z(n842) );
  OR U1961 ( .A(n843), .B(n842), .Z(n845) );
  XNOR U1962 ( .A(n843), .B(n842), .Z(n1081) );
  ANDN U1963 ( .B(b[57]), .A(n176), .Z(n1080) );
  OR U1964 ( .A(n1081), .B(n1080), .Z(n844) );
  AND U1965 ( .A(n845), .B(n844), .Z(n847) );
  OR U1966 ( .A(n846), .B(n847), .Z(n849) );
  XNOR U1967 ( .A(n847), .B(n846), .Z(n962) );
  ANDN U1968 ( .B(b[57]), .A(n21681), .Z(n963) );
  OR U1969 ( .A(n962), .B(n963), .Z(n848) );
  AND U1970 ( .A(n849), .B(n848), .Z(n850) );
  OR U1971 ( .A(n851), .B(n850), .Z(n853) );
  XNOR U1972 ( .A(n851), .B(n850), .Z(n960) );
  ANDN U1973 ( .B(b[57]), .A(n177), .Z(n961) );
  OR U1974 ( .A(n960), .B(n961), .Z(n852) );
  AND U1975 ( .A(n853), .B(n852), .Z(n854) );
  OR U1976 ( .A(n855), .B(n854), .Z(n857) );
  XNOR U1977 ( .A(n855), .B(n854), .Z(n958) );
  IV U1978 ( .A(a[23]), .Z(n21692) );
  ANDN U1979 ( .B(b[57]), .A(n21692), .Z(n959) );
  OR U1980 ( .A(n958), .B(n959), .Z(n856) );
  AND U1981 ( .A(n857), .B(n856), .Z(n888) );
  ANDN U1982 ( .B(b[58]), .A(n21692), .Z(n892) );
  OR U1983 ( .A(n859), .B(n858), .Z(n863) );
  OR U1984 ( .A(n861), .B(n860), .Z(n862) );
  AND U1985 ( .A(n863), .B(n862), .Z(n893) );
  XNOR U1986 ( .A(n892), .B(n893), .Z(n895) );
  NAND U1987 ( .A(b[61]), .B(a[20]), .Z(n906) );
  OR U1988 ( .A(n865), .B(n864), .Z(n869) );
  NANDN U1989 ( .A(n867), .B(n866), .Z(n868) );
  AND U1990 ( .A(n869), .B(n868), .Z(n904) );
  ANDN U1991 ( .B(b[63]), .A(n175), .Z(n912) );
  ANDN U1992 ( .B(a[19]), .A(n159), .Z(n910) );
  OR U1993 ( .A(n871), .B(n870), .Z(n875) );
  OR U1994 ( .A(n873), .B(n872), .Z(n874) );
  AND U1995 ( .A(n875), .B(n874), .Z(n911) );
  XNOR U1996 ( .A(n910), .B(n911), .Z(n913) );
  XNOR U1997 ( .A(n912), .B(n913), .Z(n905) );
  XNOR U1998 ( .A(n904), .B(n905), .Z(n907) );
  XOR U1999 ( .A(n906), .B(n907), .Z(n918) );
  NAND U2000 ( .A(a[21]), .B(b[60]), .Z(n917) );
  OR U2001 ( .A(n877), .B(n876), .Z(n881) );
  NANDN U2002 ( .A(n879), .B(n878), .Z(n880) );
  AND U2003 ( .A(n881), .B(n880), .Z(n916) );
  XNOR U2004 ( .A(n917), .B(n916), .Z(n919) );
  XNOR U2005 ( .A(n918), .B(n919), .Z(n898) );
  OR U2006 ( .A(n883), .B(n882), .Z(n887) );
  OR U2007 ( .A(n885), .B(n884), .Z(n886) );
  AND U2008 ( .A(n887), .B(n886), .Z(n899) );
  XNOR U2009 ( .A(n898), .B(n899), .Z(n901) );
  ANDN U2010 ( .B(b[59]), .A(n177), .Z(n900) );
  XOR U2011 ( .A(n901), .B(n900), .Z(n894) );
  NANDN U2012 ( .A(n888), .B(n889), .Z(n891) );
  XOR U2013 ( .A(n889), .B(n888), .Z(n956) );
  ANDN U2014 ( .B(b[57]), .A(n178), .Z(n957) );
  OR U2015 ( .A(n956), .B(n957), .Z(n890) );
  NAND U2016 ( .A(n891), .B(n890), .Z(n923) );
  ANDN U2017 ( .B(b[58]), .A(n178), .Z(n926) );
  OR U2018 ( .A(n893), .B(n892), .Z(n897) );
  NANDN U2019 ( .A(n895), .B(n894), .Z(n896) );
  AND U2020 ( .A(n897), .B(n896), .Z(n927) );
  XNOR U2021 ( .A(n926), .B(n927), .Z(n929) );
  OR U2022 ( .A(n899), .B(n898), .Z(n903) );
  OR U2023 ( .A(n901), .B(n900), .Z(n902) );
  AND U2024 ( .A(n903), .B(n902), .Z(n933) );
  ANDN U2025 ( .B(b[61]), .A(n21681), .Z(n940) );
  OR U2026 ( .A(n905), .B(n904), .Z(n909) );
  NANDN U2027 ( .A(n907), .B(n906), .Z(n908) );
  AND U2028 ( .A(n909), .B(n908), .Z(n938) );
  ANDN U2029 ( .B(b[63]), .A(n21670), .Z(n946) );
  ANDN U2030 ( .B(a[20]), .A(n159), .Z(n944) );
  OR U2031 ( .A(n911), .B(n910), .Z(n915) );
  OR U2032 ( .A(n913), .B(n912), .Z(n914) );
  AND U2033 ( .A(n915), .B(n914), .Z(n945) );
  XNOR U2034 ( .A(n944), .B(n945), .Z(n947) );
  XNOR U2035 ( .A(n946), .B(n947), .Z(n939) );
  XNOR U2036 ( .A(n938), .B(n939), .Z(n941) );
  XNOR U2037 ( .A(n940), .B(n941), .Z(n953) );
  ANDN U2038 ( .B(b[60]), .A(n177), .Z(n950) );
  OR U2039 ( .A(n917), .B(n916), .Z(n921) );
  NANDN U2040 ( .A(n919), .B(n918), .Z(n920) );
  NAND U2041 ( .A(n921), .B(n920), .Z(n951) );
  XOR U2042 ( .A(n950), .B(n951), .Z(n952) );
  XOR U2043 ( .A(n933), .B(n932), .Z(n935) );
  ANDN U2044 ( .B(b[59]), .A(n21692), .Z(n934) );
  XNOR U2045 ( .A(n935), .B(n934), .Z(n928) );
  XOR U2046 ( .A(n929), .B(n928), .Z(n922) );
  OR U2047 ( .A(n923), .B(n922), .Z(n925) );
  NAND U2048 ( .A(a[25]), .B(b[57]), .Z(n1103) );
  XOR U2049 ( .A(n923), .B(n922), .Z(n1102) );
  NANDN U2050 ( .A(n1103), .B(n1102), .Z(n924) );
  AND U2051 ( .A(n925), .B(n924), .Z(n1440) );
  IV U2052 ( .A(a[25]), .Z(n21703) );
  ANDN U2053 ( .B(b[58]), .A(n21703), .Z(n1470) );
  OR U2054 ( .A(n927), .B(n926), .Z(n931) );
  OR U2055 ( .A(n929), .B(n928), .Z(n930) );
  AND U2056 ( .A(n931), .B(n930), .Z(n1471) );
  XNOR U2057 ( .A(n1470), .B(n1471), .Z(n1473) );
  NANDN U2058 ( .A(n933), .B(n932), .Z(n937) );
  OR U2059 ( .A(n935), .B(n934), .Z(n936) );
  AND U2060 ( .A(n937), .B(n936), .Z(n1447) );
  ANDN U2061 ( .B(b[61]), .A(n177), .Z(n1454) );
  OR U2062 ( .A(n939), .B(n938), .Z(n943) );
  OR U2063 ( .A(n941), .B(n940), .Z(n942) );
  AND U2064 ( .A(n943), .B(n942), .Z(n1452) );
  ANDN U2065 ( .B(b[63]), .A(n176), .Z(n1460) );
  ANDN U2066 ( .B(a[21]), .A(n159), .Z(n1458) );
  OR U2067 ( .A(n945), .B(n944), .Z(n949) );
  OR U2068 ( .A(n947), .B(n946), .Z(n948) );
  AND U2069 ( .A(n949), .B(n948), .Z(n1459) );
  XNOR U2070 ( .A(n1458), .B(n1459), .Z(n1461) );
  XNOR U2071 ( .A(n1460), .B(n1461), .Z(n1453) );
  XNOR U2072 ( .A(n1452), .B(n1453), .Z(n1455) );
  XNOR U2073 ( .A(n1454), .B(n1455), .Z(n1467) );
  ANDN U2074 ( .B(b[60]), .A(n21692), .Z(n1464) );
  OR U2075 ( .A(n951), .B(n950), .Z(n955) );
  NANDN U2076 ( .A(n953), .B(n952), .Z(n954) );
  AND U2077 ( .A(n955), .B(n954), .Z(n1465) );
  XOR U2078 ( .A(n1464), .B(n1465), .Z(n1466) );
  XOR U2079 ( .A(n1447), .B(n1446), .Z(n1449) );
  ANDN U2080 ( .B(b[59]), .A(n178), .Z(n1448) );
  XNOR U2081 ( .A(n1449), .B(n1448), .Z(n1472) );
  XOR U2082 ( .A(n1473), .B(n1472), .Z(n1441) );
  XNOR U2083 ( .A(n1440), .B(n1441), .Z(n1442) );
  XOR U2084 ( .A(n1443), .B(n1442), .Z(n1478) );
  IV U2085 ( .A(a[27]), .Z(n21716) );
  ANDN U2086 ( .B(b[56]), .A(n21716), .Z(n1476) );
  XNOR U2087 ( .A(n957), .B(n956), .Z(n1098) );
  XNOR U2088 ( .A(n959), .B(n958), .Z(n1094) );
  XNOR U2089 ( .A(n961), .B(n960), .Z(n1090) );
  XNOR U2090 ( .A(n963), .B(n962), .Z(n1086) );
  XNOR U2091 ( .A(n965), .B(n964), .Z(n1071) );
  XNOR U2092 ( .A(n967), .B(n966), .Z(n1067) );
  XOR U2093 ( .A(n969), .B(n968), .Z(n1063) );
  NAND U2094 ( .A(a[15]), .B(b[56]), .Z(n972) );
  NANDN U2095 ( .A(n972), .B(n973), .Z(n1055) );
  XOR U2096 ( .A(n973), .B(n972), .Z(n1122) );
  XOR U2097 ( .A(n975), .B(n974), .Z(n1045) );
  NAND U2098 ( .A(a[12]), .B(b[56]), .Z(n978) );
  NANDN U2099 ( .A(n978), .B(n979), .Z(n1043) );
  XOR U2100 ( .A(n979), .B(n978), .Z(n1127) );
  XNOR U2101 ( .A(n981), .B(n980), .Z(n1039) );
  XOR U2102 ( .A(n983), .B(n982), .Z(n1035) );
  XOR U2103 ( .A(n985), .B(n984), .Z(n987) );
  AND U2104 ( .A(a[7]), .B(b[56]), .Z(n986) );
  NANDN U2105 ( .A(n987), .B(n986), .Z(n1021) );
  XOR U2106 ( .A(n987), .B(n986), .Z(n1136) );
  XNOR U2107 ( .A(n989), .B(n988), .Z(n1011) );
  XNOR U2108 ( .A(n991), .B(n990), .Z(n1006) );
  XNOR U2109 ( .A(n993), .B(n992), .Z(n1002) );
  NAND U2110 ( .A(b[57]), .B(a[1]), .Z(n995) );
  NAND U2111 ( .A(n995), .B(n994), .Z(n998) );
  OR U2112 ( .A(n995), .B(n1306), .Z(n1151) );
  NANDN U2113 ( .A(n997), .B(n1151), .Z(n996) );
  AND U2114 ( .A(n998), .B(n996), .Z(n1001) );
  XNOR U2115 ( .A(n1151), .B(n997), .Z(n999) );
  NAND U2116 ( .A(n999), .B(n998), .Z(n1147) );
  ANDN U2117 ( .B(b[56]), .A(n162), .Z(n1146) );
  OR U2118 ( .A(n1147), .B(n1146), .Z(n1000) );
  AND U2119 ( .A(n1001), .B(n1000), .Z(n1003) );
  OR U2120 ( .A(n1002), .B(n1003), .Z(n1005) );
  XNOR U2121 ( .A(n1003), .B(n1002), .Z(n1144) );
  ANDN U2122 ( .B(b[56]), .A(n21580), .Z(n1145) );
  OR U2123 ( .A(n1144), .B(n1145), .Z(n1004) );
  AND U2124 ( .A(n1005), .B(n1004), .Z(n1007) );
  OR U2125 ( .A(n1006), .B(n1007), .Z(n1009) );
  XNOR U2126 ( .A(n1007), .B(n1006), .Z(n1142) );
  ANDN U2127 ( .B(b[56]), .A(n163), .Z(n1143) );
  OR U2128 ( .A(n1142), .B(n1143), .Z(n1008) );
  AND U2129 ( .A(n1009), .B(n1008), .Z(n1010) );
  OR U2130 ( .A(n1011), .B(n1010), .Z(n1013) );
  XNOR U2131 ( .A(n1011), .B(n1010), .Z(n1170) );
  NAND U2132 ( .A(b[56]), .B(a[5]), .Z(n1171) );
  NANDN U2133 ( .A(n1170), .B(n1171), .Z(n1012) );
  NAND U2134 ( .A(n1013), .B(n1012), .Z(n1015) );
  AND U2135 ( .A(a[6]), .B(b[56]), .Z(n1014) );
  NANDN U2136 ( .A(n1015), .B(n1014), .Z(n1019) );
  XOR U2137 ( .A(n1015), .B(n1014), .Z(n1138) );
  XOR U2138 ( .A(n1017), .B(n1016), .Z(n1139) );
  NANDN U2139 ( .A(n1138), .B(n1139), .Z(n1018) );
  AND U2140 ( .A(n1019), .B(n1018), .Z(n1137) );
  OR U2141 ( .A(n1136), .B(n1137), .Z(n1020) );
  AND U2142 ( .A(n1021), .B(n1020), .Z(n1024) );
  XNOR U2143 ( .A(n1023), .B(n1022), .Z(n1025) );
  NANDN U2144 ( .A(n1024), .B(n1025), .Z(n1027) );
  XOR U2145 ( .A(n1025), .B(n1024), .Z(n1181) );
  NAND U2146 ( .A(a[8]), .B(b[56]), .Z(n1180) );
  OR U2147 ( .A(n1181), .B(n1180), .Z(n1026) );
  NAND U2148 ( .A(n1027), .B(n1026), .Z(n1031) );
  XOR U2149 ( .A(n1029), .B(n1028), .Z(n1030) );
  NANDN U2150 ( .A(n1031), .B(n1030), .Z(n1033) );
  ANDN U2151 ( .B(b[56]), .A(n21615), .Z(n1135) );
  XOR U2152 ( .A(n1031), .B(n1030), .Z(n1134) );
  OR U2153 ( .A(n1135), .B(n1134), .Z(n1032) );
  NAND U2154 ( .A(n1033), .B(n1032), .Z(n1034) );
  NANDN U2155 ( .A(n1035), .B(n1034), .Z(n1037) );
  ANDN U2156 ( .B(b[56]), .A(n168), .Z(n1133) );
  NANDN U2157 ( .A(n1133), .B(n1132), .Z(n1036) );
  NAND U2158 ( .A(n1037), .B(n1036), .Z(n1038) );
  NANDN U2159 ( .A(n1039), .B(n1038), .Z(n1041) );
  ANDN U2160 ( .B(b[56]), .A(n21164), .Z(n1131) );
  NANDN U2161 ( .A(n1131), .B(n1130), .Z(n1040) );
  NAND U2162 ( .A(n1041), .B(n1040), .Z(n1126) );
  OR U2163 ( .A(n1127), .B(n1126), .Z(n1042) );
  NAND U2164 ( .A(n1043), .B(n1042), .Z(n1044) );
  NANDN U2165 ( .A(n1045), .B(n1044), .Z(n1047) );
  NAND U2166 ( .A(a[13]), .B(b[56]), .Z(n1201) );
  XOR U2167 ( .A(n1045), .B(n1044), .Z(n1200) );
  OR U2168 ( .A(n1201), .B(n1200), .Z(n1046) );
  NAND U2169 ( .A(n1047), .B(n1046), .Z(n1051) );
  XOR U2170 ( .A(n1049), .B(n1048), .Z(n1050) );
  NANDN U2171 ( .A(n1051), .B(n1050), .Z(n1053) );
  ANDN U2172 ( .B(b[56]), .A(n171), .Z(n1125) );
  NANDN U2173 ( .A(n1125), .B(n1124), .Z(n1052) );
  NAND U2174 ( .A(n1053), .B(n1052), .Z(n1123) );
  OR U2175 ( .A(n1122), .B(n1123), .Z(n1054) );
  NAND U2176 ( .A(n1055), .B(n1054), .Z(n1059) );
  XOR U2177 ( .A(n1057), .B(n1056), .Z(n1058) );
  NANDN U2178 ( .A(n1059), .B(n1058), .Z(n1061) );
  ANDN U2179 ( .B(b[56]), .A(n173), .Z(n1121) );
  NANDN U2180 ( .A(n1121), .B(n1120), .Z(n1060) );
  NAND U2181 ( .A(n1061), .B(n1060), .Z(n1062) );
  NANDN U2182 ( .A(n1063), .B(n1062), .Z(n1065) );
  ANDN U2183 ( .B(b[56]), .A(n174), .Z(n1119) );
  NANDN U2184 ( .A(n1119), .B(n1118), .Z(n1064) );
  NAND U2185 ( .A(n1065), .B(n1064), .Z(n1066) );
  NANDN U2186 ( .A(n1067), .B(n1066), .Z(n1069) );
  ANDN U2187 ( .B(b[56]), .A(n175), .Z(n1223) );
  NANDN U2188 ( .A(n1223), .B(n1222), .Z(n1068) );
  NAND U2189 ( .A(n1069), .B(n1068), .Z(n1070) );
  NANDN U2190 ( .A(n1071), .B(n1070), .Z(n1073) );
  ANDN U2191 ( .B(b[56]), .A(n21670), .Z(n1116) );
  NANDN U2192 ( .A(n1116), .B(n1117), .Z(n1072) );
  NAND U2193 ( .A(n1073), .B(n1072), .Z(n1077) );
  NANDN U2194 ( .A(n1077), .B(n1076), .Z(n1079) );
  NAND U2195 ( .A(a[20]), .B(b[56]), .Z(n1232) );
  XNOR U2196 ( .A(n1077), .B(n1076), .Z(n1233) );
  NANDN U2197 ( .A(n1232), .B(n1233), .Z(n1078) );
  NAND U2198 ( .A(n1079), .B(n1078), .Z(n1083) );
  XOR U2199 ( .A(n1081), .B(n1080), .Z(n1082) );
  NANDN U2200 ( .A(n1083), .B(n1082), .Z(n1085) );
  ANDN U2201 ( .B(b[56]), .A(n21681), .Z(n1115) );
  XOR U2202 ( .A(n1083), .B(n1082), .Z(n1114) );
  OR U2203 ( .A(n1115), .B(n1114), .Z(n1084) );
  AND U2204 ( .A(n1085), .B(n1084), .Z(n1087) );
  OR U2205 ( .A(n1086), .B(n1087), .Z(n1089) );
  XNOR U2206 ( .A(n1087), .B(n1086), .Z(n1112) );
  NAND U2207 ( .A(b[56]), .B(a[22]), .Z(n1113) );
  NANDN U2208 ( .A(n1112), .B(n1113), .Z(n1088) );
  AND U2209 ( .A(n1089), .B(n1088), .Z(n1091) );
  OR U2210 ( .A(n1090), .B(n1091), .Z(n1093) );
  XNOR U2211 ( .A(n1091), .B(n1090), .Z(n1110) );
  ANDN U2212 ( .B(b[56]), .A(n21692), .Z(n1111) );
  OR U2213 ( .A(n1110), .B(n1111), .Z(n1092) );
  AND U2214 ( .A(n1093), .B(n1092), .Z(n1095) );
  OR U2215 ( .A(n1094), .B(n1095), .Z(n1097) );
  XNOR U2216 ( .A(n1095), .B(n1094), .Z(n1250) );
  NAND U2217 ( .A(b[56]), .B(a[24]), .Z(n1251) );
  NANDN U2218 ( .A(n1250), .B(n1251), .Z(n1096) );
  AND U2219 ( .A(n1097), .B(n1096), .Z(n1099) );
  OR U2220 ( .A(n1098), .B(n1099), .Z(n1101) );
  XNOR U2221 ( .A(n1099), .B(n1098), .Z(n1256) );
  ANDN U2222 ( .B(b[56]), .A(n21703), .Z(n1257) );
  OR U2223 ( .A(n1256), .B(n1257), .Z(n1100) );
  AND U2224 ( .A(n1101), .B(n1100), .Z(n1104) );
  OR U2225 ( .A(n1104), .B(n1105), .Z(n1107) );
  ANDN U2226 ( .B(b[56]), .A(n179), .Z(n1109) );
  XOR U2227 ( .A(n1105), .B(n1104), .Z(n1108) );
  NANDN U2228 ( .A(n1109), .B(n1108), .Z(n1106) );
  AND U2229 ( .A(n1107), .B(n1106), .Z(n1477) );
  XNOR U2230 ( .A(n1476), .B(n1477), .Z(n1479) );
  XOR U2231 ( .A(n1478), .B(n1479), .Z(n1434) );
  XOR U2232 ( .A(n1109), .B(n1108), .Z(n1263) );
  XNOR U2233 ( .A(n1111), .B(n1110), .Z(n1247) );
  NAND U2234 ( .A(a[23]), .B(b[55]), .Z(n1243) );
  XOR U2235 ( .A(n1113), .B(n1112), .Z(n1242) );
  NANDN U2236 ( .A(n1243), .B(n1242), .Z(n1245) );
  XNOR U2237 ( .A(n1115), .B(n1114), .Z(n1239) );
  XNOR U2238 ( .A(n1117), .B(n1116), .Z(n1229) );
  ANDN U2239 ( .B(b[55]), .A(n175), .Z(n1218) );
  XOR U2240 ( .A(n1119), .B(n1118), .Z(n1219) );
  OR U2241 ( .A(n1218), .B(n1219), .Z(n1221) );
  XOR U2242 ( .A(n1121), .B(n1120), .Z(n1215) );
  XOR U2243 ( .A(n1123), .B(n1122), .Z(n1211) );
  XOR U2244 ( .A(n1125), .B(n1124), .Z(n1207) );
  NAND U2245 ( .A(a[13]), .B(b[55]), .Z(n1129) );
  XOR U2246 ( .A(n1127), .B(n1126), .Z(n1128) );
  NANDN U2247 ( .A(n1129), .B(n1128), .Z(n1199) );
  XOR U2248 ( .A(n1129), .B(n1128), .Z(n1285) );
  XOR U2249 ( .A(n1131), .B(n1130), .Z(n1195) );
  XOR U2250 ( .A(n1133), .B(n1132), .Z(n1191) );
  XNOR U2251 ( .A(n1135), .B(n1134), .Z(n1187) );
  XNOR U2252 ( .A(n1137), .B(n1136), .Z(n1177) );
  XOR U2253 ( .A(n1139), .B(n1138), .Z(n1141) );
  AND U2254 ( .A(a[7]), .B(b[55]), .Z(n1140) );
  NANDN U2255 ( .A(n1141), .B(n1140), .Z(n1175) );
  XOR U2256 ( .A(n1141), .B(n1140), .Z(n1294) );
  XNOR U2257 ( .A(n1143), .B(n1142), .Z(n1165) );
  XNOR U2258 ( .A(n1145), .B(n1144), .Z(n1160) );
  XNOR U2259 ( .A(n1147), .B(n1146), .Z(n1156) );
  NAND U2260 ( .A(b[56]), .B(a[1]), .Z(n1149) );
  NAND U2261 ( .A(n1149), .B(n1148), .Z(n1152) );
  OR U2262 ( .A(n1149), .B(n1584), .Z(n1309) );
  NANDN U2263 ( .A(n1151), .B(n1309), .Z(n1150) );
  AND U2264 ( .A(n1152), .B(n1150), .Z(n1155) );
  XNOR U2265 ( .A(n1309), .B(n1151), .Z(n1153) );
  NAND U2266 ( .A(n1153), .B(n1152), .Z(n1305) );
  ANDN U2267 ( .B(b[55]), .A(n162), .Z(n1304) );
  OR U2268 ( .A(n1305), .B(n1304), .Z(n1154) );
  AND U2269 ( .A(n1155), .B(n1154), .Z(n1157) );
  OR U2270 ( .A(n1156), .B(n1157), .Z(n1159) );
  XNOR U2271 ( .A(n1157), .B(n1156), .Z(n1302) );
  ANDN U2272 ( .B(b[55]), .A(n21580), .Z(n1303) );
  OR U2273 ( .A(n1302), .B(n1303), .Z(n1158) );
  AND U2274 ( .A(n1159), .B(n1158), .Z(n1161) );
  OR U2275 ( .A(n1160), .B(n1161), .Z(n1163) );
  XNOR U2276 ( .A(n1161), .B(n1160), .Z(n1300) );
  ANDN U2277 ( .B(b[55]), .A(n163), .Z(n1301) );
  OR U2278 ( .A(n1300), .B(n1301), .Z(n1162) );
  AND U2279 ( .A(n1163), .B(n1162), .Z(n1164) );
  OR U2280 ( .A(n1165), .B(n1164), .Z(n1167) );
  XNOR U2281 ( .A(n1165), .B(n1164), .Z(n1328) );
  NAND U2282 ( .A(b[55]), .B(a[5]), .Z(n1329) );
  NANDN U2283 ( .A(n1328), .B(n1329), .Z(n1166) );
  NAND U2284 ( .A(n1167), .B(n1166), .Z(n1169) );
  AND U2285 ( .A(a[6]), .B(b[55]), .Z(n1168) );
  NANDN U2286 ( .A(n1169), .B(n1168), .Z(n1173) );
  XOR U2287 ( .A(n1169), .B(n1168), .Z(n1296) );
  XOR U2288 ( .A(n1171), .B(n1170), .Z(n1297) );
  NANDN U2289 ( .A(n1296), .B(n1297), .Z(n1172) );
  AND U2290 ( .A(n1173), .B(n1172), .Z(n1295) );
  OR U2291 ( .A(n1294), .B(n1295), .Z(n1174) );
  AND U2292 ( .A(n1175), .B(n1174), .Z(n1176) );
  OR U2293 ( .A(n1177), .B(n1176), .Z(n1179) );
  XNOR U2294 ( .A(n1177), .B(n1176), .Z(n1339) );
  NAND U2295 ( .A(a[8]), .B(b[55]), .Z(n1338) );
  OR U2296 ( .A(n1339), .B(n1338), .Z(n1178) );
  NAND U2297 ( .A(n1179), .B(n1178), .Z(n1182) );
  XOR U2298 ( .A(n1181), .B(n1180), .Z(n1183) );
  OR U2299 ( .A(n1182), .B(n1183), .Z(n1185) );
  ANDN U2300 ( .B(b[55]), .A(n21615), .Z(n1293) );
  XOR U2301 ( .A(n1183), .B(n1182), .Z(n1292) );
  NANDN U2302 ( .A(n1293), .B(n1292), .Z(n1184) );
  NAND U2303 ( .A(n1185), .B(n1184), .Z(n1186) );
  NANDN U2304 ( .A(n1187), .B(n1186), .Z(n1189) );
  ANDN U2305 ( .B(b[55]), .A(n168), .Z(n1291) );
  NANDN U2306 ( .A(n1291), .B(n1290), .Z(n1188) );
  NAND U2307 ( .A(n1189), .B(n1188), .Z(n1190) );
  NANDN U2308 ( .A(n1191), .B(n1190), .Z(n1193) );
  ANDN U2309 ( .B(b[55]), .A(n21164), .Z(n1289) );
  NANDN U2310 ( .A(n1289), .B(n1288), .Z(n1192) );
  NAND U2311 ( .A(n1193), .B(n1192), .Z(n1194) );
  NANDN U2312 ( .A(n1195), .B(n1194), .Z(n1197) );
  ANDN U2313 ( .B(b[55]), .A(n169), .Z(n1287) );
  NANDN U2314 ( .A(n1287), .B(n1286), .Z(n1196) );
  NAND U2315 ( .A(n1197), .B(n1196), .Z(n1284) );
  OR U2316 ( .A(n1285), .B(n1284), .Z(n1198) );
  NAND U2317 ( .A(n1199), .B(n1198), .Z(n1203) );
  XNOR U2318 ( .A(n1201), .B(n1200), .Z(n1202) );
  NANDN U2319 ( .A(n1203), .B(n1202), .Z(n1205) );
  ANDN U2320 ( .B(b[55]), .A(n171), .Z(n1283) );
  NANDN U2321 ( .A(n1283), .B(n1282), .Z(n1204) );
  NAND U2322 ( .A(n1205), .B(n1204), .Z(n1206) );
  NANDN U2323 ( .A(n1207), .B(n1206), .Z(n1209) );
  ANDN U2324 ( .B(b[55]), .A(n172), .Z(n1279) );
  NANDN U2325 ( .A(n1279), .B(n1278), .Z(n1208) );
  NAND U2326 ( .A(n1209), .B(n1208), .Z(n1210) );
  NANDN U2327 ( .A(n1211), .B(n1210), .Z(n1213) );
  ANDN U2328 ( .B(b[55]), .A(n173), .Z(n1371) );
  NANDN U2329 ( .A(n1371), .B(n1370), .Z(n1212) );
  NAND U2330 ( .A(n1213), .B(n1212), .Z(n1214) );
  NANDN U2331 ( .A(n1215), .B(n1214), .Z(n1217) );
  ANDN U2332 ( .B(b[55]), .A(n174), .Z(n1377) );
  OR U2333 ( .A(n1377), .B(n1376), .Z(n1216) );
  AND U2334 ( .A(n1217), .B(n1216), .Z(n1276) );
  XOR U2335 ( .A(n1219), .B(n1218), .Z(n1277) );
  NANDN U2336 ( .A(n1276), .B(n1277), .Z(n1220) );
  NAND U2337 ( .A(n1221), .B(n1220), .Z(n1225) );
  NANDN U2338 ( .A(n1225), .B(n1224), .Z(n1227) );
  NAND U2339 ( .A(a[19]), .B(b[55]), .Z(n1386) );
  XNOR U2340 ( .A(n1225), .B(n1224), .Z(n1387) );
  NANDN U2341 ( .A(n1386), .B(n1387), .Z(n1226) );
  NAND U2342 ( .A(n1227), .B(n1226), .Z(n1228) );
  NANDN U2343 ( .A(n1229), .B(n1228), .Z(n1231) );
  NAND U2344 ( .A(a[20]), .B(b[55]), .Z(n1392) );
  NANDN U2345 ( .A(n1392), .B(n1393), .Z(n1230) );
  NAND U2346 ( .A(n1231), .B(n1230), .Z(n1235) );
  XOR U2347 ( .A(n1233), .B(n1232), .Z(n1234) );
  NANDN U2348 ( .A(n1235), .B(n1234), .Z(n1237) );
  ANDN U2349 ( .B(b[55]), .A(n21681), .Z(n1275) );
  NANDN U2350 ( .A(n1275), .B(n1274), .Z(n1236) );
  NAND U2351 ( .A(n1237), .B(n1236), .Z(n1238) );
  NANDN U2352 ( .A(n1239), .B(n1238), .Z(n1241) );
  ANDN U2353 ( .B(b[55]), .A(n177), .Z(n1273) );
  NANDN U2354 ( .A(n1273), .B(n1272), .Z(n1240) );
  NAND U2355 ( .A(n1241), .B(n1240), .Z(n1270) );
  NANDN U2356 ( .A(n1270), .B(n1271), .Z(n1244) );
  NAND U2357 ( .A(n1245), .B(n1244), .Z(n1246) );
  OR U2358 ( .A(n1247), .B(n1246), .Z(n1249) );
  XNOR U2359 ( .A(n1247), .B(n1246), .Z(n1411) );
  ANDN U2360 ( .B(b[55]), .A(n178), .Z(n1410) );
  OR U2361 ( .A(n1411), .B(n1410), .Z(n1248) );
  NAND U2362 ( .A(n1249), .B(n1248), .Z(n1253) );
  XOR U2363 ( .A(n1251), .B(n1250), .Z(n1252) );
  NANDN U2364 ( .A(n1253), .B(n1252), .Z(n1255) );
  NAND U2365 ( .A(a[25]), .B(b[55]), .Z(n1417) );
  NANDN U2366 ( .A(n1417), .B(n1416), .Z(n1254) );
  NAND U2367 ( .A(n1255), .B(n1254), .Z(n1259) );
  XOR U2368 ( .A(n1257), .B(n1256), .Z(n1258) );
  NANDN U2369 ( .A(n1259), .B(n1258), .Z(n1261) );
  ANDN U2370 ( .B(b[55]), .A(n179), .Z(n1269) );
  NANDN U2371 ( .A(n1269), .B(n1268), .Z(n1260) );
  AND U2372 ( .A(n1261), .B(n1260), .Z(n1262) );
  OR U2373 ( .A(n1263), .B(n1262), .Z(n1265) );
  XNOR U2374 ( .A(n1263), .B(n1262), .Z(n1266) );
  ANDN U2375 ( .B(b[55]), .A(n21716), .Z(n1267) );
  OR U2376 ( .A(n1266), .B(n1267), .Z(n1264) );
  AND U2377 ( .A(n1265), .B(n1264), .Z(n1435) );
  XOR U2378 ( .A(n1434), .B(n1435), .Z(n1437) );
  XNOR U2379 ( .A(n1436), .B(n1437), .Z(n1430) );
  XNOR U2380 ( .A(n1267), .B(n1266), .Z(n1426) );
  XOR U2381 ( .A(n1269), .B(n1268), .Z(n1422) );
  XNOR U2382 ( .A(n1271), .B(n1270), .Z(n1407) );
  XOR U2383 ( .A(n1273), .B(n1272), .Z(n1403) );
  XOR U2384 ( .A(n1275), .B(n1274), .Z(n1399) );
  NAND U2385 ( .A(a[19]), .B(b[54]), .Z(n1383) );
  XOR U2386 ( .A(n1277), .B(n1276), .Z(n1382) );
  NANDN U2387 ( .A(n1383), .B(n1382), .Z(n1385) );
  ANDN U2388 ( .B(b[54]), .A(n173), .Z(n1280) );
  XOR U2389 ( .A(n1279), .B(n1278), .Z(n1281) );
  OR U2390 ( .A(n1280), .B(n1281), .Z(n1369) );
  XNOR U2391 ( .A(n1281), .B(n1280), .Z(n1556) );
  XOR U2392 ( .A(n1283), .B(n1282), .Z(n1365) );
  XOR U2393 ( .A(n1285), .B(n1284), .Z(n1361) );
  XOR U2394 ( .A(n1287), .B(n1286), .Z(n1357) );
  XOR U2395 ( .A(n1289), .B(n1288), .Z(n1353) );
  ANDN U2396 ( .B(b[54]), .A(n21164), .Z(n1349) );
  XOR U2397 ( .A(n1291), .B(n1290), .Z(n1348) );
  OR U2398 ( .A(n1349), .B(n1348), .Z(n1351) );
  XOR U2399 ( .A(n1293), .B(n1292), .Z(n1344) );
  XNOR U2400 ( .A(n1295), .B(n1294), .Z(n1335) );
  XOR U2401 ( .A(n1297), .B(n1296), .Z(n1299) );
  AND U2402 ( .A(a[7]), .B(b[54]), .Z(n1298) );
  NANDN U2403 ( .A(n1299), .B(n1298), .Z(n1333) );
  XOR U2404 ( .A(n1299), .B(n1298), .Z(n1572) );
  XNOR U2405 ( .A(n1301), .B(n1300), .Z(n1323) );
  XNOR U2406 ( .A(n1303), .B(n1302), .Z(n1318) );
  XNOR U2407 ( .A(n1305), .B(n1304), .Z(n1314) );
  NAND U2408 ( .A(b[55]), .B(a[1]), .Z(n1307) );
  NAND U2409 ( .A(n1307), .B(n1306), .Z(n1310) );
  OR U2410 ( .A(n1307), .B(n1824), .Z(n1587) );
  NANDN U2411 ( .A(n1309), .B(n1587), .Z(n1308) );
  AND U2412 ( .A(n1310), .B(n1308), .Z(n1313) );
  XNOR U2413 ( .A(n1587), .B(n1309), .Z(n1311) );
  NAND U2414 ( .A(n1311), .B(n1310), .Z(n1583) );
  ANDN U2415 ( .B(b[54]), .A(n162), .Z(n1582) );
  OR U2416 ( .A(n1583), .B(n1582), .Z(n1312) );
  AND U2417 ( .A(n1313), .B(n1312), .Z(n1315) );
  OR U2418 ( .A(n1314), .B(n1315), .Z(n1317) );
  XNOR U2419 ( .A(n1315), .B(n1314), .Z(n1580) );
  ANDN U2420 ( .B(b[54]), .A(n21580), .Z(n1581) );
  OR U2421 ( .A(n1580), .B(n1581), .Z(n1316) );
  AND U2422 ( .A(n1317), .B(n1316), .Z(n1319) );
  OR U2423 ( .A(n1318), .B(n1319), .Z(n1321) );
  XNOR U2424 ( .A(n1319), .B(n1318), .Z(n1578) );
  ANDN U2425 ( .B(b[54]), .A(n163), .Z(n1579) );
  OR U2426 ( .A(n1578), .B(n1579), .Z(n1320) );
  AND U2427 ( .A(n1321), .B(n1320), .Z(n1322) );
  OR U2428 ( .A(n1323), .B(n1322), .Z(n1325) );
  XNOR U2429 ( .A(n1323), .B(n1322), .Z(n1606) );
  NAND U2430 ( .A(b[54]), .B(a[5]), .Z(n1607) );
  NANDN U2431 ( .A(n1606), .B(n1607), .Z(n1324) );
  NAND U2432 ( .A(n1325), .B(n1324), .Z(n1327) );
  AND U2433 ( .A(a[6]), .B(b[54]), .Z(n1326) );
  NANDN U2434 ( .A(n1327), .B(n1326), .Z(n1331) );
  XOR U2435 ( .A(n1327), .B(n1326), .Z(n1574) );
  XOR U2436 ( .A(n1329), .B(n1328), .Z(n1575) );
  NANDN U2437 ( .A(n1574), .B(n1575), .Z(n1330) );
  AND U2438 ( .A(n1331), .B(n1330), .Z(n1573) );
  OR U2439 ( .A(n1572), .B(n1573), .Z(n1332) );
  AND U2440 ( .A(n1333), .B(n1332), .Z(n1334) );
  OR U2441 ( .A(n1335), .B(n1334), .Z(n1337) );
  XNOR U2442 ( .A(n1335), .B(n1334), .Z(n1617) );
  NAND U2443 ( .A(a[8]), .B(b[54]), .Z(n1616) );
  OR U2444 ( .A(n1617), .B(n1616), .Z(n1336) );
  NAND U2445 ( .A(n1337), .B(n1336), .Z(n1340) );
  XOR U2446 ( .A(n1339), .B(n1338), .Z(n1341) );
  OR U2447 ( .A(n1340), .B(n1341), .Z(n1343) );
  ANDN U2448 ( .B(b[54]), .A(n21615), .Z(n1571) );
  XOR U2449 ( .A(n1341), .B(n1340), .Z(n1570) );
  NANDN U2450 ( .A(n1571), .B(n1570), .Z(n1342) );
  AND U2451 ( .A(n1343), .B(n1342), .Z(n1345) );
  OR U2452 ( .A(n1344), .B(n1345), .Z(n1347) );
  XNOR U2453 ( .A(n1345), .B(n1344), .Z(n1568) );
  ANDN U2454 ( .B(b[54]), .A(n168), .Z(n1569) );
  OR U2455 ( .A(n1568), .B(n1569), .Z(n1346) );
  NAND U2456 ( .A(n1347), .B(n1346), .Z(n1567) );
  XOR U2457 ( .A(n1349), .B(n1348), .Z(n1566) );
  NAND U2458 ( .A(n1567), .B(n1566), .Z(n1350) );
  NAND U2459 ( .A(n1351), .B(n1350), .Z(n1352) );
  NANDN U2460 ( .A(n1353), .B(n1352), .Z(n1355) );
  ANDN U2461 ( .B(b[54]), .A(n169), .Z(n1565) );
  NANDN U2462 ( .A(n1565), .B(n1564), .Z(n1354) );
  NAND U2463 ( .A(n1355), .B(n1354), .Z(n1356) );
  NANDN U2464 ( .A(n1357), .B(n1356), .Z(n1359) );
  ANDN U2465 ( .B(b[54]), .A(n170), .Z(n1639) );
  NANDN U2466 ( .A(n1639), .B(n1638), .Z(n1358) );
  NAND U2467 ( .A(n1359), .B(n1358), .Z(n1360) );
  NANDN U2468 ( .A(n1361), .B(n1360), .Z(n1363) );
  ANDN U2469 ( .B(b[54]), .A(n171), .Z(n1563) );
  NANDN U2470 ( .A(n1563), .B(n1562), .Z(n1362) );
  NAND U2471 ( .A(n1363), .B(n1362), .Z(n1364) );
  NANDN U2472 ( .A(n1365), .B(n1364), .Z(n1367) );
  ANDN U2473 ( .B(b[54]), .A(n172), .Z(n1561) );
  NANDN U2474 ( .A(n1561), .B(n1560), .Z(n1366) );
  NAND U2475 ( .A(n1367), .B(n1366), .Z(n1557) );
  NANDN U2476 ( .A(n1556), .B(n1557), .Z(n1368) );
  NAND U2477 ( .A(n1369), .B(n1368), .Z(n1373) );
  NANDN U2478 ( .A(n1373), .B(n1372), .Z(n1375) );
  NAND U2479 ( .A(a[17]), .B(b[54]), .Z(n1654) );
  XNOR U2480 ( .A(n1373), .B(n1372), .Z(n1655) );
  NANDN U2481 ( .A(n1654), .B(n1655), .Z(n1374) );
  NAND U2482 ( .A(n1375), .B(n1374), .Z(n1379) );
  XOR U2483 ( .A(n1377), .B(n1376), .Z(n1378) );
  NANDN U2484 ( .A(n1379), .B(n1378), .Z(n1381) );
  ANDN U2485 ( .B(b[54]), .A(n175), .Z(n1661) );
  XOR U2486 ( .A(n1379), .B(n1378), .Z(n1660) );
  OR U2487 ( .A(n1661), .B(n1660), .Z(n1380) );
  NAND U2488 ( .A(n1381), .B(n1380), .Z(n1553) );
  NANDN U2489 ( .A(n1553), .B(n1552), .Z(n1384) );
  NAND U2490 ( .A(n1385), .B(n1384), .Z(n1389) );
  XOR U2491 ( .A(n1387), .B(n1386), .Z(n1388) );
  NANDN U2492 ( .A(n1389), .B(n1388), .Z(n1391) );
  ANDN U2493 ( .B(b[54]), .A(n176), .Z(n1550) );
  NANDN U2494 ( .A(n1550), .B(n1551), .Z(n1390) );
  AND U2495 ( .A(n1391), .B(n1390), .Z(n1395) );
  XOR U2496 ( .A(n1393), .B(n1392), .Z(n1394) );
  NANDN U2497 ( .A(n1395), .B(n1394), .Z(n1397) );
  ANDN U2498 ( .B(b[54]), .A(n21681), .Z(n1547) );
  NANDN U2499 ( .A(n1547), .B(n1546), .Z(n1396) );
  NAND U2500 ( .A(n1397), .B(n1396), .Z(n1398) );
  NANDN U2501 ( .A(n1399), .B(n1398), .Z(n1401) );
  ANDN U2502 ( .B(b[54]), .A(n177), .Z(n1545) );
  NANDN U2503 ( .A(n1545), .B(n1544), .Z(n1400) );
  NAND U2504 ( .A(n1401), .B(n1400), .Z(n1402) );
  NANDN U2505 ( .A(n1403), .B(n1402), .Z(n1405) );
  ANDN U2506 ( .B(b[54]), .A(n21692), .Z(n1541) );
  NANDN U2507 ( .A(n1541), .B(n1540), .Z(n1404) );
  AND U2508 ( .A(n1405), .B(n1404), .Z(n1406) );
  OR U2509 ( .A(n1407), .B(n1406), .Z(n1409) );
  ANDN U2510 ( .B(b[54]), .A(n178), .Z(n1681) );
  XNOR U2511 ( .A(n1407), .B(n1406), .Z(n1680) );
  OR U2512 ( .A(n1681), .B(n1680), .Z(n1408) );
  NAND U2513 ( .A(n1409), .B(n1408), .Z(n1413) );
  XOR U2514 ( .A(n1411), .B(n1410), .Z(n1412) );
  OR U2515 ( .A(n1413), .B(n1412), .Z(n1415) );
  NAND U2516 ( .A(a[25]), .B(b[54]), .Z(n1687) );
  XOR U2517 ( .A(n1413), .B(n1412), .Z(n1686) );
  NANDN U2518 ( .A(n1687), .B(n1686), .Z(n1414) );
  NAND U2519 ( .A(n1415), .B(n1414), .Z(n1418) );
  OR U2520 ( .A(n1418), .B(n1419), .Z(n1421) );
  ANDN U2521 ( .B(b[54]), .A(n179), .Z(n1538) );
  XOR U2522 ( .A(n1419), .B(n1418), .Z(n1539) );
  NANDN U2523 ( .A(n1538), .B(n1539), .Z(n1420) );
  AND U2524 ( .A(n1421), .B(n1420), .Z(n1423) );
  OR U2525 ( .A(n1422), .B(n1423), .Z(n1425) );
  XNOR U2526 ( .A(n1423), .B(n1422), .Z(n1696) );
  ANDN U2527 ( .B(b[54]), .A(n21716), .Z(n1697) );
  OR U2528 ( .A(n1696), .B(n1697), .Z(n1424) );
  AND U2529 ( .A(n1425), .B(n1424), .Z(n1427) );
  OR U2530 ( .A(n1426), .B(n1427), .Z(n1429) );
  XNOR U2531 ( .A(n1427), .B(n1426), .Z(n1536) );
  ANDN U2532 ( .B(b[54]), .A(n180), .Z(n1537) );
  OR U2533 ( .A(n1536), .B(n1537), .Z(n1428) );
  AND U2534 ( .A(n1429), .B(n1428), .Z(n1431) );
  OR U2535 ( .A(n1430), .B(n1431), .Z(n1433) );
  XNOR U2536 ( .A(n1431), .B(n1430), .Z(n1534) );
  IV U2537 ( .A(a[29]), .Z(n21727) );
  ANDN U2538 ( .B(b[54]), .A(n21727), .Z(n1535) );
  OR U2539 ( .A(n1534), .B(n1535), .Z(n1432) );
  AND U2540 ( .A(n1433), .B(n1432), .Z(n1482) );
  NAND U2541 ( .A(a[29]), .B(b[55]), .Z(n1531) );
  NANDN U2542 ( .A(n1435), .B(n1434), .Z(n1439) );
  OR U2543 ( .A(n1437), .B(n1436), .Z(n1438) );
  NAND U2544 ( .A(n1439), .B(n1438), .Z(n1529) );
  OR U2545 ( .A(n1441), .B(n1440), .Z(n1445) );
  OR U2546 ( .A(n1443), .B(n1442), .Z(n1444) );
  AND U2547 ( .A(n1445), .B(n1444), .Z(n1492) );
  NAND U2548 ( .A(a[25]), .B(b[59]), .Z(n1525) );
  NANDN U2549 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U2550 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U2551 ( .A(n1451), .B(n1450), .Z(n1523) );
  ANDN U2552 ( .B(b[61]), .A(n21692), .Z(n1506) );
  OR U2553 ( .A(n1453), .B(n1452), .Z(n1457) );
  OR U2554 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U2555 ( .A(n1457), .B(n1456), .Z(n1504) );
  ANDN U2556 ( .B(b[63]), .A(n21681), .Z(n1512) );
  ANDN U2557 ( .B(a[22]), .A(n159), .Z(n1510) );
  OR U2558 ( .A(n1459), .B(n1458), .Z(n1463) );
  OR U2559 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U2560 ( .A(n1463), .B(n1462), .Z(n1511) );
  XNOR U2561 ( .A(n1510), .B(n1511), .Z(n1513) );
  XNOR U2562 ( .A(n1512), .B(n1513), .Z(n1505) );
  XNOR U2563 ( .A(n1504), .B(n1505), .Z(n1507) );
  XNOR U2564 ( .A(n1506), .B(n1507), .Z(n1519) );
  ANDN U2565 ( .B(b[60]), .A(n178), .Z(n1516) );
  OR U2566 ( .A(n1465), .B(n1464), .Z(n1469) );
  NANDN U2567 ( .A(n1467), .B(n1466), .Z(n1468) );
  AND U2568 ( .A(n1469), .B(n1468), .Z(n1517) );
  XNOR U2569 ( .A(n1516), .B(n1517), .Z(n1518) );
  XOR U2570 ( .A(n1519), .B(n1518), .Z(n1522) );
  XOR U2571 ( .A(n1523), .B(n1522), .Z(n1524) );
  ANDN U2572 ( .B(b[58]), .A(n179), .Z(n1498) );
  OR U2573 ( .A(n1471), .B(n1470), .Z(n1475) );
  OR U2574 ( .A(n1473), .B(n1472), .Z(n1474) );
  AND U2575 ( .A(n1475), .B(n1474), .Z(n1499) );
  XOR U2576 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U2577 ( .A(n1501), .B(n1500), .Z(n1493) );
  XNOR U2578 ( .A(n1492), .B(n1493), .Z(n1495) );
  NAND U2579 ( .A(a[27]), .B(b[57]), .Z(n1494) );
  XOR U2580 ( .A(n1495), .B(n1494), .Z(n1489) );
  ANDN U2581 ( .B(b[56]), .A(n180), .Z(n1486) );
  OR U2582 ( .A(n1477), .B(n1476), .Z(n1481) );
  OR U2583 ( .A(n1479), .B(n1478), .Z(n1480) );
  AND U2584 ( .A(n1481), .B(n1480), .Z(n1487) );
  XOR U2585 ( .A(n1486), .B(n1487), .Z(n1488) );
  XNOR U2586 ( .A(n1489), .B(n1488), .Z(n1528) );
  XNOR U2587 ( .A(n1529), .B(n1528), .Z(n1530) );
  XOR U2588 ( .A(n1531), .B(n1530), .Z(n1483) );
  OR U2589 ( .A(n1482), .B(n1483), .Z(n1485) );
  XOR U2590 ( .A(n1483), .B(n1482), .Z(n1710) );
  NAND U2591 ( .A(b[54]), .B(a[30]), .Z(n1711) );
  NAND U2592 ( .A(n1710), .B(n1711), .Z(n1484) );
  AND U2593 ( .A(n1485), .B(n1484), .Z(n1769) );
  XNOR U2594 ( .A(n1768), .B(n1769), .Z(n1771) );
  NAND U2595 ( .A(a[29]), .B(b[56]), .Z(n1763) );
  OR U2596 ( .A(n1487), .B(n1486), .Z(n1491) );
  NANDN U2597 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U2598 ( .A(n1491), .B(n1490), .Z(n1762) );
  XNOR U2599 ( .A(n1763), .B(n1762), .Z(n1765) );
  NAND U2600 ( .A(a[28]), .B(b[57]), .Z(n1729) );
  OR U2601 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U2602 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U2603 ( .A(n1497), .B(n1496), .Z(n1726) );
  ANDN U2604 ( .B(b[58]), .A(n21716), .Z(n1732) );
  OR U2605 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U2606 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U2607 ( .A(n1503), .B(n1502), .Z(n1733) );
  XNOR U2608 ( .A(n1732), .B(n1733), .Z(n1735) );
  NAND U2609 ( .A(b[61]), .B(a[24]), .Z(n1740) );
  OR U2610 ( .A(n1505), .B(n1504), .Z(n1509) );
  OR U2611 ( .A(n1507), .B(n1506), .Z(n1508) );
  AND U2612 ( .A(n1509), .B(n1508), .Z(n1738) );
  ANDN U2613 ( .B(b[63]), .A(n177), .Z(n1746) );
  ANDN U2614 ( .B(a[23]), .A(n159), .Z(n1744) );
  OR U2615 ( .A(n1511), .B(n1510), .Z(n1515) );
  OR U2616 ( .A(n1513), .B(n1512), .Z(n1514) );
  AND U2617 ( .A(n1515), .B(n1514), .Z(n1745) );
  XNOR U2618 ( .A(n1744), .B(n1745), .Z(n1747) );
  XNOR U2619 ( .A(n1746), .B(n1747), .Z(n1739) );
  XNOR U2620 ( .A(n1738), .B(n1739), .Z(n1741) );
  XOR U2621 ( .A(n1740), .B(n1741), .Z(n1752) );
  NAND U2622 ( .A(a[25]), .B(b[60]), .Z(n1751) );
  OR U2623 ( .A(n1517), .B(n1516), .Z(n1521) );
  OR U2624 ( .A(n1519), .B(n1518), .Z(n1520) );
  NAND U2625 ( .A(n1521), .B(n1520), .Z(n1750) );
  XNOR U2626 ( .A(n1751), .B(n1750), .Z(n1753) );
  XNOR U2627 ( .A(n1752), .B(n1753), .Z(n1756) );
  OR U2628 ( .A(n1523), .B(n1522), .Z(n1527) );
  NANDN U2629 ( .A(n1525), .B(n1524), .Z(n1526) );
  NAND U2630 ( .A(n1527), .B(n1526), .Z(n1757) );
  XNOR U2631 ( .A(n1756), .B(n1757), .Z(n1759) );
  ANDN U2632 ( .B(b[59]), .A(n179), .Z(n1758) );
  XNOR U2633 ( .A(n1759), .B(n1758), .Z(n1734) );
  XOR U2634 ( .A(n1735), .B(n1734), .Z(n1727) );
  XNOR U2635 ( .A(n1726), .B(n1727), .Z(n1728) );
  XOR U2636 ( .A(n1729), .B(n1728), .Z(n1764) );
  OR U2637 ( .A(n1529), .B(n1528), .Z(n1533) );
  OR U2638 ( .A(n1531), .B(n1530), .Z(n1532) );
  NAND U2639 ( .A(n1533), .B(n1532), .Z(n1721) );
  XOR U2640 ( .A(n1720), .B(n1721), .Z(n1722) );
  ANDN U2641 ( .B(b[55]), .A(n181), .Z(n1723) );
  XOR U2642 ( .A(n1722), .B(n1723), .Z(n1770) );
  XOR U2643 ( .A(n1771), .B(n1770), .Z(n1716) );
  XNOR U2644 ( .A(n1535), .B(n1534), .Z(n1706) );
  XNOR U2645 ( .A(n1537), .B(n1536), .Z(n1702) );
  XNOR U2646 ( .A(n1539), .B(n1538), .Z(n1692) );
  NAND U2647 ( .A(a[24]), .B(b[53]), .Z(n1542) );
  NANDN U2648 ( .A(n1542), .B(n1543), .Z(n1679) );
  XOR U2649 ( .A(n1543), .B(n1542), .Z(n1781) );
  XNOR U2650 ( .A(n1545), .B(n1544), .Z(n1675) );
  NAND U2651 ( .A(a[22]), .B(b[53]), .Z(n1548) );
  NANDN U2652 ( .A(n1548), .B(n1549), .Z(n1673) );
  XOR U2653 ( .A(n1549), .B(n1548), .Z(n1787) );
  XNOR U2654 ( .A(n1551), .B(n1550), .Z(n1669) );
  NAND U2655 ( .A(b[53]), .B(a[20]), .Z(n1554) );
  XNOR U2656 ( .A(n1553), .B(n1552), .Z(n1555) );
  NANDN U2657 ( .A(n1554), .B(n1555), .Z(n1667) );
  XOR U2658 ( .A(n1555), .B(n1554), .Z(n1793) );
  NAND U2659 ( .A(a[17]), .B(b[53]), .Z(n1558) );
  XOR U2660 ( .A(n1557), .B(n1556), .Z(n1559) );
  NANDN U2661 ( .A(n1558), .B(n1559), .Z(n1653) );
  XOR U2662 ( .A(n1559), .B(n1558), .Z(n1799) );
  NAND U2663 ( .A(a[16]), .B(b[53]), .Z(n1648) );
  NANDN U2664 ( .A(n1648), .B(n1649), .Z(n1651) );
  NAND U2665 ( .A(a[15]), .B(b[53]), .Z(n1644) );
  NANDN U2666 ( .A(n1644), .B(n1645), .Z(n1647) );
  ANDN U2667 ( .B(b[53]), .A(n171), .Z(n1640) );
  XOR U2668 ( .A(n1565), .B(n1564), .Z(n1635) );
  XNOR U2669 ( .A(n1567), .B(n1566), .Z(n1631) );
  XNOR U2670 ( .A(n1569), .B(n1568), .Z(n1626) );
  XOR U2671 ( .A(n1571), .B(n1570), .Z(n1622) );
  XNOR U2672 ( .A(n1573), .B(n1572), .Z(n1613) );
  XOR U2673 ( .A(n1575), .B(n1574), .Z(n1577) );
  AND U2674 ( .A(a[7]), .B(b[53]), .Z(n1576) );
  NANDN U2675 ( .A(n1577), .B(n1576), .Z(n1611) );
  XOR U2676 ( .A(n1577), .B(n1576), .Z(n1812) );
  XNOR U2677 ( .A(n1579), .B(n1578), .Z(n1601) );
  XNOR U2678 ( .A(n1581), .B(n1580), .Z(n1596) );
  XNOR U2679 ( .A(n1583), .B(n1582), .Z(n1592) );
  NAND U2680 ( .A(b[54]), .B(a[1]), .Z(n1585) );
  NAND U2681 ( .A(n1585), .B(n1584), .Z(n1588) );
  OR U2682 ( .A(n1585), .B(n2146), .Z(n1827) );
  NANDN U2683 ( .A(n1587), .B(n1827), .Z(n1586) );
  AND U2684 ( .A(n1588), .B(n1586), .Z(n1591) );
  XNOR U2685 ( .A(n1827), .B(n1587), .Z(n1589) );
  NAND U2686 ( .A(n1589), .B(n1588), .Z(n1823) );
  ANDN U2687 ( .B(b[53]), .A(n162), .Z(n1822) );
  OR U2688 ( .A(n1823), .B(n1822), .Z(n1590) );
  AND U2689 ( .A(n1591), .B(n1590), .Z(n1593) );
  OR U2690 ( .A(n1592), .B(n1593), .Z(n1595) );
  XNOR U2691 ( .A(n1593), .B(n1592), .Z(n1820) );
  ANDN U2692 ( .B(b[53]), .A(n21580), .Z(n1821) );
  OR U2693 ( .A(n1820), .B(n1821), .Z(n1594) );
  AND U2694 ( .A(n1595), .B(n1594), .Z(n1597) );
  OR U2695 ( .A(n1596), .B(n1597), .Z(n1599) );
  XNOR U2696 ( .A(n1597), .B(n1596), .Z(n1818) );
  ANDN U2697 ( .B(b[53]), .A(n163), .Z(n1819) );
  OR U2698 ( .A(n1818), .B(n1819), .Z(n1598) );
  AND U2699 ( .A(n1599), .B(n1598), .Z(n1600) );
  OR U2700 ( .A(n1601), .B(n1600), .Z(n1603) );
  XNOR U2701 ( .A(n1601), .B(n1600), .Z(n1846) );
  NAND U2702 ( .A(b[53]), .B(a[5]), .Z(n1847) );
  NANDN U2703 ( .A(n1846), .B(n1847), .Z(n1602) );
  NAND U2704 ( .A(n1603), .B(n1602), .Z(n1605) );
  AND U2705 ( .A(a[6]), .B(b[53]), .Z(n1604) );
  NANDN U2706 ( .A(n1605), .B(n1604), .Z(n1609) );
  XOR U2707 ( .A(n1605), .B(n1604), .Z(n1814) );
  XOR U2708 ( .A(n1607), .B(n1606), .Z(n1815) );
  NANDN U2709 ( .A(n1814), .B(n1815), .Z(n1608) );
  AND U2710 ( .A(n1609), .B(n1608), .Z(n1813) );
  OR U2711 ( .A(n1812), .B(n1813), .Z(n1610) );
  AND U2712 ( .A(n1611), .B(n1610), .Z(n1612) );
  OR U2713 ( .A(n1613), .B(n1612), .Z(n1615) );
  XNOR U2714 ( .A(n1613), .B(n1612), .Z(n1857) );
  NAND U2715 ( .A(a[8]), .B(b[53]), .Z(n1856) );
  OR U2716 ( .A(n1857), .B(n1856), .Z(n1614) );
  NAND U2717 ( .A(n1615), .B(n1614), .Z(n1618) );
  XOR U2718 ( .A(n1617), .B(n1616), .Z(n1619) );
  OR U2719 ( .A(n1618), .B(n1619), .Z(n1621) );
  ANDN U2720 ( .B(b[53]), .A(n21615), .Z(n1811) );
  XOR U2721 ( .A(n1619), .B(n1618), .Z(n1810) );
  NANDN U2722 ( .A(n1811), .B(n1810), .Z(n1620) );
  AND U2723 ( .A(n1621), .B(n1620), .Z(n1623) );
  OR U2724 ( .A(n1622), .B(n1623), .Z(n1625) );
  XNOR U2725 ( .A(n1623), .B(n1622), .Z(n1808) );
  ANDN U2726 ( .B(b[53]), .A(n168), .Z(n1809) );
  OR U2727 ( .A(n1808), .B(n1809), .Z(n1624) );
  AND U2728 ( .A(n1625), .B(n1624), .Z(n1627) );
  OR U2729 ( .A(n1626), .B(n1627), .Z(n1629) );
  XNOR U2730 ( .A(n1627), .B(n1626), .Z(n1806) );
  ANDN U2731 ( .B(b[53]), .A(n21164), .Z(n1807) );
  OR U2732 ( .A(n1806), .B(n1807), .Z(n1628) );
  NAND U2733 ( .A(n1629), .B(n1628), .Z(n1630) );
  NANDN U2734 ( .A(n1631), .B(n1630), .Z(n1633) );
  ANDN U2735 ( .B(b[53]), .A(n169), .Z(n1805) );
  NANDN U2736 ( .A(n1805), .B(n1804), .Z(n1632) );
  NAND U2737 ( .A(n1633), .B(n1632), .Z(n1634) );
  NANDN U2738 ( .A(n1635), .B(n1634), .Z(n1637) );
  ANDN U2739 ( .B(b[53]), .A(n170), .Z(n1803) );
  NANDN U2740 ( .A(n1803), .B(n1802), .Z(n1636) );
  AND U2741 ( .A(n1637), .B(n1636), .Z(n1641) );
  OR U2742 ( .A(n1640), .B(n1641), .Z(n1643) );
  XOR U2743 ( .A(n1639), .B(n1638), .Z(n1801) );
  XOR U2744 ( .A(n1641), .B(n1640), .Z(n1800) );
  NANDN U2745 ( .A(n1801), .B(n1800), .Z(n1642) );
  NAND U2746 ( .A(n1643), .B(n1642), .Z(n1883) );
  XNOR U2747 ( .A(n1645), .B(n1644), .Z(n1882) );
  NANDN U2748 ( .A(n1883), .B(n1882), .Z(n1646) );
  AND U2749 ( .A(n1647), .B(n1646), .Z(n1888) );
  XNOR U2750 ( .A(n1649), .B(n1648), .Z(n1889) );
  NANDN U2751 ( .A(n1888), .B(n1889), .Z(n1650) );
  NAND U2752 ( .A(n1651), .B(n1650), .Z(n1798) );
  NANDN U2753 ( .A(n1799), .B(n1798), .Z(n1652) );
  NAND U2754 ( .A(n1653), .B(n1652), .Z(n1657) );
  XOR U2755 ( .A(n1655), .B(n1654), .Z(n1656) );
  NANDN U2756 ( .A(n1657), .B(n1656), .Z(n1659) );
  ANDN U2757 ( .B(b[53]), .A(n175), .Z(n1899) );
  NANDN U2758 ( .A(n1899), .B(n1898), .Z(n1658) );
  NAND U2759 ( .A(n1659), .B(n1658), .Z(n1663) );
  XNOR U2760 ( .A(n1661), .B(n1660), .Z(n1662) );
  NANDN U2761 ( .A(n1663), .B(n1662), .Z(n1665) );
  NAND U2762 ( .A(a[19]), .B(b[53]), .Z(n1797) );
  XNOR U2763 ( .A(n1663), .B(n1662), .Z(n1796) );
  NANDN U2764 ( .A(n1797), .B(n1796), .Z(n1664) );
  AND U2765 ( .A(n1665), .B(n1664), .Z(n1792) );
  OR U2766 ( .A(n1793), .B(n1792), .Z(n1666) );
  NAND U2767 ( .A(n1667), .B(n1666), .Z(n1668) );
  NANDN U2768 ( .A(n1669), .B(n1668), .Z(n1671) );
  NAND U2769 ( .A(b[53]), .B(a[21]), .Z(n1788) );
  NANDN U2770 ( .A(n1788), .B(n1789), .Z(n1670) );
  NAND U2771 ( .A(n1671), .B(n1670), .Z(n1786) );
  NANDN U2772 ( .A(n1787), .B(n1786), .Z(n1672) );
  NAND U2773 ( .A(n1673), .B(n1672), .Z(n1674) );
  NANDN U2774 ( .A(n1675), .B(n1674), .Z(n1677) );
  NAND U2775 ( .A(a[23]), .B(b[53]), .Z(n1783) );
  NANDN U2776 ( .A(n1783), .B(n1782), .Z(n1676) );
  NAND U2777 ( .A(n1677), .B(n1676), .Z(n1780) );
  NANDN U2778 ( .A(n1781), .B(n1780), .Z(n1678) );
  NAND U2779 ( .A(n1679), .B(n1678), .Z(n1683) );
  XOR U2780 ( .A(n1681), .B(n1680), .Z(n1682) );
  NANDN U2781 ( .A(n1683), .B(n1682), .Z(n1685) );
  ANDN U2782 ( .B(b[53]), .A(n21703), .Z(n1923) );
  XOR U2783 ( .A(n1683), .B(n1682), .Z(n1922) );
  OR U2784 ( .A(n1923), .B(n1922), .Z(n1684) );
  AND U2785 ( .A(n1685), .B(n1684), .Z(n1688) );
  NAND U2786 ( .A(n1688), .B(n1689), .Z(n1691) );
  NAND U2787 ( .A(a[26]), .B(b[53]), .Z(n1929) );
  XNOR U2788 ( .A(n1689), .B(n1688), .Z(n1928) );
  OR U2789 ( .A(n1929), .B(n1928), .Z(n1690) );
  AND U2790 ( .A(n1691), .B(n1690), .Z(n1693) );
  OR U2791 ( .A(n1692), .B(n1693), .Z(n1695) );
  XNOR U2792 ( .A(n1693), .B(n1692), .Z(n1777) );
  NAND U2793 ( .A(a[27]), .B(b[53]), .Z(n1776) );
  OR U2794 ( .A(n1777), .B(n1776), .Z(n1694) );
  NAND U2795 ( .A(n1695), .B(n1694), .Z(n1699) );
  XOR U2796 ( .A(n1697), .B(n1696), .Z(n1698) );
  NANDN U2797 ( .A(n1699), .B(n1698), .Z(n1701) );
  ANDN U2798 ( .B(b[53]), .A(n180), .Z(n1775) );
  NANDN U2799 ( .A(n1775), .B(n1774), .Z(n1700) );
  AND U2800 ( .A(n1701), .B(n1700), .Z(n1703) );
  OR U2801 ( .A(n1702), .B(n1703), .Z(n1705) );
  XNOR U2802 ( .A(n1703), .B(n1702), .Z(n1940) );
  NAND U2803 ( .A(b[53]), .B(a[29]), .Z(n1941) );
  NANDN U2804 ( .A(n1940), .B(n1941), .Z(n1704) );
  AND U2805 ( .A(n1705), .B(n1704), .Z(n1707) );
  OR U2806 ( .A(n1706), .B(n1707), .Z(n1709) );
  XNOR U2807 ( .A(n1707), .B(n1706), .Z(n1946) );
  ANDN U2808 ( .B(b[53]), .A(n181), .Z(n1947) );
  OR U2809 ( .A(n1946), .B(n1947), .Z(n1708) );
  NAND U2810 ( .A(n1709), .B(n1708), .Z(n1713) );
  NANDN U2811 ( .A(n1713), .B(n1712), .Z(n1715) );
  NAND U2812 ( .A(a[31]), .B(b[53]), .Z(n1953) );
  NANDN U2813 ( .A(n1953), .B(n1952), .Z(n1714) );
  AND U2814 ( .A(n1715), .B(n1714), .Z(n1717) );
  OR U2815 ( .A(n1716), .B(n1717), .Z(n1719) );
  XNOR U2816 ( .A(n1717), .B(n1716), .Z(n1959) );
  NAND U2817 ( .A(a[32]), .B(b[53]), .Z(n1958) );
  OR U2818 ( .A(n1959), .B(n1958), .Z(n1718) );
  NAND U2819 ( .A(n1719), .B(n1718), .Z(n1971) );
  NAND U2820 ( .A(a[31]), .B(b[55]), .Z(n2027) );
  OR U2821 ( .A(n1721), .B(n1720), .Z(n1725) );
  NANDN U2822 ( .A(n1723), .B(n1722), .Z(n1724) );
  NAND U2823 ( .A(n1725), .B(n1724), .Z(n2025) );
  NAND U2824 ( .A(a[29]), .B(b[57]), .Z(n1991) );
  OR U2825 ( .A(n1727), .B(n1726), .Z(n1731) );
  OR U2826 ( .A(n1729), .B(n1728), .Z(n1730) );
  AND U2827 ( .A(n1731), .B(n1730), .Z(n1988) );
  ANDN U2828 ( .B(b[58]), .A(n180), .Z(n1994) );
  OR U2829 ( .A(n1733), .B(n1732), .Z(n1737) );
  OR U2830 ( .A(n1735), .B(n1734), .Z(n1736) );
  AND U2831 ( .A(n1737), .B(n1736), .Z(n1995) );
  XNOR U2832 ( .A(n1994), .B(n1995), .Z(n1997) );
  NAND U2833 ( .A(b[61]), .B(a[25]), .Z(n2008) );
  OR U2834 ( .A(n1739), .B(n1738), .Z(n1743) );
  NANDN U2835 ( .A(n1741), .B(n1740), .Z(n1742) );
  AND U2836 ( .A(n1743), .B(n1742), .Z(n2006) );
  ANDN U2837 ( .B(b[63]), .A(n21692), .Z(n2014) );
  ANDN U2838 ( .B(a[24]), .A(n159), .Z(n2012) );
  OR U2839 ( .A(n1745), .B(n1744), .Z(n1749) );
  OR U2840 ( .A(n1747), .B(n1746), .Z(n1748) );
  AND U2841 ( .A(n1749), .B(n1748), .Z(n2013) );
  XNOR U2842 ( .A(n2012), .B(n2013), .Z(n2015) );
  XNOR U2843 ( .A(n2014), .B(n2015), .Z(n2007) );
  XNOR U2844 ( .A(n2006), .B(n2007), .Z(n2009) );
  XOR U2845 ( .A(n2008), .B(n2009), .Z(n2020) );
  NAND U2846 ( .A(a[26]), .B(b[60]), .Z(n2019) );
  OR U2847 ( .A(n1751), .B(n1750), .Z(n1755) );
  NANDN U2848 ( .A(n1753), .B(n1752), .Z(n1754) );
  AND U2849 ( .A(n1755), .B(n1754), .Z(n2018) );
  XNOR U2850 ( .A(n2019), .B(n2018), .Z(n2021) );
  XNOR U2851 ( .A(n2020), .B(n2021), .Z(n2000) );
  OR U2852 ( .A(n1757), .B(n1756), .Z(n1761) );
  OR U2853 ( .A(n1759), .B(n1758), .Z(n1760) );
  AND U2854 ( .A(n1761), .B(n1760), .Z(n2001) );
  XNOR U2855 ( .A(n2000), .B(n2001), .Z(n2003) );
  ANDN U2856 ( .B(b[59]), .A(n21716), .Z(n2002) );
  XNOR U2857 ( .A(n2003), .B(n2002), .Z(n1996) );
  XOR U2858 ( .A(n1997), .B(n1996), .Z(n1989) );
  XNOR U2859 ( .A(n1988), .B(n1989), .Z(n1990) );
  XOR U2860 ( .A(n1991), .B(n1990), .Z(n1985) );
  ANDN U2861 ( .B(b[56]), .A(n181), .Z(n1982) );
  OR U2862 ( .A(n1763), .B(n1762), .Z(n1767) );
  NANDN U2863 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U2864 ( .A(n1767), .B(n1766), .Z(n1983) );
  XOR U2865 ( .A(n1982), .B(n1983), .Z(n1984) );
  XNOR U2866 ( .A(n1985), .B(n1984), .Z(n2024) );
  XNOR U2867 ( .A(n2025), .B(n2024), .Z(n2026) );
  XOR U2868 ( .A(n2027), .B(n2026), .Z(n1978) );
  ANDN U2869 ( .B(b[54]), .A(n182), .Z(n1976) );
  OR U2870 ( .A(n1769), .B(n1768), .Z(n1773) );
  OR U2871 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U2872 ( .A(n1773), .B(n1772), .Z(n1977) );
  XNOR U2873 ( .A(n1976), .B(n1977), .Z(n1979) );
  XOR U2874 ( .A(n1978), .B(n1979), .Z(n1970) );
  XOR U2875 ( .A(n1973), .B(n1972), .Z(n1964) );
  XOR U2876 ( .A(n1775), .B(n1774), .Z(n1936) );
  XOR U2877 ( .A(n1777), .B(n1776), .Z(n1778) );
  ANDN U2878 ( .B(b[52]), .A(n180), .Z(n1779) );
  OR U2879 ( .A(n1778), .B(n1779), .Z(n1935) );
  XNOR U2880 ( .A(n1779), .B(n1778), .Z(n2105) );
  NAND U2881 ( .A(a[26]), .B(b[52]), .Z(n1925) );
  XOR U2882 ( .A(n1781), .B(n1780), .Z(n1919) );
  NAND U2883 ( .A(b[52]), .B(a[25]), .Z(n1918) );
  OR U2884 ( .A(n1919), .B(n1918), .Z(n1921) );
  NAND U2885 ( .A(a[24]), .B(b[52]), .Z(n1785) );
  XNOR U2886 ( .A(n1783), .B(n1782), .Z(n1784) );
  NANDN U2887 ( .A(n1785), .B(n1784), .Z(n1917) );
  XOR U2888 ( .A(n1785), .B(n1784), .Z(n2108) );
  XOR U2889 ( .A(n1787), .B(n1786), .Z(n1913) );
  NAND U2890 ( .A(a[22]), .B(b[52]), .Z(n1791) );
  XNOR U2891 ( .A(n1789), .B(n1788), .Z(n1790) );
  NANDN U2892 ( .A(n1791), .B(n1790), .Z(n1911) );
  XOR U2893 ( .A(n1791), .B(n1790), .Z(n2113) );
  NAND U2894 ( .A(a[21]), .B(b[52]), .Z(n1795) );
  XOR U2895 ( .A(n1793), .B(n1792), .Z(n1794) );
  NANDN U2896 ( .A(n1795), .B(n1794), .Z(n1909) );
  XOR U2897 ( .A(n1795), .B(n1794), .Z(n2114) );
  XOR U2898 ( .A(n1797), .B(n1796), .Z(n1905) );
  XOR U2899 ( .A(n1799), .B(n1798), .Z(n1895) );
  NAND U2900 ( .A(b[52]), .B(a[18]), .Z(n1894) );
  OR U2901 ( .A(n1895), .B(n1894), .Z(n1897) );
  XOR U2902 ( .A(n1801), .B(n1800), .Z(n2208) );
  ANDN U2903 ( .B(b[52]), .A(n172), .Z(n2209) );
  ANDN U2904 ( .B(b[52]), .A(n171), .Z(n1878) );
  XOR U2905 ( .A(n1803), .B(n1802), .Z(n1879) );
  OR U2906 ( .A(n1878), .B(n1879), .Z(n1881) );
  XOR U2907 ( .A(n1805), .B(n1804), .Z(n1875) );
  XNOR U2908 ( .A(n1807), .B(n1806), .Z(n1870) );
  XNOR U2909 ( .A(n1809), .B(n1808), .Z(n1866) );
  XOR U2910 ( .A(n1811), .B(n1810), .Z(n1862) );
  XNOR U2911 ( .A(n1813), .B(n1812), .Z(n1853) );
  XOR U2912 ( .A(n1815), .B(n1814), .Z(n1817) );
  AND U2913 ( .A(a[7]), .B(b[52]), .Z(n1816) );
  NANDN U2914 ( .A(n1817), .B(n1816), .Z(n1851) );
  XOR U2915 ( .A(n1817), .B(n1816), .Z(n2134) );
  XNOR U2916 ( .A(n1819), .B(n1818), .Z(n1841) );
  XNOR U2917 ( .A(n1821), .B(n1820), .Z(n1836) );
  XNOR U2918 ( .A(n1823), .B(n1822), .Z(n1832) );
  NAND U2919 ( .A(b[53]), .B(a[1]), .Z(n1825) );
  NAND U2920 ( .A(n1825), .B(n1824), .Z(n1828) );
  OR U2921 ( .A(n1825), .B(n2372), .Z(n2149) );
  NANDN U2922 ( .A(n1827), .B(n2149), .Z(n1826) );
  AND U2923 ( .A(n1828), .B(n1826), .Z(n1831) );
  XNOR U2924 ( .A(n2149), .B(n1827), .Z(n1829) );
  NAND U2925 ( .A(n1829), .B(n1828), .Z(n2145) );
  ANDN U2926 ( .B(b[52]), .A(n162), .Z(n2144) );
  OR U2927 ( .A(n2145), .B(n2144), .Z(n1830) );
  AND U2928 ( .A(n1831), .B(n1830), .Z(n1833) );
  OR U2929 ( .A(n1832), .B(n1833), .Z(n1835) );
  XNOR U2930 ( .A(n1833), .B(n1832), .Z(n2142) );
  ANDN U2931 ( .B(b[52]), .A(n21580), .Z(n2143) );
  OR U2932 ( .A(n2142), .B(n2143), .Z(n1834) );
  AND U2933 ( .A(n1835), .B(n1834), .Z(n1837) );
  OR U2934 ( .A(n1836), .B(n1837), .Z(n1839) );
  XNOR U2935 ( .A(n1837), .B(n1836), .Z(n2140) );
  ANDN U2936 ( .B(b[52]), .A(n163), .Z(n2141) );
  OR U2937 ( .A(n2140), .B(n2141), .Z(n1838) );
  AND U2938 ( .A(n1839), .B(n1838), .Z(n1840) );
  OR U2939 ( .A(n1841), .B(n1840), .Z(n1843) );
  XNOR U2940 ( .A(n1841), .B(n1840), .Z(n2168) );
  NAND U2941 ( .A(b[52]), .B(a[5]), .Z(n2169) );
  NANDN U2942 ( .A(n2168), .B(n2169), .Z(n1842) );
  NAND U2943 ( .A(n1843), .B(n1842), .Z(n1845) );
  AND U2944 ( .A(a[6]), .B(b[52]), .Z(n1844) );
  NANDN U2945 ( .A(n1845), .B(n1844), .Z(n1849) );
  XOR U2946 ( .A(n1845), .B(n1844), .Z(n2136) );
  XOR U2947 ( .A(n1847), .B(n1846), .Z(n2137) );
  NANDN U2948 ( .A(n2136), .B(n2137), .Z(n1848) );
  AND U2949 ( .A(n1849), .B(n1848), .Z(n2135) );
  OR U2950 ( .A(n2134), .B(n2135), .Z(n1850) );
  AND U2951 ( .A(n1851), .B(n1850), .Z(n1852) );
  OR U2952 ( .A(n1853), .B(n1852), .Z(n1855) );
  XNOR U2953 ( .A(n1853), .B(n1852), .Z(n2179) );
  NAND U2954 ( .A(a[8]), .B(b[52]), .Z(n2178) );
  OR U2955 ( .A(n2179), .B(n2178), .Z(n1854) );
  NAND U2956 ( .A(n1855), .B(n1854), .Z(n1858) );
  XOR U2957 ( .A(n1857), .B(n1856), .Z(n1859) );
  OR U2958 ( .A(n1858), .B(n1859), .Z(n1861) );
  ANDN U2959 ( .B(b[52]), .A(n21615), .Z(n2133) );
  XOR U2960 ( .A(n1859), .B(n1858), .Z(n2132) );
  NANDN U2961 ( .A(n2133), .B(n2132), .Z(n1860) );
  AND U2962 ( .A(n1861), .B(n1860), .Z(n1863) );
  OR U2963 ( .A(n1862), .B(n1863), .Z(n1865) );
  XNOR U2964 ( .A(n1863), .B(n1862), .Z(n2130) );
  ANDN U2965 ( .B(b[52]), .A(n168), .Z(n2131) );
  OR U2966 ( .A(n2130), .B(n2131), .Z(n1864) );
  AND U2967 ( .A(n1865), .B(n1864), .Z(n1867) );
  OR U2968 ( .A(n1866), .B(n1867), .Z(n1869) );
  XNOR U2969 ( .A(n1867), .B(n1866), .Z(n2128) );
  ANDN U2970 ( .B(b[52]), .A(n21164), .Z(n2129) );
  OR U2971 ( .A(n2128), .B(n2129), .Z(n1868) );
  AND U2972 ( .A(n1869), .B(n1868), .Z(n1871) );
  OR U2973 ( .A(n1870), .B(n1871), .Z(n1873) );
  XNOR U2974 ( .A(n1871), .B(n1870), .Z(n2126) );
  ANDN U2975 ( .B(b[52]), .A(n169), .Z(n2127) );
  OR U2976 ( .A(n2126), .B(n2127), .Z(n1872) );
  NAND U2977 ( .A(n1873), .B(n1872), .Z(n1874) );
  NANDN U2978 ( .A(n1875), .B(n1874), .Z(n1877) );
  ANDN U2979 ( .B(b[52]), .A(n170), .Z(n2124) );
  NANDN U2980 ( .A(n2124), .B(n2125), .Z(n1876) );
  NAND U2981 ( .A(n1877), .B(n1876), .Z(n2122) );
  XOR U2982 ( .A(n1879), .B(n1878), .Z(n2123) );
  NAND U2983 ( .A(n2122), .B(n2123), .Z(n1880) );
  AND U2984 ( .A(n1881), .B(n1880), .Z(n2211) );
  XNOR U2985 ( .A(n1883), .B(n1882), .Z(n1885) );
  NAND U2986 ( .A(n1884), .B(n1885), .Z(n1887) );
  NAND U2987 ( .A(b[52]), .B(a[16]), .Z(n2218) );
  NANDN U2988 ( .A(n2218), .B(n2219), .Z(n1886) );
  NAND U2989 ( .A(n1887), .B(n1886), .Z(n1891) );
  XOR U2990 ( .A(n1889), .B(n1888), .Z(n1890) );
  NANDN U2991 ( .A(n1891), .B(n1890), .Z(n1893) );
  ANDN U2992 ( .B(b[52]), .A(n174), .Z(n2222) );
  OR U2993 ( .A(n2222), .B(n2223), .Z(n1892) );
  NAND U2994 ( .A(n1893), .B(n1892), .Z(n2121) );
  XOR U2995 ( .A(n1895), .B(n1894), .Z(n2120) );
  NANDN U2996 ( .A(n2121), .B(n2120), .Z(n1896) );
  AND U2997 ( .A(n1897), .B(n1896), .Z(n1900) );
  NANDN U2998 ( .A(n1900), .B(n1901), .Z(n1903) );
  XOR U2999 ( .A(n1901), .B(n1900), .Z(n2118) );
  NAND U3000 ( .A(a[19]), .B(b[52]), .Z(n2119) );
  OR U3001 ( .A(n2118), .B(n2119), .Z(n1902) );
  NAND U3002 ( .A(n1903), .B(n1902), .Z(n1904) );
  NANDN U3003 ( .A(n1905), .B(n1904), .Z(n1907) );
  NAND U3004 ( .A(a[20]), .B(b[52]), .Z(n2117) );
  XOR U3005 ( .A(n1905), .B(n1904), .Z(n2116) );
  OR U3006 ( .A(n2117), .B(n2116), .Z(n1906) );
  AND U3007 ( .A(n1907), .B(n1906), .Z(n2115) );
  OR U3008 ( .A(n2114), .B(n2115), .Z(n1908) );
  NAND U3009 ( .A(n1909), .B(n1908), .Z(n2112) );
  NANDN U3010 ( .A(n2113), .B(n2112), .Z(n1910) );
  NAND U3011 ( .A(n1911), .B(n1910), .Z(n1912) );
  NANDN U3012 ( .A(n1913), .B(n1912), .Z(n1915) );
  NAND U3013 ( .A(b[52]), .B(a[23]), .Z(n2110) );
  NANDN U3014 ( .A(n2110), .B(n2111), .Z(n1914) );
  NAND U3015 ( .A(n1915), .B(n1914), .Z(n2109) );
  NANDN U3016 ( .A(n2108), .B(n2109), .Z(n1916) );
  NAND U3017 ( .A(n1917), .B(n1916), .Z(n2107) );
  XOR U3018 ( .A(n1919), .B(n1918), .Z(n2106) );
  NAND U3019 ( .A(n2107), .B(n2106), .Z(n1920) );
  NAND U3020 ( .A(n1921), .B(n1920), .Z(n1924) );
  NANDN U3021 ( .A(n1925), .B(n1924), .Z(n1927) );
  XOR U3022 ( .A(n1923), .B(n1922), .Z(n2260) );
  NANDN U3023 ( .A(n2260), .B(n2261), .Z(n1926) );
  NAND U3024 ( .A(n1927), .B(n1926), .Z(n1931) );
  XNOR U3025 ( .A(n1929), .B(n1928), .Z(n1930) );
  NANDN U3026 ( .A(n1931), .B(n1930), .Z(n1933) );
  ANDN U3027 ( .B(b[52]), .A(n21716), .Z(n2267) );
  NANDN U3028 ( .A(n2267), .B(n2266), .Z(n1932) );
  AND U3029 ( .A(n1933), .B(n1932), .Z(n2104) );
  OR U3030 ( .A(n2105), .B(n2104), .Z(n1934) );
  AND U3031 ( .A(n1935), .B(n1934), .Z(n1937) );
  OR U3032 ( .A(n1936), .B(n1937), .Z(n1939) );
  XNOR U3033 ( .A(n1937), .B(n1936), .Z(n2102) );
  ANDN U3034 ( .B(b[52]), .A(n21727), .Z(n2103) );
  OR U3035 ( .A(n2102), .B(n2103), .Z(n1938) );
  NAND U3036 ( .A(n1939), .B(n1938), .Z(n1943) );
  XOR U3037 ( .A(n1941), .B(n1940), .Z(n1942) );
  NANDN U3038 ( .A(n1943), .B(n1942), .Z(n1945) );
  NAND U3039 ( .A(a[30]), .B(b[52]), .Z(n2098) );
  NANDN U3040 ( .A(n2098), .B(n2099), .Z(n1944) );
  NAND U3041 ( .A(n1945), .B(n1944), .Z(n1949) );
  XOR U3042 ( .A(n1947), .B(n1946), .Z(n1948) );
  NANDN U3043 ( .A(n1949), .B(n1948), .Z(n1951) );
  ANDN U3044 ( .B(b[52]), .A(n21740), .Z(n2097) );
  NANDN U3045 ( .A(n2097), .B(n2096), .Z(n1950) );
  AND U3046 ( .A(n1951), .B(n1950), .Z(n1954) );
  OR U3047 ( .A(n1954), .B(n1955), .Z(n1957) );
  ANDN U3048 ( .B(b[52]), .A(n182), .Z(n2095) );
  XOR U3049 ( .A(n1955), .B(n1954), .Z(n2094) );
  NANDN U3050 ( .A(n2095), .B(n2094), .Z(n1956) );
  AND U3051 ( .A(n1957), .B(n1956), .Z(n1960) );
  XOR U3052 ( .A(n1959), .B(n1958), .Z(n1961) );
  OR U3053 ( .A(n1960), .B(n1961), .Z(n1963) );
  ANDN U3054 ( .B(b[52]), .A(n21751), .Z(n2093) );
  XOR U3055 ( .A(n1961), .B(n1960), .Z(n2092) );
  NANDN U3056 ( .A(n2093), .B(n2092), .Z(n1962) );
  AND U3057 ( .A(n1963), .B(n1962), .Z(n1965) );
  OR U3058 ( .A(n1964), .B(n1965), .Z(n1967) );
  XNOR U3059 ( .A(n1965), .B(n1964), .Z(n2294) );
  NAND U3060 ( .A(b[52]), .B(a[34]), .Z(n2295) );
  NANDN U3061 ( .A(n2294), .B(n2295), .Z(n1966) );
  NAND U3062 ( .A(n1967), .B(n1966), .Z(n1968) );
  OR U3063 ( .A(n1969), .B(n1968), .Z(n2031) );
  XNOR U3064 ( .A(n1969), .B(n1968), .Z(n2301) );
  NAND U3065 ( .A(a[34]), .B(b[53]), .Z(n2035) );
  NANDN U3066 ( .A(n1971), .B(n1970), .Z(n1975) );
  NANDN U3067 ( .A(n1973), .B(n1972), .Z(n1974) );
  NAND U3068 ( .A(n1975), .B(n1974), .Z(n2033) );
  ANDN U3069 ( .B(b[54]), .A(n21751), .Z(n2086) );
  OR U3070 ( .A(n1977), .B(n1976), .Z(n1981) );
  OR U3071 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U3072 ( .A(n1981), .B(n1980), .Z(n2087) );
  XNOR U3073 ( .A(n2086), .B(n2087), .Z(n2089) );
  NAND U3074 ( .A(a[31]), .B(b[56]), .Z(n2081) );
  OR U3075 ( .A(n1983), .B(n1982), .Z(n1987) );
  NANDN U3076 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U3077 ( .A(n1987), .B(n1986), .Z(n2080) );
  XNOR U3078 ( .A(n2081), .B(n2080), .Z(n2083) );
  NAND U3079 ( .A(a[30]), .B(b[57]), .Z(n2047) );
  OR U3080 ( .A(n1989), .B(n1988), .Z(n1993) );
  OR U3081 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U3082 ( .A(n1993), .B(n1992), .Z(n2044) );
  ANDN U3083 ( .B(b[58]), .A(n21727), .Z(n2050) );
  OR U3084 ( .A(n1995), .B(n1994), .Z(n1999) );
  OR U3085 ( .A(n1997), .B(n1996), .Z(n1998) );
  AND U3086 ( .A(n1999), .B(n1998), .Z(n2051) );
  XNOR U3087 ( .A(n2050), .B(n2051), .Z(n2053) );
  OR U3088 ( .A(n2001), .B(n2000), .Z(n2005) );
  OR U3089 ( .A(n2003), .B(n2002), .Z(n2004) );
  AND U3090 ( .A(n2005), .B(n2004), .Z(n2057) );
  ANDN U3091 ( .B(b[61]), .A(n179), .Z(n2064) );
  OR U3092 ( .A(n2007), .B(n2006), .Z(n2011) );
  NANDN U3093 ( .A(n2009), .B(n2008), .Z(n2010) );
  AND U3094 ( .A(n2011), .B(n2010), .Z(n2062) );
  ANDN U3095 ( .B(b[63]), .A(n178), .Z(n2070) );
  ANDN U3096 ( .B(a[25]), .A(n159), .Z(n2068) );
  OR U3097 ( .A(n2013), .B(n2012), .Z(n2017) );
  OR U3098 ( .A(n2015), .B(n2014), .Z(n2016) );
  AND U3099 ( .A(n2017), .B(n2016), .Z(n2069) );
  XNOR U3100 ( .A(n2068), .B(n2069), .Z(n2071) );
  XNOR U3101 ( .A(n2070), .B(n2071), .Z(n2063) );
  XNOR U3102 ( .A(n2062), .B(n2063), .Z(n2065) );
  XNOR U3103 ( .A(n2064), .B(n2065), .Z(n2077) );
  ANDN U3104 ( .B(b[60]), .A(n21716), .Z(n2074) );
  OR U3105 ( .A(n2019), .B(n2018), .Z(n2023) );
  NANDN U3106 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U3107 ( .A(n2023), .B(n2022), .Z(n2075) );
  XOR U3108 ( .A(n2074), .B(n2075), .Z(n2076) );
  XOR U3109 ( .A(n2057), .B(n2056), .Z(n2059) );
  ANDN U3110 ( .B(b[59]), .A(n180), .Z(n2058) );
  XNOR U3111 ( .A(n2059), .B(n2058), .Z(n2052) );
  XOR U3112 ( .A(n2053), .B(n2052), .Z(n2045) );
  XNOR U3113 ( .A(n2044), .B(n2045), .Z(n2046) );
  XOR U3114 ( .A(n2047), .B(n2046), .Z(n2082) );
  OR U3115 ( .A(n2025), .B(n2024), .Z(n2029) );
  OR U3116 ( .A(n2027), .B(n2026), .Z(n2028) );
  NAND U3117 ( .A(n2029), .B(n2028), .Z(n2039) );
  XOR U3118 ( .A(n2038), .B(n2039), .Z(n2040) );
  ANDN U3119 ( .B(b[55]), .A(n182), .Z(n2041) );
  XOR U3120 ( .A(n2040), .B(n2041), .Z(n2088) );
  XOR U3121 ( .A(n2089), .B(n2088), .Z(n2032) );
  XOR U3122 ( .A(n2033), .B(n2032), .Z(n2034) );
  NANDN U3123 ( .A(n2301), .B(n2300), .Z(n2030) );
  AND U3124 ( .A(n2031), .B(n2030), .Z(n2594) );
  XNOR U3125 ( .A(n2595), .B(n2594), .Z(n2597) );
  NAND U3126 ( .A(a[35]), .B(b[53]), .Z(n2537) );
  OR U3127 ( .A(n2033), .B(n2032), .Z(n2037) );
  NANDN U3128 ( .A(n2035), .B(n2034), .Z(n2036) );
  AND U3129 ( .A(n2037), .B(n2036), .Z(n2534) );
  NAND U3130 ( .A(a[33]), .B(b[55]), .Z(n2543) );
  OR U3131 ( .A(n2039), .B(n2038), .Z(n2043) );
  NANDN U3132 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U3133 ( .A(n2043), .B(n2042), .Z(n2541) );
  OR U3134 ( .A(n2045), .B(n2044), .Z(n2049) );
  OR U3135 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U3136 ( .A(n2049), .B(n2048), .Z(n2546) );
  ANDN U3137 ( .B(b[58]), .A(n181), .Z(n2552) );
  OR U3138 ( .A(n2051), .B(n2050), .Z(n2055) );
  OR U3139 ( .A(n2053), .B(n2052), .Z(n2054) );
  AND U3140 ( .A(n2055), .B(n2054), .Z(n2553) );
  XNOR U3141 ( .A(n2552), .B(n2553), .Z(n2555) );
  NANDN U3142 ( .A(n2057), .B(n2056), .Z(n2061) );
  OR U3143 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U3144 ( .A(n2061), .B(n2060), .Z(n2577) );
  ANDN U3145 ( .B(b[61]), .A(n21716), .Z(n2560) );
  OR U3146 ( .A(n2063), .B(n2062), .Z(n2067) );
  OR U3147 ( .A(n2065), .B(n2064), .Z(n2066) );
  AND U3148 ( .A(n2067), .B(n2066), .Z(n2558) );
  ANDN U3149 ( .B(b[63]), .A(n21703), .Z(n2566) );
  ANDN U3150 ( .B(a[26]), .A(n159), .Z(n2564) );
  OR U3151 ( .A(n2069), .B(n2068), .Z(n2073) );
  OR U3152 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U3153 ( .A(n2073), .B(n2072), .Z(n2565) );
  XNOR U3154 ( .A(n2564), .B(n2565), .Z(n2567) );
  XNOR U3155 ( .A(n2566), .B(n2567), .Z(n2559) );
  XNOR U3156 ( .A(n2558), .B(n2559), .Z(n2561) );
  XNOR U3157 ( .A(n2560), .B(n2561), .Z(n2573) );
  ANDN U3158 ( .B(b[60]), .A(n180), .Z(n2570) );
  OR U3159 ( .A(n2075), .B(n2074), .Z(n2079) );
  NANDN U3160 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U3161 ( .A(n2079), .B(n2078), .Z(n2571) );
  XOR U3162 ( .A(n2570), .B(n2571), .Z(n2572) );
  XOR U3163 ( .A(n2577), .B(n2576), .Z(n2579) );
  ANDN U3164 ( .B(b[59]), .A(n21727), .Z(n2578) );
  XNOR U3165 ( .A(n2579), .B(n2578), .Z(n2554) );
  XOR U3166 ( .A(n2555), .B(n2554), .Z(n2547) );
  XNOR U3167 ( .A(n2546), .B(n2547), .Z(n2549) );
  NAND U3168 ( .A(a[31]), .B(b[57]), .Z(n2548) );
  XOR U3169 ( .A(n2549), .B(n2548), .Z(n2585) );
  ANDN U3170 ( .B(b[56]), .A(n182), .Z(n2582) );
  OR U3171 ( .A(n2081), .B(n2080), .Z(n2085) );
  NANDN U3172 ( .A(n2083), .B(n2082), .Z(n2084) );
  NAND U3173 ( .A(n2085), .B(n2084), .Z(n2583) );
  XOR U3174 ( .A(n2582), .B(n2583), .Z(n2584) );
  XNOR U3175 ( .A(n2585), .B(n2584), .Z(n2540) );
  XNOR U3176 ( .A(n2541), .B(n2540), .Z(n2542) );
  XOR U3177 ( .A(n2543), .B(n2542), .Z(n2591) );
  ANDN U3178 ( .B(b[54]), .A(n183), .Z(n2588) );
  OR U3179 ( .A(n2087), .B(n2086), .Z(n2091) );
  OR U3180 ( .A(n2089), .B(n2088), .Z(n2090) );
  AND U3181 ( .A(n2091), .B(n2090), .Z(n2589) );
  XOR U3182 ( .A(n2588), .B(n2589), .Z(n2590) );
  XNOR U3183 ( .A(n2591), .B(n2590), .Z(n2535) );
  XNOR U3184 ( .A(n2534), .B(n2535), .Z(n2536) );
  XOR U3185 ( .A(n2537), .B(n2536), .Z(n2596) );
  XOR U3186 ( .A(n2093), .B(n2092), .Z(n2291) );
  XOR U3187 ( .A(n2095), .B(n2094), .Z(n2287) );
  XOR U3188 ( .A(n2097), .B(n2096), .Z(n2282) );
  XNOR U3189 ( .A(n2099), .B(n2098), .Z(n2100) );
  ANDN U3190 ( .B(b[51]), .A(n21740), .Z(n2101) );
  OR U3191 ( .A(n2100), .B(n2101), .Z(n2281) );
  XNOR U3192 ( .A(n2101), .B(n2100), .Z(n2311) );
  XNOR U3193 ( .A(n2103), .B(n2102), .Z(n2276) );
  XNOR U3194 ( .A(n2105), .B(n2104), .Z(n2273) );
  XNOR U3195 ( .A(n2107), .B(n2106), .Z(n2257) );
  XOR U3196 ( .A(n2109), .B(n2108), .Z(n2253) );
  NAND U3197 ( .A(b[51]), .B(a[25]), .Z(n2252) );
  OR U3198 ( .A(n2253), .B(n2252), .Z(n2255) );
  XOR U3199 ( .A(n2111), .B(n2110), .Z(n2249) );
  NANDN U3200 ( .A(n157), .B(a[23]), .Z(n2244) );
  NAND U3201 ( .A(n2244), .B(n2245), .Z(n2247) );
  NAND U3202 ( .A(a[22]), .B(b[51]), .Z(n2241) );
  XOR U3203 ( .A(n2115), .B(n2114), .Z(n2240) );
  NANDN U3204 ( .A(n2241), .B(n2240), .Z(n2243) );
  XOR U3205 ( .A(n2117), .B(n2116), .Z(n2237) );
  XOR U3206 ( .A(n2119), .B(n2118), .Z(n2233) );
  XNOR U3207 ( .A(n2121), .B(n2120), .Z(n2229) );
  NAND U3208 ( .A(a[17]), .B(b[51]), .Z(n2217) );
  XNOR U3209 ( .A(n2123), .B(n2122), .Z(n2205) );
  XOR U3210 ( .A(n2125), .B(n2124), .Z(n2201) );
  XNOR U3211 ( .A(n2127), .B(n2126), .Z(n2196) );
  XNOR U3212 ( .A(n2129), .B(n2128), .Z(n2192) );
  XNOR U3213 ( .A(n2131), .B(n2130), .Z(n2188) );
  XOR U3214 ( .A(n2133), .B(n2132), .Z(n2184) );
  XNOR U3215 ( .A(n2135), .B(n2134), .Z(n2175) );
  XOR U3216 ( .A(n2137), .B(n2136), .Z(n2139) );
  AND U3217 ( .A(a[7]), .B(b[51]), .Z(n2138) );
  NANDN U3218 ( .A(n2139), .B(n2138), .Z(n2173) );
  XOR U3219 ( .A(n2139), .B(n2138), .Z(n2360) );
  XNOR U3220 ( .A(n2141), .B(n2140), .Z(n2163) );
  XNOR U3221 ( .A(n2143), .B(n2142), .Z(n2158) );
  XNOR U3222 ( .A(n2145), .B(n2144), .Z(n2154) );
  NAND U3223 ( .A(b[52]), .B(a[1]), .Z(n2147) );
  NAND U3224 ( .A(n2147), .B(n2146), .Z(n2150) );
  NANDN U3225 ( .A(n157), .B(a[0]), .Z(n2662) );
  OR U3226 ( .A(n2147), .B(n2662), .Z(n2375) );
  NANDN U3227 ( .A(n2149), .B(n2375), .Z(n2148) );
  AND U3228 ( .A(n2150), .B(n2148), .Z(n2153) );
  XNOR U3229 ( .A(n2375), .B(n2149), .Z(n2151) );
  NAND U3230 ( .A(n2151), .B(n2150), .Z(n2371) );
  ANDN U3231 ( .B(b[51]), .A(n162), .Z(n2370) );
  OR U3232 ( .A(n2371), .B(n2370), .Z(n2152) );
  AND U3233 ( .A(n2153), .B(n2152), .Z(n2155) );
  OR U3234 ( .A(n2154), .B(n2155), .Z(n2157) );
  XNOR U3235 ( .A(n2155), .B(n2154), .Z(n2368) );
  ANDN U3236 ( .B(b[51]), .A(n21580), .Z(n2369) );
  OR U3237 ( .A(n2368), .B(n2369), .Z(n2156) );
  AND U3238 ( .A(n2157), .B(n2156), .Z(n2159) );
  OR U3239 ( .A(n2158), .B(n2159), .Z(n2161) );
  XNOR U3240 ( .A(n2159), .B(n2158), .Z(n2366) );
  ANDN U3241 ( .B(b[51]), .A(n163), .Z(n2367) );
  OR U3242 ( .A(n2366), .B(n2367), .Z(n2160) );
  AND U3243 ( .A(n2161), .B(n2160), .Z(n2162) );
  OR U3244 ( .A(n2163), .B(n2162), .Z(n2165) );
  XNOR U3245 ( .A(n2163), .B(n2162), .Z(n2394) );
  NAND U3246 ( .A(b[51]), .B(a[5]), .Z(n2395) );
  NANDN U3247 ( .A(n2394), .B(n2395), .Z(n2164) );
  NAND U3248 ( .A(n2165), .B(n2164), .Z(n2167) );
  AND U3249 ( .A(a[6]), .B(b[51]), .Z(n2166) );
  NANDN U3250 ( .A(n2167), .B(n2166), .Z(n2171) );
  XOR U3251 ( .A(n2167), .B(n2166), .Z(n2362) );
  XOR U3252 ( .A(n2169), .B(n2168), .Z(n2363) );
  NANDN U3253 ( .A(n2362), .B(n2363), .Z(n2170) );
  AND U3254 ( .A(n2171), .B(n2170), .Z(n2361) );
  OR U3255 ( .A(n2360), .B(n2361), .Z(n2172) );
  AND U3256 ( .A(n2173), .B(n2172), .Z(n2174) );
  OR U3257 ( .A(n2175), .B(n2174), .Z(n2177) );
  XNOR U3258 ( .A(n2175), .B(n2174), .Z(n2405) );
  NAND U3259 ( .A(a[8]), .B(b[51]), .Z(n2404) );
  OR U3260 ( .A(n2405), .B(n2404), .Z(n2176) );
  NAND U3261 ( .A(n2177), .B(n2176), .Z(n2180) );
  XOR U3262 ( .A(n2179), .B(n2178), .Z(n2181) );
  OR U3263 ( .A(n2180), .B(n2181), .Z(n2183) );
  ANDN U3264 ( .B(b[51]), .A(n21615), .Z(n2359) );
  XOR U3265 ( .A(n2181), .B(n2180), .Z(n2358) );
  NANDN U3266 ( .A(n2359), .B(n2358), .Z(n2182) );
  AND U3267 ( .A(n2183), .B(n2182), .Z(n2185) );
  OR U3268 ( .A(n2184), .B(n2185), .Z(n2187) );
  XNOR U3269 ( .A(n2185), .B(n2184), .Z(n2356) );
  ANDN U3270 ( .B(b[51]), .A(n168), .Z(n2357) );
  OR U3271 ( .A(n2356), .B(n2357), .Z(n2186) );
  AND U3272 ( .A(n2187), .B(n2186), .Z(n2189) );
  OR U3273 ( .A(n2188), .B(n2189), .Z(n2191) );
  XNOR U3274 ( .A(n2189), .B(n2188), .Z(n2354) );
  ANDN U3275 ( .B(b[51]), .A(n21164), .Z(n2355) );
  OR U3276 ( .A(n2354), .B(n2355), .Z(n2190) );
  AND U3277 ( .A(n2191), .B(n2190), .Z(n2193) );
  OR U3278 ( .A(n2192), .B(n2193), .Z(n2195) );
  XNOR U3279 ( .A(n2193), .B(n2192), .Z(n2353) );
  ANDN U3280 ( .B(b[51]), .A(n169), .Z(n2352) );
  OR U3281 ( .A(n2353), .B(n2352), .Z(n2194) );
  AND U3282 ( .A(n2195), .B(n2194), .Z(n2197) );
  OR U3283 ( .A(n2196), .B(n2197), .Z(n2199) );
  XNOR U3284 ( .A(n2197), .B(n2196), .Z(n2429) );
  ANDN U3285 ( .B(b[51]), .A(n170), .Z(n2428) );
  OR U3286 ( .A(n2429), .B(n2428), .Z(n2198) );
  NAND U3287 ( .A(n2199), .B(n2198), .Z(n2200) );
  NANDN U3288 ( .A(n2201), .B(n2200), .Z(n2203) );
  ANDN U3289 ( .B(b[51]), .A(n171), .Z(n2435) );
  NANDN U3290 ( .A(n2435), .B(n2434), .Z(n2202) );
  NAND U3291 ( .A(n2203), .B(n2202), .Z(n2204) );
  NANDN U3292 ( .A(n2205), .B(n2204), .Z(n2207) );
  ANDN U3293 ( .B(b[51]), .A(n172), .Z(n2439) );
  OR U3294 ( .A(n2439), .B(n2438), .Z(n2206) );
  NAND U3295 ( .A(n2207), .B(n2206), .Z(n2213) );
  XOR U3296 ( .A(n2209), .B(n2208), .Z(n2210) );
  XOR U3297 ( .A(n2211), .B(n2210), .Z(n2212) );
  NANDN U3298 ( .A(n2213), .B(n2212), .Z(n2215) );
  NAND U3299 ( .A(a[16]), .B(b[51]), .Z(n2351) );
  XNOR U3300 ( .A(n2213), .B(n2212), .Z(n2350) );
  NANDN U3301 ( .A(n2351), .B(n2350), .Z(n2214) );
  NAND U3302 ( .A(n2215), .B(n2214), .Z(n2216) );
  NANDN U3303 ( .A(n2217), .B(n2216), .Z(n2221) );
  XNOR U3304 ( .A(n2219), .B(n2218), .Z(n2347) );
  NAND U3305 ( .A(n2346), .B(n2347), .Z(n2220) );
  NAND U3306 ( .A(n2221), .B(n2220), .Z(n2225) );
  XOR U3307 ( .A(n2223), .B(n2222), .Z(n2224) );
  NANDN U3308 ( .A(n2225), .B(n2224), .Z(n2227) );
  ANDN U3309 ( .B(b[51]), .A(n175), .Z(n2343) );
  XOR U3310 ( .A(n2225), .B(n2224), .Z(n2342) );
  OR U3311 ( .A(n2343), .B(n2342), .Z(n2226) );
  NAND U3312 ( .A(n2227), .B(n2226), .Z(n2228) );
  NANDN U3313 ( .A(n2229), .B(n2228), .Z(n2231) );
  ANDN U3314 ( .B(b[51]), .A(n21670), .Z(n2341) );
  NANDN U3315 ( .A(n2341), .B(n2340), .Z(n2230) );
  NAND U3316 ( .A(n2231), .B(n2230), .Z(n2232) );
  NANDN U3317 ( .A(n2233), .B(n2232), .Z(n2235) );
  ANDN U3318 ( .B(b[51]), .A(n176), .Z(n2339) );
  NANDN U3319 ( .A(n2339), .B(n2338), .Z(n2234) );
  NAND U3320 ( .A(n2235), .B(n2234), .Z(n2236) );
  NANDN U3321 ( .A(n2237), .B(n2236), .Z(n2239) );
  ANDN U3322 ( .B(b[51]), .A(n21681), .Z(n2461) );
  OR U3323 ( .A(n2461), .B(n2460), .Z(n2238) );
  NAND U3324 ( .A(n2239), .B(n2238), .Z(n2335) );
  XNOR U3325 ( .A(n2241), .B(n2240), .Z(n2334) );
  NANDN U3326 ( .A(n2335), .B(n2334), .Z(n2242) );
  NAND U3327 ( .A(n2243), .B(n2242), .Z(n2330) );
  XOR U3328 ( .A(n2245), .B(n2244), .Z(n2331) );
  NANDN U3329 ( .A(n2330), .B(n2331), .Z(n2246) );
  NAND U3330 ( .A(n2247), .B(n2246), .Z(n2248) );
  OR U3331 ( .A(n2249), .B(n2248), .Z(n2251) );
  NAND U3332 ( .A(a[24]), .B(b[51]), .Z(n2327) );
  XOR U3333 ( .A(n2249), .B(n2248), .Z(n2326) );
  NANDN U3334 ( .A(n2327), .B(n2326), .Z(n2250) );
  AND U3335 ( .A(n2251), .B(n2250), .Z(n2472) );
  XOR U3336 ( .A(n2253), .B(n2252), .Z(n2473) );
  NANDN U3337 ( .A(n2472), .B(n2473), .Z(n2254) );
  NAND U3338 ( .A(n2255), .B(n2254), .Z(n2256) );
  NANDN U3339 ( .A(n2257), .B(n2256), .Z(n2259) );
  NAND U3340 ( .A(b[51]), .B(a[26]), .Z(n2322) );
  NANDN U3341 ( .A(n2322), .B(n2323), .Z(n2258) );
  NAND U3342 ( .A(n2259), .B(n2258), .Z(n2263) );
  XOR U3343 ( .A(n2261), .B(n2260), .Z(n2262) );
  NANDN U3344 ( .A(n2263), .B(n2262), .Z(n2265) );
  ANDN U3345 ( .B(b[51]), .A(n21716), .Z(n2321) );
  NANDN U3346 ( .A(n2321), .B(n2320), .Z(n2264) );
  NAND U3347 ( .A(n2265), .B(n2264), .Z(n2269) );
  NANDN U3348 ( .A(n2269), .B(n2268), .Z(n2271) );
  NAND U3349 ( .A(b[51]), .B(a[28]), .Z(n2318) );
  XNOR U3350 ( .A(n2269), .B(n2268), .Z(n2319) );
  NANDN U3351 ( .A(n2318), .B(n2319), .Z(n2270) );
  NAND U3352 ( .A(n2271), .B(n2270), .Z(n2272) );
  OR U3353 ( .A(n2273), .B(n2272), .Z(n2275) );
  XNOR U3354 ( .A(n2273), .B(n2272), .Z(n2316) );
  NAND U3355 ( .A(b[51]), .B(a[29]), .Z(n2317) );
  NANDN U3356 ( .A(n2316), .B(n2317), .Z(n2274) );
  AND U3357 ( .A(n2275), .B(n2274), .Z(n2277) );
  OR U3358 ( .A(n2276), .B(n2277), .Z(n2279) );
  XNOR U3359 ( .A(n2277), .B(n2276), .Z(n2314) );
  NAND U3360 ( .A(b[51]), .B(a[30]), .Z(n2315) );
  NANDN U3361 ( .A(n2314), .B(n2315), .Z(n2278) );
  AND U3362 ( .A(n2279), .B(n2278), .Z(n2310) );
  OR U3363 ( .A(n2311), .B(n2310), .Z(n2280) );
  AND U3364 ( .A(n2281), .B(n2280), .Z(n2283) );
  OR U3365 ( .A(n2282), .B(n2283), .Z(n2285) );
  XNOR U3366 ( .A(n2283), .B(n2282), .Z(n2498) );
  NAND U3367 ( .A(b[51]), .B(a[32]), .Z(n2499) );
  NANDN U3368 ( .A(n2498), .B(n2499), .Z(n2284) );
  AND U3369 ( .A(n2285), .B(n2284), .Z(n2286) );
  OR U3370 ( .A(n2287), .B(n2286), .Z(n2289) );
  XNOR U3371 ( .A(n2287), .B(n2286), .Z(n2506) );
  NAND U3372 ( .A(b[51]), .B(a[33]), .Z(n2507) );
  NANDN U3373 ( .A(n2506), .B(n2507), .Z(n2288) );
  AND U3374 ( .A(n2289), .B(n2288), .Z(n2290) );
  OR U3375 ( .A(n2291), .B(n2290), .Z(n2293) );
  XNOR U3376 ( .A(n2291), .B(n2290), .Z(n2308) );
  NAND U3377 ( .A(b[51]), .B(a[34]), .Z(n2309) );
  NANDN U3378 ( .A(n2308), .B(n2309), .Z(n2292) );
  NAND U3379 ( .A(n2293), .B(n2292), .Z(n2297) );
  XOR U3380 ( .A(n2295), .B(n2294), .Z(n2296) );
  NANDN U3381 ( .A(n2297), .B(n2296), .Z(n2299) );
  NAND U3382 ( .A(a[35]), .B(b[51]), .Z(n2515) );
  NANDN U3383 ( .A(n2515), .B(n2514), .Z(n2298) );
  NAND U3384 ( .A(n2299), .B(n2298), .Z(n2302) );
  OR U3385 ( .A(n2302), .B(n2303), .Z(n2305) );
  ANDN U3386 ( .B(b[51]), .A(n185), .Z(n2307) );
  XOR U3387 ( .A(n2303), .B(n2302), .Z(n2306) );
  NANDN U3388 ( .A(n2307), .B(n2306), .Z(n2304) );
  AND U3389 ( .A(n2305), .B(n2304), .Z(n2529) );
  XOR U3390 ( .A(n2528), .B(n2529), .Z(n2530) );
  IV U3391 ( .A(a[37]), .Z(n21772) );
  ANDN U3392 ( .B(b[51]), .A(n21772), .Z(n2531) );
  XOR U3393 ( .A(n2530), .B(n2531), .Z(n2525) );
  NAND U3394 ( .A(a[37]), .B(b[50]), .Z(n2520) );
  NANDN U3395 ( .A(n2520), .B(n2521), .Z(n2523) );
  NAND U3396 ( .A(a[35]), .B(b[50]), .Z(n2511) );
  XOR U3397 ( .A(n2309), .B(n2308), .Z(n2510) );
  NANDN U3398 ( .A(n2511), .B(n2510), .Z(n2513) );
  NAND U3399 ( .A(a[34]), .B(b[50]), .Z(n2504) );
  NAND U3400 ( .A(a[32]), .B(b[50]), .Z(n2312) );
  XOR U3401 ( .A(n2311), .B(n2310), .Z(n2313) );
  OR U3402 ( .A(n2312), .B(n2313), .Z(n2497) );
  XOR U3403 ( .A(n2313), .B(n2312), .Z(n2610) );
  NAND U3404 ( .A(a[31]), .B(b[50]), .Z(n2493) );
  XOR U3405 ( .A(n2315), .B(n2314), .Z(n2492) );
  NANDN U3406 ( .A(n2493), .B(n2492), .Z(n2495) );
  NAND U3407 ( .A(a[30]), .B(b[50]), .Z(n2489) );
  XOR U3408 ( .A(n2317), .B(n2316), .Z(n2488) );
  NANDN U3409 ( .A(n2489), .B(n2488), .Z(n2491) );
  XOR U3410 ( .A(n2319), .B(n2318), .Z(n2485) );
  ANDN U3411 ( .B(b[50]), .A(n180), .Z(n2480) );
  XOR U3412 ( .A(n2321), .B(n2320), .Z(n2481) );
  OR U3413 ( .A(n2480), .B(n2481), .Z(n2483) );
  NAND U3414 ( .A(b[50]), .B(a[27]), .Z(n2324) );
  XNOR U3415 ( .A(n2323), .B(n2322), .Z(n2325) );
  NANDN U3416 ( .A(n2324), .B(n2325), .Z(n2479) );
  XOR U3417 ( .A(n2325), .B(n2324), .Z(n2619) );
  NAND U3418 ( .A(a[25]), .B(b[50]), .Z(n2329) );
  XNOR U3419 ( .A(n2327), .B(n2326), .Z(n2328) );
  NANDN U3420 ( .A(n2329), .B(n2328), .Z(n2471) );
  XOR U3421 ( .A(n2329), .B(n2328), .Z(n2621) );
  NAND U3422 ( .A(a[24]), .B(b[50]), .Z(n2333) );
  XOR U3423 ( .A(n2331), .B(n2330), .Z(n2332) );
  NANDN U3424 ( .A(n2333), .B(n2332), .Z(n2469) );
  NAND U3425 ( .A(b[50]), .B(a[23]), .Z(n2336) );
  XNOR U3426 ( .A(n2335), .B(n2334), .Z(n2337) );
  NANDN U3427 ( .A(n2336), .B(n2337), .Z(n2467) );
  XOR U3428 ( .A(n2337), .B(n2336), .Z(n2623) );
  XNOR U3429 ( .A(n2339), .B(n2338), .Z(n2457) );
  XNOR U3430 ( .A(n2341), .B(n2340), .Z(n2453) );
  NAND U3431 ( .A(a[19]), .B(b[50]), .Z(n2344) );
  XNOR U3432 ( .A(n2343), .B(n2342), .Z(n2345) );
  NANDN U3433 ( .A(n2344), .B(n2345), .Z(n2451) );
  XOR U3434 ( .A(n2345), .B(n2344), .Z(n2740) );
  NAND U3435 ( .A(a[18]), .B(b[50]), .Z(n2349) );
  NANDN U3436 ( .A(n2349), .B(n2348), .Z(n2449) );
  XOR U3437 ( .A(n2349), .B(n2348), .Z(n2630) );
  XOR U3438 ( .A(n2351), .B(n2350), .Z(n2445) );
  NAND U3439 ( .A(a[15]), .B(b[50]), .Z(n2433) );
  NAND U3440 ( .A(a[14]), .B(b[50]), .Z(n2426) );
  NAND U3441 ( .A(a[13]), .B(b[50]), .Z(n2422) );
  XOR U3442 ( .A(n2353), .B(n2352), .Z(n2423) );
  OR U3443 ( .A(n2422), .B(n2423), .Z(n2425) );
  XNOR U3444 ( .A(n2355), .B(n2354), .Z(n2418) );
  XNOR U3445 ( .A(n2357), .B(n2356), .Z(n2414) );
  XOR U3446 ( .A(n2359), .B(n2358), .Z(n2410) );
  XNOR U3447 ( .A(n2361), .B(n2360), .Z(n2401) );
  XOR U3448 ( .A(n2363), .B(n2362), .Z(n2365) );
  AND U3449 ( .A(a[7]), .B(b[50]), .Z(n2364) );
  NANDN U3450 ( .A(n2365), .B(n2364), .Z(n2399) );
  XOR U3451 ( .A(n2365), .B(n2364), .Z(n2650) );
  XNOR U3452 ( .A(n2367), .B(n2366), .Z(n2389) );
  XNOR U3453 ( .A(n2369), .B(n2368), .Z(n2384) );
  XNOR U3454 ( .A(n2371), .B(n2370), .Z(n2380) );
  NAND U3455 ( .A(b[51]), .B(a[1]), .Z(n2373) );
  NAND U3456 ( .A(n2373), .B(n2372), .Z(n2376) );
  OR U3457 ( .A(n2373), .B(n2972), .Z(n2665) );
  NANDN U3458 ( .A(n2375), .B(n2665), .Z(n2374) );
  AND U3459 ( .A(n2376), .B(n2374), .Z(n2379) );
  XNOR U3460 ( .A(n2665), .B(n2375), .Z(n2377) );
  NAND U3461 ( .A(n2377), .B(n2376), .Z(n2661) );
  ANDN U3462 ( .B(b[50]), .A(n162), .Z(n2660) );
  OR U3463 ( .A(n2661), .B(n2660), .Z(n2378) );
  AND U3464 ( .A(n2379), .B(n2378), .Z(n2381) );
  OR U3465 ( .A(n2380), .B(n2381), .Z(n2383) );
  XNOR U3466 ( .A(n2381), .B(n2380), .Z(n2658) );
  ANDN U3467 ( .B(b[50]), .A(n21580), .Z(n2659) );
  OR U3468 ( .A(n2658), .B(n2659), .Z(n2382) );
  AND U3469 ( .A(n2383), .B(n2382), .Z(n2385) );
  OR U3470 ( .A(n2384), .B(n2385), .Z(n2387) );
  XNOR U3471 ( .A(n2385), .B(n2384), .Z(n2656) );
  ANDN U3472 ( .B(b[50]), .A(n163), .Z(n2657) );
  OR U3473 ( .A(n2656), .B(n2657), .Z(n2386) );
  AND U3474 ( .A(n2387), .B(n2386), .Z(n2388) );
  OR U3475 ( .A(n2389), .B(n2388), .Z(n2391) );
  XNOR U3476 ( .A(n2389), .B(n2388), .Z(n2684) );
  NAND U3477 ( .A(b[50]), .B(a[5]), .Z(n2685) );
  NANDN U3478 ( .A(n2684), .B(n2685), .Z(n2390) );
  NAND U3479 ( .A(n2391), .B(n2390), .Z(n2393) );
  AND U3480 ( .A(a[6]), .B(b[50]), .Z(n2392) );
  NANDN U3481 ( .A(n2393), .B(n2392), .Z(n2397) );
  XOR U3482 ( .A(n2393), .B(n2392), .Z(n2652) );
  XOR U3483 ( .A(n2395), .B(n2394), .Z(n2653) );
  NANDN U3484 ( .A(n2652), .B(n2653), .Z(n2396) );
  AND U3485 ( .A(n2397), .B(n2396), .Z(n2651) );
  OR U3486 ( .A(n2650), .B(n2651), .Z(n2398) );
  AND U3487 ( .A(n2399), .B(n2398), .Z(n2400) );
  OR U3488 ( .A(n2401), .B(n2400), .Z(n2403) );
  XNOR U3489 ( .A(n2401), .B(n2400), .Z(n2695) );
  NAND U3490 ( .A(a[8]), .B(b[50]), .Z(n2694) );
  OR U3491 ( .A(n2695), .B(n2694), .Z(n2402) );
  NAND U3492 ( .A(n2403), .B(n2402), .Z(n2406) );
  XOR U3493 ( .A(n2405), .B(n2404), .Z(n2407) );
  OR U3494 ( .A(n2406), .B(n2407), .Z(n2409) );
  ANDN U3495 ( .B(b[50]), .A(n21615), .Z(n2649) );
  XOR U3496 ( .A(n2407), .B(n2406), .Z(n2648) );
  NANDN U3497 ( .A(n2649), .B(n2648), .Z(n2408) );
  AND U3498 ( .A(n2409), .B(n2408), .Z(n2411) );
  OR U3499 ( .A(n2410), .B(n2411), .Z(n2413) );
  XNOR U3500 ( .A(n2411), .B(n2410), .Z(n2646) );
  ANDN U3501 ( .B(b[50]), .A(n168), .Z(n2647) );
  OR U3502 ( .A(n2646), .B(n2647), .Z(n2412) );
  AND U3503 ( .A(n2413), .B(n2412), .Z(n2415) );
  OR U3504 ( .A(n2414), .B(n2415), .Z(n2417) );
  XNOR U3505 ( .A(n2415), .B(n2414), .Z(n2644) );
  ANDN U3506 ( .B(b[50]), .A(n21164), .Z(n2645) );
  OR U3507 ( .A(n2644), .B(n2645), .Z(n2416) );
  AND U3508 ( .A(n2417), .B(n2416), .Z(n2419) );
  OR U3509 ( .A(n2418), .B(n2419), .Z(n2421) );
  XNOR U3510 ( .A(n2419), .B(n2418), .Z(n2643) );
  ANDN U3511 ( .B(b[50]), .A(n169), .Z(n2642) );
  OR U3512 ( .A(n2643), .B(n2642), .Z(n2420) );
  NAND U3513 ( .A(n2421), .B(n2420), .Z(n2640) );
  XOR U3514 ( .A(n2423), .B(n2422), .Z(n2641) );
  NANDN U3515 ( .A(n2640), .B(n2641), .Z(n2424) );
  AND U3516 ( .A(n2425), .B(n2424), .Z(n2427) );
  OR U3517 ( .A(n2426), .B(n2427), .Z(n2431) );
  XNOR U3518 ( .A(n2427), .B(n2426), .Z(n2720) );
  XOR U3519 ( .A(n2429), .B(n2428), .Z(n2721) );
  OR U3520 ( .A(n2720), .B(n2721), .Z(n2430) );
  NAND U3521 ( .A(n2431), .B(n2430), .Z(n2432) );
  NANDN U3522 ( .A(n2433), .B(n2432), .Z(n2437) );
  NAND U3523 ( .A(n2636), .B(n2637), .Z(n2436) );
  NAND U3524 ( .A(n2437), .B(n2436), .Z(n2441) );
  XOR U3525 ( .A(n2439), .B(n2438), .Z(n2440) );
  NANDN U3526 ( .A(n2441), .B(n2440), .Z(n2443) );
  ANDN U3527 ( .B(b[50]), .A(n173), .Z(n2633) );
  XOR U3528 ( .A(n2441), .B(n2440), .Z(n2632) );
  OR U3529 ( .A(n2633), .B(n2632), .Z(n2442) );
  AND U3530 ( .A(n2443), .B(n2442), .Z(n2444) );
  NANDN U3531 ( .A(n2445), .B(n2444), .Z(n2447) );
  XOR U3532 ( .A(n2445), .B(n2444), .Z(n2731) );
  NAND U3533 ( .A(b[50]), .B(a[17]), .Z(n2730) );
  OR U3534 ( .A(n2731), .B(n2730), .Z(n2446) );
  NAND U3535 ( .A(n2447), .B(n2446), .Z(n2631) );
  NANDN U3536 ( .A(n2630), .B(n2631), .Z(n2448) );
  NAND U3537 ( .A(n2449), .B(n2448), .Z(n2741) );
  NANDN U3538 ( .A(n2740), .B(n2741), .Z(n2450) );
  NAND U3539 ( .A(n2451), .B(n2450), .Z(n2452) );
  NANDN U3540 ( .A(n2453), .B(n2452), .Z(n2455) );
  NAND U3541 ( .A(a[20]), .B(b[50]), .Z(n2629) );
  NANDN U3542 ( .A(n2629), .B(n2628), .Z(n2454) );
  NAND U3543 ( .A(n2455), .B(n2454), .Z(n2456) );
  NANDN U3544 ( .A(n2457), .B(n2456), .Z(n2459) );
  NAND U3545 ( .A(a[21]), .B(b[50]), .Z(n2626) );
  NANDN U3546 ( .A(n2626), .B(n2627), .Z(n2458) );
  NAND U3547 ( .A(n2459), .B(n2458), .Z(n2463) );
  XOR U3548 ( .A(n2461), .B(n2460), .Z(n2462) );
  NANDN U3549 ( .A(n2463), .B(n2462), .Z(n2465) );
  ANDN U3550 ( .B(b[50]), .A(n177), .Z(n2755) );
  XOR U3551 ( .A(n2463), .B(n2462), .Z(n2754) );
  OR U3552 ( .A(n2755), .B(n2754), .Z(n2464) );
  NAND U3553 ( .A(n2465), .B(n2464), .Z(n2622) );
  OR U3554 ( .A(n2623), .B(n2622), .Z(n2466) );
  NAND U3555 ( .A(n2467), .B(n2466), .Z(n2763) );
  NANDN U3556 ( .A(n2762), .B(n2763), .Z(n2468) );
  AND U3557 ( .A(n2469), .B(n2468), .Z(n2620) );
  OR U3558 ( .A(n2621), .B(n2620), .Z(n2470) );
  NAND U3559 ( .A(n2471), .B(n2470), .Z(n2475) );
  XOR U3560 ( .A(n2473), .B(n2472), .Z(n2474) );
  NANDN U3561 ( .A(n2475), .B(n2474), .Z(n2477) );
  ANDN U3562 ( .B(b[50]), .A(n179), .Z(n2773) );
  NANDN U3563 ( .A(n2773), .B(n2772), .Z(n2476) );
  AND U3564 ( .A(n2477), .B(n2476), .Z(n2618) );
  NANDN U3565 ( .A(n2619), .B(n2618), .Z(n2478) );
  NAND U3566 ( .A(n2479), .B(n2478), .Z(n2617) );
  XOR U3567 ( .A(n2481), .B(n2480), .Z(n2616) );
  NANDN U3568 ( .A(n2617), .B(n2616), .Z(n2482) );
  NAND U3569 ( .A(n2483), .B(n2482), .Z(n2484) );
  OR U3570 ( .A(n2485), .B(n2484), .Z(n2487) );
  NAND U3571 ( .A(a[29]), .B(b[50]), .Z(n2789) );
  XOR U3572 ( .A(n2485), .B(n2484), .Z(n2788) );
  NANDN U3573 ( .A(n2789), .B(n2788), .Z(n2486) );
  AND U3574 ( .A(n2487), .B(n2486), .Z(n2613) );
  NANDN U3575 ( .A(n2613), .B(n2612), .Z(n2490) );
  AND U3576 ( .A(n2491), .B(n2490), .Z(n2795) );
  NANDN U3577 ( .A(n2795), .B(n2794), .Z(n2494) );
  NAND U3578 ( .A(n2495), .B(n2494), .Z(n2611) );
  NAND U3579 ( .A(n2610), .B(n2611), .Z(n2496) );
  AND U3580 ( .A(n2497), .B(n2496), .Z(n2501) );
  XOR U3581 ( .A(n2499), .B(n2498), .Z(n2500) );
  NANDN U3582 ( .A(n2501), .B(n2500), .Z(n2503) );
  NAND U3583 ( .A(a[33]), .B(b[50]), .Z(n2805) );
  NANDN U3584 ( .A(n2805), .B(n2804), .Z(n2502) );
  AND U3585 ( .A(n2503), .B(n2502), .Z(n2505) );
  OR U3586 ( .A(n2504), .B(n2505), .Z(n2509) );
  XNOR U3587 ( .A(n2505), .B(n2504), .Z(n2609) );
  XOR U3588 ( .A(n2507), .B(n2506), .Z(n2608) );
  NANDN U3589 ( .A(n2609), .B(n2608), .Z(n2508) );
  AND U3590 ( .A(n2509), .B(n2508), .Z(n2607) );
  NANDN U3591 ( .A(n2607), .B(n2606), .Z(n2512) );
  AND U3592 ( .A(n2513), .B(n2512), .Z(n2516) );
  NANDN U3593 ( .A(n2516), .B(n2517), .Z(n2519) );
  XOR U3594 ( .A(n2517), .B(n2516), .Z(n2603) );
  AND U3595 ( .A(a[36]), .B(b[50]), .Z(n2602) );
  NANDN U3596 ( .A(n2603), .B(n2602), .Z(n2518) );
  AND U3597 ( .A(n2519), .B(n2518), .Z(n2821) );
  XNOR U3598 ( .A(n2521), .B(n2520), .Z(n2820) );
  NANDN U3599 ( .A(n2821), .B(n2820), .Z(n2522) );
  NAND U3600 ( .A(n2523), .B(n2522), .Z(n2524) );
  OR U3601 ( .A(n2525), .B(n2524), .Z(n2527) );
  XNOR U3602 ( .A(n2525), .B(n2524), .Z(n2601) );
  ANDN U3603 ( .B(b[50]), .A(n186), .Z(n2600) );
  OR U3604 ( .A(n2601), .B(n2600), .Z(n2526) );
  NAND U3605 ( .A(n2527), .B(n2526), .Z(n2906) );
  XNOR U3606 ( .A(n2907), .B(n2906), .Z(n2909) );
  OR U3607 ( .A(n2529), .B(n2528), .Z(n2533) );
  NANDN U3608 ( .A(n2531), .B(n2530), .Z(n2532) );
  NAND U3609 ( .A(n2533), .B(n2532), .Z(n2835) );
  ANDN U3610 ( .B(b[53]), .A(n185), .Z(n2843) );
  OR U3611 ( .A(n2535), .B(n2534), .Z(n2539) );
  OR U3612 ( .A(n2537), .B(n2536), .Z(n2538) );
  NAND U3613 ( .A(n2539), .B(n2538), .Z(n2841) );
  OR U3614 ( .A(n2541), .B(n2540), .Z(n2545) );
  OR U3615 ( .A(n2543), .B(n2542), .Z(n2544) );
  AND U3616 ( .A(n2545), .B(n2544), .Z(n2894) );
  OR U3617 ( .A(n2547), .B(n2546), .Z(n2551) );
  OR U3618 ( .A(n2549), .B(n2548), .Z(n2550) );
  AND U3619 ( .A(n2551), .B(n2550), .Z(n2858) );
  ANDN U3620 ( .B(b[58]), .A(n21740), .Z(n2864) );
  OR U3621 ( .A(n2553), .B(n2552), .Z(n2557) );
  OR U3622 ( .A(n2555), .B(n2554), .Z(n2556) );
  AND U3623 ( .A(n2557), .B(n2556), .Z(n2865) );
  XNOR U3624 ( .A(n2864), .B(n2865), .Z(n2867) );
  NAND U3625 ( .A(b[61]), .B(a[28]), .Z(n2872) );
  OR U3626 ( .A(n2559), .B(n2558), .Z(n2563) );
  OR U3627 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U3628 ( .A(n2563), .B(n2562), .Z(n2870) );
  ANDN U3629 ( .B(b[63]), .A(n179), .Z(n2878) );
  ANDN U3630 ( .B(a[27]), .A(n159), .Z(n2876) );
  OR U3631 ( .A(n2565), .B(n2564), .Z(n2569) );
  OR U3632 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U3633 ( .A(n2569), .B(n2568), .Z(n2877) );
  XNOR U3634 ( .A(n2876), .B(n2877), .Z(n2879) );
  XNOR U3635 ( .A(n2878), .B(n2879), .Z(n2871) );
  XNOR U3636 ( .A(n2870), .B(n2871), .Z(n2873) );
  XOR U3637 ( .A(n2872), .B(n2873), .Z(n2884) );
  NAND U3638 ( .A(a[29]), .B(b[60]), .Z(n2883) );
  OR U3639 ( .A(n2571), .B(n2570), .Z(n2575) );
  NANDN U3640 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U3641 ( .A(n2575), .B(n2574), .Z(n2882) );
  XNOR U3642 ( .A(n2883), .B(n2882), .Z(n2885) );
  XNOR U3643 ( .A(n2884), .B(n2885), .Z(n2888) );
  NANDN U3644 ( .A(n2577), .B(n2576), .Z(n2581) );
  OR U3645 ( .A(n2579), .B(n2578), .Z(n2580) );
  AND U3646 ( .A(n2581), .B(n2580), .Z(n2889) );
  XNOR U3647 ( .A(n2888), .B(n2889), .Z(n2891) );
  ANDN U3648 ( .B(b[59]), .A(n181), .Z(n2890) );
  XNOR U3649 ( .A(n2891), .B(n2890), .Z(n2866) );
  XOR U3650 ( .A(n2867), .B(n2866), .Z(n2859) );
  XNOR U3651 ( .A(n2858), .B(n2859), .Z(n2861) );
  NAND U3652 ( .A(a[32]), .B(b[57]), .Z(n2860) );
  XOR U3653 ( .A(n2861), .B(n2860), .Z(n2855) );
  ANDN U3654 ( .B(b[56]), .A(n21751), .Z(n2852) );
  OR U3655 ( .A(n2583), .B(n2582), .Z(n2587) );
  NANDN U3656 ( .A(n2585), .B(n2584), .Z(n2586) );
  AND U3657 ( .A(n2587), .B(n2586), .Z(n2853) );
  XOR U3658 ( .A(n2852), .B(n2853), .Z(n2854) );
  XNOR U3659 ( .A(n2855), .B(n2854), .Z(n2895) );
  XNOR U3660 ( .A(n2894), .B(n2895), .Z(n2897) );
  NAND U3661 ( .A(a[34]), .B(b[55]), .Z(n2896) );
  XOR U3662 ( .A(n2897), .B(n2896), .Z(n2848) );
  ANDN U3663 ( .B(b[54]), .A(n184), .Z(n2846) );
  OR U3664 ( .A(n2589), .B(n2588), .Z(n2593) );
  NANDN U3665 ( .A(n2591), .B(n2590), .Z(n2592) );
  AND U3666 ( .A(n2593), .B(n2592), .Z(n2847) );
  XNOR U3667 ( .A(n2846), .B(n2847), .Z(n2849) );
  XOR U3668 ( .A(n2848), .B(n2849), .Z(n2840) );
  XOR U3669 ( .A(n2843), .B(n2842), .Z(n2903) );
  ANDN U3670 ( .B(b[52]), .A(n21772), .Z(n2900) );
  OR U3671 ( .A(n2595), .B(n2594), .Z(n2599) );
  NANDN U3672 ( .A(n2597), .B(n2596), .Z(n2598) );
  NAND U3673 ( .A(n2599), .B(n2598), .Z(n2901) );
  XNOR U3674 ( .A(n2900), .B(n2901), .Z(n2902) );
  XOR U3675 ( .A(n2903), .B(n2902), .Z(n2834) );
  XNOR U3676 ( .A(n2835), .B(n2834), .Z(n2837) );
  AND U3677 ( .A(a[38]), .B(b[51]), .Z(n2836) );
  XOR U3678 ( .A(n2837), .B(n2836), .Z(n2908) );
  XOR U3679 ( .A(n2909), .B(n2908), .Z(n2830) );
  XNOR U3680 ( .A(n2601), .B(n2600), .Z(n2827) );
  NAND U3681 ( .A(a[38]), .B(b[49]), .Z(n2822) );
  XOR U3682 ( .A(n2603), .B(n2602), .Z(n2605) );
  AND U3683 ( .A(a[37]), .B(b[49]), .Z(n2604) );
  NANDN U3684 ( .A(n2605), .B(n2604), .Z(n2819) );
  XOR U3685 ( .A(n2605), .B(n2604), .Z(n3135) );
  XOR U3686 ( .A(n2607), .B(n2606), .Z(n2815) );
  NAND U3687 ( .A(a[35]), .B(b[49]), .Z(n2811) );
  NANDN U3688 ( .A(n2811), .B(n2810), .Z(n2813) );
  ANDN U3689 ( .B(b[49]), .A(n21740), .Z(n2614) );
  OR U3690 ( .A(n2614), .B(n2615), .Z(n2793) );
  XNOR U3691 ( .A(n2615), .B(n2614), .Z(n2925) );
  NAND U3692 ( .A(a[30]), .B(b[49]), .Z(n2787) );
  NAND U3693 ( .A(a[29]), .B(b[49]), .Z(n2783) );
  XOR U3694 ( .A(n2617), .B(n2616), .Z(n2782) );
  NANDN U3695 ( .A(n2783), .B(n2782), .Z(n2785) );
  XOR U3696 ( .A(n2619), .B(n2618), .Z(n2779) );
  NAND U3697 ( .A(b[49]), .B(a[28]), .Z(n2778) );
  OR U3698 ( .A(n2779), .B(n2778), .Z(n2781) );
  XOR U3699 ( .A(n2621), .B(n2620), .Z(n2769) );
  NAND U3700 ( .A(a[24]), .B(b[49]), .Z(n2625) );
  XOR U3701 ( .A(n2623), .B(n2622), .Z(n2624) );
  NANDN U3702 ( .A(n2625), .B(n2624), .Z(n2761) );
  XOR U3703 ( .A(n2625), .B(n2624), .Z(n2936) );
  XNOR U3704 ( .A(n2627), .B(n2626), .Z(n2751) );
  XNOR U3705 ( .A(n2629), .B(n2628), .Z(n2747) );
  ANDN U3706 ( .B(b[49]), .A(n176), .Z(n2742) );
  XOR U3707 ( .A(n2631), .B(n2630), .Z(n2737) );
  NAND U3708 ( .A(a[18]), .B(b[49]), .Z(n2733) );
  NAND U3709 ( .A(a[17]), .B(b[49]), .Z(n2635) );
  XNOR U3710 ( .A(n2633), .B(n2632), .Z(n2634) );
  NANDN U3711 ( .A(n2635), .B(n2634), .Z(n2729) );
  XOR U3712 ( .A(n2635), .B(n2634), .Z(n2949) );
  NAND U3713 ( .A(b[49]), .B(a[16]), .Z(n2638) );
  NANDN U3714 ( .A(n2638), .B(n2639), .Z(n2727) );
  XOR U3715 ( .A(n2639), .B(n2638), .Z(n3043) );
  XOR U3716 ( .A(n2641), .B(n2640), .Z(n2717) );
  NAND U3717 ( .A(a[13]), .B(b[49]), .Z(n2712) );
  XOR U3718 ( .A(n2643), .B(n2642), .Z(n2713) );
  OR U3719 ( .A(n2712), .B(n2713), .Z(n2715) );
  XNOR U3720 ( .A(n2645), .B(n2644), .Z(n2708) );
  XNOR U3721 ( .A(n2647), .B(n2646), .Z(n2704) );
  XOR U3722 ( .A(n2649), .B(n2648), .Z(n2700) );
  XNOR U3723 ( .A(n2651), .B(n2650), .Z(n2691) );
  XOR U3724 ( .A(n2653), .B(n2652), .Z(n2655) );
  AND U3725 ( .A(a[7]), .B(b[49]), .Z(n2654) );
  NANDN U3726 ( .A(n2655), .B(n2654), .Z(n2689) );
  XOR U3727 ( .A(n2655), .B(n2654), .Z(n2960) );
  XNOR U3728 ( .A(n2657), .B(n2656), .Z(n2679) );
  XNOR U3729 ( .A(n2659), .B(n2658), .Z(n2674) );
  XNOR U3730 ( .A(n2661), .B(n2660), .Z(n2670) );
  NAND U3731 ( .A(b[50]), .B(a[1]), .Z(n2663) );
  NAND U3732 ( .A(n2663), .B(n2662), .Z(n2666) );
  OR U3733 ( .A(n2663), .B(n3206), .Z(n2975) );
  NANDN U3734 ( .A(n2665), .B(n2975), .Z(n2664) );
  AND U3735 ( .A(n2666), .B(n2664), .Z(n2669) );
  XNOR U3736 ( .A(n2975), .B(n2665), .Z(n2667) );
  NAND U3737 ( .A(n2667), .B(n2666), .Z(n2971) );
  ANDN U3738 ( .B(b[49]), .A(n162), .Z(n2970) );
  OR U3739 ( .A(n2971), .B(n2970), .Z(n2668) );
  AND U3740 ( .A(n2669), .B(n2668), .Z(n2671) );
  OR U3741 ( .A(n2670), .B(n2671), .Z(n2673) );
  XNOR U3742 ( .A(n2671), .B(n2670), .Z(n2968) );
  ANDN U3743 ( .B(b[49]), .A(n21580), .Z(n2969) );
  OR U3744 ( .A(n2968), .B(n2969), .Z(n2672) );
  AND U3745 ( .A(n2673), .B(n2672), .Z(n2675) );
  OR U3746 ( .A(n2674), .B(n2675), .Z(n2677) );
  XNOR U3747 ( .A(n2675), .B(n2674), .Z(n2966) );
  ANDN U3748 ( .B(b[49]), .A(n163), .Z(n2967) );
  OR U3749 ( .A(n2966), .B(n2967), .Z(n2676) );
  AND U3750 ( .A(n2677), .B(n2676), .Z(n2678) );
  OR U3751 ( .A(n2679), .B(n2678), .Z(n2681) );
  XNOR U3752 ( .A(n2679), .B(n2678), .Z(n2994) );
  NAND U3753 ( .A(b[49]), .B(a[5]), .Z(n2995) );
  NANDN U3754 ( .A(n2994), .B(n2995), .Z(n2680) );
  NAND U3755 ( .A(n2681), .B(n2680), .Z(n2683) );
  AND U3756 ( .A(a[6]), .B(b[49]), .Z(n2682) );
  NANDN U3757 ( .A(n2683), .B(n2682), .Z(n2687) );
  XOR U3758 ( .A(n2683), .B(n2682), .Z(n2962) );
  XOR U3759 ( .A(n2685), .B(n2684), .Z(n2963) );
  NANDN U3760 ( .A(n2962), .B(n2963), .Z(n2686) );
  AND U3761 ( .A(n2687), .B(n2686), .Z(n2961) );
  OR U3762 ( .A(n2960), .B(n2961), .Z(n2688) );
  AND U3763 ( .A(n2689), .B(n2688), .Z(n2690) );
  OR U3764 ( .A(n2691), .B(n2690), .Z(n2693) );
  XNOR U3765 ( .A(n2691), .B(n2690), .Z(n3005) );
  NAND U3766 ( .A(a[8]), .B(b[49]), .Z(n3004) );
  OR U3767 ( .A(n3005), .B(n3004), .Z(n2692) );
  NAND U3768 ( .A(n2693), .B(n2692), .Z(n2696) );
  XOR U3769 ( .A(n2695), .B(n2694), .Z(n2697) );
  OR U3770 ( .A(n2696), .B(n2697), .Z(n2699) );
  ANDN U3771 ( .B(b[49]), .A(n21615), .Z(n2959) );
  XOR U3772 ( .A(n2697), .B(n2696), .Z(n2958) );
  NANDN U3773 ( .A(n2959), .B(n2958), .Z(n2698) );
  AND U3774 ( .A(n2699), .B(n2698), .Z(n2701) );
  OR U3775 ( .A(n2700), .B(n2701), .Z(n2703) );
  XNOR U3776 ( .A(n2701), .B(n2700), .Z(n2956) );
  ANDN U3777 ( .B(b[49]), .A(n168), .Z(n2957) );
  OR U3778 ( .A(n2956), .B(n2957), .Z(n2702) );
  AND U3779 ( .A(n2703), .B(n2702), .Z(n2705) );
  OR U3780 ( .A(n2704), .B(n2705), .Z(n2707) );
  XNOR U3781 ( .A(n2705), .B(n2704), .Z(n2954) );
  ANDN U3782 ( .B(b[49]), .A(n21164), .Z(n2955) );
  OR U3783 ( .A(n2954), .B(n2955), .Z(n2706) );
  AND U3784 ( .A(n2707), .B(n2706), .Z(n2709) );
  OR U3785 ( .A(n2708), .B(n2709), .Z(n2711) );
  XNOR U3786 ( .A(n2709), .B(n2708), .Z(n2953) );
  ANDN U3787 ( .B(b[49]), .A(n169), .Z(n2952) );
  OR U3788 ( .A(n2953), .B(n2952), .Z(n2710) );
  NAND U3789 ( .A(n2711), .B(n2710), .Z(n3027) );
  XOR U3790 ( .A(n2713), .B(n2712), .Z(n3026) );
  NANDN U3791 ( .A(n3027), .B(n3026), .Z(n2714) );
  AND U3792 ( .A(n2715), .B(n2714), .Z(n2716) );
  OR U3793 ( .A(n2717), .B(n2716), .Z(n2719) );
  XNOR U3794 ( .A(n2717), .B(n2716), .Z(n2951) );
  AND U3795 ( .A(a[14]), .B(b[49]), .Z(n2950) );
  NANDN U3796 ( .A(n2951), .B(n2950), .Z(n2718) );
  AND U3797 ( .A(n2719), .B(n2718), .Z(n2723) );
  XOR U3798 ( .A(n2721), .B(n2720), .Z(n2722) );
  NANDN U3799 ( .A(n2723), .B(n2722), .Z(n2725) );
  NAND U3800 ( .A(a[15]), .B(b[49]), .Z(n3037) );
  NANDN U3801 ( .A(n3037), .B(n3036), .Z(n2724) );
  NAND U3802 ( .A(n2725), .B(n2724), .Z(n3042) );
  NANDN U3803 ( .A(n3043), .B(n3042), .Z(n2726) );
  AND U3804 ( .A(n2727), .B(n2726), .Z(n2948) );
  OR U3805 ( .A(n2949), .B(n2948), .Z(n2728) );
  NAND U3806 ( .A(n2729), .B(n2728), .Z(n2732) );
  NANDN U3807 ( .A(n2733), .B(n2732), .Z(n2735) );
  XOR U3808 ( .A(n2731), .B(n2730), .Z(n2946) );
  NAND U3809 ( .A(n2946), .B(n2947), .Z(n2734) );
  NAND U3810 ( .A(n2735), .B(n2734), .Z(n2736) );
  NANDN U3811 ( .A(n2737), .B(n2736), .Z(n2739) );
  NAND U3812 ( .A(a[19]), .B(b[49]), .Z(n2945) );
  NANDN U3813 ( .A(n2945), .B(n2944), .Z(n2738) );
  NAND U3814 ( .A(n2739), .B(n2738), .Z(n2743) );
  OR U3815 ( .A(n2742), .B(n2743), .Z(n2745) );
  XNOR U3816 ( .A(n2741), .B(n2740), .Z(n2942) );
  XOR U3817 ( .A(n2743), .B(n2742), .Z(n2943) );
  NANDN U3818 ( .A(n2942), .B(n2943), .Z(n2744) );
  NAND U3819 ( .A(n2745), .B(n2744), .Z(n2746) );
  NANDN U3820 ( .A(n2747), .B(n2746), .Z(n2749) );
  ANDN U3821 ( .B(b[49]), .A(n21681), .Z(n2941) );
  NANDN U3822 ( .A(n2941), .B(n2940), .Z(n2748) );
  NAND U3823 ( .A(n2749), .B(n2748), .Z(n2750) );
  NANDN U3824 ( .A(n2751), .B(n2750), .Z(n2753) );
  ANDN U3825 ( .B(b[49]), .A(n177), .Z(n3069) );
  OR U3826 ( .A(n3069), .B(n3068), .Z(n2752) );
  NAND U3827 ( .A(n2753), .B(n2752), .Z(n2757) );
  NAND U3828 ( .A(b[49]), .B(a[23]), .Z(n2756) );
  OR U3829 ( .A(n2757), .B(n2756), .Z(n2759) );
  XNOR U3830 ( .A(n2755), .B(n2754), .Z(n2939) );
  XOR U3831 ( .A(n2757), .B(n2756), .Z(n2938) );
  NAND U3832 ( .A(n2939), .B(n2938), .Z(n2758) );
  NAND U3833 ( .A(n2759), .B(n2758), .Z(n2937) );
  NANDN U3834 ( .A(n2936), .B(n2937), .Z(n2760) );
  NAND U3835 ( .A(n2761), .B(n2760), .Z(n2764) );
  XOR U3836 ( .A(n2763), .B(n2762), .Z(n2765) );
  NANDN U3837 ( .A(n2764), .B(n2765), .Z(n2767) );
  ANDN U3838 ( .B(b[49]), .A(n21703), .Z(n2935) );
  XOR U3839 ( .A(n2765), .B(n2764), .Z(n2934) );
  OR U3840 ( .A(n2935), .B(n2934), .Z(n2766) );
  NAND U3841 ( .A(n2767), .B(n2766), .Z(n2768) );
  NANDN U3842 ( .A(n2769), .B(n2768), .Z(n2771) );
  ANDN U3843 ( .B(b[49]), .A(n179), .Z(n2933) );
  NANDN U3844 ( .A(n2933), .B(n2932), .Z(n2770) );
  NAND U3845 ( .A(n2771), .B(n2770), .Z(n2775) );
  NANDN U3846 ( .A(n2775), .B(n2774), .Z(n2777) );
  XOR U3847 ( .A(n2775), .B(n2774), .Z(n2930) );
  NAND U3848 ( .A(a[27]), .B(b[49]), .Z(n2931) );
  OR U3849 ( .A(n2930), .B(n2931), .Z(n2776) );
  AND U3850 ( .A(n2777), .B(n2776), .Z(n2928) );
  XNOR U3851 ( .A(n2779), .B(n2778), .Z(n2929) );
  OR U3852 ( .A(n2928), .B(n2929), .Z(n2780) );
  NAND U3853 ( .A(n2781), .B(n2780), .Z(n2927) );
  NAND U3854 ( .A(n2927), .B(n2926), .Z(n2784) );
  NAND U3855 ( .A(n2785), .B(n2784), .Z(n2786) );
  NANDN U3856 ( .A(n2787), .B(n2786), .Z(n2791) );
  XNOR U3857 ( .A(n2789), .B(n2788), .Z(n3103) );
  NAND U3858 ( .A(n3102), .B(n3103), .Z(n2790) );
  NAND U3859 ( .A(n2791), .B(n2790), .Z(n2924) );
  OR U3860 ( .A(n2925), .B(n2924), .Z(n2792) );
  AND U3861 ( .A(n2793), .B(n2792), .Z(n2796) );
  OR U3862 ( .A(n2796), .B(n2797), .Z(n2799) );
  XOR U3863 ( .A(n2797), .B(n2796), .Z(n3112) );
  NAND U3864 ( .A(b[49]), .B(a[32]), .Z(n3113) );
  NAND U3865 ( .A(n3112), .B(n3113), .Z(n2798) );
  AND U3866 ( .A(n2799), .B(n2798), .Z(n2801) );
  OR U3867 ( .A(n2800), .B(n2801), .Z(n2803) );
  XNOR U3868 ( .A(n2801), .B(n2800), .Z(n3118) );
  ANDN U3869 ( .B(b[49]), .A(n21751), .Z(n3119) );
  OR U3870 ( .A(n3118), .B(n3119), .Z(n2802) );
  NAND U3871 ( .A(n2803), .B(n2802), .Z(n2807) );
  NANDN U3872 ( .A(n2807), .B(n2806), .Z(n2809) );
  NAND U3873 ( .A(a[34]), .B(b[49]), .Z(n2923) );
  NANDN U3874 ( .A(n2923), .B(n2922), .Z(n2808) );
  AND U3875 ( .A(n2809), .B(n2808), .Z(n2920) );
  NANDN U3876 ( .A(n2920), .B(n2921), .Z(n2812) );
  AND U3877 ( .A(n2813), .B(n2812), .Z(n2814) );
  OR U3878 ( .A(n2815), .B(n2814), .Z(n2817) );
  NAND U3879 ( .A(a[36]), .B(b[49]), .Z(n2917) );
  XNOR U3880 ( .A(n2815), .B(n2814), .Z(n2916) );
  OR U3881 ( .A(n2917), .B(n2916), .Z(n2816) );
  AND U3882 ( .A(n2817), .B(n2816), .Z(n3134) );
  OR U3883 ( .A(n3135), .B(n3134), .Z(n2818) );
  AND U3884 ( .A(n2819), .B(n2818), .Z(n2823) );
  OR U3885 ( .A(n2822), .B(n2823), .Z(n2825) );
  XOR U3886 ( .A(n2821), .B(n2820), .Z(n3141) );
  XNOR U3887 ( .A(n2823), .B(n2822), .Z(n3140) );
  OR U3888 ( .A(n3141), .B(n3140), .Z(n2824) );
  NAND U3889 ( .A(n2825), .B(n2824), .Z(n2826) );
  OR U3890 ( .A(n2827), .B(n2826), .Z(n2829) );
  XNOR U3891 ( .A(n2827), .B(n2826), .Z(n2915) );
  ANDN U3892 ( .B(b[49]), .A(n187), .Z(n2914) );
  OR U3893 ( .A(n2915), .B(n2914), .Z(n2828) );
  AND U3894 ( .A(n2829), .B(n2828), .Z(n2831) );
  OR U3895 ( .A(n2830), .B(n2831), .Z(n2833) );
  XNOR U3896 ( .A(n2831), .B(n2830), .Z(n2912) );
  NAND U3897 ( .A(b[49]), .B(a[40]), .Z(n2913) );
  NANDN U3898 ( .A(n2912), .B(n2913), .Z(n2832) );
  NAND U3899 ( .A(n2833), .B(n2832), .Z(n3407) );
  NAND U3900 ( .A(a[39]), .B(b[51]), .Z(n3415) );
  OR U3901 ( .A(n2835), .B(n2834), .Z(n2839) );
  NANDN U3902 ( .A(n2837), .B(n2836), .Z(n2838) );
  AND U3903 ( .A(n2839), .B(n2838), .Z(n3412) );
  NANDN U3904 ( .A(n2841), .B(n2840), .Z(n2845) );
  NANDN U3905 ( .A(n2843), .B(n2842), .Z(n2844) );
  NAND U3906 ( .A(n2845), .B(n2844), .Z(n3419) );
  ANDN U3907 ( .B(b[54]), .A(n185), .Z(n3472) );
  OR U3908 ( .A(n2847), .B(n2846), .Z(n2851) );
  OR U3909 ( .A(n2849), .B(n2848), .Z(n2850) );
  AND U3910 ( .A(n2851), .B(n2850), .Z(n3473) );
  XNOR U3911 ( .A(n3472), .B(n3473), .Z(n3475) );
  NAND U3912 ( .A(a[34]), .B(b[56]), .Z(n3467) );
  OR U3913 ( .A(n2853), .B(n2852), .Z(n2857) );
  NANDN U3914 ( .A(n2855), .B(n2854), .Z(n2856) );
  NAND U3915 ( .A(n2857), .B(n2856), .Z(n3466) );
  XNOR U3916 ( .A(n3467), .B(n3466), .Z(n3469) );
  NAND U3917 ( .A(a[33]), .B(b[57]), .Z(n3433) );
  OR U3918 ( .A(n2859), .B(n2858), .Z(n2863) );
  OR U3919 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U3920 ( .A(n2863), .B(n2862), .Z(n3430) );
  ANDN U3921 ( .B(b[58]), .A(n182), .Z(n3460) );
  OR U3922 ( .A(n2865), .B(n2864), .Z(n2869) );
  OR U3923 ( .A(n2867), .B(n2866), .Z(n2868) );
  AND U3924 ( .A(n2869), .B(n2868), .Z(n3461) );
  XNOR U3925 ( .A(n3460), .B(n3461), .Z(n3463) );
  NAND U3926 ( .A(b[61]), .B(a[29]), .Z(n3444) );
  OR U3927 ( .A(n2871), .B(n2870), .Z(n2875) );
  NANDN U3928 ( .A(n2873), .B(n2872), .Z(n2874) );
  AND U3929 ( .A(n2875), .B(n2874), .Z(n3442) );
  ANDN U3930 ( .B(b[63]), .A(n21716), .Z(n3450) );
  ANDN U3931 ( .B(a[28]), .A(n159), .Z(n3448) );
  OR U3932 ( .A(n2877), .B(n2876), .Z(n2881) );
  OR U3933 ( .A(n2879), .B(n2878), .Z(n2880) );
  AND U3934 ( .A(n2881), .B(n2880), .Z(n3449) );
  XNOR U3935 ( .A(n3448), .B(n3449), .Z(n3451) );
  XNOR U3936 ( .A(n3450), .B(n3451), .Z(n3443) );
  XNOR U3937 ( .A(n3442), .B(n3443), .Z(n3445) );
  XOR U3938 ( .A(n3444), .B(n3445), .Z(n3456) );
  NAND U3939 ( .A(a[30]), .B(b[60]), .Z(n3455) );
  OR U3940 ( .A(n2883), .B(n2882), .Z(n2887) );
  NANDN U3941 ( .A(n2885), .B(n2884), .Z(n2886) );
  AND U3942 ( .A(n2887), .B(n2886), .Z(n3454) );
  XNOR U3943 ( .A(n3455), .B(n3454), .Z(n3457) );
  XNOR U3944 ( .A(n3456), .B(n3457), .Z(n3436) );
  OR U3945 ( .A(n2889), .B(n2888), .Z(n2893) );
  OR U3946 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3947 ( .A(n2893), .B(n2892), .Z(n3437) );
  XNOR U3948 ( .A(n3436), .B(n3437), .Z(n3439) );
  ANDN U3949 ( .B(b[59]), .A(n21740), .Z(n3438) );
  XNOR U3950 ( .A(n3439), .B(n3438), .Z(n3462) );
  XOR U3951 ( .A(n3463), .B(n3462), .Z(n3431) );
  XNOR U3952 ( .A(n3430), .B(n3431), .Z(n3432) );
  XOR U3953 ( .A(n3433), .B(n3432), .Z(n3468) );
  OR U3954 ( .A(n2895), .B(n2894), .Z(n2899) );
  OR U3955 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U3956 ( .A(n2899), .B(n2898), .Z(n3425) );
  XOR U3957 ( .A(n3424), .B(n3425), .Z(n3426) );
  ANDN U3958 ( .B(b[55]), .A(n184), .Z(n3427) );
  XOR U3959 ( .A(n3426), .B(n3427), .Z(n3474) );
  XOR U3960 ( .A(n3475), .B(n3474), .Z(n3418) );
  XOR U3961 ( .A(n3419), .B(n3418), .Z(n3420) );
  NAND U3962 ( .A(a[37]), .B(b[53]), .Z(n3421) );
  ANDN U3963 ( .B(b[52]), .A(n186), .Z(n3478) );
  OR U3964 ( .A(n2901), .B(n2900), .Z(n2905) );
  OR U3965 ( .A(n2903), .B(n2902), .Z(n2904) );
  AND U3966 ( .A(n2905), .B(n2904), .Z(n3479) );
  XOR U3967 ( .A(n3478), .B(n3479), .Z(n3480) );
  XNOR U3968 ( .A(n3481), .B(n3480), .Z(n3413) );
  XNOR U3969 ( .A(n3412), .B(n3413), .Z(n3414) );
  XOR U3970 ( .A(n3415), .B(n3414), .Z(n3487) );
  ANDN U3971 ( .B(b[50]), .A(n188), .Z(n3484) );
  OR U3972 ( .A(n2907), .B(n2906), .Z(n2911) );
  OR U3973 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U3974 ( .A(n2911), .B(n2910), .Z(n3485) );
  XOR U3975 ( .A(n3484), .B(n3485), .Z(n3486) );
  XNOR U3976 ( .A(n3487), .B(n3486), .Z(n3406) );
  XNOR U3977 ( .A(n3407), .B(n3406), .Z(n3408) );
  XOR U3978 ( .A(n3409), .B(n3408), .Z(n3490) );
  NAND U3979 ( .A(a[41]), .B(b[48]), .Z(n3151) );
  XOR U3980 ( .A(n2913), .B(n2912), .Z(n3150) );
  NANDN U3981 ( .A(n3151), .B(n3150), .Z(n3153) );
  XOR U3982 ( .A(n2915), .B(n2914), .Z(n3146) );
  XNOR U3983 ( .A(n2917), .B(n2916), .Z(n2919) );
  AND U3984 ( .A(a[37]), .B(b[48]), .Z(n2918) );
  NANDN U3985 ( .A(n2919), .B(n2918), .Z(n3133) );
  XOR U3986 ( .A(n2919), .B(n2918), .Z(n3378) );
  XOR U3987 ( .A(n2921), .B(n2920), .Z(n3129) );
  AND U3988 ( .A(a[36]), .B(b[48]), .Z(n3128) );
  NANDN U3989 ( .A(n3129), .B(n3128), .Z(n3131) );
  XNOR U3990 ( .A(n2923), .B(n2922), .Z(n3124) );
  NAND U3991 ( .A(a[32]), .B(b[48]), .Z(n3108) );
  XOR U3992 ( .A(n2925), .B(n2924), .Z(n3109) );
  OR U3993 ( .A(n3108), .B(n3109), .Z(n3111) );
  XNOR U3994 ( .A(n2927), .B(n2926), .Z(n3099) );
  NAND U3995 ( .A(b[48]), .B(a[30]), .Z(n3098) );
  OR U3996 ( .A(n3099), .B(n3098), .Z(n3101) );
  NAND U3997 ( .A(a[29]), .B(b[48]), .Z(n3095) );
  XOR U3998 ( .A(n2929), .B(n2928), .Z(n3094) );
  NANDN U3999 ( .A(n3095), .B(n3094), .Z(n3097) );
  ANDN U4000 ( .B(b[48]), .A(n180), .Z(n3091) );
  XOR U4001 ( .A(n2931), .B(n2930), .Z(n3090) );
  OR U4002 ( .A(n3091), .B(n3090), .Z(n3093) );
  XOR U4003 ( .A(n2933), .B(n2932), .Z(n3087) );
  XNOR U4004 ( .A(n2935), .B(n2934), .Z(n3083) );
  XNOR U4005 ( .A(n2937), .B(n2936), .Z(n3079) );
  XOR U4006 ( .A(n2939), .B(n2938), .Z(n3075) );
  XNOR U4007 ( .A(n2941), .B(n2940), .Z(n3065) );
  NAND U4008 ( .A(a[21]), .B(b[48]), .Z(n3061) );
  XOR U4009 ( .A(n2943), .B(n2942), .Z(n3060) );
  NANDN U4010 ( .A(n3061), .B(n3060), .Z(n3063) );
  XNOR U4011 ( .A(n2945), .B(n2944), .Z(n3057) );
  XOR U4012 ( .A(n2947), .B(n2946), .Z(n3053) );
  XOR U4013 ( .A(n2949), .B(n2948), .Z(n3049) );
  NAND U4014 ( .A(a[15]), .B(b[48]), .Z(n3033) );
  XNOR U4015 ( .A(n2951), .B(n2950), .Z(n3032) );
  NANDN U4016 ( .A(n3033), .B(n3032), .Z(n3035) );
  NAND U4017 ( .A(a[13]), .B(b[48]), .Z(n3022) );
  XOR U4018 ( .A(n2953), .B(n2952), .Z(n3023) );
  OR U4019 ( .A(n3022), .B(n3023), .Z(n3025) );
  XNOR U4020 ( .A(n2955), .B(n2954), .Z(n3018) );
  XNOR U4021 ( .A(n2957), .B(n2956), .Z(n3014) );
  XOR U4022 ( .A(n2959), .B(n2958), .Z(n3010) );
  XNOR U4023 ( .A(n2961), .B(n2960), .Z(n3001) );
  XOR U4024 ( .A(n2963), .B(n2962), .Z(n2965) );
  AND U4025 ( .A(a[7]), .B(b[48]), .Z(n2964) );
  NANDN U4026 ( .A(n2965), .B(n2964), .Z(n2999) );
  XOR U4027 ( .A(n2965), .B(n2964), .Z(n3194) );
  XNOR U4028 ( .A(n2967), .B(n2966), .Z(n2989) );
  XNOR U4029 ( .A(n2969), .B(n2968), .Z(n2984) );
  XNOR U4030 ( .A(n2971), .B(n2970), .Z(n2980) );
  NAND U4031 ( .A(b[49]), .B(a[1]), .Z(n2973) );
  NAND U4032 ( .A(n2973), .B(n2972), .Z(n2976) );
  OR U4033 ( .A(n2973), .B(n3752), .Z(n3209) );
  NANDN U4034 ( .A(n2975), .B(n3209), .Z(n2974) );
  AND U4035 ( .A(n2976), .B(n2974), .Z(n2979) );
  XNOR U4036 ( .A(n3209), .B(n2975), .Z(n2977) );
  NAND U4037 ( .A(n2977), .B(n2976), .Z(n3205) );
  ANDN U4038 ( .B(b[48]), .A(n162), .Z(n3204) );
  OR U4039 ( .A(n3205), .B(n3204), .Z(n2978) );
  AND U4040 ( .A(n2979), .B(n2978), .Z(n2981) );
  OR U4041 ( .A(n2980), .B(n2981), .Z(n2983) );
  XNOR U4042 ( .A(n2981), .B(n2980), .Z(n3202) );
  ANDN U4043 ( .B(b[48]), .A(n21580), .Z(n3203) );
  OR U4044 ( .A(n3202), .B(n3203), .Z(n2982) );
  AND U4045 ( .A(n2983), .B(n2982), .Z(n2985) );
  OR U4046 ( .A(n2984), .B(n2985), .Z(n2987) );
  XNOR U4047 ( .A(n2985), .B(n2984), .Z(n3200) );
  ANDN U4048 ( .B(b[48]), .A(n163), .Z(n3201) );
  OR U4049 ( .A(n3200), .B(n3201), .Z(n2986) );
  AND U4050 ( .A(n2987), .B(n2986), .Z(n2988) );
  OR U4051 ( .A(n2989), .B(n2988), .Z(n2991) );
  XNOR U4052 ( .A(n2989), .B(n2988), .Z(n3228) );
  NAND U4053 ( .A(b[48]), .B(a[5]), .Z(n3229) );
  NANDN U4054 ( .A(n3228), .B(n3229), .Z(n2990) );
  NAND U4055 ( .A(n2991), .B(n2990), .Z(n2993) );
  AND U4056 ( .A(a[6]), .B(b[48]), .Z(n2992) );
  NANDN U4057 ( .A(n2993), .B(n2992), .Z(n2997) );
  XOR U4058 ( .A(n2993), .B(n2992), .Z(n3196) );
  XOR U4059 ( .A(n2995), .B(n2994), .Z(n3197) );
  NANDN U4060 ( .A(n3196), .B(n3197), .Z(n2996) );
  AND U4061 ( .A(n2997), .B(n2996), .Z(n3195) );
  OR U4062 ( .A(n3194), .B(n3195), .Z(n2998) );
  AND U4063 ( .A(n2999), .B(n2998), .Z(n3000) );
  OR U4064 ( .A(n3001), .B(n3000), .Z(n3003) );
  XNOR U4065 ( .A(n3001), .B(n3000), .Z(n3239) );
  NAND U4066 ( .A(a[8]), .B(b[48]), .Z(n3238) );
  OR U4067 ( .A(n3239), .B(n3238), .Z(n3002) );
  NAND U4068 ( .A(n3003), .B(n3002), .Z(n3006) );
  XOR U4069 ( .A(n3005), .B(n3004), .Z(n3007) );
  OR U4070 ( .A(n3006), .B(n3007), .Z(n3009) );
  ANDN U4071 ( .B(b[48]), .A(n21615), .Z(n3193) );
  XOR U4072 ( .A(n3007), .B(n3006), .Z(n3192) );
  NANDN U4073 ( .A(n3193), .B(n3192), .Z(n3008) );
  AND U4074 ( .A(n3009), .B(n3008), .Z(n3011) );
  OR U4075 ( .A(n3010), .B(n3011), .Z(n3013) );
  XNOR U4076 ( .A(n3011), .B(n3010), .Z(n3190) );
  ANDN U4077 ( .B(b[48]), .A(n168), .Z(n3191) );
  OR U4078 ( .A(n3190), .B(n3191), .Z(n3012) );
  AND U4079 ( .A(n3013), .B(n3012), .Z(n3015) );
  OR U4080 ( .A(n3014), .B(n3015), .Z(n3017) );
  XNOR U4081 ( .A(n3015), .B(n3014), .Z(n3188) );
  ANDN U4082 ( .B(b[48]), .A(n21164), .Z(n3189) );
  OR U4083 ( .A(n3188), .B(n3189), .Z(n3016) );
  AND U4084 ( .A(n3017), .B(n3016), .Z(n3019) );
  OR U4085 ( .A(n3018), .B(n3019), .Z(n3021) );
  XNOR U4086 ( .A(n3019), .B(n3018), .Z(n3186) );
  NAND U4087 ( .A(b[48]), .B(a[12]), .Z(n3187) );
  NANDN U4088 ( .A(n3186), .B(n3187), .Z(n3020) );
  NAND U4089 ( .A(n3021), .B(n3020), .Z(n3261) );
  XOR U4090 ( .A(n3023), .B(n3022), .Z(n3260) );
  NANDN U4091 ( .A(n3261), .B(n3260), .Z(n3024) );
  AND U4092 ( .A(n3025), .B(n3024), .Z(n3028) );
  NANDN U4093 ( .A(n3028), .B(n3029), .Z(n3031) );
  XOR U4094 ( .A(n3029), .B(n3028), .Z(n3267) );
  AND U4095 ( .A(a[14]), .B(b[48]), .Z(n3266) );
  NANDN U4096 ( .A(n3267), .B(n3266), .Z(n3030) );
  AND U4097 ( .A(n3031), .B(n3030), .Z(n3272) );
  NANDN U4098 ( .A(n3272), .B(n3273), .Z(n3034) );
  AND U4099 ( .A(n3035), .B(n3034), .Z(n3039) );
  NANDN U4100 ( .A(n3039), .B(n3038), .Z(n3041) );
  NAND U4101 ( .A(a[16]), .B(b[48]), .Z(n3279) );
  NANDN U4102 ( .A(n3279), .B(n3278), .Z(n3040) );
  NAND U4103 ( .A(n3041), .B(n3040), .Z(n3044) );
  NANDN U4104 ( .A(n3044), .B(n3045), .Z(n3047) );
  ANDN U4105 ( .B(b[48]), .A(n174), .Z(n3285) );
  XOR U4106 ( .A(n3045), .B(n3044), .Z(n3284) );
  OR U4107 ( .A(n3285), .B(n3284), .Z(n3046) );
  NAND U4108 ( .A(n3047), .B(n3046), .Z(n3048) );
  NANDN U4109 ( .A(n3049), .B(n3048), .Z(n3051) );
  ANDN U4110 ( .B(b[48]), .A(n175), .Z(n3185) );
  NANDN U4111 ( .A(n3185), .B(n3184), .Z(n3050) );
  NAND U4112 ( .A(n3051), .B(n3050), .Z(n3052) );
  NANDN U4113 ( .A(n3053), .B(n3052), .Z(n3055) );
  ANDN U4114 ( .B(b[48]), .A(n21670), .Z(n3183) );
  NANDN U4115 ( .A(n3183), .B(n3182), .Z(n3054) );
  NAND U4116 ( .A(n3055), .B(n3054), .Z(n3056) );
  NANDN U4117 ( .A(n3057), .B(n3056), .Z(n3059) );
  ANDN U4118 ( .B(b[48]), .A(n176), .Z(n3299) );
  NANDN U4119 ( .A(n3299), .B(n3298), .Z(n3058) );
  NAND U4120 ( .A(n3059), .B(n3058), .Z(n3181) );
  NANDN U4121 ( .A(n3181), .B(n3180), .Z(n3062) );
  NAND U4122 ( .A(n3063), .B(n3062), .Z(n3064) );
  NANDN U4123 ( .A(n3065), .B(n3064), .Z(n3067) );
  NAND U4124 ( .A(b[48]), .B(a[22]), .Z(n3178) );
  NANDN U4125 ( .A(n3178), .B(n3179), .Z(n3066) );
  NAND U4126 ( .A(n3067), .B(n3066), .Z(n3071) );
  XOR U4127 ( .A(n3069), .B(n3068), .Z(n3070) );
  NANDN U4128 ( .A(n3071), .B(n3070), .Z(n3073) );
  ANDN U4129 ( .B(b[48]), .A(n21692), .Z(n3175) );
  XOR U4130 ( .A(n3071), .B(n3070), .Z(n3174) );
  OR U4131 ( .A(n3175), .B(n3174), .Z(n3072) );
  NAND U4132 ( .A(n3073), .B(n3072), .Z(n3074) );
  NANDN U4133 ( .A(n3075), .B(n3074), .Z(n3077) );
  ANDN U4134 ( .B(b[48]), .A(n178), .Z(n3317) );
  NANDN U4135 ( .A(n3317), .B(n3316), .Z(n3076) );
  NAND U4136 ( .A(n3077), .B(n3076), .Z(n3078) );
  NANDN U4137 ( .A(n3079), .B(n3078), .Z(n3081) );
  ANDN U4138 ( .B(b[48]), .A(n21703), .Z(n3321) );
  OR U4139 ( .A(n3321), .B(n3320), .Z(n3080) );
  NAND U4140 ( .A(n3081), .B(n3080), .Z(n3082) );
  NANDN U4141 ( .A(n3083), .B(n3082), .Z(n3085) );
  ANDN U4142 ( .B(b[48]), .A(n179), .Z(n3173) );
  NANDN U4143 ( .A(n3173), .B(n3172), .Z(n3084) );
  NAND U4144 ( .A(n3085), .B(n3084), .Z(n3086) );
  NANDN U4145 ( .A(n3087), .B(n3086), .Z(n3089) );
  ANDN U4146 ( .B(b[48]), .A(n21716), .Z(n3171) );
  NANDN U4147 ( .A(n3171), .B(n3170), .Z(n3088) );
  AND U4148 ( .A(n3089), .B(n3088), .Z(n3334) );
  XOR U4149 ( .A(n3091), .B(n3090), .Z(n3335) );
  NANDN U4150 ( .A(n3334), .B(n3335), .Z(n3092) );
  NAND U4151 ( .A(n3093), .B(n3092), .Z(n3341) );
  XNOR U4152 ( .A(n3095), .B(n3094), .Z(n3340) );
  NANDN U4153 ( .A(n3341), .B(n3340), .Z(n3096) );
  NAND U4154 ( .A(n3097), .B(n3096), .Z(n3168) );
  XOR U4155 ( .A(n3099), .B(n3098), .Z(n3169) );
  NAND U4156 ( .A(n3168), .B(n3169), .Z(n3100) );
  NAND U4157 ( .A(n3101), .B(n3100), .Z(n3104) );
  NAND U4158 ( .A(n3104), .B(n3105), .Z(n3107) );
  NAND U4159 ( .A(a[31]), .B(b[48]), .Z(n3351) );
  XNOR U4160 ( .A(n3105), .B(n3104), .Z(n3350) );
  OR U4161 ( .A(n3351), .B(n3350), .Z(n3106) );
  AND U4162 ( .A(n3107), .B(n3106), .Z(n3357) );
  XNOR U4163 ( .A(n3109), .B(n3108), .Z(n3356) );
  OR U4164 ( .A(n3357), .B(n3356), .Z(n3110) );
  AND U4165 ( .A(n3111), .B(n3110), .Z(n3115) );
  NANDN U4166 ( .A(n3115), .B(n3114), .Z(n3117) );
  NAND U4167 ( .A(a[33]), .B(b[48]), .Z(n3165) );
  NANDN U4168 ( .A(n3165), .B(n3164), .Z(n3116) );
  NAND U4169 ( .A(n3117), .B(n3116), .Z(n3121) );
  XOR U4170 ( .A(n3119), .B(n3118), .Z(n3120) );
  NANDN U4171 ( .A(n3121), .B(n3120), .Z(n3123) );
  NAND U4172 ( .A(b[48]), .B(a[34]), .Z(n3365) );
  NAND U4173 ( .A(n3364), .B(n3365), .Z(n3122) );
  AND U4174 ( .A(n3123), .B(n3122), .Z(n3125) );
  OR U4175 ( .A(n3124), .B(n3125), .Z(n3127) );
  XNOR U4176 ( .A(n3125), .B(n3124), .Z(n3160) );
  NAND U4177 ( .A(b[48]), .B(a[35]), .Z(n3161) );
  NANDN U4178 ( .A(n3160), .B(n3161), .Z(n3126) );
  NAND U4179 ( .A(n3127), .B(n3126), .Z(n3373) );
  XNOR U4180 ( .A(n3129), .B(n3128), .Z(n3372) );
  NANDN U4181 ( .A(n3373), .B(n3372), .Z(n3130) );
  AND U4182 ( .A(n3131), .B(n3130), .Z(n3379) );
  OR U4183 ( .A(n3378), .B(n3379), .Z(n3132) );
  NAND U4184 ( .A(n3133), .B(n3132), .Z(n3136) );
  XOR U4185 ( .A(n3135), .B(n3134), .Z(n3137) );
  OR U4186 ( .A(n3136), .B(n3137), .Z(n3139) );
  XOR U4187 ( .A(n3137), .B(n3136), .Z(n3158) );
  NAND U4188 ( .A(b[48]), .B(a[38]), .Z(n3159) );
  NAND U4189 ( .A(n3158), .B(n3159), .Z(n3138) );
  NAND U4190 ( .A(n3139), .B(n3138), .Z(n3143) );
  XOR U4191 ( .A(n3141), .B(n3140), .Z(n3142) );
  NANDN U4192 ( .A(n3143), .B(n3142), .Z(n3145) );
  NAND U4193 ( .A(a[39]), .B(b[48]), .Z(n3389) );
  NANDN U4194 ( .A(n3389), .B(n3388), .Z(n3144) );
  AND U4195 ( .A(n3145), .B(n3144), .Z(n3147) );
  OR U4196 ( .A(n3146), .B(n3147), .Z(n3149) );
  XNOR U4197 ( .A(n3147), .B(n3146), .Z(n3157) );
  NAND U4198 ( .A(a[40]), .B(b[48]), .Z(n3156) );
  OR U4199 ( .A(n3157), .B(n3156), .Z(n3148) );
  AND U4200 ( .A(n3149), .B(n3148), .Z(n3154) );
  NANDN U4201 ( .A(n3154), .B(n3155), .Z(n3152) );
  AND U4202 ( .A(n3153), .B(n3152), .Z(n3491) );
  XOR U4203 ( .A(n3490), .B(n3491), .Z(n3493) );
  NAND U4204 ( .A(a[42]), .B(b[48]), .Z(n3492) );
  XOR U4205 ( .A(n3493), .B(n3492), .Z(n3402) );
  XNOR U4206 ( .A(n3155), .B(n3154), .Z(n3398) );
  XOR U4207 ( .A(n3157), .B(n3156), .Z(n3394) );
  NAND U4208 ( .A(a[39]), .B(b[47]), .Z(n3385) );
  NANDN U4209 ( .A(n3385), .B(n3384), .Z(n3387) );
  NAND U4210 ( .A(a[36]), .B(b[47]), .Z(n3163) );
  XOR U4211 ( .A(n3161), .B(n3160), .Z(n3162) );
  NANDN U4212 ( .A(n3163), .B(n3162), .Z(n3371) );
  NAND U4213 ( .A(a[34]), .B(b[47]), .Z(n3167) );
  NANDN U4214 ( .A(n3167), .B(n3166), .Z(n3363) );
  XOR U4215 ( .A(n3167), .B(n3166), .Z(n3701) );
  XNOR U4216 ( .A(n3169), .B(n3168), .Z(n3347) );
  NAND U4217 ( .A(b[47]), .B(a[31]), .Z(n3346) );
  OR U4218 ( .A(n3347), .B(n3346), .Z(n3349) );
  ANDN U4219 ( .B(b[47]), .A(n180), .Z(n3331) );
  XOR U4220 ( .A(n3171), .B(n3170), .Z(n3330) );
  OR U4221 ( .A(n3331), .B(n3330), .Z(n3333) );
  XOR U4222 ( .A(n3173), .B(n3172), .Z(n3327) );
  NAND U4223 ( .A(a[25]), .B(b[47]), .Z(n3315) );
  NAND U4224 ( .A(a[24]), .B(b[47]), .Z(n3176) );
  XNOR U4225 ( .A(n3175), .B(n3174), .Z(n3177) );
  NANDN U4226 ( .A(n3176), .B(n3177), .Z(n3313) );
  XOR U4227 ( .A(n3177), .B(n3176), .Z(n3719) );
  NAND U4228 ( .A(b[47]), .B(a[23]), .Z(n3308) );
  XNOR U4229 ( .A(n3179), .B(n3178), .Z(n3309) );
  NANDN U4230 ( .A(n3308), .B(n3309), .Z(n3311) );
  XOR U4231 ( .A(n3181), .B(n3180), .Z(n3305) );
  XOR U4232 ( .A(n3183), .B(n3182), .Z(n3295) );
  XOR U4233 ( .A(n3185), .B(n3184), .Z(n3291) );
  NAND U4234 ( .A(a[16]), .B(b[47]), .Z(n3274) );
  NAND U4235 ( .A(a[13]), .B(b[47]), .Z(n3257) );
  XOR U4236 ( .A(n3187), .B(n3186), .Z(n3256) );
  NANDN U4237 ( .A(n3257), .B(n3256), .Z(n3259) );
  XNOR U4238 ( .A(n3189), .B(n3188), .Z(n3252) );
  XNOR U4239 ( .A(n3191), .B(n3190), .Z(n3248) );
  XOR U4240 ( .A(n3193), .B(n3192), .Z(n3244) );
  XNOR U4241 ( .A(n3195), .B(n3194), .Z(n3235) );
  XOR U4242 ( .A(n3197), .B(n3196), .Z(n3199) );
  AND U4243 ( .A(a[7]), .B(b[47]), .Z(n3198) );
  NANDN U4244 ( .A(n3199), .B(n3198), .Z(n3233) );
  XOR U4245 ( .A(n3199), .B(n3198), .Z(n3740) );
  XNOR U4246 ( .A(n3201), .B(n3200), .Z(n3223) );
  XNOR U4247 ( .A(n3203), .B(n3202), .Z(n3218) );
  XNOR U4248 ( .A(n3205), .B(n3204), .Z(n3214) );
  NAND U4249 ( .A(b[48]), .B(a[1]), .Z(n3207) );
  NAND U4250 ( .A(n3207), .B(n3206), .Z(n3210) );
  OR U4251 ( .A(n3207), .B(n4012), .Z(n3755) );
  NANDN U4252 ( .A(n3209), .B(n3755), .Z(n3208) );
  AND U4253 ( .A(n3210), .B(n3208), .Z(n3213) );
  XNOR U4254 ( .A(n3755), .B(n3209), .Z(n3211) );
  NAND U4255 ( .A(n3211), .B(n3210), .Z(n3751) );
  ANDN U4256 ( .B(b[47]), .A(n162), .Z(n3750) );
  OR U4257 ( .A(n3751), .B(n3750), .Z(n3212) );
  AND U4258 ( .A(n3213), .B(n3212), .Z(n3215) );
  OR U4259 ( .A(n3214), .B(n3215), .Z(n3217) );
  XNOR U4260 ( .A(n3215), .B(n3214), .Z(n3748) );
  ANDN U4261 ( .B(b[47]), .A(n21580), .Z(n3749) );
  OR U4262 ( .A(n3748), .B(n3749), .Z(n3216) );
  AND U4263 ( .A(n3217), .B(n3216), .Z(n3219) );
  OR U4264 ( .A(n3218), .B(n3219), .Z(n3221) );
  XNOR U4265 ( .A(n3219), .B(n3218), .Z(n3746) );
  ANDN U4266 ( .B(b[47]), .A(n163), .Z(n3747) );
  OR U4267 ( .A(n3746), .B(n3747), .Z(n3220) );
  AND U4268 ( .A(n3221), .B(n3220), .Z(n3222) );
  OR U4269 ( .A(n3223), .B(n3222), .Z(n3225) );
  XNOR U4270 ( .A(n3223), .B(n3222), .Z(n3774) );
  NAND U4271 ( .A(b[47]), .B(a[5]), .Z(n3775) );
  NANDN U4272 ( .A(n3774), .B(n3775), .Z(n3224) );
  NAND U4273 ( .A(n3225), .B(n3224), .Z(n3227) );
  AND U4274 ( .A(a[6]), .B(b[47]), .Z(n3226) );
  NANDN U4275 ( .A(n3227), .B(n3226), .Z(n3231) );
  XOR U4276 ( .A(n3227), .B(n3226), .Z(n3742) );
  XOR U4277 ( .A(n3229), .B(n3228), .Z(n3743) );
  NANDN U4278 ( .A(n3742), .B(n3743), .Z(n3230) );
  AND U4279 ( .A(n3231), .B(n3230), .Z(n3741) );
  OR U4280 ( .A(n3740), .B(n3741), .Z(n3232) );
  AND U4281 ( .A(n3233), .B(n3232), .Z(n3234) );
  OR U4282 ( .A(n3235), .B(n3234), .Z(n3237) );
  XNOR U4283 ( .A(n3235), .B(n3234), .Z(n3785) );
  NAND U4284 ( .A(a[8]), .B(b[47]), .Z(n3784) );
  OR U4285 ( .A(n3785), .B(n3784), .Z(n3236) );
  NAND U4286 ( .A(n3237), .B(n3236), .Z(n3240) );
  XOR U4287 ( .A(n3239), .B(n3238), .Z(n3241) );
  OR U4288 ( .A(n3240), .B(n3241), .Z(n3243) );
  ANDN U4289 ( .B(b[47]), .A(n21615), .Z(n3739) );
  XOR U4290 ( .A(n3241), .B(n3240), .Z(n3738) );
  NANDN U4291 ( .A(n3739), .B(n3738), .Z(n3242) );
  AND U4292 ( .A(n3243), .B(n3242), .Z(n3245) );
  OR U4293 ( .A(n3244), .B(n3245), .Z(n3247) );
  XNOR U4294 ( .A(n3245), .B(n3244), .Z(n3736) );
  ANDN U4295 ( .B(b[47]), .A(n168), .Z(n3737) );
  OR U4296 ( .A(n3736), .B(n3737), .Z(n3246) );
  AND U4297 ( .A(n3247), .B(n3246), .Z(n3249) );
  OR U4298 ( .A(n3248), .B(n3249), .Z(n3251) );
  XNOR U4299 ( .A(n3249), .B(n3248), .Z(n3734) );
  ANDN U4300 ( .B(b[47]), .A(n21164), .Z(n3735) );
  OR U4301 ( .A(n3734), .B(n3735), .Z(n3250) );
  AND U4302 ( .A(n3251), .B(n3250), .Z(n3253) );
  OR U4303 ( .A(n3252), .B(n3253), .Z(n3255) );
  XNOR U4304 ( .A(n3253), .B(n3252), .Z(n3733) );
  ANDN U4305 ( .B(b[47]), .A(n169), .Z(n3732) );
  OR U4306 ( .A(n3733), .B(n3732), .Z(n3254) );
  NAND U4307 ( .A(n3255), .B(n3254), .Z(n3807) );
  NANDN U4308 ( .A(n3807), .B(n3806), .Z(n3258) );
  AND U4309 ( .A(n3259), .B(n3258), .Z(n3262) );
  NANDN U4310 ( .A(n3262), .B(n3263), .Z(n3265) );
  XOR U4311 ( .A(n3263), .B(n3262), .Z(n3813) );
  AND U4312 ( .A(a[14]), .B(b[47]), .Z(n3812) );
  NANDN U4313 ( .A(n3813), .B(n3812), .Z(n3264) );
  AND U4314 ( .A(n3265), .B(n3264), .Z(n3268) );
  XNOR U4315 ( .A(n3267), .B(n3266), .Z(n3269) );
  NANDN U4316 ( .A(n3268), .B(n3269), .Z(n3271) );
  XOR U4317 ( .A(n3269), .B(n3268), .Z(n3821) );
  AND U4318 ( .A(a[15]), .B(b[47]), .Z(n3820) );
  NANDN U4319 ( .A(n3821), .B(n3820), .Z(n3270) );
  AND U4320 ( .A(n3271), .B(n3270), .Z(n3275) );
  OR U4321 ( .A(n3274), .B(n3275), .Z(n3277) );
  XOR U4322 ( .A(n3273), .B(n3272), .Z(n3729) );
  XNOR U4323 ( .A(n3275), .B(n3274), .Z(n3728) );
  OR U4324 ( .A(n3729), .B(n3728), .Z(n3276) );
  AND U4325 ( .A(n3277), .B(n3276), .Z(n3280) );
  NANDN U4326 ( .A(n3280), .B(n3281), .Z(n3283) );
  XOR U4327 ( .A(n3281), .B(n3280), .Z(n3827) );
  AND U4328 ( .A(a[17]), .B(b[47]), .Z(n3826) );
  NANDN U4329 ( .A(n3827), .B(n3826), .Z(n3282) );
  NAND U4330 ( .A(n3283), .B(n3282), .Z(n3287) );
  XOR U4331 ( .A(n3285), .B(n3284), .Z(n3286) );
  NANDN U4332 ( .A(n3287), .B(n3286), .Z(n3289) );
  ANDN U4333 ( .B(b[47]), .A(n175), .Z(n3833) );
  XOR U4334 ( .A(n3287), .B(n3286), .Z(n3832) );
  OR U4335 ( .A(n3833), .B(n3832), .Z(n3288) );
  NAND U4336 ( .A(n3289), .B(n3288), .Z(n3290) );
  NANDN U4337 ( .A(n3291), .B(n3290), .Z(n3293) );
  ANDN U4338 ( .B(b[47]), .A(n21670), .Z(n3839) );
  NANDN U4339 ( .A(n3839), .B(n3838), .Z(n3292) );
  NAND U4340 ( .A(n3293), .B(n3292), .Z(n3294) );
  NANDN U4341 ( .A(n3295), .B(n3294), .Z(n3297) );
  ANDN U4342 ( .B(b[47]), .A(n176), .Z(n3725) );
  NANDN U4343 ( .A(n3725), .B(n3724), .Z(n3296) );
  NAND U4344 ( .A(n3297), .B(n3296), .Z(n3300) );
  NANDN U4345 ( .A(n3300), .B(n3301), .Z(n3303) );
  NAND U4346 ( .A(a[21]), .B(b[47]), .Z(n3721) );
  XNOR U4347 ( .A(n3301), .B(n3300), .Z(n3720) );
  NANDN U4348 ( .A(n3721), .B(n3720), .Z(n3302) );
  NAND U4349 ( .A(n3303), .B(n3302), .Z(n3304) );
  NANDN U4350 ( .A(n3305), .B(n3304), .Z(n3307) );
  XOR U4351 ( .A(n3305), .B(n3304), .Z(n3849) );
  NAND U4352 ( .A(b[47]), .B(a[22]), .Z(n3848) );
  OR U4353 ( .A(n3849), .B(n3848), .Z(n3306) );
  AND U4354 ( .A(n3307), .B(n3306), .Z(n3854) );
  XNOR U4355 ( .A(n3309), .B(n3308), .Z(n3855) );
  NANDN U4356 ( .A(n3854), .B(n3855), .Z(n3310) );
  AND U4357 ( .A(n3311), .B(n3310), .Z(n3718) );
  OR U4358 ( .A(n3719), .B(n3718), .Z(n3312) );
  NAND U4359 ( .A(n3313), .B(n3312), .Z(n3314) );
  NANDN U4360 ( .A(n3315), .B(n3314), .Z(n3319) );
  NAND U4361 ( .A(n3716), .B(n3717), .Z(n3318) );
  NAND U4362 ( .A(n3319), .B(n3318), .Z(n3323) );
  XOR U4363 ( .A(n3321), .B(n3320), .Z(n3322) );
  NANDN U4364 ( .A(n3323), .B(n3322), .Z(n3325) );
  ANDN U4365 ( .B(b[47]), .A(n179), .Z(n3869) );
  XOR U4366 ( .A(n3323), .B(n3322), .Z(n3868) );
  OR U4367 ( .A(n3869), .B(n3868), .Z(n3324) );
  NAND U4368 ( .A(n3325), .B(n3324), .Z(n3326) );
  NANDN U4369 ( .A(n3327), .B(n3326), .Z(n3329) );
  ANDN U4370 ( .B(b[47]), .A(n21716), .Z(n3715) );
  NANDN U4371 ( .A(n3715), .B(n3714), .Z(n3328) );
  NAND U4372 ( .A(n3329), .B(n3328), .Z(n3712) );
  XOR U4373 ( .A(n3331), .B(n3330), .Z(n3713) );
  NAND U4374 ( .A(n3712), .B(n3713), .Z(n3332) );
  NAND U4375 ( .A(n3333), .B(n3332), .Z(n3337) );
  XOR U4376 ( .A(n3335), .B(n3334), .Z(n3336) );
  NANDN U4377 ( .A(n3337), .B(n3336), .Z(n3339) );
  NAND U4378 ( .A(a[29]), .B(b[47]), .Z(n3709) );
  NANDN U4379 ( .A(n3709), .B(n3708), .Z(n3338) );
  NAND U4380 ( .A(n3339), .B(n3338), .Z(n3343) );
  XOR U4381 ( .A(n3341), .B(n3340), .Z(n3342) );
  NANDN U4382 ( .A(n3343), .B(n3342), .Z(n3345) );
  ANDN U4383 ( .B(b[47]), .A(n181), .Z(n3884) );
  OR U4384 ( .A(n3884), .B(n3885), .Z(n3344) );
  NAND U4385 ( .A(n3345), .B(n3344), .Z(n3707) );
  XOR U4386 ( .A(n3347), .B(n3346), .Z(n3706) );
  NANDN U4387 ( .A(n3707), .B(n3706), .Z(n3348) );
  NAND U4388 ( .A(n3349), .B(n3348), .Z(n3353) );
  XNOR U4389 ( .A(n3351), .B(n3350), .Z(n3352) );
  NANDN U4390 ( .A(n3353), .B(n3352), .Z(n3355) );
  ANDN U4391 ( .B(b[47]), .A(n182), .Z(n3705) );
  NANDN U4392 ( .A(n3705), .B(n3704), .Z(n3354) );
  NAND U4393 ( .A(n3355), .B(n3354), .Z(n3359) );
  XOR U4394 ( .A(n3357), .B(n3356), .Z(n3358) );
  NANDN U4395 ( .A(n3359), .B(n3358), .Z(n3361) );
  XOR U4396 ( .A(n3359), .B(n3358), .Z(n3703) );
  NAND U4397 ( .A(a[33]), .B(b[47]), .Z(n3702) );
  OR U4398 ( .A(n3703), .B(n3702), .Z(n3360) );
  AND U4399 ( .A(n3361), .B(n3360), .Z(n3700) );
  OR U4400 ( .A(n3701), .B(n3700), .Z(n3362) );
  AND U4401 ( .A(n3363), .B(n3362), .Z(n3367) );
  OR U4402 ( .A(n3367), .B(n3366), .Z(n3369) );
  NAND U4403 ( .A(a[35]), .B(b[47]), .Z(n3699) );
  XOR U4404 ( .A(n3367), .B(n3366), .Z(n3698) );
  NANDN U4405 ( .A(n3699), .B(n3698), .Z(n3368) );
  NAND U4406 ( .A(n3369), .B(n3368), .Z(n3911) );
  NAND U4407 ( .A(n3910), .B(n3911), .Z(n3370) );
  NAND U4408 ( .A(n3371), .B(n3370), .Z(n3374) );
  OR U4409 ( .A(n3374), .B(n3375), .Z(n3377) );
  ANDN U4410 ( .B(b[47]), .A(n21772), .Z(n3697) );
  XOR U4411 ( .A(n3375), .B(n3374), .Z(n3696) );
  NANDN U4412 ( .A(n3697), .B(n3696), .Z(n3376) );
  NAND U4413 ( .A(n3377), .B(n3376), .Z(n3381) );
  XOR U4414 ( .A(n3379), .B(n3378), .Z(n3380) );
  NANDN U4415 ( .A(n3381), .B(n3380), .Z(n3383) );
  NAND U4416 ( .A(a[38]), .B(b[47]), .Z(n3695) );
  NANDN U4417 ( .A(n3695), .B(n3694), .Z(n3382) );
  AND U4418 ( .A(n3383), .B(n3382), .Z(n3692) );
  NANDN U4419 ( .A(n3692), .B(n3693), .Z(n3386) );
  NAND U4420 ( .A(n3387), .B(n3386), .Z(n3390) );
  OR U4421 ( .A(n3390), .B(n3391), .Z(n3393) );
  ANDN U4422 ( .B(b[47]), .A(n188), .Z(n3691) );
  XOR U4423 ( .A(n3391), .B(n3390), .Z(n3690) );
  NANDN U4424 ( .A(n3691), .B(n3690), .Z(n3392) );
  AND U4425 ( .A(n3393), .B(n3392), .Z(n3395) );
  OR U4426 ( .A(n3394), .B(n3395), .Z(n3397) );
  XNOR U4427 ( .A(n3395), .B(n3394), .Z(n3688) );
  ANDN U4428 ( .B(b[47]), .A(n189), .Z(n3689) );
  OR U4429 ( .A(n3688), .B(n3689), .Z(n3396) );
  AND U4430 ( .A(n3397), .B(n3396), .Z(n3399) );
  OR U4431 ( .A(n3398), .B(n3399), .Z(n3401) );
  XNOR U4432 ( .A(n3399), .B(n3398), .Z(n3686) );
  NAND U4433 ( .A(b[47]), .B(a[42]), .Z(n3687) );
  NANDN U4434 ( .A(n3686), .B(n3687), .Z(n3400) );
  AND U4435 ( .A(n3401), .B(n3400), .Z(n3403) );
  OR U4436 ( .A(n3402), .B(n3403), .Z(n3405) );
  XNOR U4437 ( .A(n3403), .B(n3402), .Z(n3941) );
  ANDN U4438 ( .B(b[47]), .A(n191), .Z(n3940) );
  OR U4439 ( .A(n3941), .B(n3940), .Z(n3404) );
  AND U4440 ( .A(n3405), .B(n3404), .Z(n3497) );
  NAND U4441 ( .A(a[42]), .B(b[49]), .Z(n3503) );
  OR U4442 ( .A(n3407), .B(n3406), .Z(n3411) );
  OR U4443 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U4444 ( .A(n3411), .B(n3410), .Z(n3500) );
  ANDN U4445 ( .B(b[51]), .A(n188), .Z(n3509) );
  OR U4446 ( .A(n3413), .B(n3412), .Z(n3417) );
  OR U4447 ( .A(n3415), .B(n3414), .Z(n3416) );
  NAND U4448 ( .A(n3417), .B(n3416), .Z(n3507) );
  NAND U4449 ( .A(a[38]), .B(b[53]), .Z(n3515) );
  OR U4450 ( .A(n3419), .B(n3418), .Z(n3423) );
  NANDN U4451 ( .A(n3421), .B(n3420), .Z(n3422) );
  AND U4452 ( .A(n3423), .B(n3422), .Z(n3512) );
  NAND U4453 ( .A(a[36]), .B(b[55]), .Z(n3521) );
  OR U4454 ( .A(n3425), .B(n3424), .Z(n3429) );
  NANDN U4455 ( .A(n3427), .B(n3426), .Z(n3428) );
  NAND U4456 ( .A(n3429), .B(n3428), .Z(n3519) );
  NAND U4457 ( .A(a[34]), .B(b[57]), .Z(n3527) );
  OR U4458 ( .A(n3431), .B(n3430), .Z(n3435) );
  OR U4459 ( .A(n3433), .B(n3432), .Z(n3434) );
  AND U4460 ( .A(n3435), .B(n3434), .Z(n3524) );
  NAND U4461 ( .A(a[32]), .B(b[59]), .Z(n3533) );
  OR U4462 ( .A(n3437), .B(n3436), .Z(n3441) );
  OR U4463 ( .A(n3439), .B(n3438), .Z(n3440) );
  NAND U4464 ( .A(n3441), .B(n3440), .Z(n3531) );
  ANDN U4465 ( .B(b[61]), .A(n181), .Z(n3538) );
  OR U4466 ( .A(n3443), .B(n3442), .Z(n3447) );
  NANDN U4467 ( .A(n3445), .B(n3444), .Z(n3446) );
  AND U4468 ( .A(n3447), .B(n3446), .Z(n3536) );
  ANDN U4469 ( .B(b[63]), .A(n180), .Z(n3544) );
  ANDN U4470 ( .B(a[29]), .A(n159), .Z(n3542) );
  OR U4471 ( .A(n3449), .B(n3448), .Z(n3453) );
  OR U4472 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U4473 ( .A(n3453), .B(n3452), .Z(n3543) );
  XNOR U4474 ( .A(n3542), .B(n3543), .Z(n3545) );
  XNOR U4475 ( .A(n3544), .B(n3545), .Z(n3537) );
  XNOR U4476 ( .A(n3536), .B(n3537), .Z(n3539) );
  XNOR U4477 ( .A(n3538), .B(n3539), .Z(n3551) );
  ANDN U4478 ( .B(b[60]), .A(n21740), .Z(n3548) );
  OR U4479 ( .A(n3455), .B(n3454), .Z(n3459) );
  NANDN U4480 ( .A(n3457), .B(n3456), .Z(n3458) );
  NAND U4481 ( .A(n3459), .B(n3458), .Z(n3549) );
  XNOR U4482 ( .A(n3548), .B(n3549), .Z(n3550) );
  XOR U4483 ( .A(n3551), .B(n3550), .Z(n3530) );
  XOR U4484 ( .A(n3531), .B(n3530), .Z(n3532) );
  ANDN U4485 ( .B(b[58]), .A(n21751), .Z(n3554) );
  OR U4486 ( .A(n3461), .B(n3460), .Z(n3465) );
  OR U4487 ( .A(n3463), .B(n3462), .Z(n3464) );
  AND U4488 ( .A(n3465), .B(n3464), .Z(n3555) );
  XOR U4489 ( .A(n3554), .B(n3555), .Z(n3556) );
  XNOR U4490 ( .A(n3557), .B(n3556), .Z(n3525) );
  XNOR U4491 ( .A(n3524), .B(n3525), .Z(n3526) );
  XOR U4492 ( .A(n3527), .B(n3526), .Z(n3563) );
  ANDN U4493 ( .B(b[56]), .A(n184), .Z(n3560) );
  OR U4494 ( .A(n3467), .B(n3466), .Z(n3471) );
  NANDN U4495 ( .A(n3469), .B(n3468), .Z(n3470) );
  NAND U4496 ( .A(n3471), .B(n3470), .Z(n3561) );
  XOR U4497 ( .A(n3560), .B(n3561), .Z(n3562) );
  XNOR U4498 ( .A(n3563), .B(n3562), .Z(n3518) );
  XNOR U4499 ( .A(n3519), .B(n3518), .Z(n3520) );
  XOR U4500 ( .A(n3521), .B(n3520), .Z(n3569) );
  ANDN U4501 ( .B(b[54]), .A(n21772), .Z(n3566) );
  OR U4502 ( .A(n3473), .B(n3472), .Z(n3477) );
  OR U4503 ( .A(n3475), .B(n3474), .Z(n3476) );
  AND U4504 ( .A(n3477), .B(n3476), .Z(n3567) );
  XOR U4505 ( .A(n3566), .B(n3567), .Z(n3568) );
  XNOR U4506 ( .A(n3569), .B(n3568), .Z(n3513) );
  XNOR U4507 ( .A(n3512), .B(n3513), .Z(n3514) );
  XOR U4508 ( .A(n3515), .B(n3514), .Z(n3574) );
  ANDN U4509 ( .B(b[52]), .A(n187), .Z(n3572) );
  OR U4510 ( .A(n3479), .B(n3478), .Z(n3483) );
  NANDN U4511 ( .A(n3481), .B(n3480), .Z(n3482) );
  AND U4512 ( .A(n3483), .B(n3482), .Z(n3573) );
  XNOR U4513 ( .A(n3572), .B(n3573), .Z(n3575) );
  XOR U4514 ( .A(n3574), .B(n3575), .Z(n3506) );
  XOR U4515 ( .A(n3509), .B(n3508), .Z(n3581) );
  ANDN U4516 ( .B(b[50]), .A(n189), .Z(n3578) );
  OR U4517 ( .A(n3485), .B(n3484), .Z(n3489) );
  NANDN U4518 ( .A(n3487), .B(n3486), .Z(n3488) );
  AND U4519 ( .A(n3489), .B(n3488), .Z(n3579) );
  XNOR U4520 ( .A(n3578), .B(n3579), .Z(n3580) );
  XOR U4521 ( .A(n3581), .B(n3580), .Z(n3501) );
  XNOR U4522 ( .A(n3500), .B(n3501), .Z(n3502) );
  XOR U4523 ( .A(n3503), .B(n3502), .Z(n3586) );
  ANDN U4524 ( .B(b[48]), .A(n191), .Z(n3584) );
  NANDN U4525 ( .A(n3491), .B(n3490), .Z(n3495) );
  OR U4526 ( .A(n3493), .B(n3492), .Z(n3494) );
  NAND U4527 ( .A(n3495), .B(n3494), .Z(n3585) );
  XNOR U4528 ( .A(n3584), .B(n3585), .Z(n3587) );
  XOR U4529 ( .A(n3586), .B(n3587), .Z(n3496) );
  NANDN U4530 ( .A(n3497), .B(n3496), .Z(n3499) );
  NAND U4531 ( .A(b[47]), .B(a[44]), .Z(n3947) );
  NAND U4532 ( .A(n3946), .B(n3947), .Z(n3498) );
  AND U4533 ( .A(n3499), .B(n3498), .Z(n3591) );
  ANDN U4534 ( .B(b[49]), .A(n191), .Z(n3597) );
  OR U4535 ( .A(n3501), .B(n3500), .Z(n3505) );
  OR U4536 ( .A(n3503), .B(n3502), .Z(n3504) );
  NAND U4537 ( .A(n3505), .B(n3504), .Z(n3595) );
  ANDN U4538 ( .B(b[51]), .A(n189), .Z(n3602) );
  NANDN U4539 ( .A(n3507), .B(n3506), .Z(n3511) );
  NANDN U4540 ( .A(n3509), .B(n3508), .Z(n3510) );
  AND U4541 ( .A(n3511), .B(n3510), .Z(n3601) );
  ANDN U4542 ( .B(b[53]), .A(n187), .Z(n3609) );
  OR U4543 ( .A(n3513), .B(n3512), .Z(n3517) );
  OR U4544 ( .A(n3515), .B(n3514), .Z(n3516) );
  NAND U4545 ( .A(n3517), .B(n3516), .Z(n3607) );
  NAND U4546 ( .A(a[37]), .B(b[55]), .Z(n3615) );
  OR U4547 ( .A(n3519), .B(n3518), .Z(n3523) );
  OR U4548 ( .A(n3521), .B(n3520), .Z(n3522) );
  AND U4549 ( .A(n3523), .B(n3522), .Z(n3612) );
  NAND U4550 ( .A(a[35]), .B(b[57]), .Z(n3621) );
  OR U4551 ( .A(n3525), .B(n3524), .Z(n3529) );
  OR U4552 ( .A(n3527), .B(n3526), .Z(n3528) );
  AND U4553 ( .A(n3529), .B(n3528), .Z(n3618) );
  ANDN U4554 ( .B(b[59]), .A(n21751), .Z(n3627) );
  OR U4555 ( .A(n3531), .B(n3530), .Z(n3535) );
  NANDN U4556 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U4557 ( .A(n3535), .B(n3534), .Z(n3625) );
  ANDN U4558 ( .B(b[61]), .A(n21740), .Z(n3632) );
  OR U4559 ( .A(n3537), .B(n3536), .Z(n3541) );
  OR U4560 ( .A(n3539), .B(n3538), .Z(n3540) );
  AND U4561 ( .A(n3541), .B(n3540), .Z(n3630) );
  ANDN U4562 ( .B(b[63]), .A(n21727), .Z(n3638) );
  ANDN U4563 ( .B(a[30]), .A(n159), .Z(n3636) );
  OR U4564 ( .A(n3543), .B(n3542), .Z(n3547) );
  OR U4565 ( .A(n3545), .B(n3544), .Z(n3546) );
  AND U4566 ( .A(n3547), .B(n3546), .Z(n3637) );
  XNOR U4567 ( .A(n3636), .B(n3637), .Z(n3639) );
  XNOR U4568 ( .A(n3638), .B(n3639), .Z(n3631) );
  XNOR U4569 ( .A(n3630), .B(n3631), .Z(n3633) );
  XNOR U4570 ( .A(n3632), .B(n3633), .Z(n3645) );
  ANDN U4571 ( .B(b[60]), .A(n182), .Z(n3642) );
  OR U4572 ( .A(n3549), .B(n3548), .Z(n3553) );
  OR U4573 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U4574 ( .A(n3553), .B(n3552), .Z(n3643) );
  XOR U4575 ( .A(n3642), .B(n3643), .Z(n3644) );
  XOR U4576 ( .A(n3627), .B(n3626), .Z(n3651) );
  ANDN U4577 ( .B(b[58]), .A(n183), .Z(n3648) );
  OR U4578 ( .A(n3555), .B(n3554), .Z(n3559) );
  NANDN U4579 ( .A(n3557), .B(n3556), .Z(n3558) );
  AND U4580 ( .A(n3559), .B(n3558), .Z(n3649) );
  XNOR U4581 ( .A(n3648), .B(n3649), .Z(n3650) );
  XOR U4582 ( .A(n3651), .B(n3650), .Z(n3619) );
  XNOR U4583 ( .A(n3618), .B(n3619), .Z(n3620) );
  XOR U4584 ( .A(n3621), .B(n3620), .Z(n3657) );
  ANDN U4585 ( .B(b[56]), .A(n185), .Z(n3654) );
  OR U4586 ( .A(n3561), .B(n3560), .Z(n3565) );
  NANDN U4587 ( .A(n3563), .B(n3562), .Z(n3564) );
  AND U4588 ( .A(n3565), .B(n3564), .Z(n3655) );
  XOR U4589 ( .A(n3654), .B(n3655), .Z(n3656) );
  XNOR U4590 ( .A(n3657), .B(n3656), .Z(n3613) );
  XNOR U4591 ( .A(n3612), .B(n3613), .Z(n3614) );
  XOR U4592 ( .A(n3615), .B(n3614), .Z(n3662) );
  ANDN U4593 ( .B(b[54]), .A(n186), .Z(n3660) );
  OR U4594 ( .A(n3567), .B(n3566), .Z(n3571) );
  NANDN U4595 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U4596 ( .A(n3571), .B(n3570), .Z(n3661) );
  XNOR U4597 ( .A(n3660), .B(n3661), .Z(n3663) );
  XOR U4598 ( .A(n3662), .B(n3663), .Z(n3606) );
  XOR U4599 ( .A(n3609), .B(n3608), .Z(n3669) );
  ANDN U4600 ( .B(b[52]), .A(n188), .Z(n3666) );
  OR U4601 ( .A(n3573), .B(n3572), .Z(n3577) );
  OR U4602 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U4603 ( .A(n3577), .B(n3576), .Z(n3667) );
  XOR U4604 ( .A(n3666), .B(n3667), .Z(n3668) );
  XOR U4605 ( .A(n3601), .B(n3600), .Z(n3603) );
  XNOR U4606 ( .A(n3602), .B(n3603), .Z(n3675) );
  ANDN U4607 ( .B(b[50]), .A(n190), .Z(n3672) );
  OR U4608 ( .A(n3579), .B(n3578), .Z(n3583) );
  OR U4609 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U4610 ( .A(n3583), .B(n3582), .Z(n3673) );
  XOR U4611 ( .A(n3672), .B(n3673), .Z(n3674) );
  XOR U4612 ( .A(n3597), .B(n3596), .Z(n3681) );
  ANDN U4613 ( .B(b[48]), .A(n192), .Z(n3678) );
  OR U4614 ( .A(n3585), .B(n3584), .Z(n3589) );
  OR U4615 ( .A(n3587), .B(n3586), .Z(n3588) );
  AND U4616 ( .A(n3589), .B(n3588), .Z(n3679) );
  XOR U4617 ( .A(n3678), .B(n3679), .Z(n3680) );
  NANDN U4618 ( .A(n3591), .B(n3590), .Z(n3593) );
  XOR U4619 ( .A(n3591), .B(n3590), .Z(n3684) );
  ANDN U4620 ( .B(b[47]), .A(n193), .Z(n3685) );
  OR U4621 ( .A(n3684), .B(n3685), .Z(n3592) );
  AND U4622 ( .A(n3593), .B(n3592), .Z(n4819) );
  ANDN U4623 ( .B(b[49]), .A(n192), .Z(n4826) );
  NANDN U4624 ( .A(n3595), .B(n3594), .Z(n3599) );
  NANDN U4625 ( .A(n3597), .B(n3596), .Z(n3598) );
  AND U4626 ( .A(n3599), .B(n3598), .Z(n4825) );
  NAND U4627 ( .A(a[42]), .B(b[51]), .Z(n4905) );
  NANDN U4628 ( .A(n3601), .B(n3600), .Z(n3605) );
  OR U4629 ( .A(n3603), .B(n3602), .Z(n3604) );
  NAND U4630 ( .A(n3605), .B(n3604), .Z(n4903) );
  ANDN U4631 ( .B(b[53]), .A(n188), .Z(n4844) );
  NANDN U4632 ( .A(n3607), .B(n3606), .Z(n3611) );
  NANDN U4633 ( .A(n3609), .B(n3608), .Z(n3610) );
  AND U4634 ( .A(n3611), .B(n3610), .Z(n4843) );
  NAND U4635 ( .A(a[38]), .B(b[55]), .Z(n4851) );
  OR U4636 ( .A(n3613), .B(n3612), .Z(n3617) );
  OR U4637 ( .A(n3615), .B(n3614), .Z(n3616) );
  AND U4638 ( .A(n3617), .B(n3616), .Z(n4848) );
  NAND U4639 ( .A(a[36]), .B(b[57]), .Z(n4893) );
  OR U4640 ( .A(n3619), .B(n3618), .Z(n3623) );
  OR U4641 ( .A(n3621), .B(n3620), .Z(n3622) );
  AND U4642 ( .A(n3623), .B(n3622), .Z(n4890) );
  NAND U4643 ( .A(a[34]), .B(b[59]), .Z(n4863) );
  NANDN U4644 ( .A(n3625), .B(n3624), .Z(n3629) );
  NANDN U4645 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U4646 ( .A(n3629), .B(n3628), .Z(n4861) );
  ANDN U4647 ( .B(b[61]), .A(n182), .Z(n4868) );
  OR U4648 ( .A(n3631), .B(n3630), .Z(n3635) );
  OR U4649 ( .A(n3633), .B(n3632), .Z(n3634) );
  AND U4650 ( .A(n3635), .B(n3634), .Z(n4866) );
  ANDN U4651 ( .B(b[63]), .A(n181), .Z(n4874) );
  ANDN U4652 ( .B(a[31]), .A(n159), .Z(n4872) );
  OR U4653 ( .A(n3637), .B(n3636), .Z(n3641) );
  OR U4654 ( .A(n3639), .B(n3638), .Z(n3640) );
  AND U4655 ( .A(n3641), .B(n3640), .Z(n4873) );
  XNOR U4656 ( .A(n4872), .B(n4873), .Z(n4875) );
  XNOR U4657 ( .A(n4874), .B(n4875), .Z(n4867) );
  XNOR U4658 ( .A(n4866), .B(n4867), .Z(n4869) );
  XNOR U4659 ( .A(n4868), .B(n4869), .Z(n4881) );
  ANDN U4660 ( .B(b[60]), .A(n21751), .Z(n4878) );
  OR U4661 ( .A(n3643), .B(n3642), .Z(n3647) );
  NANDN U4662 ( .A(n3645), .B(n3644), .Z(n3646) );
  AND U4663 ( .A(n3647), .B(n3646), .Z(n4879) );
  XNOR U4664 ( .A(n4878), .B(n4879), .Z(n4880) );
  XOR U4665 ( .A(n4881), .B(n4880), .Z(n4860) );
  XOR U4666 ( .A(n4861), .B(n4860), .Z(n4862) );
  ANDN U4667 ( .B(b[58]), .A(n184), .Z(n4884) );
  OR U4668 ( .A(n3649), .B(n3648), .Z(n3653) );
  OR U4669 ( .A(n3651), .B(n3650), .Z(n3652) );
  AND U4670 ( .A(n3653), .B(n3652), .Z(n4885) );
  XOR U4671 ( .A(n4884), .B(n4885), .Z(n4886) );
  XNOR U4672 ( .A(n4887), .B(n4886), .Z(n4891) );
  XNOR U4673 ( .A(n4890), .B(n4891), .Z(n4892) );
  XOR U4674 ( .A(n4893), .B(n4892), .Z(n4857) );
  ANDN U4675 ( .B(b[56]), .A(n21772), .Z(n4854) );
  OR U4676 ( .A(n3655), .B(n3654), .Z(n3659) );
  NANDN U4677 ( .A(n3657), .B(n3656), .Z(n3658) );
  AND U4678 ( .A(n3659), .B(n3658), .Z(n4855) );
  XOR U4679 ( .A(n4854), .B(n4855), .Z(n4856) );
  XNOR U4680 ( .A(n4857), .B(n4856), .Z(n4849) );
  XNOR U4681 ( .A(n4848), .B(n4849), .Z(n4850) );
  XOR U4682 ( .A(n4851), .B(n4850), .Z(n4898) );
  ANDN U4683 ( .B(b[54]), .A(n187), .Z(n4896) );
  OR U4684 ( .A(n3661), .B(n3660), .Z(n3665) );
  OR U4685 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U4686 ( .A(n3665), .B(n3664), .Z(n4897) );
  XNOR U4687 ( .A(n4896), .B(n4897), .Z(n4899) );
  XOR U4688 ( .A(n4898), .B(n4899), .Z(n4842) );
  XOR U4689 ( .A(n4843), .B(n4842), .Z(n4845) );
  XNOR U4690 ( .A(n4844), .B(n4845), .Z(n4839) );
  ANDN U4691 ( .B(b[52]), .A(n189), .Z(n4836) );
  OR U4692 ( .A(n3667), .B(n3666), .Z(n3671) );
  NANDN U4693 ( .A(n3669), .B(n3668), .Z(n3670) );
  AND U4694 ( .A(n3671), .B(n3670), .Z(n4837) );
  XNOR U4695 ( .A(n4836), .B(n4837), .Z(n4838) );
  XOR U4696 ( .A(n4839), .B(n4838), .Z(n4902) );
  XOR U4697 ( .A(n4903), .B(n4902), .Z(n4904) );
  ANDN U4698 ( .B(b[50]), .A(n191), .Z(n4830) );
  OR U4699 ( .A(n3673), .B(n3672), .Z(n3677) );
  NANDN U4700 ( .A(n3675), .B(n3674), .Z(n3676) );
  AND U4701 ( .A(n3677), .B(n3676), .Z(n4831) );
  XNOR U4702 ( .A(n4830), .B(n4831), .Z(n4833) );
  XOR U4703 ( .A(n4832), .B(n4833), .Z(n4824) );
  XOR U4704 ( .A(n4825), .B(n4824), .Z(n4827) );
  XNOR U4705 ( .A(n4826), .B(n4827), .Z(n4911) );
  ANDN U4706 ( .B(b[48]), .A(n193), .Z(n4908) );
  OR U4707 ( .A(n3679), .B(n3678), .Z(n3683) );
  NANDN U4708 ( .A(n3681), .B(n3680), .Z(n3682) );
  AND U4709 ( .A(n3683), .B(n3682), .Z(n4909) );
  XOR U4710 ( .A(n4908), .B(n4909), .Z(n4910) );
  XOR U4711 ( .A(n4819), .B(n4818), .Z(n4821) );
  XNOR U4712 ( .A(n4820), .B(n4821), .Z(n4917) );
  ANDN U4713 ( .B(b[46]), .A(n195), .Z(n4914) );
  XNOR U4714 ( .A(n3685), .B(n3684), .Z(n3953) );
  NAND U4715 ( .A(a[43]), .B(b[46]), .Z(n3937) );
  XOR U4716 ( .A(n3687), .B(n3686), .Z(n3936) );
  NANDN U4717 ( .A(n3937), .B(n3936), .Z(n3939) );
  XNOR U4718 ( .A(n3689), .B(n3688), .Z(n3932) );
  XOR U4719 ( .A(n3691), .B(n3690), .Z(n3928) );
  XNOR U4720 ( .A(n3693), .B(n3692), .Z(n3924) );
  XNOR U4721 ( .A(n3695), .B(n3694), .Z(n3920) );
  XOR U4722 ( .A(n3697), .B(n3696), .Z(n3916) );
  NAND U4723 ( .A(a[36]), .B(b[46]), .Z(n3907) );
  XNOR U4724 ( .A(n3699), .B(n3698), .Z(n3906) );
  NANDN U4725 ( .A(n3907), .B(n3906), .Z(n3909) );
  NAND U4726 ( .A(a[35]), .B(b[46]), .Z(n3903) );
  XOR U4727 ( .A(n3701), .B(n3700), .Z(n3902) );
  NANDN U4728 ( .A(n3903), .B(n3902), .Z(n3905) );
  XOR U4729 ( .A(n3703), .B(n3702), .Z(n3899) );
  XOR U4730 ( .A(n3705), .B(n3704), .Z(n3895) );
  XNOR U4731 ( .A(n3707), .B(n3706), .Z(n3891) );
  NAND U4732 ( .A(b[46]), .B(a[30]), .Z(n3710) );
  XNOR U4733 ( .A(n3709), .B(n3708), .Z(n3711) );
  NANDN U4734 ( .A(n3710), .B(n3711), .Z(n3883) );
  XOR U4735 ( .A(n3711), .B(n3710), .Z(n4147) );
  ANDN U4736 ( .B(b[46]), .A(n21727), .Z(n3879) );
  XNOR U4737 ( .A(n3713), .B(n3712), .Z(n3878) );
  OR U4738 ( .A(n3879), .B(n3878), .Z(n3881) );
  NAND U4739 ( .A(a[28]), .B(b[46]), .Z(n3875) );
  NANDN U4740 ( .A(n3875), .B(n3874), .Z(n3877) );
  NAND U4741 ( .A(b[46]), .B(a[26]), .Z(n3864) );
  NANDN U4742 ( .A(n3864), .B(n3865), .Z(n3867) );
  XOR U4743 ( .A(n3719), .B(n3718), .Z(n3861) );
  NAND U4744 ( .A(a[22]), .B(b[46]), .Z(n3723) );
  XNOR U4745 ( .A(n3721), .B(n3720), .Z(n3722) );
  NANDN U4746 ( .A(n3723), .B(n3722), .Z(n3847) );
  XOR U4747 ( .A(n3723), .B(n3722), .Z(n4109) );
  NAND U4748 ( .A(a[21]), .B(b[46]), .Z(n3726) );
  NANDN U4749 ( .A(n3726), .B(n3727), .Z(n3845) );
  XOR U4750 ( .A(n3727), .B(n3726), .Z(n4105) );
  XNOR U4751 ( .A(n3729), .B(n3728), .Z(n3731) );
  AND U4752 ( .A(a[17]), .B(b[46]), .Z(n3730) );
  NANDN U4753 ( .A(n3731), .B(n3730), .Z(n3825) );
  XOR U4754 ( .A(n3731), .B(n3730), .Z(n3986) );
  NAND U4755 ( .A(a[16]), .B(b[46]), .Z(n3818) );
  NAND U4756 ( .A(a[13]), .B(b[46]), .Z(n3802) );
  XOR U4757 ( .A(n3733), .B(n3732), .Z(n3803) );
  OR U4758 ( .A(n3802), .B(n3803), .Z(n3805) );
  XNOR U4759 ( .A(n3735), .B(n3734), .Z(n3798) );
  XNOR U4760 ( .A(n3737), .B(n3736), .Z(n3794) );
  XOR U4761 ( .A(n3739), .B(n3738), .Z(n3790) );
  XNOR U4762 ( .A(n3741), .B(n3740), .Z(n3781) );
  XOR U4763 ( .A(n3743), .B(n3742), .Z(n3745) );
  AND U4764 ( .A(a[7]), .B(b[46]), .Z(n3744) );
  NANDN U4765 ( .A(n3745), .B(n3744), .Z(n3779) );
  XOR U4766 ( .A(n3745), .B(n3744), .Z(n4000) );
  XNOR U4767 ( .A(n3747), .B(n3746), .Z(n3769) );
  XNOR U4768 ( .A(n3749), .B(n3748), .Z(n3764) );
  XNOR U4769 ( .A(n3751), .B(n3750), .Z(n3760) );
  NAND U4770 ( .A(b[47]), .B(a[1]), .Z(n3753) );
  NAND U4771 ( .A(n3753), .B(n3752), .Z(n3756) );
  OR U4772 ( .A(n3753), .B(n4320), .Z(n4015) );
  NANDN U4773 ( .A(n3755), .B(n4015), .Z(n3754) );
  AND U4774 ( .A(n3756), .B(n3754), .Z(n3759) );
  XNOR U4775 ( .A(n4015), .B(n3755), .Z(n3757) );
  NAND U4776 ( .A(n3757), .B(n3756), .Z(n4011) );
  ANDN U4777 ( .B(b[46]), .A(n162), .Z(n4010) );
  OR U4778 ( .A(n4011), .B(n4010), .Z(n3758) );
  AND U4779 ( .A(n3759), .B(n3758), .Z(n3761) );
  OR U4780 ( .A(n3760), .B(n3761), .Z(n3763) );
  XNOR U4781 ( .A(n3761), .B(n3760), .Z(n4008) );
  ANDN U4782 ( .B(b[46]), .A(n21580), .Z(n4009) );
  OR U4783 ( .A(n4008), .B(n4009), .Z(n3762) );
  AND U4784 ( .A(n3763), .B(n3762), .Z(n3765) );
  OR U4785 ( .A(n3764), .B(n3765), .Z(n3767) );
  XNOR U4786 ( .A(n3765), .B(n3764), .Z(n4006) );
  ANDN U4787 ( .B(b[46]), .A(n163), .Z(n4007) );
  OR U4788 ( .A(n4006), .B(n4007), .Z(n3766) );
  AND U4789 ( .A(n3767), .B(n3766), .Z(n3768) );
  OR U4790 ( .A(n3769), .B(n3768), .Z(n3771) );
  XNOR U4791 ( .A(n3769), .B(n3768), .Z(n4034) );
  NAND U4792 ( .A(b[46]), .B(a[5]), .Z(n4035) );
  NANDN U4793 ( .A(n4034), .B(n4035), .Z(n3770) );
  NAND U4794 ( .A(n3771), .B(n3770), .Z(n3773) );
  AND U4795 ( .A(a[6]), .B(b[46]), .Z(n3772) );
  NANDN U4796 ( .A(n3773), .B(n3772), .Z(n3777) );
  XOR U4797 ( .A(n3773), .B(n3772), .Z(n4002) );
  XOR U4798 ( .A(n3775), .B(n3774), .Z(n4003) );
  NANDN U4799 ( .A(n4002), .B(n4003), .Z(n3776) );
  AND U4800 ( .A(n3777), .B(n3776), .Z(n4001) );
  OR U4801 ( .A(n4000), .B(n4001), .Z(n3778) );
  AND U4802 ( .A(n3779), .B(n3778), .Z(n3780) );
  OR U4803 ( .A(n3781), .B(n3780), .Z(n3783) );
  XNOR U4804 ( .A(n3781), .B(n3780), .Z(n4045) );
  NAND U4805 ( .A(a[8]), .B(b[46]), .Z(n4044) );
  OR U4806 ( .A(n4045), .B(n4044), .Z(n3782) );
  NAND U4807 ( .A(n3783), .B(n3782), .Z(n3786) );
  XOR U4808 ( .A(n3785), .B(n3784), .Z(n3787) );
  OR U4809 ( .A(n3786), .B(n3787), .Z(n3789) );
  ANDN U4810 ( .B(b[46]), .A(n21615), .Z(n3999) );
  XOR U4811 ( .A(n3787), .B(n3786), .Z(n3998) );
  NANDN U4812 ( .A(n3999), .B(n3998), .Z(n3788) );
  AND U4813 ( .A(n3789), .B(n3788), .Z(n3791) );
  OR U4814 ( .A(n3790), .B(n3791), .Z(n3793) );
  XNOR U4815 ( .A(n3791), .B(n3790), .Z(n3996) );
  ANDN U4816 ( .B(b[46]), .A(n168), .Z(n3997) );
  OR U4817 ( .A(n3996), .B(n3997), .Z(n3792) );
  AND U4818 ( .A(n3793), .B(n3792), .Z(n3795) );
  OR U4819 ( .A(n3794), .B(n3795), .Z(n3797) );
  XNOR U4820 ( .A(n3795), .B(n3794), .Z(n3994) );
  ANDN U4821 ( .B(b[46]), .A(n21164), .Z(n3995) );
  OR U4822 ( .A(n3994), .B(n3995), .Z(n3796) );
  AND U4823 ( .A(n3797), .B(n3796), .Z(n3799) );
  OR U4824 ( .A(n3798), .B(n3799), .Z(n3801) );
  XNOR U4825 ( .A(n3799), .B(n3798), .Z(n3993) );
  ANDN U4826 ( .B(b[46]), .A(n169), .Z(n3992) );
  OR U4827 ( .A(n3993), .B(n3992), .Z(n3800) );
  NAND U4828 ( .A(n3801), .B(n3800), .Z(n4067) );
  XOR U4829 ( .A(n3803), .B(n3802), .Z(n4066) );
  NANDN U4830 ( .A(n4067), .B(n4066), .Z(n3804) );
  AND U4831 ( .A(n3805), .B(n3804), .Z(n3808) );
  NANDN U4832 ( .A(n3808), .B(n3809), .Z(n3811) );
  XOR U4833 ( .A(n3809), .B(n3808), .Z(n4073) );
  AND U4834 ( .A(a[14]), .B(b[46]), .Z(n4072) );
  NANDN U4835 ( .A(n4073), .B(n4072), .Z(n3810) );
  AND U4836 ( .A(n3811), .B(n3810), .Z(n3815) );
  XNOR U4837 ( .A(n3813), .B(n3812), .Z(n3814) );
  NANDN U4838 ( .A(n3815), .B(n3814), .Z(n3817) );
  NAND U4839 ( .A(a[15]), .B(b[46]), .Z(n4081) );
  NANDN U4840 ( .A(n4081), .B(n4080), .Z(n3816) );
  AND U4841 ( .A(n3817), .B(n3816), .Z(n3819) );
  OR U4842 ( .A(n3818), .B(n3819), .Z(n3823) );
  XNOR U4843 ( .A(n3819), .B(n3818), .Z(n3989) );
  XNOR U4844 ( .A(n3821), .B(n3820), .Z(n3988) );
  NANDN U4845 ( .A(n3989), .B(n3988), .Z(n3822) );
  AND U4846 ( .A(n3823), .B(n3822), .Z(n3987) );
  OR U4847 ( .A(n3986), .B(n3987), .Z(n3824) );
  AND U4848 ( .A(n3825), .B(n3824), .Z(n3828) );
  XNOR U4849 ( .A(n3827), .B(n3826), .Z(n3829) );
  NANDN U4850 ( .A(n3828), .B(n3829), .Z(n3831) );
  XOR U4851 ( .A(n3829), .B(n3828), .Z(n4091) );
  NAND U4852 ( .A(a[18]), .B(b[46]), .Z(n4090) );
  OR U4853 ( .A(n4091), .B(n4090), .Z(n3830) );
  NAND U4854 ( .A(n3831), .B(n3830), .Z(n3835) );
  XOR U4855 ( .A(n3833), .B(n3832), .Z(n3834) );
  NANDN U4856 ( .A(n3835), .B(n3834), .Z(n3837) );
  ANDN U4857 ( .B(b[46]), .A(n21670), .Z(n3983) );
  XOR U4858 ( .A(n3835), .B(n3834), .Z(n3982) );
  OR U4859 ( .A(n3983), .B(n3982), .Z(n3836) );
  NAND U4860 ( .A(n3837), .B(n3836), .Z(n3841) );
  NANDN U4861 ( .A(n3841), .B(n3840), .Z(n3843) );
  XOR U4862 ( .A(n3841), .B(n3840), .Z(n3980) );
  NAND U4863 ( .A(a[20]), .B(b[46]), .Z(n3981) );
  OR U4864 ( .A(n3980), .B(n3981), .Z(n3842) );
  NAND U4865 ( .A(n3843), .B(n3842), .Z(n4104) );
  NANDN U4866 ( .A(n4105), .B(n4104), .Z(n3844) );
  NAND U4867 ( .A(n3845), .B(n3844), .Z(n4108) );
  NANDN U4868 ( .A(n4109), .B(n4108), .Z(n3846) );
  NAND U4869 ( .A(n3847), .B(n3846), .Z(n3850) );
  XOR U4870 ( .A(n3849), .B(n3848), .Z(n3851) );
  NAND U4871 ( .A(n3850), .B(n3851), .Z(n3853) );
  XNOR U4872 ( .A(n3851), .B(n3850), .Z(n3979) );
  NAND U4873 ( .A(a[23]), .B(b[46]), .Z(n3978) );
  OR U4874 ( .A(n3979), .B(n3978), .Z(n3852) );
  NAND U4875 ( .A(n3853), .B(n3852), .Z(n3857) );
  XOR U4876 ( .A(n3855), .B(n3854), .Z(n3856) );
  NANDN U4877 ( .A(n3857), .B(n3856), .Z(n3859) );
  ANDN U4878 ( .B(b[46]), .A(n178), .Z(n3977) );
  NANDN U4879 ( .A(n3977), .B(n3976), .Z(n3858) );
  NAND U4880 ( .A(n3859), .B(n3858), .Z(n3860) );
  NANDN U4881 ( .A(n3861), .B(n3860), .Z(n3863) );
  ANDN U4882 ( .B(b[46]), .A(n21703), .Z(n3975) );
  NANDN U4883 ( .A(n3975), .B(n3974), .Z(n3862) );
  NAND U4884 ( .A(n3863), .B(n3862), .Z(n4127) );
  XNOR U4885 ( .A(n3865), .B(n3864), .Z(n4126) );
  NANDN U4886 ( .A(n4127), .B(n4126), .Z(n3866) );
  NAND U4887 ( .A(n3867), .B(n3866), .Z(n3871) );
  XOR U4888 ( .A(n3869), .B(n3868), .Z(n3870) );
  NANDN U4889 ( .A(n3871), .B(n3870), .Z(n3873) );
  ANDN U4890 ( .B(b[46]), .A(n21716), .Z(n3973) );
  XOR U4891 ( .A(n3871), .B(n3870), .Z(n3972) );
  OR U4892 ( .A(n3973), .B(n3972), .Z(n3872) );
  NAND U4893 ( .A(n3873), .B(n3872), .Z(n4137) );
  XNOR U4894 ( .A(n3875), .B(n3874), .Z(n4136) );
  NANDN U4895 ( .A(n4137), .B(n4136), .Z(n3876) );
  AND U4896 ( .A(n3877), .B(n3876), .Z(n3970) );
  XOR U4897 ( .A(n3879), .B(n3878), .Z(n3971) );
  NAND U4898 ( .A(n3970), .B(n3971), .Z(n3880) );
  NAND U4899 ( .A(n3881), .B(n3880), .Z(n4146) );
  OR U4900 ( .A(n4147), .B(n4146), .Z(n3882) );
  NAND U4901 ( .A(n3883), .B(n3882), .Z(n3887) );
  XOR U4902 ( .A(n3885), .B(n3884), .Z(n3886) );
  NANDN U4903 ( .A(n3887), .B(n3886), .Z(n3889) );
  ANDN U4904 ( .B(b[46]), .A(n21740), .Z(n3969) );
  XOR U4905 ( .A(n3887), .B(n3886), .Z(n3968) );
  OR U4906 ( .A(n3969), .B(n3968), .Z(n3888) );
  NAND U4907 ( .A(n3889), .B(n3888), .Z(n3890) );
  NANDN U4908 ( .A(n3891), .B(n3890), .Z(n3893) );
  ANDN U4909 ( .B(b[46]), .A(n182), .Z(n3967) );
  NANDN U4910 ( .A(n3967), .B(n3966), .Z(n3892) );
  NAND U4911 ( .A(n3893), .B(n3892), .Z(n3894) );
  NANDN U4912 ( .A(n3895), .B(n3894), .Z(n3897) );
  ANDN U4913 ( .B(b[46]), .A(n21751), .Z(n3965) );
  NANDN U4914 ( .A(n3965), .B(n3964), .Z(n3896) );
  NAND U4915 ( .A(n3897), .B(n3896), .Z(n3898) );
  NANDN U4916 ( .A(n3899), .B(n3898), .Z(n3901) );
  ANDN U4917 ( .B(b[46]), .A(n183), .Z(n4165) );
  NANDN U4918 ( .A(n4165), .B(n4164), .Z(n3900) );
  NAND U4919 ( .A(n3901), .B(n3900), .Z(n3963) );
  XNOR U4920 ( .A(n3903), .B(n3902), .Z(n3962) );
  NANDN U4921 ( .A(n3963), .B(n3962), .Z(n3904) );
  AND U4922 ( .A(n3905), .B(n3904), .Z(n4174) );
  XNOR U4923 ( .A(n3907), .B(n3906), .Z(n4175) );
  NANDN U4924 ( .A(n4174), .B(n4175), .Z(n3908) );
  NAND U4925 ( .A(n3909), .B(n3908), .Z(n3912) );
  OR U4926 ( .A(n3912), .B(n3913), .Z(n3915) );
  ANDN U4927 ( .B(b[46]), .A(n21772), .Z(n3961) );
  XOR U4928 ( .A(n3913), .B(n3912), .Z(n3960) );
  NANDN U4929 ( .A(n3961), .B(n3960), .Z(n3914) );
  AND U4930 ( .A(n3915), .B(n3914), .Z(n3917) );
  OR U4931 ( .A(n3916), .B(n3917), .Z(n3919) );
  XNOR U4932 ( .A(n3917), .B(n3916), .Z(n3958) );
  ANDN U4933 ( .B(b[46]), .A(n186), .Z(n3959) );
  OR U4934 ( .A(n3958), .B(n3959), .Z(n3918) );
  AND U4935 ( .A(n3919), .B(n3918), .Z(n3921) );
  OR U4936 ( .A(n3920), .B(n3921), .Z(n3923) );
  XNOR U4937 ( .A(n3921), .B(n3920), .Z(n4188) );
  NAND U4938 ( .A(b[46]), .B(a[39]), .Z(n4189) );
  NANDN U4939 ( .A(n4188), .B(n4189), .Z(n3922) );
  AND U4940 ( .A(n3923), .B(n3922), .Z(n3925) );
  OR U4941 ( .A(n3924), .B(n3925), .Z(n3927) );
  XNOR U4942 ( .A(n3925), .B(n3924), .Z(n4194) );
  ANDN U4943 ( .B(b[46]), .A(n188), .Z(n4195) );
  OR U4944 ( .A(n4194), .B(n4195), .Z(n3926) );
  AND U4945 ( .A(n3927), .B(n3926), .Z(n3929) );
  OR U4946 ( .A(n3928), .B(n3929), .Z(n3931) );
  XNOR U4947 ( .A(n3929), .B(n3928), .Z(n4200) );
  NAND U4948 ( .A(b[46]), .B(a[41]), .Z(n4201) );
  NANDN U4949 ( .A(n4200), .B(n4201), .Z(n3930) );
  AND U4950 ( .A(n3931), .B(n3930), .Z(n3933) );
  OR U4951 ( .A(n3932), .B(n3933), .Z(n3935) );
  XNOR U4952 ( .A(n3933), .B(n3932), .Z(n4206) );
  ANDN U4953 ( .B(b[46]), .A(n190), .Z(n4207) );
  OR U4954 ( .A(n4206), .B(n4207), .Z(n3934) );
  NAND U4955 ( .A(n3935), .B(n3934), .Z(n3957) );
  NANDN U4956 ( .A(n3957), .B(n3956), .Z(n3938) );
  NAND U4957 ( .A(n3939), .B(n3938), .Z(n3943) );
  XOR U4958 ( .A(n3941), .B(n3940), .Z(n3942) );
  NANDN U4959 ( .A(n3943), .B(n3942), .Z(n3945) );
  NAND U4960 ( .A(b[46]), .B(a[44]), .Z(n4217) );
  NAND U4961 ( .A(n4216), .B(n4217), .Z(n3944) );
  NAND U4962 ( .A(n3945), .B(n3944), .Z(n3949) );
  NANDN U4963 ( .A(n3949), .B(n3948), .Z(n3951) );
  NAND U4964 ( .A(a[45]), .B(b[46]), .Z(n4223) );
  NANDN U4965 ( .A(n4223), .B(n4222), .Z(n3950) );
  NAND U4966 ( .A(n3951), .B(n3950), .Z(n3952) );
  OR U4967 ( .A(n3953), .B(n3952), .Z(n3955) );
  XNOR U4968 ( .A(n3953), .B(n3952), .Z(n4228) );
  NAND U4969 ( .A(b[46]), .B(a[46]), .Z(n4229) );
  NANDN U4970 ( .A(n4228), .B(n4229), .Z(n3954) );
  AND U4971 ( .A(n3955), .B(n3954), .Z(n4915) );
  XOR U4972 ( .A(n4914), .B(n4915), .Z(n4916) );
  XNOR U4973 ( .A(n3957), .B(n3956), .Z(n4212) );
  XNOR U4974 ( .A(n3959), .B(n3958), .Z(n4184) );
  XOR U4975 ( .A(n3961), .B(n3960), .Z(n4181) );
  XOR U4976 ( .A(n3963), .B(n3962), .Z(n4171) );
  XOR U4977 ( .A(n3965), .B(n3964), .Z(n4161) );
  XOR U4978 ( .A(n3967), .B(n3966), .Z(n4157) );
  ANDN U4979 ( .B(b[45]), .A(n182), .Z(n4152) );
  XNOR U4980 ( .A(n3969), .B(n3968), .Z(n4153) );
  OR U4981 ( .A(n4152), .B(n4153), .Z(n4155) );
  XNOR U4982 ( .A(n3971), .B(n3970), .Z(n4143) );
  XOR U4983 ( .A(n3973), .B(n3972), .Z(n4133) );
  XOR U4984 ( .A(n3975), .B(n3974), .Z(n4123) );
  XOR U4985 ( .A(n3977), .B(n3976), .Z(n4119) );
  XOR U4986 ( .A(n3979), .B(n3978), .Z(n4115) );
  ANDN U4987 ( .B(b[45]), .A(n177), .Z(n4103) );
  ANDN U4988 ( .B(b[45]), .A(n21681), .Z(n4099) );
  XOR U4989 ( .A(n3981), .B(n3980), .Z(n4098) );
  OR U4990 ( .A(n4099), .B(n4098), .Z(n4101) );
  NAND U4991 ( .A(a[20]), .B(b[45]), .Z(n3984) );
  XNOR U4992 ( .A(n3983), .B(n3982), .Z(n3985) );
  NANDN U4993 ( .A(n3984), .B(n3985), .Z(n4097) );
  XOR U4994 ( .A(n3985), .B(n3984), .Z(n4291) );
  XNOR U4995 ( .A(n3987), .B(n3986), .Z(n4087) );
  AND U4996 ( .A(a[17]), .B(b[45]), .Z(n3990) );
  NANDN U4997 ( .A(n3991), .B(n3990), .Z(n4085) );
  XOR U4998 ( .A(n3991), .B(n3990), .Z(n4294) );
  NAND U4999 ( .A(a[16]), .B(b[45]), .Z(n4078) );
  NAND U5000 ( .A(a[13]), .B(b[45]), .Z(n4062) );
  XOR U5001 ( .A(n3993), .B(n3992), .Z(n4063) );
  OR U5002 ( .A(n4062), .B(n4063), .Z(n4065) );
  XNOR U5003 ( .A(n3995), .B(n3994), .Z(n4058) );
  XNOR U5004 ( .A(n3997), .B(n3996), .Z(n4054) );
  XOR U5005 ( .A(n3999), .B(n3998), .Z(n4050) );
  XNOR U5006 ( .A(n4001), .B(n4000), .Z(n4041) );
  XOR U5007 ( .A(n4003), .B(n4002), .Z(n4005) );
  AND U5008 ( .A(a[7]), .B(b[45]), .Z(n4004) );
  NANDN U5009 ( .A(n4005), .B(n4004), .Z(n4039) );
  XOR U5010 ( .A(n4005), .B(n4004), .Z(n4308) );
  XNOR U5011 ( .A(n4007), .B(n4006), .Z(n4029) );
  XNOR U5012 ( .A(n4009), .B(n4008), .Z(n4024) );
  XNOR U5013 ( .A(n4011), .B(n4010), .Z(n4020) );
  NAND U5014 ( .A(b[46]), .B(a[1]), .Z(n4013) );
  NAND U5015 ( .A(n4013), .B(n4012), .Z(n4016) );
  OR U5016 ( .A(n4013), .B(n4580), .Z(n4323) );
  NANDN U5017 ( .A(n4015), .B(n4323), .Z(n4014) );
  AND U5018 ( .A(n4016), .B(n4014), .Z(n4019) );
  XNOR U5019 ( .A(n4323), .B(n4015), .Z(n4017) );
  NAND U5020 ( .A(n4017), .B(n4016), .Z(n4319) );
  ANDN U5021 ( .B(b[45]), .A(n162), .Z(n4318) );
  OR U5022 ( .A(n4319), .B(n4318), .Z(n4018) );
  AND U5023 ( .A(n4019), .B(n4018), .Z(n4021) );
  OR U5024 ( .A(n4020), .B(n4021), .Z(n4023) );
  XNOR U5025 ( .A(n4021), .B(n4020), .Z(n4316) );
  ANDN U5026 ( .B(b[45]), .A(n21580), .Z(n4317) );
  OR U5027 ( .A(n4316), .B(n4317), .Z(n4022) );
  AND U5028 ( .A(n4023), .B(n4022), .Z(n4025) );
  OR U5029 ( .A(n4024), .B(n4025), .Z(n4027) );
  XNOR U5030 ( .A(n4025), .B(n4024), .Z(n4314) );
  ANDN U5031 ( .B(b[45]), .A(n163), .Z(n4315) );
  OR U5032 ( .A(n4314), .B(n4315), .Z(n4026) );
  AND U5033 ( .A(n4027), .B(n4026), .Z(n4028) );
  OR U5034 ( .A(n4029), .B(n4028), .Z(n4031) );
  XNOR U5035 ( .A(n4029), .B(n4028), .Z(n4342) );
  NAND U5036 ( .A(b[45]), .B(a[5]), .Z(n4343) );
  NANDN U5037 ( .A(n4342), .B(n4343), .Z(n4030) );
  NAND U5038 ( .A(n4031), .B(n4030), .Z(n4033) );
  AND U5039 ( .A(a[6]), .B(b[45]), .Z(n4032) );
  NANDN U5040 ( .A(n4033), .B(n4032), .Z(n4037) );
  XOR U5041 ( .A(n4033), .B(n4032), .Z(n4310) );
  XOR U5042 ( .A(n4035), .B(n4034), .Z(n4311) );
  NANDN U5043 ( .A(n4310), .B(n4311), .Z(n4036) );
  AND U5044 ( .A(n4037), .B(n4036), .Z(n4309) );
  OR U5045 ( .A(n4308), .B(n4309), .Z(n4038) );
  AND U5046 ( .A(n4039), .B(n4038), .Z(n4040) );
  OR U5047 ( .A(n4041), .B(n4040), .Z(n4043) );
  XNOR U5048 ( .A(n4041), .B(n4040), .Z(n4353) );
  NAND U5049 ( .A(a[8]), .B(b[45]), .Z(n4352) );
  OR U5050 ( .A(n4353), .B(n4352), .Z(n4042) );
  NAND U5051 ( .A(n4043), .B(n4042), .Z(n4046) );
  XOR U5052 ( .A(n4045), .B(n4044), .Z(n4047) );
  OR U5053 ( .A(n4046), .B(n4047), .Z(n4049) );
  ANDN U5054 ( .B(b[45]), .A(n21615), .Z(n4307) );
  XOR U5055 ( .A(n4047), .B(n4046), .Z(n4306) );
  NANDN U5056 ( .A(n4307), .B(n4306), .Z(n4048) );
  AND U5057 ( .A(n4049), .B(n4048), .Z(n4051) );
  OR U5058 ( .A(n4050), .B(n4051), .Z(n4053) );
  XNOR U5059 ( .A(n4051), .B(n4050), .Z(n4304) );
  ANDN U5060 ( .B(b[45]), .A(n168), .Z(n4305) );
  OR U5061 ( .A(n4304), .B(n4305), .Z(n4052) );
  AND U5062 ( .A(n4053), .B(n4052), .Z(n4055) );
  OR U5063 ( .A(n4054), .B(n4055), .Z(n4057) );
  XNOR U5064 ( .A(n4055), .B(n4054), .Z(n4302) );
  ANDN U5065 ( .B(b[45]), .A(n21164), .Z(n4303) );
  OR U5066 ( .A(n4302), .B(n4303), .Z(n4056) );
  AND U5067 ( .A(n4057), .B(n4056), .Z(n4059) );
  OR U5068 ( .A(n4058), .B(n4059), .Z(n4061) );
  XNOR U5069 ( .A(n4059), .B(n4058), .Z(n4301) );
  ANDN U5070 ( .B(b[45]), .A(n169), .Z(n4300) );
  OR U5071 ( .A(n4301), .B(n4300), .Z(n4060) );
  NAND U5072 ( .A(n4061), .B(n4060), .Z(n4375) );
  XOR U5073 ( .A(n4063), .B(n4062), .Z(n4374) );
  NANDN U5074 ( .A(n4375), .B(n4374), .Z(n4064) );
  AND U5075 ( .A(n4065), .B(n4064), .Z(n4068) );
  NANDN U5076 ( .A(n4068), .B(n4069), .Z(n4071) );
  XOR U5077 ( .A(n4069), .B(n4068), .Z(n4381) );
  AND U5078 ( .A(a[14]), .B(b[45]), .Z(n4380) );
  NANDN U5079 ( .A(n4381), .B(n4380), .Z(n4070) );
  AND U5080 ( .A(n4071), .B(n4070), .Z(n4074) );
  XNOR U5081 ( .A(n4073), .B(n4072), .Z(n4075) );
  NANDN U5082 ( .A(n4074), .B(n4075), .Z(n4077) );
  XOR U5083 ( .A(n4075), .B(n4074), .Z(n4389) );
  AND U5084 ( .A(a[15]), .B(b[45]), .Z(n4388) );
  NANDN U5085 ( .A(n4389), .B(n4388), .Z(n4076) );
  AND U5086 ( .A(n4077), .B(n4076), .Z(n4079) );
  OR U5087 ( .A(n4078), .B(n4079), .Z(n4083) );
  XNOR U5088 ( .A(n4079), .B(n4078), .Z(n4297) );
  NANDN U5089 ( .A(n4297), .B(n4296), .Z(n4082) );
  AND U5090 ( .A(n4083), .B(n4082), .Z(n4295) );
  OR U5091 ( .A(n4294), .B(n4295), .Z(n4084) );
  AND U5092 ( .A(n4085), .B(n4084), .Z(n4086) );
  OR U5093 ( .A(n4087), .B(n4086), .Z(n4089) );
  XNOR U5094 ( .A(n4087), .B(n4086), .Z(n4399) );
  AND U5095 ( .A(a[18]), .B(b[45]), .Z(n4398) );
  NANDN U5096 ( .A(n4399), .B(n4398), .Z(n4088) );
  NAND U5097 ( .A(n4089), .B(n4088), .Z(n4092) );
  XOR U5098 ( .A(n4091), .B(n4090), .Z(n4093) );
  OR U5099 ( .A(n4092), .B(n4093), .Z(n4095) );
  XOR U5100 ( .A(n4093), .B(n4092), .Z(n4406) );
  NAND U5101 ( .A(b[45]), .B(a[19]), .Z(n4407) );
  NAND U5102 ( .A(n4406), .B(n4407), .Z(n4094) );
  NAND U5103 ( .A(n4095), .B(n4094), .Z(n4290) );
  OR U5104 ( .A(n4291), .B(n4290), .Z(n4096) );
  NAND U5105 ( .A(n4097), .B(n4096), .Z(n4413) );
  XOR U5106 ( .A(n4099), .B(n4098), .Z(n4412) );
  NANDN U5107 ( .A(n4413), .B(n4412), .Z(n4100) );
  NAND U5108 ( .A(n4101), .B(n4100), .Z(n4102) );
  NANDN U5109 ( .A(n4103), .B(n4102), .Z(n4107) );
  NANDN U5110 ( .A(n4288), .B(n4289), .Z(n4106) );
  AND U5111 ( .A(n4107), .B(n4106), .Z(n4110) );
  NANDN U5112 ( .A(n4110), .B(n4111), .Z(n4113) );
  ANDN U5113 ( .B(b[45]), .A(n21692), .Z(n4423) );
  XOR U5114 ( .A(n4111), .B(n4110), .Z(n4422) );
  OR U5115 ( .A(n4423), .B(n4422), .Z(n4112) );
  NAND U5116 ( .A(n4113), .B(n4112), .Z(n4114) );
  NANDN U5117 ( .A(n4115), .B(n4114), .Z(n4117) );
  ANDN U5118 ( .B(b[45]), .A(n178), .Z(n4285) );
  NANDN U5119 ( .A(n4285), .B(n4284), .Z(n4116) );
  NAND U5120 ( .A(n4117), .B(n4116), .Z(n4118) );
  NANDN U5121 ( .A(n4119), .B(n4118), .Z(n4121) );
  ANDN U5122 ( .B(b[45]), .A(n21703), .Z(n4283) );
  NANDN U5123 ( .A(n4283), .B(n4282), .Z(n4120) );
  NAND U5124 ( .A(n4121), .B(n4120), .Z(n4122) );
  NANDN U5125 ( .A(n4123), .B(n4122), .Z(n4125) );
  ANDN U5126 ( .B(b[45]), .A(n179), .Z(n4281) );
  NANDN U5127 ( .A(n4281), .B(n4280), .Z(n4124) );
  NAND U5128 ( .A(n4125), .B(n4124), .Z(n4129) );
  XNOR U5129 ( .A(n4127), .B(n4126), .Z(n4128) );
  NANDN U5130 ( .A(n4129), .B(n4128), .Z(n4131) );
  NAND U5131 ( .A(a[27]), .B(b[45]), .Z(n4277) );
  XNOR U5132 ( .A(n4129), .B(n4128), .Z(n4276) );
  NANDN U5133 ( .A(n4277), .B(n4276), .Z(n4130) );
  NAND U5134 ( .A(n4131), .B(n4130), .Z(n4132) );
  NANDN U5135 ( .A(n4133), .B(n4132), .Z(n4135) );
  NAND U5136 ( .A(a[28]), .B(b[45]), .Z(n4275) );
  NANDN U5137 ( .A(n4275), .B(n4274), .Z(n4134) );
  NAND U5138 ( .A(n4135), .B(n4134), .Z(n4139) );
  XOR U5139 ( .A(n4137), .B(n4136), .Z(n4138) );
  NANDN U5140 ( .A(n4139), .B(n4138), .Z(n4141) );
  ANDN U5141 ( .B(b[45]), .A(n21727), .Z(n4445) );
  OR U5142 ( .A(n4445), .B(n4444), .Z(n4140) );
  NAND U5143 ( .A(n4141), .B(n4140), .Z(n4142) );
  NANDN U5144 ( .A(n4143), .B(n4142), .Z(n4145) );
  ANDN U5145 ( .B(b[45]), .A(n181), .Z(n4273) );
  NANDN U5146 ( .A(n4273), .B(n4272), .Z(n4144) );
  NAND U5147 ( .A(n4145), .B(n4144), .Z(n4149) );
  XOR U5148 ( .A(n4147), .B(n4146), .Z(n4148) );
  NANDN U5149 ( .A(n4149), .B(n4148), .Z(n4151) );
  NAND U5150 ( .A(a[31]), .B(b[45]), .Z(n4269) );
  XNOR U5151 ( .A(n4149), .B(n4148), .Z(n4268) );
  NANDN U5152 ( .A(n4269), .B(n4268), .Z(n4150) );
  AND U5153 ( .A(n4151), .B(n4150), .Z(n4266) );
  XOR U5154 ( .A(n4153), .B(n4152), .Z(n4267) );
  NAND U5155 ( .A(n4266), .B(n4267), .Z(n4154) );
  NAND U5156 ( .A(n4155), .B(n4154), .Z(n4156) );
  NANDN U5157 ( .A(n4157), .B(n4156), .Z(n4159) );
  ANDN U5158 ( .B(b[45]), .A(n21751), .Z(n4265) );
  NANDN U5159 ( .A(n4265), .B(n4264), .Z(n4158) );
  NAND U5160 ( .A(n4159), .B(n4158), .Z(n4160) );
  NANDN U5161 ( .A(n4161), .B(n4160), .Z(n4163) );
  ANDN U5162 ( .B(b[45]), .A(n183), .Z(n4263) );
  NANDN U5163 ( .A(n4263), .B(n4262), .Z(n4162) );
  NAND U5164 ( .A(n4163), .B(n4162), .Z(n4167) );
  NANDN U5165 ( .A(n4167), .B(n4166), .Z(n4169) );
  NAND U5166 ( .A(a[35]), .B(b[45]), .Z(n4259) );
  XNOR U5167 ( .A(n4167), .B(n4166), .Z(n4258) );
  NANDN U5168 ( .A(n4259), .B(n4258), .Z(n4168) );
  NAND U5169 ( .A(n4169), .B(n4168), .Z(n4170) );
  NANDN U5170 ( .A(n4171), .B(n4170), .Z(n4173) );
  XOR U5171 ( .A(n4171), .B(n4170), .Z(n4255) );
  NAND U5172 ( .A(b[45]), .B(a[36]), .Z(n4254) );
  OR U5173 ( .A(n4255), .B(n4254), .Z(n4172) );
  NAND U5174 ( .A(n4173), .B(n4172), .Z(n4177) );
  XOR U5175 ( .A(n4175), .B(n4174), .Z(n4176) );
  NANDN U5176 ( .A(n4177), .B(n4176), .Z(n4179) );
  ANDN U5177 ( .B(b[45]), .A(n21772), .Z(n4251) );
  NANDN U5178 ( .A(n4251), .B(n4250), .Z(n4178) );
  NAND U5179 ( .A(n4179), .B(n4178), .Z(n4180) );
  NANDN U5180 ( .A(n4181), .B(n4180), .Z(n4183) );
  ANDN U5181 ( .B(b[45]), .A(n186), .Z(n4249) );
  NANDN U5182 ( .A(n4249), .B(n4248), .Z(n4182) );
  AND U5183 ( .A(n4183), .B(n4182), .Z(n4185) );
  OR U5184 ( .A(n4184), .B(n4185), .Z(n4187) );
  XNOR U5185 ( .A(n4185), .B(n4184), .Z(n4246) );
  ANDN U5186 ( .B(b[45]), .A(n187), .Z(n4247) );
  OR U5187 ( .A(n4246), .B(n4247), .Z(n4186) );
  NAND U5188 ( .A(n4187), .B(n4186), .Z(n4191) );
  XOR U5189 ( .A(n4189), .B(n4188), .Z(n4190) );
  NANDN U5190 ( .A(n4191), .B(n4190), .Z(n4193) );
  NAND U5191 ( .A(a[40]), .B(b[45]), .Z(n4244) );
  NANDN U5192 ( .A(n4244), .B(n4245), .Z(n4192) );
  NAND U5193 ( .A(n4193), .B(n4192), .Z(n4197) );
  XOR U5194 ( .A(n4195), .B(n4194), .Z(n4196) );
  NANDN U5195 ( .A(n4197), .B(n4196), .Z(n4199) );
  ANDN U5196 ( .B(b[45]), .A(n189), .Z(n4243) );
  NANDN U5197 ( .A(n4243), .B(n4242), .Z(n4198) );
  NAND U5198 ( .A(n4199), .B(n4198), .Z(n4203) );
  XOR U5199 ( .A(n4201), .B(n4200), .Z(n4202) );
  NANDN U5200 ( .A(n4203), .B(n4202), .Z(n4205) );
  AND U5201 ( .A(a[42]), .B(b[45]), .Z(n4240) );
  NANDN U5202 ( .A(n4241), .B(n4240), .Z(n4204) );
  NAND U5203 ( .A(n4205), .B(n4204), .Z(n4209) );
  XOR U5204 ( .A(n4207), .B(n4206), .Z(n4208) );
  NANDN U5205 ( .A(n4209), .B(n4208), .Z(n4211) );
  ANDN U5206 ( .B(b[45]), .A(n191), .Z(n4495) );
  NANDN U5207 ( .A(n4495), .B(n4494), .Z(n4210) );
  AND U5208 ( .A(n4211), .B(n4210), .Z(n4213) );
  OR U5209 ( .A(n4212), .B(n4213), .Z(n4215) );
  XNOR U5210 ( .A(n4213), .B(n4212), .Z(n4238) );
  ANDN U5211 ( .B(b[45]), .A(n192), .Z(n4239) );
  OR U5212 ( .A(n4238), .B(n4239), .Z(n4214) );
  NAND U5213 ( .A(n4215), .B(n4214), .Z(n4219) );
  NANDN U5214 ( .A(n4219), .B(n4218), .Z(n4221) );
  NAND U5215 ( .A(a[45]), .B(b[45]), .Z(n4237) );
  NANDN U5216 ( .A(n4237), .B(n4236), .Z(n4220) );
  NAND U5217 ( .A(n4221), .B(n4220), .Z(n4224) );
  OR U5218 ( .A(n4224), .B(n4225), .Z(n4227) );
  ANDN U5219 ( .B(b[45]), .A(n194), .Z(n4235) );
  XOR U5220 ( .A(n4225), .B(n4224), .Z(n4234) );
  NANDN U5221 ( .A(n4235), .B(n4234), .Z(n4226) );
  NAND U5222 ( .A(n4227), .B(n4226), .Z(n4231) );
  XOR U5223 ( .A(n4229), .B(n4228), .Z(n4230) );
  NANDN U5224 ( .A(n4231), .B(n4230), .Z(n4233) );
  NAND U5225 ( .A(a[47]), .B(b[45]), .Z(n4513) );
  NANDN U5226 ( .A(n4513), .B(n4512), .Z(n4232) );
  NAND U5227 ( .A(n4233), .B(n4232), .Z(n4921) );
  XOR U5228 ( .A(n4235), .B(n4234), .Z(n4508) );
  XNOR U5229 ( .A(n4237), .B(n4236), .Z(n4504) );
  XNOR U5230 ( .A(n4239), .B(n4238), .Z(n4500) );
  XOR U5231 ( .A(n4241), .B(n4240), .Z(n4491) );
  AND U5232 ( .A(a[43]), .B(b[44]), .Z(n4490) );
  NANDN U5233 ( .A(n4491), .B(n4490), .Z(n4493) );
  XOR U5234 ( .A(n4243), .B(n4242), .Z(n4486) );
  XNOR U5235 ( .A(n4245), .B(n4244), .Z(n4482) );
  XNOR U5236 ( .A(n4247), .B(n4246), .Z(n4479) );
  ANDN U5237 ( .B(b[44]), .A(n187), .Z(n4474) );
  XOR U5238 ( .A(n4249), .B(n4248), .Z(n4475) );
  OR U5239 ( .A(n4474), .B(n4475), .Z(n4477) );
  NAND U5240 ( .A(a[38]), .B(b[44]), .Z(n4252) );
  NANDN U5241 ( .A(n4252), .B(n4253), .Z(n4473) );
  XOR U5242 ( .A(n4253), .B(n4252), .Z(n4532) );
  NAND U5243 ( .A(a[37]), .B(b[44]), .Z(n4257) );
  XOR U5244 ( .A(n4255), .B(n4254), .Z(n4256) );
  NANDN U5245 ( .A(n4257), .B(n4256), .Z(n4471) );
  XOR U5246 ( .A(n4257), .B(n4256), .Z(n4753) );
  ANDN U5247 ( .B(b[44]), .A(n185), .Z(n4260) );
  XOR U5248 ( .A(n4259), .B(n4258), .Z(n4261) );
  NANDN U5249 ( .A(n4260), .B(n4261), .Z(n4469) );
  XOR U5250 ( .A(n4261), .B(n4260), .Z(n4747) );
  ANDN U5251 ( .B(b[44]), .A(n184), .Z(n4465) );
  XOR U5252 ( .A(n4263), .B(n4262), .Z(n4464) );
  OR U5253 ( .A(n4465), .B(n4464), .Z(n4467) );
  XOR U5254 ( .A(n4265), .B(n4264), .Z(n4461) );
  XNOR U5255 ( .A(n4267), .B(n4266), .Z(n4457) );
  ANDN U5256 ( .B(b[44]), .A(n182), .Z(n4271) );
  XOR U5257 ( .A(n4269), .B(n4268), .Z(n4270) );
  NANDN U5258 ( .A(n4271), .B(n4270), .Z(n4455) );
  XOR U5259 ( .A(n4273), .B(n4272), .Z(n4451) );
  NAND U5260 ( .A(a[29]), .B(b[44]), .Z(n4441) );
  XNOR U5261 ( .A(n4275), .B(n4274), .Z(n4440) );
  NANDN U5262 ( .A(n4441), .B(n4440), .Z(n4443) );
  NAND U5263 ( .A(a[28]), .B(b[44]), .Z(n4279) );
  XNOR U5264 ( .A(n4277), .B(n4276), .Z(n4278) );
  NANDN U5265 ( .A(n4279), .B(n4278), .Z(n4439) );
  XOR U5266 ( .A(n4279), .B(n4278), .Z(n4543) );
  XNOR U5267 ( .A(n4281), .B(n4280), .Z(n4435) );
  XNOR U5268 ( .A(n4283), .B(n4282), .Z(n4431) );
  NAND U5269 ( .A(a[25]), .B(b[44]), .Z(n4287) );
  NANDN U5270 ( .A(n4287), .B(n4286), .Z(n4429) );
  XOR U5271 ( .A(n4287), .B(n4286), .Z(n4547) );
  NAND U5272 ( .A(a[23]), .B(b[44]), .Z(n4418) );
  XNOR U5273 ( .A(n4289), .B(n4288), .Z(n4419) );
  OR U5274 ( .A(n4418), .B(n4419), .Z(n4421) );
  NAND U5275 ( .A(a[21]), .B(b[44]), .Z(n4293) );
  XOR U5276 ( .A(n4291), .B(n4290), .Z(n4292) );
  NANDN U5277 ( .A(n4293), .B(n4292), .Z(n4411) );
  XOR U5278 ( .A(n4293), .B(n4292), .Z(n4675) );
  NAND U5279 ( .A(a[20]), .B(b[44]), .Z(n4404) );
  XNOR U5280 ( .A(n4295), .B(n4294), .Z(n4395) );
  AND U5281 ( .A(a[17]), .B(b[44]), .Z(n4298) );
  NANDN U5282 ( .A(n4299), .B(n4298), .Z(n4393) );
  XOR U5283 ( .A(n4299), .B(n4298), .Z(n4554) );
  NAND U5284 ( .A(a[16]), .B(b[44]), .Z(n4386) );
  NAND U5285 ( .A(a[13]), .B(b[44]), .Z(n4370) );
  XOR U5286 ( .A(n4301), .B(n4300), .Z(n4371) );
  OR U5287 ( .A(n4370), .B(n4371), .Z(n4373) );
  XNOR U5288 ( .A(n4303), .B(n4302), .Z(n4366) );
  XNOR U5289 ( .A(n4305), .B(n4304), .Z(n4362) );
  XOR U5290 ( .A(n4307), .B(n4306), .Z(n4358) );
  XNOR U5291 ( .A(n4309), .B(n4308), .Z(n4349) );
  XOR U5292 ( .A(n4311), .B(n4310), .Z(n4313) );
  AND U5293 ( .A(a[7]), .B(b[44]), .Z(n4312) );
  NANDN U5294 ( .A(n4313), .B(n4312), .Z(n4347) );
  XOR U5295 ( .A(n4313), .B(n4312), .Z(n4568) );
  XNOR U5296 ( .A(n4315), .B(n4314), .Z(n4337) );
  XNOR U5297 ( .A(n4317), .B(n4316), .Z(n4332) );
  XNOR U5298 ( .A(n4319), .B(n4318), .Z(n4328) );
  NAND U5299 ( .A(b[45]), .B(a[1]), .Z(n4321) );
  NAND U5300 ( .A(n4321), .B(n4320), .Z(n4324) );
  OR U5301 ( .A(n4321), .B(n5002), .Z(n4583) );
  NANDN U5302 ( .A(n4323), .B(n4583), .Z(n4322) );
  AND U5303 ( .A(n4324), .B(n4322), .Z(n4327) );
  XNOR U5304 ( .A(n4583), .B(n4323), .Z(n4325) );
  NAND U5305 ( .A(n4325), .B(n4324), .Z(n4579) );
  ANDN U5306 ( .B(b[44]), .A(n162), .Z(n4578) );
  OR U5307 ( .A(n4579), .B(n4578), .Z(n4326) );
  AND U5308 ( .A(n4327), .B(n4326), .Z(n4329) );
  OR U5309 ( .A(n4328), .B(n4329), .Z(n4331) );
  XNOR U5310 ( .A(n4329), .B(n4328), .Z(n4576) );
  ANDN U5311 ( .B(b[44]), .A(n21580), .Z(n4577) );
  OR U5312 ( .A(n4576), .B(n4577), .Z(n4330) );
  AND U5313 ( .A(n4331), .B(n4330), .Z(n4333) );
  OR U5314 ( .A(n4332), .B(n4333), .Z(n4335) );
  XNOR U5315 ( .A(n4333), .B(n4332), .Z(n4574) );
  ANDN U5316 ( .B(b[44]), .A(n163), .Z(n4575) );
  OR U5317 ( .A(n4574), .B(n4575), .Z(n4334) );
  AND U5318 ( .A(n4335), .B(n4334), .Z(n4336) );
  OR U5319 ( .A(n4337), .B(n4336), .Z(n4339) );
  XNOR U5320 ( .A(n4337), .B(n4336), .Z(n4602) );
  NAND U5321 ( .A(b[44]), .B(a[5]), .Z(n4603) );
  NANDN U5322 ( .A(n4602), .B(n4603), .Z(n4338) );
  NAND U5323 ( .A(n4339), .B(n4338), .Z(n4341) );
  AND U5324 ( .A(a[6]), .B(b[44]), .Z(n4340) );
  NANDN U5325 ( .A(n4341), .B(n4340), .Z(n4345) );
  XOR U5326 ( .A(n4341), .B(n4340), .Z(n4570) );
  XOR U5327 ( .A(n4343), .B(n4342), .Z(n4571) );
  NANDN U5328 ( .A(n4570), .B(n4571), .Z(n4344) );
  AND U5329 ( .A(n4345), .B(n4344), .Z(n4569) );
  OR U5330 ( .A(n4568), .B(n4569), .Z(n4346) );
  AND U5331 ( .A(n4347), .B(n4346), .Z(n4348) );
  OR U5332 ( .A(n4349), .B(n4348), .Z(n4351) );
  XNOR U5333 ( .A(n4349), .B(n4348), .Z(n4613) );
  NAND U5334 ( .A(a[8]), .B(b[44]), .Z(n4612) );
  OR U5335 ( .A(n4613), .B(n4612), .Z(n4350) );
  NAND U5336 ( .A(n4351), .B(n4350), .Z(n4354) );
  XOR U5337 ( .A(n4353), .B(n4352), .Z(n4355) );
  OR U5338 ( .A(n4354), .B(n4355), .Z(n4357) );
  ANDN U5339 ( .B(b[44]), .A(n21615), .Z(n4567) );
  XOR U5340 ( .A(n4355), .B(n4354), .Z(n4566) );
  NANDN U5341 ( .A(n4567), .B(n4566), .Z(n4356) );
  AND U5342 ( .A(n4357), .B(n4356), .Z(n4359) );
  OR U5343 ( .A(n4358), .B(n4359), .Z(n4361) );
  XNOR U5344 ( .A(n4359), .B(n4358), .Z(n4564) );
  ANDN U5345 ( .B(b[44]), .A(n168), .Z(n4565) );
  OR U5346 ( .A(n4564), .B(n4565), .Z(n4360) );
  AND U5347 ( .A(n4361), .B(n4360), .Z(n4363) );
  OR U5348 ( .A(n4362), .B(n4363), .Z(n4365) );
  XNOR U5349 ( .A(n4363), .B(n4362), .Z(n4562) );
  ANDN U5350 ( .B(b[44]), .A(n21164), .Z(n4563) );
  OR U5351 ( .A(n4562), .B(n4563), .Z(n4364) );
  AND U5352 ( .A(n4365), .B(n4364), .Z(n4367) );
  OR U5353 ( .A(n4366), .B(n4367), .Z(n4369) );
  XNOR U5354 ( .A(n4367), .B(n4366), .Z(n4561) );
  ANDN U5355 ( .B(b[44]), .A(n169), .Z(n4560) );
  OR U5356 ( .A(n4561), .B(n4560), .Z(n4368) );
  NAND U5357 ( .A(n4369), .B(n4368), .Z(n4635) );
  XOR U5358 ( .A(n4371), .B(n4370), .Z(n4634) );
  NANDN U5359 ( .A(n4635), .B(n4634), .Z(n4372) );
  AND U5360 ( .A(n4373), .B(n4372), .Z(n4376) );
  NANDN U5361 ( .A(n4376), .B(n4377), .Z(n4379) );
  XOR U5362 ( .A(n4377), .B(n4376), .Z(n4641) );
  AND U5363 ( .A(a[14]), .B(b[44]), .Z(n4640) );
  NANDN U5364 ( .A(n4641), .B(n4640), .Z(n4378) );
  AND U5365 ( .A(n4379), .B(n4378), .Z(n4383) );
  XNOR U5366 ( .A(n4381), .B(n4380), .Z(n4382) );
  NANDN U5367 ( .A(n4383), .B(n4382), .Z(n4385) );
  NAND U5368 ( .A(a[15]), .B(b[44]), .Z(n4649) );
  NANDN U5369 ( .A(n4649), .B(n4648), .Z(n4384) );
  AND U5370 ( .A(n4385), .B(n4384), .Z(n4387) );
  OR U5371 ( .A(n4386), .B(n4387), .Z(n4391) );
  XNOR U5372 ( .A(n4387), .B(n4386), .Z(n4557) );
  XNOR U5373 ( .A(n4389), .B(n4388), .Z(n4556) );
  NANDN U5374 ( .A(n4557), .B(n4556), .Z(n4390) );
  AND U5375 ( .A(n4391), .B(n4390), .Z(n4555) );
  OR U5376 ( .A(n4554), .B(n4555), .Z(n4392) );
  AND U5377 ( .A(n4393), .B(n4392), .Z(n4394) );
  OR U5378 ( .A(n4395), .B(n4394), .Z(n4397) );
  XNOR U5379 ( .A(n4395), .B(n4394), .Z(n4553) );
  AND U5380 ( .A(a[18]), .B(b[44]), .Z(n4552) );
  NANDN U5381 ( .A(n4553), .B(n4552), .Z(n4396) );
  AND U5382 ( .A(n4397), .B(n4396), .Z(n4401) );
  XNOR U5383 ( .A(n4399), .B(n4398), .Z(n4400) );
  NANDN U5384 ( .A(n4401), .B(n4400), .Z(n4403) );
  XOR U5385 ( .A(n4401), .B(n4400), .Z(n4663) );
  AND U5386 ( .A(a[19]), .B(b[44]), .Z(n4662) );
  NANDN U5387 ( .A(n4663), .B(n4662), .Z(n4402) );
  AND U5388 ( .A(n4403), .B(n4402), .Z(n4405) );
  OR U5389 ( .A(n4404), .B(n4405), .Z(n4409) );
  XNOR U5390 ( .A(n4405), .B(n4404), .Z(n4668) );
  NANDN U5391 ( .A(n4668), .B(n4669), .Z(n4408) );
  AND U5392 ( .A(n4409), .B(n4408), .Z(n4674) );
  OR U5393 ( .A(n4675), .B(n4674), .Z(n4410) );
  NAND U5394 ( .A(n4411), .B(n4410), .Z(n4415) );
  XNOR U5395 ( .A(n4413), .B(n4412), .Z(n4414) );
  NANDN U5396 ( .A(n4415), .B(n4414), .Z(n4417) );
  ANDN U5397 ( .B(b[44]), .A(n177), .Z(n4551) );
  XOR U5398 ( .A(n4415), .B(n4414), .Z(n4550) );
  OR U5399 ( .A(n4551), .B(n4550), .Z(n4416) );
  NAND U5400 ( .A(n4417), .B(n4416), .Z(n4684) );
  XOR U5401 ( .A(n4419), .B(n4418), .Z(n4685) );
  NANDN U5402 ( .A(n4684), .B(n4685), .Z(n4420) );
  AND U5403 ( .A(n4421), .B(n4420), .Z(n4424) );
  XNOR U5404 ( .A(n4423), .B(n4422), .Z(n4425) );
  NANDN U5405 ( .A(n4424), .B(n4425), .Z(n4427) );
  XOR U5406 ( .A(n4425), .B(n4424), .Z(n4548) );
  NAND U5407 ( .A(a[24]), .B(b[44]), .Z(n4549) );
  OR U5408 ( .A(n4548), .B(n4549), .Z(n4426) );
  AND U5409 ( .A(n4427), .B(n4426), .Z(n4546) );
  OR U5410 ( .A(n4547), .B(n4546), .Z(n4428) );
  NAND U5411 ( .A(n4429), .B(n4428), .Z(n4430) );
  NANDN U5412 ( .A(n4431), .B(n4430), .Z(n4433) );
  NAND U5413 ( .A(a[26]), .B(b[44]), .Z(n4699) );
  NANDN U5414 ( .A(n4699), .B(n4698), .Z(n4432) );
  NAND U5415 ( .A(n4433), .B(n4432), .Z(n4434) );
  NANDN U5416 ( .A(n4435), .B(n4434), .Z(n4437) );
  NAND U5417 ( .A(b[44]), .B(a[27]), .Z(n4544) );
  NANDN U5418 ( .A(n4544), .B(n4545), .Z(n4436) );
  NAND U5419 ( .A(n4437), .B(n4436), .Z(n4542) );
  NANDN U5420 ( .A(n4543), .B(n4542), .Z(n4438) );
  AND U5421 ( .A(n4439), .B(n4438), .Z(n4712) );
  XNOR U5422 ( .A(n4441), .B(n4440), .Z(n4713) );
  NANDN U5423 ( .A(n4712), .B(n4713), .Z(n4442) );
  NAND U5424 ( .A(n4443), .B(n4442), .Z(n4447) );
  XOR U5425 ( .A(n4445), .B(n4444), .Z(n4446) );
  NANDN U5426 ( .A(n4447), .B(n4446), .Z(n4449) );
  ANDN U5427 ( .B(b[44]), .A(n181), .Z(n4541) );
  XOR U5428 ( .A(n4447), .B(n4446), .Z(n4540) );
  OR U5429 ( .A(n4541), .B(n4540), .Z(n4448) );
  NAND U5430 ( .A(n4449), .B(n4448), .Z(n4450) );
  NANDN U5431 ( .A(n4451), .B(n4450), .Z(n4453) );
  ANDN U5432 ( .B(b[44]), .A(n21740), .Z(n4539) );
  NANDN U5433 ( .A(n4539), .B(n4538), .Z(n4452) );
  NAND U5434 ( .A(n4453), .B(n4452), .Z(n4728) );
  NANDN U5435 ( .A(n4729), .B(n4728), .Z(n4454) );
  NAND U5436 ( .A(n4455), .B(n4454), .Z(n4456) );
  NANDN U5437 ( .A(n4457), .B(n4456), .Z(n4459) );
  ANDN U5438 ( .B(b[44]), .A(n21751), .Z(n4733) );
  OR U5439 ( .A(n4733), .B(n4732), .Z(n4458) );
  NAND U5440 ( .A(n4459), .B(n4458), .Z(n4460) );
  NANDN U5441 ( .A(n4461), .B(n4460), .Z(n4463) );
  ANDN U5442 ( .B(b[44]), .A(n183), .Z(n4537) );
  NANDN U5443 ( .A(n4537), .B(n4536), .Z(n4462) );
  NAND U5444 ( .A(n4463), .B(n4462), .Z(n4535) );
  XOR U5445 ( .A(n4465), .B(n4464), .Z(n4534) );
  NAND U5446 ( .A(n4535), .B(n4534), .Z(n4466) );
  NAND U5447 ( .A(n4467), .B(n4466), .Z(n4746) );
  NANDN U5448 ( .A(n4747), .B(n4746), .Z(n4468) );
  NAND U5449 ( .A(n4469), .B(n4468), .Z(n4752) );
  OR U5450 ( .A(n4753), .B(n4752), .Z(n4470) );
  NAND U5451 ( .A(n4471), .B(n4470), .Z(n4533) );
  NANDN U5452 ( .A(n4532), .B(n4533), .Z(n4472) );
  NAND U5453 ( .A(n4473), .B(n4472), .Z(n4531) );
  XOR U5454 ( .A(n4475), .B(n4474), .Z(n4530) );
  NANDN U5455 ( .A(n4531), .B(n4530), .Z(n4476) );
  NAND U5456 ( .A(n4477), .B(n4476), .Z(n4478) );
  NANDN U5457 ( .A(n4479), .B(n4478), .Z(n4481) );
  ANDN U5458 ( .B(b[44]), .A(n188), .Z(n4767) );
  OR U5459 ( .A(n4767), .B(n4766), .Z(n4480) );
  AND U5460 ( .A(n4481), .B(n4480), .Z(n4483) );
  OR U5461 ( .A(n4482), .B(n4483), .Z(n4485) );
  XNOR U5462 ( .A(n4483), .B(n4482), .Z(n4528) );
  NAND U5463 ( .A(b[44]), .B(a[41]), .Z(n4529) );
  NANDN U5464 ( .A(n4528), .B(n4529), .Z(n4484) );
  AND U5465 ( .A(n4485), .B(n4484), .Z(n4487) );
  OR U5466 ( .A(n4486), .B(n4487), .Z(n4489) );
  XNOR U5467 ( .A(n4487), .B(n4486), .Z(n4776) );
  ANDN U5468 ( .B(b[44]), .A(n190), .Z(n4777) );
  OR U5469 ( .A(n4776), .B(n4777), .Z(n4488) );
  NAND U5470 ( .A(n4489), .B(n4488), .Z(n4527) );
  XOR U5471 ( .A(n4491), .B(n4490), .Z(n4526) );
  OR U5472 ( .A(n4527), .B(n4526), .Z(n4492) );
  NAND U5473 ( .A(n4493), .B(n4492), .Z(n4497) );
  OR U5474 ( .A(n4497), .B(n4496), .Z(n4499) );
  ANDN U5475 ( .B(b[44]), .A(n192), .Z(n4525) );
  XOR U5476 ( .A(n4497), .B(n4496), .Z(n4524) );
  NANDN U5477 ( .A(n4525), .B(n4524), .Z(n4498) );
  AND U5478 ( .A(n4499), .B(n4498), .Z(n4501) );
  OR U5479 ( .A(n4500), .B(n4501), .Z(n4503) );
  XNOR U5480 ( .A(n4501), .B(n4500), .Z(n4790) );
  NAND U5481 ( .A(b[44]), .B(a[45]), .Z(n4791) );
  NANDN U5482 ( .A(n4790), .B(n4791), .Z(n4502) );
  AND U5483 ( .A(n4503), .B(n4502), .Z(n4505) );
  OR U5484 ( .A(n4504), .B(n4505), .Z(n4507) );
  XNOR U5485 ( .A(n4505), .B(n4504), .Z(n4520) );
  ANDN U5486 ( .B(b[44]), .A(n194), .Z(n4521) );
  OR U5487 ( .A(n4520), .B(n4521), .Z(n4506) );
  AND U5488 ( .A(n4507), .B(n4506), .Z(n4509) );
  OR U5489 ( .A(n4508), .B(n4509), .Z(n4511) );
  XNOR U5490 ( .A(n4509), .B(n4508), .Z(n4518) );
  ANDN U5491 ( .B(b[44]), .A(n195), .Z(n4519) );
  OR U5492 ( .A(n4518), .B(n4519), .Z(n4510) );
  AND U5493 ( .A(n4511), .B(n4510), .Z(n4514) );
  OR U5494 ( .A(n4514), .B(n4515), .Z(n4517) );
  XOR U5495 ( .A(n4515), .B(n4514), .Z(n4802) );
  NAND U5496 ( .A(b[44]), .B(a[48]), .Z(n4803) );
  NAND U5497 ( .A(n4802), .B(n4803), .Z(n4516) );
  NAND U5498 ( .A(n4517), .B(n4516), .Z(n4813) );
  NAND U5499 ( .A(a[49]), .B(b[44]), .Z(n4815) );
  XNOR U5500 ( .A(n4814), .B(n4815), .Z(n4808) );
  ANDN U5501 ( .B(b[43]), .A(n198), .Z(n4809) );
  OR U5502 ( .A(n4808), .B(n4809), .Z(n4811) );
  XNOR U5503 ( .A(n4519), .B(n4518), .Z(n4798) );
  XNOR U5504 ( .A(n4521), .B(n4520), .Z(n4522) );
  ANDN U5505 ( .B(b[43]), .A(n195), .Z(n4523) );
  OR U5506 ( .A(n4522), .B(n4523), .Z(n4797) );
  XNOR U5507 ( .A(n4523), .B(n4522), .Z(n4931) );
  XOR U5508 ( .A(n4525), .B(n4524), .Z(n4786) );
  XOR U5509 ( .A(n4527), .B(n4526), .Z(n4783) );
  NAND U5510 ( .A(a[42]), .B(b[43]), .Z(n4773) );
  XOR U5511 ( .A(n4529), .B(n4528), .Z(n4772) );
  NANDN U5512 ( .A(n4773), .B(n4772), .Z(n4775) );
  NAND U5513 ( .A(a[40]), .B(b[43]), .Z(n4763) );
  XOR U5514 ( .A(n4531), .B(n4530), .Z(n4762) );
  NANDN U5515 ( .A(n4763), .B(n4762), .Z(n4765) );
  ANDN U5516 ( .B(b[43]), .A(n187), .Z(n4759) );
  XNOR U5517 ( .A(n4533), .B(n4532), .Z(n4758) );
  OR U5518 ( .A(n4759), .B(n4758), .Z(n4761) );
  XNOR U5519 ( .A(n4535), .B(n4534), .Z(n4743) );
  XOR U5520 ( .A(n4537), .B(n4536), .Z(n4739) );
  ANDN U5521 ( .B(b[43]), .A(n182), .Z(n4723) );
  XOR U5522 ( .A(n4539), .B(n4538), .Z(n4722) );
  OR U5523 ( .A(n4723), .B(n4722), .Z(n4725) );
  XNOR U5524 ( .A(n4541), .B(n4540), .Z(n4719) );
  XOR U5525 ( .A(n4543), .B(n4542), .Z(n4709) );
  NAND U5526 ( .A(b[43]), .B(a[29]), .Z(n4708) );
  OR U5527 ( .A(n4709), .B(n4708), .Z(n4711) );
  XOR U5528 ( .A(n4545), .B(n4544), .Z(n4705) );
  XOR U5529 ( .A(n4547), .B(n4546), .Z(n4695) );
  XOR U5530 ( .A(n4549), .B(n4548), .Z(n4691) );
  XOR U5531 ( .A(n4551), .B(n4550), .Z(n4681) );
  NAND U5532 ( .A(a[19]), .B(b[43]), .Z(n4659) );
  XNOR U5533 ( .A(n4553), .B(n4552), .Z(n4658) );
  NANDN U5534 ( .A(n4659), .B(n4658), .Z(n4661) );
  XNOR U5535 ( .A(n4555), .B(n4554), .Z(n4655) );
  AND U5536 ( .A(a[17]), .B(b[43]), .Z(n4558) );
  NANDN U5537 ( .A(n4559), .B(n4558), .Z(n4653) );
  XOR U5538 ( .A(n4559), .B(n4558), .Z(n4974) );
  NAND U5539 ( .A(a[16]), .B(b[43]), .Z(n4646) );
  NAND U5540 ( .A(a[13]), .B(b[43]), .Z(n4630) );
  XOR U5541 ( .A(n4561), .B(n4560), .Z(n4631) );
  OR U5542 ( .A(n4630), .B(n4631), .Z(n4633) );
  XNOR U5543 ( .A(n4563), .B(n4562), .Z(n4626) );
  XNOR U5544 ( .A(n4565), .B(n4564), .Z(n4622) );
  XOR U5545 ( .A(n4567), .B(n4566), .Z(n4618) );
  XNOR U5546 ( .A(n4569), .B(n4568), .Z(n4609) );
  XOR U5547 ( .A(n4571), .B(n4570), .Z(n4573) );
  AND U5548 ( .A(a[7]), .B(b[43]), .Z(n4572) );
  NANDN U5549 ( .A(n4573), .B(n4572), .Z(n4607) );
  XOR U5550 ( .A(n4573), .B(n4572), .Z(n4990) );
  XNOR U5551 ( .A(n4575), .B(n4574), .Z(n4597) );
  XNOR U5552 ( .A(n4577), .B(n4576), .Z(n4592) );
  XNOR U5553 ( .A(n4579), .B(n4578), .Z(n4588) );
  NAND U5554 ( .A(b[44]), .B(a[1]), .Z(n4581) );
  NAND U5555 ( .A(n4581), .B(n4580), .Z(n4584) );
  NANDN U5556 ( .A(n156), .B(a[0]), .Z(n5312) );
  OR U5557 ( .A(n4581), .B(n5312), .Z(n5005) );
  NANDN U5558 ( .A(n4583), .B(n5005), .Z(n4582) );
  AND U5559 ( .A(n4584), .B(n4582), .Z(n4587) );
  XNOR U5560 ( .A(n5005), .B(n4583), .Z(n4585) );
  NAND U5561 ( .A(n4585), .B(n4584), .Z(n5001) );
  ANDN U5562 ( .B(b[43]), .A(n162), .Z(n5000) );
  OR U5563 ( .A(n5001), .B(n5000), .Z(n4586) );
  AND U5564 ( .A(n4587), .B(n4586), .Z(n4589) );
  OR U5565 ( .A(n4588), .B(n4589), .Z(n4591) );
  XNOR U5566 ( .A(n4589), .B(n4588), .Z(n4998) );
  ANDN U5567 ( .B(b[43]), .A(n21580), .Z(n4999) );
  OR U5568 ( .A(n4998), .B(n4999), .Z(n4590) );
  AND U5569 ( .A(n4591), .B(n4590), .Z(n4593) );
  OR U5570 ( .A(n4592), .B(n4593), .Z(n4595) );
  XNOR U5571 ( .A(n4593), .B(n4592), .Z(n4996) );
  ANDN U5572 ( .B(b[43]), .A(n163), .Z(n4997) );
  OR U5573 ( .A(n4996), .B(n4997), .Z(n4594) );
  AND U5574 ( .A(n4595), .B(n4594), .Z(n4596) );
  OR U5575 ( .A(n4597), .B(n4596), .Z(n4599) );
  XNOR U5576 ( .A(n4597), .B(n4596), .Z(n5024) );
  NAND U5577 ( .A(b[43]), .B(a[5]), .Z(n5025) );
  NANDN U5578 ( .A(n5024), .B(n5025), .Z(n4598) );
  NAND U5579 ( .A(n4599), .B(n4598), .Z(n4601) );
  AND U5580 ( .A(a[6]), .B(b[43]), .Z(n4600) );
  NANDN U5581 ( .A(n4601), .B(n4600), .Z(n4605) );
  XOR U5582 ( .A(n4601), .B(n4600), .Z(n4992) );
  XOR U5583 ( .A(n4603), .B(n4602), .Z(n4993) );
  NANDN U5584 ( .A(n4992), .B(n4993), .Z(n4604) );
  AND U5585 ( .A(n4605), .B(n4604), .Z(n4991) );
  OR U5586 ( .A(n4990), .B(n4991), .Z(n4606) );
  AND U5587 ( .A(n4607), .B(n4606), .Z(n4608) );
  OR U5588 ( .A(n4609), .B(n4608), .Z(n4611) );
  XNOR U5589 ( .A(n4609), .B(n4608), .Z(n5035) );
  NAND U5590 ( .A(a[8]), .B(b[43]), .Z(n5034) );
  OR U5591 ( .A(n5035), .B(n5034), .Z(n4610) );
  NAND U5592 ( .A(n4611), .B(n4610), .Z(n4614) );
  XOR U5593 ( .A(n4613), .B(n4612), .Z(n4615) );
  OR U5594 ( .A(n4614), .B(n4615), .Z(n4617) );
  ANDN U5595 ( .B(b[43]), .A(n21615), .Z(n4989) );
  XOR U5596 ( .A(n4615), .B(n4614), .Z(n4988) );
  NANDN U5597 ( .A(n4989), .B(n4988), .Z(n4616) );
  AND U5598 ( .A(n4617), .B(n4616), .Z(n4619) );
  OR U5599 ( .A(n4618), .B(n4619), .Z(n4621) );
  XNOR U5600 ( .A(n4619), .B(n4618), .Z(n4986) );
  ANDN U5601 ( .B(b[43]), .A(n168), .Z(n4987) );
  OR U5602 ( .A(n4986), .B(n4987), .Z(n4620) );
  AND U5603 ( .A(n4621), .B(n4620), .Z(n4623) );
  OR U5604 ( .A(n4622), .B(n4623), .Z(n4625) );
  XNOR U5605 ( .A(n4623), .B(n4622), .Z(n4984) );
  ANDN U5606 ( .B(b[43]), .A(n21164), .Z(n4985) );
  OR U5607 ( .A(n4984), .B(n4985), .Z(n4624) );
  AND U5608 ( .A(n4625), .B(n4624), .Z(n4627) );
  OR U5609 ( .A(n4626), .B(n4627), .Z(n4629) );
  XNOR U5610 ( .A(n4627), .B(n4626), .Z(n4982) );
  NAND U5611 ( .A(b[43]), .B(a[12]), .Z(n4983) );
  NANDN U5612 ( .A(n4982), .B(n4983), .Z(n4628) );
  NAND U5613 ( .A(n4629), .B(n4628), .Z(n5057) );
  XOR U5614 ( .A(n4631), .B(n4630), .Z(n5056) );
  NANDN U5615 ( .A(n5057), .B(n5056), .Z(n4632) );
  AND U5616 ( .A(n4633), .B(n4632), .Z(n4636) );
  NANDN U5617 ( .A(n4636), .B(n4637), .Z(n4639) );
  XOR U5618 ( .A(n4637), .B(n4636), .Z(n4981) );
  AND U5619 ( .A(a[14]), .B(b[43]), .Z(n4980) );
  NANDN U5620 ( .A(n4981), .B(n4980), .Z(n4638) );
  AND U5621 ( .A(n4639), .B(n4638), .Z(n4642) );
  XNOR U5622 ( .A(n4641), .B(n4640), .Z(n4643) );
  NANDN U5623 ( .A(n4642), .B(n4643), .Z(n4645) );
  XOR U5624 ( .A(n4643), .B(n4642), .Z(n5069) );
  AND U5625 ( .A(a[15]), .B(b[43]), .Z(n5068) );
  NANDN U5626 ( .A(n5069), .B(n5068), .Z(n4644) );
  AND U5627 ( .A(n4645), .B(n4644), .Z(n4647) );
  OR U5628 ( .A(n4646), .B(n4647), .Z(n4651) );
  XNOR U5629 ( .A(n4647), .B(n4646), .Z(n4977) );
  NANDN U5630 ( .A(n4977), .B(n4976), .Z(n4650) );
  AND U5631 ( .A(n4651), .B(n4650), .Z(n4975) );
  OR U5632 ( .A(n4974), .B(n4975), .Z(n4652) );
  AND U5633 ( .A(n4653), .B(n4652), .Z(n4654) );
  OR U5634 ( .A(n4655), .B(n4654), .Z(n4657) );
  XNOR U5635 ( .A(n4655), .B(n4654), .Z(n4973) );
  AND U5636 ( .A(a[18]), .B(b[43]), .Z(n4972) );
  NANDN U5637 ( .A(n4973), .B(n4972), .Z(n4656) );
  AND U5638 ( .A(n4657), .B(n4656), .Z(n4970) );
  NANDN U5639 ( .A(n4970), .B(n4971), .Z(n4660) );
  AND U5640 ( .A(n4661), .B(n4660), .Z(n4665) );
  XNOR U5641 ( .A(n4663), .B(n4662), .Z(n4664) );
  NANDN U5642 ( .A(n4665), .B(n4664), .Z(n4667) );
  NAND U5643 ( .A(a[20]), .B(b[43]), .Z(n4969) );
  NANDN U5644 ( .A(n4969), .B(n4968), .Z(n4666) );
  NAND U5645 ( .A(n4667), .B(n4666), .Z(n4670) );
  XNOR U5646 ( .A(n4669), .B(n4668), .Z(n4671) );
  OR U5647 ( .A(n4670), .B(n4671), .Z(n4673) );
  XNOR U5648 ( .A(n4671), .B(n4670), .Z(n5090) );
  NAND U5649 ( .A(b[43]), .B(a[21]), .Z(n5091) );
  NANDN U5650 ( .A(n5090), .B(n5091), .Z(n4672) );
  NAND U5651 ( .A(n4673), .B(n4672), .Z(n4677) );
  XOR U5652 ( .A(n4675), .B(n4674), .Z(n4676) );
  NANDN U5653 ( .A(n4677), .B(n4676), .Z(n4679) );
  NAND U5654 ( .A(a[22]), .B(b[43]), .Z(n4967) );
  XNOR U5655 ( .A(n4677), .B(n4676), .Z(n4966) );
  NANDN U5656 ( .A(n4967), .B(n4966), .Z(n4678) );
  NAND U5657 ( .A(n4679), .B(n4678), .Z(n4680) );
  NANDN U5658 ( .A(n4681), .B(n4680), .Z(n4683) );
  NAND U5659 ( .A(b[43]), .B(a[23]), .Z(n5102) );
  NANDN U5660 ( .A(n5102), .B(n5103), .Z(n4682) );
  NAND U5661 ( .A(n4683), .B(n4682), .Z(n4687) );
  XOR U5662 ( .A(n4685), .B(n4684), .Z(n4686) );
  NANDN U5663 ( .A(n4687), .B(n4686), .Z(n4689) );
  ANDN U5664 ( .B(b[43]), .A(n178), .Z(n5107) );
  OR U5665 ( .A(n5107), .B(n5106), .Z(n4688) );
  NAND U5666 ( .A(n4689), .B(n4688), .Z(n4690) );
  NANDN U5667 ( .A(n4691), .B(n4690), .Z(n4693) );
  ANDN U5668 ( .B(b[43]), .A(n21703), .Z(n5113) );
  NANDN U5669 ( .A(n5113), .B(n5112), .Z(n4692) );
  NAND U5670 ( .A(n4693), .B(n4692), .Z(n4694) );
  NANDN U5671 ( .A(n4695), .B(n4694), .Z(n4697) );
  ANDN U5672 ( .B(b[43]), .A(n179), .Z(n4963) );
  NANDN U5673 ( .A(n4963), .B(n4962), .Z(n4696) );
  NAND U5674 ( .A(n4697), .B(n4696), .Z(n4701) );
  XNOR U5675 ( .A(n4699), .B(n4698), .Z(n4700) );
  NANDN U5676 ( .A(n4701), .B(n4700), .Z(n4703) );
  NAND U5677 ( .A(b[43]), .B(a[27]), .Z(n5120) );
  XNOR U5678 ( .A(n4701), .B(n4700), .Z(n5121) );
  NANDN U5679 ( .A(n5120), .B(n5121), .Z(n4702) );
  NAND U5680 ( .A(n4703), .B(n4702), .Z(n4704) );
  NANDN U5681 ( .A(n4705), .B(n4704), .Z(n4707) );
  XOR U5682 ( .A(n4705), .B(n4704), .Z(n5127) );
  NAND U5683 ( .A(b[43]), .B(a[28]), .Z(n5126) );
  OR U5684 ( .A(n5127), .B(n5126), .Z(n4706) );
  AND U5685 ( .A(n4707), .B(n4706), .Z(n5132) );
  XOR U5686 ( .A(n4709), .B(n4708), .Z(n5133) );
  NANDN U5687 ( .A(n5132), .B(n5133), .Z(n4710) );
  NAND U5688 ( .A(n4711), .B(n4710), .Z(n4715) );
  XOR U5689 ( .A(n4713), .B(n4712), .Z(n4714) );
  NANDN U5690 ( .A(n4715), .B(n4714), .Z(n4717) );
  ANDN U5691 ( .B(b[43]), .A(n181), .Z(n4961) );
  NANDN U5692 ( .A(n4961), .B(n4960), .Z(n4716) );
  NAND U5693 ( .A(n4717), .B(n4716), .Z(n4718) );
  NANDN U5694 ( .A(n4719), .B(n4718), .Z(n4721) );
  ANDN U5695 ( .B(b[43]), .A(n21740), .Z(n4958) );
  NANDN U5696 ( .A(n4958), .B(n4959), .Z(n4720) );
  NAND U5697 ( .A(n4721), .B(n4720), .Z(n4956) );
  XOR U5698 ( .A(n4723), .B(n4722), .Z(n4957) );
  NAND U5699 ( .A(n4956), .B(n4957), .Z(n4724) );
  NAND U5700 ( .A(n4725), .B(n4724), .Z(n4727) );
  NAND U5701 ( .A(b[43]), .B(a[33]), .Z(n4726) );
  OR U5702 ( .A(n4727), .B(n4726), .Z(n4731) );
  XOR U5703 ( .A(n4727), .B(n4726), .Z(n4954) );
  NAND U5704 ( .A(n4954), .B(n4955), .Z(n4730) );
  NAND U5705 ( .A(n4731), .B(n4730), .Z(n4735) );
  XOR U5706 ( .A(n4733), .B(n4732), .Z(n4734) );
  NANDN U5707 ( .A(n4735), .B(n4734), .Z(n4737) );
  ANDN U5708 ( .B(b[43]), .A(n183), .Z(n5155) );
  XOR U5709 ( .A(n4735), .B(n4734), .Z(n5154) );
  OR U5710 ( .A(n5155), .B(n5154), .Z(n4736) );
  NAND U5711 ( .A(n4737), .B(n4736), .Z(n4738) );
  NANDN U5712 ( .A(n4739), .B(n4738), .Z(n4741) );
  ANDN U5713 ( .B(b[43]), .A(n184), .Z(n4953) );
  NANDN U5714 ( .A(n4953), .B(n4952), .Z(n4740) );
  NAND U5715 ( .A(n4741), .B(n4740), .Z(n4742) );
  NANDN U5716 ( .A(n4743), .B(n4742), .Z(n4745) );
  ANDN U5717 ( .B(b[43]), .A(n185), .Z(n4951) );
  NANDN U5718 ( .A(n4951), .B(n4950), .Z(n4744) );
  NAND U5719 ( .A(n4745), .B(n4744), .Z(n4749) );
  NAND U5720 ( .A(n4749), .B(n4748), .Z(n4751) );
  ANDN U5721 ( .B(b[43]), .A(n21772), .Z(n4949) );
  XNOR U5722 ( .A(n4749), .B(n4748), .Z(n4948) );
  OR U5723 ( .A(n4949), .B(n4948), .Z(n4750) );
  NAND U5724 ( .A(n4751), .B(n4750), .Z(n4755) );
  XOR U5725 ( .A(n4753), .B(n4752), .Z(n4754) );
  NANDN U5726 ( .A(n4755), .B(n4754), .Z(n4757) );
  XOR U5727 ( .A(n4755), .B(n4754), .Z(n4946) );
  NAND U5728 ( .A(a[38]), .B(b[43]), .Z(n4947) );
  OR U5729 ( .A(n4946), .B(n4947), .Z(n4756) );
  AND U5730 ( .A(n4757), .B(n4756), .Z(n4944) );
  XOR U5731 ( .A(n4759), .B(n4758), .Z(n4945) );
  NAND U5732 ( .A(n4944), .B(n4945), .Z(n4760) );
  NAND U5733 ( .A(n4761), .B(n4760), .Z(n4942) );
  NANDN U5734 ( .A(n4942), .B(n4943), .Z(n4764) );
  NAND U5735 ( .A(n4765), .B(n4764), .Z(n4769) );
  XOR U5736 ( .A(n4767), .B(n4766), .Z(n4768) );
  NANDN U5737 ( .A(n4769), .B(n4768), .Z(n4771) );
  ANDN U5738 ( .B(b[43]), .A(n189), .Z(n4941) );
  XOR U5739 ( .A(n4769), .B(n4768), .Z(n4940) );
  OR U5740 ( .A(n4941), .B(n4940), .Z(n4770) );
  NAND U5741 ( .A(n4771), .B(n4770), .Z(n5189) );
  XNOR U5742 ( .A(n4773), .B(n4772), .Z(n5188) );
  NANDN U5743 ( .A(n5189), .B(n5188), .Z(n4774) );
  NAND U5744 ( .A(n4775), .B(n4774), .Z(n4779) );
  XOR U5745 ( .A(n4777), .B(n4776), .Z(n4778) );
  NANDN U5746 ( .A(n4779), .B(n4778), .Z(n4781) );
  ANDN U5747 ( .B(b[43]), .A(n191), .Z(n4939) );
  XOR U5748 ( .A(n4779), .B(n4778), .Z(n4938) );
  OR U5749 ( .A(n4939), .B(n4938), .Z(n4780) );
  NAND U5750 ( .A(n4781), .B(n4780), .Z(n4782) );
  NANDN U5751 ( .A(n4783), .B(n4782), .Z(n4785) );
  ANDN U5752 ( .B(b[43]), .A(n192), .Z(n4937) );
  NANDN U5753 ( .A(n4937), .B(n4936), .Z(n4784) );
  AND U5754 ( .A(n4785), .B(n4784), .Z(n4787) );
  OR U5755 ( .A(n4786), .B(n4787), .Z(n4789) );
  XNOR U5756 ( .A(n4787), .B(n4786), .Z(n4934) );
  ANDN U5757 ( .B(b[43]), .A(n193), .Z(n4935) );
  OR U5758 ( .A(n4934), .B(n4935), .Z(n4788) );
  NAND U5759 ( .A(n4789), .B(n4788), .Z(n4793) );
  XOR U5760 ( .A(n4791), .B(n4790), .Z(n4792) );
  NANDN U5761 ( .A(n4793), .B(n4792), .Z(n4795) );
  NAND U5762 ( .A(a[46]), .B(b[43]), .Z(n4933) );
  NANDN U5763 ( .A(n4933), .B(n4932), .Z(n4794) );
  NAND U5764 ( .A(n4795), .B(n4794), .Z(n4930) );
  OR U5765 ( .A(n4931), .B(n4930), .Z(n4796) );
  AND U5766 ( .A(n4797), .B(n4796), .Z(n4799) );
  OR U5767 ( .A(n4798), .B(n4799), .Z(n4801) );
  XNOR U5768 ( .A(n4799), .B(n4798), .Z(n4928) );
  ANDN U5769 ( .B(b[43]), .A(n196), .Z(n4929) );
  OR U5770 ( .A(n4928), .B(n4929), .Z(n4800) );
  NAND U5771 ( .A(n4801), .B(n4800), .Z(n4805) );
  NANDN U5772 ( .A(n4805), .B(n4804), .Z(n4807) );
  NAND U5773 ( .A(a[49]), .B(b[43]), .Z(n4926) );
  NANDN U5774 ( .A(n4926), .B(n4927), .Z(n4806) );
  NAND U5775 ( .A(n4807), .B(n4806), .Z(n5223) );
  XOR U5776 ( .A(n4809), .B(n4808), .Z(n5222) );
  NANDN U5777 ( .A(n5223), .B(n5222), .Z(n4810) );
  NAND U5778 ( .A(n4811), .B(n4810), .Z(n5663) );
  NANDN U5779 ( .A(n4813), .B(n4812), .Z(n4817) );
  NANDN U5780 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U5781 ( .A(n4817), .B(n4816), .Z(n5549) );
  NAND U5782 ( .A(b[47]), .B(a[47]), .Z(n5562) );
  NANDN U5783 ( .A(n4819), .B(n4818), .Z(n4823) );
  OR U5784 ( .A(n4821), .B(n4820), .Z(n4822) );
  AND U5785 ( .A(n4823), .B(n4822), .Z(n5561) );
  NANDN U5786 ( .A(n4825), .B(n4824), .Z(n4829) );
  OR U5787 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5788 ( .A(n4829), .B(n4828), .Z(n5567) );
  ANDN U5789 ( .B(b[50]), .A(n192), .Z(n5644) );
  OR U5790 ( .A(n4831), .B(n4830), .Z(n4835) );
  OR U5791 ( .A(n4833), .B(n4832), .Z(n4834) );
  AND U5792 ( .A(n4835), .B(n4834), .Z(n5645) );
  XNOR U5793 ( .A(n5644), .B(n5645), .Z(n5647) );
  NAND U5794 ( .A(a[42]), .B(b[52]), .Z(n5639) );
  OR U5795 ( .A(n4837), .B(n4836), .Z(n4841) );
  OR U5796 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5797 ( .A(n4841), .B(n4840), .Z(n5638) );
  XNOR U5798 ( .A(n5639), .B(n5638), .Z(n5641) );
  NAND U5799 ( .A(a[41]), .B(b[53]), .Z(n5581) );
  NANDN U5800 ( .A(n4843), .B(n4842), .Z(n4847) );
  OR U5801 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5802 ( .A(n4847), .B(n4846), .Z(n5579) );
  NAND U5803 ( .A(a[39]), .B(b[55]), .Z(n5587) );
  OR U5804 ( .A(n4849), .B(n4848), .Z(n4853) );
  OR U5805 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U5806 ( .A(n4853), .B(n4852), .Z(n5584) );
  ANDN U5807 ( .B(b[56]), .A(n186), .Z(n5626) );
  OR U5808 ( .A(n4855), .B(n4854), .Z(n4859) );
  NANDN U5809 ( .A(n4857), .B(n4856), .Z(n4858) );
  AND U5810 ( .A(n4859), .B(n4858), .Z(n5627) );
  XNOR U5811 ( .A(n5626), .B(n5627), .Z(n5629) );
  NAND U5812 ( .A(b[59]), .B(a[35]), .Z(n5598) );
  OR U5813 ( .A(n4861), .B(n4860), .Z(n4865) );
  NANDN U5814 ( .A(n4863), .B(n4862), .Z(n4864) );
  NAND U5815 ( .A(n4865), .B(n4864), .Z(n5597) );
  ANDN U5816 ( .B(b[61]), .A(n21751), .Z(n5604) );
  OR U5817 ( .A(n4867), .B(n4866), .Z(n4871) );
  OR U5818 ( .A(n4869), .B(n4868), .Z(n4870) );
  AND U5819 ( .A(n4871), .B(n4870), .Z(n5602) );
  ANDN U5820 ( .B(b[63]), .A(n21740), .Z(n5610) );
  ANDN U5821 ( .B(a[32]), .A(n159), .Z(n5608) );
  OR U5822 ( .A(n4873), .B(n4872), .Z(n4877) );
  OR U5823 ( .A(n4875), .B(n4874), .Z(n4876) );
  AND U5824 ( .A(n4877), .B(n4876), .Z(n5609) );
  XNOR U5825 ( .A(n5608), .B(n5609), .Z(n5611) );
  XNOR U5826 ( .A(n5610), .B(n5611), .Z(n5603) );
  XNOR U5827 ( .A(n5602), .B(n5603), .Z(n5605) );
  XNOR U5828 ( .A(n5604), .B(n5605), .Z(n5617) );
  ANDN U5829 ( .B(b[60]), .A(n183), .Z(n5614) );
  OR U5830 ( .A(n4879), .B(n4878), .Z(n4883) );
  OR U5831 ( .A(n4881), .B(n4880), .Z(n4882) );
  AND U5832 ( .A(n4883), .B(n4882), .Z(n5615) );
  XOR U5833 ( .A(n5614), .B(n5615), .Z(n5616) );
  NAND U5834 ( .A(a[36]), .B(b[58]), .Z(n5621) );
  OR U5835 ( .A(n4885), .B(n4884), .Z(n4889) );
  NANDN U5836 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5837 ( .A(n4889), .B(n4888), .Z(n5620) );
  XNOR U5838 ( .A(n5621), .B(n5620), .Z(n5623) );
  XNOR U5839 ( .A(n5622), .B(n5623), .Z(n5590) );
  OR U5840 ( .A(n4891), .B(n4890), .Z(n4895) );
  OR U5841 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U5842 ( .A(n4895), .B(n4894), .Z(n5591) );
  XNOR U5843 ( .A(n5590), .B(n5591), .Z(n5593) );
  ANDN U5844 ( .B(b[57]), .A(n21772), .Z(n5592) );
  XNOR U5845 ( .A(n5593), .B(n5592), .Z(n5628) );
  XOR U5846 ( .A(n5629), .B(n5628), .Z(n5585) );
  XNOR U5847 ( .A(n5584), .B(n5585), .Z(n5586) );
  XOR U5848 ( .A(n5587), .B(n5586), .Z(n5635) );
  ANDN U5849 ( .B(b[54]), .A(n188), .Z(n5632) );
  OR U5850 ( .A(n4897), .B(n4896), .Z(n4901) );
  OR U5851 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U5852 ( .A(n4901), .B(n4900), .Z(n5633) );
  XOR U5853 ( .A(n5632), .B(n5633), .Z(n5634) );
  XNOR U5854 ( .A(n5635), .B(n5634), .Z(n5578) );
  XNOR U5855 ( .A(n5579), .B(n5578), .Z(n5580) );
  XOR U5856 ( .A(n5581), .B(n5580), .Z(n5640) );
  OR U5857 ( .A(n4903), .B(n4902), .Z(n4907) );
  NANDN U5858 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U5859 ( .A(n4907), .B(n4906), .Z(n5573) );
  XOR U5860 ( .A(n5572), .B(n5573), .Z(n5574) );
  ANDN U5861 ( .B(b[51]), .A(n191), .Z(n5575) );
  XOR U5862 ( .A(n5574), .B(n5575), .Z(n5646) );
  XOR U5863 ( .A(n5647), .B(n5646), .Z(n5566) );
  XOR U5864 ( .A(n5567), .B(n5566), .Z(n5568) );
  NAND U5865 ( .A(a[45]), .B(b[49]), .Z(n5569) );
  ANDN U5866 ( .B(b[48]), .A(n194), .Z(n5650) );
  OR U5867 ( .A(n4909), .B(n4908), .Z(n4913) );
  NANDN U5868 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U5869 ( .A(n4913), .B(n4912), .Z(n5651) );
  XNOR U5870 ( .A(n5650), .B(n5651), .Z(n5653) );
  XOR U5871 ( .A(n5652), .B(n5653), .Z(n5560) );
  NAND U5872 ( .A(a[48]), .B(b[46]), .Z(n5657) );
  OR U5873 ( .A(n4915), .B(n4914), .Z(n4919) );
  NANDN U5874 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U5875 ( .A(n4919), .B(n4918), .Z(n5656) );
  XNOR U5876 ( .A(n5657), .B(n5656), .Z(n5659) );
  XNOR U5877 ( .A(n5658), .B(n5659), .Z(n5554) );
  NANDN U5878 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U5879 ( .A(n4923), .B(n4922), .Z(n4924) );
  AND U5880 ( .A(n4925), .B(n4924), .Z(n5555) );
  XNOR U5881 ( .A(n5554), .B(n5555), .Z(n5557) );
  ANDN U5882 ( .B(b[45]), .A(n197), .Z(n5556) );
  XOR U5883 ( .A(n5557), .B(n5556), .Z(n5548) );
  ANDN U5884 ( .B(b[44]), .A(n198), .Z(n5551) );
  XNOR U5885 ( .A(n5663), .B(n5662), .Z(n5664) );
  XNOR U5886 ( .A(n4927), .B(n4926), .Z(n5218) );
  XNOR U5887 ( .A(n4929), .B(n4928), .Z(n5214) );
  XNOR U5888 ( .A(n4931), .B(n4930), .Z(n5210) );
  XNOR U5889 ( .A(n4933), .B(n4932), .Z(n5207) );
  XNOR U5890 ( .A(n4935), .B(n4934), .Z(n5203) );
  XOR U5891 ( .A(n4937), .B(n4936), .Z(n5199) );
  XNOR U5892 ( .A(n4939), .B(n4938), .Z(n5195) );
  NAND U5893 ( .A(a[42]), .B(b[42]), .Z(n5184) );
  XNOR U5894 ( .A(n4941), .B(n4940), .Z(n5185) );
  NANDN U5895 ( .A(n5184), .B(n5185), .Z(n5187) );
  XNOR U5896 ( .A(n4943), .B(n4942), .Z(n5181) );
  XNOR U5897 ( .A(n4945), .B(n4944), .Z(n5177) );
  XOR U5898 ( .A(n4947), .B(n4946), .Z(n5173) );
  XNOR U5899 ( .A(n4949), .B(n4948), .Z(n5168) );
  ANDN U5900 ( .B(b[42]), .A(n21772), .Z(n5165) );
  XOR U5901 ( .A(n4951), .B(n4950), .Z(n5164) );
  OR U5902 ( .A(n5165), .B(n5164), .Z(n5167) );
  XOR U5903 ( .A(n4953), .B(n4952), .Z(n5161) );
  NAND U5904 ( .A(a[34]), .B(b[42]), .Z(n5151) );
  NANDN U5905 ( .A(n5151), .B(n5150), .Z(n5153) );
  XNOR U5906 ( .A(n4957), .B(n4956), .Z(n5147) );
  ANDN U5907 ( .B(b[42]), .A(n182), .Z(n5143) );
  XOR U5908 ( .A(n4959), .B(n4958), .Z(n5142) );
  OR U5909 ( .A(n5143), .B(n5142), .Z(n5145) );
  XOR U5910 ( .A(n4961), .B(n4960), .Z(n5139) );
  NAND U5911 ( .A(a[29]), .B(b[42]), .Z(n5129) );
  NAND U5912 ( .A(a[28]), .B(b[42]), .Z(n5123) );
  NAND U5913 ( .A(a[27]), .B(b[42]), .Z(n4965) );
  NANDN U5914 ( .A(n4965), .B(n4964), .Z(n5119) );
  XOR U5915 ( .A(n4965), .B(n4964), .Z(n5271) );
  NAND U5916 ( .A(a[24]), .B(b[42]), .Z(n5101) );
  XOR U5917 ( .A(n4967), .B(n4966), .Z(n5097) );
  NAND U5918 ( .A(a[21]), .B(b[42]), .Z(n5087) );
  NANDN U5919 ( .A(n5087), .B(n5086), .Z(n5089) );
  XOR U5920 ( .A(n4971), .B(n4970), .Z(n5083) );
  NAND U5921 ( .A(a[19]), .B(b[42]), .Z(n5079) );
  XNOR U5922 ( .A(n4973), .B(n4972), .Z(n5078) );
  NANDN U5923 ( .A(n5079), .B(n5078), .Z(n5081) );
  XNOR U5924 ( .A(n4975), .B(n4974), .Z(n5075) );
  AND U5925 ( .A(a[17]), .B(b[42]), .Z(n4978) );
  NANDN U5926 ( .A(n4979), .B(n4978), .Z(n5073) );
  XOR U5927 ( .A(n4979), .B(n4978), .Z(n5284) );
  NAND U5928 ( .A(a[16]), .B(b[42]), .Z(n5066) );
  NAND U5929 ( .A(a[15]), .B(b[42]), .Z(n5063) );
  XNOR U5930 ( .A(n4981), .B(n4980), .Z(n5062) );
  NANDN U5931 ( .A(n5063), .B(n5062), .Z(n5065) );
  NAND U5932 ( .A(a[13]), .B(b[42]), .Z(n5053) );
  XOR U5933 ( .A(n4983), .B(n4982), .Z(n5052) );
  NANDN U5934 ( .A(n5053), .B(n5052), .Z(n5055) );
  XNOR U5935 ( .A(n4985), .B(n4984), .Z(n5048) );
  XNOR U5936 ( .A(n4987), .B(n4986), .Z(n5044) );
  XOR U5937 ( .A(n4989), .B(n4988), .Z(n5040) );
  XNOR U5938 ( .A(n4991), .B(n4990), .Z(n5031) );
  XOR U5939 ( .A(n4993), .B(n4992), .Z(n4995) );
  AND U5940 ( .A(a[7]), .B(b[42]), .Z(n4994) );
  NANDN U5941 ( .A(n4995), .B(n4994), .Z(n5029) );
  XOR U5942 ( .A(n4995), .B(n4994), .Z(n5300) );
  XNOR U5943 ( .A(n4997), .B(n4996), .Z(n5019) );
  XNOR U5944 ( .A(n4999), .B(n4998), .Z(n5014) );
  XNOR U5945 ( .A(n5001), .B(n5000), .Z(n5010) );
  NAND U5946 ( .A(b[43]), .B(a[1]), .Z(n5003) );
  NAND U5947 ( .A(n5003), .B(n5002), .Z(n5006) );
  NANDN U5948 ( .A(n155), .B(a[0]), .Z(n5892) );
  OR U5949 ( .A(n5003), .B(n5892), .Z(n5315) );
  NANDN U5950 ( .A(n5005), .B(n5315), .Z(n5004) );
  AND U5951 ( .A(n5006), .B(n5004), .Z(n5009) );
  XNOR U5952 ( .A(n5315), .B(n5005), .Z(n5007) );
  NAND U5953 ( .A(n5007), .B(n5006), .Z(n5311) );
  ANDN U5954 ( .B(b[42]), .A(n162), .Z(n5310) );
  OR U5955 ( .A(n5311), .B(n5310), .Z(n5008) );
  AND U5956 ( .A(n5009), .B(n5008), .Z(n5011) );
  OR U5957 ( .A(n5010), .B(n5011), .Z(n5013) );
  XNOR U5958 ( .A(n5011), .B(n5010), .Z(n5308) );
  ANDN U5959 ( .B(b[42]), .A(n21580), .Z(n5309) );
  OR U5960 ( .A(n5308), .B(n5309), .Z(n5012) );
  AND U5961 ( .A(n5013), .B(n5012), .Z(n5015) );
  OR U5962 ( .A(n5014), .B(n5015), .Z(n5017) );
  XNOR U5963 ( .A(n5015), .B(n5014), .Z(n5306) );
  ANDN U5964 ( .B(b[42]), .A(n163), .Z(n5307) );
  OR U5965 ( .A(n5306), .B(n5307), .Z(n5016) );
  AND U5966 ( .A(n5017), .B(n5016), .Z(n5018) );
  OR U5967 ( .A(n5019), .B(n5018), .Z(n5021) );
  XNOR U5968 ( .A(n5019), .B(n5018), .Z(n5334) );
  NAND U5969 ( .A(b[42]), .B(a[5]), .Z(n5335) );
  NANDN U5970 ( .A(n5334), .B(n5335), .Z(n5020) );
  NAND U5971 ( .A(n5021), .B(n5020), .Z(n5023) );
  AND U5972 ( .A(a[6]), .B(b[42]), .Z(n5022) );
  NANDN U5973 ( .A(n5023), .B(n5022), .Z(n5027) );
  XOR U5974 ( .A(n5023), .B(n5022), .Z(n5302) );
  XOR U5975 ( .A(n5025), .B(n5024), .Z(n5303) );
  NANDN U5976 ( .A(n5302), .B(n5303), .Z(n5026) );
  AND U5977 ( .A(n5027), .B(n5026), .Z(n5301) );
  OR U5978 ( .A(n5300), .B(n5301), .Z(n5028) );
  AND U5979 ( .A(n5029), .B(n5028), .Z(n5030) );
  OR U5980 ( .A(n5031), .B(n5030), .Z(n5033) );
  XNOR U5981 ( .A(n5031), .B(n5030), .Z(n5345) );
  NAND U5982 ( .A(a[8]), .B(b[42]), .Z(n5344) );
  OR U5983 ( .A(n5345), .B(n5344), .Z(n5032) );
  NAND U5984 ( .A(n5033), .B(n5032), .Z(n5036) );
  XOR U5985 ( .A(n5035), .B(n5034), .Z(n5037) );
  OR U5986 ( .A(n5036), .B(n5037), .Z(n5039) );
  ANDN U5987 ( .B(b[42]), .A(n21615), .Z(n5299) );
  XOR U5988 ( .A(n5037), .B(n5036), .Z(n5298) );
  NANDN U5989 ( .A(n5299), .B(n5298), .Z(n5038) );
  AND U5990 ( .A(n5039), .B(n5038), .Z(n5041) );
  OR U5991 ( .A(n5040), .B(n5041), .Z(n5043) );
  XNOR U5992 ( .A(n5041), .B(n5040), .Z(n5296) );
  ANDN U5993 ( .B(b[42]), .A(n168), .Z(n5297) );
  OR U5994 ( .A(n5296), .B(n5297), .Z(n5042) );
  AND U5995 ( .A(n5043), .B(n5042), .Z(n5045) );
  OR U5996 ( .A(n5044), .B(n5045), .Z(n5047) );
  XNOR U5997 ( .A(n5045), .B(n5044), .Z(n5292) );
  ANDN U5998 ( .B(b[42]), .A(n21164), .Z(n5293) );
  OR U5999 ( .A(n5292), .B(n5293), .Z(n5046) );
  AND U6000 ( .A(n5047), .B(n5046), .Z(n5049) );
  OR U6001 ( .A(n5048), .B(n5049), .Z(n5051) );
  XNOR U6002 ( .A(n5049), .B(n5048), .Z(n5291) );
  ANDN U6003 ( .B(b[42]), .A(n169), .Z(n5290) );
  OR U6004 ( .A(n5291), .B(n5290), .Z(n5050) );
  NAND U6005 ( .A(n5051), .B(n5050), .Z(n5365) );
  NANDN U6006 ( .A(n5365), .B(n5364), .Z(n5054) );
  AND U6007 ( .A(n5055), .B(n5054), .Z(n5058) );
  NANDN U6008 ( .A(n5058), .B(n5059), .Z(n5061) );
  XOR U6009 ( .A(n5059), .B(n5058), .Z(n5371) );
  AND U6010 ( .A(a[14]), .B(b[42]), .Z(n5370) );
  NANDN U6011 ( .A(n5371), .B(n5370), .Z(n5060) );
  AND U6012 ( .A(n5061), .B(n5060), .Z(n5376) );
  NANDN U6013 ( .A(n5376), .B(n5377), .Z(n5064) );
  AND U6014 ( .A(n5065), .B(n5064), .Z(n5067) );
  OR U6015 ( .A(n5066), .B(n5067), .Z(n5071) );
  XNOR U6016 ( .A(n5067), .B(n5066), .Z(n5287) );
  XNOR U6017 ( .A(n5069), .B(n5068), .Z(n5286) );
  NANDN U6018 ( .A(n5287), .B(n5286), .Z(n5070) );
  AND U6019 ( .A(n5071), .B(n5070), .Z(n5285) );
  OR U6020 ( .A(n5284), .B(n5285), .Z(n5072) );
  AND U6021 ( .A(n5073), .B(n5072), .Z(n5074) );
  OR U6022 ( .A(n5075), .B(n5074), .Z(n5077) );
  XNOR U6023 ( .A(n5075), .B(n5074), .Z(n5283) );
  AND U6024 ( .A(a[18]), .B(b[42]), .Z(n5282) );
  NANDN U6025 ( .A(n5283), .B(n5282), .Z(n5076) );
  AND U6026 ( .A(n5077), .B(n5076), .Z(n5280) );
  NANDN U6027 ( .A(n5280), .B(n5281), .Z(n5080) );
  AND U6028 ( .A(n5081), .B(n5080), .Z(n5082) );
  OR U6029 ( .A(n5083), .B(n5082), .Z(n5085) );
  NAND U6030 ( .A(a[20]), .B(b[42]), .Z(n5397) );
  XNOR U6031 ( .A(n5083), .B(n5082), .Z(n5396) );
  OR U6032 ( .A(n5397), .B(n5396), .Z(n5084) );
  AND U6033 ( .A(n5085), .B(n5084), .Z(n5278) );
  NANDN U6034 ( .A(n5278), .B(n5279), .Z(n5088) );
  AND U6035 ( .A(n5089), .B(n5088), .Z(n5093) );
  XOR U6036 ( .A(n5091), .B(n5090), .Z(n5092) );
  NANDN U6037 ( .A(n5093), .B(n5092), .Z(n5095) );
  XOR U6038 ( .A(n5093), .B(n5092), .Z(n5407) );
  NAND U6039 ( .A(a[22]), .B(b[42]), .Z(n5406) );
  OR U6040 ( .A(n5407), .B(n5406), .Z(n5094) );
  AND U6041 ( .A(n5095), .B(n5094), .Z(n5096) );
  OR U6042 ( .A(n5097), .B(n5096), .Z(n5099) );
  NAND U6043 ( .A(a[23]), .B(b[42]), .Z(n5413) );
  XOR U6044 ( .A(n5097), .B(n5096), .Z(n5412) );
  NANDN U6045 ( .A(n5413), .B(n5412), .Z(n5098) );
  NAND U6046 ( .A(n5099), .B(n5098), .Z(n5100) );
  NANDN U6047 ( .A(n5101), .B(n5100), .Z(n5105) );
  XNOR U6048 ( .A(n5103), .B(n5102), .Z(n5421) );
  NAND U6049 ( .A(n5420), .B(n5421), .Z(n5104) );
  NAND U6050 ( .A(n5105), .B(n5104), .Z(n5109) );
  XOR U6051 ( .A(n5107), .B(n5106), .Z(n5108) );
  NANDN U6052 ( .A(n5109), .B(n5108), .Z(n5111) );
  ANDN U6053 ( .B(b[42]), .A(n21703), .Z(n5277) );
  XOR U6054 ( .A(n5109), .B(n5108), .Z(n5276) );
  OR U6055 ( .A(n5277), .B(n5276), .Z(n5110) );
  NAND U6056 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U6057 ( .A(n5115), .B(n5114), .Z(n5117) );
  NAND U6058 ( .A(a[26]), .B(b[42]), .Z(n5273) );
  XNOR U6059 ( .A(n5115), .B(n5114), .Z(n5272) );
  NANDN U6060 ( .A(n5273), .B(n5272), .Z(n5116) );
  NAND U6061 ( .A(n5117), .B(n5116), .Z(n5270) );
  NANDN U6062 ( .A(n5271), .B(n5270), .Z(n5118) );
  NAND U6063 ( .A(n5119), .B(n5118), .Z(n5122) );
  NANDN U6064 ( .A(n5123), .B(n5122), .Z(n5125) );
  XOR U6065 ( .A(n5121), .B(n5120), .Z(n5435) );
  NANDN U6066 ( .A(n5435), .B(n5434), .Z(n5124) );
  NAND U6067 ( .A(n5125), .B(n5124), .Z(n5128) );
  NANDN U6068 ( .A(n5129), .B(n5128), .Z(n5131) );
  XOR U6069 ( .A(n5127), .B(n5126), .Z(n5268) );
  NAND U6070 ( .A(n5268), .B(n5269), .Z(n5130) );
  NAND U6071 ( .A(n5131), .B(n5130), .Z(n5135) );
  XOR U6072 ( .A(n5133), .B(n5132), .Z(n5134) );
  NANDN U6073 ( .A(n5135), .B(n5134), .Z(n5137) );
  ANDN U6074 ( .B(b[42]), .A(n181), .Z(n5267) );
  NANDN U6075 ( .A(n5267), .B(n5266), .Z(n5136) );
  NAND U6076 ( .A(n5137), .B(n5136), .Z(n5138) );
  NANDN U6077 ( .A(n5139), .B(n5138), .Z(n5141) );
  ANDN U6078 ( .B(b[42]), .A(n21740), .Z(n5265) );
  NANDN U6079 ( .A(n5265), .B(n5264), .Z(n5140) );
  NAND U6080 ( .A(n5141), .B(n5140), .Z(n5262) );
  XOR U6081 ( .A(n5143), .B(n5142), .Z(n5263) );
  NAND U6082 ( .A(n5262), .B(n5263), .Z(n5144) );
  NAND U6083 ( .A(n5145), .B(n5144), .Z(n5146) );
  NANDN U6084 ( .A(n5147), .B(n5146), .Z(n5149) );
  ANDN U6085 ( .B(b[42]), .A(n21751), .Z(n5261) );
  NANDN U6086 ( .A(n5261), .B(n5260), .Z(n5148) );
  NAND U6087 ( .A(n5149), .B(n5148), .Z(n5259) );
  XNOR U6088 ( .A(n5151), .B(n5150), .Z(n5258) );
  NANDN U6089 ( .A(n5259), .B(n5258), .Z(n5152) );
  NAND U6090 ( .A(n5153), .B(n5152), .Z(n5157) );
  XOR U6091 ( .A(n5155), .B(n5154), .Z(n5156) );
  NANDN U6092 ( .A(n5157), .B(n5156), .Z(n5159) );
  ANDN U6093 ( .B(b[42]), .A(n184), .Z(n5257) );
  XOR U6094 ( .A(n5157), .B(n5156), .Z(n5256) );
  OR U6095 ( .A(n5257), .B(n5256), .Z(n5158) );
  NAND U6096 ( .A(n5159), .B(n5158), .Z(n5160) );
  NANDN U6097 ( .A(n5161), .B(n5160), .Z(n5163) );
  ANDN U6098 ( .B(b[42]), .A(n185), .Z(n5255) );
  NANDN U6099 ( .A(n5255), .B(n5254), .Z(n5162) );
  NAND U6100 ( .A(n5163), .B(n5162), .Z(n5252) );
  XOR U6101 ( .A(n5165), .B(n5164), .Z(n5253) );
  NAND U6102 ( .A(n5252), .B(n5253), .Z(n5166) );
  NAND U6103 ( .A(n5167), .B(n5166), .Z(n5169) );
  NANDN U6104 ( .A(n5168), .B(n5169), .Z(n5171) );
  ANDN U6105 ( .B(b[42]), .A(n186), .Z(n5477) );
  XOR U6106 ( .A(n5169), .B(n5168), .Z(n5476) );
  OR U6107 ( .A(n5477), .B(n5476), .Z(n5170) );
  NAND U6108 ( .A(n5171), .B(n5170), .Z(n5172) );
  NANDN U6109 ( .A(n5173), .B(n5172), .Z(n5175) );
  ANDN U6110 ( .B(b[42]), .A(n187), .Z(n5251) );
  NANDN U6111 ( .A(n5251), .B(n5250), .Z(n5174) );
  NAND U6112 ( .A(n5175), .B(n5174), .Z(n5176) );
  NANDN U6113 ( .A(n5177), .B(n5176), .Z(n5179) );
  ANDN U6114 ( .B(b[42]), .A(n188), .Z(n5247) );
  NANDN U6115 ( .A(n5247), .B(n5246), .Z(n5178) );
  NAND U6116 ( .A(n5179), .B(n5178), .Z(n5180) );
  NANDN U6117 ( .A(n5181), .B(n5180), .Z(n5183) );
  ANDN U6118 ( .B(b[42]), .A(n189), .Z(n5245) );
  NANDN U6119 ( .A(n5245), .B(n5244), .Z(n5182) );
  NAND U6120 ( .A(n5183), .B(n5182), .Z(n5241) );
  XNOR U6121 ( .A(n5185), .B(n5184), .Z(n5240) );
  NANDN U6122 ( .A(n5241), .B(n5240), .Z(n5186) );
  NAND U6123 ( .A(n5187), .B(n5186), .Z(n5191) );
  XOR U6124 ( .A(n5189), .B(n5188), .Z(n5190) );
  NANDN U6125 ( .A(n5191), .B(n5190), .Z(n5193) );
  ANDN U6126 ( .B(b[42]), .A(n191), .Z(n5239) );
  NANDN U6127 ( .A(n5239), .B(n5238), .Z(n5192) );
  NAND U6128 ( .A(n5193), .B(n5192), .Z(n5194) );
  NANDN U6129 ( .A(n5195), .B(n5194), .Z(n5197) );
  ANDN U6130 ( .B(b[42]), .A(n192), .Z(n5237) );
  NANDN U6131 ( .A(n5237), .B(n5236), .Z(n5196) );
  NAND U6132 ( .A(n5197), .B(n5196), .Z(n5198) );
  NANDN U6133 ( .A(n5199), .B(n5198), .Z(n5201) );
  ANDN U6134 ( .B(b[42]), .A(n193), .Z(n5503) );
  NANDN U6135 ( .A(n5503), .B(n5502), .Z(n5200) );
  NAND U6136 ( .A(n5201), .B(n5200), .Z(n5202) );
  NANDN U6137 ( .A(n5203), .B(n5202), .Z(n5205) );
  ANDN U6138 ( .B(b[42]), .A(n194), .Z(n5509) );
  NANDN U6139 ( .A(n5509), .B(n5508), .Z(n5204) );
  NAND U6140 ( .A(n5205), .B(n5204), .Z(n5206) );
  NANDN U6141 ( .A(n5207), .B(n5206), .Z(n5209) );
  NANDN U6142 ( .A(n155), .B(a[47]), .Z(n5235) );
  NAND U6143 ( .A(n5234), .B(n5235), .Z(n5208) );
  AND U6144 ( .A(n5209), .B(n5208), .Z(n5211) );
  OR U6145 ( .A(n5210), .B(n5211), .Z(n5213) );
  XNOR U6146 ( .A(n5211), .B(n5210), .Z(n5230) );
  NAND U6147 ( .A(b[42]), .B(a[48]), .Z(n5231) );
  NANDN U6148 ( .A(n5230), .B(n5231), .Z(n5212) );
  AND U6149 ( .A(n5213), .B(n5212), .Z(n5215) );
  OR U6150 ( .A(n5214), .B(n5215), .Z(n5217) );
  XNOR U6151 ( .A(n5215), .B(n5214), .Z(n5520) );
  ANDN U6152 ( .B(b[42]), .A(n197), .Z(n5521) );
  OR U6153 ( .A(n5520), .B(n5521), .Z(n5216) );
  AND U6154 ( .A(n5217), .B(n5216), .Z(n5219) );
  OR U6155 ( .A(n5218), .B(n5219), .Z(n5221) );
  XNOR U6156 ( .A(n5219), .B(n5218), .Z(n5228) );
  ANDN U6157 ( .B(b[42]), .A(n198), .Z(n5229) );
  OR U6158 ( .A(n5228), .B(n5229), .Z(n5220) );
  AND U6159 ( .A(n5221), .B(n5220), .Z(n5225) );
  NANDN U6160 ( .A(n5225), .B(n5224), .Z(n5227) );
  NAND U6161 ( .A(b[42]), .B(a[51]), .Z(n5531) );
  NAND U6162 ( .A(n5530), .B(n5531), .Z(n5226) );
  AND U6163 ( .A(n5227), .B(n5226), .Z(n5543) );
  XOR U6164 ( .A(n5542), .B(n5543), .Z(n5545) );
  NANDN U6165 ( .A(n5537), .B(n5536), .Z(n5539) );
  XNOR U6166 ( .A(n5229), .B(n5228), .Z(n5526) );
  NAND U6167 ( .A(a[49]), .B(b[41]), .Z(n5233) );
  XOR U6168 ( .A(n5231), .B(n5230), .Z(n5232) );
  NANDN U6169 ( .A(n5233), .B(n5232), .Z(n5519) );
  XOR U6170 ( .A(n5233), .B(n5232), .Z(n5807) );
  NAND U6171 ( .A(a[48]), .B(b[41]), .Z(n5514) );
  OR U6172 ( .A(n5515), .B(n5514), .Z(n5517) );
  NAND U6173 ( .A(a[45]), .B(b[41]), .Z(n5499) );
  NANDN U6174 ( .A(n5499), .B(n5498), .Z(n5501) );
  XOR U6175 ( .A(n5239), .B(n5238), .Z(n5495) );
  NAND U6176 ( .A(a[43]), .B(b[41]), .Z(n5243) );
  XNOR U6177 ( .A(n5241), .B(n5240), .Z(n5242) );
  NANDN U6178 ( .A(n5243), .B(n5242), .Z(n5493) );
  XOR U6179 ( .A(n5243), .B(n5242), .Z(n5818) );
  ANDN U6180 ( .B(b[41]), .A(n190), .Z(n5488) );
  XOR U6181 ( .A(n5245), .B(n5244), .Z(n5489) );
  OR U6182 ( .A(n5488), .B(n5489), .Z(n5491) );
  NAND U6183 ( .A(a[41]), .B(b[41]), .Z(n5249) );
  NANDN U6184 ( .A(n5249), .B(n5248), .Z(n5487) );
  XOR U6185 ( .A(n5249), .B(n5248), .Z(n5821) );
  XNOR U6186 ( .A(n5251), .B(n5250), .Z(n5483) );
  XNOR U6187 ( .A(n5253), .B(n5252), .Z(n5473) );
  XNOR U6188 ( .A(n5255), .B(n5254), .Z(n5469) );
  NAND U6189 ( .A(a[36]), .B(b[41]), .Z(n5465) );
  XNOR U6190 ( .A(n5257), .B(n5256), .Z(n5464) );
  NANDN U6191 ( .A(n5465), .B(n5464), .Z(n5467) );
  NAND U6192 ( .A(b[41]), .B(a[35]), .Z(n5460) );
  XNOR U6193 ( .A(n5259), .B(n5258), .Z(n5461) );
  NANDN U6194 ( .A(n5460), .B(n5461), .Z(n5463) );
  XOR U6195 ( .A(n5261), .B(n5260), .Z(n5457) );
  XNOR U6196 ( .A(n5263), .B(n5262), .Z(n5453) );
  XOR U6197 ( .A(n5265), .B(n5264), .Z(n5449) );
  XOR U6198 ( .A(n5267), .B(n5266), .Z(n5445) );
  XOR U6199 ( .A(n5271), .B(n5270), .Z(n5431) );
  NAND U6200 ( .A(a[27]), .B(b[41]), .Z(n5275) );
  XNOR U6201 ( .A(n5273), .B(n5272), .Z(n5274) );
  NANDN U6202 ( .A(n5275), .B(n5274), .Z(n5429) );
  XOR U6203 ( .A(n5275), .B(n5274), .Z(n5847) );
  ANDN U6204 ( .B(b[41]), .A(n179), .Z(n5424) );
  XNOR U6205 ( .A(n5277), .B(n5276), .Z(n5425) );
  OR U6206 ( .A(n5424), .B(n5425), .Z(n5427) );
  NAND U6207 ( .A(a[25]), .B(b[41]), .Z(n5419) );
  NAND U6208 ( .A(a[24]), .B(b[41]), .Z(n5415) );
  XOR U6209 ( .A(n5279), .B(n5278), .Z(n5403) );
  XOR U6210 ( .A(n5281), .B(n5280), .Z(n5393) );
  NAND U6211 ( .A(a[19]), .B(b[41]), .Z(n5389) );
  XNOR U6212 ( .A(n5283), .B(n5282), .Z(n5388) );
  NANDN U6213 ( .A(n5389), .B(n5388), .Z(n5391) );
  XNOR U6214 ( .A(n5285), .B(n5284), .Z(n5385) );
  AND U6215 ( .A(a[17]), .B(b[41]), .Z(n5288) );
  NANDN U6216 ( .A(n5289), .B(n5288), .Z(n5383) );
  XOR U6217 ( .A(n5289), .B(n5288), .Z(n5864) );
  NAND U6218 ( .A(a[16]), .B(b[41]), .Z(n5378) );
  NAND U6219 ( .A(a[13]), .B(b[41]), .Z(n5360) );
  XOR U6220 ( .A(n5291), .B(n5290), .Z(n5361) );
  OR U6221 ( .A(n5360), .B(n5361), .Z(n5363) );
  XNOR U6222 ( .A(n5293), .B(n5292), .Z(n5294) );
  ANDN U6223 ( .B(b[41]), .A(n169), .Z(n5295) );
  OR U6224 ( .A(n5294), .B(n5295), .Z(n5359) );
  XNOR U6225 ( .A(n5295), .B(n5294), .Z(n5871) );
  XNOR U6226 ( .A(n5297), .B(n5296), .Z(n5354) );
  XOR U6227 ( .A(n5299), .B(n5298), .Z(n5350) );
  XNOR U6228 ( .A(n5301), .B(n5300), .Z(n5341) );
  XOR U6229 ( .A(n5303), .B(n5302), .Z(n5305) );
  AND U6230 ( .A(a[7]), .B(b[41]), .Z(n5304) );
  NANDN U6231 ( .A(n5305), .B(n5304), .Z(n5339) );
  XOR U6232 ( .A(n5305), .B(n5304), .Z(n5880) );
  XNOR U6233 ( .A(n5307), .B(n5306), .Z(n5329) );
  XNOR U6234 ( .A(n5309), .B(n5308), .Z(n5324) );
  XNOR U6235 ( .A(n5311), .B(n5310), .Z(n5320) );
  NAND U6236 ( .A(b[42]), .B(a[1]), .Z(n5313) );
  NAND U6237 ( .A(n5313), .B(n5312), .Z(n5316) );
  OR U6238 ( .A(n5313), .B(n6336), .Z(n5895) );
  NANDN U6239 ( .A(n5315), .B(n5895), .Z(n5314) );
  AND U6240 ( .A(n5316), .B(n5314), .Z(n5319) );
  XNOR U6241 ( .A(n5895), .B(n5315), .Z(n5317) );
  NAND U6242 ( .A(n5317), .B(n5316), .Z(n5891) );
  ANDN U6243 ( .B(b[41]), .A(n162), .Z(n5890) );
  OR U6244 ( .A(n5891), .B(n5890), .Z(n5318) );
  AND U6245 ( .A(n5319), .B(n5318), .Z(n5321) );
  OR U6246 ( .A(n5320), .B(n5321), .Z(n5323) );
  XNOR U6247 ( .A(n5321), .B(n5320), .Z(n5888) );
  ANDN U6248 ( .B(b[41]), .A(n21580), .Z(n5889) );
  OR U6249 ( .A(n5888), .B(n5889), .Z(n5322) );
  AND U6250 ( .A(n5323), .B(n5322), .Z(n5325) );
  OR U6251 ( .A(n5324), .B(n5325), .Z(n5327) );
  XNOR U6252 ( .A(n5325), .B(n5324), .Z(n5886) );
  ANDN U6253 ( .B(b[41]), .A(n163), .Z(n5887) );
  OR U6254 ( .A(n5886), .B(n5887), .Z(n5326) );
  AND U6255 ( .A(n5327), .B(n5326), .Z(n5328) );
  OR U6256 ( .A(n5329), .B(n5328), .Z(n5331) );
  XNOR U6257 ( .A(n5329), .B(n5328), .Z(n5914) );
  NAND U6258 ( .A(b[41]), .B(a[5]), .Z(n5915) );
  NANDN U6259 ( .A(n5914), .B(n5915), .Z(n5330) );
  NAND U6260 ( .A(n5331), .B(n5330), .Z(n5333) );
  AND U6261 ( .A(a[6]), .B(b[41]), .Z(n5332) );
  NANDN U6262 ( .A(n5333), .B(n5332), .Z(n5337) );
  XOR U6263 ( .A(n5333), .B(n5332), .Z(n5882) );
  XOR U6264 ( .A(n5335), .B(n5334), .Z(n5883) );
  NANDN U6265 ( .A(n5882), .B(n5883), .Z(n5336) );
  AND U6266 ( .A(n5337), .B(n5336), .Z(n5881) );
  OR U6267 ( .A(n5880), .B(n5881), .Z(n5338) );
  AND U6268 ( .A(n5339), .B(n5338), .Z(n5340) );
  OR U6269 ( .A(n5341), .B(n5340), .Z(n5343) );
  XNOR U6270 ( .A(n5341), .B(n5340), .Z(n5925) );
  NAND U6271 ( .A(a[8]), .B(b[41]), .Z(n5924) );
  OR U6272 ( .A(n5925), .B(n5924), .Z(n5342) );
  NAND U6273 ( .A(n5343), .B(n5342), .Z(n5346) );
  XOR U6274 ( .A(n5345), .B(n5344), .Z(n5347) );
  OR U6275 ( .A(n5346), .B(n5347), .Z(n5349) );
  ANDN U6276 ( .B(b[41]), .A(n21615), .Z(n5879) );
  XOR U6277 ( .A(n5347), .B(n5346), .Z(n5878) );
  NANDN U6278 ( .A(n5879), .B(n5878), .Z(n5348) );
  AND U6279 ( .A(n5349), .B(n5348), .Z(n5351) );
  OR U6280 ( .A(n5350), .B(n5351), .Z(n5353) );
  XNOR U6281 ( .A(n5351), .B(n5350), .Z(n5876) );
  ANDN U6282 ( .B(b[41]), .A(n168), .Z(n5877) );
  OR U6283 ( .A(n5876), .B(n5877), .Z(n5352) );
  AND U6284 ( .A(n5353), .B(n5352), .Z(n5355) );
  OR U6285 ( .A(n5354), .B(n5355), .Z(n5357) );
  XNOR U6286 ( .A(n5355), .B(n5354), .Z(n5872) );
  ANDN U6287 ( .B(b[41]), .A(n21164), .Z(n5873) );
  OR U6288 ( .A(n5872), .B(n5873), .Z(n5356) );
  AND U6289 ( .A(n5357), .B(n5356), .Z(n5870) );
  OR U6290 ( .A(n5871), .B(n5870), .Z(n5358) );
  NAND U6291 ( .A(n5359), .B(n5358), .Z(n5945) );
  XOR U6292 ( .A(n5361), .B(n5360), .Z(n5944) );
  NANDN U6293 ( .A(n5945), .B(n5944), .Z(n5362) );
  AND U6294 ( .A(n5363), .B(n5362), .Z(n5366) );
  NANDN U6295 ( .A(n5366), .B(n5367), .Z(n5369) );
  XOR U6296 ( .A(n5367), .B(n5366), .Z(n5951) );
  AND U6297 ( .A(a[14]), .B(b[41]), .Z(n5950) );
  NANDN U6298 ( .A(n5951), .B(n5950), .Z(n5368) );
  AND U6299 ( .A(n5369), .B(n5368), .Z(n5373) );
  XNOR U6300 ( .A(n5371), .B(n5370), .Z(n5372) );
  NANDN U6301 ( .A(n5373), .B(n5372), .Z(n5375) );
  NAND U6302 ( .A(a[15]), .B(b[41]), .Z(n5959) );
  NANDN U6303 ( .A(n5959), .B(n5958), .Z(n5374) );
  AND U6304 ( .A(n5375), .B(n5374), .Z(n5379) );
  OR U6305 ( .A(n5378), .B(n5379), .Z(n5381) );
  XOR U6306 ( .A(n5377), .B(n5376), .Z(n5867) );
  XNOR U6307 ( .A(n5379), .B(n5378), .Z(n5866) );
  OR U6308 ( .A(n5867), .B(n5866), .Z(n5380) );
  AND U6309 ( .A(n5381), .B(n5380), .Z(n5865) );
  OR U6310 ( .A(n5864), .B(n5865), .Z(n5382) );
  AND U6311 ( .A(n5383), .B(n5382), .Z(n5384) );
  OR U6312 ( .A(n5385), .B(n5384), .Z(n5387) );
  XNOR U6313 ( .A(n5385), .B(n5384), .Z(n5969) );
  AND U6314 ( .A(a[18]), .B(b[41]), .Z(n5968) );
  NANDN U6315 ( .A(n5969), .B(n5968), .Z(n5386) );
  AND U6316 ( .A(n5387), .B(n5386), .Z(n5862) );
  NANDN U6317 ( .A(n5862), .B(n5863), .Z(n5390) );
  AND U6318 ( .A(n5391), .B(n5390), .Z(n5392) );
  OR U6319 ( .A(n5393), .B(n5392), .Z(n5395) );
  NAND U6320 ( .A(a[20]), .B(b[41]), .Z(n5979) );
  XNOR U6321 ( .A(n5393), .B(n5392), .Z(n5978) );
  OR U6322 ( .A(n5979), .B(n5978), .Z(n5394) );
  NAND U6323 ( .A(n5395), .B(n5394), .Z(n5398) );
  XOR U6324 ( .A(n5397), .B(n5396), .Z(n5399) );
  OR U6325 ( .A(n5398), .B(n5399), .Z(n5401) );
  ANDN U6326 ( .B(b[41]), .A(n21681), .Z(n5861) );
  XOR U6327 ( .A(n5399), .B(n5398), .Z(n5860) );
  NANDN U6328 ( .A(n5861), .B(n5860), .Z(n5400) );
  NAND U6329 ( .A(n5401), .B(n5400), .Z(n5402) );
  OR U6330 ( .A(n5403), .B(n5402), .Z(n5405) );
  NAND U6331 ( .A(a[22]), .B(b[41]), .Z(n5859) );
  XNOR U6332 ( .A(n5403), .B(n5402), .Z(n5858) );
  OR U6333 ( .A(n5859), .B(n5858), .Z(n5404) );
  NAND U6334 ( .A(n5405), .B(n5404), .Z(n5408) );
  XOR U6335 ( .A(n5407), .B(n5406), .Z(n5409) );
  OR U6336 ( .A(n5408), .B(n5409), .Z(n5411) );
  ANDN U6337 ( .B(b[41]), .A(n21692), .Z(n5856) );
  XOR U6338 ( .A(n5409), .B(n5408), .Z(n5857) );
  NANDN U6339 ( .A(n5856), .B(n5857), .Z(n5410) );
  AND U6340 ( .A(n5411), .B(n5410), .Z(n5414) );
  NANDN U6341 ( .A(n5415), .B(n5414), .Z(n5417) );
  XOR U6342 ( .A(n5413), .B(n5412), .Z(n5855) );
  NANDN U6343 ( .A(n5855), .B(n5854), .Z(n5416) );
  NAND U6344 ( .A(n5417), .B(n5416), .Z(n5418) );
  NANDN U6345 ( .A(n5419), .B(n5418), .Z(n5423) );
  NAND U6346 ( .A(n5850), .B(n5851), .Z(n5422) );
  AND U6347 ( .A(n5423), .B(n5422), .Z(n5848) );
  XOR U6348 ( .A(n5425), .B(n5424), .Z(n5849) );
  NAND U6349 ( .A(n5848), .B(n5849), .Z(n5426) );
  NAND U6350 ( .A(n5427), .B(n5426), .Z(n5846) );
  OR U6351 ( .A(n5847), .B(n5846), .Z(n5428) );
  NAND U6352 ( .A(n5429), .B(n5428), .Z(n5430) );
  NANDN U6353 ( .A(n5431), .B(n5430), .Z(n5433) );
  NAND U6354 ( .A(a[28]), .B(b[41]), .Z(n5844) );
  NANDN U6355 ( .A(n5844), .B(n5845), .Z(n5432) );
  NAND U6356 ( .A(n5433), .B(n5432), .Z(n5436) );
  XNOR U6357 ( .A(n5435), .B(n5434), .Z(n5437) );
  NAND U6358 ( .A(n5436), .B(n5437), .Z(n5439) );
  XNOR U6359 ( .A(n5437), .B(n5436), .Z(n5843) );
  NAND U6360 ( .A(a[29]), .B(b[41]), .Z(n5842) );
  OR U6361 ( .A(n5843), .B(n5842), .Z(n5438) );
  NAND U6362 ( .A(n5439), .B(n5438), .Z(n5440) );
  OR U6363 ( .A(n5441), .B(n5440), .Z(n5443) );
  ANDN U6364 ( .B(b[41]), .A(n181), .Z(n5841) );
  XOR U6365 ( .A(n5441), .B(n5440), .Z(n5840) );
  NANDN U6366 ( .A(n5841), .B(n5840), .Z(n5442) );
  NAND U6367 ( .A(n5443), .B(n5442), .Z(n5444) );
  NANDN U6368 ( .A(n5445), .B(n5444), .Z(n5447) );
  ANDN U6369 ( .B(b[41]), .A(n21740), .Z(n5837) );
  NANDN U6370 ( .A(n5837), .B(n5836), .Z(n5446) );
  NAND U6371 ( .A(n5447), .B(n5446), .Z(n5448) );
  NANDN U6372 ( .A(n5449), .B(n5448), .Z(n5451) );
  ANDN U6373 ( .B(b[41]), .A(n182), .Z(n6025) );
  NANDN U6374 ( .A(n6025), .B(n6024), .Z(n5450) );
  NAND U6375 ( .A(n5451), .B(n5450), .Z(n5452) );
  NANDN U6376 ( .A(n5453), .B(n5452), .Z(n5455) );
  ANDN U6377 ( .B(b[41]), .A(n21751), .Z(n5833) );
  NANDN U6378 ( .A(n5833), .B(n5832), .Z(n5454) );
  NAND U6379 ( .A(n5455), .B(n5454), .Z(n5456) );
  NANDN U6380 ( .A(n5457), .B(n5456), .Z(n5459) );
  ANDN U6381 ( .B(b[41]), .A(n183), .Z(n5831) );
  NANDN U6382 ( .A(n5831), .B(n5830), .Z(n5458) );
  NAND U6383 ( .A(n5459), .B(n5458), .Z(n6039) );
  XNOR U6384 ( .A(n5461), .B(n5460), .Z(n6038) );
  NANDN U6385 ( .A(n6039), .B(n6038), .Z(n5462) );
  AND U6386 ( .A(n5463), .B(n5462), .Z(n5826) );
  XNOR U6387 ( .A(n5465), .B(n5464), .Z(n5827) );
  NANDN U6388 ( .A(n5826), .B(n5827), .Z(n5466) );
  NAND U6389 ( .A(n5467), .B(n5466), .Z(n5468) );
  NANDN U6390 ( .A(n5469), .B(n5468), .Z(n5471) );
  NAND U6391 ( .A(a[37]), .B(b[41]), .Z(n6044) );
  NANDN U6392 ( .A(n6044), .B(n6045), .Z(n5470) );
  AND U6393 ( .A(n5471), .B(n5470), .Z(n5472) );
  NANDN U6394 ( .A(n5473), .B(n5472), .Z(n5475) );
  ANDN U6395 ( .B(b[41]), .A(n186), .Z(n5825) );
  NANDN U6396 ( .A(n5825), .B(n5824), .Z(n5474) );
  NAND U6397 ( .A(n5475), .B(n5474), .Z(n5479) );
  XNOR U6398 ( .A(n5477), .B(n5476), .Z(n5478) );
  NANDN U6399 ( .A(n5479), .B(n5478), .Z(n5481) );
  NAND U6400 ( .A(a[39]), .B(b[41]), .Z(n6055) );
  XNOR U6401 ( .A(n5479), .B(n5478), .Z(n6054) );
  NANDN U6402 ( .A(n6055), .B(n6054), .Z(n5480) );
  NAND U6403 ( .A(n5481), .B(n5480), .Z(n5482) );
  NANDN U6404 ( .A(n5483), .B(n5482), .Z(n5485) );
  NAND U6405 ( .A(a[40]), .B(b[41]), .Z(n5823) );
  NANDN U6406 ( .A(n5823), .B(n5822), .Z(n5484) );
  NAND U6407 ( .A(n5485), .B(n5484), .Z(n5820) );
  NANDN U6408 ( .A(n5821), .B(n5820), .Z(n5486) );
  NAND U6409 ( .A(n5487), .B(n5486), .Z(n6068) );
  XNOR U6410 ( .A(n5489), .B(n5488), .Z(n6069) );
  OR U6411 ( .A(n6068), .B(n6069), .Z(n5490) );
  NAND U6412 ( .A(n5491), .B(n5490), .Z(n5819) );
  OR U6413 ( .A(n5818), .B(n5819), .Z(n5492) );
  AND U6414 ( .A(n5493), .B(n5492), .Z(n5494) );
  NANDN U6415 ( .A(n5495), .B(n5494), .Z(n5497) );
  ANDN U6416 ( .B(b[41]), .A(n192), .Z(n5817) );
  NANDN U6417 ( .A(n5817), .B(n5816), .Z(n5496) );
  NAND U6418 ( .A(n5497), .B(n5496), .Z(n5813) );
  XNOR U6419 ( .A(n5499), .B(n5498), .Z(n5812) );
  NANDN U6420 ( .A(n5813), .B(n5812), .Z(n5500) );
  AND U6421 ( .A(n5501), .B(n5500), .Z(n5504) );
  NANDN U6422 ( .A(n5504), .B(n5505), .Z(n5507) );
  NAND U6423 ( .A(a[46]), .B(b[41]), .Z(n5811) );
  XNOR U6424 ( .A(n5505), .B(n5504), .Z(n5810) );
  NANDN U6425 ( .A(n5811), .B(n5810), .Z(n5506) );
  AND U6426 ( .A(n5507), .B(n5506), .Z(n5510) );
  NANDN U6427 ( .A(n5510), .B(n5511), .Z(n5513) );
  NAND U6428 ( .A(a[47]), .B(b[41]), .Z(n5809) );
  XNOR U6429 ( .A(n5511), .B(n5510), .Z(n5808) );
  NANDN U6430 ( .A(n5809), .B(n5808), .Z(n5512) );
  AND U6431 ( .A(n5513), .B(n5512), .Z(n6092) );
  XOR U6432 ( .A(n5515), .B(n5514), .Z(n6093) );
  NANDN U6433 ( .A(n6092), .B(n6093), .Z(n5516) );
  AND U6434 ( .A(n5517), .B(n5516), .Z(n5806) );
  OR U6435 ( .A(n5807), .B(n5806), .Z(n5518) );
  NAND U6436 ( .A(n5519), .B(n5518), .Z(n5523) );
  XOR U6437 ( .A(n5521), .B(n5520), .Z(n5522) );
  NANDN U6438 ( .A(n5523), .B(n5522), .Z(n5525) );
  ANDN U6439 ( .B(b[41]), .A(n198), .Z(n5805) );
  XOR U6440 ( .A(n5523), .B(n5522), .Z(n5804) );
  OR U6441 ( .A(n5805), .B(n5804), .Z(n5524) );
  AND U6442 ( .A(n5525), .B(n5524), .Z(n5527) );
  OR U6443 ( .A(n5526), .B(n5527), .Z(n5529) );
  XNOR U6444 ( .A(n5527), .B(n5526), .Z(n5800) );
  ANDN U6445 ( .B(b[41]), .A(n199), .Z(n5801) );
  OR U6446 ( .A(n5800), .B(n5801), .Z(n5528) );
  NAND U6447 ( .A(n5529), .B(n5528), .Z(n5533) );
  NANDN U6448 ( .A(n5533), .B(n5532), .Z(n5535) );
  NAND U6449 ( .A(a[52]), .B(b[41]), .Z(n6111) );
  NANDN U6450 ( .A(n6111), .B(n6110), .Z(n5534) );
  AND U6451 ( .A(n5535), .B(n5534), .Z(n6115) );
  NANDN U6452 ( .A(n6115), .B(n6114), .Z(n5538) );
  AND U6453 ( .A(n5539), .B(n5538), .Z(n5541) );
  OR U6454 ( .A(n5540), .B(n5541), .Z(n5669) );
  XNOR U6455 ( .A(n5541), .B(n5540), .Z(n5798) );
  OR U6456 ( .A(n5543), .B(n5542), .Z(n5547) );
  NAND U6457 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U6458 ( .A(n5547), .B(n5546), .Z(n5670) );
  NAND U6459 ( .A(a[52]), .B(b[43]), .Z(n5679) );
  NAND U6460 ( .A(a[51]), .B(b[44]), .Z(n5683) );
  NANDN U6461 ( .A(n5549), .B(n5548), .Z(n5553) );
  NANDN U6462 ( .A(n5551), .B(n5550), .Z(n5552) );
  NAND U6463 ( .A(n5553), .B(n5552), .Z(n5682) );
  XNOR U6464 ( .A(n5683), .B(n5682), .Z(n5685) );
  NAND U6465 ( .A(a[50]), .B(b[45]), .Z(n5793) );
  OR U6466 ( .A(n5555), .B(n5554), .Z(n5559) );
  OR U6467 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U6468 ( .A(n5559), .B(n5558), .Z(n5791) );
  ANDN U6469 ( .B(b[47]), .A(n196), .Z(n5690) );
  NANDN U6470 ( .A(n5561), .B(n5560), .Z(n5565) );
  NAND U6471 ( .A(n5563), .B(n5562), .Z(n5564) );
  AND U6472 ( .A(n5565), .B(n5564), .Z(n5689) );
  NAND U6473 ( .A(a[46]), .B(b[49]), .Z(n5697) );
  OR U6474 ( .A(n5567), .B(n5566), .Z(n5571) );
  NANDN U6475 ( .A(n5569), .B(n5568), .Z(n5570) );
  AND U6476 ( .A(n5571), .B(n5570), .Z(n5694) );
  NAND U6477 ( .A(a[44]), .B(b[51]), .Z(n5775) );
  OR U6478 ( .A(n5573), .B(n5572), .Z(n5577) );
  NANDN U6479 ( .A(n5575), .B(n5574), .Z(n5576) );
  NAND U6480 ( .A(n5577), .B(n5576), .Z(n5773) );
  NAND U6481 ( .A(a[42]), .B(b[53]), .Z(n5709) );
  OR U6482 ( .A(n5579), .B(n5578), .Z(n5583) );
  OR U6483 ( .A(n5581), .B(n5580), .Z(n5582) );
  AND U6484 ( .A(n5583), .B(n5582), .Z(n5706) );
  NAND U6485 ( .A(a[40]), .B(b[55]), .Z(n5763) );
  OR U6486 ( .A(n5585), .B(n5584), .Z(n5589) );
  OR U6487 ( .A(n5587), .B(n5586), .Z(n5588) );
  AND U6488 ( .A(n5589), .B(n5588), .Z(n5760) );
  NAND U6489 ( .A(a[38]), .B(b[57]), .Z(n5727) );
  OR U6490 ( .A(n5591), .B(n5590), .Z(n5595) );
  OR U6491 ( .A(n5593), .B(n5592), .Z(n5594) );
  NAND U6492 ( .A(n5595), .B(n5594), .Z(n5725) );
  NAND U6493 ( .A(a[36]), .B(b[59]), .Z(n5757) );
  NANDN U6494 ( .A(n5597), .B(n5596), .Z(n5601) );
  NAND U6495 ( .A(n5599), .B(n5598), .Z(n5600) );
  NAND U6496 ( .A(n5601), .B(n5600), .Z(n5755) );
  ANDN U6497 ( .B(b[61]), .A(n183), .Z(n5738) );
  OR U6498 ( .A(n5603), .B(n5602), .Z(n5607) );
  OR U6499 ( .A(n5605), .B(n5604), .Z(n5606) );
  AND U6500 ( .A(n5607), .B(n5606), .Z(n5736) );
  ANDN U6501 ( .B(b[63]), .A(n182), .Z(n5744) );
  ANDN U6502 ( .B(a[33]), .A(n159), .Z(n5742) );
  OR U6503 ( .A(n5609), .B(n5608), .Z(n5613) );
  OR U6504 ( .A(n5611), .B(n5610), .Z(n5612) );
  AND U6505 ( .A(n5613), .B(n5612), .Z(n5743) );
  XNOR U6506 ( .A(n5742), .B(n5743), .Z(n5745) );
  XNOR U6507 ( .A(n5744), .B(n5745), .Z(n5737) );
  XNOR U6508 ( .A(n5736), .B(n5737), .Z(n5739) );
  XNOR U6509 ( .A(n5738), .B(n5739), .Z(n5751) );
  ANDN U6510 ( .B(b[60]), .A(n184), .Z(n5748) );
  OR U6511 ( .A(n5615), .B(n5614), .Z(n5619) );
  NANDN U6512 ( .A(n5617), .B(n5616), .Z(n5618) );
  AND U6513 ( .A(n5619), .B(n5618), .Z(n5749) );
  XNOR U6514 ( .A(n5748), .B(n5749), .Z(n5750) );
  XOR U6515 ( .A(n5751), .B(n5750), .Z(n5754) );
  XOR U6516 ( .A(n5755), .B(n5754), .Z(n5756) );
  ANDN U6517 ( .B(b[58]), .A(n21772), .Z(n5730) );
  OR U6518 ( .A(n5621), .B(n5620), .Z(n5625) );
  NANDN U6519 ( .A(n5623), .B(n5622), .Z(n5624) );
  NAND U6520 ( .A(n5625), .B(n5624), .Z(n5731) );
  XOR U6521 ( .A(n5730), .B(n5731), .Z(n5732) );
  XNOR U6522 ( .A(n5733), .B(n5732), .Z(n5724) );
  XNOR U6523 ( .A(n5725), .B(n5724), .Z(n5726) );
  XOR U6524 ( .A(n5727), .B(n5726), .Z(n5721) );
  ANDN U6525 ( .B(b[56]), .A(n187), .Z(n5718) );
  OR U6526 ( .A(n5627), .B(n5626), .Z(n5631) );
  OR U6527 ( .A(n5629), .B(n5628), .Z(n5630) );
  AND U6528 ( .A(n5631), .B(n5630), .Z(n5719) );
  XOR U6529 ( .A(n5718), .B(n5719), .Z(n5720) );
  XNOR U6530 ( .A(n5721), .B(n5720), .Z(n5761) );
  XNOR U6531 ( .A(n5760), .B(n5761), .Z(n5762) );
  XOR U6532 ( .A(n5763), .B(n5762), .Z(n5715) );
  ANDN U6533 ( .B(b[54]), .A(n189), .Z(n5712) );
  OR U6534 ( .A(n5633), .B(n5632), .Z(n5637) );
  NANDN U6535 ( .A(n5635), .B(n5634), .Z(n5636) );
  AND U6536 ( .A(n5637), .B(n5636), .Z(n5713) );
  XOR U6537 ( .A(n5712), .B(n5713), .Z(n5714) );
  XNOR U6538 ( .A(n5715), .B(n5714), .Z(n5707) );
  XNOR U6539 ( .A(n5706), .B(n5707), .Z(n5708) );
  XOR U6540 ( .A(n5709), .B(n5708), .Z(n5769) );
  ANDN U6541 ( .B(b[52]), .A(n191), .Z(n5766) );
  OR U6542 ( .A(n5639), .B(n5638), .Z(n5643) );
  NANDN U6543 ( .A(n5641), .B(n5640), .Z(n5642) );
  NAND U6544 ( .A(n5643), .B(n5642), .Z(n5767) );
  XOR U6545 ( .A(n5766), .B(n5767), .Z(n5768) );
  XNOR U6546 ( .A(n5769), .B(n5768), .Z(n5772) );
  XNOR U6547 ( .A(n5773), .B(n5772), .Z(n5774) );
  XOR U6548 ( .A(n5775), .B(n5774), .Z(n5703) );
  ANDN U6549 ( .B(b[50]), .A(n193), .Z(n5700) );
  OR U6550 ( .A(n5645), .B(n5644), .Z(n5649) );
  OR U6551 ( .A(n5647), .B(n5646), .Z(n5648) );
  AND U6552 ( .A(n5649), .B(n5648), .Z(n5701) );
  XOR U6553 ( .A(n5700), .B(n5701), .Z(n5702) );
  XNOR U6554 ( .A(n5703), .B(n5702), .Z(n5695) );
  XNOR U6555 ( .A(n5694), .B(n5695), .Z(n5696) );
  XOR U6556 ( .A(n5697), .B(n5696), .Z(n5780) );
  ANDN U6557 ( .B(b[48]), .A(n195), .Z(n5778) );
  OR U6558 ( .A(n5651), .B(n5650), .Z(n5655) );
  OR U6559 ( .A(n5653), .B(n5652), .Z(n5654) );
  AND U6560 ( .A(n5655), .B(n5654), .Z(n5779) );
  XNOR U6561 ( .A(n5778), .B(n5779), .Z(n5781) );
  XOR U6562 ( .A(n5780), .B(n5781), .Z(n5688) );
  XOR U6563 ( .A(n5689), .B(n5688), .Z(n5691) );
  XNOR U6564 ( .A(n5690), .B(n5691), .Z(n5787) );
  ANDN U6565 ( .B(b[46]), .A(n197), .Z(n5784) );
  OR U6566 ( .A(n5657), .B(n5656), .Z(n5661) );
  NANDN U6567 ( .A(n5659), .B(n5658), .Z(n5660) );
  NAND U6568 ( .A(n5661), .B(n5660), .Z(n5785) );
  XNOR U6569 ( .A(n5784), .B(n5785), .Z(n5786) );
  XOR U6570 ( .A(n5787), .B(n5786), .Z(n5790) );
  XOR U6571 ( .A(n5791), .B(n5790), .Z(n5792) );
  NANDN U6572 ( .A(n5663), .B(n5662), .Z(n5667) );
  NANDN U6573 ( .A(n5665), .B(n5664), .Z(n5666) );
  AND U6574 ( .A(n5667), .B(n5666), .Z(n5677) );
  XOR U6575 ( .A(n5676), .B(n5677), .Z(n5678) );
  XOR U6576 ( .A(n5679), .B(n5678), .Z(n5671) );
  XNOR U6577 ( .A(n5670), .B(n5671), .Z(n5673) );
  ANDN U6578 ( .B(b[42]), .A(n201), .Z(n5672) );
  XOR U6579 ( .A(n5673), .B(n5672), .Z(n5799) );
  OR U6580 ( .A(n5798), .B(n5799), .Z(n5668) );
  NAND U6581 ( .A(n5669), .B(n5668), .Z(n6128) );
  OR U6582 ( .A(n5671), .B(n5670), .Z(n5675) );
  OR U6583 ( .A(n5673), .B(n5672), .Z(n5674) );
  AND U6584 ( .A(n5675), .B(n5674), .Z(n6252) );
  NANDN U6585 ( .A(n5677), .B(n5676), .Z(n5681) );
  OR U6586 ( .A(n5679), .B(n5678), .Z(n5680) );
  AND U6587 ( .A(n5681), .B(n5680), .Z(n6132) );
  ANDN U6588 ( .B(b[44]), .A(n200), .Z(n6246) );
  OR U6589 ( .A(n5683), .B(n5682), .Z(n5687) );
  NANDN U6590 ( .A(n5685), .B(n5684), .Z(n5686) );
  NAND U6591 ( .A(n5687), .B(n5686), .Z(n6247) );
  XNOR U6592 ( .A(n6246), .B(n6247), .Z(n6249) );
  ANDN U6593 ( .B(b[47]), .A(n197), .Z(n6146) );
  NANDN U6594 ( .A(n5689), .B(n5688), .Z(n5693) );
  OR U6595 ( .A(n5691), .B(n5690), .Z(n5692) );
  AND U6596 ( .A(n5693), .B(n5692), .Z(n6145) );
  NAND U6597 ( .A(a[47]), .B(b[49]), .Z(n6153) );
  OR U6598 ( .A(n5695), .B(n5694), .Z(n5699) );
  OR U6599 ( .A(n5697), .B(n5696), .Z(n5698) );
  AND U6600 ( .A(n5699), .B(n5698), .Z(n6150) );
  ANDN U6601 ( .B(b[50]), .A(n194), .Z(n6228) );
  OR U6602 ( .A(n5701), .B(n5700), .Z(n5705) );
  NANDN U6603 ( .A(n5703), .B(n5702), .Z(n5704) );
  AND U6604 ( .A(n5705), .B(n5704), .Z(n6229) );
  XNOR U6605 ( .A(n6228), .B(n6229), .Z(n6231) );
  NAND U6606 ( .A(a[43]), .B(b[53]), .Z(n6165) );
  OR U6607 ( .A(n5707), .B(n5706), .Z(n5711) );
  OR U6608 ( .A(n5709), .B(n5708), .Z(n5710) );
  AND U6609 ( .A(n5711), .B(n5710), .Z(n6162) );
  ANDN U6610 ( .B(b[54]), .A(n190), .Z(n6216) );
  OR U6611 ( .A(n5713), .B(n5712), .Z(n5717) );
  NANDN U6612 ( .A(n5715), .B(n5714), .Z(n5716) );
  AND U6613 ( .A(n5717), .B(n5716), .Z(n6217) );
  XNOR U6614 ( .A(n6216), .B(n6217), .Z(n6219) );
  NAND U6615 ( .A(a[40]), .B(b[56]), .Z(n6211) );
  OR U6616 ( .A(n5719), .B(n5718), .Z(n5723) );
  NANDN U6617 ( .A(n5721), .B(n5720), .Z(n5722) );
  NAND U6618 ( .A(n5723), .B(n5722), .Z(n6210) );
  XNOR U6619 ( .A(n6211), .B(n6210), .Z(n6213) );
  NAND U6620 ( .A(a[39]), .B(b[57]), .Z(n6177) );
  OR U6621 ( .A(n5725), .B(n5724), .Z(n5729) );
  OR U6622 ( .A(n5727), .B(n5726), .Z(n5728) );
  AND U6623 ( .A(n5729), .B(n5728), .Z(n6174) );
  ANDN U6624 ( .B(b[58]), .A(n186), .Z(n6204) );
  OR U6625 ( .A(n5731), .B(n5730), .Z(n5735) );
  NANDN U6626 ( .A(n5733), .B(n5732), .Z(n5734) );
  AND U6627 ( .A(n5735), .B(n5734), .Z(n6205) );
  XNOR U6628 ( .A(n6204), .B(n6205), .Z(n6207) );
  NAND U6629 ( .A(b[61]), .B(a[35]), .Z(n6188) );
  OR U6630 ( .A(n5737), .B(n5736), .Z(n5741) );
  OR U6631 ( .A(n5739), .B(n5738), .Z(n5740) );
  AND U6632 ( .A(n5741), .B(n5740), .Z(n6186) );
  ANDN U6633 ( .B(b[63]), .A(n21751), .Z(n6194) );
  ANDN U6634 ( .B(a[34]), .A(n159), .Z(n6192) );
  OR U6635 ( .A(n5743), .B(n5742), .Z(n5747) );
  OR U6636 ( .A(n5745), .B(n5744), .Z(n5746) );
  AND U6637 ( .A(n5747), .B(n5746), .Z(n6193) );
  XNOR U6638 ( .A(n6192), .B(n6193), .Z(n6195) );
  XNOR U6639 ( .A(n6194), .B(n6195), .Z(n6187) );
  XNOR U6640 ( .A(n6186), .B(n6187), .Z(n6189) );
  XOR U6641 ( .A(n6188), .B(n6189), .Z(n6200) );
  NAND U6642 ( .A(a[36]), .B(b[60]), .Z(n6199) );
  OR U6643 ( .A(n5749), .B(n5748), .Z(n5753) );
  OR U6644 ( .A(n5751), .B(n5750), .Z(n5752) );
  NAND U6645 ( .A(n5753), .B(n5752), .Z(n6198) );
  XNOR U6646 ( .A(n6199), .B(n6198), .Z(n6201) );
  XNOR U6647 ( .A(n6200), .B(n6201), .Z(n6180) );
  OR U6648 ( .A(n5755), .B(n5754), .Z(n5759) );
  NANDN U6649 ( .A(n5757), .B(n5756), .Z(n5758) );
  NAND U6650 ( .A(n5759), .B(n5758), .Z(n6181) );
  XNOR U6651 ( .A(n6180), .B(n6181), .Z(n6183) );
  ANDN U6652 ( .B(b[59]), .A(n21772), .Z(n6182) );
  XNOR U6653 ( .A(n6183), .B(n6182), .Z(n6206) );
  XOR U6654 ( .A(n6207), .B(n6206), .Z(n6175) );
  XNOR U6655 ( .A(n6174), .B(n6175), .Z(n6176) );
  XOR U6656 ( .A(n6177), .B(n6176), .Z(n6212) );
  OR U6657 ( .A(n5761), .B(n5760), .Z(n5765) );
  OR U6658 ( .A(n5763), .B(n5762), .Z(n5764) );
  NAND U6659 ( .A(n5765), .B(n5764), .Z(n6169) );
  XOR U6660 ( .A(n6168), .B(n6169), .Z(n6170) );
  ANDN U6661 ( .B(b[55]), .A(n189), .Z(n6171) );
  XOR U6662 ( .A(n6170), .B(n6171), .Z(n6218) );
  XOR U6663 ( .A(n6219), .B(n6218), .Z(n6163) );
  XNOR U6664 ( .A(n6162), .B(n6163), .Z(n6164) );
  XOR U6665 ( .A(n6165), .B(n6164), .Z(n6224) );
  OR U6666 ( .A(n5767), .B(n5766), .Z(n5771) );
  NANDN U6667 ( .A(n5769), .B(n5768), .Z(n5770) );
  AND U6668 ( .A(n5771), .B(n5770), .Z(n6222) );
  ANDN U6669 ( .B(b[52]), .A(n192), .Z(n6223) );
  XNOR U6670 ( .A(n6222), .B(n6223), .Z(n6225) );
  XOR U6671 ( .A(n6224), .B(n6225), .Z(n6156) );
  OR U6672 ( .A(n5773), .B(n5772), .Z(n5777) );
  OR U6673 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U6674 ( .A(n5777), .B(n5776), .Z(n6157) );
  XOR U6675 ( .A(n6156), .B(n6157), .Z(n6159) );
  ANDN U6676 ( .B(b[51]), .A(n193), .Z(n6158) );
  XNOR U6677 ( .A(n6159), .B(n6158), .Z(n6230) );
  XOR U6678 ( .A(n6231), .B(n6230), .Z(n6151) );
  XNOR U6679 ( .A(n6150), .B(n6151), .Z(n6152) );
  XOR U6680 ( .A(n6153), .B(n6152), .Z(n6236) );
  ANDN U6681 ( .B(b[48]), .A(n196), .Z(n6234) );
  OR U6682 ( .A(n5779), .B(n5778), .Z(n5783) );
  OR U6683 ( .A(n5781), .B(n5780), .Z(n5782) );
  AND U6684 ( .A(n5783), .B(n5782), .Z(n6235) );
  XNOR U6685 ( .A(n6234), .B(n6235), .Z(n6237) );
  XOR U6686 ( .A(n6236), .B(n6237), .Z(n6144) );
  XOR U6687 ( .A(n6145), .B(n6144), .Z(n6147) );
  XNOR U6688 ( .A(n6146), .B(n6147), .Z(n6243) );
  ANDN U6689 ( .B(b[46]), .A(n198), .Z(n6240) );
  OR U6690 ( .A(n5785), .B(n5784), .Z(n5789) );
  OR U6691 ( .A(n5787), .B(n5786), .Z(n5788) );
  AND U6692 ( .A(n5789), .B(n5788), .Z(n6241) );
  XOR U6693 ( .A(n6240), .B(n6241), .Z(n6242) );
  OR U6694 ( .A(n5791), .B(n5790), .Z(n5795) );
  NANDN U6695 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U6696 ( .A(n5795), .B(n5794), .Z(n6139) );
  XOR U6697 ( .A(n6138), .B(n6139), .Z(n6141) );
  ANDN U6698 ( .B(b[45]), .A(n199), .Z(n6140) );
  XNOR U6699 ( .A(n6141), .B(n6140), .Z(n6248) );
  XOR U6700 ( .A(n6249), .B(n6248), .Z(n6133) );
  XNOR U6701 ( .A(n6132), .B(n6133), .Z(n6135) );
  NAND U6702 ( .A(a[53]), .B(b[43]), .Z(n6134) );
  XOR U6703 ( .A(n6135), .B(n6134), .Z(n6253) );
  XNOR U6704 ( .A(n6252), .B(n6253), .Z(n6255) );
  ANDN U6705 ( .B(b[42]), .A(n202), .Z(n6254) );
  XOR U6706 ( .A(n6255), .B(n6254), .Z(n6126) );
  NAND U6707 ( .A(a[55]), .B(b[41]), .Z(n6127) );
  XOR U6708 ( .A(n6126), .B(n6127), .Z(n6129) );
  OR U6709 ( .A(n5796), .B(n5797), .Z(n6125) );
  XNOR U6710 ( .A(n5797), .B(n5796), .Z(n6595) );
  NAND U6711 ( .A(a[55]), .B(b[40]), .Z(n6121) );
  XOR U6712 ( .A(n5799), .B(n5798), .Z(n6120) );
  NANDN U6713 ( .A(n6121), .B(n6120), .Z(n6123) );
  ANDN U6714 ( .B(b[40]), .A(n201), .Z(n6108) );
  XNOR U6715 ( .A(n5801), .B(n5800), .Z(n5802) );
  ANDN U6716 ( .B(b[40]), .A(n200), .Z(n5803) );
  OR U6717 ( .A(n5802), .B(n5803), .Z(n6107) );
  XNOR U6718 ( .A(n5803), .B(n5802), .Z(n6263) );
  XNOR U6719 ( .A(n5805), .B(n5804), .Z(n6103) );
  XOR U6720 ( .A(n5807), .B(n5806), .Z(n6099) );
  XOR U6721 ( .A(n5809), .B(n5808), .Z(n6089) );
  NAND U6722 ( .A(a[47]), .B(b[40]), .Z(n6085) );
  XNOR U6723 ( .A(n5811), .B(n5810), .Z(n6084) );
  NANDN U6724 ( .A(n6085), .B(n6084), .Z(n6087) );
  ANDN U6725 ( .B(b[40]), .A(n194), .Z(n5814) );
  XOR U6726 ( .A(n5813), .B(n5812), .Z(n5815) );
  NANDN U6727 ( .A(n5814), .B(n5815), .Z(n6083) );
  XOR U6728 ( .A(n5815), .B(n5814), .Z(n6545) );
  XOR U6729 ( .A(n5817), .B(n5816), .Z(n6079) );
  XOR U6730 ( .A(n5819), .B(n5818), .Z(n6075) );
  XOR U6731 ( .A(n5821), .B(n5820), .Z(n6065) );
  NAND U6732 ( .A(b[40]), .B(a[42]), .Z(n6064) );
  OR U6733 ( .A(n6065), .B(n6064), .Z(n6067) );
  XNOR U6734 ( .A(n5823), .B(n5822), .Z(n6061) );
  ANDN U6735 ( .B(b[40]), .A(n187), .Z(n6051) );
  XOR U6736 ( .A(n5825), .B(n5824), .Z(n6050) );
  OR U6737 ( .A(n6051), .B(n6050), .Z(n6053) );
  ANDN U6738 ( .B(b[40]), .A(n21772), .Z(n5828) );
  XOR U6739 ( .A(n5827), .B(n5826), .Z(n5829) );
  NANDN U6740 ( .A(n5828), .B(n5829), .Z(n6043) );
  XOR U6741 ( .A(n5829), .B(n5828), .Z(n6279) );
  NAND U6742 ( .A(a[36]), .B(b[40]), .Z(n6037) );
  XNOR U6743 ( .A(n5831), .B(n5830), .Z(n6033) );
  NAND U6744 ( .A(a[34]), .B(b[40]), .Z(n5835) );
  NANDN U6745 ( .A(n5835), .B(n5834), .Z(n6031) );
  XOR U6746 ( .A(n5835), .B(n5834), .Z(n6288) );
  NAND U6747 ( .A(a[32]), .B(b[40]), .Z(n5838) );
  NANDN U6748 ( .A(n5838), .B(n5839), .Z(n6023) );
  XOR U6749 ( .A(n5839), .B(n5838), .Z(n6483) );
  NAND U6750 ( .A(a[31]), .B(b[40]), .Z(n6018) );
  NANDN U6751 ( .A(n6018), .B(n6019), .Z(n6021) );
  XOR U6752 ( .A(n5843), .B(n5842), .Z(n6015) );
  XNOR U6753 ( .A(n5845), .B(n5844), .Z(n6011) );
  XOR U6754 ( .A(n5847), .B(n5846), .Z(n6007) );
  XNOR U6755 ( .A(n5849), .B(n5848), .Z(n6003) );
  ANDN U6756 ( .B(b[40]), .A(n179), .Z(n5852) );
  OR U6757 ( .A(n5853), .B(n5852), .Z(n6001) );
  XNOR U6758 ( .A(n5853), .B(n5852), .Z(n6297) );
  XNOR U6759 ( .A(n5855), .B(n5854), .Z(n5997) );
  XNOR U6760 ( .A(n5857), .B(n5856), .Z(n5992) );
  NAND U6761 ( .A(a[23]), .B(b[40]), .Z(n5989) );
  XOR U6762 ( .A(n5859), .B(n5858), .Z(n5988) );
  NANDN U6763 ( .A(n5989), .B(n5988), .Z(n5991) );
  XOR U6764 ( .A(n5861), .B(n5860), .Z(n5984) );
  XOR U6765 ( .A(n5863), .B(n5862), .Z(n5975) );
  XNOR U6766 ( .A(n5865), .B(n5864), .Z(n5965) );
  XNOR U6767 ( .A(n5867), .B(n5866), .Z(n5869) );
  AND U6768 ( .A(a[17]), .B(b[40]), .Z(n5868) );
  NANDN U6769 ( .A(n5869), .B(n5868), .Z(n5963) );
  XOR U6770 ( .A(n5869), .B(n5868), .Z(n6308) );
  NAND U6771 ( .A(a[16]), .B(b[40]), .Z(n5956) );
  NAND U6772 ( .A(a[13]), .B(b[40]), .Z(n5940) );
  XOR U6773 ( .A(n5871), .B(n5870), .Z(n5941) );
  OR U6774 ( .A(n5940), .B(n5941), .Z(n5943) );
  XNOR U6775 ( .A(n5873), .B(n5872), .Z(n5874) );
  ANDN U6776 ( .B(b[40]), .A(n169), .Z(n5875) );
  OR U6777 ( .A(n5874), .B(n5875), .Z(n5939) );
  XOR U6778 ( .A(n5875), .B(n5874), .Z(n6314) );
  XNOR U6779 ( .A(n5877), .B(n5876), .Z(n5934) );
  XOR U6780 ( .A(n5879), .B(n5878), .Z(n5930) );
  XNOR U6781 ( .A(n5881), .B(n5880), .Z(n5921) );
  XOR U6782 ( .A(n5883), .B(n5882), .Z(n5885) );
  AND U6783 ( .A(a[7]), .B(b[40]), .Z(n5884) );
  NANDN U6784 ( .A(n5885), .B(n5884), .Z(n5919) );
  XOR U6785 ( .A(n5885), .B(n5884), .Z(n6324) );
  XNOR U6786 ( .A(n5887), .B(n5886), .Z(n5909) );
  XNOR U6787 ( .A(n5889), .B(n5888), .Z(n5904) );
  XNOR U6788 ( .A(n5891), .B(n5890), .Z(n5900) );
  NAND U6789 ( .A(b[41]), .B(a[1]), .Z(n5893) );
  NAND U6790 ( .A(n5893), .B(n5892), .Z(n5896) );
  NANDN U6791 ( .A(n154), .B(a[0]), .Z(n7140) );
  OR U6792 ( .A(n5893), .B(n7140), .Z(n6339) );
  NANDN U6793 ( .A(n5895), .B(n6339), .Z(n5894) );
  AND U6794 ( .A(n5896), .B(n5894), .Z(n5899) );
  XNOR U6795 ( .A(n6339), .B(n5895), .Z(n5897) );
  NAND U6796 ( .A(n5897), .B(n5896), .Z(n6335) );
  ANDN U6797 ( .B(b[40]), .A(n162), .Z(n6334) );
  OR U6798 ( .A(n6335), .B(n6334), .Z(n5898) );
  AND U6799 ( .A(n5899), .B(n5898), .Z(n5901) );
  OR U6800 ( .A(n5900), .B(n5901), .Z(n5903) );
  XNOR U6801 ( .A(n5901), .B(n5900), .Z(n6332) );
  ANDN U6802 ( .B(b[40]), .A(n21580), .Z(n6333) );
  OR U6803 ( .A(n6332), .B(n6333), .Z(n5902) );
  AND U6804 ( .A(n5903), .B(n5902), .Z(n5905) );
  OR U6805 ( .A(n5904), .B(n5905), .Z(n5907) );
  XNOR U6806 ( .A(n5905), .B(n5904), .Z(n6330) );
  ANDN U6807 ( .B(b[40]), .A(n163), .Z(n6331) );
  OR U6808 ( .A(n6330), .B(n6331), .Z(n5906) );
  AND U6809 ( .A(n5907), .B(n5906), .Z(n5908) );
  OR U6810 ( .A(n5909), .B(n5908), .Z(n5911) );
  XNOR U6811 ( .A(n5909), .B(n5908), .Z(n6358) );
  NAND U6812 ( .A(b[40]), .B(a[5]), .Z(n6359) );
  NANDN U6813 ( .A(n6358), .B(n6359), .Z(n5910) );
  NAND U6814 ( .A(n5911), .B(n5910), .Z(n5913) );
  AND U6815 ( .A(a[6]), .B(b[40]), .Z(n5912) );
  NANDN U6816 ( .A(n5913), .B(n5912), .Z(n5917) );
  XOR U6817 ( .A(n5913), .B(n5912), .Z(n6326) );
  XOR U6818 ( .A(n5915), .B(n5914), .Z(n6327) );
  NANDN U6819 ( .A(n6326), .B(n6327), .Z(n5916) );
  AND U6820 ( .A(n5917), .B(n5916), .Z(n6325) );
  OR U6821 ( .A(n6324), .B(n6325), .Z(n5918) );
  AND U6822 ( .A(n5919), .B(n5918), .Z(n5920) );
  OR U6823 ( .A(n5921), .B(n5920), .Z(n5923) );
  XNOR U6824 ( .A(n5921), .B(n5920), .Z(n6369) );
  NAND U6825 ( .A(a[8]), .B(b[40]), .Z(n6368) );
  OR U6826 ( .A(n6369), .B(n6368), .Z(n5922) );
  NAND U6827 ( .A(n5923), .B(n5922), .Z(n5926) );
  XOR U6828 ( .A(n5925), .B(n5924), .Z(n5927) );
  OR U6829 ( .A(n5926), .B(n5927), .Z(n5929) );
  ANDN U6830 ( .B(b[40]), .A(n21615), .Z(n6323) );
  XOR U6831 ( .A(n5927), .B(n5926), .Z(n6322) );
  NANDN U6832 ( .A(n6323), .B(n6322), .Z(n5928) );
  AND U6833 ( .A(n5929), .B(n5928), .Z(n5931) );
  OR U6834 ( .A(n5930), .B(n5931), .Z(n5933) );
  XNOR U6835 ( .A(n5931), .B(n5930), .Z(n6320) );
  ANDN U6836 ( .B(b[40]), .A(n168), .Z(n6321) );
  OR U6837 ( .A(n6320), .B(n6321), .Z(n5932) );
  AND U6838 ( .A(n5933), .B(n5932), .Z(n5935) );
  OR U6839 ( .A(n5934), .B(n5935), .Z(n5937) );
  XNOR U6840 ( .A(n5935), .B(n5934), .Z(n6316) );
  ANDN U6841 ( .B(b[40]), .A(n21164), .Z(n6317) );
  OR U6842 ( .A(n6316), .B(n6317), .Z(n5936) );
  NAND U6843 ( .A(n5937), .B(n5936), .Z(n6315) );
  NAND U6844 ( .A(n6314), .B(n6315), .Z(n5938) );
  NAND U6845 ( .A(n5939), .B(n5938), .Z(n6389) );
  XOR U6846 ( .A(n5941), .B(n5940), .Z(n6388) );
  NANDN U6847 ( .A(n6389), .B(n6388), .Z(n5942) );
  AND U6848 ( .A(n5943), .B(n5942), .Z(n5946) );
  NANDN U6849 ( .A(n5946), .B(n5947), .Z(n5949) );
  XOR U6850 ( .A(n5947), .B(n5946), .Z(n6395) );
  AND U6851 ( .A(a[14]), .B(b[40]), .Z(n6394) );
  NANDN U6852 ( .A(n6395), .B(n6394), .Z(n5948) );
  AND U6853 ( .A(n5949), .B(n5948), .Z(n5953) );
  XNOR U6854 ( .A(n5951), .B(n5950), .Z(n5952) );
  NANDN U6855 ( .A(n5953), .B(n5952), .Z(n5955) );
  NAND U6856 ( .A(a[15]), .B(b[40]), .Z(n6403) );
  NANDN U6857 ( .A(n6403), .B(n6402), .Z(n5954) );
  AND U6858 ( .A(n5955), .B(n5954), .Z(n5957) );
  OR U6859 ( .A(n5956), .B(n5957), .Z(n5961) );
  XNOR U6860 ( .A(n5957), .B(n5956), .Z(n6311) );
  NANDN U6861 ( .A(n6311), .B(n6310), .Z(n5960) );
  AND U6862 ( .A(n5961), .B(n5960), .Z(n6309) );
  OR U6863 ( .A(n6308), .B(n6309), .Z(n5962) );
  AND U6864 ( .A(n5963), .B(n5962), .Z(n5964) );
  OR U6865 ( .A(n5965), .B(n5964), .Z(n5967) );
  XNOR U6866 ( .A(n5965), .B(n5964), .Z(n6307) );
  AND U6867 ( .A(a[18]), .B(b[40]), .Z(n6306) );
  NANDN U6868 ( .A(n6307), .B(n6306), .Z(n5966) );
  AND U6869 ( .A(n5967), .B(n5966), .Z(n5970) );
  XNOR U6870 ( .A(n5969), .B(n5968), .Z(n5971) );
  NANDN U6871 ( .A(n5970), .B(n5971), .Z(n5973) );
  NAND U6872 ( .A(a[19]), .B(b[40]), .Z(n6417) );
  XOR U6873 ( .A(n5971), .B(n5970), .Z(n6416) );
  OR U6874 ( .A(n6417), .B(n6416), .Z(n5972) );
  AND U6875 ( .A(n5973), .B(n5972), .Z(n5974) );
  OR U6876 ( .A(n5975), .B(n5974), .Z(n5977) );
  NAND U6877 ( .A(a[20]), .B(b[40]), .Z(n6305) );
  XNOR U6878 ( .A(n5975), .B(n5974), .Z(n6304) );
  OR U6879 ( .A(n6305), .B(n6304), .Z(n5976) );
  NAND U6880 ( .A(n5977), .B(n5976), .Z(n5980) );
  XOR U6881 ( .A(n5979), .B(n5978), .Z(n5981) );
  OR U6882 ( .A(n5980), .B(n5981), .Z(n5983) );
  ANDN U6883 ( .B(b[40]), .A(n21681), .Z(n6303) );
  XOR U6884 ( .A(n5981), .B(n5980), .Z(n6302) );
  NANDN U6885 ( .A(n6303), .B(n6302), .Z(n5982) );
  AND U6886 ( .A(n5983), .B(n5982), .Z(n5985) );
  OR U6887 ( .A(n5984), .B(n5985), .Z(n5987) );
  XNOR U6888 ( .A(n5985), .B(n5984), .Z(n6300) );
  NAND U6889 ( .A(b[40]), .B(a[22]), .Z(n6301) );
  NANDN U6890 ( .A(n6300), .B(n6301), .Z(n5986) );
  NAND U6891 ( .A(n5987), .B(n5986), .Z(n6435) );
  NANDN U6892 ( .A(n6435), .B(n6434), .Z(n5990) );
  AND U6893 ( .A(n5991), .B(n5990), .Z(n5993) );
  OR U6894 ( .A(n5992), .B(n5993), .Z(n5995) );
  NAND U6895 ( .A(a[24]), .B(b[40]), .Z(n6441) );
  XNOR U6896 ( .A(n5993), .B(n5992), .Z(n6440) );
  OR U6897 ( .A(n6441), .B(n6440), .Z(n5994) );
  NAND U6898 ( .A(n5995), .B(n5994), .Z(n5996) );
  OR U6899 ( .A(n5997), .B(n5996), .Z(n5999) );
  ANDN U6900 ( .B(b[40]), .A(n21703), .Z(n6299) );
  XOR U6901 ( .A(n5997), .B(n5996), .Z(n6298) );
  NANDN U6902 ( .A(n6299), .B(n6298), .Z(n5998) );
  AND U6903 ( .A(n5999), .B(n5998), .Z(n6296) );
  OR U6904 ( .A(n6297), .B(n6296), .Z(n6000) );
  NAND U6905 ( .A(n6001), .B(n6000), .Z(n6002) );
  NANDN U6906 ( .A(n6003), .B(n6002), .Z(n6005) );
  ANDN U6907 ( .B(b[40]), .A(n21716), .Z(n6455) );
  OR U6908 ( .A(n6455), .B(n6454), .Z(n6004) );
  NAND U6909 ( .A(n6005), .B(n6004), .Z(n6006) );
  NANDN U6910 ( .A(n6007), .B(n6006), .Z(n6009) );
  ANDN U6911 ( .B(b[40]), .A(n180), .Z(n6461) );
  NANDN U6912 ( .A(n6461), .B(n6460), .Z(n6008) );
  NAND U6913 ( .A(n6009), .B(n6008), .Z(n6010) );
  NANDN U6914 ( .A(n6011), .B(n6010), .Z(n6013) );
  ANDN U6915 ( .B(b[40]), .A(n21727), .Z(n6467) );
  OR U6916 ( .A(n6467), .B(n6466), .Z(n6012) );
  NAND U6917 ( .A(n6013), .B(n6012), .Z(n6014) );
  NANDN U6918 ( .A(n6015), .B(n6014), .Z(n6017) );
  ANDN U6919 ( .B(b[40]), .A(n181), .Z(n6473) );
  NANDN U6920 ( .A(n6473), .B(n6472), .Z(n6016) );
  NAND U6921 ( .A(n6017), .B(n6016), .Z(n6295) );
  XNOR U6922 ( .A(n6019), .B(n6018), .Z(n6294) );
  NANDN U6923 ( .A(n6295), .B(n6294), .Z(n6020) );
  NAND U6924 ( .A(n6021), .B(n6020), .Z(n6482) );
  NANDN U6925 ( .A(n6483), .B(n6482), .Z(n6022) );
  AND U6926 ( .A(n6023), .B(n6022), .Z(n6026) );
  NANDN U6927 ( .A(n6026), .B(n6027), .Z(n6029) );
  XOR U6928 ( .A(n6027), .B(n6026), .Z(n6293) );
  NAND U6929 ( .A(a[33]), .B(b[40]), .Z(n6292) );
  OR U6930 ( .A(n6293), .B(n6292), .Z(n6028) );
  AND U6931 ( .A(n6029), .B(n6028), .Z(n6289) );
  OR U6932 ( .A(n6288), .B(n6289), .Z(n6030) );
  NAND U6933 ( .A(n6031), .B(n6030), .Z(n6032) );
  NANDN U6934 ( .A(n6033), .B(n6032), .Z(n6035) );
  NAND U6935 ( .A(b[40]), .B(a[35]), .Z(n6284) );
  NANDN U6936 ( .A(n6284), .B(n6285), .Z(n6034) );
  NAND U6937 ( .A(n6035), .B(n6034), .Z(n6036) );
  NANDN U6938 ( .A(n6037), .B(n6036), .Z(n6041) );
  XNOR U6939 ( .A(n6039), .B(n6038), .Z(n6281) );
  NAND U6940 ( .A(n6280), .B(n6281), .Z(n6040) );
  NAND U6941 ( .A(n6041), .B(n6040), .Z(n6278) );
  OR U6942 ( .A(n6279), .B(n6278), .Z(n6042) );
  AND U6943 ( .A(n6043), .B(n6042), .Z(n6047) );
  XOR U6944 ( .A(n6045), .B(n6044), .Z(n6046) );
  NANDN U6945 ( .A(n6047), .B(n6046), .Z(n6049) );
  ANDN U6946 ( .B(b[40]), .A(n186), .Z(n6277) );
  NANDN U6947 ( .A(n6277), .B(n6276), .Z(n6048) );
  NAND U6948 ( .A(n6049), .B(n6048), .Z(n6507) );
  XOR U6949 ( .A(n6051), .B(n6050), .Z(n6506) );
  NAND U6950 ( .A(n6507), .B(n6506), .Z(n6052) );
  AND U6951 ( .A(n6053), .B(n6052), .Z(n6057) );
  XOR U6952 ( .A(n6055), .B(n6054), .Z(n6056) );
  NANDN U6953 ( .A(n6057), .B(n6056), .Z(n6059) );
  ANDN U6954 ( .B(b[40]), .A(n188), .Z(n6513) );
  OR U6955 ( .A(n6513), .B(n6512), .Z(n6058) );
  NAND U6956 ( .A(n6059), .B(n6058), .Z(n6060) );
  NANDN U6957 ( .A(n6061), .B(n6060), .Z(n6063) );
  NANDN U6958 ( .A(n154), .B(a[41]), .Z(n6275) );
  NAND U6959 ( .A(n6274), .B(n6275), .Z(n6062) );
  NAND U6960 ( .A(n6063), .B(n6062), .Z(n6523) );
  XOR U6961 ( .A(n6065), .B(n6064), .Z(n6522) );
  NANDN U6962 ( .A(n6523), .B(n6522), .Z(n6066) );
  NAND U6963 ( .A(n6067), .B(n6066), .Z(n6071) );
  XOR U6964 ( .A(n6069), .B(n6068), .Z(n6070) );
  NANDN U6965 ( .A(n6071), .B(n6070), .Z(n6073) );
  ANDN U6966 ( .B(b[40]), .A(n191), .Z(n6529) );
  XOR U6967 ( .A(n6071), .B(n6070), .Z(n6528) );
  OR U6968 ( .A(n6529), .B(n6528), .Z(n6072) );
  NAND U6969 ( .A(n6073), .B(n6072), .Z(n6074) );
  NANDN U6970 ( .A(n6075), .B(n6074), .Z(n6077) );
  ANDN U6971 ( .B(b[40]), .A(n192), .Z(n6535) );
  NANDN U6972 ( .A(n6535), .B(n6534), .Z(n6076) );
  NAND U6973 ( .A(n6077), .B(n6076), .Z(n6078) );
  NANDN U6974 ( .A(n6079), .B(n6078), .Z(n6081) );
  ANDN U6975 ( .B(b[40]), .A(n193), .Z(n6273) );
  NANDN U6976 ( .A(n6273), .B(n6272), .Z(n6080) );
  NAND U6977 ( .A(n6081), .B(n6080), .Z(n6544) );
  NANDN U6978 ( .A(n6545), .B(n6544), .Z(n6082) );
  NAND U6979 ( .A(n6083), .B(n6082), .Z(n6551) );
  XNOR U6980 ( .A(n6085), .B(n6084), .Z(n6550) );
  NANDN U6981 ( .A(n6551), .B(n6550), .Z(n6086) );
  NAND U6982 ( .A(n6087), .B(n6086), .Z(n6088) );
  NANDN U6983 ( .A(n6089), .B(n6088), .Z(n6091) );
  XOR U6984 ( .A(n6089), .B(n6088), .Z(n6557) );
  NAND U6985 ( .A(b[40]), .B(a[48]), .Z(n6556) );
  OR U6986 ( .A(n6557), .B(n6556), .Z(n6090) );
  NAND U6987 ( .A(n6091), .B(n6090), .Z(n6095) );
  XOR U6988 ( .A(n6093), .B(n6092), .Z(n6094) );
  NANDN U6989 ( .A(n6095), .B(n6094), .Z(n6097) );
  ANDN U6990 ( .B(b[40]), .A(n197), .Z(n6269) );
  NANDN U6991 ( .A(n6269), .B(n6268), .Z(n6096) );
  NAND U6992 ( .A(n6097), .B(n6096), .Z(n6098) );
  NANDN U6993 ( .A(n6099), .B(n6098), .Z(n6101) );
  ANDN U6994 ( .B(b[40]), .A(n198), .Z(n6267) );
  NANDN U6995 ( .A(n6267), .B(n6266), .Z(n6100) );
  NAND U6996 ( .A(n6101), .B(n6100), .Z(n6102) );
  NANDN U6997 ( .A(n6103), .B(n6102), .Z(n6105) );
  ANDN U6998 ( .B(b[40]), .A(n199), .Z(n6569) );
  OR U6999 ( .A(n6569), .B(n6568), .Z(n6104) );
  AND U7000 ( .A(n6105), .B(n6104), .Z(n6262) );
  OR U7001 ( .A(n6263), .B(n6262), .Z(n6106) );
  AND U7002 ( .A(n6107), .B(n6106), .Z(n6109) );
  OR U7003 ( .A(n6108), .B(n6109), .Z(n6113) );
  XNOR U7004 ( .A(n6109), .B(n6108), .Z(n6577) );
  OR U7005 ( .A(n6577), .B(n6576), .Z(n6112) );
  NAND U7006 ( .A(n6113), .B(n6112), .Z(n6117) );
  AND U7007 ( .A(a[54]), .B(b[40]), .Z(n6116) );
  NANDN U7008 ( .A(n6117), .B(n6116), .Z(n6119) );
  XOR U7009 ( .A(n6115), .B(n6114), .Z(n6583) );
  XNOR U7010 ( .A(n6117), .B(n6116), .Z(n6582) );
  NANDN U7011 ( .A(n6583), .B(n6582), .Z(n6118) );
  AND U7012 ( .A(n6119), .B(n6118), .Z(n6260) );
  NANDN U7013 ( .A(n6260), .B(n6261), .Z(n6122) );
  NAND U7014 ( .A(n6123), .B(n6122), .Z(n6594) );
  OR U7015 ( .A(n6595), .B(n6594), .Z(n6124) );
  NAND U7016 ( .A(n6125), .B(n6124), .Z(n6733) );
  OR U7017 ( .A(n6127), .B(n6126), .Z(n6131) );
  NAND U7018 ( .A(n6129), .B(n6128), .Z(n6130) );
  NAND U7019 ( .A(n6131), .B(n6130), .Z(n6601) );
  ANDN U7020 ( .B(b[43]), .A(n202), .Z(n6609) );
  OR U7021 ( .A(n6133), .B(n6132), .Z(n6137) );
  OR U7022 ( .A(n6135), .B(n6134), .Z(n6136) );
  NAND U7023 ( .A(n6137), .B(n6136), .Z(n6607) );
  NAND U7024 ( .A(a[52]), .B(b[45]), .Z(n6615) );
  NANDN U7025 ( .A(n6139), .B(n6138), .Z(n6143) );
  OR U7026 ( .A(n6141), .B(n6140), .Z(n6142) );
  NAND U7027 ( .A(n6143), .B(n6142), .Z(n6613) );
  ANDN U7028 ( .B(b[47]), .A(n198), .Z(n6620) );
  NANDN U7029 ( .A(n6145), .B(n6144), .Z(n6149) );
  OR U7030 ( .A(n6147), .B(n6146), .Z(n6148) );
  AND U7031 ( .A(n6149), .B(n6148), .Z(n6619) );
  ANDN U7032 ( .B(b[49]), .A(n196), .Z(n6627) );
  OR U7033 ( .A(n6151), .B(n6150), .Z(n6155) );
  OR U7034 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U7035 ( .A(n6155), .B(n6154), .Z(n6625) );
  NAND U7036 ( .A(a[46]), .B(b[51]), .Z(n6633) );
  NANDN U7037 ( .A(n6157), .B(n6156), .Z(n6161) );
  OR U7038 ( .A(n6159), .B(n6158), .Z(n6160) );
  NAND U7039 ( .A(n6161), .B(n6160), .Z(n6631) );
  ANDN U7040 ( .B(b[53]), .A(n192), .Z(n6639) );
  OR U7041 ( .A(n6163), .B(n6162), .Z(n6167) );
  OR U7042 ( .A(n6165), .B(n6164), .Z(n6166) );
  NAND U7043 ( .A(n6167), .B(n6166), .Z(n6637) );
  NAND U7044 ( .A(a[42]), .B(b[55]), .Z(n6645) );
  OR U7045 ( .A(n6169), .B(n6168), .Z(n6173) );
  NANDN U7046 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U7047 ( .A(n6173), .B(n6172), .Z(n6643) );
  NAND U7048 ( .A(a[40]), .B(b[57]), .Z(n6651) );
  OR U7049 ( .A(n6175), .B(n6174), .Z(n6179) );
  OR U7050 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U7051 ( .A(n6179), .B(n6178), .Z(n6648) );
  NAND U7052 ( .A(a[38]), .B(b[59]), .Z(n6657) );
  OR U7053 ( .A(n6181), .B(n6180), .Z(n6185) );
  OR U7054 ( .A(n6183), .B(n6182), .Z(n6184) );
  NAND U7055 ( .A(n6185), .B(n6184), .Z(n6655) );
  ANDN U7056 ( .B(b[61]), .A(n185), .Z(n6662) );
  OR U7057 ( .A(n6187), .B(n6186), .Z(n6191) );
  NANDN U7058 ( .A(n6189), .B(n6188), .Z(n6190) );
  AND U7059 ( .A(n6191), .B(n6190), .Z(n6660) );
  ANDN U7060 ( .B(b[63]), .A(n183), .Z(n6668) );
  ANDN U7061 ( .B(a[35]), .A(n159), .Z(n6666) );
  OR U7062 ( .A(n6193), .B(n6192), .Z(n6197) );
  OR U7063 ( .A(n6195), .B(n6194), .Z(n6196) );
  AND U7064 ( .A(n6197), .B(n6196), .Z(n6667) );
  XNOR U7065 ( .A(n6666), .B(n6667), .Z(n6669) );
  XNOR U7066 ( .A(n6668), .B(n6669), .Z(n6661) );
  XNOR U7067 ( .A(n6660), .B(n6661), .Z(n6663) );
  XNOR U7068 ( .A(n6662), .B(n6663), .Z(n6675) );
  ANDN U7069 ( .B(b[60]), .A(n21772), .Z(n6672) );
  OR U7070 ( .A(n6199), .B(n6198), .Z(n6203) );
  NANDN U7071 ( .A(n6201), .B(n6200), .Z(n6202) );
  NAND U7072 ( .A(n6203), .B(n6202), .Z(n6673) );
  XNOR U7073 ( .A(n6672), .B(n6673), .Z(n6674) );
  XOR U7074 ( .A(n6675), .B(n6674), .Z(n6654) );
  XOR U7075 ( .A(n6655), .B(n6654), .Z(n6656) );
  ANDN U7076 ( .B(b[58]), .A(n187), .Z(n6678) );
  OR U7077 ( .A(n6205), .B(n6204), .Z(n6209) );
  OR U7078 ( .A(n6207), .B(n6206), .Z(n6208) );
  AND U7079 ( .A(n6209), .B(n6208), .Z(n6679) );
  XOR U7080 ( .A(n6678), .B(n6679), .Z(n6680) );
  XNOR U7081 ( .A(n6681), .B(n6680), .Z(n6649) );
  XNOR U7082 ( .A(n6648), .B(n6649), .Z(n6650) );
  XOR U7083 ( .A(n6651), .B(n6650), .Z(n6687) );
  ANDN U7084 ( .B(b[56]), .A(n189), .Z(n6684) );
  OR U7085 ( .A(n6211), .B(n6210), .Z(n6215) );
  NANDN U7086 ( .A(n6213), .B(n6212), .Z(n6214) );
  NAND U7087 ( .A(n6215), .B(n6214), .Z(n6685) );
  XOR U7088 ( .A(n6684), .B(n6685), .Z(n6686) );
  XNOR U7089 ( .A(n6687), .B(n6686), .Z(n6642) );
  XNOR U7090 ( .A(n6643), .B(n6642), .Z(n6644) );
  XOR U7091 ( .A(n6645), .B(n6644), .Z(n6692) );
  ANDN U7092 ( .B(b[54]), .A(n191), .Z(n6690) );
  OR U7093 ( .A(n6217), .B(n6216), .Z(n6221) );
  OR U7094 ( .A(n6219), .B(n6218), .Z(n6220) );
  AND U7095 ( .A(n6221), .B(n6220), .Z(n6691) );
  XNOR U7096 ( .A(n6690), .B(n6691), .Z(n6693) );
  XOR U7097 ( .A(n6692), .B(n6693), .Z(n6636) );
  XOR U7098 ( .A(n6639), .B(n6638), .Z(n6699) );
  ANDN U7099 ( .B(b[52]), .A(n193), .Z(n6696) );
  OR U7100 ( .A(n6223), .B(n6222), .Z(n6227) );
  OR U7101 ( .A(n6225), .B(n6224), .Z(n6226) );
  AND U7102 ( .A(n6227), .B(n6226), .Z(n6697) );
  XNOR U7103 ( .A(n6696), .B(n6697), .Z(n6698) );
  XOR U7104 ( .A(n6699), .B(n6698), .Z(n6630) );
  XOR U7105 ( .A(n6631), .B(n6630), .Z(n6632) );
  ANDN U7106 ( .B(b[50]), .A(n195), .Z(n6702) );
  OR U7107 ( .A(n6229), .B(n6228), .Z(n6233) );
  OR U7108 ( .A(n6231), .B(n6230), .Z(n6232) );
  AND U7109 ( .A(n6233), .B(n6232), .Z(n6703) );
  XNOR U7110 ( .A(n6702), .B(n6703), .Z(n6705) );
  XOR U7111 ( .A(n6704), .B(n6705), .Z(n6624) );
  XOR U7112 ( .A(n6627), .B(n6626), .Z(n6711) );
  ANDN U7113 ( .B(b[48]), .A(n197), .Z(n6708) );
  OR U7114 ( .A(n6235), .B(n6234), .Z(n6239) );
  OR U7115 ( .A(n6237), .B(n6236), .Z(n6238) );
  AND U7116 ( .A(n6239), .B(n6238), .Z(n6709) );
  XOR U7117 ( .A(n6708), .B(n6709), .Z(n6710) );
  XOR U7118 ( .A(n6619), .B(n6618), .Z(n6621) );
  XNOR U7119 ( .A(n6620), .B(n6621), .Z(n6717) );
  ANDN U7120 ( .B(b[46]), .A(n199), .Z(n6714) );
  OR U7121 ( .A(n6241), .B(n6240), .Z(n6245) );
  NANDN U7122 ( .A(n6243), .B(n6242), .Z(n6244) );
  AND U7123 ( .A(n6245), .B(n6244), .Z(n6715) );
  XNOR U7124 ( .A(n6714), .B(n6715), .Z(n6716) );
  XOR U7125 ( .A(n6717), .B(n6716), .Z(n6612) );
  XOR U7126 ( .A(n6613), .B(n6612), .Z(n6614) );
  ANDN U7127 ( .B(b[44]), .A(n201), .Z(n6720) );
  OR U7128 ( .A(n6247), .B(n6246), .Z(n6251) );
  OR U7129 ( .A(n6249), .B(n6248), .Z(n6250) );
  AND U7130 ( .A(n6251), .B(n6250), .Z(n6721) );
  XNOR U7131 ( .A(n6720), .B(n6721), .Z(n6723) );
  XOR U7132 ( .A(n6722), .B(n6723), .Z(n6606) );
  XOR U7133 ( .A(n6609), .B(n6608), .Z(n6729) );
  ANDN U7134 ( .B(b[42]), .A(n203), .Z(n6726) );
  OR U7135 ( .A(n6253), .B(n6252), .Z(n6257) );
  OR U7136 ( .A(n6255), .B(n6254), .Z(n6256) );
  AND U7137 ( .A(n6257), .B(n6256), .Z(n6727) );
  XOR U7138 ( .A(n6726), .B(n6727), .Z(n6728) );
  ANDN U7139 ( .B(b[41]), .A(n204), .Z(n6603) );
  XNOR U7140 ( .A(n6733), .B(n6732), .Z(n6734) );
  AND U7141 ( .A(a[58]), .B(b[39]), .Z(n6258) );
  NANDN U7142 ( .A(n6259), .B(n6258), .Z(n6599) );
  XOR U7143 ( .A(n6259), .B(n6258), .Z(n7026) );
  NAND U7144 ( .A(a[57]), .B(b[39]), .Z(n6593) );
  XOR U7145 ( .A(n6261), .B(n6260), .Z(n6589) );
  NAND U7146 ( .A(a[53]), .B(b[39]), .Z(n6265) );
  XNOR U7147 ( .A(n6263), .B(n6262), .Z(n6264) );
  NANDN U7148 ( .A(n6265), .B(n6264), .Z(n6575) );
  XOR U7149 ( .A(n6265), .B(n6264), .Z(n7036) );
  XNOR U7150 ( .A(n6267), .B(n6266), .Z(n6565) );
  NAND U7151 ( .A(a[50]), .B(b[39]), .Z(n6271) );
  NANDN U7152 ( .A(n6271), .B(n6270), .Z(n6563) );
  XOR U7153 ( .A(n6271), .B(n6270), .Z(n7043) );
  XNOR U7154 ( .A(n6273), .B(n6272), .Z(n6541) );
  ANDN U7155 ( .B(b[39]), .A(n192), .Z(n6531) );
  NAND U7156 ( .A(a[43]), .B(b[39]), .Z(n6525) );
  NAND U7157 ( .A(a[40]), .B(b[39]), .Z(n6509) );
  XNOR U7158 ( .A(n6277), .B(n6276), .Z(n6503) );
  NAND U7159 ( .A(a[38]), .B(b[39]), .Z(n6499) );
  XNOR U7160 ( .A(n6279), .B(n6278), .Z(n6498) );
  NANDN U7161 ( .A(n6499), .B(n6498), .Z(n6501) );
  NAND U7162 ( .A(b[39]), .B(a[37]), .Z(n6282) );
  NANDN U7163 ( .A(n6282), .B(n6283), .Z(n6497) );
  XOR U7164 ( .A(n6283), .B(n6282), .Z(n7069) );
  NAND U7165 ( .A(b[39]), .B(a[36]), .Z(n6286) );
  XNOR U7166 ( .A(n6285), .B(n6284), .Z(n6287) );
  NANDN U7167 ( .A(n6286), .B(n6287), .Z(n6495) );
  XOR U7168 ( .A(n6287), .B(n6286), .Z(n7071) );
  NAND U7169 ( .A(a[35]), .B(b[39]), .Z(n6291) );
  XOR U7170 ( .A(n6289), .B(n6288), .Z(n6290) );
  NANDN U7171 ( .A(n6291), .B(n6290), .Z(n6493) );
  XOR U7172 ( .A(n6291), .B(n6290), .Z(n7072) );
  XOR U7173 ( .A(n6293), .B(n6292), .Z(n6489) );
  XOR U7174 ( .A(n6295), .B(n6294), .Z(n6479) );
  NAND U7175 ( .A(a[27]), .B(b[39]), .Z(n6451) );
  XNOR U7176 ( .A(n6297), .B(n6296), .Z(n6450) );
  NANDN U7177 ( .A(n6451), .B(n6450), .Z(n6453) );
  XOR U7178 ( .A(n6299), .B(n6298), .Z(n6447) );
  NAND U7179 ( .A(a[23]), .B(b[39]), .Z(n6431) );
  XOR U7180 ( .A(n6301), .B(n6300), .Z(n6430) );
  NANDN U7181 ( .A(n6431), .B(n6430), .Z(n6433) );
  XOR U7182 ( .A(n6303), .B(n6302), .Z(n6426) );
  XOR U7183 ( .A(n6305), .B(n6304), .Z(n6422) );
  NAND U7184 ( .A(a[19]), .B(b[39]), .Z(n6413) );
  XNOR U7185 ( .A(n6307), .B(n6306), .Z(n6412) );
  NANDN U7186 ( .A(n6413), .B(n6412), .Z(n6415) );
  XNOR U7187 ( .A(n6309), .B(n6308), .Z(n6409) );
  AND U7188 ( .A(a[17]), .B(b[39]), .Z(n6312) );
  NANDN U7189 ( .A(n6313), .B(n6312), .Z(n6407) );
  XOR U7190 ( .A(n6313), .B(n6312), .Z(n7108) );
  NAND U7191 ( .A(a[16]), .B(b[39]), .Z(n6400) );
  NAND U7192 ( .A(a[13]), .B(b[39]), .Z(n6384) );
  OR U7193 ( .A(n6384), .B(n6385), .Z(n6387) );
  XNOR U7194 ( .A(n6317), .B(n6316), .Z(n6318) );
  ANDN U7195 ( .B(b[39]), .A(n169), .Z(n6319) );
  OR U7196 ( .A(n6318), .B(n6319), .Z(n6383) );
  XNOR U7197 ( .A(n6319), .B(n6318), .Z(n7118) );
  XNOR U7198 ( .A(n6321), .B(n6320), .Z(n6378) );
  XOR U7199 ( .A(n6323), .B(n6322), .Z(n6374) );
  XNOR U7200 ( .A(n6325), .B(n6324), .Z(n6365) );
  XOR U7201 ( .A(n6327), .B(n6326), .Z(n6329) );
  AND U7202 ( .A(a[7]), .B(b[39]), .Z(n6328) );
  NANDN U7203 ( .A(n6329), .B(n6328), .Z(n6363) );
  XOR U7204 ( .A(n6329), .B(n6328), .Z(n7128) );
  XNOR U7205 ( .A(n6331), .B(n6330), .Z(n6353) );
  XNOR U7206 ( .A(n6333), .B(n6332), .Z(n6348) );
  XNOR U7207 ( .A(n6335), .B(n6334), .Z(n6344) );
  NAND U7208 ( .A(b[40]), .B(a[1]), .Z(n6337) );
  NAND U7209 ( .A(n6337), .B(n6336), .Z(n6340) );
  OR U7210 ( .A(n6337), .B(n7536), .Z(n7143) );
  NANDN U7211 ( .A(n6339), .B(n7143), .Z(n6338) );
  AND U7212 ( .A(n6340), .B(n6338), .Z(n6343) );
  XNOR U7213 ( .A(n7143), .B(n6339), .Z(n6341) );
  NAND U7214 ( .A(n6341), .B(n6340), .Z(n7139) );
  ANDN U7215 ( .B(b[39]), .A(n162), .Z(n7138) );
  OR U7216 ( .A(n7139), .B(n7138), .Z(n6342) );
  AND U7217 ( .A(n6343), .B(n6342), .Z(n6345) );
  OR U7218 ( .A(n6344), .B(n6345), .Z(n6347) );
  XNOR U7219 ( .A(n6345), .B(n6344), .Z(n7136) );
  ANDN U7220 ( .B(b[39]), .A(n21580), .Z(n7137) );
  OR U7221 ( .A(n7136), .B(n7137), .Z(n6346) );
  AND U7222 ( .A(n6347), .B(n6346), .Z(n6349) );
  OR U7223 ( .A(n6348), .B(n6349), .Z(n6351) );
  XNOR U7224 ( .A(n6349), .B(n6348), .Z(n7134) );
  ANDN U7225 ( .B(b[39]), .A(n163), .Z(n7135) );
  OR U7226 ( .A(n7134), .B(n7135), .Z(n6350) );
  AND U7227 ( .A(n6351), .B(n6350), .Z(n6352) );
  OR U7228 ( .A(n6353), .B(n6352), .Z(n6355) );
  XNOR U7229 ( .A(n6353), .B(n6352), .Z(n7132) );
  ANDN U7230 ( .B(b[39]), .A(n164), .Z(n7133) );
  OR U7231 ( .A(n7132), .B(n7133), .Z(n6354) );
  NAND U7232 ( .A(n6355), .B(n6354), .Z(n6357) );
  AND U7233 ( .A(a[6]), .B(b[39]), .Z(n6356) );
  NANDN U7234 ( .A(n6357), .B(n6356), .Z(n6361) );
  XNOR U7235 ( .A(n6357), .B(n6356), .Z(n7130) );
  XOR U7236 ( .A(n6359), .B(n6358), .Z(n7131) );
  NAND U7237 ( .A(n7130), .B(n7131), .Z(n6360) );
  NAND U7238 ( .A(n6361), .B(n6360), .Z(n7129) );
  NANDN U7239 ( .A(n7128), .B(n7129), .Z(n6362) );
  AND U7240 ( .A(n6363), .B(n6362), .Z(n6364) );
  OR U7241 ( .A(n6365), .B(n6364), .Z(n6367) );
  XNOR U7242 ( .A(n6365), .B(n6364), .Z(n7127) );
  NAND U7243 ( .A(a[8]), .B(b[39]), .Z(n7126) );
  OR U7244 ( .A(n7127), .B(n7126), .Z(n6366) );
  NAND U7245 ( .A(n6367), .B(n6366), .Z(n6370) );
  XOR U7246 ( .A(n6369), .B(n6368), .Z(n6371) );
  OR U7247 ( .A(n6370), .B(n6371), .Z(n6373) );
  ANDN U7248 ( .B(b[39]), .A(n21615), .Z(n7125) );
  XOR U7249 ( .A(n6371), .B(n6370), .Z(n7124) );
  NANDN U7250 ( .A(n7125), .B(n7124), .Z(n6372) );
  AND U7251 ( .A(n6373), .B(n6372), .Z(n6375) );
  OR U7252 ( .A(n6374), .B(n6375), .Z(n6377) );
  XNOR U7253 ( .A(n6375), .B(n6374), .Z(n7122) );
  ANDN U7254 ( .B(b[39]), .A(n168), .Z(n7123) );
  OR U7255 ( .A(n7122), .B(n7123), .Z(n6376) );
  AND U7256 ( .A(n6377), .B(n6376), .Z(n6379) );
  OR U7257 ( .A(n6378), .B(n6379), .Z(n6381) );
  XNOR U7258 ( .A(n6379), .B(n6378), .Z(n7120) );
  ANDN U7259 ( .B(b[39]), .A(n21164), .Z(n7121) );
  OR U7260 ( .A(n7120), .B(n7121), .Z(n6380) );
  AND U7261 ( .A(n6381), .B(n6380), .Z(n7119) );
  OR U7262 ( .A(n7118), .B(n7119), .Z(n6382) );
  NAND U7263 ( .A(n6383), .B(n6382), .Z(n7117) );
  XOR U7264 ( .A(n6385), .B(n6384), .Z(n7116) );
  NANDN U7265 ( .A(n7117), .B(n7116), .Z(n6386) );
  AND U7266 ( .A(n6387), .B(n6386), .Z(n6390) );
  NANDN U7267 ( .A(n6390), .B(n6391), .Z(n6393) );
  XOR U7268 ( .A(n6391), .B(n6390), .Z(n7115) );
  NAND U7269 ( .A(a[14]), .B(b[39]), .Z(n7114) );
  OR U7270 ( .A(n7115), .B(n7114), .Z(n6392) );
  AND U7271 ( .A(n6393), .B(n6392), .Z(n6396) );
  XNOR U7272 ( .A(n6395), .B(n6394), .Z(n6397) );
  NANDN U7273 ( .A(n6396), .B(n6397), .Z(n6399) );
  NAND U7274 ( .A(a[15]), .B(b[39]), .Z(n7113) );
  XOR U7275 ( .A(n6397), .B(n6396), .Z(n7112) );
  OR U7276 ( .A(n7113), .B(n7112), .Z(n6398) );
  AND U7277 ( .A(n6399), .B(n6398), .Z(n6401) );
  OR U7278 ( .A(n6400), .B(n6401), .Z(n6405) );
  XNOR U7279 ( .A(n6401), .B(n6400), .Z(n7110) );
  NANDN U7280 ( .A(n7110), .B(n7111), .Z(n6404) );
  NAND U7281 ( .A(n6405), .B(n6404), .Z(n7109) );
  NANDN U7282 ( .A(n7108), .B(n7109), .Z(n6406) );
  AND U7283 ( .A(n6407), .B(n6406), .Z(n6408) );
  OR U7284 ( .A(n6409), .B(n6408), .Z(n6411) );
  XNOR U7285 ( .A(n6409), .B(n6408), .Z(n7107) );
  NAND U7286 ( .A(a[18]), .B(b[39]), .Z(n7106) );
  OR U7287 ( .A(n7107), .B(n7106), .Z(n6410) );
  AND U7288 ( .A(n6411), .B(n6410), .Z(n7104) );
  NANDN U7289 ( .A(n7104), .B(n7105), .Z(n6414) );
  NAND U7290 ( .A(n6415), .B(n6414), .Z(n6418) );
  XOR U7291 ( .A(n6417), .B(n6416), .Z(n6419) );
  OR U7292 ( .A(n6418), .B(n6419), .Z(n6421) );
  ANDN U7293 ( .B(b[39]), .A(n176), .Z(n7102) );
  XOR U7294 ( .A(n6419), .B(n6418), .Z(n7103) );
  NANDN U7295 ( .A(n7102), .B(n7103), .Z(n6420) );
  AND U7296 ( .A(n6421), .B(n6420), .Z(n6423) );
  OR U7297 ( .A(n6422), .B(n6423), .Z(n6425) );
  XNOR U7298 ( .A(n6423), .B(n6422), .Z(n7100) );
  ANDN U7299 ( .B(b[39]), .A(n21681), .Z(n7101) );
  OR U7300 ( .A(n7100), .B(n7101), .Z(n6424) );
  AND U7301 ( .A(n6425), .B(n6424), .Z(n6427) );
  OR U7302 ( .A(n6426), .B(n6427), .Z(n6429) );
  XNOR U7303 ( .A(n6427), .B(n6426), .Z(n7098) );
  ANDN U7304 ( .B(b[39]), .A(n177), .Z(n7099) );
  OR U7305 ( .A(n7098), .B(n7099), .Z(n6428) );
  NAND U7306 ( .A(n6429), .B(n6428), .Z(n7096) );
  NANDN U7307 ( .A(n7096), .B(n7097), .Z(n6432) );
  AND U7308 ( .A(n6433), .B(n6432), .Z(n6436) );
  NANDN U7309 ( .A(n6436), .B(n6437), .Z(n6439) );
  XOR U7310 ( .A(n6437), .B(n6436), .Z(n7095) );
  NAND U7311 ( .A(a[24]), .B(b[39]), .Z(n7094) );
  OR U7312 ( .A(n7095), .B(n7094), .Z(n6438) );
  NAND U7313 ( .A(n6439), .B(n6438), .Z(n6442) );
  XOR U7314 ( .A(n6441), .B(n6440), .Z(n6443) );
  OR U7315 ( .A(n6442), .B(n6443), .Z(n6445) );
  ANDN U7316 ( .B(b[39]), .A(n21703), .Z(n7093) );
  XOR U7317 ( .A(n6443), .B(n6442), .Z(n7092) );
  NANDN U7318 ( .A(n7093), .B(n7092), .Z(n6444) );
  NAND U7319 ( .A(n6445), .B(n6444), .Z(n6446) );
  NANDN U7320 ( .A(n6447), .B(n6446), .Z(n6449) );
  ANDN U7321 ( .B(b[39]), .A(n179), .Z(n7091) );
  NANDN U7322 ( .A(n7091), .B(n7090), .Z(n6448) );
  NAND U7323 ( .A(n6449), .B(n6448), .Z(n7089) );
  NANDN U7324 ( .A(n7089), .B(n7088), .Z(n6452) );
  NAND U7325 ( .A(n6453), .B(n6452), .Z(n6457) );
  XOR U7326 ( .A(n6455), .B(n6454), .Z(n6456) );
  NANDN U7327 ( .A(n6457), .B(n6456), .Z(n6459) );
  ANDN U7328 ( .B(b[39]), .A(n180), .Z(n7087) );
  XOR U7329 ( .A(n6457), .B(n6456), .Z(n7086) );
  OR U7330 ( .A(n7087), .B(n7086), .Z(n6458) );
  NAND U7331 ( .A(n6459), .B(n6458), .Z(n6463) );
  NAND U7332 ( .A(b[39]), .B(a[29]), .Z(n6462) );
  OR U7333 ( .A(n6463), .B(n6462), .Z(n6465) );
  XOR U7334 ( .A(n6463), .B(n6462), .Z(n7084) );
  NAND U7335 ( .A(n7085), .B(n7084), .Z(n6464) );
  NAND U7336 ( .A(n6465), .B(n6464), .Z(n6469) );
  XOR U7337 ( .A(n6467), .B(n6466), .Z(n6468) );
  NANDN U7338 ( .A(n6469), .B(n6468), .Z(n6471) );
  ANDN U7339 ( .B(b[39]), .A(n181), .Z(n7083) );
  XOR U7340 ( .A(n6469), .B(n6468), .Z(n7082) );
  OR U7341 ( .A(n7083), .B(n7082), .Z(n6470) );
  NAND U7342 ( .A(n6471), .B(n6470), .Z(n6475) );
  NANDN U7343 ( .A(n6475), .B(n6474), .Z(n6477) );
  XOR U7344 ( .A(n6475), .B(n6474), .Z(n7080) );
  NAND U7345 ( .A(a[31]), .B(b[39]), .Z(n7081) );
  OR U7346 ( .A(n7080), .B(n7081), .Z(n6476) );
  NAND U7347 ( .A(n6477), .B(n6476), .Z(n6478) );
  NANDN U7348 ( .A(n6479), .B(n6478), .Z(n6481) );
  XOR U7349 ( .A(n6479), .B(n6478), .Z(n7079) );
  NAND U7350 ( .A(a[32]), .B(b[39]), .Z(n7078) );
  OR U7351 ( .A(n7079), .B(n7078), .Z(n6480) );
  NAND U7352 ( .A(n6481), .B(n6480), .Z(n6484) );
  NANDN U7353 ( .A(n6484), .B(n6485), .Z(n6487) );
  ANDN U7354 ( .B(b[39]), .A(n21751), .Z(n7077) );
  XOR U7355 ( .A(n6485), .B(n6484), .Z(n7076) );
  OR U7356 ( .A(n7077), .B(n7076), .Z(n6486) );
  NAND U7357 ( .A(n6487), .B(n6486), .Z(n6488) );
  NANDN U7358 ( .A(n6489), .B(n6488), .Z(n6491) );
  ANDN U7359 ( .B(b[39]), .A(n183), .Z(n7075) );
  NANDN U7360 ( .A(n7075), .B(n7074), .Z(n6490) );
  NAND U7361 ( .A(n6491), .B(n6490), .Z(n7073) );
  OR U7362 ( .A(n7072), .B(n7073), .Z(n6492) );
  AND U7363 ( .A(n6493), .B(n6492), .Z(n7070) );
  OR U7364 ( .A(n7071), .B(n7070), .Z(n6494) );
  AND U7365 ( .A(n6495), .B(n6494), .Z(n7068) );
  OR U7366 ( .A(n7069), .B(n7068), .Z(n6496) );
  AND U7367 ( .A(n6497), .B(n6496), .Z(n7066) );
  NANDN U7368 ( .A(n7066), .B(n7067), .Z(n6500) );
  NAND U7369 ( .A(n6501), .B(n6500), .Z(n6502) );
  NANDN U7370 ( .A(n6503), .B(n6502), .Z(n6505) );
  NAND U7371 ( .A(a[39]), .B(b[39]), .Z(n7065) );
  NANDN U7372 ( .A(n7065), .B(n7064), .Z(n6504) );
  NAND U7373 ( .A(n6505), .B(n6504), .Z(n6508) );
  NANDN U7374 ( .A(n6509), .B(n6508), .Z(n6511) );
  XOR U7375 ( .A(n6507), .B(n6506), .Z(n7062) );
  NANDN U7376 ( .A(n7062), .B(n7063), .Z(n6510) );
  NAND U7377 ( .A(n6511), .B(n6510), .Z(n6515) );
  XOR U7378 ( .A(n6513), .B(n6512), .Z(n6514) );
  NANDN U7379 ( .A(n6515), .B(n6514), .Z(n6517) );
  ANDN U7380 ( .B(b[39]), .A(n189), .Z(n7061) );
  XOR U7381 ( .A(n6515), .B(n6514), .Z(n7060) );
  OR U7382 ( .A(n7061), .B(n7060), .Z(n6516) );
  NAND U7383 ( .A(n6517), .B(n6516), .Z(n6519) );
  OR U7384 ( .A(n6518), .B(n6519), .Z(n6521) );
  NAND U7385 ( .A(a[42]), .B(b[39]), .Z(n7059) );
  XOR U7386 ( .A(n6519), .B(n6518), .Z(n7058) );
  NANDN U7387 ( .A(n7059), .B(n7058), .Z(n6520) );
  NAND U7388 ( .A(n6521), .B(n6520), .Z(n6524) );
  NANDN U7389 ( .A(n6525), .B(n6524), .Z(n6527) );
  XOR U7390 ( .A(n6523), .B(n6522), .Z(n7056) );
  NANDN U7391 ( .A(n7056), .B(n7057), .Z(n6526) );
  NAND U7392 ( .A(n6527), .B(n6526), .Z(n6530) );
  OR U7393 ( .A(n6531), .B(n6530), .Z(n6533) );
  XNOR U7394 ( .A(n6529), .B(n6528), .Z(n7055) );
  XOR U7395 ( .A(n6531), .B(n6530), .Z(n7054) );
  NANDN U7396 ( .A(n7055), .B(n7054), .Z(n6532) );
  NAND U7397 ( .A(n6533), .B(n6532), .Z(n6537) );
  NANDN U7398 ( .A(n6537), .B(n6536), .Z(n6539) );
  XOR U7399 ( .A(n6537), .B(n6536), .Z(n7052) );
  NAND U7400 ( .A(a[45]), .B(b[39]), .Z(n7053) );
  OR U7401 ( .A(n7052), .B(n7053), .Z(n6538) );
  NAND U7402 ( .A(n6539), .B(n6538), .Z(n6540) );
  NANDN U7403 ( .A(n6541), .B(n6540), .Z(n6543) );
  NAND U7404 ( .A(a[46]), .B(b[39]), .Z(n7050) );
  NANDN U7405 ( .A(n7050), .B(n7051), .Z(n6542) );
  AND U7406 ( .A(n6543), .B(n6542), .Z(n6546) );
  NAND U7407 ( .A(n6546), .B(n6547), .Z(n6549) );
  ANDN U7408 ( .B(b[39]), .A(n195), .Z(n7049) );
  XNOR U7409 ( .A(n6547), .B(n6546), .Z(n7048) );
  OR U7410 ( .A(n7049), .B(n7048), .Z(n6548) );
  NAND U7411 ( .A(n6549), .B(n6548), .Z(n6553) );
  XNOR U7412 ( .A(n6551), .B(n6550), .Z(n6552) );
  NANDN U7413 ( .A(n6553), .B(n6552), .Z(n6555) );
  XOR U7414 ( .A(n6553), .B(n6552), .Z(n7046) );
  NAND U7415 ( .A(a[48]), .B(b[39]), .Z(n7047) );
  OR U7416 ( .A(n7046), .B(n7047), .Z(n6554) );
  NAND U7417 ( .A(n6555), .B(n6554), .Z(n6558) );
  XOR U7418 ( .A(n6557), .B(n6556), .Z(n6559) );
  NAND U7419 ( .A(n6558), .B(n6559), .Z(n6561) );
  XNOR U7420 ( .A(n6559), .B(n6558), .Z(n7045) );
  NAND U7421 ( .A(a[49]), .B(b[39]), .Z(n7044) );
  OR U7422 ( .A(n7045), .B(n7044), .Z(n6560) );
  AND U7423 ( .A(n6561), .B(n6560), .Z(n7042) );
  OR U7424 ( .A(n7043), .B(n7042), .Z(n6562) );
  NAND U7425 ( .A(n6563), .B(n6562), .Z(n6564) );
  NANDN U7426 ( .A(n6565), .B(n6564), .Z(n6567) );
  NAND U7427 ( .A(a[51]), .B(b[39]), .Z(n7040) );
  NANDN U7428 ( .A(n7040), .B(n7041), .Z(n6566) );
  NAND U7429 ( .A(n6567), .B(n6566), .Z(n6571) );
  XOR U7430 ( .A(n6569), .B(n6568), .Z(n6570) );
  NANDN U7431 ( .A(n6571), .B(n6570), .Z(n6573) );
  ANDN U7432 ( .B(b[39]), .A(n200), .Z(n7039) );
  XOR U7433 ( .A(n6571), .B(n6570), .Z(n7038) );
  OR U7434 ( .A(n7039), .B(n7038), .Z(n6572) );
  NAND U7435 ( .A(n6573), .B(n6572), .Z(n7037) );
  OR U7436 ( .A(n7036), .B(n7037), .Z(n6574) );
  NAND U7437 ( .A(n6575), .B(n6574), .Z(n6579) );
  XOR U7438 ( .A(n6577), .B(n6576), .Z(n6578) );
  NANDN U7439 ( .A(n6579), .B(n6578), .Z(n6581) );
  ANDN U7440 ( .B(b[39]), .A(n202), .Z(n7035) );
  NANDN U7441 ( .A(n7035), .B(n7034), .Z(n6580) );
  NAND U7442 ( .A(n6581), .B(n6580), .Z(n6584) );
  NANDN U7443 ( .A(n6584), .B(n6585), .Z(n6587) );
  NAND U7444 ( .A(a[55]), .B(b[39]), .Z(n7033) );
  XOR U7445 ( .A(n6585), .B(n6584), .Z(n7032) );
  OR U7446 ( .A(n7033), .B(n7032), .Z(n6586) );
  AND U7447 ( .A(n6587), .B(n6586), .Z(n6588) );
  OR U7448 ( .A(n6589), .B(n6588), .Z(n6591) );
  XNOR U7449 ( .A(n6589), .B(n6588), .Z(n7031) );
  NAND U7450 ( .A(a[56]), .B(b[39]), .Z(n7030) );
  OR U7451 ( .A(n7031), .B(n7030), .Z(n6590) );
  AND U7452 ( .A(n6591), .B(n6590), .Z(n6592) );
  OR U7453 ( .A(n6593), .B(n6592), .Z(n6597) );
  XNOR U7454 ( .A(n6593), .B(n6592), .Z(n7028) );
  XOR U7455 ( .A(n6595), .B(n6594), .Z(n7029) );
  OR U7456 ( .A(n7028), .B(n7029), .Z(n6596) );
  NAND U7457 ( .A(n6597), .B(n6596), .Z(n7027) );
  NANDN U7458 ( .A(n7026), .B(n7027), .Z(n6598) );
  AND U7459 ( .A(n6599), .B(n6598), .Z(n6739) );
  NAND U7460 ( .A(b[40]), .B(a[58]), .Z(n6876) );
  ANDN U7461 ( .B(b[41]), .A(n205), .Z(n6744) );
  NANDN U7462 ( .A(n6601), .B(n6600), .Z(n6605) );
  NANDN U7463 ( .A(n6603), .B(n6602), .Z(n6604) );
  AND U7464 ( .A(n6605), .B(n6604), .Z(n6743) );
  ANDN U7465 ( .B(b[43]), .A(n203), .Z(n6750) );
  NANDN U7466 ( .A(n6607), .B(n6606), .Z(n6611) );
  NANDN U7467 ( .A(n6609), .B(n6608), .Z(n6610) );
  AND U7468 ( .A(n6611), .B(n6610), .Z(n6749) );
  NAND U7469 ( .A(a[53]), .B(b[45]), .Z(n6757) );
  OR U7470 ( .A(n6613), .B(n6612), .Z(n6617) );
  NANDN U7471 ( .A(n6615), .B(n6614), .Z(n6616) );
  AND U7472 ( .A(n6617), .B(n6616), .Z(n6754) );
  ANDN U7473 ( .B(b[47]), .A(n199), .Z(n6762) );
  NANDN U7474 ( .A(n6619), .B(n6618), .Z(n6623) );
  OR U7475 ( .A(n6621), .B(n6620), .Z(n6622) );
  AND U7476 ( .A(n6623), .B(n6622), .Z(n6761) );
  ANDN U7477 ( .B(b[49]), .A(n197), .Z(n6768) );
  NANDN U7478 ( .A(n6625), .B(n6624), .Z(n6629) );
  NANDN U7479 ( .A(n6627), .B(n6626), .Z(n6628) );
  AND U7480 ( .A(n6629), .B(n6628), .Z(n6767) );
  NAND U7481 ( .A(a[47]), .B(b[51]), .Z(n6775) );
  OR U7482 ( .A(n6631), .B(n6630), .Z(n6635) );
  NANDN U7483 ( .A(n6633), .B(n6632), .Z(n6634) );
  AND U7484 ( .A(n6635), .B(n6634), .Z(n6772) );
  ANDN U7485 ( .B(b[53]), .A(n193), .Z(n6780) );
  NANDN U7486 ( .A(n6637), .B(n6636), .Z(n6641) );
  NANDN U7487 ( .A(n6639), .B(n6638), .Z(n6640) );
  AND U7488 ( .A(n6641), .B(n6640), .Z(n6779) );
  NAND U7489 ( .A(a[43]), .B(b[55]), .Z(n6787) );
  OR U7490 ( .A(n6643), .B(n6642), .Z(n6647) );
  OR U7491 ( .A(n6645), .B(n6644), .Z(n6646) );
  AND U7492 ( .A(n6647), .B(n6646), .Z(n6784) );
  NAND U7493 ( .A(a[41]), .B(b[57]), .Z(n6793) );
  OR U7494 ( .A(n6649), .B(n6648), .Z(n6653) );
  OR U7495 ( .A(n6651), .B(n6650), .Z(n6652) );
  AND U7496 ( .A(n6653), .B(n6652), .Z(n6790) );
  ANDN U7497 ( .B(b[59]), .A(n187), .Z(n6799) );
  OR U7498 ( .A(n6655), .B(n6654), .Z(n6659) );
  NANDN U7499 ( .A(n6657), .B(n6656), .Z(n6658) );
  NAND U7500 ( .A(n6659), .B(n6658), .Z(n6797) );
  ANDN U7501 ( .B(b[61]), .A(n21772), .Z(n6804) );
  OR U7502 ( .A(n6661), .B(n6660), .Z(n6665) );
  OR U7503 ( .A(n6663), .B(n6662), .Z(n6664) );
  AND U7504 ( .A(n6665), .B(n6664), .Z(n6802) );
  ANDN U7505 ( .B(b[63]), .A(n184), .Z(n6810) );
  ANDN U7506 ( .B(a[36]), .A(n159), .Z(n6808) );
  OR U7507 ( .A(n6667), .B(n6666), .Z(n6671) );
  OR U7508 ( .A(n6669), .B(n6668), .Z(n6670) );
  AND U7509 ( .A(n6671), .B(n6670), .Z(n6809) );
  XNOR U7510 ( .A(n6808), .B(n6809), .Z(n6811) );
  XNOR U7511 ( .A(n6810), .B(n6811), .Z(n6803) );
  XNOR U7512 ( .A(n6802), .B(n6803), .Z(n6805) );
  XNOR U7513 ( .A(n6804), .B(n6805), .Z(n6817) );
  ANDN U7514 ( .B(b[60]), .A(n186), .Z(n6814) );
  OR U7515 ( .A(n6673), .B(n6672), .Z(n6677) );
  OR U7516 ( .A(n6675), .B(n6674), .Z(n6676) );
  AND U7517 ( .A(n6677), .B(n6676), .Z(n6815) );
  XOR U7518 ( .A(n6814), .B(n6815), .Z(n6816) );
  XOR U7519 ( .A(n6799), .B(n6798), .Z(n6823) );
  ANDN U7520 ( .B(b[58]), .A(n188), .Z(n6820) );
  OR U7521 ( .A(n6679), .B(n6678), .Z(n6683) );
  NANDN U7522 ( .A(n6681), .B(n6680), .Z(n6682) );
  AND U7523 ( .A(n6683), .B(n6682), .Z(n6821) );
  XNOR U7524 ( .A(n6820), .B(n6821), .Z(n6822) );
  XOR U7525 ( .A(n6823), .B(n6822), .Z(n6791) );
  XNOR U7526 ( .A(n6790), .B(n6791), .Z(n6792) );
  XOR U7527 ( .A(n6793), .B(n6792), .Z(n6829) );
  ANDN U7528 ( .B(b[56]), .A(n190), .Z(n6826) );
  OR U7529 ( .A(n6685), .B(n6684), .Z(n6689) );
  NANDN U7530 ( .A(n6687), .B(n6686), .Z(n6688) );
  AND U7531 ( .A(n6689), .B(n6688), .Z(n6827) );
  XOR U7532 ( .A(n6826), .B(n6827), .Z(n6828) );
  XNOR U7533 ( .A(n6829), .B(n6828), .Z(n6785) );
  XNOR U7534 ( .A(n6784), .B(n6785), .Z(n6786) );
  XOR U7535 ( .A(n6787), .B(n6786), .Z(n6834) );
  ANDN U7536 ( .B(b[54]), .A(n192), .Z(n6832) );
  OR U7537 ( .A(n6691), .B(n6690), .Z(n6695) );
  OR U7538 ( .A(n6693), .B(n6692), .Z(n6694) );
  AND U7539 ( .A(n6695), .B(n6694), .Z(n6833) );
  XNOR U7540 ( .A(n6832), .B(n6833), .Z(n6835) );
  XOR U7541 ( .A(n6834), .B(n6835), .Z(n6778) );
  XOR U7542 ( .A(n6779), .B(n6778), .Z(n6781) );
  XNOR U7543 ( .A(n6780), .B(n6781), .Z(n6841) );
  ANDN U7544 ( .B(b[52]), .A(n194), .Z(n6838) );
  OR U7545 ( .A(n6697), .B(n6696), .Z(n6701) );
  OR U7546 ( .A(n6699), .B(n6698), .Z(n6700) );
  AND U7547 ( .A(n6701), .B(n6700), .Z(n6839) );
  XNOR U7548 ( .A(n6838), .B(n6839), .Z(n6840) );
  XOR U7549 ( .A(n6841), .B(n6840), .Z(n6773) );
  XNOR U7550 ( .A(n6772), .B(n6773), .Z(n6774) );
  XOR U7551 ( .A(n6775), .B(n6774), .Z(n6846) );
  ANDN U7552 ( .B(b[50]), .A(n196), .Z(n6844) );
  OR U7553 ( .A(n6703), .B(n6702), .Z(n6707) );
  OR U7554 ( .A(n6705), .B(n6704), .Z(n6706) );
  AND U7555 ( .A(n6707), .B(n6706), .Z(n6845) );
  XNOR U7556 ( .A(n6844), .B(n6845), .Z(n6847) );
  XOR U7557 ( .A(n6846), .B(n6847), .Z(n6766) );
  XOR U7558 ( .A(n6767), .B(n6766), .Z(n6769) );
  XNOR U7559 ( .A(n6768), .B(n6769), .Z(n6853) );
  ANDN U7560 ( .B(b[48]), .A(n198), .Z(n6850) );
  OR U7561 ( .A(n6709), .B(n6708), .Z(n6713) );
  NANDN U7562 ( .A(n6711), .B(n6710), .Z(n6712) );
  AND U7563 ( .A(n6713), .B(n6712), .Z(n6851) );
  XOR U7564 ( .A(n6850), .B(n6851), .Z(n6852) );
  XOR U7565 ( .A(n6761), .B(n6760), .Z(n6763) );
  XNOR U7566 ( .A(n6762), .B(n6763), .Z(n6859) );
  ANDN U7567 ( .B(b[46]), .A(n200), .Z(n6856) );
  OR U7568 ( .A(n6715), .B(n6714), .Z(n6719) );
  OR U7569 ( .A(n6717), .B(n6716), .Z(n6718) );
  AND U7570 ( .A(n6719), .B(n6718), .Z(n6857) );
  XNOR U7571 ( .A(n6856), .B(n6857), .Z(n6858) );
  XOR U7572 ( .A(n6859), .B(n6858), .Z(n6755) );
  XNOR U7573 ( .A(n6754), .B(n6755), .Z(n6756) );
  XOR U7574 ( .A(n6757), .B(n6756), .Z(n6864) );
  ANDN U7575 ( .B(b[44]), .A(n202), .Z(n6862) );
  OR U7576 ( .A(n6721), .B(n6720), .Z(n6725) );
  OR U7577 ( .A(n6723), .B(n6722), .Z(n6724) );
  AND U7578 ( .A(n6725), .B(n6724), .Z(n6863) );
  XNOR U7579 ( .A(n6862), .B(n6863), .Z(n6865) );
  XOR U7580 ( .A(n6864), .B(n6865), .Z(n6748) );
  XOR U7581 ( .A(n6749), .B(n6748), .Z(n6751) );
  XNOR U7582 ( .A(n6750), .B(n6751), .Z(n6871) );
  ANDN U7583 ( .B(b[42]), .A(n204), .Z(n6868) );
  OR U7584 ( .A(n6727), .B(n6726), .Z(n6731) );
  NANDN U7585 ( .A(n6729), .B(n6728), .Z(n6730) );
  AND U7586 ( .A(n6731), .B(n6730), .Z(n6869) );
  XOR U7587 ( .A(n6868), .B(n6869), .Z(n6870) );
  XOR U7588 ( .A(n6743), .B(n6742), .Z(n6745) );
  XNOR U7589 ( .A(n6744), .B(n6745), .Z(n6875) );
  NANDN U7590 ( .A(n6733), .B(n6732), .Z(n6737) );
  NANDN U7591 ( .A(n6735), .B(n6734), .Z(n6736) );
  NAND U7592 ( .A(n6737), .B(n6736), .Z(n6874) );
  XNOR U7593 ( .A(n6875), .B(n6874), .Z(n6877) );
  XOR U7594 ( .A(n6876), .B(n6877), .Z(n6738) );
  NANDN U7595 ( .A(n6739), .B(n6738), .Z(n6741) );
  NAND U7596 ( .A(a[59]), .B(b[39]), .Z(n7025) );
  XOR U7597 ( .A(n6739), .B(n6738), .Z(n7024) );
  OR U7598 ( .A(n7025), .B(n7024), .Z(n6740) );
  NAND U7599 ( .A(n6741), .B(n6740), .Z(n6881) );
  NAND U7600 ( .A(a[58]), .B(b[41]), .Z(n6887) );
  NANDN U7601 ( .A(n6743), .B(n6742), .Z(n6747) );
  OR U7602 ( .A(n6745), .B(n6744), .Z(n6746) );
  NAND U7603 ( .A(n6747), .B(n6746), .Z(n6885) );
  NAND U7604 ( .A(a[56]), .B(b[43]), .Z(n6893) );
  NANDN U7605 ( .A(n6749), .B(n6748), .Z(n6753) );
  OR U7606 ( .A(n6751), .B(n6750), .Z(n6752) );
  NAND U7607 ( .A(n6753), .B(n6752), .Z(n6891) );
  ANDN U7608 ( .B(b[45]), .A(n202), .Z(n7007) );
  OR U7609 ( .A(n6755), .B(n6754), .Z(n6759) );
  OR U7610 ( .A(n6757), .B(n6756), .Z(n6758) );
  NAND U7611 ( .A(n6759), .B(n6758), .Z(n7005) );
  ANDN U7612 ( .B(b[47]), .A(n200), .Z(n6910) );
  NANDN U7613 ( .A(n6761), .B(n6760), .Z(n6765) );
  OR U7614 ( .A(n6763), .B(n6762), .Z(n6764) );
  AND U7615 ( .A(n6765), .B(n6764), .Z(n6909) );
  NAND U7616 ( .A(a[50]), .B(b[49]), .Z(n7001) );
  NANDN U7617 ( .A(n6767), .B(n6766), .Z(n6771) );
  OR U7618 ( .A(n6769), .B(n6768), .Z(n6770) );
  NAND U7619 ( .A(n6771), .B(n6770), .Z(n6999) );
  ANDN U7620 ( .B(b[51]), .A(n196), .Z(n6923) );
  OR U7621 ( .A(n6773), .B(n6772), .Z(n6777) );
  OR U7622 ( .A(n6775), .B(n6774), .Z(n6776) );
  NAND U7623 ( .A(n6777), .B(n6776), .Z(n6921) );
  NAND U7624 ( .A(a[46]), .B(b[53]), .Z(n6929) );
  NANDN U7625 ( .A(n6779), .B(n6778), .Z(n6783) );
  OR U7626 ( .A(n6781), .B(n6780), .Z(n6782) );
  NAND U7627 ( .A(n6783), .B(n6782), .Z(n6927) );
  NAND U7628 ( .A(a[44]), .B(b[55]), .Z(n6983) );
  OR U7629 ( .A(n6785), .B(n6784), .Z(n6789) );
  OR U7630 ( .A(n6787), .B(n6786), .Z(n6788) );
  AND U7631 ( .A(n6789), .B(n6788), .Z(n6980) );
  NAND U7632 ( .A(a[42]), .B(b[57]), .Z(n6947) );
  OR U7633 ( .A(n6791), .B(n6790), .Z(n6795) );
  OR U7634 ( .A(n6793), .B(n6792), .Z(n6794) );
  AND U7635 ( .A(n6795), .B(n6794), .Z(n6944) );
  NAND U7636 ( .A(a[40]), .B(b[59]), .Z(n6977) );
  NANDN U7637 ( .A(n6797), .B(n6796), .Z(n6801) );
  NANDN U7638 ( .A(n6799), .B(n6798), .Z(n6800) );
  NAND U7639 ( .A(n6801), .B(n6800), .Z(n6975) );
  ANDN U7640 ( .B(b[61]), .A(n186), .Z(n6958) );
  OR U7641 ( .A(n6803), .B(n6802), .Z(n6807) );
  OR U7642 ( .A(n6805), .B(n6804), .Z(n6806) );
  AND U7643 ( .A(n6807), .B(n6806), .Z(n6956) );
  ANDN U7644 ( .B(b[63]), .A(n185), .Z(n6964) );
  ANDN U7645 ( .B(a[37]), .A(n159), .Z(n6962) );
  OR U7646 ( .A(n6809), .B(n6808), .Z(n6813) );
  OR U7647 ( .A(n6811), .B(n6810), .Z(n6812) );
  AND U7648 ( .A(n6813), .B(n6812), .Z(n6963) );
  XNOR U7649 ( .A(n6962), .B(n6963), .Z(n6965) );
  XNOR U7650 ( .A(n6964), .B(n6965), .Z(n6957) );
  XNOR U7651 ( .A(n6956), .B(n6957), .Z(n6959) );
  XNOR U7652 ( .A(n6958), .B(n6959), .Z(n6971) );
  ANDN U7653 ( .B(b[60]), .A(n187), .Z(n6968) );
  OR U7654 ( .A(n6815), .B(n6814), .Z(n6819) );
  NANDN U7655 ( .A(n6817), .B(n6816), .Z(n6818) );
  AND U7656 ( .A(n6819), .B(n6818), .Z(n6969) );
  XNOR U7657 ( .A(n6968), .B(n6969), .Z(n6970) );
  XOR U7658 ( .A(n6971), .B(n6970), .Z(n6974) );
  XOR U7659 ( .A(n6975), .B(n6974), .Z(n6976) );
  ANDN U7660 ( .B(b[58]), .A(n189), .Z(n6950) );
  OR U7661 ( .A(n6821), .B(n6820), .Z(n6825) );
  OR U7662 ( .A(n6823), .B(n6822), .Z(n6824) );
  AND U7663 ( .A(n6825), .B(n6824), .Z(n6951) );
  XOR U7664 ( .A(n6950), .B(n6951), .Z(n6952) );
  XNOR U7665 ( .A(n6953), .B(n6952), .Z(n6945) );
  XNOR U7666 ( .A(n6944), .B(n6945), .Z(n6946) );
  XOR U7667 ( .A(n6947), .B(n6946), .Z(n6941) );
  ANDN U7668 ( .B(b[56]), .A(n191), .Z(n6938) );
  OR U7669 ( .A(n6827), .B(n6826), .Z(n6831) );
  NANDN U7670 ( .A(n6829), .B(n6828), .Z(n6830) );
  AND U7671 ( .A(n6831), .B(n6830), .Z(n6939) );
  XOR U7672 ( .A(n6938), .B(n6939), .Z(n6940) );
  XNOR U7673 ( .A(n6941), .B(n6940), .Z(n6981) );
  XNOR U7674 ( .A(n6980), .B(n6981), .Z(n6982) );
  XOR U7675 ( .A(n6983), .B(n6982), .Z(n6935) );
  ANDN U7676 ( .B(b[54]), .A(n193), .Z(n6932) );
  OR U7677 ( .A(n6833), .B(n6832), .Z(n6837) );
  OR U7678 ( .A(n6835), .B(n6834), .Z(n6836) );
  AND U7679 ( .A(n6837), .B(n6836), .Z(n6933) );
  XOR U7680 ( .A(n6932), .B(n6933), .Z(n6934) );
  XNOR U7681 ( .A(n6935), .B(n6934), .Z(n6926) );
  XNOR U7682 ( .A(n6927), .B(n6926), .Z(n6928) );
  XOR U7683 ( .A(n6929), .B(n6928), .Z(n6988) );
  ANDN U7684 ( .B(b[52]), .A(n195), .Z(n6986) );
  OR U7685 ( .A(n6839), .B(n6838), .Z(n6843) );
  OR U7686 ( .A(n6841), .B(n6840), .Z(n6842) );
  AND U7687 ( .A(n6843), .B(n6842), .Z(n6987) );
  XNOR U7688 ( .A(n6986), .B(n6987), .Z(n6989) );
  XOR U7689 ( .A(n6988), .B(n6989), .Z(n6920) );
  XOR U7690 ( .A(n6923), .B(n6922), .Z(n6995) );
  ANDN U7691 ( .B(b[50]), .A(n197), .Z(n6992) );
  OR U7692 ( .A(n6845), .B(n6844), .Z(n6849) );
  OR U7693 ( .A(n6847), .B(n6846), .Z(n6848) );
  AND U7694 ( .A(n6849), .B(n6848), .Z(n6993) );
  XNOR U7695 ( .A(n6992), .B(n6993), .Z(n6994) );
  XOR U7696 ( .A(n6995), .B(n6994), .Z(n6998) );
  XOR U7697 ( .A(n6999), .B(n6998), .Z(n7000) );
  ANDN U7698 ( .B(b[48]), .A(n199), .Z(n6914) );
  OR U7699 ( .A(n6851), .B(n6850), .Z(n6855) );
  NANDN U7700 ( .A(n6853), .B(n6852), .Z(n6854) );
  AND U7701 ( .A(n6855), .B(n6854), .Z(n6915) );
  XNOR U7702 ( .A(n6914), .B(n6915), .Z(n6917) );
  XOR U7703 ( .A(n6916), .B(n6917), .Z(n6908) );
  XOR U7704 ( .A(n6909), .B(n6908), .Z(n6911) );
  XNOR U7705 ( .A(n6910), .B(n6911), .Z(n6905) );
  ANDN U7706 ( .B(b[46]), .A(n201), .Z(n6902) );
  OR U7707 ( .A(n6857), .B(n6856), .Z(n6861) );
  OR U7708 ( .A(n6859), .B(n6858), .Z(n6860) );
  AND U7709 ( .A(n6861), .B(n6860), .Z(n6903) );
  XOR U7710 ( .A(n6902), .B(n6903), .Z(n6904) );
  XOR U7711 ( .A(n7007), .B(n7006), .Z(n6899) );
  ANDN U7712 ( .B(b[44]), .A(n203), .Z(n6896) );
  OR U7713 ( .A(n6863), .B(n6862), .Z(n6867) );
  OR U7714 ( .A(n6865), .B(n6864), .Z(n6866) );
  AND U7715 ( .A(n6867), .B(n6866), .Z(n6897) );
  XNOR U7716 ( .A(n6896), .B(n6897), .Z(n6898) );
  XOR U7717 ( .A(n6899), .B(n6898), .Z(n6890) );
  XOR U7718 ( .A(n6891), .B(n6890), .Z(n6892) );
  ANDN U7719 ( .B(b[42]), .A(n205), .Z(n7010) );
  OR U7720 ( .A(n6869), .B(n6868), .Z(n6873) );
  NANDN U7721 ( .A(n6871), .B(n6870), .Z(n6872) );
  AND U7722 ( .A(n6873), .B(n6872), .Z(n7011) );
  XOR U7723 ( .A(n7010), .B(n7011), .Z(n7012) );
  XNOR U7724 ( .A(n7013), .B(n7012), .Z(n6884) );
  XNOR U7725 ( .A(n6885), .B(n6884), .Z(n6886) );
  XOR U7726 ( .A(n6887), .B(n6886), .Z(n7018) );
  ANDN U7727 ( .B(b[40]), .A(n207), .Z(n7016) );
  OR U7728 ( .A(n6875), .B(n6874), .Z(n6879) );
  NANDN U7729 ( .A(n6877), .B(n6876), .Z(n6878) );
  AND U7730 ( .A(n6879), .B(n6878), .Z(n7017) );
  XNOR U7731 ( .A(n7016), .B(n7017), .Z(n7019) );
  XOR U7732 ( .A(n7018), .B(n7019), .Z(n6880) );
  NANDN U7733 ( .A(n6881), .B(n6880), .Z(n6883) );
  ANDN U7734 ( .B(b[39]), .A(n208), .Z(n7023) );
  NANDN U7735 ( .A(n7023), .B(n7022), .Z(n6882) );
  NAND U7736 ( .A(n6883), .B(n6882), .Z(n7527) );
  NAND U7737 ( .A(a[59]), .B(b[41]), .Z(n7397) );
  OR U7738 ( .A(n6885), .B(n6884), .Z(n6889) );
  OR U7739 ( .A(n6887), .B(n6886), .Z(n6888) );
  AND U7740 ( .A(n6889), .B(n6888), .Z(n7394) );
  OR U7741 ( .A(n6891), .B(n6890), .Z(n6895) );
  NANDN U7742 ( .A(n6893), .B(n6892), .Z(n6894) );
  AND U7743 ( .A(n6895), .B(n6894), .Z(n7520) );
  ANDN U7744 ( .B(b[44]), .A(n204), .Z(n7406) );
  OR U7745 ( .A(n6897), .B(n6896), .Z(n6901) );
  OR U7746 ( .A(n6899), .B(n6898), .Z(n6900) );
  AND U7747 ( .A(n6901), .B(n6900), .Z(n7407) );
  XNOR U7748 ( .A(n7406), .B(n7407), .Z(n7409) );
  NAND U7749 ( .A(a[54]), .B(b[46]), .Z(n7515) );
  OR U7750 ( .A(n6903), .B(n6902), .Z(n6907) );
  NANDN U7751 ( .A(n6905), .B(n6904), .Z(n6906) );
  NAND U7752 ( .A(n6907), .B(n6906), .Z(n7514) );
  XNOR U7753 ( .A(n7515), .B(n7514), .Z(n7517) );
  NAND U7754 ( .A(a[53]), .B(b[47]), .Z(n7421) );
  NANDN U7755 ( .A(n6909), .B(n6908), .Z(n6913) );
  OR U7756 ( .A(n6911), .B(n6910), .Z(n6912) );
  NAND U7757 ( .A(n6913), .B(n6912), .Z(n7419) );
  ANDN U7758 ( .B(b[48]), .A(n200), .Z(n7508) );
  OR U7759 ( .A(n6915), .B(n6914), .Z(n6919) );
  OR U7760 ( .A(n6917), .B(n6916), .Z(n6918) );
  AND U7761 ( .A(n6919), .B(n6918), .Z(n7509) );
  XNOR U7762 ( .A(n7508), .B(n7509), .Z(n7511) );
  NAND U7763 ( .A(b[51]), .B(a[49]), .Z(n7504) );
  NANDN U7764 ( .A(n6921), .B(n6920), .Z(n6925) );
  NANDN U7765 ( .A(n6923), .B(n6922), .Z(n6924) );
  AND U7766 ( .A(n6925), .B(n6924), .Z(n7503) );
  NAND U7767 ( .A(a[47]), .B(b[53]), .Z(n7445) );
  OR U7768 ( .A(n6927), .B(n6926), .Z(n6931) );
  OR U7769 ( .A(n6929), .B(n6928), .Z(n6930) );
  AND U7770 ( .A(n6931), .B(n6930), .Z(n7442) );
  ANDN U7771 ( .B(b[54]), .A(n194), .Z(n7448) );
  OR U7772 ( .A(n6933), .B(n6932), .Z(n6937) );
  NANDN U7773 ( .A(n6935), .B(n6934), .Z(n6936) );
  AND U7774 ( .A(n6937), .B(n6936), .Z(n7449) );
  XNOR U7775 ( .A(n7448), .B(n7449), .Z(n7451) );
  NAND U7776 ( .A(a[44]), .B(b[56]), .Z(n7455) );
  OR U7777 ( .A(n6939), .B(n6938), .Z(n6943) );
  NANDN U7778 ( .A(n6941), .B(n6940), .Z(n6942) );
  NAND U7779 ( .A(n6943), .B(n6942), .Z(n7454) );
  XNOR U7780 ( .A(n7455), .B(n7454), .Z(n7457) );
  NAND U7781 ( .A(a[43]), .B(b[57]), .Z(n7463) );
  OR U7782 ( .A(n6945), .B(n6944), .Z(n6949) );
  OR U7783 ( .A(n6947), .B(n6946), .Z(n6948) );
  AND U7784 ( .A(n6949), .B(n6948), .Z(n7460) );
  ANDN U7785 ( .B(b[58]), .A(n190), .Z(n7490) );
  OR U7786 ( .A(n6951), .B(n6950), .Z(n6955) );
  NANDN U7787 ( .A(n6953), .B(n6952), .Z(n6954) );
  AND U7788 ( .A(n6955), .B(n6954), .Z(n7491) );
  XNOR U7789 ( .A(n7490), .B(n7491), .Z(n7493) );
  NAND U7790 ( .A(b[61]), .B(a[39]), .Z(n7474) );
  OR U7791 ( .A(n6957), .B(n6956), .Z(n6961) );
  OR U7792 ( .A(n6959), .B(n6958), .Z(n6960) );
  AND U7793 ( .A(n6961), .B(n6960), .Z(n7472) );
  ANDN U7794 ( .B(b[63]), .A(n21772), .Z(n7480) );
  ANDN U7795 ( .B(a[38]), .A(n159), .Z(n7478) );
  OR U7796 ( .A(n6963), .B(n6962), .Z(n6967) );
  OR U7797 ( .A(n6965), .B(n6964), .Z(n6966) );
  AND U7798 ( .A(n6967), .B(n6966), .Z(n7479) );
  XNOR U7799 ( .A(n7478), .B(n7479), .Z(n7481) );
  XNOR U7800 ( .A(n7480), .B(n7481), .Z(n7473) );
  XNOR U7801 ( .A(n7472), .B(n7473), .Z(n7475) );
  XOR U7802 ( .A(n7474), .B(n7475), .Z(n7486) );
  NAND U7803 ( .A(a[40]), .B(b[60]), .Z(n7485) );
  OR U7804 ( .A(n6969), .B(n6968), .Z(n6973) );
  OR U7805 ( .A(n6971), .B(n6970), .Z(n6972) );
  NAND U7806 ( .A(n6973), .B(n6972), .Z(n7484) );
  XNOR U7807 ( .A(n7485), .B(n7484), .Z(n7487) );
  XNOR U7808 ( .A(n7486), .B(n7487), .Z(n7466) );
  OR U7809 ( .A(n6975), .B(n6974), .Z(n6979) );
  NANDN U7810 ( .A(n6977), .B(n6976), .Z(n6978) );
  NAND U7811 ( .A(n6979), .B(n6978), .Z(n7467) );
  XNOR U7812 ( .A(n7466), .B(n7467), .Z(n7469) );
  ANDN U7813 ( .B(b[59]), .A(n189), .Z(n7468) );
  XNOR U7814 ( .A(n7469), .B(n7468), .Z(n7492) );
  XOR U7815 ( .A(n7493), .B(n7492), .Z(n7461) );
  XNOR U7816 ( .A(n7460), .B(n7461), .Z(n7462) );
  XOR U7817 ( .A(n7463), .B(n7462), .Z(n7456) );
  OR U7818 ( .A(n6981), .B(n6980), .Z(n6985) );
  OR U7819 ( .A(n6983), .B(n6982), .Z(n6984) );
  NAND U7820 ( .A(n6985), .B(n6984), .Z(n7497) );
  XOR U7821 ( .A(n7496), .B(n7497), .Z(n7498) );
  ANDN U7822 ( .B(b[55]), .A(n193), .Z(n7499) );
  XOR U7823 ( .A(n7498), .B(n7499), .Z(n7450) );
  XOR U7824 ( .A(n7451), .B(n7450), .Z(n7443) );
  XNOR U7825 ( .A(n7442), .B(n7443), .Z(n7444) );
  XOR U7826 ( .A(n7445), .B(n7444), .Z(n7438) );
  ANDN U7827 ( .B(b[52]), .A(n196), .Z(n7436) );
  OR U7828 ( .A(n6987), .B(n6986), .Z(n6991) );
  OR U7829 ( .A(n6989), .B(n6988), .Z(n6990) );
  AND U7830 ( .A(n6991), .B(n6990), .Z(n7437) );
  XNOR U7831 ( .A(n7436), .B(n7437), .Z(n7439) );
  XOR U7832 ( .A(n7438), .B(n7439), .Z(n7502) );
  NAND U7833 ( .A(a[50]), .B(b[50]), .Z(n7431) );
  OR U7834 ( .A(n6993), .B(n6992), .Z(n6997) );
  OR U7835 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U7836 ( .A(n6997), .B(n6996), .Z(n7430) );
  XNOR U7837 ( .A(n7431), .B(n7430), .Z(n7433) );
  XNOR U7838 ( .A(n7432), .B(n7433), .Z(n7424) );
  OR U7839 ( .A(n6999), .B(n6998), .Z(n7003) );
  NANDN U7840 ( .A(n7001), .B(n7000), .Z(n7002) );
  NAND U7841 ( .A(n7003), .B(n7002), .Z(n7425) );
  XNOR U7842 ( .A(n7424), .B(n7425), .Z(n7427) );
  ANDN U7843 ( .B(b[49]), .A(n199), .Z(n7426) );
  XNOR U7844 ( .A(n7427), .B(n7426), .Z(n7510) );
  XOR U7845 ( .A(n7511), .B(n7510), .Z(n7418) );
  XOR U7846 ( .A(n7419), .B(n7418), .Z(n7420) );
  NANDN U7847 ( .A(n7005), .B(n7004), .Z(n7009) );
  NANDN U7848 ( .A(n7007), .B(n7006), .Z(n7008) );
  AND U7849 ( .A(n7009), .B(n7008), .Z(n7413) );
  XOR U7850 ( .A(n7412), .B(n7413), .Z(n7414) );
  ANDN U7851 ( .B(b[45]), .A(n203), .Z(n7415) );
  XOR U7852 ( .A(n7414), .B(n7415), .Z(n7408) );
  XOR U7853 ( .A(n7409), .B(n7408), .Z(n7521) );
  XNOR U7854 ( .A(n7520), .B(n7521), .Z(n7523) );
  NAND U7855 ( .A(a[57]), .B(b[43]), .Z(n7522) );
  XOR U7856 ( .A(n7523), .B(n7522), .Z(n7403) );
  ANDN U7857 ( .B(b[42]), .A(n206), .Z(n7400) );
  OR U7858 ( .A(n7011), .B(n7010), .Z(n7015) );
  NANDN U7859 ( .A(n7013), .B(n7012), .Z(n7014) );
  AND U7860 ( .A(n7015), .B(n7014), .Z(n7401) );
  XOR U7861 ( .A(n7400), .B(n7401), .Z(n7402) );
  XNOR U7862 ( .A(n7403), .B(n7402), .Z(n7395) );
  XNOR U7863 ( .A(n7394), .B(n7395), .Z(n7396) );
  XOR U7864 ( .A(n7397), .B(n7396), .Z(n7391) );
  ANDN U7865 ( .B(b[40]), .A(n208), .Z(n7388) );
  OR U7866 ( .A(n7017), .B(n7016), .Z(n7021) );
  OR U7867 ( .A(n7019), .B(n7018), .Z(n7020) );
  AND U7868 ( .A(n7021), .B(n7020), .Z(n7389) );
  XOR U7869 ( .A(n7388), .B(n7389), .Z(n7390) );
  XNOR U7870 ( .A(n7391), .B(n7390), .Z(n7526) );
  XNOR U7871 ( .A(n7527), .B(n7526), .Z(n7529) );
  NAND U7872 ( .A(a[61]), .B(b[39]), .Z(n7528) );
  XOR U7873 ( .A(n7529), .B(n7528), .Z(n7384) );
  XOR U7874 ( .A(n7023), .B(n7022), .Z(n7380) );
  XOR U7875 ( .A(n7025), .B(n7024), .Z(n7377) );
  XNOR U7876 ( .A(n7027), .B(n7026), .Z(n7373) );
  XOR U7877 ( .A(n7029), .B(n7028), .Z(n7369) );
  XOR U7878 ( .A(n7031), .B(n7030), .Z(n7365) );
  XOR U7879 ( .A(n7033), .B(n7032), .Z(n7361) );
  XOR U7880 ( .A(n7035), .B(n7034), .Z(n7357) );
  XOR U7881 ( .A(n7037), .B(n7036), .Z(n7353) );
  XNOR U7882 ( .A(n7039), .B(n7038), .Z(n7349) );
  XNOR U7883 ( .A(n7041), .B(n7040), .Z(n7345) );
  XOR U7884 ( .A(n7043), .B(n7042), .Z(n7341) );
  XOR U7885 ( .A(n7045), .B(n7044), .Z(n7337) );
  XOR U7886 ( .A(n7047), .B(n7046), .Z(n7333) );
  XNOR U7887 ( .A(n7049), .B(n7048), .Z(n7328) );
  XNOR U7888 ( .A(n7051), .B(n7050), .Z(n7325) );
  XOR U7889 ( .A(n7053), .B(n7052), .Z(n7321) );
  XOR U7890 ( .A(n7055), .B(n7054), .Z(n7317) );
  XNOR U7891 ( .A(n7057), .B(n7056), .Z(n7313) );
  XNOR U7892 ( .A(n7059), .B(n7058), .Z(n7309) );
  XNOR U7893 ( .A(n7061), .B(n7060), .Z(n7305) );
  XNOR U7894 ( .A(n7063), .B(n7062), .Z(n7301) );
  XNOR U7895 ( .A(n7065), .B(n7064), .Z(n7297) );
  XNOR U7896 ( .A(n7067), .B(n7066), .Z(n7293) );
  XOR U7897 ( .A(n7069), .B(n7068), .Z(n7289) );
  XOR U7898 ( .A(n7071), .B(n7070), .Z(n7285) );
  XOR U7899 ( .A(n7073), .B(n7072), .Z(n7281) );
  XOR U7900 ( .A(n7075), .B(n7074), .Z(n7277) );
  XNOR U7901 ( .A(n7077), .B(n7076), .Z(n7273) );
  XOR U7902 ( .A(n7079), .B(n7078), .Z(n7269) );
  XOR U7903 ( .A(n7081), .B(n7080), .Z(n7265) );
  XNOR U7904 ( .A(n7083), .B(n7082), .Z(n7261) );
  XOR U7905 ( .A(n7085), .B(n7084), .Z(n7257) );
  XNOR U7906 ( .A(n7087), .B(n7086), .Z(n7253) );
  XNOR U7907 ( .A(n7089), .B(n7088), .Z(n7249) );
  XOR U7908 ( .A(n7091), .B(n7090), .Z(n7245) );
  XOR U7909 ( .A(n7093), .B(n7092), .Z(n7240) );
  XOR U7910 ( .A(n7095), .B(n7094), .Z(n7236) );
  XNOR U7911 ( .A(n7097), .B(n7096), .Z(n7232) );
  XNOR U7912 ( .A(n7099), .B(n7098), .Z(n7228) );
  XNOR U7913 ( .A(n7101), .B(n7100), .Z(n7224) );
  XOR U7914 ( .A(n7103), .B(n7102), .Z(n7220) );
  XNOR U7915 ( .A(n7105), .B(n7104), .Z(n7216) );
  XOR U7916 ( .A(n7107), .B(n7106), .Z(n7212) );
  XNOR U7917 ( .A(n7109), .B(n7108), .Z(n7208) );
  XNOR U7918 ( .A(n7111), .B(n7110), .Z(n7204) );
  XOR U7919 ( .A(n7113), .B(n7112), .Z(n7200) );
  XOR U7920 ( .A(n7115), .B(n7114), .Z(n7196) );
  XNOR U7921 ( .A(n7117), .B(n7116), .Z(n7192) );
  XNOR U7922 ( .A(n7119), .B(n7118), .Z(n7188) );
  XNOR U7923 ( .A(n7121), .B(n7120), .Z(n7184) );
  XNOR U7924 ( .A(n7123), .B(n7122), .Z(n7180) );
  XOR U7925 ( .A(n7125), .B(n7124), .Z(n7176) );
  XOR U7926 ( .A(n7127), .B(n7126), .Z(n7172) );
  XNOR U7927 ( .A(n7129), .B(n7128), .Z(n7168) );
  XOR U7928 ( .A(n7131), .B(n7130), .Z(n7164) );
  XNOR U7929 ( .A(n7133), .B(n7132), .Z(n7160) );
  XNOR U7930 ( .A(n7135), .B(n7134), .Z(n7156) );
  XNOR U7931 ( .A(n7137), .B(n7136), .Z(n7152) );
  XNOR U7932 ( .A(n7139), .B(n7138), .Z(n7148) );
  NAND U7933 ( .A(b[39]), .B(a[1]), .Z(n7141) );
  NAND U7934 ( .A(n7141), .B(n7140), .Z(n7144) );
  AND U7935 ( .A(b[38]), .B(a[0]), .Z(n7912) );
  NANDN U7936 ( .A(n7141), .B(n7912), .Z(n7539) );
  NANDN U7937 ( .A(n7143), .B(n7539), .Z(n7142) );
  AND U7938 ( .A(n7144), .B(n7142), .Z(n7147) );
  XNOR U7939 ( .A(n7539), .B(n7143), .Z(n7145) );
  NAND U7940 ( .A(n7145), .B(n7144), .Z(n7547) );
  AND U7941 ( .A(b[38]), .B(a[2]), .Z(n7548) );
  OR U7942 ( .A(n7547), .B(n7548), .Z(n7146) );
  AND U7943 ( .A(n7147), .B(n7146), .Z(n7149) );
  OR U7944 ( .A(n7148), .B(n7149), .Z(n7151) );
  XNOR U7945 ( .A(n7149), .B(n7148), .Z(n7534) );
  AND U7946 ( .A(b[38]), .B(a[3]), .Z(n7535) );
  OR U7947 ( .A(n7534), .B(n7535), .Z(n7150) );
  AND U7948 ( .A(n7151), .B(n7150), .Z(n7153) );
  OR U7949 ( .A(n7152), .B(n7153), .Z(n7155) );
  XNOR U7950 ( .A(n7153), .B(n7152), .Z(n7557) );
  AND U7951 ( .A(b[38]), .B(a[4]), .Z(n7558) );
  OR U7952 ( .A(n7557), .B(n7558), .Z(n7154) );
  AND U7953 ( .A(n7155), .B(n7154), .Z(n7157) );
  OR U7954 ( .A(n7156), .B(n7157), .Z(n7159) );
  XNOR U7955 ( .A(n7157), .B(n7156), .Z(n7561) );
  NAND U7956 ( .A(a[5]), .B(b[38]), .Z(n7562) );
  NANDN U7957 ( .A(n7561), .B(n7562), .Z(n7158) );
  AND U7958 ( .A(n7159), .B(n7158), .Z(n7161) );
  OR U7959 ( .A(n7160), .B(n7161), .Z(n7163) );
  XNOR U7960 ( .A(n7161), .B(n7160), .Z(n7569) );
  AND U7961 ( .A(b[38]), .B(a[6]), .Z(n7570) );
  OR U7962 ( .A(n7569), .B(n7570), .Z(n7162) );
  AND U7963 ( .A(n7163), .B(n7162), .Z(n7165) );
  OR U7964 ( .A(n7164), .B(n7165), .Z(n7167) );
  XNOR U7965 ( .A(n7165), .B(n7164), .Z(n7575) );
  NAND U7966 ( .A(a[7]), .B(b[38]), .Z(n7576) );
  NANDN U7967 ( .A(n7575), .B(n7576), .Z(n7166) );
  AND U7968 ( .A(n7167), .B(n7166), .Z(n7169) );
  OR U7969 ( .A(n7168), .B(n7169), .Z(n7171) );
  XNOR U7970 ( .A(n7169), .B(n7168), .Z(n7581) );
  AND U7971 ( .A(b[38]), .B(a[8]), .Z(n7582) );
  OR U7972 ( .A(n7581), .B(n7582), .Z(n7170) );
  AND U7973 ( .A(n7171), .B(n7170), .Z(n7173) );
  OR U7974 ( .A(n7172), .B(n7173), .Z(n7175) );
  XNOR U7975 ( .A(n7173), .B(n7172), .Z(n7585) );
  NAND U7976 ( .A(a[9]), .B(b[38]), .Z(n7586) );
  NANDN U7977 ( .A(n7585), .B(n7586), .Z(n7174) );
  AND U7978 ( .A(n7175), .B(n7174), .Z(n7177) );
  OR U7979 ( .A(n7176), .B(n7177), .Z(n7179) );
  XNOR U7980 ( .A(n7177), .B(n7176), .Z(n7593) );
  AND U7981 ( .A(b[38]), .B(a[10]), .Z(n7594) );
  OR U7982 ( .A(n7593), .B(n7594), .Z(n7178) );
  AND U7983 ( .A(n7179), .B(n7178), .Z(n7181) );
  OR U7984 ( .A(n7180), .B(n7181), .Z(n7183) );
  XNOR U7985 ( .A(n7181), .B(n7180), .Z(n7599) );
  NAND U7986 ( .A(a[11]), .B(b[38]), .Z(n7600) );
  NANDN U7987 ( .A(n7599), .B(n7600), .Z(n7182) );
  AND U7988 ( .A(n7183), .B(n7182), .Z(n7185) );
  OR U7989 ( .A(n7184), .B(n7185), .Z(n7187) );
  XNOR U7990 ( .A(n7185), .B(n7184), .Z(n7605) );
  AND U7991 ( .A(b[38]), .B(a[12]), .Z(n7606) );
  OR U7992 ( .A(n7605), .B(n7606), .Z(n7186) );
  AND U7993 ( .A(n7187), .B(n7186), .Z(n7189) );
  OR U7994 ( .A(n7188), .B(n7189), .Z(n7191) );
  XNOR U7995 ( .A(n7189), .B(n7188), .Z(n7609) );
  NAND U7996 ( .A(a[13]), .B(b[38]), .Z(n7610) );
  NANDN U7997 ( .A(n7609), .B(n7610), .Z(n7190) );
  AND U7998 ( .A(n7191), .B(n7190), .Z(n7193) );
  OR U7999 ( .A(n7192), .B(n7193), .Z(n7195) );
  XNOR U8000 ( .A(n7193), .B(n7192), .Z(n7617) );
  AND U8001 ( .A(b[38]), .B(a[14]), .Z(n7618) );
  OR U8002 ( .A(n7617), .B(n7618), .Z(n7194) );
  AND U8003 ( .A(n7195), .B(n7194), .Z(n7197) );
  OR U8004 ( .A(n7196), .B(n7197), .Z(n7199) );
  XNOR U8005 ( .A(n7197), .B(n7196), .Z(n7621) );
  NAND U8006 ( .A(a[15]), .B(b[38]), .Z(n7622) );
  NANDN U8007 ( .A(n7621), .B(n7622), .Z(n7198) );
  AND U8008 ( .A(n7199), .B(n7198), .Z(n7201) );
  OR U8009 ( .A(n7200), .B(n7201), .Z(n7203) );
  XNOR U8010 ( .A(n7201), .B(n7200), .Z(n7629) );
  AND U8011 ( .A(b[38]), .B(a[16]), .Z(n7630) );
  OR U8012 ( .A(n7629), .B(n7630), .Z(n7202) );
  AND U8013 ( .A(n7203), .B(n7202), .Z(n7205) );
  OR U8014 ( .A(n7204), .B(n7205), .Z(n7207) );
  XNOR U8015 ( .A(n7205), .B(n7204), .Z(n7633) );
  NAND U8016 ( .A(a[17]), .B(b[38]), .Z(n7634) );
  NANDN U8017 ( .A(n7633), .B(n7634), .Z(n7206) );
  AND U8018 ( .A(n7207), .B(n7206), .Z(n7209) );
  OR U8019 ( .A(n7208), .B(n7209), .Z(n7211) );
  XNOR U8020 ( .A(n7209), .B(n7208), .Z(n7641) );
  AND U8021 ( .A(b[38]), .B(a[18]), .Z(n7642) );
  OR U8022 ( .A(n7641), .B(n7642), .Z(n7210) );
  AND U8023 ( .A(n7211), .B(n7210), .Z(n7213) );
  OR U8024 ( .A(n7212), .B(n7213), .Z(n7215) );
  XNOR U8025 ( .A(n7213), .B(n7212), .Z(n7645) );
  NAND U8026 ( .A(a[19]), .B(b[38]), .Z(n7646) );
  NANDN U8027 ( .A(n7645), .B(n7646), .Z(n7214) );
  AND U8028 ( .A(n7215), .B(n7214), .Z(n7217) );
  OR U8029 ( .A(n7216), .B(n7217), .Z(n7219) );
  XNOR U8030 ( .A(n7217), .B(n7216), .Z(n7653) );
  NAND U8031 ( .A(a[20]), .B(b[38]), .Z(n7654) );
  NANDN U8032 ( .A(n7653), .B(n7654), .Z(n7218) );
  AND U8033 ( .A(n7219), .B(n7218), .Z(n7221) );
  OR U8034 ( .A(n7220), .B(n7221), .Z(n7223) );
  XNOR U8035 ( .A(n7221), .B(n7220), .Z(n7657) );
  NAND U8036 ( .A(a[21]), .B(b[38]), .Z(n7658) );
  NANDN U8037 ( .A(n7657), .B(n7658), .Z(n7222) );
  AND U8038 ( .A(n7223), .B(n7222), .Z(n7225) );
  OR U8039 ( .A(n7224), .B(n7225), .Z(n7227) );
  XNOR U8040 ( .A(n7225), .B(n7224), .Z(n7665) );
  AND U8041 ( .A(b[38]), .B(a[22]), .Z(n7666) );
  OR U8042 ( .A(n7665), .B(n7666), .Z(n7226) );
  AND U8043 ( .A(n7227), .B(n7226), .Z(n7229) );
  OR U8044 ( .A(n7228), .B(n7229), .Z(n7231) );
  XNOR U8045 ( .A(n7229), .B(n7228), .Z(n7669) );
  NAND U8046 ( .A(a[23]), .B(b[38]), .Z(n7670) );
  NANDN U8047 ( .A(n7669), .B(n7670), .Z(n7230) );
  AND U8048 ( .A(n7231), .B(n7230), .Z(n7233) );
  OR U8049 ( .A(n7232), .B(n7233), .Z(n7235) );
  XNOR U8050 ( .A(n7233), .B(n7232), .Z(n7677) );
  AND U8051 ( .A(b[38]), .B(a[24]), .Z(n7678) );
  OR U8052 ( .A(n7677), .B(n7678), .Z(n7234) );
  AND U8053 ( .A(n7235), .B(n7234), .Z(n7237) );
  OR U8054 ( .A(n7236), .B(n7237), .Z(n7239) );
  XNOR U8055 ( .A(n7237), .B(n7236), .Z(n7681) );
  NAND U8056 ( .A(a[25]), .B(b[38]), .Z(n7682) );
  NANDN U8057 ( .A(n7681), .B(n7682), .Z(n7238) );
  AND U8058 ( .A(n7239), .B(n7238), .Z(n7241) );
  OR U8059 ( .A(n7240), .B(n7241), .Z(n7243) );
  XNOR U8060 ( .A(n7241), .B(n7240), .Z(n7689) );
  AND U8061 ( .A(b[38]), .B(a[26]), .Z(n7690) );
  OR U8062 ( .A(n7689), .B(n7690), .Z(n7242) );
  NAND U8063 ( .A(n7243), .B(n7242), .Z(n7244) );
  NANDN U8064 ( .A(n7245), .B(n7244), .Z(n7247) );
  AND U8065 ( .A(b[38]), .B(a[27]), .Z(n7696) );
  NANDN U8066 ( .A(n7696), .B(n7695), .Z(n7246) );
  NAND U8067 ( .A(n7247), .B(n7246), .Z(n7248) );
  NANDN U8068 ( .A(n7249), .B(n7248), .Z(n7251) );
  AND U8069 ( .A(b[38]), .B(a[28]), .Z(n7702) );
  NANDN U8070 ( .A(n7702), .B(n7701), .Z(n7250) );
  NAND U8071 ( .A(n7251), .B(n7250), .Z(n7252) );
  NANDN U8072 ( .A(n7253), .B(n7252), .Z(n7255) );
  AND U8073 ( .A(b[38]), .B(a[29]), .Z(n7706) );
  NANDN U8074 ( .A(n7706), .B(n7705), .Z(n7254) );
  NAND U8075 ( .A(n7255), .B(n7254), .Z(n7256) );
  NANDN U8076 ( .A(n7257), .B(n7256), .Z(n7259) );
  AND U8077 ( .A(b[38]), .B(a[30]), .Z(n7714) );
  NANDN U8078 ( .A(n7714), .B(n7713), .Z(n7258) );
  NAND U8079 ( .A(n7259), .B(n7258), .Z(n7260) );
  NANDN U8080 ( .A(n7261), .B(n7260), .Z(n7263) );
  AND U8081 ( .A(b[38]), .B(a[31]), .Z(n7718) );
  NANDN U8082 ( .A(n7718), .B(n7717), .Z(n7262) );
  NAND U8083 ( .A(n7263), .B(n7262), .Z(n7264) );
  NANDN U8084 ( .A(n7265), .B(n7264), .Z(n7267) );
  AND U8085 ( .A(b[38]), .B(a[32]), .Z(n7726) );
  NANDN U8086 ( .A(n7726), .B(n7725), .Z(n7266) );
  NAND U8087 ( .A(n7267), .B(n7266), .Z(n7268) );
  NANDN U8088 ( .A(n7269), .B(n7268), .Z(n7271) );
  AND U8089 ( .A(b[38]), .B(a[33]), .Z(n7730) );
  NANDN U8090 ( .A(n7730), .B(n7729), .Z(n7270) );
  NAND U8091 ( .A(n7271), .B(n7270), .Z(n7272) );
  NANDN U8092 ( .A(n7273), .B(n7272), .Z(n7275) );
  AND U8093 ( .A(b[38]), .B(a[34]), .Z(n7738) );
  NANDN U8094 ( .A(n7738), .B(n7737), .Z(n7274) );
  NAND U8095 ( .A(n7275), .B(n7274), .Z(n7276) );
  NANDN U8096 ( .A(n7277), .B(n7276), .Z(n7279) );
  AND U8097 ( .A(b[38]), .B(a[35]), .Z(n7742) );
  NANDN U8098 ( .A(n7742), .B(n7741), .Z(n7278) );
  NAND U8099 ( .A(n7279), .B(n7278), .Z(n7280) );
  NANDN U8100 ( .A(n7281), .B(n7280), .Z(n7283) );
  AND U8101 ( .A(b[38]), .B(a[36]), .Z(n7750) );
  NANDN U8102 ( .A(n7750), .B(n7749), .Z(n7282) );
  NAND U8103 ( .A(n7283), .B(n7282), .Z(n7284) );
  NANDN U8104 ( .A(n7285), .B(n7284), .Z(n7287) );
  AND U8105 ( .A(b[38]), .B(a[37]), .Z(n7754) );
  NANDN U8106 ( .A(n7754), .B(n7753), .Z(n7286) );
  NAND U8107 ( .A(n7287), .B(n7286), .Z(n7288) );
  NANDN U8108 ( .A(n7289), .B(n7288), .Z(n7291) );
  AND U8109 ( .A(b[38]), .B(a[38]), .Z(n7762) );
  NANDN U8110 ( .A(n7762), .B(n7761), .Z(n7290) );
  NAND U8111 ( .A(n7291), .B(n7290), .Z(n7292) );
  NANDN U8112 ( .A(n7293), .B(n7292), .Z(n7295) );
  AND U8113 ( .A(b[38]), .B(a[39]), .Z(n7766) );
  NANDN U8114 ( .A(n7766), .B(n7765), .Z(n7294) );
  NAND U8115 ( .A(n7295), .B(n7294), .Z(n7296) );
  NANDN U8116 ( .A(n7297), .B(n7296), .Z(n7299) );
  AND U8117 ( .A(b[38]), .B(a[40]), .Z(n7774) );
  NANDN U8118 ( .A(n7774), .B(n7773), .Z(n7298) );
  NAND U8119 ( .A(n7299), .B(n7298), .Z(n7300) );
  NANDN U8120 ( .A(n7301), .B(n7300), .Z(n7303) );
  AND U8121 ( .A(b[38]), .B(a[41]), .Z(n7778) );
  NANDN U8122 ( .A(n7778), .B(n7777), .Z(n7302) );
  NAND U8123 ( .A(n7303), .B(n7302), .Z(n7304) );
  NANDN U8124 ( .A(n7305), .B(n7304), .Z(n7307) );
  AND U8125 ( .A(b[38]), .B(a[42]), .Z(n7786) );
  NANDN U8126 ( .A(n7786), .B(n7785), .Z(n7306) );
  NAND U8127 ( .A(n7307), .B(n7306), .Z(n7308) );
  NANDN U8128 ( .A(n7309), .B(n7308), .Z(n7311) );
  AND U8129 ( .A(b[38]), .B(a[43]), .Z(n7790) );
  NANDN U8130 ( .A(n7790), .B(n7789), .Z(n7310) );
  NAND U8131 ( .A(n7311), .B(n7310), .Z(n7312) );
  NANDN U8132 ( .A(n7313), .B(n7312), .Z(n7315) );
  AND U8133 ( .A(b[38]), .B(a[44]), .Z(n7798) );
  NANDN U8134 ( .A(n7798), .B(n7797), .Z(n7314) );
  NAND U8135 ( .A(n7315), .B(n7314), .Z(n7316) );
  NANDN U8136 ( .A(n7317), .B(n7316), .Z(n7319) );
  AND U8137 ( .A(b[38]), .B(a[45]), .Z(n7802) );
  OR U8138 ( .A(n7802), .B(n7801), .Z(n7318) );
  NAND U8139 ( .A(n7319), .B(n7318), .Z(n7320) );
  NANDN U8140 ( .A(n7321), .B(n7320), .Z(n7323) );
  AND U8141 ( .A(b[38]), .B(a[46]), .Z(n7810) );
  NANDN U8142 ( .A(n7810), .B(n7809), .Z(n7322) );
  NAND U8143 ( .A(n7323), .B(n7322), .Z(n7324) );
  NANDN U8144 ( .A(n7325), .B(n7324), .Z(n7327) );
  AND U8145 ( .A(b[38]), .B(a[47]), .Z(n7814) );
  NANDN U8146 ( .A(n7814), .B(n7813), .Z(n7326) );
  NAND U8147 ( .A(n7327), .B(n7326), .Z(n7329) );
  NANDN U8148 ( .A(n7328), .B(n7329), .Z(n7331) );
  AND U8149 ( .A(b[38]), .B(a[48]), .Z(n7822) );
  XOR U8150 ( .A(n7329), .B(n7328), .Z(n7821) );
  OR U8151 ( .A(n7822), .B(n7821), .Z(n7330) );
  NAND U8152 ( .A(n7331), .B(n7330), .Z(n7332) );
  NANDN U8153 ( .A(n7333), .B(n7332), .Z(n7335) );
  AND U8154 ( .A(b[38]), .B(a[49]), .Z(n7826) );
  NANDN U8155 ( .A(n7826), .B(n7825), .Z(n7334) );
  NAND U8156 ( .A(n7335), .B(n7334), .Z(n7336) );
  NANDN U8157 ( .A(n7337), .B(n7336), .Z(n7339) );
  AND U8158 ( .A(b[38]), .B(a[50]), .Z(n7834) );
  NANDN U8159 ( .A(n7834), .B(n7833), .Z(n7338) );
  NAND U8160 ( .A(n7339), .B(n7338), .Z(n7340) );
  NANDN U8161 ( .A(n7341), .B(n7340), .Z(n7343) );
  AND U8162 ( .A(b[38]), .B(a[51]), .Z(n7838) );
  NANDN U8163 ( .A(n7838), .B(n7837), .Z(n7342) );
  NAND U8164 ( .A(n7343), .B(n7342), .Z(n7344) );
  NANDN U8165 ( .A(n7345), .B(n7344), .Z(n7347) );
  AND U8166 ( .A(b[38]), .B(a[52]), .Z(n7846) );
  NANDN U8167 ( .A(n7846), .B(n7845), .Z(n7346) );
  NAND U8168 ( .A(n7347), .B(n7346), .Z(n7348) );
  NANDN U8169 ( .A(n7349), .B(n7348), .Z(n7351) );
  AND U8170 ( .A(b[38]), .B(a[53]), .Z(n7850) );
  NANDN U8171 ( .A(n7850), .B(n7849), .Z(n7350) );
  NAND U8172 ( .A(n7351), .B(n7350), .Z(n7352) );
  NANDN U8173 ( .A(n7353), .B(n7352), .Z(n7355) );
  AND U8174 ( .A(b[38]), .B(a[54]), .Z(n7858) );
  NANDN U8175 ( .A(n7858), .B(n7857), .Z(n7354) );
  NAND U8176 ( .A(n7355), .B(n7354), .Z(n7356) );
  NANDN U8177 ( .A(n7357), .B(n7356), .Z(n7359) );
  AND U8178 ( .A(b[38]), .B(a[55]), .Z(n7862) );
  NANDN U8179 ( .A(n7862), .B(n7861), .Z(n7358) );
  NAND U8180 ( .A(n7359), .B(n7358), .Z(n7360) );
  NANDN U8181 ( .A(n7361), .B(n7360), .Z(n7363) );
  AND U8182 ( .A(b[38]), .B(a[56]), .Z(n7870) );
  NANDN U8183 ( .A(n7870), .B(n7869), .Z(n7362) );
  NAND U8184 ( .A(n7363), .B(n7362), .Z(n7364) );
  NANDN U8185 ( .A(n7365), .B(n7364), .Z(n7367) );
  AND U8186 ( .A(b[38]), .B(a[57]), .Z(n7874) );
  NANDN U8187 ( .A(n7874), .B(n7873), .Z(n7366) );
  NAND U8188 ( .A(n7367), .B(n7366), .Z(n7368) );
  NANDN U8189 ( .A(n7369), .B(n7368), .Z(n7371) );
  AND U8190 ( .A(b[38]), .B(a[58]), .Z(n7882) );
  NANDN U8191 ( .A(n7882), .B(n7881), .Z(n7370) );
  NAND U8192 ( .A(n7371), .B(n7370), .Z(n7372) );
  NANDN U8193 ( .A(n7373), .B(n7372), .Z(n7375) );
  AND U8194 ( .A(b[38]), .B(a[59]), .Z(n7886) );
  OR U8195 ( .A(n7886), .B(n7885), .Z(n7374) );
  NAND U8196 ( .A(n7375), .B(n7374), .Z(n7376) );
  NANDN U8197 ( .A(n7377), .B(n7376), .Z(n7379) );
  AND U8198 ( .A(b[38]), .B(a[60]), .Z(n7894) );
  NANDN U8199 ( .A(n7894), .B(n7893), .Z(n7378) );
  AND U8200 ( .A(n7379), .B(n7378), .Z(n7381) );
  OR U8201 ( .A(n7380), .B(n7381), .Z(n7383) );
  XNOR U8202 ( .A(n7381), .B(n7380), .Z(n7899) );
  NAND U8203 ( .A(a[61]), .B(b[38]), .Z(n7900) );
  NANDN U8204 ( .A(n7899), .B(n7900), .Z(n7382) );
  AND U8205 ( .A(n7383), .B(n7382), .Z(n7385) );
  OR U8206 ( .A(n7384), .B(n7385), .Z(n7387) );
  XNOR U8207 ( .A(n7385), .B(n7384), .Z(n7532) );
  AND U8208 ( .A(b[38]), .B(a[62]), .Z(n7533) );
  OR U8209 ( .A(n7532), .B(n7533), .Z(n7386) );
  AND U8210 ( .A(n7387), .B(n7386), .Z(n22151) );
  AND U8211 ( .A(b[38]), .B(a[63]), .Z(n22152) );
  XNOR U8212 ( .A(n22151), .B(n22152), .Z(n22154) );
  NAND U8213 ( .A(a[61]), .B(b[40]), .Z(n22140) );
  OR U8214 ( .A(n7389), .B(n7388), .Z(n7393) );
  NANDN U8215 ( .A(n7391), .B(n7390), .Z(n7392) );
  NAND U8216 ( .A(n7393), .B(n7392), .Z(n22139) );
  XNOR U8217 ( .A(n22140), .B(n22139), .Z(n22142) );
  OR U8218 ( .A(n7395), .B(n7394), .Z(n7399) );
  OR U8219 ( .A(n7397), .B(n7396), .Z(n7398) );
  AND U8220 ( .A(n7399), .B(n7398), .Z(n22133) );
  ANDN U8221 ( .B(b[42]), .A(n207), .Z(n22127) );
  OR U8222 ( .A(n7401), .B(n7400), .Z(n7405) );
  NANDN U8223 ( .A(n7403), .B(n7402), .Z(n7404) );
  AND U8224 ( .A(n7405), .B(n7404), .Z(n22128) );
  XNOR U8225 ( .A(n22127), .B(n22128), .Z(n22130) );
  NAND U8226 ( .A(a[57]), .B(b[44]), .Z(n22122) );
  OR U8227 ( .A(n7407), .B(n7406), .Z(n7411) );
  OR U8228 ( .A(n7409), .B(n7408), .Z(n7410) );
  NAND U8229 ( .A(n7411), .B(n7410), .Z(n22121) );
  XNOR U8230 ( .A(n22122), .B(n22121), .Z(n22124) );
  OR U8231 ( .A(n7413), .B(n7412), .Z(n7417) );
  NANDN U8232 ( .A(n7415), .B(n7414), .Z(n7416) );
  NAND U8233 ( .A(n7417), .B(n7416), .Z(n22014) );
  ANDN U8234 ( .B(b[47]), .A(n202), .Z(n22112) );
  OR U8235 ( .A(n7419), .B(n7418), .Z(n7423) );
  NANDN U8236 ( .A(n7421), .B(n7420), .Z(n7422) );
  NAND U8237 ( .A(n7423), .B(n7422), .Z(n22110) );
  OR U8238 ( .A(n7425), .B(n7424), .Z(n7429) );
  OR U8239 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U8240 ( .A(n7429), .B(n7428), .Z(n22020) );
  ANDN U8241 ( .B(b[50]), .A(n199), .Z(n22097) );
  OR U8242 ( .A(n7431), .B(n7430), .Z(n7435) );
  NANDN U8243 ( .A(n7433), .B(n7432), .Z(n7434) );
  NAND U8244 ( .A(n7435), .B(n7434), .Z(n22098) );
  XNOR U8245 ( .A(n22097), .B(n22098), .Z(n22100) );
  NAND U8246 ( .A(a[49]), .B(b[52]), .Z(n22092) );
  OR U8247 ( .A(n7437), .B(n7436), .Z(n7441) );
  OR U8248 ( .A(n7439), .B(n7438), .Z(n7440) );
  NAND U8249 ( .A(n7441), .B(n7440), .Z(n22091) );
  XNOR U8250 ( .A(n22092), .B(n22091), .Z(n22094) );
  OR U8251 ( .A(n7443), .B(n7442), .Z(n7447) );
  OR U8252 ( .A(n7445), .B(n7444), .Z(n7446) );
  AND U8253 ( .A(n7447), .B(n7446), .Z(n22085) );
  ANDN U8254 ( .B(b[54]), .A(n195), .Z(n22079) );
  OR U8255 ( .A(n7449), .B(n7448), .Z(n7453) );
  OR U8256 ( .A(n7451), .B(n7450), .Z(n7452) );
  AND U8257 ( .A(n7453), .B(n7452), .Z(n22080) );
  XNOR U8258 ( .A(n22079), .B(n22080), .Z(n22082) );
  NAND U8259 ( .A(a[45]), .B(b[56]), .Z(n22074) );
  OR U8260 ( .A(n7455), .B(n7454), .Z(n7459) );
  NANDN U8261 ( .A(n7457), .B(n7456), .Z(n7458) );
  AND U8262 ( .A(n7459), .B(n7458), .Z(n22073) );
  XNOR U8263 ( .A(n22074), .B(n22073), .Z(n22076) );
  OR U8264 ( .A(n7461), .B(n7460), .Z(n7465) );
  OR U8265 ( .A(n7463), .B(n7462), .Z(n7464) );
  AND U8266 ( .A(n7465), .B(n7464), .Z(n22067) );
  OR U8267 ( .A(n7467), .B(n7466), .Z(n7471) );
  OR U8268 ( .A(n7469), .B(n7468), .Z(n7470) );
  NAND U8269 ( .A(n7471), .B(n7470), .Z(n22038) );
  ANDN U8270 ( .B(b[61]), .A(n188), .Z(n22051) );
  OR U8271 ( .A(n7473), .B(n7472), .Z(n7477) );
  NANDN U8272 ( .A(n7475), .B(n7474), .Z(n7476) );
  AND U8273 ( .A(n7477), .B(n7476), .Z(n22049) );
  ANDN U8274 ( .B(b[63]), .A(n186), .Z(n22045) );
  ANDN U8275 ( .B(a[39]), .A(n159), .Z(n22043) );
  OR U8276 ( .A(n7479), .B(n7478), .Z(n7483) );
  OR U8277 ( .A(n7481), .B(n7480), .Z(n7482) );
  AND U8278 ( .A(n7483), .B(n7482), .Z(n22044) );
  XNOR U8279 ( .A(n22043), .B(n22044), .Z(n22046) );
  XNOR U8280 ( .A(n22045), .B(n22046), .Z(n22050) );
  XNOR U8281 ( .A(n22049), .B(n22050), .Z(n22052) );
  XNOR U8282 ( .A(n22051), .B(n22052), .Z(n22058) );
  ANDN U8283 ( .B(b[60]), .A(n189), .Z(n22055) );
  OR U8284 ( .A(n7485), .B(n7484), .Z(n7489) );
  NANDN U8285 ( .A(n7487), .B(n7486), .Z(n7488) );
  NAND U8286 ( .A(n7489), .B(n7488), .Z(n22056) );
  XNOR U8287 ( .A(n22055), .B(n22056), .Z(n22057) );
  XOR U8288 ( .A(n22058), .B(n22057), .Z(n22037) );
  XOR U8289 ( .A(n22038), .B(n22037), .Z(n22039) );
  NAND U8290 ( .A(a[42]), .B(b[59]), .Z(n22040) );
  ANDN U8291 ( .B(b[58]), .A(n191), .Z(n22061) );
  OR U8292 ( .A(n7491), .B(n7490), .Z(n7495) );
  OR U8293 ( .A(n7493), .B(n7492), .Z(n7494) );
  AND U8294 ( .A(n7495), .B(n7494), .Z(n22062) );
  XOR U8295 ( .A(n22061), .B(n22062), .Z(n22063) );
  XNOR U8296 ( .A(n22064), .B(n22063), .Z(n22068) );
  XNOR U8297 ( .A(n22067), .B(n22068), .Z(n22070) );
  AND U8298 ( .A(a[44]), .B(b[57]), .Z(n22069) );
  XNOR U8299 ( .A(n22070), .B(n22069), .Z(n22075) );
  OR U8300 ( .A(n7497), .B(n7496), .Z(n7501) );
  NANDN U8301 ( .A(n7499), .B(n7498), .Z(n7500) );
  AND U8302 ( .A(n7501), .B(n7500), .Z(n22032) );
  XOR U8303 ( .A(n22031), .B(n22032), .Z(n22033) );
  ANDN U8304 ( .B(b[55]), .A(n194), .Z(n22034) );
  XOR U8305 ( .A(n22033), .B(n22034), .Z(n22081) );
  XOR U8306 ( .A(n22082), .B(n22081), .Z(n22086) );
  XNOR U8307 ( .A(n22085), .B(n22086), .Z(n22088) );
  AND U8308 ( .A(a[48]), .B(b[53]), .Z(n22087) );
  XNOR U8309 ( .A(n22088), .B(n22087), .Z(n22093) );
  NANDN U8310 ( .A(n7503), .B(n7502), .Z(n7507) );
  NAND U8311 ( .A(n7505), .B(n7504), .Z(n7506) );
  AND U8312 ( .A(n7507), .B(n7506), .Z(n22026) );
  XOR U8313 ( .A(n22025), .B(n22026), .Z(n22027) );
  ANDN U8314 ( .B(b[51]), .A(n198), .Z(n22028) );
  XOR U8315 ( .A(n22027), .B(n22028), .Z(n22099) );
  XOR U8316 ( .A(n22100), .B(n22099), .Z(n22019) );
  XOR U8317 ( .A(n22020), .B(n22019), .Z(n22021) );
  NAND U8318 ( .A(a[52]), .B(b[49]), .Z(n22022) );
  ANDN U8319 ( .B(b[48]), .A(n201), .Z(n22103) );
  OR U8320 ( .A(n7509), .B(n7508), .Z(n7513) );
  OR U8321 ( .A(n7511), .B(n7510), .Z(n7512) );
  AND U8322 ( .A(n7513), .B(n7512), .Z(n22104) );
  XNOR U8323 ( .A(n22103), .B(n22104), .Z(n22106) );
  XOR U8324 ( .A(n22105), .B(n22106), .Z(n22109) );
  XOR U8325 ( .A(n22112), .B(n22111), .Z(n22118) );
  ANDN U8326 ( .B(b[46]), .A(n203), .Z(n22115) );
  OR U8327 ( .A(n7515), .B(n7514), .Z(n7519) );
  NANDN U8328 ( .A(n7517), .B(n7516), .Z(n7518) );
  NAND U8329 ( .A(n7519), .B(n7518), .Z(n22116) );
  XNOR U8330 ( .A(n22115), .B(n22116), .Z(n22117) );
  XOR U8331 ( .A(n22118), .B(n22117), .Z(n22013) );
  XNOR U8332 ( .A(n22014), .B(n22013), .Z(n22016) );
  AND U8333 ( .A(a[56]), .B(b[45]), .Z(n22015) );
  XOR U8334 ( .A(n22016), .B(n22015), .Z(n22123) );
  XOR U8335 ( .A(n22124), .B(n22123), .Z(n22007) );
  OR U8336 ( .A(n7521), .B(n7520), .Z(n7525) );
  OR U8337 ( .A(n7523), .B(n7522), .Z(n7524) );
  NAND U8338 ( .A(n7525), .B(n7524), .Z(n22008) );
  XOR U8339 ( .A(n22007), .B(n22008), .Z(n22009) );
  ANDN U8340 ( .B(b[43]), .A(n206), .Z(n22010) );
  XOR U8341 ( .A(n22009), .B(n22010), .Z(n22129) );
  XOR U8342 ( .A(n22130), .B(n22129), .Z(n22134) );
  XNOR U8343 ( .A(n22133), .B(n22134), .Z(n22136) );
  AND U8344 ( .A(a[60]), .B(b[41]), .Z(n22135) );
  XNOR U8345 ( .A(n22136), .B(n22135), .Z(n22141) );
  OR U8346 ( .A(n7527), .B(n7526), .Z(n7531) );
  OR U8347 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U8348 ( .A(n7531), .B(n7530), .Z(n22146) );
  XOR U8349 ( .A(n22145), .B(n22146), .Z(n22147) );
  XOR U8350 ( .A(n22147), .B(n22148), .Z(n22153) );
  XOR U8351 ( .A(n22154), .B(n22153), .Z(n22005) );
  XNOR U8352 ( .A(n7533), .B(n7532), .Z(n7904) );
  NAND U8353 ( .A(a[62]), .B(b[37]), .Z(n7897) );
  NAND U8354 ( .A(a[61]), .B(b[37]), .Z(n7892) );
  NAND U8355 ( .A(a[60]), .B(b[37]), .Z(n7888) );
  NAND U8356 ( .A(a[59]), .B(b[37]), .Z(n7880) );
  NAND U8357 ( .A(a[58]), .B(b[37]), .Z(n7876) );
  NAND U8358 ( .A(a[57]), .B(b[37]), .Z(n7868) );
  NAND U8359 ( .A(a[56]), .B(b[37]), .Z(n7864) );
  NAND U8360 ( .A(a[55]), .B(b[37]), .Z(n7856) );
  NAND U8361 ( .A(a[54]), .B(b[37]), .Z(n7852) );
  NAND U8362 ( .A(a[53]), .B(b[37]), .Z(n7844) );
  NAND U8363 ( .A(a[52]), .B(b[37]), .Z(n7840) );
  NAND U8364 ( .A(a[51]), .B(b[37]), .Z(n7832) );
  NAND U8365 ( .A(a[50]), .B(b[37]), .Z(n7828) );
  NAND U8366 ( .A(a[49]), .B(b[37]), .Z(n7820) );
  NAND U8367 ( .A(a[48]), .B(b[37]), .Z(n7816) );
  NAND U8368 ( .A(a[47]), .B(b[37]), .Z(n7808) );
  NAND U8369 ( .A(a[46]), .B(b[37]), .Z(n7804) );
  NAND U8370 ( .A(a[45]), .B(b[37]), .Z(n7796) );
  NAND U8371 ( .A(a[44]), .B(b[37]), .Z(n7792) );
  NAND U8372 ( .A(a[43]), .B(b[37]), .Z(n7784) );
  NAND U8373 ( .A(a[42]), .B(b[37]), .Z(n7780) );
  NAND U8374 ( .A(a[41]), .B(b[37]), .Z(n7772) );
  NAND U8375 ( .A(a[40]), .B(b[37]), .Z(n7768) );
  NAND U8376 ( .A(a[39]), .B(b[37]), .Z(n7760) );
  NAND U8377 ( .A(a[38]), .B(b[37]), .Z(n7756) );
  NAND U8378 ( .A(a[37]), .B(b[37]), .Z(n7748) );
  NAND U8379 ( .A(a[36]), .B(b[37]), .Z(n7744) );
  NAND U8380 ( .A(a[35]), .B(b[37]), .Z(n7736) );
  NAND U8381 ( .A(a[34]), .B(b[37]), .Z(n7732) );
  NAND U8382 ( .A(a[33]), .B(b[37]), .Z(n7724) );
  NAND U8383 ( .A(a[32]), .B(b[37]), .Z(n7720) );
  NAND U8384 ( .A(a[31]), .B(b[37]), .Z(n7712) );
  NAND U8385 ( .A(a[30]), .B(b[37]), .Z(n7708) );
  NAND U8386 ( .A(a[29]), .B(b[37]), .Z(n7700) );
  NAND U8387 ( .A(a[21]), .B(b[37]), .Z(n7651) );
  ANDN U8388 ( .B(b[37]), .A(n164), .Z(n7555) );
  XNOR U8389 ( .A(n7535), .B(n7534), .Z(n7551) );
  ANDN U8390 ( .B(b[37]), .A(n21580), .Z(n7545) );
  NAND U8391 ( .A(a[1]), .B(b[38]), .Z(n7537) );
  NAND U8392 ( .A(n7537), .B(n7536), .Z(n7541) );
  AND U8393 ( .A(b[37]), .B(a[0]), .Z(n8290) );
  ANDN U8394 ( .B(n8290), .A(n7537), .Z(n7540) );
  OR U8395 ( .A(n7540), .B(n7539), .Z(n7538) );
  AND U8396 ( .A(n7541), .B(n7538), .Z(n7544) );
  XOR U8397 ( .A(n7540), .B(n7539), .Z(n7542) );
  NAND U8398 ( .A(n7542), .B(n7541), .Z(n7920) );
  ANDN U8399 ( .B(b[37]), .A(n162), .Z(n7921) );
  OR U8400 ( .A(n7920), .B(n7921), .Z(n7543) );
  AND U8401 ( .A(n7544), .B(n7543), .Z(n7546) );
  OR U8402 ( .A(n7545), .B(n7546), .Z(n7550) );
  XNOR U8403 ( .A(n7546), .B(n7545), .Z(n7925) );
  XNOR U8404 ( .A(n7548), .B(n7547), .Z(n7924) );
  OR U8405 ( .A(n7925), .B(n7924), .Z(n7549) );
  AND U8406 ( .A(n7550), .B(n7549), .Z(n7552) );
  OR U8407 ( .A(n7551), .B(n7552), .Z(n7554) );
  XNOR U8408 ( .A(n7552), .B(n7551), .Z(n7932) );
  ANDN U8409 ( .B(b[37]), .A(n163), .Z(n7933) );
  OR U8410 ( .A(n7932), .B(n7933), .Z(n7553) );
  AND U8411 ( .A(n7554), .B(n7553), .Z(n7556) );
  OR U8412 ( .A(n7555), .B(n7556), .Z(n7560) );
  XNOR U8413 ( .A(n7556), .B(n7555), .Z(n7937) );
  XNOR U8414 ( .A(n7558), .B(n7557), .Z(n7936) );
  OR U8415 ( .A(n7937), .B(n7936), .Z(n7559) );
  NAND U8416 ( .A(n7560), .B(n7559), .Z(n7564) );
  XOR U8417 ( .A(n7562), .B(n7561), .Z(n7563) );
  NANDN U8418 ( .A(n7564), .B(n7563), .Z(n7566) );
  NAND U8419 ( .A(a[6]), .B(b[37]), .Z(n7945) );
  NANDN U8420 ( .A(n7945), .B(n7944), .Z(n7565) );
  NAND U8421 ( .A(n7566), .B(n7565), .Z(n7567) );
  ANDN U8422 ( .B(b[37]), .A(n166), .Z(n7568) );
  OR U8423 ( .A(n7567), .B(n7568), .Z(n7572) );
  XNOR U8424 ( .A(n7568), .B(n7567), .Z(n7949) );
  XOR U8425 ( .A(n7570), .B(n7569), .Z(n7948) );
  NANDN U8426 ( .A(n7949), .B(n7948), .Z(n7571) );
  NAND U8427 ( .A(n7572), .B(n7571), .Z(n7574) );
  AND U8428 ( .A(b[37]), .B(a[8]), .Z(n7573) );
  NANDN U8429 ( .A(n7574), .B(n7573), .Z(n7578) );
  XOR U8430 ( .A(n7574), .B(n7573), .Z(n7956) );
  XOR U8431 ( .A(n7576), .B(n7575), .Z(n7957) );
  NANDN U8432 ( .A(n7956), .B(n7957), .Z(n7577) );
  NAND U8433 ( .A(n7578), .B(n7577), .Z(n7579) );
  ANDN U8434 ( .B(b[37]), .A(n21615), .Z(n7580) );
  OR U8435 ( .A(n7579), .B(n7580), .Z(n7584) );
  XNOR U8436 ( .A(n7580), .B(n7579), .Z(n7961) );
  XNOR U8437 ( .A(n7582), .B(n7581), .Z(n7960) );
  OR U8438 ( .A(n7961), .B(n7960), .Z(n7583) );
  NAND U8439 ( .A(n7584), .B(n7583), .Z(n7588) );
  XOR U8440 ( .A(n7586), .B(n7585), .Z(n7587) );
  NANDN U8441 ( .A(n7588), .B(n7587), .Z(n7590) );
  NAND U8442 ( .A(a[10]), .B(b[37]), .Z(n7967) );
  NANDN U8443 ( .A(n7967), .B(n7966), .Z(n7589) );
  NAND U8444 ( .A(n7590), .B(n7589), .Z(n7591) );
  ANDN U8445 ( .B(b[37]), .A(n21164), .Z(n7592) );
  OR U8446 ( .A(n7591), .B(n7592), .Z(n7596) );
  XNOR U8447 ( .A(n7592), .B(n7591), .Z(n7973) );
  XNOR U8448 ( .A(n7594), .B(n7593), .Z(n7972) );
  OR U8449 ( .A(n7973), .B(n7972), .Z(n7595) );
  NAND U8450 ( .A(n7596), .B(n7595), .Z(n7598) );
  AND U8451 ( .A(b[37]), .B(a[12]), .Z(n7597) );
  NANDN U8452 ( .A(n7598), .B(n7597), .Z(n7602) );
  XOR U8453 ( .A(n7598), .B(n7597), .Z(n7980) );
  XOR U8454 ( .A(n7600), .B(n7599), .Z(n7981) );
  NANDN U8455 ( .A(n7980), .B(n7981), .Z(n7601) );
  NAND U8456 ( .A(n7602), .B(n7601), .Z(n7603) );
  ANDN U8457 ( .B(b[37]), .A(n170), .Z(n7604) );
  OR U8458 ( .A(n7603), .B(n7604), .Z(n7608) );
  XNOR U8459 ( .A(n7604), .B(n7603), .Z(n7985) );
  XOR U8460 ( .A(n7606), .B(n7605), .Z(n7984) );
  NANDN U8461 ( .A(n7985), .B(n7984), .Z(n7607) );
  NAND U8462 ( .A(n7608), .B(n7607), .Z(n7612) );
  XOR U8463 ( .A(n7610), .B(n7609), .Z(n7611) );
  NANDN U8464 ( .A(n7612), .B(n7611), .Z(n7614) );
  NAND U8465 ( .A(a[14]), .B(b[37]), .Z(n7993) );
  NANDN U8466 ( .A(n7993), .B(n7992), .Z(n7613) );
  NAND U8467 ( .A(n7614), .B(n7613), .Z(n7615) );
  ANDN U8468 ( .B(b[37]), .A(n172), .Z(n7616) );
  OR U8469 ( .A(n7615), .B(n7616), .Z(n7620) );
  XNOR U8470 ( .A(n7616), .B(n7615), .Z(n7997) );
  XNOR U8471 ( .A(n7618), .B(n7617), .Z(n7996) );
  OR U8472 ( .A(n7997), .B(n7996), .Z(n7619) );
  NAND U8473 ( .A(n7620), .B(n7619), .Z(n7624) );
  XOR U8474 ( .A(n7622), .B(n7621), .Z(n7623) );
  NANDN U8475 ( .A(n7624), .B(n7623), .Z(n7626) );
  NAND U8476 ( .A(a[16]), .B(b[37]), .Z(n8003) );
  NANDN U8477 ( .A(n8003), .B(n8002), .Z(n7625) );
  NAND U8478 ( .A(n7626), .B(n7625), .Z(n7627) );
  ANDN U8479 ( .B(b[37]), .A(n174), .Z(n7628) );
  OR U8480 ( .A(n7627), .B(n7628), .Z(n7632) );
  XNOR U8481 ( .A(n7628), .B(n7627), .Z(n8009) );
  XOR U8482 ( .A(n7630), .B(n7629), .Z(n8008) );
  NANDN U8483 ( .A(n8009), .B(n8008), .Z(n7631) );
  NAND U8484 ( .A(n7632), .B(n7631), .Z(n7636) );
  XOR U8485 ( .A(n7634), .B(n7633), .Z(n7635) );
  NANDN U8486 ( .A(n7636), .B(n7635), .Z(n7638) );
  NAND U8487 ( .A(a[18]), .B(b[37]), .Z(n8015) );
  NANDN U8488 ( .A(n8015), .B(n8014), .Z(n7637) );
  NAND U8489 ( .A(n7638), .B(n7637), .Z(n7639) );
  ANDN U8490 ( .B(b[37]), .A(n21670), .Z(n7640) );
  OR U8491 ( .A(n7639), .B(n7640), .Z(n7644) );
  XNOR U8492 ( .A(n7640), .B(n7639), .Z(n8021) );
  XNOR U8493 ( .A(n7642), .B(n7641), .Z(n8020) );
  OR U8494 ( .A(n8021), .B(n8020), .Z(n7643) );
  NAND U8495 ( .A(n7644), .B(n7643), .Z(n7648) );
  XOR U8496 ( .A(n7646), .B(n7645), .Z(n7647) );
  NANDN U8497 ( .A(n7648), .B(n7647), .Z(n7650) );
  NAND U8498 ( .A(a[20]), .B(b[37]), .Z(n8027) );
  NANDN U8499 ( .A(n8027), .B(n8026), .Z(n7649) );
  AND U8500 ( .A(n7650), .B(n7649), .Z(n7652) );
  OR U8501 ( .A(n7651), .B(n7652), .Z(n7656) );
  XNOR U8502 ( .A(n7652), .B(n7651), .Z(n8032) );
  XOR U8503 ( .A(n7654), .B(n7653), .Z(n8033) );
  NANDN U8504 ( .A(n8032), .B(n8033), .Z(n7655) );
  AND U8505 ( .A(n7656), .B(n7655), .Z(n7660) );
  XOR U8506 ( .A(n7658), .B(n7657), .Z(n7659) );
  NANDN U8507 ( .A(n7660), .B(n7659), .Z(n7662) );
  AND U8508 ( .A(b[37]), .B(a[22]), .Z(n8040) );
  NANDN U8509 ( .A(n8041), .B(n8040), .Z(n7661) );
  NAND U8510 ( .A(n7662), .B(n7661), .Z(n7663) );
  ANDN U8511 ( .B(b[37]), .A(n21692), .Z(n7664) );
  OR U8512 ( .A(n7663), .B(n7664), .Z(n7668) );
  XNOR U8513 ( .A(n7664), .B(n7663), .Z(n8045) );
  XNOR U8514 ( .A(n7666), .B(n7665), .Z(n8044) );
  OR U8515 ( .A(n8045), .B(n8044), .Z(n7667) );
  NAND U8516 ( .A(n7668), .B(n7667), .Z(n7672) );
  XOR U8517 ( .A(n7670), .B(n7669), .Z(n7671) );
  NANDN U8518 ( .A(n7672), .B(n7671), .Z(n7674) );
  AND U8519 ( .A(b[37]), .B(a[24]), .Z(n8052) );
  NANDN U8520 ( .A(n8053), .B(n8052), .Z(n7673) );
  NAND U8521 ( .A(n7674), .B(n7673), .Z(n7675) );
  ANDN U8522 ( .B(b[37]), .A(n21703), .Z(n7676) );
  OR U8523 ( .A(n7675), .B(n7676), .Z(n7680) );
  XNOR U8524 ( .A(n7676), .B(n7675), .Z(n8057) );
  XNOR U8525 ( .A(n7678), .B(n7677), .Z(n8056) );
  OR U8526 ( .A(n8057), .B(n8056), .Z(n7679) );
  NAND U8527 ( .A(n7680), .B(n7679), .Z(n7684) );
  XOR U8528 ( .A(n7682), .B(n7681), .Z(n7683) );
  NANDN U8529 ( .A(n7684), .B(n7683), .Z(n7686) );
  AND U8530 ( .A(b[37]), .B(a[26]), .Z(n8064) );
  NANDN U8531 ( .A(n8065), .B(n8064), .Z(n7685) );
  NAND U8532 ( .A(n7686), .B(n7685), .Z(n7687) );
  ANDN U8533 ( .B(b[37]), .A(n21716), .Z(n7688) );
  OR U8534 ( .A(n7687), .B(n7688), .Z(n7692) );
  XNOR U8535 ( .A(n7688), .B(n7687), .Z(n8071) );
  XNOR U8536 ( .A(n7690), .B(n7689), .Z(n8070) );
  OR U8537 ( .A(n8071), .B(n8070), .Z(n7691) );
  NAND U8538 ( .A(n7692), .B(n7691), .Z(n7694) );
  NAND U8539 ( .A(a[28]), .B(b[37]), .Z(n7693) );
  OR U8540 ( .A(n7694), .B(n7693), .Z(n7698) );
  XOR U8541 ( .A(n7694), .B(n7693), .Z(n8074) );
  NAND U8542 ( .A(n8074), .B(n8075), .Z(n7697) );
  NAND U8543 ( .A(n7698), .B(n7697), .Z(n7699) );
  NANDN U8544 ( .A(n7700), .B(n7699), .Z(n7704) );
  NAND U8545 ( .A(n8082), .B(n8083), .Z(n7703) );
  NAND U8546 ( .A(n7704), .B(n7703), .Z(n7707) );
  NANDN U8547 ( .A(n7708), .B(n7707), .Z(n7710) );
  NAND U8548 ( .A(n8087), .B(n8086), .Z(n7709) );
  NAND U8549 ( .A(n7710), .B(n7709), .Z(n7711) );
  NANDN U8550 ( .A(n7712), .B(n7711), .Z(n7716) );
  NAND U8551 ( .A(n8094), .B(n8095), .Z(n7715) );
  NAND U8552 ( .A(n7716), .B(n7715), .Z(n7719) );
  NANDN U8553 ( .A(n7720), .B(n7719), .Z(n7722) );
  NAND U8554 ( .A(n8099), .B(n8098), .Z(n7721) );
  NAND U8555 ( .A(n7722), .B(n7721), .Z(n7723) );
  NANDN U8556 ( .A(n7724), .B(n7723), .Z(n7728) );
  NAND U8557 ( .A(n8106), .B(n8107), .Z(n7727) );
  NAND U8558 ( .A(n7728), .B(n7727), .Z(n7731) );
  NANDN U8559 ( .A(n7732), .B(n7731), .Z(n7734) );
  NAND U8560 ( .A(n8111), .B(n8110), .Z(n7733) );
  NAND U8561 ( .A(n7734), .B(n7733), .Z(n7735) );
  NANDN U8562 ( .A(n7736), .B(n7735), .Z(n7740) );
  NAND U8563 ( .A(n8118), .B(n8119), .Z(n7739) );
  NAND U8564 ( .A(n7740), .B(n7739), .Z(n7743) );
  NANDN U8565 ( .A(n7744), .B(n7743), .Z(n7746) );
  NAND U8566 ( .A(n8123), .B(n8122), .Z(n7745) );
  NAND U8567 ( .A(n7746), .B(n7745), .Z(n7747) );
  NANDN U8568 ( .A(n7748), .B(n7747), .Z(n7752) );
  NAND U8569 ( .A(n8130), .B(n8131), .Z(n7751) );
  NAND U8570 ( .A(n7752), .B(n7751), .Z(n7755) );
  NANDN U8571 ( .A(n7756), .B(n7755), .Z(n7758) );
  NAND U8572 ( .A(n8135), .B(n8134), .Z(n7757) );
  NAND U8573 ( .A(n7758), .B(n7757), .Z(n7759) );
  NANDN U8574 ( .A(n7760), .B(n7759), .Z(n7764) );
  NAND U8575 ( .A(n8142), .B(n8143), .Z(n7763) );
  NAND U8576 ( .A(n7764), .B(n7763), .Z(n7767) );
  NANDN U8577 ( .A(n7768), .B(n7767), .Z(n7770) );
  NAND U8578 ( .A(n8147), .B(n8146), .Z(n7769) );
  NAND U8579 ( .A(n7770), .B(n7769), .Z(n7771) );
  NANDN U8580 ( .A(n7772), .B(n7771), .Z(n7776) );
  NAND U8581 ( .A(n8154), .B(n8155), .Z(n7775) );
  NAND U8582 ( .A(n7776), .B(n7775), .Z(n7779) );
  NANDN U8583 ( .A(n7780), .B(n7779), .Z(n7782) );
  NAND U8584 ( .A(n8159), .B(n8158), .Z(n7781) );
  NAND U8585 ( .A(n7782), .B(n7781), .Z(n7783) );
  NANDN U8586 ( .A(n7784), .B(n7783), .Z(n7788) );
  NAND U8587 ( .A(n8166), .B(n8167), .Z(n7787) );
  NAND U8588 ( .A(n7788), .B(n7787), .Z(n7791) );
  NANDN U8589 ( .A(n7792), .B(n7791), .Z(n7794) );
  NAND U8590 ( .A(n8171), .B(n8170), .Z(n7793) );
  NAND U8591 ( .A(n7794), .B(n7793), .Z(n7795) );
  NANDN U8592 ( .A(n7796), .B(n7795), .Z(n7800) );
  NAND U8593 ( .A(n8178), .B(n8179), .Z(n7799) );
  NAND U8594 ( .A(n7800), .B(n7799), .Z(n7803) );
  NANDN U8595 ( .A(n7804), .B(n7803), .Z(n7806) );
  XNOR U8596 ( .A(n7802), .B(n7801), .Z(n8183) );
  NAND U8597 ( .A(n8183), .B(n8182), .Z(n7805) );
  NAND U8598 ( .A(n7806), .B(n7805), .Z(n7807) );
  NANDN U8599 ( .A(n7808), .B(n7807), .Z(n7812) );
  NAND U8600 ( .A(n8190), .B(n8191), .Z(n7811) );
  NAND U8601 ( .A(n7812), .B(n7811), .Z(n7815) );
  NANDN U8602 ( .A(n7816), .B(n7815), .Z(n7818) );
  NAND U8603 ( .A(n8195), .B(n8194), .Z(n7817) );
  NAND U8604 ( .A(n7818), .B(n7817), .Z(n7819) );
  NANDN U8605 ( .A(n7820), .B(n7819), .Z(n7824) );
  XNOR U8606 ( .A(n7822), .B(n7821), .Z(n8203) );
  NAND U8607 ( .A(n8202), .B(n8203), .Z(n7823) );
  NAND U8608 ( .A(n7824), .B(n7823), .Z(n7827) );
  NANDN U8609 ( .A(n7828), .B(n7827), .Z(n7830) );
  NAND U8610 ( .A(n8207), .B(n8206), .Z(n7829) );
  NAND U8611 ( .A(n7830), .B(n7829), .Z(n7831) );
  NANDN U8612 ( .A(n7832), .B(n7831), .Z(n7836) );
  NAND U8613 ( .A(n8214), .B(n8215), .Z(n7835) );
  NAND U8614 ( .A(n7836), .B(n7835), .Z(n7839) );
  NANDN U8615 ( .A(n7840), .B(n7839), .Z(n7842) );
  NAND U8616 ( .A(n8219), .B(n8218), .Z(n7841) );
  NAND U8617 ( .A(n7842), .B(n7841), .Z(n7843) );
  NANDN U8618 ( .A(n7844), .B(n7843), .Z(n7848) );
  NAND U8619 ( .A(n8226), .B(n8227), .Z(n7847) );
  NAND U8620 ( .A(n7848), .B(n7847), .Z(n7851) );
  NANDN U8621 ( .A(n7852), .B(n7851), .Z(n7854) );
  NAND U8622 ( .A(n8231), .B(n8230), .Z(n7853) );
  NAND U8623 ( .A(n7854), .B(n7853), .Z(n7855) );
  NANDN U8624 ( .A(n7856), .B(n7855), .Z(n7860) );
  NAND U8625 ( .A(n8238), .B(n8239), .Z(n7859) );
  NAND U8626 ( .A(n7860), .B(n7859), .Z(n7863) );
  NANDN U8627 ( .A(n7864), .B(n7863), .Z(n7866) );
  NAND U8628 ( .A(n8243), .B(n8242), .Z(n7865) );
  NAND U8629 ( .A(n7866), .B(n7865), .Z(n7867) );
  NANDN U8630 ( .A(n7868), .B(n7867), .Z(n7872) );
  NAND U8631 ( .A(n8250), .B(n8251), .Z(n7871) );
  NAND U8632 ( .A(n7872), .B(n7871), .Z(n7875) );
  NANDN U8633 ( .A(n7876), .B(n7875), .Z(n7878) );
  NAND U8634 ( .A(n8255), .B(n8254), .Z(n7877) );
  NAND U8635 ( .A(n7878), .B(n7877), .Z(n7879) );
  NANDN U8636 ( .A(n7880), .B(n7879), .Z(n7884) );
  NAND U8637 ( .A(n8262), .B(n8263), .Z(n7883) );
  NAND U8638 ( .A(n7884), .B(n7883), .Z(n7887) );
  NANDN U8639 ( .A(n7888), .B(n7887), .Z(n7890) );
  XNOR U8640 ( .A(n7886), .B(n7885), .Z(n8267) );
  NAND U8641 ( .A(n8267), .B(n8266), .Z(n7889) );
  NAND U8642 ( .A(n7890), .B(n7889), .Z(n7891) );
  NANDN U8643 ( .A(n7892), .B(n7891), .Z(n7896) );
  NAND U8644 ( .A(n8274), .B(n8275), .Z(n7895) );
  AND U8645 ( .A(n7896), .B(n7895), .Z(n7898) );
  OR U8646 ( .A(n7897), .B(n7898), .Z(n7902) );
  XNOR U8647 ( .A(n7898), .B(n7897), .Z(n8281) );
  XOR U8648 ( .A(n7900), .B(n7899), .Z(n8280) );
  NANDN U8649 ( .A(n8281), .B(n8280), .Z(n7901) );
  NAND U8650 ( .A(n7902), .B(n7901), .Z(n7903) );
  OR U8651 ( .A(n7904), .B(n7903), .Z(n7906) );
  XNOR U8652 ( .A(n7904), .B(n7903), .Z(n7908) );
  ANDN U8653 ( .B(b[37]), .A(n210), .Z(n7907) );
  OR U8654 ( .A(n7908), .B(n7907), .Z(n7905) );
  NAND U8655 ( .A(n7906), .B(n7905), .Z(n22006) );
  XOR U8656 ( .A(n22005), .B(n22006), .Z(n24210) );
  XOR U8657 ( .A(n7908), .B(n7907), .Z(n8663) );
  ANDN U8658 ( .B(b[36]), .A(n209), .Z(n8269) );
  ANDN U8659 ( .B(b[36]), .A(n207), .Z(n8257) );
  ANDN U8660 ( .B(b[36]), .A(n205), .Z(n8245) );
  ANDN U8661 ( .B(b[36]), .A(n203), .Z(n8233) );
  ANDN U8662 ( .B(b[36]), .A(n201), .Z(n8221) );
  ANDN U8663 ( .B(b[36]), .A(n199), .Z(n8209) );
  ANDN U8664 ( .B(b[36]), .A(n197), .Z(n8197) );
  ANDN U8665 ( .B(b[36]), .A(n195), .Z(n8185) );
  ANDN U8666 ( .B(b[36]), .A(n193), .Z(n8173) );
  ANDN U8667 ( .B(b[36]), .A(n191), .Z(n8161) );
  ANDN U8668 ( .B(b[36]), .A(n189), .Z(n8149) );
  ANDN U8669 ( .B(b[36]), .A(n187), .Z(n8137) );
  ANDN U8670 ( .B(b[36]), .A(n21772), .Z(n8125) );
  ANDN U8671 ( .B(b[36]), .A(n184), .Z(n8113) );
  ANDN U8672 ( .B(b[36]), .A(n21751), .Z(n8101) );
  ANDN U8673 ( .B(b[36]), .A(n21740), .Z(n8089) );
  NAND U8674 ( .A(a[30]), .B(b[36]), .Z(n8081) );
  NAND U8675 ( .A(a[28]), .B(b[36]), .Z(n8068) );
  NAND U8676 ( .A(a[27]), .B(b[36]), .Z(n8062) );
  NAND U8677 ( .A(a[25]), .B(b[36]), .Z(n8050) );
  NAND U8678 ( .A(a[23]), .B(b[36]), .Z(n8039) );
  ANDN U8679 ( .B(b[36]), .A(n21670), .Z(n8016) );
  ANDN U8680 ( .B(b[36]), .A(n172), .Z(n7990) );
  ANDN U8681 ( .B(b[36]), .A(n21615), .Z(n7954) );
  ANDN U8682 ( .B(b[36]), .A(n21580), .Z(n7918) );
  NAND U8683 ( .A(b[37]), .B(a[1]), .Z(n7913) );
  NANDN U8684 ( .A(n7913), .B(a[0]), .Z(n7909) );
  XNOR U8685 ( .A(a[2]), .B(n7909), .Z(n7910) );
  NAND U8686 ( .A(b[36]), .B(n7910), .Z(n8298) );
  AND U8687 ( .A(a[1]), .B(b[37]), .Z(n7911) );
  XOR U8688 ( .A(n7912), .B(n7911), .Z(n8299) );
  OR U8689 ( .A(n8298), .B(n8299), .Z(n7917) );
  AND U8690 ( .A(b[36]), .B(a[0]), .Z(n8671) );
  NANDN U8691 ( .A(n7913), .B(n8671), .Z(n7915) );
  NAND U8692 ( .A(a[2]), .B(b[36]), .Z(n7914) );
  AND U8693 ( .A(n7915), .B(n7914), .Z(n7916) );
  ANDN U8694 ( .B(n7917), .A(n7916), .Z(n7919) );
  OR U8695 ( .A(n7918), .B(n7919), .Z(n7923) );
  XNOR U8696 ( .A(n7919), .B(n7918), .Z(n8303) );
  XNOR U8697 ( .A(n7921), .B(n7920), .Z(n8302) );
  OR U8698 ( .A(n8303), .B(n8302), .Z(n7922) );
  NAND U8699 ( .A(n7923), .B(n7922), .Z(n7926) );
  XOR U8700 ( .A(n7925), .B(n7924), .Z(n7927) );
  OR U8701 ( .A(n7926), .B(n7927), .Z(n7929) );
  XNOR U8702 ( .A(n7927), .B(n7926), .Z(n8311) );
  AND U8703 ( .A(b[36]), .B(a[4]), .Z(n8310) );
  NANDN U8704 ( .A(n8311), .B(n8310), .Z(n7928) );
  NAND U8705 ( .A(n7929), .B(n7928), .Z(n7930) );
  ANDN U8706 ( .B(b[36]), .A(n164), .Z(n7931) );
  OR U8707 ( .A(n7930), .B(n7931), .Z(n7935) );
  XNOR U8708 ( .A(n7931), .B(n7930), .Z(n8315) );
  XNOR U8709 ( .A(n7933), .B(n7932), .Z(n8314) );
  OR U8710 ( .A(n8315), .B(n8314), .Z(n7934) );
  NAND U8711 ( .A(n7935), .B(n7934), .Z(n7938) );
  XOR U8712 ( .A(n7937), .B(n7936), .Z(n7939) );
  OR U8713 ( .A(n7938), .B(n7939), .Z(n7941) );
  XNOR U8714 ( .A(n7939), .B(n7938), .Z(n8323) );
  AND U8715 ( .A(b[36]), .B(a[6]), .Z(n8322) );
  NANDN U8716 ( .A(n8323), .B(n8322), .Z(n7940) );
  NAND U8717 ( .A(n7941), .B(n7940), .Z(n7942) );
  ANDN U8718 ( .B(b[36]), .A(n166), .Z(n7943) );
  OR U8719 ( .A(n7942), .B(n7943), .Z(n7947) );
  XNOR U8720 ( .A(n7943), .B(n7942), .Z(n8326) );
  OR U8721 ( .A(n8326), .B(n8327), .Z(n7946) );
  AND U8722 ( .A(n7947), .B(n7946), .Z(n7951) );
  NANDN U8723 ( .A(n7951), .B(n7950), .Z(n7953) );
  XOR U8724 ( .A(n7951), .B(n7950), .Z(n8332) );
  ANDN U8725 ( .B(b[36]), .A(n167), .Z(n8333) );
  OR U8726 ( .A(n8332), .B(n8333), .Z(n7952) );
  AND U8727 ( .A(n7953), .B(n7952), .Z(n7955) );
  OR U8728 ( .A(n7954), .B(n7955), .Z(n7959) );
  XOR U8729 ( .A(n7955), .B(n7954), .Z(n8338) );
  XOR U8730 ( .A(n7957), .B(n7956), .Z(n8339) );
  NAND U8731 ( .A(n8338), .B(n8339), .Z(n7958) );
  NAND U8732 ( .A(n7959), .B(n7958), .Z(n7962) );
  XOR U8733 ( .A(n7961), .B(n7960), .Z(n7963) );
  OR U8734 ( .A(n7962), .B(n7963), .Z(n7965) );
  NAND U8735 ( .A(a[10]), .B(b[36]), .Z(n8345) );
  XOR U8736 ( .A(n7963), .B(n7962), .Z(n8344) );
  NANDN U8737 ( .A(n8345), .B(n8344), .Z(n7964) );
  NAND U8738 ( .A(n7965), .B(n7964), .Z(n7968) );
  ANDN U8739 ( .B(b[36]), .A(n21164), .Z(n7969) );
  OR U8740 ( .A(n7968), .B(n7969), .Z(n7971) );
  XOR U8741 ( .A(n7969), .B(n7968), .Z(n8350) );
  NANDN U8742 ( .A(n8351), .B(n8350), .Z(n7970) );
  NAND U8743 ( .A(n7971), .B(n7970), .Z(n7974) );
  XOR U8744 ( .A(n7973), .B(n7972), .Z(n7975) );
  OR U8745 ( .A(n7974), .B(n7975), .Z(n7977) );
  XNOR U8746 ( .A(n7975), .B(n7974), .Z(n8359) );
  AND U8747 ( .A(b[36]), .B(a[12]), .Z(n8358) );
  NANDN U8748 ( .A(n8359), .B(n8358), .Z(n7976) );
  NAND U8749 ( .A(n7977), .B(n7976), .Z(n7978) );
  ANDN U8750 ( .B(b[36]), .A(n170), .Z(n7979) );
  OR U8751 ( .A(n7978), .B(n7979), .Z(n7983) );
  XOR U8752 ( .A(n7979), .B(n7978), .Z(n8362) );
  XOR U8753 ( .A(n7981), .B(n7980), .Z(n8363) );
  NAND U8754 ( .A(n8362), .B(n8363), .Z(n7982) );
  AND U8755 ( .A(n7983), .B(n7982), .Z(n7987) );
  NANDN U8756 ( .A(n7987), .B(n7986), .Z(n7989) );
  XOR U8757 ( .A(n7987), .B(n7986), .Z(n8368) );
  ANDN U8758 ( .B(b[36]), .A(n171), .Z(n8369) );
  OR U8759 ( .A(n8368), .B(n8369), .Z(n7988) );
  AND U8760 ( .A(n7989), .B(n7988), .Z(n7991) );
  OR U8761 ( .A(n7990), .B(n7991), .Z(n7995) );
  XNOR U8762 ( .A(n7991), .B(n7990), .Z(n8374) );
  OR U8763 ( .A(n8374), .B(n8375), .Z(n7994) );
  NAND U8764 ( .A(n7995), .B(n7994), .Z(n7998) );
  XOR U8765 ( .A(n7997), .B(n7996), .Z(n7999) );
  OR U8766 ( .A(n7998), .B(n7999), .Z(n8001) );
  NAND U8767 ( .A(a[16]), .B(b[36]), .Z(n8381) );
  XOR U8768 ( .A(n7999), .B(n7998), .Z(n8380) );
  NANDN U8769 ( .A(n8381), .B(n8380), .Z(n8000) );
  NAND U8770 ( .A(n8001), .B(n8000), .Z(n8004) );
  ANDN U8771 ( .B(b[36]), .A(n174), .Z(n8005) );
  OR U8772 ( .A(n8004), .B(n8005), .Z(n8007) );
  XOR U8773 ( .A(n8005), .B(n8004), .Z(n8386) );
  NANDN U8774 ( .A(n8387), .B(n8386), .Z(n8006) );
  AND U8775 ( .A(n8007), .B(n8006), .Z(n8011) );
  NANDN U8776 ( .A(n8011), .B(n8010), .Z(n8013) );
  XOR U8777 ( .A(n8011), .B(n8010), .Z(n8392) );
  ANDN U8778 ( .B(b[36]), .A(n175), .Z(n8393) );
  OR U8779 ( .A(n8392), .B(n8393), .Z(n8012) );
  AND U8780 ( .A(n8013), .B(n8012), .Z(n8017) );
  OR U8781 ( .A(n8016), .B(n8017), .Z(n8019) );
  XOR U8782 ( .A(n8017), .B(n8016), .Z(n8398) );
  NANDN U8783 ( .A(n8399), .B(n8398), .Z(n8018) );
  NAND U8784 ( .A(n8019), .B(n8018), .Z(n8022) );
  XOR U8785 ( .A(n8021), .B(n8020), .Z(n8023) );
  OR U8786 ( .A(n8022), .B(n8023), .Z(n8025) );
  NAND U8787 ( .A(a[20]), .B(b[36]), .Z(n8407) );
  XOR U8788 ( .A(n8023), .B(n8022), .Z(n8406) );
  NANDN U8789 ( .A(n8407), .B(n8406), .Z(n8024) );
  NAND U8790 ( .A(n8025), .B(n8024), .Z(n8028) );
  ANDN U8791 ( .B(b[36]), .A(n21681), .Z(n8029) );
  OR U8792 ( .A(n8028), .B(n8029), .Z(n8031) );
  XOR U8793 ( .A(n8029), .B(n8028), .Z(n8410) );
  NANDN U8794 ( .A(n8411), .B(n8410), .Z(n8030) );
  AND U8795 ( .A(n8031), .B(n8030), .Z(n8034) );
  XNOR U8796 ( .A(n8033), .B(n8032), .Z(n8035) );
  OR U8797 ( .A(n8034), .B(n8035), .Z(n8037) );
  XNOR U8798 ( .A(n8035), .B(n8034), .Z(n8418) );
  ANDN U8799 ( .B(b[36]), .A(n177), .Z(n8419) );
  OR U8800 ( .A(n8418), .B(n8419), .Z(n8036) );
  NAND U8801 ( .A(n8037), .B(n8036), .Z(n8038) );
  OR U8802 ( .A(n8039), .B(n8038), .Z(n8043) );
  XNOR U8803 ( .A(n8039), .B(n8038), .Z(n8423) );
  XOR U8804 ( .A(n8041), .B(n8040), .Z(n8422) );
  OR U8805 ( .A(n8423), .B(n8422), .Z(n8042) );
  AND U8806 ( .A(n8043), .B(n8042), .Z(n8046) );
  XOR U8807 ( .A(n8045), .B(n8044), .Z(n8047) );
  OR U8808 ( .A(n8046), .B(n8047), .Z(n8049) );
  NAND U8809 ( .A(a[24]), .B(b[36]), .Z(n8429) );
  XOR U8810 ( .A(n8047), .B(n8046), .Z(n8428) );
  NANDN U8811 ( .A(n8429), .B(n8428), .Z(n8048) );
  AND U8812 ( .A(n8049), .B(n8048), .Z(n8051) );
  OR U8813 ( .A(n8050), .B(n8051), .Z(n8055) );
  XNOR U8814 ( .A(n8051), .B(n8050), .Z(n8435) );
  XOR U8815 ( .A(n8053), .B(n8052), .Z(n8434) );
  OR U8816 ( .A(n8435), .B(n8434), .Z(n8054) );
  AND U8817 ( .A(n8055), .B(n8054), .Z(n8058) );
  XOR U8818 ( .A(n8057), .B(n8056), .Z(n8059) );
  OR U8819 ( .A(n8058), .B(n8059), .Z(n8061) );
  NAND U8820 ( .A(a[26]), .B(b[36]), .Z(n8441) );
  XOR U8821 ( .A(n8059), .B(n8058), .Z(n8440) );
  NANDN U8822 ( .A(n8441), .B(n8440), .Z(n8060) );
  AND U8823 ( .A(n8061), .B(n8060), .Z(n8063) );
  OR U8824 ( .A(n8062), .B(n8063), .Z(n8067) );
  XNOR U8825 ( .A(n8063), .B(n8062), .Z(n8447) );
  XOR U8826 ( .A(n8065), .B(n8064), .Z(n8446) );
  OR U8827 ( .A(n8447), .B(n8446), .Z(n8066) );
  AND U8828 ( .A(n8067), .B(n8066), .Z(n8069) );
  OR U8829 ( .A(n8068), .B(n8069), .Z(n8073) );
  XNOR U8830 ( .A(n8069), .B(n8068), .Z(n8454) );
  XOR U8831 ( .A(n8071), .B(n8070), .Z(n8455) );
  OR U8832 ( .A(n8454), .B(n8455), .Z(n8072) );
  NAND U8833 ( .A(n8073), .B(n8072), .Z(n8077) );
  NAND U8834 ( .A(n8077), .B(n8076), .Z(n8079) );
  XNOR U8835 ( .A(n8077), .B(n8076), .Z(n8459) );
  NAND U8836 ( .A(a[29]), .B(b[36]), .Z(n8458) );
  OR U8837 ( .A(n8459), .B(n8458), .Z(n8078) );
  NAND U8838 ( .A(n8079), .B(n8078), .Z(n8080) );
  NANDN U8839 ( .A(n8081), .B(n8080), .Z(n8085) );
  NAND U8840 ( .A(n8464), .B(n8465), .Z(n8084) );
  NAND U8841 ( .A(n8085), .B(n8084), .Z(n8088) );
  OR U8842 ( .A(n8089), .B(n8088), .Z(n8091) );
  XOR U8843 ( .A(n8087), .B(n8086), .Z(n8471) );
  XOR U8844 ( .A(n8089), .B(n8088), .Z(n8470) );
  NANDN U8845 ( .A(n8471), .B(n8470), .Z(n8090) );
  NAND U8846 ( .A(n8091), .B(n8090), .Z(n8093) );
  NAND U8847 ( .A(a[32]), .B(b[36]), .Z(n8092) );
  OR U8848 ( .A(n8093), .B(n8092), .Z(n8097) );
  XOR U8849 ( .A(n8093), .B(n8092), .Z(n8476) );
  NAND U8850 ( .A(n8476), .B(n8477), .Z(n8096) );
  NAND U8851 ( .A(n8097), .B(n8096), .Z(n8100) );
  OR U8852 ( .A(n8101), .B(n8100), .Z(n8103) );
  XOR U8853 ( .A(n8099), .B(n8098), .Z(n8483) );
  XOR U8854 ( .A(n8101), .B(n8100), .Z(n8482) );
  NANDN U8855 ( .A(n8483), .B(n8482), .Z(n8102) );
  NAND U8856 ( .A(n8103), .B(n8102), .Z(n8105) );
  NAND U8857 ( .A(a[34]), .B(b[36]), .Z(n8104) );
  OR U8858 ( .A(n8105), .B(n8104), .Z(n8109) );
  XOR U8859 ( .A(n8105), .B(n8104), .Z(n8488) );
  NAND U8860 ( .A(n8488), .B(n8489), .Z(n8108) );
  NAND U8861 ( .A(n8109), .B(n8108), .Z(n8112) );
  OR U8862 ( .A(n8113), .B(n8112), .Z(n8115) );
  XOR U8863 ( .A(n8111), .B(n8110), .Z(n8495) );
  XOR U8864 ( .A(n8113), .B(n8112), .Z(n8494) );
  NANDN U8865 ( .A(n8495), .B(n8494), .Z(n8114) );
  NAND U8866 ( .A(n8115), .B(n8114), .Z(n8117) );
  NAND U8867 ( .A(a[36]), .B(b[36]), .Z(n8116) );
  OR U8868 ( .A(n8117), .B(n8116), .Z(n8121) );
  XOR U8869 ( .A(n8117), .B(n8116), .Z(n8500) );
  NAND U8870 ( .A(n8500), .B(n8501), .Z(n8120) );
  NAND U8871 ( .A(n8121), .B(n8120), .Z(n8124) );
  OR U8872 ( .A(n8125), .B(n8124), .Z(n8127) );
  XOR U8873 ( .A(n8123), .B(n8122), .Z(n8507) );
  XOR U8874 ( .A(n8125), .B(n8124), .Z(n8506) );
  NANDN U8875 ( .A(n8507), .B(n8506), .Z(n8126) );
  NAND U8876 ( .A(n8127), .B(n8126), .Z(n8129) );
  NAND U8877 ( .A(a[38]), .B(b[36]), .Z(n8128) );
  OR U8878 ( .A(n8129), .B(n8128), .Z(n8133) );
  XOR U8879 ( .A(n8129), .B(n8128), .Z(n8512) );
  NAND U8880 ( .A(n8512), .B(n8513), .Z(n8132) );
  NAND U8881 ( .A(n8133), .B(n8132), .Z(n8136) );
  OR U8882 ( .A(n8137), .B(n8136), .Z(n8139) );
  XOR U8883 ( .A(n8135), .B(n8134), .Z(n8519) );
  XOR U8884 ( .A(n8137), .B(n8136), .Z(n8518) );
  NANDN U8885 ( .A(n8519), .B(n8518), .Z(n8138) );
  NAND U8886 ( .A(n8139), .B(n8138), .Z(n8141) );
  NAND U8887 ( .A(a[40]), .B(b[36]), .Z(n8140) );
  OR U8888 ( .A(n8141), .B(n8140), .Z(n8145) );
  XOR U8889 ( .A(n8141), .B(n8140), .Z(n8524) );
  NAND U8890 ( .A(n8524), .B(n8525), .Z(n8144) );
  NAND U8891 ( .A(n8145), .B(n8144), .Z(n8148) );
  OR U8892 ( .A(n8149), .B(n8148), .Z(n8151) );
  XOR U8893 ( .A(n8147), .B(n8146), .Z(n8531) );
  XOR U8894 ( .A(n8149), .B(n8148), .Z(n8530) );
  NANDN U8895 ( .A(n8531), .B(n8530), .Z(n8150) );
  NAND U8896 ( .A(n8151), .B(n8150), .Z(n8153) );
  NAND U8897 ( .A(a[42]), .B(b[36]), .Z(n8152) );
  OR U8898 ( .A(n8153), .B(n8152), .Z(n8157) );
  XOR U8899 ( .A(n8153), .B(n8152), .Z(n8536) );
  NAND U8900 ( .A(n8536), .B(n8537), .Z(n8156) );
  NAND U8901 ( .A(n8157), .B(n8156), .Z(n8160) );
  OR U8902 ( .A(n8161), .B(n8160), .Z(n8163) );
  XOR U8903 ( .A(n8159), .B(n8158), .Z(n8543) );
  XOR U8904 ( .A(n8161), .B(n8160), .Z(n8542) );
  NANDN U8905 ( .A(n8543), .B(n8542), .Z(n8162) );
  NAND U8906 ( .A(n8163), .B(n8162), .Z(n8165) );
  NAND U8907 ( .A(a[44]), .B(b[36]), .Z(n8164) );
  OR U8908 ( .A(n8165), .B(n8164), .Z(n8169) );
  XOR U8909 ( .A(n8165), .B(n8164), .Z(n8548) );
  NAND U8910 ( .A(n8548), .B(n8549), .Z(n8168) );
  NAND U8911 ( .A(n8169), .B(n8168), .Z(n8172) );
  OR U8912 ( .A(n8173), .B(n8172), .Z(n8175) );
  XOR U8913 ( .A(n8171), .B(n8170), .Z(n8555) );
  XOR U8914 ( .A(n8173), .B(n8172), .Z(n8554) );
  NANDN U8915 ( .A(n8555), .B(n8554), .Z(n8174) );
  NAND U8916 ( .A(n8175), .B(n8174), .Z(n8177) );
  NAND U8917 ( .A(a[46]), .B(b[36]), .Z(n8176) );
  OR U8918 ( .A(n8177), .B(n8176), .Z(n8181) );
  XOR U8919 ( .A(n8177), .B(n8176), .Z(n8560) );
  NAND U8920 ( .A(n8560), .B(n8561), .Z(n8180) );
  NAND U8921 ( .A(n8181), .B(n8180), .Z(n8184) );
  OR U8922 ( .A(n8185), .B(n8184), .Z(n8187) );
  XOR U8923 ( .A(n8183), .B(n8182), .Z(n8567) );
  XOR U8924 ( .A(n8185), .B(n8184), .Z(n8566) );
  NANDN U8925 ( .A(n8567), .B(n8566), .Z(n8186) );
  NAND U8926 ( .A(n8187), .B(n8186), .Z(n8189) );
  NAND U8927 ( .A(a[48]), .B(b[36]), .Z(n8188) );
  OR U8928 ( .A(n8189), .B(n8188), .Z(n8193) );
  XOR U8929 ( .A(n8189), .B(n8188), .Z(n8572) );
  NAND U8930 ( .A(n8572), .B(n8573), .Z(n8192) );
  NAND U8931 ( .A(n8193), .B(n8192), .Z(n8196) );
  OR U8932 ( .A(n8197), .B(n8196), .Z(n8199) );
  XOR U8933 ( .A(n8195), .B(n8194), .Z(n8579) );
  XOR U8934 ( .A(n8197), .B(n8196), .Z(n8578) );
  NANDN U8935 ( .A(n8579), .B(n8578), .Z(n8198) );
  NAND U8936 ( .A(n8199), .B(n8198), .Z(n8201) );
  NAND U8937 ( .A(a[50]), .B(b[36]), .Z(n8200) );
  OR U8938 ( .A(n8201), .B(n8200), .Z(n8205) );
  XOR U8939 ( .A(n8201), .B(n8200), .Z(n8584) );
  NAND U8940 ( .A(n8584), .B(n8585), .Z(n8204) );
  NAND U8941 ( .A(n8205), .B(n8204), .Z(n8208) );
  OR U8942 ( .A(n8209), .B(n8208), .Z(n8211) );
  XOR U8943 ( .A(n8207), .B(n8206), .Z(n8591) );
  XOR U8944 ( .A(n8209), .B(n8208), .Z(n8590) );
  NANDN U8945 ( .A(n8591), .B(n8590), .Z(n8210) );
  NAND U8946 ( .A(n8211), .B(n8210), .Z(n8213) );
  NAND U8947 ( .A(a[52]), .B(b[36]), .Z(n8212) );
  OR U8948 ( .A(n8213), .B(n8212), .Z(n8217) );
  XOR U8949 ( .A(n8213), .B(n8212), .Z(n8596) );
  NAND U8950 ( .A(n8596), .B(n8597), .Z(n8216) );
  NAND U8951 ( .A(n8217), .B(n8216), .Z(n8220) );
  OR U8952 ( .A(n8221), .B(n8220), .Z(n8223) );
  XOR U8953 ( .A(n8219), .B(n8218), .Z(n8603) );
  XOR U8954 ( .A(n8221), .B(n8220), .Z(n8602) );
  NANDN U8955 ( .A(n8603), .B(n8602), .Z(n8222) );
  NAND U8956 ( .A(n8223), .B(n8222), .Z(n8225) );
  NAND U8957 ( .A(a[54]), .B(b[36]), .Z(n8224) );
  OR U8958 ( .A(n8225), .B(n8224), .Z(n8229) );
  XOR U8959 ( .A(n8225), .B(n8224), .Z(n8608) );
  NAND U8960 ( .A(n8608), .B(n8609), .Z(n8228) );
  NAND U8961 ( .A(n8229), .B(n8228), .Z(n8232) );
  OR U8962 ( .A(n8233), .B(n8232), .Z(n8235) );
  XOR U8963 ( .A(n8231), .B(n8230), .Z(n8615) );
  XOR U8964 ( .A(n8233), .B(n8232), .Z(n8614) );
  NANDN U8965 ( .A(n8615), .B(n8614), .Z(n8234) );
  NAND U8966 ( .A(n8235), .B(n8234), .Z(n8237) );
  NAND U8967 ( .A(a[56]), .B(b[36]), .Z(n8236) );
  OR U8968 ( .A(n8237), .B(n8236), .Z(n8241) );
  XOR U8969 ( .A(n8237), .B(n8236), .Z(n8620) );
  NAND U8970 ( .A(n8620), .B(n8621), .Z(n8240) );
  NAND U8971 ( .A(n8241), .B(n8240), .Z(n8244) );
  OR U8972 ( .A(n8245), .B(n8244), .Z(n8247) );
  XOR U8973 ( .A(n8243), .B(n8242), .Z(n8627) );
  XOR U8974 ( .A(n8245), .B(n8244), .Z(n8626) );
  NANDN U8975 ( .A(n8627), .B(n8626), .Z(n8246) );
  NAND U8976 ( .A(n8247), .B(n8246), .Z(n8249) );
  NAND U8977 ( .A(a[58]), .B(b[36]), .Z(n8248) );
  OR U8978 ( .A(n8249), .B(n8248), .Z(n8253) );
  XOR U8979 ( .A(n8249), .B(n8248), .Z(n8632) );
  NAND U8980 ( .A(n8632), .B(n8633), .Z(n8252) );
  NAND U8981 ( .A(n8253), .B(n8252), .Z(n8256) );
  OR U8982 ( .A(n8257), .B(n8256), .Z(n8259) );
  XOR U8983 ( .A(n8255), .B(n8254), .Z(n8639) );
  XOR U8984 ( .A(n8257), .B(n8256), .Z(n8638) );
  NANDN U8985 ( .A(n8639), .B(n8638), .Z(n8258) );
  NAND U8986 ( .A(n8259), .B(n8258), .Z(n8261) );
  NAND U8987 ( .A(a[60]), .B(b[36]), .Z(n8260) );
  OR U8988 ( .A(n8261), .B(n8260), .Z(n8265) );
  XOR U8989 ( .A(n8261), .B(n8260), .Z(n8644) );
  NAND U8990 ( .A(n8644), .B(n8645), .Z(n8264) );
  NAND U8991 ( .A(n8265), .B(n8264), .Z(n8268) );
  OR U8992 ( .A(n8269), .B(n8268), .Z(n8271) );
  XOR U8993 ( .A(n8267), .B(n8266), .Z(n8651) );
  XOR U8994 ( .A(n8269), .B(n8268), .Z(n8650) );
  NANDN U8995 ( .A(n8651), .B(n8650), .Z(n8270) );
  NAND U8996 ( .A(n8271), .B(n8270), .Z(n8273) );
  NAND U8997 ( .A(a[62]), .B(b[36]), .Z(n8272) );
  OR U8998 ( .A(n8273), .B(n8272), .Z(n8277) );
  XOR U8999 ( .A(n8273), .B(n8272), .Z(n8656) );
  NAND U9000 ( .A(n8656), .B(n8657), .Z(n8276) );
  NAND U9001 ( .A(n8277), .B(n8276), .Z(n8278) );
  ANDN U9002 ( .B(b[36]), .A(n210), .Z(n8279) );
  OR U9003 ( .A(n8278), .B(n8279), .Z(n8283) );
  XOR U9004 ( .A(n8279), .B(n8278), .Z(n8285) );
  NAND U9005 ( .A(n8285), .B(n8286), .Z(n8282) );
  AND U9006 ( .A(n8283), .B(n8282), .Z(n8662) );
  NANDN U9007 ( .A(n8663), .B(n8662), .Z(n8284) );
  NANDN U9008 ( .A(n24210), .B(n8284), .Z(n22004) );
  IV U9009 ( .A(n8284), .Z(n24211) );
  AND U9010 ( .A(n24210), .B(n24211), .Z(n22002) );
  NAND U9011 ( .A(a[63]), .B(b[35]), .Z(n8658) );
  NAND U9012 ( .A(a[54]), .B(b[35]), .Z(n8604) );
  NAND U9013 ( .A(a[53]), .B(b[35]), .Z(n8598) );
  NAND U9014 ( .A(a[46]), .B(b[35]), .Z(n8556) );
  NAND U9015 ( .A(a[45]), .B(b[35]), .Z(n8550) );
  NAND U9016 ( .A(a[42]), .B(b[35]), .Z(n8532) );
  NAND U9017 ( .A(a[41]), .B(b[35]), .Z(n8526) );
  NAND U9018 ( .A(a[38]), .B(b[35]), .Z(n8508) );
  NAND U9019 ( .A(a[36]), .B(b[35]), .Z(n8496) );
  NAND U9020 ( .A(a[34]), .B(b[35]), .Z(n8484) );
  NAND U9021 ( .A(a[32]), .B(b[35]), .Z(n8472) );
  ANDN U9022 ( .B(b[35]), .A(n21727), .Z(n8452) );
  ANDN U9023 ( .B(b[35]), .A(n21716), .Z(n8442) );
  ANDN U9024 ( .B(b[35]), .A(n21703), .Z(n8430) );
  ANDN U9025 ( .B(b[35]), .A(n174), .Z(n8382) );
  NAND U9026 ( .A(a[13]), .B(b[35]), .Z(n8356) );
  ANDN U9027 ( .B(b[35]), .A(n21615), .Z(n8334) );
  NAND U9028 ( .A(a[7]), .B(b[35]), .Z(n8320) );
  NAND U9029 ( .A(a[5]), .B(b[35]), .Z(n8308) );
  ANDN U9030 ( .B(b[35]), .A(n21580), .Z(n8296) );
  NAND U9031 ( .A(b[36]), .B(a[1]), .Z(n8291) );
  NANDN U9032 ( .A(n8291), .B(a[0]), .Z(n8287) );
  XNOR U9033 ( .A(a[2]), .B(n8287), .Z(n8288) );
  NAND U9034 ( .A(b[35]), .B(n8288), .Z(n8679) );
  AND U9035 ( .A(a[1]), .B(b[36]), .Z(n8289) );
  XOR U9036 ( .A(n8290), .B(n8289), .Z(n8680) );
  OR U9037 ( .A(n8679), .B(n8680), .Z(n8295) );
  AND U9038 ( .A(b[35]), .B(a[0]), .Z(n9052) );
  NANDN U9039 ( .A(n8291), .B(n9052), .Z(n8293) );
  NAND U9040 ( .A(a[2]), .B(b[35]), .Z(n8292) );
  AND U9041 ( .A(n8293), .B(n8292), .Z(n8294) );
  ANDN U9042 ( .B(n8295), .A(n8294), .Z(n8297) );
  OR U9043 ( .A(n8296), .B(n8297), .Z(n8301) );
  XNOR U9044 ( .A(n8297), .B(n8296), .Z(n8684) );
  XNOR U9045 ( .A(n8299), .B(n8298), .Z(n8683) );
  OR U9046 ( .A(n8684), .B(n8683), .Z(n8300) );
  NAND U9047 ( .A(n8301), .B(n8300), .Z(n8304) );
  XOR U9048 ( .A(n8303), .B(n8302), .Z(n8305) );
  OR U9049 ( .A(n8304), .B(n8305), .Z(n8307) );
  NAND U9050 ( .A(a[4]), .B(b[35]), .Z(n8692) );
  XOR U9051 ( .A(n8305), .B(n8304), .Z(n8691) );
  NANDN U9052 ( .A(n8692), .B(n8691), .Z(n8306) );
  AND U9053 ( .A(n8307), .B(n8306), .Z(n8309) );
  OR U9054 ( .A(n8308), .B(n8309), .Z(n8313) );
  XNOR U9055 ( .A(n8309), .B(n8308), .Z(n8696) );
  XOR U9056 ( .A(n8311), .B(n8310), .Z(n8695) );
  OR U9057 ( .A(n8696), .B(n8695), .Z(n8312) );
  AND U9058 ( .A(n8313), .B(n8312), .Z(n8316) );
  XOR U9059 ( .A(n8315), .B(n8314), .Z(n8317) );
  OR U9060 ( .A(n8316), .B(n8317), .Z(n8319) );
  NAND U9061 ( .A(a[6]), .B(b[35]), .Z(n8702) );
  XOR U9062 ( .A(n8317), .B(n8316), .Z(n8701) );
  NANDN U9063 ( .A(n8702), .B(n8701), .Z(n8318) );
  AND U9064 ( .A(n8319), .B(n8318), .Z(n8321) );
  OR U9065 ( .A(n8320), .B(n8321), .Z(n8325) );
  XNOR U9066 ( .A(n8321), .B(n8320), .Z(n8708) );
  XOR U9067 ( .A(n8323), .B(n8322), .Z(n8707) );
  OR U9068 ( .A(n8708), .B(n8707), .Z(n8324) );
  NAND U9069 ( .A(n8325), .B(n8324), .Z(n8328) );
  XOR U9070 ( .A(n8327), .B(n8326), .Z(n8329) );
  NANDN U9071 ( .A(n8328), .B(n8329), .Z(n8331) );
  XOR U9072 ( .A(n8329), .B(n8328), .Z(n8715) );
  ANDN U9073 ( .B(b[35]), .A(n167), .Z(n8716) );
  OR U9074 ( .A(n8715), .B(n8716), .Z(n8330) );
  AND U9075 ( .A(n8331), .B(n8330), .Z(n8335) );
  OR U9076 ( .A(n8334), .B(n8335), .Z(n8337) );
  XNOR U9077 ( .A(n8333), .B(n8332), .Z(n8720) );
  XNOR U9078 ( .A(n8335), .B(n8334), .Z(n8719) );
  OR U9079 ( .A(n8720), .B(n8719), .Z(n8336) );
  NAND U9080 ( .A(n8337), .B(n8336), .Z(n8340) );
  OR U9081 ( .A(n8340), .B(n8341), .Z(n8343) );
  NAND U9082 ( .A(a[10]), .B(b[35]), .Z(n8728) );
  XOR U9083 ( .A(n8341), .B(n8340), .Z(n8727) );
  NANDN U9084 ( .A(n8728), .B(n8727), .Z(n8342) );
  NAND U9085 ( .A(n8343), .B(n8342), .Z(n8346) );
  ANDN U9086 ( .B(b[35]), .A(n21164), .Z(n8347) );
  OR U9087 ( .A(n8346), .B(n8347), .Z(n8349) );
  XOR U9088 ( .A(n8347), .B(n8346), .Z(n8731) );
  NANDN U9089 ( .A(n8732), .B(n8731), .Z(n8348) );
  NAND U9090 ( .A(n8349), .B(n8348), .Z(n8352) );
  XNOR U9091 ( .A(n8351), .B(n8350), .Z(n8353) );
  OR U9092 ( .A(n8352), .B(n8353), .Z(n8355) );
  XNOR U9093 ( .A(n8353), .B(n8352), .Z(n8738) );
  NAND U9094 ( .A(a[12]), .B(b[35]), .Z(n8737) );
  OR U9095 ( .A(n8738), .B(n8737), .Z(n8354) );
  AND U9096 ( .A(n8355), .B(n8354), .Z(n8357) );
  OR U9097 ( .A(n8356), .B(n8357), .Z(n8361) );
  XNOR U9098 ( .A(n8357), .B(n8356), .Z(n8744) );
  XOR U9099 ( .A(n8359), .B(n8358), .Z(n8743) );
  OR U9100 ( .A(n8744), .B(n8743), .Z(n8360) );
  AND U9101 ( .A(n8361), .B(n8360), .Z(n8364) );
  OR U9102 ( .A(n8364), .B(n8365), .Z(n8367) );
  NAND U9103 ( .A(a[14]), .B(b[35]), .Z(n8750) );
  XOR U9104 ( .A(n8365), .B(n8364), .Z(n8749) );
  NANDN U9105 ( .A(n8750), .B(n8749), .Z(n8366) );
  NAND U9106 ( .A(n8367), .B(n8366), .Z(n8370) );
  ANDN U9107 ( .B(b[35]), .A(n172), .Z(n8371) );
  OR U9108 ( .A(n8370), .B(n8371), .Z(n8373) );
  XNOR U9109 ( .A(n8369), .B(n8368), .Z(n8756) );
  XNOR U9110 ( .A(n8371), .B(n8370), .Z(n8755) );
  OR U9111 ( .A(n8756), .B(n8755), .Z(n8372) );
  AND U9112 ( .A(n8373), .B(n8372), .Z(n8377) );
  XOR U9113 ( .A(n8375), .B(n8374), .Z(n8376) );
  NANDN U9114 ( .A(n8377), .B(n8376), .Z(n8379) );
  XOR U9115 ( .A(n8377), .B(n8376), .Z(n8763) );
  ANDN U9116 ( .B(b[35]), .A(n173), .Z(n8764) );
  OR U9117 ( .A(n8763), .B(n8764), .Z(n8378) );
  AND U9118 ( .A(n8379), .B(n8378), .Z(n8383) );
  OR U9119 ( .A(n8382), .B(n8383), .Z(n8385) );
  XOR U9120 ( .A(n8383), .B(n8382), .Z(n8767) );
  NANDN U9121 ( .A(n8768), .B(n8767), .Z(n8384) );
  NAND U9122 ( .A(n8385), .B(n8384), .Z(n8388) );
  XNOR U9123 ( .A(n8387), .B(n8386), .Z(n8389) );
  OR U9124 ( .A(n8388), .B(n8389), .Z(n8391) );
  XNOR U9125 ( .A(n8389), .B(n8388), .Z(n8774) );
  NAND U9126 ( .A(a[18]), .B(b[35]), .Z(n8773) );
  OR U9127 ( .A(n8774), .B(n8773), .Z(n8390) );
  NAND U9128 ( .A(n8391), .B(n8390), .Z(n8394) );
  ANDN U9129 ( .B(b[35]), .A(n21670), .Z(n8395) );
  OR U9130 ( .A(n8394), .B(n8395), .Z(n8397) );
  XNOR U9131 ( .A(n8393), .B(n8392), .Z(n8780) );
  XOR U9132 ( .A(n8395), .B(n8394), .Z(n8779) );
  NANDN U9133 ( .A(n8780), .B(n8779), .Z(n8396) );
  NAND U9134 ( .A(n8397), .B(n8396), .Z(n8400) );
  XNOR U9135 ( .A(n8399), .B(n8398), .Z(n8401) );
  OR U9136 ( .A(n8400), .B(n8401), .Z(n8403) );
  XNOR U9137 ( .A(n8401), .B(n8400), .Z(n8788) );
  AND U9138 ( .A(b[35]), .B(a[20]), .Z(n8787) );
  NANDN U9139 ( .A(n8788), .B(n8787), .Z(n8402) );
  NAND U9140 ( .A(n8403), .B(n8402), .Z(n8404) );
  ANDN U9141 ( .B(b[35]), .A(n21681), .Z(n8405) );
  OR U9142 ( .A(n8404), .B(n8405), .Z(n8409) );
  XNOR U9143 ( .A(n8405), .B(n8404), .Z(n8791) );
  OR U9144 ( .A(n8791), .B(n8792), .Z(n8408) );
  NAND U9145 ( .A(n8409), .B(n8408), .Z(n8412) );
  XNOR U9146 ( .A(n8411), .B(n8410), .Z(n8413) );
  OR U9147 ( .A(n8412), .B(n8413), .Z(n8415) );
  XNOR U9148 ( .A(n8413), .B(n8412), .Z(n8800) );
  NAND U9149 ( .A(a[22]), .B(b[35]), .Z(n8799) );
  OR U9150 ( .A(n8800), .B(n8799), .Z(n8414) );
  NAND U9151 ( .A(n8415), .B(n8414), .Z(n8416) );
  ANDN U9152 ( .B(b[35]), .A(n21692), .Z(n8417) );
  OR U9153 ( .A(n8416), .B(n8417), .Z(n8421) );
  XNOR U9154 ( .A(n8417), .B(n8416), .Z(n8804) );
  XNOR U9155 ( .A(n8419), .B(n8418), .Z(n8803) );
  OR U9156 ( .A(n8804), .B(n8803), .Z(n8420) );
  AND U9157 ( .A(n8421), .B(n8420), .Z(n8424) );
  XOR U9158 ( .A(n8423), .B(n8422), .Z(n8425) );
  OR U9159 ( .A(n8424), .B(n8425), .Z(n8427) );
  ANDN U9160 ( .B(b[35]), .A(n178), .Z(n8812) );
  XOR U9161 ( .A(n8425), .B(n8424), .Z(n8811) );
  NANDN U9162 ( .A(n8812), .B(n8811), .Z(n8426) );
  AND U9163 ( .A(n8427), .B(n8426), .Z(n8431) );
  OR U9164 ( .A(n8430), .B(n8431), .Z(n8433) );
  XOR U9165 ( .A(n8431), .B(n8430), .Z(n8815) );
  NANDN U9166 ( .A(n8816), .B(n8815), .Z(n8432) );
  AND U9167 ( .A(n8433), .B(n8432), .Z(n8436) );
  XOR U9168 ( .A(n8435), .B(n8434), .Z(n8437) );
  OR U9169 ( .A(n8436), .B(n8437), .Z(n8439) );
  ANDN U9170 ( .B(b[35]), .A(n179), .Z(n8824) );
  XOR U9171 ( .A(n8437), .B(n8436), .Z(n8823) );
  NANDN U9172 ( .A(n8824), .B(n8823), .Z(n8438) );
  AND U9173 ( .A(n8439), .B(n8438), .Z(n8443) );
  OR U9174 ( .A(n8442), .B(n8443), .Z(n8445) );
  XOR U9175 ( .A(n8443), .B(n8442), .Z(n8827) );
  NANDN U9176 ( .A(n8828), .B(n8827), .Z(n8444) );
  AND U9177 ( .A(n8445), .B(n8444), .Z(n8448) );
  XOR U9178 ( .A(n8447), .B(n8446), .Z(n8449) );
  OR U9179 ( .A(n8448), .B(n8449), .Z(n8451) );
  ANDN U9180 ( .B(b[35]), .A(n180), .Z(n8836) );
  XOR U9181 ( .A(n8449), .B(n8448), .Z(n8835) );
  NANDN U9182 ( .A(n8836), .B(n8835), .Z(n8450) );
  AND U9183 ( .A(n8451), .B(n8450), .Z(n8453) );
  OR U9184 ( .A(n8452), .B(n8453), .Z(n8457) );
  XOR U9185 ( .A(n8453), .B(n8452), .Z(n8839) );
  XNOR U9186 ( .A(n8455), .B(n8454), .Z(n8840) );
  NAND U9187 ( .A(n8839), .B(n8840), .Z(n8456) );
  NAND U9188 ( .A(n8457), .B(n8456), .Z(n8461) );
  NAND U9189 ( .A(a[30]), .B(b[35]), .Z(n8460) );
  OR U9190 ( .A(n8461), .B(n8460), .Z(n8463) );
  XOR U9191 ( .A(n8459), .B(n8458), .Z(n8845) );
  XOR U9192 ( .A(n8461), .B(n8460), .Z(n8846) );
  NAND U9193 ( .A(n8845), .B(n8846), .Z(n8462) );
  NAND U9194 ( .A(n8463), .B(n8462), .Z(n8467) );
  NAND U9195 ( .A(n8467), .B(n8466), .Z(n8469) );
  XNOR U9196 ( .A(n8467), .B(n8466), .Z(n8852) );
  NAND U9197 ( .A(a[31]), .B(b[35]), .Z(n8851) );
  OR U9198 ( .A(n8852), .B(n8851), .Z(n8468) );
  NAND U9199 ( .A(n8469), .B(n8468), .Z(n8473) );
  NANDN U9200 ( .A(n8472), .B(n8473), .Z(n8475) );
  XNOR U9201 ( .A(n8471), .B(n8470), .Z(n8858) );
  XNOR U9202 ( .A(n8473), .B(n8472), .Z(n8857) );
  NANDN U9203 ( .A(n8858), .B(n8857), .Z(n8474) );
  NAND U9204 ( .A(n8475), .B(n8474), .Z(n8479) );
  NAND U9205 ( .A(n8479), .B(n8478), .Z(n8481) );
  XNOR U9206 ( .A(n8479), .B(n8478), .Z(n8864) );
  NAND U9207 ( .A(a[33]), .B(b[35]), .Z(n8863) );
  OR U9208 ( .A(n8864), .B(n8863), .Z(n8480) );
  NAND U9209 ( .A(n8481), .B(n8480), .Z(n8485) );
  NANDN U9210 ( .A(n8484), .B(n8485), .Z(n8487) );
  XNOR U9211 ( .A(n8483), .B(n8482), .Z(n8870) );
  XNOR U9212 ( .A(n8485), .B(n8484), .Z(n8869) );
  NANDN U9213 ( .A(n8870), .B(n8869), .Z(n8486) );
  NAND U9214 ( .A(n8487), .B(n8486), .Z(n8491) );
  NAND U9215 ( .A(n8491), .B(n8490), .Z(n8493) );
  XNOR U9216 ( .A(n8491), .B(n8490), .Z(n8876) );
  NAND U9217 ( .A(a[35]), .B(b[35]), .Z(n8875) );
  OR U9218 ( .A(n8876), .B(n8875), .Z(n8492) );
  NAND U9219 ( .A(n8493), .B(n8492), .Z(n8497) );
  NANDN U9220 ( .A(n8496), .B(n8497), .Z(n8499) );
  XNOR U9221 ( .A(n8495), .B(n8494), .Z(n8882) );
  XNOR U9222 ( .A(n8497), .B(n8496), .Z(n8881) );
  NANDN U9223 ( .A(n8882), .B(n8881), .Z(n8498) );
  NAND U9224 ( .A(n8499), .B(n8498), .Z(n8503) );
  NAND U9225 ( .A(n8503), .B(n8502), .Z(n8505) );
  XNOR U9226 ( .A(n8503), .B(n8502), .Z(n8888) );
  NAND U9227 ( .A(a[37]), .B(b[35]), .Z(n8887) );
  OR U9228 ( .A(n8888), .B(n8887), .Z(n8504) );
  NAND U9229 ( .A(n8505), .B(n8504), .Z(n8509) );
  NANDN U9230 ( .A(n8508), .B(n8509), .Z(n8511) );
  XNOR U9231 ( .A(n8507), .B(n8506), .Z(n8894) );
  XNOR U9232 ( .A(n8509), .B(n8508), .Z(n8893) );
  NANDN U9233 ( .A(n8894), .B(n8893), .Z(n8510) );
  NAND U9234 ( .A(n8511), .B(n8510), .Z(n8514) );
  AND U9235 ( .A(b[35]), .B(a[39]), .Z(n8515) );
  OR U9236 ( .A(n8514), .B(n8515), .Z(n8517) );
  XOR U9237 ( .A(n8515), .B(n8514), .Z(n8899) );
  NANDN U9238 ( .A(n8900), .B(n8899), .Z(n8516) );
  NAND U9239 ( .A(n8517), .B(n8516), .Z(n8521) );
  NAND U9240 ( .A(a[40]), .B(b[35]), .Z(n8520) );
  OR U9241 ( .A(n8521), .B(n8520), .Z(n8523) );
  XNOR U9242 ( .A(n8519), .B(n8518), .Z(n8906) );
  XOR U9243 ( .A(n8521), .B(n8520), .Z(n8905) );
  NANDN U9244 ( .A(n8906), .B(n8905), .Z(n8522) );
  NAND U9245 ( .A(n8523), .B(n8522), .Z(n8527) );
  NANDN U9246 ( .A(n8526), .B(n8527), .Z(n8529) );
  XNOR U9247 ( .A(n8527), .B(n8526), .Z(n8912) );
  NAND U9248 ( .A(n8911), .B(n8912), .Z(n8528) );
  NAND U9249 ( .A(n8529), .B(n8528), .Z(n8533) );
  NANDN U9250 ( .A(n8532), .B(n8533), .Z(n8535) );
  XNOR U9251 ( .A(n8531), .B(n8530), .Z(n8918) );
  XNOR U9252 ( .A(n8533), .B(n8532), .Z(n8917) );
  NANDN U9253 ( .A(n8918), .B(n8917), .Z(n8534) );
  NAND U9254 ( .A(n8535), .B(n8534), .Z(n8538) );
  AND U9255 ( .A(b[35]), .B(a[43]), .Z(n8539) );
  OR U9256 ( .A(n8538), .B(n8539), .Z(n8541) );
  XOR U9257 ( .A(n8539), .B(n8538), .Z(n8923) );
  NANDN U9258 ( .A(n8924), .B(n8923), .Z(n8540) );
  NAND U9259 ( .A(n8541), .B(n8540), .Z(n8545) );
  NAND U9260 ( .A(a[44]), .B(b[35]), .Z(n8544) );
  OR U9261 ( .A(n8545), .B(n8544), .Z(n8547) );
  XNOR U9262 ( .A(n8543), .B(n8542), .Z(n8930) );
  XOR U9263 ( .A(n8545), .B(n8544), .Z(n8929) );
  NANDN U9264 ( .A(n8930), .B(n8929), .Z(n8546) );
  NAND U9265 ( .A(n8547), .B(n8546), .Z(n8551) );
  NANDN U9266 ( .A(n8550), .B(n8551), .Z(n8553) );
  XNOR U9267 ( .A(n8551), .B(n8550), .Z(n8938) );
  NAND U9268 ( .A(n8937), .B(n8938), .Z(n8552) );
  NAND U9269 ( .A(n8553), .B(n8552), .Z(n8557) );
  NANDN U9270 ( .A(n8556), .B(n8557), .Z(n8559) );
  XNOR U9271 ( .A(n8555), .B(n8554), .Z(n8942) );
  XNOR U9272 ( .A(n8557), .B(n8556), .Z(n8941) );
  NANDN U9273 ( .A(n8942), .B(n8941), .Z(n8558) );
  NAND U9274 ( .A(n8559), .B(n8558), .Z(n8562) );
  AND U9275 ( .A(b[35]), .B(a[47]), .Z(n8563) );
  OR U9276 ( .A(n8562), .B(n8563), .Z(n8565) );
  XOR U9277 ( .A(n8563), .B(n8562), .Z(n8947) );
  NANDN U9278 ( .A(n8948), .B(n8947), .Z(n8564) );
  NAND U9279 ( .A(n8565), .B(n8564), .Z(n8569) );
  NAND U9280 ( .A(a[48]), .B(b[35]), .Z(n8568) );
  OR U9281 ( .A(n8569), .B(n8568), .Z(n8571) );
  XNOR U9282 ( .A(n8567), .B(n8566), .Z(n8954) );
  XOR U9283 ( .A(n8569), .B(n8568), .Z(n8953) );
  NANDN U9284 ( .A(n8954), .B(n8953), .Z(n8570) );
  NAND U9285 ( .A(n8571), .B(n8570), .Z(n8574) );
  AND U9286 ( .A(b[35]), .B(a[49]), .Z(n8575) );
  OR U9287 ( .A(n8574), .B(n8575), .Z(n8577) );
  XOR U9288 ( .A(n8575), .B(n8574), .Z(n8959) );
  NANDN U9289 ( .A(n8960), .B(n8959), .Z(n8576) );
  NAND U9290 ( .A(n8577), .B(n8576), .Z(n8581) );
  NAND U9291 ( .A(a[50]), .B(b[35]), .Z(n8580) );
  OR U9292 ( .A(n8581), .B(n8580), .Z(n8583) );
  XNOR U9293 ( .A(n8579), .B(n8578), .Z(n8966) );
  XOR U9294 ( .A(n8581), .B(n8580), .Z(n8965) );
  NANDN U9295 ( .A(n8966), .B(n8965), .Z(n8582) );
  NAND U9296 ( .A(n8583), .B(n8582), .Z(n8586) );
  AND U9297 ( .A(b[35]), .B(a[51]), .Z(n8587) );
  OR U9298 ( .A(n8586), .B(n8587), .Z(n8589) );
  XOR U9299 ( .A(n8587), .B(n8586), .Z(n8971) );
  NANDN U9300 ( .A(n8972), .B(n8971), .Z(n8588) );
  NAND U9301 ( .A(n8589), .B(n8588), .Z(n8593) );
  NAND U9302 ( .A(a[52]), .B(b[35]), .Z(n8592) );
  OR U9303 ( .A(n8593), .B(n8592), .Z(n8595) );
  XNOR U9304 ( .A(n8591), .B(n8590), .Z(n8978) );
  XOR U9305 ( .A(n8593), .B(n8592), .Z(n8977) );
  NANDN U9306 ( .A(n8978), .B(n8977), .Z(n8594) );
  NAND U9307 ( .A(n8595), .B(n8594), .Z(n8599) );
  NANDN U9308 ( .A(n8598), .B(n8599), .Z(n8601) );
  XNOR U9309 ( .A(n8599), .B(n8598), .Z(n8986) );
  NAND U9310 ( .A(n8985), .B(n8986), .Z(n8600) );
  NAND U9311 ( .A(n8601), .B(n8600), .Z(n8605) );
  NANDN U9312 ( .A(n8604), .B(n8605), .Z(n8607) );
  XNOR U9313 ( .A(n8603), .B(n8602), .Z(n8990) );
  XNOR U9314 ( .A(n8605), .B(n8604), .Z(n8989) );
  NANDN U9315 ( .A(n8990), .B(n8989), .Z(n8606) );
  NAND U9316 ( .A(n8607), .B(n8606), .Z(n8610) );
  AND U9317 ( .A(b[35]), .B(a[55]), .Z(n8611) );
  OR U9318 ( .A(n8610), .B(n8611), .Z(n8613) );
  XOR U9319 ( .A(n8611), .B(n8610), .Z(n8995) );
  NANDN U9320 ( .A(n8996), .B(n8995), .Z(n8612) );
  NAND U9321 ( .A(n8613), .B(n8612), .Z(n8617) );
  NAND U9322 ( .A(a[56]), .B(b[35]), .Z(n8616) );
  OR U9323 ( .A(n8617), .B(n8616), .Z(n8619) );
  XNOR U9324 ( .A(n8615), .B(n8614), .Z(n9002) );
  XOR U9325 ( .A(n8617), .B(n8616), .Z(n9001) );
  NANDN U9326 ( .A(n9002), .B(n9001), .Z(n8618) );
  NAND U9327 ( .A(n8619), .B(n8618), .Z(n8622) );
  AND U9328 ( .A(b[35]), .B(a[57]), .Z(n8623) );
  OR U9329 ( .A(n8622), .B(n8623), .Z(n8625) );
  XOR U9330 ( .A(n8623), .B(n8622), .Z(n9007) );
  NANDN U9331 ( .A(n9008), .B(n9007), .Z(n8624) );
  NAND U9332 ( .A(n8625), .B(n8624), .Z(n8629) );
  NAND U9333 ( .A(a[58]), .B(b[35]), .Z(n8628) );
  OR U9334 ( .A(n8629), .B(n8628), .Z(n8631) );
  XNOR U9335 ( .A(n8627), .B(n8626), .Z(n9014) );
  XOR U9336 ( .A(n8629), .B(n8628), .Z(n9013) );
  NANDN U9337 ( .A(n9014), .B(n9013), .Z(n8630) );
  NAND U9338 ( .A(n8631), .B(n8630), .Z(n8634) );
  AND U9339 ( .A(b[35]), .B(a[59]), .Z(n8635) );
  OR U9340 ( .A(n8634), .B(n8635), .Z(n8637) );
  XOR U9341 ( .A(n8635), .B(n8634), .Z(n9019) );
  NANDN U9342 ( .A(n9020), .B(n9019), .Z(n8636) );
  NAND U9343 ( .A(n8637), .B(n8636), .Z(n8641) );
  NAND U9344 ( .A(a[60]), .B(b[35]), .Z(n8640) );
  OR U9345 ( .A(n8641), .B(n8640), .Z(n8643) );
  XNOR U9346 ( .A(n8639), .B(n8638), .Z(n9026) );
  XOR U9347 ( .A(n8641), .B(n8640), .Z(n9025) );
  NANDN U9348 ( .A(n9026), .B(n9025), .Z(n8642) );
  NAND U9349 ( .A(n8643), .B(n8642), .Z(n8646) );
  AND U9350 ( .A(b[35]), .B(a[61]), .Z(n8647) );
  OR U9351 ( .A(n8646), .B(n8647), .Z(n8649) );
  XOR U9352 ( .A(n8647), .B(n8646), .Z(n9031) );
  NANDN U9353 ( .A(n9032), .B(n9031), .Z(n8648) );
  NAND U9354 ( .A(n8649), .B(n8648), .Z(n8653) );
  NAND U9355 ( .A(a[62]), .B(b[35]), .Z(n8652) );
  OR U9356 ( .A(n8653), .B(n8652), .Z(n8655) );
  XNOR U9357 ( .A(n8651), .B(n8650), .Z(n9038) );
  XOR U9358 ( .A(n8653), .B(n8652), .Z(n9037) );
  NANDN U9359 ( .A(n9038), .B(n9037), .Z(n8654) );
  NAND U9360 ( .A(n8655), .B(n8654), .Z(n8659) );
  NANDN U9361 ( .A(n8658), .B(n8659), .Z(n8661) );
  XNOR U9362 ( .A(n8659), .B(n8658), .Z(n9044) );
  NAND U9363 ( .A(n9043), .B(n9044), .Z(n8660) );
  NAND U9364 ( .A(n8661), .B(n8660), .Z(n8666) );
  NANDN U9365 ( .A(n8667), .B(n8666), .Z(n8665) );
  XOR U9366 ( .A(n8663), .B(n8662), .Z(n8664) );
  NAND U9367 ( .A(n8665), .B(n8664), .Z(n22001) );
  XNOR U9368 ( .A(n8665), .B(n8664), .Z(n24209) );
  XNOR U9369 ( .A(n8667), .B(n8666), .Z(n21998) );
  NAND U9370 ( .A(a[32]), .B(b[34]), .Z(n8853) );
  ANDN U9371 ( .B(b[34]), .A(n21692), .Z(n8797) );
  NAND U9372 ( .A(a[21]), .B(b[34]), .Z(n8786) );
  ANDN U9373 ( .B(b[34]), .A(n172), .Z(n8751) );
  ANDN U9374 ( .B(b[34]), .A(n21615), .Z(n8713) );
  ANDN U9375 ( .B(b[34]), .A(n166), .Z(n8703) );
  ANDN U9376 ( .B(b[34]), .A(n21580), .Z(n8677) );
  NAND U9377 ( .A(b[35]), .B(a[1]), .Z(n8672) );
  NANDN U9378 ( .A(n8672), .B(a[0]), .Z(n8668) );
  XNOR U9379 ( .A(a[2]), .B(n8668), .Z(n8669) );
  NAND U9380 ( .A(b[34]), .B(n8669), .Z(n9060) );
  AND U9381 ( .A(a[1]), .B(b[35]), .Z(n8670) );
  XOR U9382 ( .A(n8671), .B(n8670), .Z(n9061) );
  OR U9383 ( .A(n9060), .B(n9061), .Z(n8676) );
  AND U9384 ( .A(b[34]), .B(a[0]), .Z(n9429) );
  NANDN U9385 ( .A(n8672), .B(n9429), .Z(n8674) );
  NAND U9386 ( .A(a[2]), .B(b[34]), .Z(n8673) );
  AND U9387 ( .A(n8674), .B(n8673), .Z(n8675) );
  ANDN U9388 ( .B(n8676), .A(n8675), .Z(n8678) );
  OR U9389 ( .A(n8677), .B(n8678), .Z(n8682) );
  XNOR U9390 ( .A(n8678), .B(n8677), .Z(n9065) );
  XNOR U9391 ( .A(n8680), .B(n8679), .Z(n9064) );
  OR U9392 ( .A(n9065), .B(n9064), .Z(n8681) );
  NAND U9393 ( .A(n8682), .B(n8681), .Z(n8685) );
  XOR U9394 ( .A(n8684), .B(n8683), .Z(n8686) );
  OR U9395 ( .A(n8685), .B(n8686), .Z(n8688) );
  NAND U9396 ( .A(a[4]), .B(b[34]), .Z(n9073) );
  XOR U9397 ( .A(n8686), .B(n8685), .Z(n9072) );
  NANDN U9398 ( .A(n9073), .B(n9072), .Z(n8687) );
  NAND U9399 ( .A(n8688), .B(n8687), .Z(n8689) );
  ANDN U9400 ( .B(b[34]), .A(n164), .Z(n8690) );
  OR U9401 ( .A(n8689), .B(n8690), .Z(n8694) );
  XNOR U9402 ( .A(n8690), .B(n8689), .Z(n9076) );
  OR U9403 ( .A(n9076), .B(n9077), .Z(n8693) );
  AND U9404 ( .A(n8694), .B(n8693), .Z(n8697) );
  XOR U9405 ( .A(n8696), .B(n8695), .Z(n8698) );
  OR U9406 ( .A(n8697), .B(n8698), .Z(n8700) );
  ANDN U9407 ( .B(b[34]), .A(n165), .Z(n9085) );
  XOR U9408 ( .A(n8698), .B(n8697), .Z(n9084) );
  NANDN U9409 ( .A(n9085), .B(n9084), .Z(n8699) );
  AND U9410 ( .A(n8700), .B(n8699), .Z(n8704) );
  OR U9411 ( .A(n8703), .B(n8704), .Z(n8706) );
  XOR U9412 ( .A(n8704), .B(n8703), .Z(n9088) );
  NANDN U9413 ( .A(n9089), .B(n9088), .Z(n8705) );
  AND U9414 ( .A(n8706), .B(n8705), .Z(n8709) );
  XOR U9415 ( .A(n8708), .B(n8707), .Z(n8710) );
  OR U9416 ( .A(n8709), .B(n8710), .Z(n8712) );
  ANDN U9417 ( .B(b[34]), .A(n167), .Z(n9097) );
  XOR U9418 ( .A(n8710), .B(n8709), .Z(n9096) );
  NANDN U9419 ( .A(n9097), .B(n9096), .Z(n8711) );
  AND U9420 ( .A(n8712), .B(n8711), .Z(n8714) );
  OR U9421 ( .A(n8713), .B(n8714), .Z(n8718) );
  XNOR U9422 ( .A(n8714), .B(n8713), .Z(n9101) );
  XNOR U9423 ( .A(n8716), .B(n8715), .Z(n9100) );
  OR U9424 ( .A(n9101), .B(n9100), .Z(n8717) );
  NAND U9425 ( .A(n8718), .B(n8717), .Z(n8721) );
  XOR U9426 ( .A(n8720), .B(n8719), .Z(n8722) );
  OR U9427 ( .A(n8721), .B(n8722), .Z(n8724) );
  NAND U9428 ( .A(a[10]), .B(b[34]), .Z(n9107) );
  XOR U9429 ( .A(n8722), .B(n8721), .Z(n9106) );
  NANDN U9430 ( .A(n9107), .B(n9106), .Z(n8723) );
  NAND U9431 ( .A(n8724), .B(n8723), .Z(n8725) );
  ANDN U9432 ( .B(b[34]), .A(n21164), .Z(n8726) );
  OR U9433 ( .A(n8725), .B(n8726), .Z(n8730) );
  XNOR U9434 ( .A(n8726), .B(n8725), .Z(n9112) );
  OR U9435 ( .A(n9112), .B(n9113), .Z(n8729) );
  NAND U9436 ( .A(n8730), .B(n8729), .Z(n8733) );
  XNOR U9437 ( .A(n8732), .B(n8731), .Z(n8734) );
  OR U9438 ( .A(n8733), .B(n8734), .Z(n8736) );
  XNOR U9439 ( .A(n8734), .B(n8733), .Z(n9121) );
  AND U9440 ( .A(b[34]), .B(a[12]), .Z(n9120) );
  NANDN U9441 ( .A(n9121), .B(n9120), .Z(n8735) );
  NAND U9442 ( .A(n8736), .B(n8735), .Z(n8739) );
  ANDN U9443 ( .B(b[34]), .A(n170), .Z(n8740) );
  OR U9444 ( .A(n8739), .B(n8740), .Z(n8742) );
  XOR U9445 ( .A(n8738), .B(n8737), .Z(n9125) );
  XOR U9446 ( .A(n8740), .B(n8739), .Z(n9124) );
  NANDN U9447 ( .A(n9125), .B(n9124), .Z(n8741) );
  AND U9448 ( .A(n8742), .B(n8741), .Z(n8745) );
  XOR U9449 ( .A(n8744), .B(n8743), .Z(n8746) );
  OR U9450 ( .A(n8745), .B(n8746), .Z(n8748) );
  ANDN U9451 ( .B(b[34]), .A(n171), .Z(n9133) );
  XOR U9452 ( .A(n8746), .B(n8745), .Z(n9132) );
  NANDN U9453 ( .A(n9133), .B(n9132), .Z(n8747) );
  AND U9454 ( .A(n8748), .B(n8747), .Z(n8752) );
  OR U9455 ( .A(n8751), .B(n8752), .Z(n8754) );
  XOR U9456 ( .A(n8752), .B(n8751), .Z(n9136) );
  NANDN U9457 ( .A(n9137), .B(n9136), .Z(n8753) );
  NAND U9458 ( .A(n8754), .B(n8753), .Z(n8757) );
  XOR U9459 ( .A(n8756), .B(n8755), .Z(n8758) );
  OR U9460 ( .A(n8757), .B(n8758), .Z(n8760) );
  NAND U9461 ( .A(a[16]), .B(b[34]), .Z(n9143) );
  XOR U9462 ( .A(n8758), .B(n8757), .Z(n9142) );
  NANDN U9463 ( .A(n9143), .B(n9142), .Z(n8759) );
  NAND U9464 ( .A(n8760), .B(n8759), .Z(n8761) );
  ANDN U9465 ( .B(b[34]), .A(n174), .Z(n8762) );
  OR U9466 ( .A(n8761), .B(n8762), .Z(n8766) );
  XNOR U9467 ( .A(n8762), .B(n8761), .Z(n9149) );
  XNOR U9468 ( .A(n8764), .B(n8763), .Z(n9148) );
  OR U9469 ( .A(n9149), .B(n9148), .Z(n8765) );
  NAND U9470 ( .A(n8766), .B(n8765), .Z(n8769) );
  XNOR U9471 ( .A(n8768), .B(n8767), .Z(n8770) );
  OR U9472 ( .A(n8769), .B(n8770), .Z(n8772) );
  XNOR U9473 ( .A(n8770), .B(n8769), .Z(n9155) );
  NAND U9474 ( .A(a[18]), .B(b[34]), .Z(n9154) );
  OR U9475 ( .A(n9155), .B(n9154), .Z(n8771) );
  NAND U9476 ( .A(n8772), .B(n8771), .Z(n8775) );
  ANDN U9477 ( .B(b[34]), .A(n21670), .Z(n8776) );
  OR U9478 ( .A(n8775), .B(n8776), .Z(n8778) );
  XOR U9479 ( .A(n8774), .B(n8773), .Z(n9161) );
  XOR U9480 ( .A(n8776), .B(n8775), .Z(n9160) );
  NANDN U9481 ( .A(n9161), .B(n9160), .Z(n8777) );
  AND U9482 ( .A(n8778), .B(n8777), .Z(n8782) );
  NANDN U9483 ( .A(n8782), .B(n8781), .Z(n8784) );
  XOR U9484 ( .A(n8782), .B(n8781), .Z(n9168) );
  ANDN U9485 ( .B(b[34]), .A(n176), .Z(n9169) );
  OR U9486 ( .A(n9168), .B(n9169), .Z(n8783) );
  NAND U9487 ( .A(n8784), .B(n8783), .Z(n8785) );
  OR U9488 ( .A(n8786), .B(n8785), .Z(n8790) );
  XNOR U9489 ( .A(n8786), .B(n8785), .Z(n9173) );
  XNOR U9490 ( .A(n8788), .B(n8787), .Z(n9172) );
  NANDN U9491 ( .A(n9173), .B(n9172), .Z(n8789) );
  NAND U9492 ( .A(n8790), .B(n8789), .Z(n8793) );
  XOR U9493 ( .A(n8792), .B(n8791), .Z(n8794) );
  NANDN U9494 ( .A(n8793), .B(n8794), .Z(n8796) );
  XOR U9495 ( .A(n8794), .B(n8793), .Z(n9180) );
  ANDN U9496 ( .B(b[34]), .A(n177), .Z(n9181) );
  OR U9497 ( .A(n9180), .B(n9181), .Z(n8795) );
  AND U9498 ( .A(n8796), .B(n8795), .Z(n8798) );
  OR U9499 ( .A(n8797), .B(n8798), .Z(n8802) );
  XNOR U9500 ( .A(n8798), .B(n8797), .Z(n9184) );
  XOR U9501 ( .A(n8800), .B(n8799), .Z(n9185) );
  OR U9502 ( .A(n9184), .B(n9185), .Z(n8801) );
  NAND U9503 ( .A(n8802), .B(n8801), .Z(n8805) );
  XOR U9504 ( .A(n8804), .B(n8803), .Z(n8806) );
  OR U9505 ( .A(n8805), .B(n8806), .Z(n8808) );
  NAND U9506 ( .A(a[24]), .B(b[34]), .Z(n9191) );
  XOR U9507 ( .A(n8806), .B(n8805), .Z(n9190) );
  NANDN U9508 ( .A(n9191), .B(n9190), .Z(n8807) );
  NAND U9509 ( .A(n8808), .B(n8807), .Z(n8809) );
  ANDN U9510 ( .B(b[34]), .A(n21703), .Z(n8810) );
  OR U9511 ( .A(n8809), .B(n8810), .Z(n8814) );
  XNOR U9512 ( .A(n8810), .B(n8809), .Z(n9197) );
  XOR U9513 ( .A(n8812), .B(n8811), .Z(n9196) );
  OR U9514 ( .A(n9197), .B(n9196), .Z(n8813) );
  NAND U9515 ( .A(n8814), .B(n8813), .Z(n8817) );
  XNOR U9516 ( .A(n8816), .B(n8815), .Z(n8818) );
  OR U9517 ( .A(n8817), .B(n8818), .Z(n8820) );
  XNOR U9518 ( .A(n8818), .B(n8817), .Z(n9203) );
  NAND U9519 ( .A(a[26]), .B(b[34]), .Z(n9202) );
  OR U9520 ( .A(n9203), .B(n9202), .Z(n8819) );
  NAND U9521 ( .A(n8820), .B(n8819), .Z(n8821) );
  ANDN U9522 ( .B(b[34]), .A(n21716), .Z(n8822) );
  OR U9523 ( .A(n8821), .B(n8822), .Z(n8826) );
  XNOR U9524 ( .A(n8822), .B(n8821), .Z(n9209) );
  OR U9525 ( .A(n9209), .B(n9208), .Z(n8825) );
  NAND U9526 ( .A(n8826), .B(n8825), .Z(n8829) );
  XNOR U9527 ( .A(n8828), .B(n8827), .Z(n8830) );
  OR U9528 ( .A(n8829), .B(n8830), .Z(n8832) );
  XNOR U9529 ( .A(n8830), .B(n8829), .Z(n9215) );
  NAND U9530 ( .A(a[28]), .B(b[34]), .Z(n9214) );
  OR U9531 ( .A(n9215), .B(n9214), .Z(n8831) );
  NAND U9532 ( .A(n8832), .B(n8831), .Z(n8833) );
  ANDN U9533 ( .B(b[34]), .A(n21727), .Z(n8834) );
  OR U9534 ( .A(n8833), .B(n8834), .Z(n8838) );
  XNOR U9535 ( .A(n8834), .B(n8833), .Z(n9221) );
  XOR U9536 ( .A(n8836), .B(n8835), .Z(n9220) );
  OR U9537 ( .A(n9221), .B(n9220), .Z(n8837) );
  NAND U9538 ( .A(n8838), .B(n8837), .Z(n8842) );
  AND U9539 ( .A(b[34]), .B(a[30]), .Z(n8841) );
  NANDN U9540 ( .A(n8842), .B(n8841), .Z(n8844) );
  XNOR U9541 ( .A(n8842), .B(n8841), .Z(n9228) );
  NANDN U9542 ( .A(n9229), .B(n9228), .Z(n8843) );
  NAND U9543 ( .A(n8844), .B(n8843), .Z(n8848) );
  XOR U9544 ( .A(n8846), .B(n8845), .Z(n8847) );
  NAND U9545 ( .A(n8848), .B(n8847), .Z(n8850) );
  XNOR U9546 ( .A(n8848), .B(n8847), .Z(n9233) );
  NAND U9547 ( .A(a[31]), .B(b[34]), .Z(n9232) );
  OR U9548 ( .A(n9233), .B(n9232), .Z(n8849) );
  NAND U9549 ( .A(n8850), .B(n8849), .Z(n8854) );
  NANDN U9550 ( .A(n8853), .B(n8854), .Z(n8856) );
  XOR U9551 ( .A(n8852), .B(n8851), .Z(n9238) );
  XNOR U9552 ( .A(n8854), .B(n8853), .Z(n9239) );
  NAND U9553 ( .A(n9238), .B(n9239), .Z(n8855) );
  NAND U9554 ( .A(n8856), .B(n8855), .Z(n8859) );
  AND U9555 ( .A(b[34]), .B(a[33]), .Z(n8860) );
  OR U9556 ( .A(n8859), .B(n8860), .Z(n8862) );
  XNOR U9557 ( .A(n8858), .B(n8857), .Z(n9245) );
  XOR U9558 ( .A(n8860), .B(n8859), .Z(n9244) );
  NANDN U9559 ( .A(n9245), .B(n9244), .Z(n8861) );
  NAND U9560 ( .A(n8862), .B(n8861), .Z(n8866) );
  NAND U9561 ( .A(a[34]), .B(b[34]), .Z(n8865) );
  OR U9562 ( .A(n8866), .B(n8865), .Z(n8868) );
  XOR U9563 ( .A(n8864), .B(n8863), .Z(n9250) );
  XOR U9564 ( .A(n8866), .B(n8865), .Z(n9251) );
  NAND U9565 ( .A(n9250), .B(n9251), .Z(n8867) );
  NAND U9566 ( .A(n8868), .B(n8867), .Z(n8871) );
  AND U9567 ( .A(b[34]), .B(a[35]), .Z(n8872) );
  OR U9568 ( .A(n8871), .B(n8872), .Z(n8874) );
  XNOR U9569 ( .A(n8870), .B(n8869), .Z(n9257) );
  XOR U9570 ( .A(n8872), .B(n8871), .Z(n9256) );
  NANDN U9571 ( .A(n9257), .B(n9256), .Z(n8873) );
  NAND U9572 ( .A(n8874), .B(n8873), .Z(n8878) );
  NAND U9573 ( .A(a[36]), .B(b[34]), .Z(n8877) );
  OR U9574 ( .A(n8878), .B(n8877), .Z(n8880) );
  XOR U9575 ( .A(n8876), .B(n8875), .Z(n9262) );
  XOR U9576 ( .A(n8878), .B(n8877), .Z(n9263) );
  NAND U9577 ( .A(n9262), .B(n9263), .Z(n8879) );
  NAND U9578 ( .A(n8880), .B(n8879), .Z(n8883) );
  AND U9579 ( .A(b[34]), .B(a[37]), .Z(n8884) );
  OR U9580 ( .A(n8883), .B(n8884), .Z(n8886) );
  XNOR U9581 ( .A(n8882), .B(n8881), .Z(n9269) );
  XOR U9582 ( .A(n8884), .B(n8883), .Z(n9268) );
  NANDN U9583 ( .A(n9269), .B(n9268), .Z(n8885) );
  NAND U9584 ( .A(n8886), .B(n8885), .Z(n8890) );
  NAND U9585 ( .A(a[38]), .B(b[34]), .Z(n8889) );
  OR U9586 ( .A(n8890), .B(n8889), .Z(n8892) );
  XOR U9587 ( .A(n8888), .B(n8887), .Z(n9274) );
  XOR U9588 ( .A(n8890), .B(n8889), .Z(n9275) );
  NAND U9589 ( .A(n9274), .B(n9275), .Z(n8891) );
  NAND U9590 ( .A(n8892), .B(n8891), .Z(n8895) );
  AND U9591 ( .A(b[34]), .B(a[39]), .Z(n8896) );
  OR U9592 ( .A(n8895), .B(n8896), .Z(n8898) );
  XNOR U9593 ( .A(n8894), .B(n8893), .Z(n9281) );
  XOR U9594 ( .A(n8896), .B(n8895), .Z(n9280) );
  NANDN U9595 ( .A(n9281), .B(n9280), .Z(n8897) );
  NAND U9596 ( .A(n8898), .B(n8897), .Z(n8902) );
  NAND U9597 ( .A(a[40]), .B(b[34]), .Z(n8901) );
  OR U9598 ( .A(n8902), .B(n8901), .Z(n8904) );
  XOR U9599 ( .A(n8900), .B(n8899), .Z(n9287) );
  XOR U9600 ( .A(n8902), .B(n8901), .Z(n9286) );
  NAND U9601 ( .A(n9287), .B(n9286), .Z(n8903) );
  NAND U9602 ( .A(n8904), .B(n8903), .Z(n8907) );
  AND U9603 ( .A(b[34]), .B(a[41]), .Z(n8908) );
  OR U9604 ( .A(n8907), .B(n8908), .Z(n8910) );
  XNOR U9605 ( .A(n8906), .B(n8905), .Z(n9293) );
  XOR U9606 ( .A(n8908), .B(n8907), .Z(n9292) );
  NANDN U9607 ( .A(n9293), .B(n9292), .Z(n8909) );
  NAND U9608 ( .A(n8910), .B(n8909), .Z(n8914) );
  NAND U9609 ( .A(a[42]), .B(b[34]), .Z(n8913) );
  OR U9610 ( .A(n8914), .B(n8913), .Z(n8916) );
  XOR U9611 ( .A(n8912), .B(n8911), .Z(n9298) );
  XOR U9612 ( .A(n8914), .B(n8913), .Z(n9299) );
  NAND U9613 ( .A(n9298), .B(n9299), .Z(n8915) );
  NAND U9614 ( .A(n8916), .B(n8915), .Z(n8919) );
  AND U9615 ( .A(b[34]), .B(a[43]), .Z(n8920) );
  OR U9616 ( .A(n8919), .B(n8920), .Z(n8922) );
  XNOR U9617 ( .A(n8918), .B(n8917), .Z(n9305) );
  XOR U9618 ( .A(n8920), .B(n8919), .Z(n9304) );
  NANDN U9619 ( .A(n9305), .B(n9304), .Z(n8921) );
  NAND U9620 ( .A(n8922), .B(n8921), .Z(n8926) );
  NAND U9621 ( .A(a[44]), .B(b[34]), .Z(n8925) );
  OR U9622 ( .A(n8926), .B(n8925), .Z(n8928) );
  XOR U9623 ( .A(n8924), .B(n8923), .Z(n9311) );
  XOR U9624 ( .A(n8926), .B(n8925), .Z(n9310) );
  NAND U9625 ( .A(n9311), .B(n9310), .Z(n8927) );
  NAND U9626 ( .A(n8928), .B(n8927), .Z(n8931) );
  AND U9627 ( .A(b[34]), .B(a[45]), .Z(n8932) );
  OR U9628 ( .A(n8931), .B(n8932), .Z(n8934) );
  XNOR U9629 ( .A(n8930), .B(n8929), .Z(n9317) );
  XOR U9630 ( .A(n8932), .B(n8931), .Z(n9316) );
  NANDN U9631 ( .A(n9317), .B(n9316), .Z(n8933) );
  NAND U9632 ( .A(n8934), .B(n8933), .Z(n8936) );
  NAND U9633 ( .A(a[46]), .B(b[34]), .Z(n8935) );
  OR U9634 ( .A(n8936), .B(n8935), .Z(n8940) );
  XOR U9635 ( .A(n8936), .B(n8935), .Z(n9322) );
  XOR U9636 ( .A(n8938), .B(n8937), .Z(n9323) );
  NAND U9637 ( .A(n9322), .B(n9323), .Z(n8939) );
  NAND U9638 ( .A(n8940), .B(n8939), .Z(n8943) );
  AND U9639 ( .A(b[34]), .B(a[47]), .Z(n8944) );
  OR U9640 ( .A(n8943), .B(n8944), .Z(n8946) );
  XNOR U9641 ( .A(n8942), .B(n8941), .Z(n9329) );
  XOR U9642 ( .A(n8944), .B(n8943), .Z(n9328) );
  NANDN U9643 ( .A(n9329), .B(n9328), .Z(n8945) );
  NAND U9644 ( .A(n8946), .B(n8945), .Z(n8950) );
  NAND U9645 ( .A(a[48]), .B(b[34]), .Z(n8949) );
  OR U9646 ( .A(n8950), .B(n8949), .Z(n8952) );
  XOR U9647 ( .A(n8948), .B(n8947), .Z(n9335) );
  XOR U9648 ( .A(n8950), .B(n8949), .Z(n9334) );
  NAND U9649 ( .A(n9335), .B(n9334), .Z(n8951) );
  NAND U9650 ( .A(n8952), .B(n8951), .Z(n8955) );
  AND U9651 ( .A(b[34]), .B(a[49]), .Z(n8956) );
  OR U9652 ( .A(n8955), .B(n8956), .Z(n8958) );
  XNOR U9653 ( .A(n8954), .B(n8953), .Z(n9341) );
  XOR U9654 ( .A(n8956), .B(n8955), .Z(n9340) );
  NANDN U9655 ( .A(n9341), .B(n9340), .Z(n8957) );
  NAND U9656 ( .A(n8958), .B(n8957), .Z(n8962) );
  NAND U9657 ( .A(a[50]), .B(b[34]), .Z(n8961) );
  OR U9658 ( .A(n8962), .B(n8961), .Z(n8964) );
  XOR U9659 ( .A(n8960), .B(n8959), .Z(n9347) );
  XOR U9660 ( .A(n8962), .B(n8961), .Z(n9346) );
  NAND U9661 ( .A(n9347), .B(n9346), .Z(n8963) );
  NAND U9662 ( .A(n8964), .B(n8963), .Z(n8967) );
  AND U9663 ( .A(b[34]), .B(a[51]), .Z(n8968) );
  OR U9664 ( .A(n8967), .B(n8968), .Z(n8970) );
  XNOR U9665 ( .A(n8966), .B(n8965), .Z(n9353) );
  XOR U9666 ( .A(n8968), .B(n8967), .Z(n9352) );
  NANDN U9667 ( .A(n9353), .B(n9352), .Z(n8969) );
  NAND U9668 ( .A(n8970), .B(n8969), .Z(n8974) );
  NAND U9669 ( .A(a[52]), .B(b[34]), .Z(n8973) );
  OR U9670 ( .A(n8974), .B(n8973), .Z(n8976) );
  XOR U9671 ( .A(n8972), .B(n8971), .Z(n9359) );
  XOR U9672 ( .A(n8974), .B(n8973), .Z(n9358) );
  NAND U9673 ( .A(n9359), .B(n9358), .Z(n8975) );
  NAND U9674 ( .A(n8976), .B(n8975), .Z(n8979) );
  AND U9675 ( .A(b[34]), .B(a[53]), .Z(n8980) );
  OR U9676 ( .A(n8979), .B(n8980), .Z(n8982) );
  XNOR U9677 ( .A(n8978), .B(n8977), .Z(n9365) );
  XOR U9678 ( .A(n8980), .B(n8979), .Z(n9364) );
  NANDN U9679 ( .A(n9365), .B(n9364), .Z(n8981) );
  NAND U9680 ( .A(n8982), .B(n8981), .Z(n8984) );
  NAND U9681 ( .A(a[54]), .B(b[34]), .Z(n8983) );
  OR U9682 ( .A(n8984), .B(n8983), .Z(n8988) );
  XOR U9683 ( .A(n8984), .B(n8983), .Z(n9370) );
  XOR U9684 ( .A(n8986), .B(n8985), .Z(n9371) );
  NAND U9685 ( .A(n9370), .B(n9371), .Z(n8987) );
  NAND U9686 ( .A(n8988), .B(n8987), .Z(n8991) );
  AND U9687 ( .A(b[34]), .B(a[55]), .Z(n8992) );
  OR U9688 ( .A(n8991), .B(n8992), .Z(n8994) );
  XNOR U9689 ( .A(n8990), .B(n8989), .Z(n9377) );
  XOR U9690 ( .A(n8992), .B(n8991), .Z(n9376) );
  NANDN U9691 ( .A(n9377), .B(n9376), .Z(n8993) );
  NAND U9692 ( .A(n8994), .B(n8993), .Z(n8998) );
  NAND U9693 ( .A(a[56]), .B(b[34]), .Z(n8997) );
  OR U9694 ( .A(n8998), .B(n8997), .Z(n9000) );
  XOR U9695 ( .A(n8996), .B(n8995), .Z(n9383) );
  XOR U9696 ( .A(n8998), .B(n8997), .Z(n9382) );
  NAND U9697 ( .A(n9383), .B(n9382), .Z(n8999) );
  NAND U9698 ( .A(n9000), .B(n8999), .Z(n9003) );
  AND U9699 ( .A(b[34]), .B(a[57]), .Z(n9004) );
  OR U9700 ( .A(n9003), .B(n9004), .Z(n9006) );
  XNOR U9701 ( .A(n9002), .B(n9001), .Z(n9389) );
  XOR U9702 ( .A(n9004), .B(n9003), .Z(n9388) );
  NANDN U9703 ( .A(n9389), .B(n9388), .Z(n9005) );
  NAND U9704 ( .A(n9006), .B(n9005), .Z(n9010) );
  NAND U9705 ( .A(a[58]), .B(b[34]), .Z(n9009) );
  OR U9706 ( .A(n9010), .B(n9009), .Z(n9012) );
  XOR U9707 ( .A(n9008), .B(n9007), .Z(n9395) );
  XOR U9708 ( .A(n9010), .B(n9009), .Z(n9394) );
  NAND U9709 ( .A(n9395), .B(n9394), .Z(n9011) );
  NAND U9710 ( .A(n9012), .B(n9011), .Z(n9015) );
  AND U9711 ( .A(b[34]), .B(a[59]), .Z(n9016) );
  OR U9712 ( .A(n9015), .B(n9016), .Z(n9018) );
  XNOR U9713 ( .A(n9014), .B(n9013), .Z(n9401) );
  XOR U9714 ( .A(n9016), .B(n9015), .Z(n9400) );
  NANDN U9715 ( .A(n9401), .B(n9400), .Z(n9017) );
  NAND U9716 ( .A(n9018), .B(n9017), .Z(n9022) );
  NAND U9717 ( .A(a[60]), .B(b[34]), .Z(n9021) );
  OR U9718 ( .A(n9022), .B(n9021), .Z(n9024) );
  XOR U9719 ( .A(n9020), .B(n9019), .Z(n9407) );
  XOR U9720 ( .A(n9022), .B(n9021), .Z(n9406) );
  NAND U9721 ( .A(n9407), .B(n9406), .Z(n9023) );
  NAND U9722 ( .A(n9024), .B(n9023), .Z(n9027) );
  AND U9723 ( .A(b[34]), .B(a[61]), .Z(n9028) );
  OR U9724 ( .A(n9027), .B(n9028), .Z(n9030) );
  XNOR U9725 ( .A(n9026), .B(n9025), .Z(n9413) );
  XOR U9726 ( .A(n9028), .B(n9027), .Z(n9412) );
  NANDN U9727 ( .A(n9413), .B(n9412), .Z(n9029) );
  NAND U9728 ( .A(n9030), .B(n9029), .Z(n9034) );
  NAND U9729 ( .A(a[62]), .B(b[34]), .Z(n9033) );
  OR U9730 ( .A(n9034), .B(n9033), .Z(n9036) );
  XOR U9731 ( .A(n9032), .B(n9031), .Z(n9419) );
  XOR U9732 ( .A(n9034), .B(n9033), .Z(n9418) );
  NAND U9733 ( .A(n9419), .B(n9418), .Z(n9035) );
  NAND U9734 ( .A(n9036), .B(n9035), .Z(n9039) );
  AND U9735 ( .A(b[34]), .B(a[63]), .Z(n9040) );
  OR U9736 ( .A(n9039), .B(n9040), .Z(n9042) );
  XNOR U9737 ( .A(n9038), .B(n9037), .Z(n9048) );
  XOR U9738 ( .A(n9040), .B(n9039), .Z(n9047) );
  NANDN U9739 ( .A(n9048), .B(n9047), .Z(n9041) );
  AND U9740 ( .A(n9042), .B(n9041), .Z(n9045) );
  XOR U9741 ( .A(n9044), .B(n9043), .Z(n9046) );
  AND U9742 ( .A(n9045), .B(n9046), .Z(n21999) );
  XNOR U9743 ( .A(n9046), .B(n9045), .Z(n21995) );
  XNOR U9744 ( .A(n9048), .B(n9047), .Z(n9425) );
  NAND U9745 ( .A(a[62]), .B(b[33]), .Z(n9414) );
  NAND U9746 ( .A(a[60]), .B(b[33]), .Z(n9402) );
  NAND U9747 ( .A(a[59]), .B(b[33]), .Z(n9396) );
  NAND U9748 ( .A(a[58]), .B(b[33]), .Z(n9390) );
  NAND U9749 ( .A(a[57]), .B(b[33]), .Z(n9384) );
  NAND U9750 ( .A(a[56]), .B(b[33]), .Z(n9378) );
  NAND U9751 ( .A(a[55]), .B(b[33]), .Z(n9372) );
  NAND U9752 ( .A(a[54]), .B(b[33]), .Z(n9366) );
  NAND U9753 ( .A(a[53]), .B(b[33]), .Z(n9360) );
  NAND U9754 ( .A(a[52]), .B(b[33]), .Z(n9354) );
  NAND U9755 ( .A(a[51]), .B(b[33]), .Z(n9348) );
  NAND U9756 ( .A(a[50]), .B(b[33]), .Z(n9342) );
  NAND U9757 ( .A(a[49]), .B(b[33]), .Z(n9336) );
  NAND U9758 ( .A(a[48]), .B(b[33]), .Z(n9330) );
  NAND U9759 ( .A(a[46]), .B(b[33]), .Z(n9318) );
  NAND U9760 ( .A(a[44]), .B(b[33]), .Z(n9306) );
  NAND U9761 ( .A(a[42]), .B(b[33]), .Z(n9294) );
  NAND U9762 ( .A(a[40]), .B(b[33]), .Z(n9282) );
  NAND U9763 ( .A(a[38]), .B(b[33]), .Z(n9270) );
  NAND U9764 ( .A(a[36]), .B(b[33]), .Z(n9258) );
  NAND U9765 ( .A(a[34]), .B(b[33]), .Z(n9246) );
  ANDN U9766 ( .B(b[33]), .A(n21727), .Z(n9216) );
  ANDN U9767 ( .B(b[33]), .A(n21703), .Z(n9192) );
  ANDN U9768 ( .B(b[33]), .A(n21692), .Z(n9178) );
  NAND U9769 ( .A(a[13]), .B(b[33]), .Z(n9119) );
  ANDN U9770 ( .B(b[33]), .A(n166), .Z(n9082) );
  ANDN U9771 ( .B(b[33]), .A(n21580), .Z(n9058) );
  NAND U9772 ( .A(b[34]), .B(a[1]), .Z(n9053) );
  NANDN U9773 ( .A(n9053), .B(a[0]), .Z(n9049) );
  XNOR U9774 ( .A(a[2]), .B(n9049), .Z(n9050) );
  NAND U9775 ( .A(b[33]), .B(n9050), .Z(n9437) );
  AND U9776 ( .A(a[1]), .B(b[34]), .Z(n9051) );
  XOR U9777 ( .A(n9052), .B(n9051), .Z(n9438) );
  OR U9778 ( .A(n9437), .B(n9438), .Z(n9057) );
  AND U9779 ( .A(b[33]), .B(a[0]), .Z(n9811) );
  NANDN U9780 ( .A(n9053), .B(n9811), .Z(n9055) );
  NAND U9781 ( .A(a[2]), .B(b[33]), .Z(n9054) );
  AND U9782 ( .A(n9055), .B(n9054), .Z(n9056) );
  ANDN U9783 ( .B(n9057), .A(n9056), .Z(n9059) );
  OR U9784 ( .A(n9058), .B(n9059), .Z(n9063) );
  XNOR U9785 ( .A(n9059), .B(n9058), .Z(n9442) );
  XNOR U9786 ( .A(n9061), .B(n9060), .Z(n9441) );
  OR U9787 ( .A(n9442), .B(n9441), .Z(n9062) );
  NAND U9788 ( .A(n9063), .B(n9062), .Z(n9066) );
  XOR U9789 ( .A(n9065), .B(n9064), .Z(n9067) );
  OR U9790 ( .A(n9066), .B(n9067), .Z(n9069) );
  NAND U9791 ( .A(a[4]), .B(b[33]), .Z(n9450) );
  XOR U9792 ( .A(n9067), .B(n9066), .Z(n9449) );
  NANDN U9793 ( .A(n9450), .B(n9449), .Z(n9068) );
  NAND U9794 ( .A(n9069), .B(n9068), .Z(n9070) );
  ANDN U9795 ( .B(b[33]), .A(n164), .Z(n9071) );
  OR U9796 ( .A(n9070), .B(n9071), .Z(n9075) );
  XNOR U9797 ( .A(n9071), .B(n9070), .Z(n9453) );
  OR U9798 ( .A(n9453), .B(n9454), .Z(n9074) );
  AND U9799 ( .A(n9075), .B(n9074), .Z(n9079) );
  XOR U9800 ( .A(n9077), .B(n9076), .Z(n9078) );
  NANDN U9801 ( .A(n9079), .B(n9078), .Z(n9081) );
  XOR U9802 ( .A(n9079), .B(n9078), .Z(n9461) );
  ANDN U9803 ( .B(b[33]), .A(n165), .Z(n9462) );
  OR U9804 ( .A(n9461), .B(n9462), .Z(n9080) );
  AND U9805 ( .A(n9081), .B(n9080), .Z(n9083) );
  OR U9806 ( .A(n9082), .B(n9083), .Z(n9087) );
  XNOR U9807 ( .A(n9083), .B(n9082), .Z(n9466) );
  XOR U9808 ( .A(n9085), .B(n9084), .Z(n9465) );
  OR U9809 ( .A(n9466), .B(n9465), .Z(n9086) );
  NAND U9810 ( .A(n9087), .B(n9086), .Z(n9090) );
  XNOR U9811 ( .A(n9089), .B(n9088), .Z(n9091) );
  OR U9812 ( .A(n9090), .B(n9091), .Z(n9093) );
  XNOR U9813 ( .A(n9091), .B(n9090), .Z(n9472) );
  NAND U9814 ( .A(a[8]), .B(b[33]), .Z(n9471) );
  OR U9815 ( .A(n9472), .B(n9471), .Z(n9092) );
  NAND U9816 ( .A(n9093), .B(n9092), .Z(n9094) );
  ANDN U9817 ( .B(b[33]), .A(n21615), .Z(n9095) );
  OR U9818 ( .A(n9094), .B(n9095), .Z(n9099) );
  XNOR U9819 ( .A(n9095), .B(n9094), .Z(n9478) );
  XOR U9820 ( .A(n9097), .B(n9096), .Z(n9477) );
  OR U9821 ( .A(n9478), .B(n9477), .Z(n9098) );
  NAND U9822 ( .A(n9099), .B(n9098), .Z(n9102) );
  XOR U9823 ( .A(n9101), .B(n9100), .Z(n9103) );
  OR U9824 ( .A(n9102), .B(n9103), .Z(n9105) );
  NAND U9825 ( .A(a[10]), .B(b[33]), .Z(n9484) );
  XOR U9826 ( .A(n9103), .B(n9102), .Z(n9483) );
  NANDN U9827 ( .A(n9484), .B(n9483), .Z(n9104) );
  NAND U9828 ( .A(n9105), .B(n9104), .Z(n9108) );
  ANDN U9829 ( .B(b[33]), .A(n21164), .Z(n9109) );
  OR U9830 ( .A(n9108), .B(n9109), .Z(n9111) );
  XOR U9831 ( .A(n9109), .B(n9108), .Z(n9489) );
  NANDN U9832 ( .A(n9490), .B(n9489), .Z(n9110) );
  AND U9833 ( .A(n9111), .B(n9110), .Z(n9115) );
  XOR U9834 ( .A(n9113), .B(n9112), .Z(n9114) );
  NANDN U9835 ( .A(n9115), .B(n9114), .Z(n9117) );
  XOR U9836 ( .A(n9115), .B(n9114), .Z(n9497) );
  ANDN U9837 ( .B(b[33]), .A(n169), .Z(n9498) );
  OR U9838 ( .A(n9497), .B(n9498), .Z(n9116) );
  NAND U9839 ( .A(n9117), .B(n9116), .Z(n9118) );
  OR U9840 ( .A(n9119), .B(n9118), .Z(n9123) );
  XNOR U9841 ( .A(n9119), .B(n9118), .Z(n9502) );
  XNOR U9842 ( .A(n9121), .B(n9120), .Z(n9501) );
  NANDN U9843 ( .A(n9502), .B(n9501), .Z(n9122) );
  AND U9844 ( .A(n9123), .B(n9122), .Z(n9126) );
  XNOR U9845 ( .A(n9125), .B(n9124), .Z(n9127) );
  OR U9846 ( .A(n9126), .B(n9127), .Z(n9129) );
  XNOR U9847 ( .A(n9127), .B(n9126), .Z(n9508) );
  NAND U9848 ( .A(a[14]), .B(b[33]), .Z(n9507) );
  OR U9849 ( .A(n9508), .B(n9507), .Z(n9128) );
  NAND U9850 ( .A(n9129), .B(n9128), .Z(n9130) );
  ANDN U9851 ( .B(b[33]), .A(n172), .Z(n9131) );
  OR U9852 ( .A(n9130), .B(n9131), .Z(n9135) );
  XNOR U9853 ( .A(n9131), .B(n9130), .Z(n9514) );
  XOR U9854 ( .A(n9133), .B(n9132), .Z(n9513) );
  OR U9855 ( .A(n9514), .B(n9513), .Z(n9134) );
  NAND U9856 ( .A(n9135), .B(n9134), .Z(n9138) );
  XNOR U9857 ( .A(n9137), .B(n9136), .Z(n9139) );
  OR U9858 ( .A(n9138), .B(n9139), .Z(n9141) );
  XNOR U9859 ( .A(n9139), .B(n9138), .Z(n9520) );
  NAND U9860 ( .A(a[16]), .B(b[33]), .Z(n9519) );
  OR U9861 ( .A(n9520), .B(n9519), .Z(n9140) );
  NAND U9862 ( .A(n9141), .B(n9140), .Z(n9144) );
  ANDN U9863 ( .B(b[33]), .A(n174), .Z(n9145) );
  OR U9864 ( .A(n9144), .B(n9145), .Z(n9147) );
  XOR U9865 ( .A(n9145), .B(n9144), .Z(n9525) );
  NANDN U9866 ( .A(n9526), .B(n9525), .Z(n9146) );
  NAND U9867 ( .A(n9147), .B(n9146), .Z(n9150) );
  XOR U9868 ( .A(n9149), .B(n9148), .Z(n9151) );
  OR U9869 ( .A(n9150), .B(n9151), .Z(n9153) );
  NAND U9870 ( .A(a[18]), .B(b[33]), .Z(n9532) );
  XOR U9871 ( .A(n9151), .B(n9150), .Z(n9531) );
  NANDN U9872 ( .A(n9532), .B(n9531), .Z(n9152) );
  NAND U9873 ( .A(n9153), .B(n9152), .Z(n9156) );
  ANDN U9874 ( .B(b[33]), .A(n21670), .Z(n9157) );
  OR U9875 ( .A(n9156), .B(n9157), .Z(n9159) );
  XOR U9876 ( .A(n9155), .B(n9154), .Z(n9538) );
  XOR U9877 ( .A(n9157), .B(n9156), .Z(n9537) );
  NANDN U9878 ( .A(n9538), .B(n9537), .Z(n9158) );
  NAND U9879 ( .A(n9159), .B(n9158), .Z(n9162) );
  XNOR U9880 ( .A(n9161), .B(n9160), .Z(n9163) );
  OR U9881 ( .A(n9162), .B(n9163), .Z(n9165) );
  XNOR U9882 ( .A(n9163), .B(n9162), .Z(n9544) );
  NAND U9883 ( .A(a[20]), .B(b[33]), .Z(n9543) );
  OR U9884 ( .A(n9544), .B(n9543), .Z(n9164) );
  NAND U9885 ( .A(n9165), .B(n9164), .Z(n9166) );
  ANDN U9886 ( .B(b[33]), .A(n21681), .Z(n9167) );
  OR U9887 ( .A(n9166), .B(n9167), .Z(n9171) );
  XNOR U9888 ( .A(n9167), .B(n9166), .Z(n9550) );
  XOR U9889 ( .A(n9169), .B(n9168), .Z(n9549) );
  NANDN U9890 ( .A(n9550), .B(n9549), .Z(n9170) );
  AND U9891 ( .A(n9171), .B(n9170), .Z(n9174) );
  OR U9892 ( .A(n9174), .B(n9175), .Z(n9177) );
  ANDN U9893 ( .B(b[33]), .A(n177), .Z(n9558) );
  XOR U9894 ( .A(n9175), .B(n9174), .Z(n9557) );
  NANDN U9895 ( .A(n9558), .B(n9557), .Z(n9176) );
  AND U9896 ( .A(n9177), .B(n9176), .Z(n9179) );
  OR U9897 ( .A(n9178), .B(n9179), .Z(n9183) );
  XNOR U9898 ( .A(n9179), .B(n9178), .Z(n9562) );
  XNOR U9899 ( .A(n9181), .B(n9180), .Z(n9561) );
  OR U9900 ( .A(n9562), .B(n9561), .Z(n9182) );
  AND U9901 ( .A(n9183), .B(n9182), .Z(n9187) );
  XOR U9902 ( .A(n9185), .B(n9184), .Z(n9186) );
  NANDN U9903 ( .A(n9187), .B(n9186), .Z(n9189) );
  XOR U9904 ( .A(n9187), .B(n9186), .Z(n9569) );
  ANDN U9905 ( .B(b[33]), .A(n178), .Z(n9570) );
  OR U9906 ( .A(n9569), .B(n9570), .Z(n9188) );
  AND U9907 ( .A(n9189), .B(n9188), .Z(n9193) );
  OR U9908 ( .A(n9192), .B(n9193), .Z(n9195) );
  XOR U9909 ( .A(n9193), .B(n9192), .Z(n9573) );
  NANDN U9910 ( .A(n9574), .B(n9573), .Z(n9194) );
  NAND U9911 ( .A(n9195), .B(n9194), .Z(n9198) );
  XOR U9912 ( .A(n9197), .B(n9196), .Z(n9199) );
  OR U9913 ( .A(n9198), .B(n9199), .Z(n9201) );
  NAND U9914 ( .A(a[26]), .B(b[33]), .Z(n9580) );
  XOR U9915 ( .A(n9199), .B(n9198), .Z(n9579) );
  NANDN U9916 ( .A(n9580), .B(n9579), .Z(n9200) );
  NAND U9917 ( .A(n9201), .B(n9200), .Z(n9204) );
  ANDN U9918 ( .B(b[33]), .A(n21716), .Z(n9205) );
  OR U9919 ( .A(n9204), .B(n9205), .Z(n9207) );
  XOR U9920 ( .A(n9203), .B(n9202), .Z(n9586) );
  XOR U9921 ( .A(n9205), .B(n9204), .Z(n9585) );
  NANDN U9922 ( .A(n9586), .B(n9585), .Z(n9206) );
  AND U9923 ( .A(n9207), .B(n9206), .Z(n9211) );
  XOR U9924 ( .A(n9209), .B(n9208), .Z(n9210) );
  NANDN U9925 ( .A(n9211), .B(n9210), .Z(n9213) );
  XOR U9926 ( .A(n9211), .B(n9210), .Z(n9591) );
  ANDN U9927 ( .B(b[33]), .A(n180), .Z(n9592) );
  OR U9928 ( .A(n9591), .B(n9592), .Z(n9212) );
  AND U9929 ( .A(n9213), .B(n9212), .Z(n9217) );
  OR U9930 ( .A(n9216), .B(n9217), .Z(n9219) );
  XOR U9931 ( .A(n9215), .B(n9214), .Z(n9598) );
  XOR U9932 ( .A(n9217), .B(n9216), .Z(n9597) );
  NANDN U9933 ( .A(n9598), .B(n9597), .Z(n9218) );
  NAND U9934 ( .A(n9219), .B(n9218), .Z(n9222) );
  XOR U9935 ( .A(n9221), .B(n9220), .Z(n9223) );
  OR U9936 ( .A(n9222), .B(n9223), .Z(n9225) );
  NAND U9937 ( .A(a[30]), .B(b[33]), .Z(n9604) );
  XOR U9938 ( .A(n9223), .B(n9222), .Z(n9603) );
  NANDN U9939 ( .A(n9604), .B(n9603), .Z(n9224) );
  NAND U9940 ( .A(n9225), .B(n9224), .Z(n9226) );
  ANDN U9941 ( .B(b[33]), .A(n21740), .Z(n9227) );
  OR U9942 ( .A(n9226), .B(n9227), .Z(n9231) );
  XOR U9943 ( .A(n9227), .B(n9226), .Z(n9609) );
  NAND U9944 ( .A(n9609), .B(n9610), .Z(n9230) );
  NAND U9945 ( .A(n9231), .B(n9230), .Z(n9235) );
  NAND U9946 ( .A(a[32]), .B(b[33]), .Z(n9234) );
  OR U9947 ( .A(n9235), .B(n9234), .Z(n9237) );
  XOR U9948 ( .A(n9233), .B(n9232), .Z(n9615) );
  XOR U9949 ( .A(n9235), .B(n9234), .Z(n9616) );
  NAND U9950 ( .A(n9615), .B(n9616), .Z(n9236) );
  NAND U9951 ( .A(n9237), .B(n9236), .Z(n9241) );
  XOR U9952 ( .A(n9239), .B(n9238), .Z(n9240) );
  NAND U9953 ( .A(n9241), .B(n9240), .Z(n9243) );
  XNOR U9954 ( .A(n9241), .B(n9240), .Z(n9622) );
  NAND U9955 ( .A(a[33]), .B(b[33]), .Z(n9621) );
  OR U9956 ( .A(n9622), .B(n9621), .Z(n9242) );
  NAND U9957 ( .A(n9243), .B(n9242), .Z(n9247) );
  NANDN U9958 ( .A(n9246), .B(n9247), .Z(n9249) );
  XNOR U9959 ( .A(n9245), .B(n9244), .Z(n9628) );
  XNOR U9960 ( .A(n9247), .B(n9246), .Z(n9627) );
  NANDN U9961 ( .A(n9628), .B(n9627), .Z(n9248) );
  NAND U9962 ( .A(n9249), .B(n9248), .Z(n9253) );
  XOR U9963 ( .A(n9251), .B(n9250), .Z(n9252) );
  NAND U9964 ( .A(n9253), .B(n9252), .Z(n9255) );
  XNOR U9965 ( .A(n9253), .B(n9252), .Z(n9634) );
  NAND U9966 ( .A(a[35]), .B(b[33]), .Z(n9633) );
  OR U9967 ( .A(n9634), .B(n9633), .Z(n9254) );
  NAND U9968 ( .A(n9255), .B(n9254), .Z(n9259) );
  NANDN U9969 ( .A(n9258), .B(n9259), .Z(n9261) );
  XNOR U9970 ( .A(n9257), .B(n9256), .Z(n9640) );
  XNOR U9971 ( .A(n9259), .B(n9258), .Z(n9639) );
  NANDN U9972 ( .A(n9640), .B(n9639), .Z(n9260) );
  NAND U9973 ( .A(n9261), .B(n9260), .Z(n9265) );
  XOR U9974 ( .A(n9263), .B(n9262), .Z(n9264) );
  NAND U9975 ( .A(n9265), .B(n9264), .Z(n9267) );
  XNOR U9976 ( .A(n9265), .B(n9264), .Z(n9646) );
  NAND U9977 ( .A(a[37]), .B(b[33]), .Z(n9645) );
  OR U9978 ( .A(n9646), .B(n9645), .Z(n9266) );
  NAND U9979 ( .A(n9267), .B(n9266), .Z(n9271) );
  NANDN U9980 ( .A(n9270), .B(n9271), .Z(n9273) );
  XNOR U9981 ( .A(n9269), .B(n9268), .Z(n9652) );
  XNOR U9982 ( .A(n9271), .B(n9270), .Z(n9651) );
  NANDN U9983 ( .A(n9652), .B(n9651), .Z(n9272) );
  NAND U9984 ( .A(n9273), .B(n9272), .Z(n9277) );
  XOR U9985 ( .A(n9275), .B(n9274), .Z(n9276) );
  NAND U9986 ( .A(n9277), .B(n9276), .Z(n9279) );
  XNOR U9987 ( .A(n9277), .B(n9276), .Z(n9658) );
  NAND U9988 ( .A(a[39]), .B(b[33]), .Z(n9657) );
  OR U9989 ( .A(n9658), .B(n9657), .Z(n9278) );
  NAND U9990 ( .A(n9279), .B(n9278), .Z(n9283) );
  NANDN U9991 ( .A(n9282), .B(n9283), .Z(n9285) );
  XNOR U9992 ( .A(n9281), .B(n9280), .Z(n9664) );
  XNOR U9993 ( .A(n9283), .B(n9282), .Z(n9663) );
  NANDN U9994 ( .A(n9664), .B(n9663), .Z(n9284) );
  NAND U9995 ( .A(n9285), .B(n9284), .Z(n9289) );
  XOR U9996 ( .A(n9287), .B(n9286), .Z(n9288) );
  NAND U9997 ( .A(n9289), .B(n9288), .Z(n9291) );
  XNOR U9998 ( .A(n9289), .B(n9288), .Z(n9670) );
  NAND U9999 ( .A(a[41]), .B(b[33]), .Z(n9669) );
  OR U10000 ( .A(n9670), .B(n9669), .Z(n9290) );
  NAND U10001 ( .A(n9291), .B(n9290), .Z(n9295) );
  NANDN U10002 ( .A(n9294), .B(n9295), .Z(n9297) );
  XNOR U10003 ( .A(n9293), .B(n9292), .Z(n9676) );
  XNOR U10004 ( .A(n9295), .B(n9294), .Z(n9675) );
  NANDN U10005 ( .A(n9676), .B(n9675), .Z(n9296) );
  NAND U10006 ( .A(n9297), .B(n9296), .Z(n9301) );
  XOR U10007 ( .A(n9299), .B(n9298), .Z(n9300) );
  NAND U10008 ( .A(n9301), .B(n9300), .Z(n9303) );
  XNOR U10009 ( .A(n9301), .B(n9300), .Z(n9682) );
  NAND U10010 ( .A(a[43]), .B(b[33]), .Z(n9681) );
  OR U10011 ( .A(n9682), .B(n9681), .Z(n9302) );
  NAND U10012 ( .A(n9303), .B(n9302), .Z(n9307) );
  NANDN U10013 ( .A(n9306), .B(n9307), .Z(n9309) );
  XNOR U10014 ( .A(n9305), .B(n9304), .Z(n9688) );
  XNOR U10015 ( .A(n9307), .B(n9306), .Z(n9687) );
  NANDN U10016 ( .A(n9688), .B(n9687), .Z(n9308) );
  NAND U10017 ( .A(n9309), .B(n9308), .Z(n9313) );
  XOR U10018 ( .A(n9311), .B(n9310), .Z(n9312) );
  NAND U10019 ( .A(n9313), .B(n9312), .Z(n9315) );
  XNOR U10020 ( .A(n9313), .B(n9312), .Z(n9694) );
  NAND U10021 ( .A(a[45]), .B(b[33]), .Z(n9693) );
  OR U10022 ( .A(n9694), .B(n9693), .Z(n9314) );
  NAND U10023 ( .A(n9315), .B(n9314), .Z(n9319) );
  NANDN U10024 ( .A(n9318), .B(n9319), .Z(n9321) );
  XNOR U10025 ( .A(n9317), .B(n9316), .Z(n9700) );
  XNOR U10026 ( .A(n9319), .B(n9318), .Z(n9699) );
  NANDN U10027 ( .A(n9700), .B(n9699), .Z(n9320) );
  NAND U10028 ( .A(n9321), .B(n9320), .Z(n9325) );
  XOR U10029 ( .A(n9323), .B(n9322), .Z(n9324) );
  NAND U10030 ( .A(n9325), .B(n9324), .Z(n9327) );
  XNOR U10031 ( .A(n9325), .B(n9324), .Z(n9706) );
  NAND U10032 ( .A(a[47]), .B(b[33]), .Z(n9705) );
  OR U10033 ( .A(n9706), .B(n9705), .Z(n9326) );
  NAND U10034 ( .A(n9327), .B(n9326), .Z(n9331) );
  NANDN U10035 ( .A(n9330), .B(n9331), .Z(n9333) );
  XNOR U10036 ( .A(n9329), .B(n9328), .Z(n9712) );
  XNOR U10037 ( .A(n9331), .B(n9330), .Z(n9711) );
  NANDN U10038 ( .A(n9712), .B(n9711), .Z(n9332) );
  NAND U10039 ( .A(n9333), .B(n9332), .Z(n9337) );
  NANDN U10040 ( .A(n9336), .B(n9337), .Z(n9339) );
  XOR U10041 ( .A(n9335), .B(n9334), .Z(n9717) );
  XNOR U10042 ( .A(n9337), .B(n9336), .Z(n9718) );
  NAND U10043 ( .A(n9717), .B(n9718), .Z(n9338) );
  NAND U10044 ( .A(n9339), .B(n9338), .Z(n9343) );
  NANDN U10045 ( .A(n9342), .B(n9343), .Z(n9345) );
  XNOR U10046 ( .A(n9341), .B(n9340), .Z(n9724) );
  XNOR U10047 ( .A(n9343), .B(n9342), .Z(n9723) );
  NANDN U10048 ( .A(n9724), .B(n9723), .Z(n9344) );
  NAND U10049 ( .A(n9345), .B(n9344), .Z(n9349) );
  NANDN U10050 ( .A(n9348), .B(n9349), .Z(n9351) );
  XOR U10051 ( .A(n9347), .B(n9346), .Z(n9729) );
  XNOR U10052 ( .A(n9349), .B(n9348), .Z(n9730) );
  NAND U10053 ( .A(n9729), .B(n9730), .Z(n9350) );
  NAND U10054 ( .A(n9351), .B(n9350), .Z(n9355) );
  NANDN U10055 ( .A(n9354), .B(n9355), .Z(n9357) );
  XNOR U10056 ( .A(n9353), .B(n9352), .Z(n9736) );
  XNOR U10057 ( .A(n9355), .B(n9354), .Z(n9735) );
  NANDN U10058 ( .A(n9736), .B(n9735), .Z(n9356) );
  NAND U10059 ( .A(n9357), .B(n9356), .Z(n9361) );
  NANDN U10060 ( .A(n9360), .B(n9361), .Z(n9363) );
  XOR U10061 ( .A(n9359), .B(n9358), .Z(n9741) );
  XNOR U10062 ( .A(n9361), .B(n9360), .Z(n9742) );
  NAND U10063 ( .A(n9741), .B(n9742), .Z(n9362) );
  NAND U10064 ( .A(n9363), .B(n9362), .Z(n9367) );
  NANDN U10065 ( .A(n9366), .B(n9367), .Z(n9369) );
  XNOR U10066 ( .A(n9365), .B(n9364), .Z(n9748) );
  XNOR U10067 ( .A(n9367), .B(n9366), .Z(n9747) );
  NANDN U10068 ( .A(n9748), .B(n9747), .Z(n9368) );
  NAND U10069 ( .A(n9369), .B(n9368), .Z(n9373) );
  NANDN U10070 ( .A(n9372), .B(n9373), .Z(n9375) );
  XOR U10071 ( .A(n9371), .B(n9370), .Z(n9753) );
  XNOR U10072 ( .A(n9373), .B(n9372), .Z(n9754) );
  NAND U10073 ( .A(n9753), .B(n9754), .Z(n9374) );
  NAND U10074 ( .A(n9375), .B(n9374), .Z(n9379) );
  NANDN U10075 ( .A(n9378), .B(n9379), .Z(n9381) );
  XNOR U10076 ( .A(n9377), .B(n9376), .Z(n9760) );
  XNOR U10077 ( .A(n9379), .B(n9378), .Z(n9759) );
  NANDN U10078 ( .A(n9760), .B(n9759), .Z(n9380) );
  NAND U10079 ( .A(n9381), .B(n9380), .Z(n9385) );
  NANDN U10080 ( .A(n9384), .B(n9385), .Z(n9387) );
  XOR U10081 ( .A(n9383), .B(n9382), .Z(n9765) );
  XNOR U10082 ( .A(n9385), .B(n9384), .Z(n9766) );
  NAND U10083 ( .A(n9765), .B(n9766), .Z(n9386) );
  NAND U10084 ( .A(n9387), .B(n9386), .Z(n9391) );
  NANDN U10085 ( .A(n9390), .B(n9391), .Z(n9393) );
  XNOR U10086 ( .A(n9389), .B(n9388), .Z(n9772) );
  XNOR U10087 ( .A(n9391), .B(n9390), .Z(n9771) );
  NANDN U10088 ( .A(n9772), .B(n9771), .Z(n9392) );
  NAND U10089 ( .A(n9393), .B(n9392), .Z(n9397) );
  NANDN U10090 ( .A(n9396), .B(n9397), .Z(n9399) );
  XOR U10091 ( .A(n9395), .B(n9394), .Z(n9777) );
  XNOR U10092 ( .A(n9397), .B(n9396), .Z(n9778) );
  NAND U10093 ( .A(n9777), .B(n9778), .Z(n9398) );
  NAND U10094 ( .A(n9399), .B(n9398), .Z(n9403) );
  NANDN U10095 ( .A(n9402), .B(n9403), .Z(n9405) );
  XNOR U10096 ( .A(n9401), .B(n9400), .Z(n9784) );
  XNOR U10097 ( .A(n9403), .B(n9402), .Z(n9783) );
  NANDN U10098 ( .A(n9784), .B(n9783), .Z(n9404) );
  NAND U10099 ( .A(n9405), .B(n9404), .Z(n9409) );
  XOR U10100 ( .A(n9407), .B(n9406), .Z(n9408) );
  NAND U10101 ( .A(n9409), .B(n9408), .Z(n9411) );
  XNOR U10102 ( .A(n9409), .B(n9408), .Z(n9790) );
  NAND U10103 ( .A(a[61]), .B(b[33]), .Z(n9789) );
  OR U10104 ( .A(n9790), .B(n9789), .Z(n9410) );
  NAND U10105 ( .A(n9411), .B(n9410), .Z(n9415) );
  NANDN U10106 ( .A(n9414), .B(n9415), .Z(n9417) );
  XNOR U10107 ( .A(n9413), .B(n9412), .Z(n9796) );
  XNOR U10108 ( .A(n9415), .B(n9414), .Z(n9795) );
  NANDN U10109 ( .A(n9796), .B(n9795), .Z(n9416) );
  NAND U10110 ( .A(n9417), .B(n9416), .Z(n9420) );
  XOR U10111 ( .A(n9419), .B(n9418), .Z(n9421) );
  OR U10112 ( .A(n9420), .B(n9421), .Z(n9423) );
  AND U10113 ( .A(b[33]), .B(a[63]), .Z(n9802) );
  XOR U10114 ( .A(n9421), .B(n9420), .Z(n9801) );
  NANDN U10115 ( .A(n9802), .B(n9801), .Z(n9422) );
  AND U10116 ( .A(n9423), .B(n9422), .Z(n9424) );
  NANDN U10117 ( .A(n9425), .B(n9424), .Z(n21994) );
  OR U10118 ( .A(n21995), .B(n21994), .Z(n21997) );
  XNOR U10119 ( .A(n9425), .B(n9424), .Z(n21992) );
  NAND U10120 ( .A(a[34]), .B(b[32]), .Z(n9623) );
  ANDN U10121 ( .B(b[32]), .A(n21692), .Z(n9555) );
  ANDN U10122 ( .B(b[32]), .A(n172), .Z(n9509) );
  ANDN U10123 ( .B(b[32]), .A(n166), .Z(n9459) );
  ANDN U10124 ( .B(b[32]), .A(n21580), .Z(n9435) );
  NAND U10125 ( .A(b[33]), .B(a[1]), .Z(n9430) );
  NANDN U10126 ( .A(n9430), .B(a[0]), .Z(n9426) );
  XNOR U10127 ( .A(a[2]), .B(n9426), .Z(n9427) );
  NAND U10128 ( .A(b[32]), .B(n9427), .Z(n9817) );
  AND U10129 ( .A(a[1]), .B(b[33]), .Z(n9428) );
  XNOR U10130 ( .A(n9429), .B(n9428), .Z(n9816) );
  NANDN U10131 ( .A(n9817), .B(n9816), .Z(n9434) );
  AND U10132 ( .A(b[32]), .B(a[0]), .Z(n10186) );
  NANDN U10133 ( .A(n9430), .B(n10186), .Z(n9432) );
  NAND U10134 ( .A(a[2]), .B(b[32]), .Z(n9431) );
  AND U10135 ( .A(n9432), .B(n9431), .Z(n9433) );
  ANDN U10136 ( .B(n9434), .A(n9433), .Z(n9436) );
  OR U10137 ( .A(n9435), .B(n9436), .Z(n9440) );
  XNOR U10138 ( .A(n9436), .B(n9435), .Z(n9821) );
  XNOR U10139 ( .A(n9438), .B(n9437), .Z(n9820) );
  OR U10140 ( .A(n9821), .B(n9820), .Z(n9439) );
  NAND U10141 ( .A(n9440), .B(n9439), .Z(n9443) );
  XOR U10142 ( .A(n9442), .B(n9441), .Z(n9444) );
  OR U10143 ( .A(n9443), .B(n9444), .Z(n9446) );
  NAND U10144 ( .A(a[4]), .B(b[32]), .Z(n9829) );
  XOR U10145 ( .A(n9444), .B(n9443), .Z(n9828) );
  NANDN U10146 ( .A(n9829), .B(n9828), .Z(n9445) );
  NAND U10147 ( .A(n9446), .B(n9445), .Z(n9447) );
  ANDN U10148 ( .B(b[32]), .A(n164), .Z(n9448) );
  OR U10149 ( .A(n9447), .B(n9448), .Z(n9452) );
  XNOR U10150 ( .A(n9448), .B(n9447), .Z(n9832) );
  OR U10151 ( .A(n9832), .B(n9833), .Z(n9451) );
  AND U10152 ( .A(n9452), .B(n9451), .Z(n9456) );
  XOR U10153 ( .A(n9454), .B(n9453), .Z(n9455) );
  NANDN U10154 ( .A(n9456), .B(n9455), .Z(n9458) );
  XOR U10155 ( .A(n9456), .B(n9455), .Z(n9840) );
  ANDN U10156 ( .B(b[32]), .A(n165), .Z(n9841) );
  OR U10157 ( .A(n9840), .B(n9841), .Z(n9457) );
  AND U10158 ( .A(n9458), .B(n9457), .Z(n9460) );
  OR U10159 ( .A(n9459), .B(n9460), .Z(n9464) );
  XNOR U10160 ( .A(n9460), .B(n9459), .Z(n9845) );
  XNOR U10161 ( .A(n9462), .B(n9461), .Z(n9844) );
  OR U10162 ( .A(n9845), .B(n9844), .Z(n9463) );
  NAND U10163 ( .A(n9464), .B(n9463), .Z(n9467) );
  XOR U10164 ( .A(n9466), .B(n9465), .Z(n9468) );
  OR U10165 ( .A(n9467), .B(n9468), .Z(n9470) );
  NAND U10166 ( .A(a[8]), .B(b[32]), .Z(n9851) );
  XOR U10167 ( .A(n9468), .B(n9467), .Z(n9850) );
  NANDN U10168 ( .A(n9851), .B(n9850), .Z(n9469) );
  NAND U10169 ( .A(n9470), .B(n9469), .Z(n9473) );
  ANDN U10170 ( .B(b[32]), .A(n21615), .Z(n9474) );
  OR U10171 ( .A(n9473), .B(n9474), .Z(n9476) );
  XOR U10172 ( .A(n9472), .B(n9471), .Z(n9857) );
  XOR U10173 ( .A(n9474), .B(n9473), .Z(n9856) );
  NANDN U10174 ( .A(n9857), .B(n9856), .Z(n9475) );
  NAND U10175 ( .A(n9476), .B(n9475), .Z(n9479) );
  XOR U10176 ( .A(n9478), .B(n9477), .Z(n9480) );
  OR U10177 ( .A(n9479), .B(n9480), .Z(n9482) );
  NAND U10178 ( .A(a[10]), .B(b[32]), .Z(n9863) );
  XOR U10179 ( .A(n9480), .B(n9479), .Z(n9862) );
  NANDN U10180 ( .A(n9863), .B(n9862), .Z(n9481) );
  NAND U10181 ( .A(n9482), .B(n9481), .Z(n9485) );
  ANDN U10182 ( .B(b[32]), .A(n21164), .Z(n9486) );
  OR U10183 ( .A(n9485), .B(n9486), .Z(n9488) );
  XOR U10184 ( .A(n9486), .B(n9485), .Z(n9868) );
  NANDN U10185 ( .A(n9869), .B(n9868), .Z(n9487) );
  NAND U10186 ( .A(n9488), .B(n9487), .Z(n9491) );
  XNOR U10187 ( .A(n9490), .B(n9489), .Z(n9492) );
  OR U10188 ( .A(n9491), .B(n9492), .Z(n9494) );
  XNOR U10189 ( .A(n9492), .B(n9491), .Z(n9875) );
  NAND U10190 ( .A(a[12]), .B(b[32]), .Z(n9874) );
  OR U10191 ( .A(n9875), .B(n9874), .Z(n9493) );
  NAND U10192 ( .A(n9494), .B(n9493), .Z(n9495) );
  ANDN U10193 ( .B(b[32]), .A(n170), .Z(n9496) );
  OR U10194 ( .A(n9495), .B(n9496), .Z(n9500) );
  XNOR U10195 ( .A(n9496), .B(n9495), .Z(n9881) );
  XNOR U10196 ( .A(n9498), .B(n9497), .Z(n9880) );
  OR U10197 ( .A(n9881), .B(n9880), .Z(n9499) );
  AND U10198 ( .A(n9500), .B(n9499), .Z(n9503) );
  OR U10199 ( .A(n9503), .B(n9504), .Z(n9506) );
  ANDN U10200 ( .B(b[32]), .A(n171), .Z(n9889) );
  XOR U10201 ( .A(n9504), .B(n9503), .Z(n9888) );
  NANDN U10202 ( .A(n9889), .B(n9888), .Z(n9505) );
  AND U10203 ( .A(n9506), .B(n9505), .Z(n9510) );
  OR U10204 ( .A(n9509), .B(n9510), .Z(n9512) );
  XOR U10205 ( .A(n9508), .B(n9507), .Z(n9893) );
  XOR U10206 ( .A(n9510), .B(n9509), .Z(n9892) );
  NANDN U10207 ( .A(n9893), .B(n9892), .Z(n9511) );
  NAND U10208 ( .A(n9512), .B(n9511), .Z(n9515) );
  XOR U10209 ( .A(n9514), .B(n9513), .Z(n9516) );
  OR U10210 ( .A(n9515), .B(n9516), .Z(n9518) );
  NAND U10211 ( .A(a[16]), .B(b[32]), .Z(n9899) );
  XOR U10212 ( .A(n9516), .B(n9515), .Z(n9898) );
  NANDN U10213 ( .A(n9899), .B(n9898), .Z(n9517) );
  NAND U10214 ( .A(n9518), .B(n9517), .Z(n9521) );
  ANDN U10215 ( .B(b[32]), .A(n174), .Z(n9522) );
  OR U10216 ( .A(n9521), .B(n9522), .Z(n9524) );
  XOR U10217 ( .A(n9520), .B(n9519), .Z(n9905) );
  XOR U10218 ( .A(n9522), .B(n9521), .Z(n9904) );
  NANDN U10219 ( .A(n9905), .B(n9904), .Z(n9523) );
  NAND U10220 ( .A(n9524), .B(n9523), .Z(n9527) );
  XNOR U10221 ( .A(n9526), .B(n9525), .Z(n9528) );
  OR U10222 ( .A(n9527), .B(n9528), .Z(n9530) );
  XNOR U10223 ( .A(n9528), .B(n9527), .Z(n9911) );
  NAND U10224 ( .A(a[18]), .B(b[32]), .Z(n9910) );
  OR U10225 ( .A(n9911), .B(n9910), .Z(n9529) );
  NAND U10226 ( .A(n9530), .B(n9529), .Z(n9533) );
  ANDN U10227 ( .B(b[32]), .A(n21670), .Z(n9534) );
  OR U10228 ( .A(n9533), .B(n9534), .Z(n9536) );
  XOR U10229 ( .A(n9534), .B(n9533), .Z(n9916) );
  NANDN U10230 ( .A(n9917), .B(n9916), .Z(n9535) );
  NAND U10231 ( .A(n9536), .B(n9535), .Z(n9539) );
  XNOR U10232 ( .A(n9538), .B(n9537), .Z(n9540) );
  OR U10233 ( .A(n9539), .B(n9540), .Z(n9542) );
  XNOR U10234 ( .A(n9540), .B(n9539), .Z(n9923) );
  NAND U10235 ( .A(a[20]), .B(b[32]), .Z(n9922) );
  OR U10236 ( .A(n9923), .B(n9922), .Z(n9541) );
  NAND U10237 ( .A(n9542), .B(n9541), .Z(n9545) );
  ANDN U10238 ( .B(b[32]), .A(n21681), .Z(n9546) );
  OR U10239 ( .A(n9545), .B(n9546), .Z(n9548) );
  XOR U10240 ( .A(n9544), .B(n9543), .Z(n9929) );
  XOR U10241 ( .A(n9546), .B(n9545), .Z(n9928) );
  NANDN U10242 ( .A(n9929), .B(n9928), .Z(n9547) );
  AND U10243 ( .A(n9548), .B(n9547), .Z(n9552) );
  NANDN U10244 ( .A(n9552), .B(n9551), .Z(n9554) );
  XOR U10245 ( .A(n9552), .B(n9551), .Z(n9934) );
  ANDN U10246 ( .B(b[32]), .A(n177), .Z(n9935) );
  OR U10247 ( .A(n9934), .B(n9935), .Z(n9553) );
  AND U10248 ( .A(n9554), .B(n9553), .Z(n9556) );
  OR U10249 ( .A(n9555), .B(n9556), .Z(n9560) );
  XNOR U10250 ( .A(n9556), .B(n9555), .Z(n9941) );
  OR U10251 ( .A(n9941), .B(n9940), .Z(n9559) );
  NAND U10252 ( .A(n9560), .B(n9559), .Z(n9563) );
  XOR U10253 ( .A(n9562), .B(n9561), .Z(n9564) );
  OR U10254 ( .A(n9563), .B(n9564), .Z(n9566) );
  NAND U10255 ( .A(a[24]), .B(b[32]), .Z(n9949) );
  XOR U10256 ( .A(n9564), .B(n9563), .Z(n9948) );
  NANDN U10257 ( .A(n9949), .B(n9948), .Z(n9565) );
  NAND U10258 ( .A(n9566), .B(n9565), .Z(n9567) );
  ANDN U10259 ( .B(b[32]), .A(n21703), .Z(n9568) );
  OR U10260 ( .A(n9567), .B(n9568), .Z(n9572) );
  XNOR U10261 ( .A(n9568), .B(n9567), .Z(n9953) );
  XNOR U10262 ( .A(n9570), .B(n9569), .Z(n9952) );
  OR U10263 ( .A(n9953), .B(n9952), .Z(n9571) );
  NAND U10264 ( .A(n9572), .B(n9571), .Z(n9575) );
  XNOR U10265 ( .A(n9574), .B(n9573), .Z(n9576) );
  OR U10266 ( .A(n9575), .B(n9576), .Z(n9578) );
  XNOR U10267 ( .A(n9576), .B(n9575), .Z(n9961) );
  NAND U10268 ( .A(a[26]), .B(b[32]), .Z(n9960) );
  OR U10269 ( .A(n9961), .B(n9960), .Z(n9577) );
  NAND U10270 ( .A(n9578), .B(n9577), .Z(n9581) );
  ANDN U10271 ( .B(b[32]), .A(n21716), .Z(n9582) );
  OR U10272 ( .A(n9581), .B(n9582), .Z(n9584) );
  XOR U10273 ( .A(n9582), .B(n9581), .Z(n9964) );
  NANDN U10274 ( .A(n9965), .B(n9964), .Z(n9583) );
  NAND U10275 ( .A(n9584), .B(n9583), .Z(n9587) );
  XNOR U10276 ( .A(n9586), .B(n9585), .Z(n9588) );
  OR U10277 ( .A(n9587), .B(n9588), .Z(n9590) );
  XNOR U10278 ( .A(n9588), .B(n9587), .Z(n9971) );
  NAND U10279 ( .A(a[28]), .B(b[32]), .Z(n9970) );
  OR U10280 ( .A(n9971), .B(n9970), .Z(n9589) );
  NAND U10281 ( .A(n9590), .B(n9589), .Z(n9593) );
  ANDN U10282 ( .B(b[32]), .A(n21727), .Z(n9594) );
  OR U10283 ( .A(n9593), .B(n9594), .Z(n9596) );
  XNOR U10284 ( .A(n9592), .B(n9591), .Z(n9977) );
  XNOR U10285 ( .A(n9594), .B(n9593), .Z(n9976) );
  OR U10286 ( .A(n9977), .B(n9976), .Z(n9595) );
  NAND U10287 ( .A(n9596), .B(n9595), .Z(n9599) );
  XNOR U10288 ( .A(n9598), .B(n9597), .Z(n9600) );
  OR U10289 ( .A(n9599), .B(n9600), .Z(n9602) );
  XNOR U10290 ( .A(n9600), .B(n9599), .Z(n9983) );
  NAND U10291 ( .A(a[30]), .B(b[32]), .Z(n9982) );
  OR U10292 ( .A(n9983), .B(n9982), .Z(n9601) );
  NAND U10293 ( .A(n9602), .B(n9601), .Z(n9605) );
  ANDN U10294 ( .B(b[32]), .A(n21740), .Z(n9606) );
  OR U10295 ( .A(n9605), .B(n9606), .Z(n9608) );
  XOR U10296 ( .A(n9606), .B(n9605), .Z(n9988) );
  NANDN U10297 ( .A(n9989), .B(n9988), .Z(n9607) );
  NAND U10298 ( .A(n9608), .B(n9607), .Z(n9612) );
  AND U10299 ( .A(b[32]), .B(a[32]), .Z(n9611) );
  NANDN U10300 ( .A(n9612), .B(n9611), .Z(n9614) );
  XNOR U10301 ( .A(n9612), .B(n9611), .Z(n9996) );
  NANDN U10302 ( .A(n9997), .B(n9996), .Z(n9613) );
  NAND U10303 ( .A(n9614), .B(n9613), .Z(n9618) );
  XOR U10304 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U10305 ( .A(n9618), .B(n9617), .Z(n9620) );
  XNOR U10306 ( .A(n9618), .B(n9617), .Z(n10001) );
  NAND U10307 ( .A(a[33]), .B(b[32]), .Z(n10000) );
  OR U10308 ( .A(n10001), .B(n10000), .Z(n9619) );
  NAND U10309 ( .A(n9620), .B(n9619), .Z(n9624) );
  NANDN U10310 ( .A(n9623), .B(n9624), .Z(n9626) );
  XOR U10311 ( .A(n9622), .B(n9621), .Z(n10006) );
  XNOR U10312 ( .A(n9624), .B(n9623), .Z(n10007) );
  NAND U10313 ( .A(n10006), .B(n10007), .Z(n9625) );
  NAND U10314 ( .A(n9626), .B(n9625), .Z(n9629) );
  AND U10315 ( .A(b[32]), .B(a[35]), .Z(n9630) );
  OR U10316 ( .A(n9629), .B(n9630), .Z(n9632) );
  XNOR U10317 ( .A(n9628), .B(n9627), .Z(n10013) );
  XOR U10318 ( .A(n9630), .B(n9629), .Z(n10012) );
  NANDN U10319 ( .A(n10013), .B(n10012), .Z(n9631) );
  NAND U10320 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U10321 ( .A(a[36]), .B(b[32]), .Z(n9635) );
  OR U10322 ( .A(n9636), .B(n9635), .Z(n9638) );
  XOR U10323 ( .A(n9634), .B(n9633), .Z(n10018) );
  XOR U10324 ( .A(n9636), .B(n9635), .Z(n10019) );
  NAND U10325 ( .A(n10018), .B(n10019), .Z(n9637) );
  NAND U10326 ( .A(n9638), .B(n9637), .Z(n9641) );
  AND U10327 ( .A(b[32]), .B(a[37]), .Z(n9642) );
  OR U10328 ( .A(n9641), .B(n9642), .Z(n9644) );
  XNOR U10329 ( .A(n9640), .B(n9639), .Z(n10025) );
  XOR U10330 ( .A(n9642), .B(n9641), .Z(n10024) );
  NANDN U10331 ( .A(n10025), .B(n10024), .Z(n9643) );
  NAND U10332 ( .A(n9644), .B(n9643), .Z(n9648) );
  NAND U10333 ( .A(a[38]), .B(b[32]), .Z(n9647) );
  OR U10334 ( .A(n9648), .B(n9647), .Z(n9650) );
  XOR U10335 ( .A(n9646), .B(n9645), .Z(n10030) );
  XOR U10336 ( .A(n9648), .B(n9647), .Z(n10031) );
  NAND U10337 ( .A(n10030), .B(n10031), .Z(n9649) );
  NAND U10338 ( .A(n9650), .B(n9649), .Z(n9653) );
  AND U10339 ( .A(b[32]), .B(a[39]), .Z(n9654) );
  OR U10340 ( .A(n9653), .B(n9654), .Z(n9656) );
  XNOR U10341 ( .A(n9652), .B(n9651), .Z(n10037) );
  XOR U10342 ( .A(n9654), .B(n9653), .Z(n10036) );
  NANDN U10343 ( .A(n10037), .B(n10036), .Z(n9655) );
  NAND U10344 ( .A(n9656), .B(n9655), .Z(n9660) );
  NAND U10345 ( .A(a[40]), .B(b[32]), .Z(n9659) );
  OR U10346 ( .A(n9660), .B(n9659), .Z(n9662) );
  XOR U10347 ( .A(n9658), .B(n9657), .Z(n10042) );
  XOR U10348 ( .A(n9660), .B(n9659), .Z(n10043) );
  NAND U10349 ( .A(n10042), .B(n10043), .Z(n9661) );
  NAND U10350 ( .A(n9662), .B(n9661), .Z(n9665) );
  AND U10351 ( .A(b[32]), .B(a[41]), .Z(n9666) );
  OR U10352 ( .A(n9665), .B(n9666), .Z(n9668) );
  XNOR U10353 ( .A(n9664), .B(n9663), .Z(n10049) );
  XOR U10354 ( .A(n9666), .B(n9665), .Z(n10048) );
  NANDN U10355 ( .A(n10049), .B(n10048), .Z(n9667) );
  NAND U10356 ( .A(n9668), .B(n9667), .Z(n9672) );
  NAND U10357 ( .A(a[42]), .B(b[32]), .Z(n9671) );
  OR U10358 ( .A(n9672), .B(n9671), .Z(n9674) );
  XOR U10359 ( .A(n9670), .B(n9669), .Z(n10054) );
  XOR U10360 ( .A(n9672), .B(n9671), .Z(n10055) );
  NAND U10361 ( .A(n10054), .B(n10055), .Z(n9673) );
  NAND U10362 ( .A(n9674), .B(n9673), .Z(n9677) );
  AND U10363 ( .A(b[32]), .B(a[43]), .Z(n9678) );
  OR U10364 ( .A(n9677), .B(n9678), .Z(n9680) );
  XNOR U10365 ( .A(n9676), .B(n9675), .Z(n10061) );
  XOR U10366 ( .A(n9678), .B(n9677), .Z(n10060) );
  NANDN U10367 ( .A(n10061), .B(n10060), .Z(n9679) );
  NAND U10368 ( .A(n9680), .B(n9679), .Z(n9684) );
  NAND U10369 ( .A(a[44]), .B(b[32]), .Z(n9683) );
  OR U10370 ( .A(n9684), .B(n9683), .Z(n9686) );
  XOR U10371 ( .A(n9682), .B(n9681), .Z(n10066) );
  XOR U10372 ( .A(n9684), .B(n9683), .Z(n10067) );
  NAND U10373 ( .A(n10066), .B(n10067), .Z(n9685) );
  NAND U10374 ( .A(n9686), .B(n9685), .Z(n9689) );
  AND U10375 ( .A(b[32]), .B(a[45]), .Z(n9690) );
  OR U10376 ( .A(n9689), .B(n9690), .Z(n9692) );
  XNOR U10377 ( .A(n9688), .B(n9687), .Z(n10073) );
  XOR U10378 ( .A(n9690), .B(n9689), .Z(n10072) );
  NANDN U10379 ( .A(n10073), .B(n10072), .Z(n9691) );
  NAND U10380 ( .A(n9692), .B(n9691), .Z(n9696) );
  NAND U10381 ( .A(a[46]), .B(b[32]), .Z(n9695) );
  OR U10382 ( .A(n9696), .B(n9695), .Z(n9698) );
  XOR U10383 ( .A(n9694), .B(n9693), .Z(n10078) );
  XOR U10384 ( .A(n9696), .B(n9695), .Z(n10079) );
  NAND U10385 ( .A(n10078), .B(n10079), .Z(n9697) );
  NAND U10386 ( .A(n9698), .B(n9697), .Z(n9701) );
  AND U10387 ( .A(b[32]), .B(a[47]), .Z(n9702) );
  OR U10388 ( .A(n9701), .B(n9702), .Z(n9704) );
  XNOR U10389 ( .A(n9700), .B(n9699), .Z(n10085) );
  XOR U10390 ( .A(n9702), .B(n9701), .Z(n10084) );
  NANDN U10391 ( .A(n10085), .B(n10084), .Z(n9703) );
  NAND U10392 ( .A(n9704), .B(n9703), .Z(n9708) );
  NAND U10393 ( .A(a[48]), .B(b[32]), .Z(n9707) );
  OR U10394 ( .A(n9708), .B(n9707), .Z(n9710) );
  XOR U10395 ( .A(n9706), .B(n9705), .Z(n10090) );
  XOR U10396 ( .A(n9708), .B(n9707), .Z(n10091) );
  NAND U10397 ( .A(n10090), .B(n10091), .Z(n9709) );
  NAND U10398 ( .A(n9710), .B(n9709), .Z(n9713) );
  AND U10399 ( .A(b[32]), .B(a[49]), .Z(n9714) );
  OR U10400 ( .A(n9713), .B(n9714), .Z(n9716) );
  XNOR U10401 ( .A(n9712), .B(n9711), .Z(n10097) );
  XOR U10402 ( .A(n9714), .B(n9713), .Z(n10096) );
  NANDN U10403 ( .A(n10097), .B(n10096), .Z(n9715) );
  NAND U10404 ( .A(n9716), .B(n9715), .Z(n9720) );
  NAND U10405 ( .A(a[50]), .B(b[32]), .Z(n9719) );
  OR U10406 ( .A(n9720), .B(n9719), .Z(n9722) );
  XOR U10407 ( .A(n9718), .B(n9717), .Z(n10102) );
  XOR U10408 ( .A(n9720), .B(n9719), .Z(n10103) );
  NAND U10409 ( .A(n10102), .B(n10103), .Z(n9721) );
  NAND U10410 ( .A(n9722), .B(n9721), .Z(n9725) );
  AND U10411 ( .A(b[32]), .B(a[51]), .Z(n9726) );
  OR U10412 ( .A(n9725), .B(n9726), .Z(n9728) );
  XNOR U10413 ( .A(n9724), .B(n9723), .Z(n10109) );
  XOR U10414 ( .A(n9726), .B(n9725), .Z(n10108) );
  NANDN U10415 ( .A(n10109), .B(n10108), .Z(n9727) );
  NAND U10416 ( .A(n9728), .B(n9727), .Z(n9732) );
  NAND U10417 ( .A(a[52]), .B(b[32]), .Z(n9731) );
  OR U10418 ( .A(n9732), .B(n9731), .Z(n9734) );
  XOR U10419 ( .A(n9730), .B(n9729), .Z(n10114) );
  XOR U10420 ( .A(n9732), .B(n9731), .Z(n10115) );
  NAND U10421 ( .A(n10114), .B(n10115), .Z(n9733) );
  NAND U10422 ( .A(n9734), .B(n9733), .Z(n9737) );
  AND U10423 ( .A(b[32]), .B(a[53]), .Z(n9738) );
  OR U10424 ( .A(n9737), .B(n9738), .Z(n9740) );
  XNOR U10425 ( .A(n9736), .B(n9735), .Z(n10121) );
  XOR U10426 ( .A(n9738), .B(n9737), .Z(n10120) );
  NANDN U10427 ( .A(n10121), .B(n10120), .Z(n9739) );
  NAND U10428 ( .A(n9740), .B(n9739), .Z(n9744) );
  NAND U10429 ( .A(a[54]), .B(b[32]), .Z(n9743) );
  OR U10430 ( .A(n9744), .B(n9743), .Z(n9746) );
  XOR U10431 ( .A(n9742), .B(n9741), .Z(n10126) );
  XOR U10432 ( .A(n9744), .B(n9743), .Z(n10127) );
  NAND U10433 ( .A(n10126), .B(n10127), .Z(n9745) );
  NAND U10434 ( .A(n9746), .B(n9745), .Z(n9749) );
  AND U10435 ( .A(b[32]), .B(a[55]), .Z(n9750) );
  OR U10436 ( .A(n9749), .B(n9750), .Z(n9752) );
  XNOR U10437 ( .A(n9748), .B(n9747), .Z(n10133) );
  XOR U10438 ( .A(n9750), .B(n9749), .Z(n10132) );
  NANDN U10439 ( .A(n10133), .B(n10132), .Z(n9751) );
  NAND U10440 ( .A(n9752), .B(n9751), .Z(n9756) );
  NAND U10441 ( .A(a[56]), .B(b[32]), .Z(n9755) );
  OR U10442 ( .A(n9756), .B(n9755), .Z(n9758) );
  XOR U10443 ( .A(n9754), .B(n9753), .Z(n10138) );
  XOR U10444 ( .A(n9756), .B(n9755), .Z(n10139) );
  NAND U10445 ( .A(n10138), .B(n10139), .Z(n9757) );
  NAND U10446 ( .A(n9758), .B(n9757), .Z(n9761) );
  AND U10447 ( .A(b[32]), .B(a[57]), .Z(n9762) );
  OR U10448 ( .A(n9761), .B(n9762), .Z(n9764) );
  XNOR U10449 ( .A(n9760), .B(n9759), .Z(n10145) );
  XOR U10450 ( .A(n9762), .B(n9761), .Z(n10144) );
  NANDN U10451 ( .A(n10145), .B(n10144), .Z(n9763) );
  NAND U10452 ( .A(n9764), .B(n9763), .Z(n9768) );
  NAND U10453 ( .A(a[58]), .B(b[32]), .Z(n9767) );
  OR U10454 ( .A(n9768), .B(n9767), .Z(n9770) );
  XOR U10455 ( .A(n9766), .B(n9765), .Z(n10150) );
  XOR U10456 ( .A(n9768), .B(n9767), .Z(n10151) );
  NAND U10457 ( .A(n10150), .B(n10151), .Z(n9769) );
  NAND U10458 ( .A(n9770), .B(n9769), .Z(n9773) );
  AND U10459 ( .A(b[32]), .B(a[59]), .Z(n9774) );
  OR U10460 ( .A(n9773), .B(n9774), .Z(n9776) );
  XNOR U10461 ( .A(n9772), .B(n9771), .Z(n10155) );
  XOR U10462 ( .A(n9774), .B(n9773), .Z(n10154) );
  NANDN U10463 ( .A(n10155), .B(n10154), .Z(n9775) );
  NAND U10464 ( .A(n9776), .B(n9775), .Z(n9780) );
  NAND U10465 ( .A(a[60]), .B(b[32]), .Z(n9779) );
  OR U10466 ( .A(n9780), .B(n9779), .Z(n9782) );
  XOR U10467 ( .A(n9778), .B(n9777), .Z(n10160) );
  XOR U10468 ( .A(n9780), .B(n9779), .Z(n10161) );
  NAND U10469 ( .A(n10160), .B(n10161), .Z(n9781) );
  NAND U10470 ( .A(n9782), .B(n9781), .Z(n9785) );
  AND U10471 ( .A(b[32]), .B(a[61]), .Z(n9786) );
  OR U10472 ( .A(n9785), .B(n9786), .Z(n9788) );
  XNOR U10473 ( .A(n9784), .B(n9783), .Z(n10167) );
  XOR U10474 ( .A(n9786), .B(n9785), .Z(n10166) );
  NANDN U10475 ( .A(n10167), .B(n10166), .Z(n9787) );
  NAND U10476 ( .A(n9788), .B(n9787), .Z(n9792) );
  NAND U10477 ( .A(a[62]), .B(b[32]), .Z(n9791) );
  OR U10478 ( .A(n9792), .B(n9791), .Z(n9794) );
  XOR U10479 ( .A(n9790), .B(n9789), .Z(n10172) );
  XOR U10480 ( .A(n9792), .B(n9791), .Z(n10173) );
  NAND U10481 ( .A(n10172), .B(n10173), .Z(n9793) );
  NAND U10482 ( .A(n9794), .B(n9793), .Z(n9797) );
  AND U10483 ( .A(b[32]), .B(a[63]), .Z(n9798) );
  OR U10484 ( .A(n9797), .B(n9798), .Z(n9800) );
  XNOR U10485 ( .A(n9796), .B(n9795), .Z(n10177) );
  XOR U10486 ( .A(n9798), .B(n9797), .Z(n10176) );
  NANDN U10487 ( .A(n10177), .B(n10176), .Z(n9799) );
  AND U10488 ( .A(n9800), .B(n9799), .Z(n9803) );
  XOR U10489 ( .A(n9802), .B(n9801), .Z(n9804) );
  AND U10490 ( .A(n9803), .B(n9804), .Z(n21993) );
  XOR U10491 ( .A(n9804), .B(n9803), .Z(n21988) );
  NAND U10492 ( .A(a[62]), .B(b[31]), .Z(n10168) );
  NAND U10493 ( .A(a[61]), .B(b[31]), .Z(n10162) );
  NAND U10494 ( .A(a[58]), .B(b[31]), .Z(n10146) );
  NAND U10495 ( .A(a[56]), .B(b[31]), .Z(n10134) );
  NAND U10496 ( .A(a[54]), .B(b[31]), .Z(n10122) );
  NAND U10497 ( .A(a[52]), .B(b[31]), .Z(n10110) );
  NAND U10498 ( .A(a[50]), .B(b[31]), .Z(n10098) );
  NAND U10499 ( .A(a[48]), .B(b[31]), .Z(n10086) );
  NAND U10500 ( .A(a[46]), .B(b[31]), .Z(n10074) );
  NAND U10501 ( .A(a[44]), .B(b[31]), .Z(n10062) );
  NAND U10502 ( .A(a[42]), .B(b[31]), .Z(n10050) );
  NAND U10503 ( .A(a[40]), .B(b[31]), .Z(n10038) );
  NAND U10504 ( .A(a[38]), .B(b[31]), .Z(n10026) );
  NAND U10505 ( .A(a[36]), .B(b[31]), .Z(n10014) );
  ANDN U10506 ( .B(b[31]), .A(n21703), .Z(n9946) );
  ANDN U10507 ( .B(b[31]), .A(n166), .Z(n9838) );
  ANDN U10508 ( .B(b[31]), .A(n21580), .Z(n9814) );
  NAND U10509 ( .A(b[32]), .B(a[1]), .Z(n9807) );
  AND U10510 ( .A(b[31]), .B(a[0]), .Z(n10569) );
  NANDN U10511 ( .A(n9807), .B(n10569), .Z(n9806) );
  NAND U10512 ( .A(a[2]), .B(b[31]), .Z(n9805) );
  AND U10513 ( .A(n9806), .B(n9805), .Z(n9813) );
  NANDN U10514 ( .A(n9807), .B(a[0]), .Z(n9808) );
  XNOR U10515 ( .A(a[2]), .B(n9808), .Z(n9809) );
  NAND U10516 ( .A(b[31]), .B(n9809), .Z(n10192) );
  AND U10517 ( .A(a[1]), .B(b[32]), .Z(n9810) );
  XNOR U10518 ( .A(n9811), .B(n9810), .Z(n10191) );
  NANDN U10519 ( .A(n10192), .B(n10191), .Z(n9812) );
  NANDN U10520 ( .A(n9813), .B(n9812), .Z(n9815) );
  NANDN U10521 ( .A(n9814), .B(n9815), .Z(n9819) );
  XOR U10522 ( .A(n9815), .B(n9814), .Z(n10196) );
  NANDN U10523 ( .A(n10196), .B(n10195), .Z(n9818) );
  NAND U10524 ( .A(n9819), .B(n9818), .Z(n9822) );
  XOR U10525 ( .A(n9821), .B(n9820), .Z(n9823) );
  OR U10526 ( .A(n9822), .B(n9823), .Z(n9825) );
  NAND U10527 ( .A(a[4]), .B(b[31]), .Z(n10204) );
  XOR U10528 ( .A(n9823), .B(n9822), .Z(n10203) );
  NANDN U10529 ( .A(n10204), .B(n10203), .Z(n9824) );
  NAND U10530 ( .A(n9825), .B(n9824), .Z(n9826) );
  ANDN U10531 ( .B(b[31]), .A(n164), .Z(n9827) );
  OR U10532 ( .A(n9826), .B(n9827), .Z(n9831) );
  XNOR U10533 ( .A(n9827), .B(n9826), .Z(n10207) );
  OR U10534 ( .A(n10207), .B(n10208), .Z(n9830) );
  AND U10535 ( .A(n9831), .B(n9830), .Z(n9835) );
  XOR U10536 ( .A(n9833), .B(n9832), .Z(n9834) );
  NANDN U10537 ( .A(n9835), .B(n9834), .Z(n9837) );
  XOR U10538 ( .A(n9835), .B(n9834), .Z(n10215) );
  ANDN U10539 ( .B(b[31]), .A(n165), .Z(n10216) );
  OR U10540 ( .A(n10215), .B(n10216), .Z(n9836) );
  AND U10541 ( .A(n9837), .B(n9836), .Z(n9839) );
  OR U10542 ( .A(n9838), .B(n9839), .Z(n9843) );
  XNOR U10543 ( .A(n9839), .B(n9838), .Z(n10220) );
  XNOR U10544 ( .A(n9841), .B(n9840), .Z(n10219) );
  OR U10545 ( .A(n10220), .B(n10219), .Z(n9842) );
  NAND U10546 ( .A(n9843), .B(n9842), .Z(n9846) );
  XOR U10547 ( .A(n9845), .B(n9844), .Z(n9847) );
  OR U10548 ( .A(n9846), .B(n9847), .Z(n9849) );
  NAND U10549 ( .A(a[8]), .B(b[31]), .Z(n10226) );
  XOR U10550 ( .A(n9847), .B(n9846), .Z(n10225) );
  NANDN U10551 ( .A(n10226), .B(n10225), .Z(n9848) );
  NAND U10552 ( .A(n9849), .B(n9848), .Z(n9852) );
  ANDN U10553 ( .B(b[31]), .A(n21615), .Z(n9853) );
  OR U10554 ( .A(n9852), .B(n9853), .Z(n9855) );
  XOR U10555 ( .A(n9853), .B(n9852), .Z(n10231) );
  NANDN U10556 ( .A(n10232), .B(n10231), .Z(n9854) );
  NAND U10557 ( .A(n9855), .B(n9854), .Z(n9858) );
  XNOR U10558 ( .A(n9857), .B(n9856), .Z(n9859) );
  OR U10559 ( .A(n9858), .B(n9859), .Z(n9861) );
  XNOR U10560 ( .A(n9859), .B(n9858), .Z(n10238) );
  NAND U10561 ( .A(a[10]), .B(b[31]), .Z(n10237) );
  OR U10562 ( .A(n10238), .B(n10237), .Z(n9860) );
  NAND U10563 ( .A(n9861), .B(n9860), .Z(n9864) );
  ANDN U10564 ( .B(b[31]), .A(n21164), .Z(n9865) );
  OR U10565 ( .A(n9864), .B(n9865), .Z(n9867) );
  XOR U10566 ( .A(n9865), .B(n9864), .Z(n10243) );
  NANDN U10567 ( .A(n10244), .B(n10243), .Z(n9866) );
  NAND U10568 ( .A(n9867), .B(n9866), .Z(n9870) );
  XNOR U10569 ( .A(n9869), .B(n9868), .Z(n9871) );
  OR U10570 ( .A(n9870), .B(n9871), .Z(n9873) );
  XNOR U10571 ( .A(n9871), .B(n9870), .Z(n10250) );
  NAND U10572 ( .A(a[12]), .B(b[31]), .Z(n10249) );
  OR U10573 ( .A(n10250), .B(n10249), .Z(n9872) );
  NAND U10574 ( .A(n9873), .B(n9872), .Z(n9876) );
  ANDN U10575 ( .B(b[31]), .A(n170), .Z(n9877) );
  OR U10576 ( .A(n9876), .B(n9877), .Z(n9879) );
  XOR U10577 ( .A(n9875), .B(n9874), .Z(n10256) );
  XOR U10578 ( .A(n9877), .B(n9876), .Z(n10255) );
  NANDN U10579 ( .A(n10256), .B(n10255), .Z(n9878) );
  NAND U10580 ( .A(n9879), .B(n9878), .Z(n9882) );
  XOR U10581 ( .A(n9881), .B(n9880), .Z(n9883) );
  OR U10582 ( .A(n9882), .B(n9883), .Z(n9885) );
  NAND U10583 ( .A(a[14]), .B(b[31]), .Z(n10262) );
  XOR U10584 ( .A(n9883), .B(n9882), .Z(n10261) );
  NANDN U10585 ( .A(n10262), .B(n10261), .Z(n9884) );
  NAND U10586 ( .A(n9885), .B(n9884), .Z(n9886) );
  ANDN U10587 ( .B(b[31]), .A(n172), .Z(n9887) );
  OR U10588 ( .A(n9886), .B(n9887), .Z(n9891) );
  XNOR U10589 ( .A(n9887), .B(n9886), .Z(n10268) );
  XOR U10590 ( .A(n9889), .B(n9888), .Z(n10267) );
  OR U10591 ( .A(n10268), .B(n10267), .Z(n9890) );
  NAND U10592 ( .A(n9891), .B(n9890), .Z(n9894) );
  XNOR U10593 ( .A(n9893), .B(n9892), .Z(n9895) );
  OR U10594 ( .A(n9894), .B(n9895), .Z(n9897) );
  XNOR U10595 ( .A(n9895), .B(n9894), .Z(n10274) );
  NAND U10596 ( .A(a[16]), .B(b[31]), .Z(n10273) );
  OR U10597 ( .A(n10274), .B(n10273), .Z(n9896) );
  NAND U10598 ( .A(n9897), .B(n9896), .Z(n9900) );
  ANDN U10599 ( .B(b[31]), .A(n174), .Z(n9901) );
  OR U10600 ( .A(n9900), .B(n9901), .Z(n9903) );
  XOR U10601 ( .A(n9901), .B(n9900), .Z(n10279) );
  NANDN U10602 ( .A(n10280), .B(n10279), .Z(n9902) );
  NAND U10603 ( .A(n9903), .B(n9902), .Z(n9906) );
  XNOR U10604 ( .A(n9905), .B(n9904), .Z(n9907) );
  OR U10605 ( .A(n9906), .B(n9907), .Z(n9909) );
  XNOR U10606 ( .A(n9907), .B(n9906), .Z(n10286) );
  NAND U10607 ( .A(a[18]), .B(b[31]), .Z(n10285) );
  OR U10608 ( .A(n10286), .B(n10285), .Z(n9908) );
  NAND U10609 ( .A(n9909), .B(n9908), .Z(n9912) );
  ANDN U10610 ( .B(b[31]), .A(n21670), .Z(n9913) );
  OR U10611 ( .A(n9912), .B(n9913), .Z(n9915) );
  XOR U10612 ( .A(n9911), .B(n9910), .Z(n10292) );
  XOR U10613 ( .A(n9913), .B(n9912), .Z(n10291) );
  NANDN U10614 ( .A(n10292), .B(n10291), .Z(n9914) );
  NAND U10615 ( .A(n9915), .B(n9914), .Z(n9918) );
  XNOR U10616 ( .A(n9917), .B(n9916), .Z(n9919) );
  OR U10617 ( .A(n9918), .B(n9919), .Z(n9921) );
  XNOR U10618 ( .A(n9919), .B(n9918), .Z(n10298) );
  NAND U10619 ( .A(a[20]), .B(b[31]), .Z(n10297) );
  OR U10620 ( .A(n10298), .B(n10297), .Z(n9920) );
  NAND U10621 ( .A(n9921), .B(n9920), .Z(n9924) );
  ANDN U10622 ( .B(b[31]), .A(n21681), .Z(n9925) );
  OR U10623 ( .A(n9924), .B(n9925), .Z(n9927) );
  XOR U10624 ( .A(n9923), .B(n9922), .Z(n10304) );
  XOR U10625 ( .A(n9925), .B(n9924), .Z(n10303) );
  NANDN U10626 ( .A(n10304), .B(n10303), .Z(n9926) );
  NAND U10627 ( .A(n9927), .B(n9926), .Z(n9930) );
  XNOR U10628 ( .A(n9929), .B(n9928), .Z(n9931) );
  OR U10629 ( .A(n9930), .B(n9931), .Z(n9933) );
  XNOR U10630 ( .A(n9931), .B(n9930), .Z(n10310) );
  NAND U10631 ( .A(a[22]), .B(b[31]), .Z(n10309) );
  OR U10632 ( .A(n10310), .B(n10309), .Z(n9932) );
  NAND U10633 ( .A(n9933), .B(n9932), .Z(n9936) );
  ANDN U10634 ( .B(b[31]), .A(n21692), .Z(n9937) );
  OR U10635 ( .A(n9936), .B(n9937), .Z(n9939) );
  XNOR U10636 ( .A(n9935), .B(n9934), .Z(n10316) );
  XNOR U10637 ( .A(n9937), .B(n9936), .Z(n10315) );
  OR U10638 ( .A(n10316), .B(n10315), .Z(n9938) );
  AND U10639 ( .A(n9939), .B(n9938), .Z(n9943) );
  XOR U10640 ( .A(n9941), .B(n9940), .Z(n9942) );
  NANDN U10641 ( .A(n9943), .B(n9942), .Z(n9945) );
  XOR U10642 ( .A(n9943), .B(n9942), .Z(n10321) );
  ANDN U10643 ( .B(b[31]), .A(n178), .Z(n10322) );
  OR U10644 ( .A(n10321), .B(n10322), .Z(n9944) );
  AND U10645 ( .A(n9945), .B(n9944), .Z(n9947) );
  OR U10646 ( .A(n9946), .B(n9947), .Z(n9951) );
  XNOR U10647 ( .A(n9947), .B(n9946), .Z(n10327) );
  OR U10648 ( .A(n10327), .B(n10328), .Z(n9950) );
  NAND U10649 ( .A(n9951), .B(n9950), .Z(n9954) );
  XOR U10650 ( .A(n9953), .B(n9952), .Z(n9955) );
  OR U10651 ( .A(n9954), .B(n9955), .Z(n9957) );
  XNOR U10652 ( .A(n9955), .B(n9954), .Z(n10336) );
  AND U10653 ( .A(b[31]), .B(a[26]), .Z(n10335) );
  NANDN U10654 ( .A(n10336), .B(n10335), .Z(n9956) );
  NAND U10655 ( .A(n9957), .B(n9956), .Z(n9958) );
  ANDN U10656 ( .B(b[31]), .A(n21716), .Z(n9959) );
  OR U10657 ( .A(n9958), .B(n9959), .Z(n9963) );
  XNOR U10658 ( .A(n9959), .B(n9958), .Z(n10339) );
  XOR U10659 ( .A(n9961), .B(n9960), .Z(n10340) );
  OR U10660 ( .A(n10339), .B(n10340), .Z(n9962) );
  NAND U10661 ( .A(n9963), .B(n9962), .Z(n9966) );
  XNOR U10662 ( .A(n9965), .B(n9964), .Z(n9967) );
  OR U10663 ( .A(n9966), .B(n9967), .Z(n9969) );
  XNOR U10664 ( .A(n9967), .B(n9966), .Z(n10346) );
  NAND U10665 ( .A(a[28]), .B(b[31]), .Z(n10345) );
  OR U10666 ( .A(n10346), .B(n10345), .Z(n9968) );
  NAND U10667 ( .A(n9969), .B(n9968), .Z(n9972) );
  ANDN U10668 ( .B(b[31]), .A(n21727), .Z(n9973) );
  OR U10669 ( .A(n9972), .B(n9973), .Z(n9975) );
  XOR U10670 ( .A(n9971), .B(n9970), .Z(n10352) );
  XOR U10671 ( .A(n9973), .B(n9972), .Z(n10351) );
  NANDN U10672 ( .A(n10352), .B(n10351), .Z(n9974) );
  NAND U10673 ( .A(n9975), .B(n9974), .Z(n9978) );
  XOR U10674 ( .A(n9977), .B(n9976), .Z(n9979) );
  OR U10675 ( .A(n9978), .B(n9979), .Z(n9981) );
  NAND U10676 ( .A(a[30]), .B(b[31]), .Z(n10358) );
  XOR U10677 ( .A(n9979), .B(n9978), .Z(n10357) );
  NANDN U10678 ( .A(n10358), .B(n10357), .Z(n9980) );
  NAND U10679 ( .A(n9981), .B(n9980), .Z(n9984) );
  ANDN U10680 ( .B(b[31]), .A(n21740), .Z(n9985) );
  OR U10681 ( .A(n9984), .B(n9985), .Z(n9987) );
  XOR U10682 ( .A(n9983), .B(n9982), .Z(n10364) );
  XOR U10683 ( .A(n9985), .B(n9984), .Z(n10363) );
  NANDN U10684 ( .A(n10364), .B(n10363), .Z(n9986) );
  NAND U10685 ( .A(n9987), .B(n9986), .Z(n9990) );
  XNOR U10686 ( .A(n9989), .B(n9988), .Z(n9991) );
  OR U10687 ( .A(n9990), .B(n9991), .Z(n9993) );
  XNOR U10688 ( .A(n9991), .B(n9990), .Z(n10370) );
  NAND U10689 ( .A(a[32]), .B(b[31]), .Z(n10369) );
  OR U10690 ( .A(n10370), .B(n10369), .Z(n9992) );
  NAND U10691 ( .A(n9993), .B(n9992), .Z(n9994) );
  ANDN U10692 ( .B(b[31]), .A(n21751), .Z(n9995) );
  OR U10693 ( .A(n9994), .B(n9995), .Z(n9999) );
  XOR U10694 ( .A(n9995), .B(n9994), .Z(n10375) );
  NAND U10695 ( .A(n10375), .B(n10376), .Z(n9998) );
  NAND U10696 ( .A(n9999), .B(n9998), .Z(n10003) );
  NAND U10697 ( .A(a[34]), .B(b[31]), .Z(n10002) );
  OR U10698 ( .A(n10003), .B(n10002), .Z(n10005) );
  XOR U10699 ( .A(n10001), .B(n10000), .Z(n10381) );
  XOR U10700 ( .A(n10003), .B(n10002), .Z(n10382) );
  NAND U10701 ( .A(n10381), .B(n10382), .Z(n10004) );
  NAND U10702 ( .A(n10005), .B(n10004), .Z(n10009) );
  XOR U10703 ( .A(n10007), .B(n10006), .Z(n10008) );
  NAND U10704 ( .A(n10009), .B(n10008), .Z(n10011) );
  XNOR U10705 ( .A(n10009), .B(n10008), .Z(n10388) );
  NAND U10706 ( .A(a[35]), .B(b[31]), .Z(n10387) );
  OR U10707 ( .A(n10388), .B(n10387), .Z(n10010) );
  NAND U10708 ( .A(n10011), .B(n10010), .Z(n10015) );
  NANDN U10709 ( .A(n10014), .B(n10015), .Z(n10017) );
  XNOR U10710 ( .A(n10013), .B(n10012), .Z(n10394) );
  XNOR U10711 ( .A(n10015), .B(n10014), .Z(n10393) );
  NANDN U10712 ( .A(n10394), .B(n10393), .Z(n10016) );
  NAND U10713 ( .A(n10017), .B(n10016), .Z(n10021) );
  XOR U10714 ( .A(n10019), .B(n10018), .Z(n10020) );
  NAND U10715 ( .A(n10021), .B(n10020), .Z(n10023) );
  XNOR U10716 ( .A(n10021), .B(n10020), .Z(n10400) );
  NAND U10717 ( .A(a[37]), .B(b[31]), .Z(n10399) );
  OR U10718 ( .A(n10400), .B(n10399), .Z(n10022) );
  NAND U10719 ( .A(n10023), .B(n10022), .Z(n10027) );
  NANDN U10720 ( .A(n10026), .B(n10027), .Z(n10029) );
  XNOR U10721 ( .A(n10025), .B(n10024), .Z(n10406) );
  XNOR U10722 ( .A(n10027), .B(n10026), .Z(n10405) );
  NANDN U10723 ( .A(n10406), .B(n10405), .Z(n10028) );
  NAND U10724 ( .A(n10029), .B(n10028), .Z(n10033) );
  XOR U10725 ( .A(n10031), .B(n10030), .Z(n10032) );
  NAND U10726 ( .A(n10033), .B(n10032), .Z(n10035) );
  XNOR U10727 ( .A(n10033), .B(n10032), .Z(n10412) );
  NAND U10728 ( .A(a[39]), .B(b[31]), .Z(n10411) );
  OR U10729 ( .A(n10412), .B(n10411), .Z(n10034) );
  NAND U10730 ( .A(n10035), .B(n10034), .Z(n10039) );
  NANDN U10731 ( .A(n10038), .B(n10039), .Z(n10041) );
  XNOR U10732 ( .A(n10037), .B(n10036), .Z(n10418) );
  XNOR U10733 ( .A(n10039), .B(n10038), .Z(n10417) );
  NANDN U10734 ( .A(n10418), .B(n10417), .Z(n10040) );
  NAND U10735 ( .A(n10041), .B(n10040), .Z(n10045) );
  XOR U10736 ( .A(n10043), .B(n10042), .Z(n10044) );
  NAND U10737 ( .A(n10045), .B(n10044), .Z(n10047) );
  XNOR U10738 ( .A(n10045), .B(n10044), .Z(n10424) );
  NAND U10739 ( .A(a[41]), .B(b[31]), .Z(n10423) );
  OR U10740 ( .A(n10424), .B(n10423), .Z(n10046) );
  NAND U10741 ( .A(n10047), .B(n10046), .Z(n10051) );
  NANDN U10742 ( .A(n10050), .B(n10051), .Z(n10053) );
  XNOR U10743 ( .A(n10049), .B(n10048), .Z(n10430) );
  XNOR U10744 ( .A(n10051), .B(n10050), .Z(n10429) );
  NANDN U10745 ( .A(n10430), .B(n10429), .Z(n10052) );
  NAND U10746 ( .A(n10053), .B(n10052), .Z(n10057) );
  XOR U10747 ( .A(n10055), .B(n10054), .Z(n10056) );
  NAND U10748 ( .A(n10057), .B(n10056), .Z(n10059) );
  XNOR U10749 ( .A(n10057), .B(n10056), .Z(n10436) );
  NAND U10750 ( .A(a[43]), .B(b[31]), .Z(n10435) );
  OR U10751 ( .A(n10436), .B(n10435), .Z(n10058) );
  NAND U10752 ( .A(n10059), .B(n10058), .Z(n10063) );
  NANDN U10753 ( .A(n10062), .B(n10063), .Z(n10065) );
  XNOR U10754 ( .A(n10061), .B(n10060), .Z(n10442) );
  XNOR U10755 ( .A(n10063), .B(n10062), .Z(n10441) );
  NANDN U10756 ( .A(n10442), .B(n10441), .Z(n10064) );
  NAND U10757 ( .A(n10065), .B(n10064), .Z(n10069) );
  XOR U10758 ( .A(n10067), .B(n10066), .Z(n10068) );
  NAND U10759 ( .A(n10069), .B(n10068), .Z(n10071) );
  XNOR U10760 ( .A(n10069), .B(n10068), .Z(n10448) );
  NAND U10761 ( .A(a[45]), .B(b[31]), .Z(n10447) );
  OR U10762 ( .A(n10448), .B(n10447), .Z(n10070) );
  NAND U10763 ( .A(n10071), .B(n10070), .Z(n10075) );
  NANDN U10764 ( .A(n10074), .B(n10075), .Z(n10077) );
  XNOR U10765 ( .A(n10073), .B(n10072), .Z(n10454) );
  XNOR U10766 ( .A(n10075), .B(n10074), .Z(n10453) );
  NANDN U10767 ( .A(n10454), .B(n10453), .Z(n10076) );
  NAND U10768 ( .A(n10077), .B(n10076), .Z(n10081) );
  XOR U10769 ( .A(n10079), .B(n10078), .Z(n10080) );
  NAND U10770 ( .A(n10081), .B(n10080), .Z(n10083) );
  XNOR U10771 ( .A(n10081), .B(n10080), .Z(n10460) );
  NAND U10772 ( .A(a[47]), .B(b[31]), .Z(n10459) );
  OR U10773 ( .A(n10460), .B(n10459), .Z(n10082) );
  NAND U10774 ( .A(n10083), .B(n10082), .Z(n10087) );
  NANDN U10775 ( .A(n10086), .B(n10087), .Z(n10089) );
  XNOR U10776 ( .A(n10085), .B(n10084), .Z(n10466) );
  XNOR U10777 ( .A(n10087), .B(n10086), .Z(n10465) );
  NANDN U10778 ( .A(n10466), .B(n10465), .Z(n10088) );
  NAND U10779 ( .A(n10089), .B(n10088), .Z(n10093) );
  XOR U10780 ( .A(n10091), .B(n10090), .Z(n10092) );
  NAND U10781 ( .A(n10093), .B(n10092), .Z(n10095) );
  XNOR U10782 ( .A(n10093), .B(n10092), .Z(n10472) );
  NAND U10783 ( .A(a[49]), .B(b[31]), .Z(n10471) );
  OR U10784 ( .A(n10472), .B(n10471), .Z(n10094) );
  NAND U10785 ( .A(n10095), .B(n10094), .Z(n10099) );
  NANDN U10786 ( .A(n10098), .B(n10099), .Z(n10101) );
  XNOR U10787 ( .A(n10097), .B(n10096), .Z(n10478) );
  XNOR U10788 ( .A(n10099), .B(n10098), .Z(n10477) );
  NANDN U10789 ( .A(n10478), .B(n10477), .Z(n10100) );
  NAND U10790 ( .A(n10101), .B(n10100), .Z(n10105) );
  XOR U10791 ( .A(n10103), .B(n10102), .Z(n10104) );
  NAND U10792 ( .A(n10105), .B(n10104), .Z(n10107) );
  XNOR U10793 ( .A(n10105), .B(n10104), .Z(n10484) );
  NAND U10794 ( .A(a[51]), .B(b[31]), .Z(n10483) );
  OR U10795 ( .A(n10484), .B(n10483), .Z(n10106) );
  NAND U10796 ( .A(n10107), .B(n10106), .Z(n10111) );
  NANDN U10797 ( .A(n10110), .B(n10111), .Z(n10113) );
  XNOR U10798 ( .A(n10109), .B(n10108), .Z(n10490) );
  XNOR U10799 ( .A(n10111), .B(n10110), .Z(n10489) );
  NANDN U10800 ( .A(n10490), .B(n10489), .Z(n10112) );
  NAND U10801 ( .A(n10113), .B(n10112), .Z(n10117) );
  XOR U10802 ( .A(n10115), .B(n10114), .Z(n10116) );
  NAND U10803 ( .A(n10117), .B(n10116), .Z(n10119) );
  XNOR U10804 ( .A(n10117), .B(n10116), .Z(n10496) );
  NAND U10805 ( .A(a[53]), .B(b[31]), .Z(n10495) );
  OR U10806 ( .A(n10496), .B(n10495), .Z(n10118) );
  NAND U10807 ( .A(n10119), .B(n10118), .Z(n10123) );
  NANDN U10808 ( .A(n10122), .B(n10123), .Z(n10125) );
  XNOR U10809 ( .A(n10121), .B(n10120), .Z(n10502) );
  XNOR U10810 ( .A(n10123), .B(n10122), .Z(n10501) );
  NANDN U10811 ( .A(n10502), .B(n10501), .Z(n10124) );
  NAND U10812 ( .A(n10125), .B(n10124), .Z(n10129) );
  XOR U10813 ( .A(n10127), .B(n10126), .Z(n10128) );
  NAND U10814 ( .A(n10129), .B(n10128), .Z(n10131) );
  XNOR U10815 ( .A(n10129), .B(n10128), .Z(n10508) );
  NAND U10816 ( .A(a[55]), .B(b[31]), .Z(n10507) );
  OR U10817 ( .A(n10508), .B(n10507), .Z(n10130) );
  NAND U10818 ( .A(n10131), .B(n10130), .Z(n10135) );
  NANDN U10819 ( .A(n10134), .B(n10135), .Z(n10137) );
  XNOR U10820 ( .A(n10133), .B(n10132), .Z(n10514) );
  XNOR U10821 ( .A(n10135), .B(n10134), .Z(n10513) );
  NANDN U10822 ( .A(n10514), .B(n10513), .Z(n10136) );
  NAND U10823 ( .A(n10137), .B(n10136), .Z(n10141) );
  XOR U10824 ( .A(n10139), .B(n10138), .Z(n10140) );
  NAND U10825 ( .A(n10141), .B(n10140), .Z(n10143) );
  XNOR U10826 ( .A(n10141), .B(n10140), .Z(n10520) );
  NAND U10827 ( .A(a[57]), .B(b[31]), .Z(n10519) );
  OR U10828 ( .A(n10520), .B(n10519), .Z(n10142) );
  NAND U10829 ( .A(n10143), .B(n10142), .Z(n10147) );
  NANDN U10830 ( .A(n10146), .B(n10147), .Z(n10149) );
  XNOR U10831 ( .A(n10145), .B(n10144), .Z(n10526) );
  XNOR U10832 ( .A(n10147), .B(n10146), .Z(n10525) );
  NANDN U10833 ( .A(n10526), .B(n10525), .Z(n10148) );
  NAND U10834 ( .A(n10149), .B(n10148), .Z(n10152) );
  AND U10835 ( .A(b[31]), .B(a[59]), .Z(n10153) );
  XOR U10836 ( .A(n10151), .B(n10150), .Z(n10532) );
  XOR U10837 ( .A(n10153), .B(n10152), .Z(n10531) );
  NAND U10838 ( .A(a[60]), .B(b[31]), .Z(n10156) );
  OR U10839 ( .A(n10157), .B(n10156), .Z(n10159) );
  XNOR U10840 ( .A(n10155), .B(n10154), .Z(n10538) );
  XOR U10841 ( .A(n10157), .B(n10156), .Z(n10537) );
  NANDN U10842 ( .A(n10538), .B(n10537), .Z(n10158) );
  NAND U10843 ( .A(n10159), .B(n10158), .Z(n10163) );
  NANDN U10844 ( .A(n10162), .B(n10163), .Z(n10165) );
  XOR U10845 ( .A(n10161), .B(n10160), .Z(n10543) );
  XNOR U10846 ( .A(n10163), .B(n10162), .Z(n10544) );
  NAND U10847 ( .A(n10543), .B(n10544), .Z(n10164) );
  NAND U10848 ( .A(n10165), .B(n10164), .Z(n10169) );
  NANDN U10849 ( .A(n10168), .B(n10169), .Z(n10171) );
  XNOR U10850 ( .A(n10167), .B(n10166), .Z(n10550) );
  XNOR U10851 ( .A(n10169), .B(n10168), .Z(n10549) );
  NANDN U10852 ( .A(n10550), .B(n10549), .Z(n10170) );
  NAND U10853 ( .A(n10171), .B(n10170), .Z(n10174) );
  XOR U10854 ( .A(n10173), .B(n10172), .Z(n10175) );
  AND U10855 ( .A(b[31]), .B(a[63]), .Z(n10179) );
  XOR U10856 ( .A(n10175), .B(n10174), .Z(n10178) );
  XNOR U10857 ( .A(n10177), .B(n10176), .Z(n10556) );
  OR U10858 ( .A(n10555), .B(n10556), .Z(n21989) );
  NANDN U10859 ( .A(n21988), .B(n21989), .Z(n21991) );
  XOR U10860 ( .A(n10179), .B(n10178), .Z(n10560) );
  NAND U10861 ( .A(a[36]), .B(b[30]), .Z(n10389) );
  ANDN U10862 ( .B(b[30]), .A(n21727), .Z(n10347) );
  NAND U10863 ( .A(a[27]), .B(b[30]), .Z(n10334) );
  ANDN U10864 ( .B(b[30]), .A(n166), .Z(n10213) );
  ANDN U10865 ( .B(b[30]), .A(n21580), .Z(n10189) );
  NAND U10866 ( .A(b[31]), .B(a[1]), .Z(n10182) );
  AND U10867 ( .A(b[30]), .B(a[0]), .Z(n10948) );
  NANDN U10868 ( .A(n10182), .B(n10948), .Z(n10181) );
  NAND U10869 ( .A(a[2]), .B(b[30]), .Z(n10180) );
  AND U10870 ( .A(n10181), .B(n10180), .Z(n10188) );
  NANDN U10871 ( .A(n10182), .B(a[0]), .Z(n10183) );
  XNOR U10872 ( .A(a[2]), .B(n10183), .Z(n10184) );
  NAND U10873 ( .A(b[30]), .B(n10184), .Z(n10575) );
  AND U10874 ( .A(a[1]), .B(b[31]), .Z(n10185) );
  XNOR U10875 ( .A(n10186), .B(n10185), .Z(n10574) );
  NANDN U10876 ( .A(n10575), .B(n10574), .Z(n10187) );
  NANDN U10877 ( .A(n10188), .B(n10187), .Z(n10190) );
  NANDN U10878 ( .A(n10189), .B(n10190), .Z(n10194) );
  XOR U10879 ( .A(n10190), .B(n10189), .Z(n10579) );
  NANDN U10880 ( .A(n10579), .B(n10578), .Z(n10193) );
  NAND U10881 ( .A(n10194), .B(n10193), .Z(n10198) );
  XOR U10882 ( .A(n10196), .B(n10195), .Z(n10197) );
  NANDN U10883 ( .A(n10198), .B(n10197), .Z(n10200) );
  NAND U10884 ( .A(a[4]), .B(b[30]), .Z(n10584) );
  NANDN U10885 ( .A(n10584), .B(n10585), .Z(n10199) );
  NAND U10886 ( .A(n10200), .B(n10199), .Z(n10201) );
  ANDN U10887 ( .B(b[30]), .A(n164), .Z(n10202) );
  OR U10888 ( .A(n10201), .B(n10202), .Z(n10206) );
  XNOR U10889 ( .A(n10202), .B(n10201), .Z(n10590) );
  OR U10890 ( .A(n10590), .B(n10591), .Z(n10205) );
  AND U10891 ( .A(n10206), .B(n10205), .Z(n10210) );
  XOR U10892 ( .A(n10208), .B(n10207), .Z(n10209) );
  NANDN U10893 ( .A(n10210), .B(n10209), .Z(n10212) );
  XOR U10894 ( .A(n10210), .B(n10209), .Z(n10598) );
  ANDN U10895 ( .B(b[30]), .A(n165), .Z(n10599) );
  OR U10896 ( .A(n10598), .B(n10599), .Z(n10211) );
  AND U10897 ( .A(n10212), .B(n10211), .Z(n10214) );
  OR U10898 ( .A(n10213), .B(n10214), .Z(n10218) );
  XNOR U10899 ( .A(n10214), .B(n10213), .Z(n10603) );
  XNOR U10900 ( .A(n10216), .B(n10215), .Z(n10602) );
  OR U10901 ( .A(n10603), .B(n10602), .Z(n10217) );
  NAND U10902 ( .A(n10218), .B(n10217), .Z(n10221) );
  XOR U10903 ( .A(n10220), .B(n10219), .Z(n10222) );
  OR U10904 ( .A(n10221), .B(n10222), .Z(n10224) );
  NAND U10905 ( .A(a[8]), .B(b[30]), .Z(n10611) );
  XOR U10906 ( .A(n10222), .B(n10221), .Z(n10610) );
  NANDN U10907 ( .A(n10611), .B(n10610), .Z(n10223) );
  NAND U10908 ( .A(n10224), .B(n10223), .Z(n10227) );
  ANDN U10909 ( .B(b[30]), .A(n21615), .Z(n10228) );
  OR U10910 ( .A(n10227), .B(n10228), .Z(n10230) );
  XOR U10911 ( .A(n10228), .B(n10227), .Z(n10614) );
  NANDN U10912 ( .A(n10615), .B(n10614), .Z(n10229) );
  NAND U10913 ( .A(n10230), .B(n10229), .Z(n10233) );
  XNOR U10914 ( .A(n10232), .B(n10231), .Z(n10234) );
  OR U10915 ( .A(n10233), .B(n10234), .Z(n10236) );
  XNOR U10916 ( .A(n10234), .B(n10233), .Z(n10621) );
  NAND U10917 ( .A(a[10]), .B(b[30]), .Z(n10620) );
  OR U10918 ( .A(n10621), .B(n10620), .Z(n10235) );
  NAND U10919 ( .A(n10236), .B(n10235), .Z(n10239) );
  ANDN U10920 ( .B(b[30]), .A(n21164), .Z(n10240) );
  OR U10921 ( .A(n10239), .B(n10240), .Z(n10242) );
  XOR U10922 ( .A(n10238), .B(n10237), .Z(n10627) );
  XOR U10923 ( .A(n10240), .B(n10239), .Z(n10626) );
  NANDN U10924 ( .A(n10627), .B(n10626), .Z(n10241) );
  NAND U10925 ( .A(n10242), .B(n10241), .Z(n10245) );
  XNOR U10926 ( .A(n10244), .B(n10243), .Z(n10246) );
  OR U10927 ( .A(n10245), .B(n10246), .Z(n10248) );
  XNOR U10928 ( .A(n10246), .B(n10245), .Z(n10633) );
  NAND U10929 ( .A(a[12]), .B(b[30]), .Z(n10632) );
  OR U10930 ( .A(n10633), .B(n10632), .Z(n10247) );
  NAND U10931 ( .A(n10248), .B(n10247), .Z(n10251) );
  ANDN U10932 ( .B(b[30]), .A(n170), .Z(n10252) );
  OR U10933 ( .A(n10251), .B(n10252), .Z(n10254) );
  XOR U10934 ( .A(n10250), .B(n10249), .Z(n10639) );
  XOR U10935 ( .A(n10252), .B(n10251), .Z(n10638) );
  NANDN U10936 ( .A(n10639), .B(n10638), .Z(n10253) );
  NAND U10937 ( .A(n10254), .B(n10253), .Z(n10257) );
  XNOR U10938 ( .A(n10256), .B(n10255), .Z(n10258) );
  OR U10939 ( .A(n10257), .B(n10258), .Z(n10260) );
  XNOR U10940 ( .A(n10258), .B(n10257), .Z(n10645) );
  NAND U10941 ( .A(a[14]), .B(b[30]), .Z(n10644) );
  OR U10942 ( .A(n10645), .B(n10644), .Z(n10259) );
  NAND U10943 ( .A(n10260), .B(n10259), .Z(n10263) );
  ANDN U10944 ( .B(b[30]), .A(n172), .Z(n10264) );
  OR U10945 ( .A(n10263), .B(n10264), .Z(n10266) );
  XOR U10946 ( .A(n10264), .B(n10263), .Z(n10650) );
  NANDN U10947 ( .A(n10651), .B(n10650), .Z(n10265) );
  NAND U10948 ( .A(n10266), .B(n10265), .Z(n10269) );
  XOR U10949 ( .A(n10268), .B(n10267), .Z(n10270) );
  OR U10950 ( .A(n10269), .B(n10270), .Z(n10272) );
  NAND U10951 ( .A(a[16]), .B(b[30]), .Z(n10657) );
  XOR U10952 ( .A(n10270), .B(n10269), .Z(n10656) );
  NANDN U10953 ( .A(n10657), .B(n10656), .Z(n10271) );
  NAND U10954 ( .A(n10272), .B(n10271), .Z(n10275) );
  ANDN U10955 ( .B(b[30]), .A(n174), .Z(n10276) );
  OR U10956 ( .A(n10275), .B(n10276), .Z(n10278) );
  XOR U10957 ( .A(n10274), .B(n10273), .Z(n10663) );
  XOR U10958 ( .A(n10276), .B(n10275), .Z(n10662) );
  NANDN U10959 ( .A(n10663), .B(n10662), .Z(n10277) );
  NAND U10960 ( .A(n10278), .B(n10277), .Z(n10281) );
  XNOR U10961 ( .A(n10280), .B(n10279), .Z(n10282) );
  OR U10962 ( .A(n10281), .B(n10282), .Z(n10284) );
  XNOR U10963 ( .A(n10282), .B(n10281), .Z(n10669) );
  NAND U10964 ( .A(a[18]), .B(b[30]), .Z(n10668) );
  OR U10965 ( .A(n10669), .B(n10668), .Z(n10283) );
  NAND U10966 ( .A(n10284), .B(n10283), .Z(n10287) );
  ANDN U10967 ( .B(b[30]), .A(n21670), .Z(n10288) );
  OR U10968 ( .A(n10287), .B(n10288), .Z(n10290) );
  XOR U10969 ( .A(n10286), .B(n10285), .Z(n10675) );
  XOR U10970 ( .A(n10288), .B(n10287), .Z(n10674) );
  NANDN U10971 ( .A(n10675), .B(n10674), .Z(n10289) );
  NAND U10972 ( .A(n10290), .B(n10289), .Z(n10293) );
  XNOR U10973 ( .A(n10292), .B(n10291), .Z(n10294) );
  OR U10974 ( .A(n10293), .B(n10294), .Z(n10296) );
  XNOR U10975 ( .A(n10294), .B(n10293), .Z(n10681) );
  NAND U10976 ( .A(a[20]), .B(b[30]), .Z(n10680) );
  OR U10977 ( .A(n10681), .B(n10680), .Z(n10295) );
  NAND U10978 ( .A(n10296), .B(n10295), .Z(n10299) );
  ANDN U10979 ( .B(b[30]), .A(n21681), .Z(n10300) );
  OR U10980 ( .A(n10299), .B(n10300), .Z(n10302) );
  XOR U10981 ( .A(n10298), .B(n10297), .Z(n10687) );
  XOR U10982 ( .A(n10300), .B(n10299), .Z(n10686) );
  NANDN U10983 ( .A(n10687), .B(n10686), .Z(n10301) );
  NAND U10984 ( .A(n10302), .B(n10301), .Z(n10305) );
  XNOR U10985 ( .A(n10304), .B(n10303), .Z(n10306) );
  OR U10986 ( .A(n10305), .B(n10306), .Z(n10308) );
  XNOR U10987 ( .A(n10306), .B(n10305), .Z(n10693) );
  NAND U10988 ( .A(a[22]), .B(b[30]), .Z(n10692) );
  OR U10989 ( .A(n10693), .B(n10692), .Z(n10307) );
  NAND U10990 ( .A(n10308), .B(n10307), .Z(n10311) );
  ANDN U10991 ( .B(b[30]), .A(n21692), .Z(n10312) );
  OR U10992 ( .A(n10311), .B(n10312), .Z(n10314) );
  XOR U10993 ( .A(n10310), .B(n10309), .Z(n10699) );
  XOR U10994 ( .A(n10312), .B(n10311), .Z(n10698) );
  NANDN U10995 ( .A(n10699), .B(n10698), .Z(n10313) );
  NAND U10996 ( .A(n10314), .B(n10313), .Z(n10317) );
  XOR U10997 ( .A(n10316), .B(n10315), .Z(n10318) );
  OR U10998 ( .A(n10317), .B(n10318), .Z(n10320) );
  NAND U10999 ( .A(a[24]), .B(b[30]), .Z(n10705) );
  XOR U11000 ( .A(n10318), .B(n10317), .Z(n10704) );
  NANDN U11001 ( .A(n10705), .B(n10704), .Z(n10319) );
  NAND U11002 ( .A(n10320), .B(n10319), .Z(n10323) );
  ANDN U11003 ( .B(b[30]), .A(n21703), .Z(n10324) );
  OR U11004 ( .A(n10323), .B(n10324), .Z(n10326) );
  XNOR U11005 ( .A(n10322), .B(n10321), .Z(n10711) );
  XNOR U11006 ( .A(n10324), .B(n10323), .Z(n10710) );
  OR U11007 ( .A(n10711), .B(n10710), .Z(n10325) );
  AND U11008 ( .A(n10326), .B(n10325), .Z(n10330) );
  XOR U11009 ( .A(n10328), .B(n10327), .Z(n10329) );
  NANDN U11010 ( .A(n10330), .B(n10329), .Z(n10332) );
  XOR U11011 ( .A(n10330), .B(n10329), .Z(n10718) );
  ANDN U11012 ( .B(b[30]), .A(n179), .Z(n10719) );
  OR U11013 ( .A(n10718), .B(n10719), .Z(n10331) );
  NAND U11014 ( .A(n10332), .B(n10331), .Z(n10333) );
  OR U11015 ( .A(n10334), .B(n10333), .Z(n10338) );
  XNOR U11016 ( .A(n10334), .B(n10333), .Z(n10723) );
  XOR U11017 ( .A(n10336), .B(n10335), .Z(n10722) );
  OR U11018 ( .A(n10723), .B(n10722), .Z(n10337) );
  NAND U11019 ( .A(n10338), .B(n10337), .Z(n10341) );
  XOR U11020 ( .A(n10340), .B(n10339), .Z(n10342) );
  NANDN U11021 ( .A(n10341), .B(n10342), .Z(n10344) );
  XOR U11022 ( .A(n10342), .B(n10341), .Z(n10730) );
  ANDN U11023 ( .B(b[30]), .A(n180), .Z(n10731) );
  OR U11024 ( .A(n10730), .B(n10731), .Z(n10343) );
  AND U11025 ( .A(n10344), .B(n10343), .Z(n10348) );
  OR U11026 ( .A(n10347), .B(n10348), .Z(n10350) );
  XOR U11027 ( .A(n10346), .B(n10345), .Z(n10735) );
  XOR U11028 ( .A(n10348), .B(n10347), .Z(n10734) );
  NANDN U11029 ( .A(n10735), .B(n10734), .Z(n10349) );
  NAND U11030 ( .A(n10350), .B(n10349), .Z(n10353) );
  XNOR U11031 ( .A(n10352), .B(n10351), .Z(n10354) );
  OR U11032 ( .A(n10353), .B(n10354), .Z(n10356) );
  XNOR U11033 ( .A(n10354), .B(n10353), .Z(n10741) );
  NAND U11034 ( .A(a[30]), .B(b[30]), .Z(n10740) );
  OR U11035 ( .A(n10741), .B(n10740), .Z(n10355) );
  NAND U11036 ( .A(n10356), .B(n10355), .Z(n10359) );
  ANDN U11037 ( .B(b[30]), .A(n21740), .Z(n10360) );
  OR U11038 ( .A(n10359), .B(n10360), .Z(n10362) );
  XOR U11039 ( .A(n10360), .B(n10359), .Z(n10746) );
  NANDN U11040 ( .A(n10747), .B(n10746), .Z(n10361) );
  NAND U11041 ( .A(n10362), .B(n10361), .Z(n10365) );
  XNOR U11042 ( .A(n10364), .B(n10363), .Z(n10366) );
  OR U11043 ( .A(n10365), .B(n10366), .Z(n10368) );
  XNOR U11044 ( .A(n10366), .B(n10365), .Z(n10753) );
  NAND U11045 ( .A(a[32]), .B(b[30]), .Z(n10752) );
  OR U11046 ( .A(n10753), .B(n10752), .Z(n10367) );
  NAND U11047 ( .A(n10368), .B(n10367), .Z(n10371) );
  ANDN U11048 ( .B(b[30]), .A(n21751), .Z(n10372) );
  OR U11049 ( .A(n10371), .B(n10372), .Z(n10374) );
  XOR U11050 ( .A(n10370), .B(n10369), .Z(n10759) );
  XOR U11051 ( .A(n10372), .B(n10371), .Z(n10758) );
  NANDN U11052 ( .A(n10759), .B(n10758), .Z(n10373) );
  NAND U11053 ( .A(n10374), .B(n10373), .Z(n10378) );
  AND U11054 ( .A(b[30]), .B(a[34]), .Z(n10377) );
  NANDN U11055 ( .A(n10378), .B(n10377), .Z(n10380) );
  XNOR U11056 ( .A(n10378), .B(n10377), .Z(n10766) );
  NANDN U11057 ( .A(n10767), .B(n10766), .Z(n10379) );
  NAND U11058 ( .A(n10380), .B(n10379), .Z(n10384) );
  XOR U11059 ( .A(n10382), .B(n10381), .Z(n10383) );
  NAND U11060 ( .A(n10384), .B(n10383), .Z(n10386) );
  XNOR U11061 ( .A(n10384), .B(n10383), .Z(n10771) );
  NAND U11062 ( .A(a[35]), .B(b[30]), .Z(n10770) );
  OR U11063 ( .A(n10771), .B(n10770), .Z(n10385) );
  NAND U11064 ( .A(n10386), .B(n10385), .Z(n10390) );
  NANDN U11065 ( .A(n10389), .B(n10390), .Z(n10392) );
  XOR U11066 ( .A(n10388), .B(n10387), .Z(n10776) );
  XNOR U11067 ( .A(n10390), .B(n10389), .Z(n10777) );
  NAND U11068 ( .A(n10776), .B(n10777), .Z(n10391) );
  NAND U11069 ( .A(n10392), .B(n10391), .Z(n10395) );
  AND U11070 ( .A(b[30]), .B(a[37]), .Z(n10396) );
  OR U11071 ( .A(n10395), .B(n10396), .Z(n10398) );
  XNOR U11072 ( .A(n10394), .B(n10393), .Z(n10783) );
  XOR U11073 ( .A(n10396), .B(n10395), .Z(n10782) );
  NANDN U11074 ( .A(n10783), .B(n10782), .Z(n10397) );
  NAND U11075 ( .A(n10398), .B(n10397), .Z(n10402) );
  NAND U11076 ( .A(a[38]), .B(b[30]), .Z(n10401) );
  OR U11077 ( .A(n10402), .B(n10401), .Z(n10404) );
  XOR U11078 ( .A(n10400), .B(n10399), .Z(n10788) );
  XOR U11079 ( .A(n10402), .B(n10401), .Z(n10789) );
  NAND U11080 ( .A(n10788), .B(n10789), .Z(n10403) );
  NAND U11081 ( .A(n10404), .B(n10403), .Z(n10407) );
  AND U11082 ( .A(b[30]), .B(a[39]), .Z(n10408) );
  OR U11083 ( .A(n10407), .B(n10408), .Z(n10410) );
  XNOR U11084 ( .A(n10406), .B(n10405), .Z(n10795) );
  XOR U11085 ( .A(n10408), .B(n10407), .Z(n10794) );
  NANDN U11086 ( .A(n10795), .B(n10794), .Z(n10409) );
  NAND U11087 ( .A(n10410), .B(n10409), .Z(n10414) );
  NAND U11088 ( .A(a[40]), .B(b[30]), .Z(n10413) );
  OR U11089 ( .A(n10414), .B(n10413), .Z(n10416) );
  XOR U11090 ( .A(n10412), .B(n10411), .Z(n10800) );
  XOR U11091 ( .A(n10414), .B(n10413), .Z(n10801) );
  NAND U11092 ( .A(n10800), .B(n10801), .Z(n10415) );
  NAND U11093 ( .A(n10416), .B(n10415), .Z(n10419) );
  AND U11094 ( .A(b[30]), .B(a[41]), .Z(n10420) );
  OR U11095 ( .A(n10419), .B(n10420), .Z(n10422) );
  XNOR U11096 ( .A(n10418), .B(n10417), .Z(n10807) );
  XOR U11097 ( .A(n10420), .B(n10419), .Z(n10806) );
  NANDN U11098 ( .A(n10807), .B(n10806), .Z(n10421) );
  NAND U11099 ( .A(n10422), .B(n10421), .Z(n10426) );
  NAND U11100 ( .A(a[42]), .B(b[30]), .Z(n10425) );
  OR U11101 ( .A(n10426), .B(n10425), .Z(n10428) );
  XOR U11102 ( .A(n10424), .B(n10423), .Z(n10812) );
  XOR U11103 ( .A(n10426), .B(n10425), .Z(n10813) );
  NAND U11104 ( .A(n10812), .B(n10813), .Z(n10427) );
  NAND U11105 ( .A(n10428), .B(n10427), .Z(n10431) );
  AND U11106 ( .A(b[30]), .B(a[43]), .Z(n10432) );
  OR U11107 ( .A(n10431), .B(n10432), .Z(n10434) );
  XNOR U11108 ( .A(n10430), .B(n10429), .Z(n10819) );
  XOR U11109 ( .A(n10432), .B(n10431), .Z(n10818) );
  NANDN U11110 ( .A(n10819), .B(n10818), .Z(n10433) );
  NAND U11111 ( .A(n10434), .B(n10433), .Z(n10438) );
  NAND U11112 ( .A(a[44]), .B(b[30]), .Z(n10437) );
  OR U11113 ( .A(n10438), .B(n10437), .Z(n10440) );
  XOR U11114 ( .A(n10436), .B(n10435), .Z(n10824) );
  XOR U11115 ( .A(n10438), .B(n10437), .Z(n10825) );
  NAND U11116 ( .A(n10824), .B(n10825), .Z(n10439) );
  NAND U11117 ( .A(n10440), .B(n10439), .Z(n10443) );
  AND U11118 ( .A(b[30]), .B(a[45]), .Z(n10444) );
  OR U11119 ( .A(n10443), .B(n10444), .Z(n10446) );
  XNOR U11120 ( .A(n10442), .B(n10441), .Z(n10831) );
  XOR U11121 ( .A(n10444), .B(n10443), .Z(n10830) );
  NANDN U11122 ( .A(n10831), .B(n10830), .Z(n10445) );
  NAND U11123 ( .A(n10446), .B(n10445), .Z(n10450) );
  NAND U11124 ( .A(a[46]), .B(b[30]), .Z(n10449) );
  OR U11125 ( .A(n10450), .B(n10449), .Z(n10452) );
  XOR U11126 ( .A(n10448), .B(n10447), .Z(n10836) );
  XOR U11127 ( .A(n10450), .B(n10449), .Z(n10837) );
  NAND U11128 ( .A(n10836), .B(n10837), .Z(n10451) );
  NAND U11129 ( .A(n10452), .B(n10451), .Z(n10455) );
  AND U11130 ( .A(b[30]), .B(a[47]), .Z(n10456) );
  OR U11131 ( .A(n10455), .B(n10456), .Z(n10458) );
  XNOR U11132 ( .A(n10454), .B(n10453), .Z(n10843) );
  XOR U11133 ( .A(n10456), .B(n10455), .Z(n10842) );
  NANDN U11134 ( .A(n10843), .B(n10842), .Z(n10457) );
  NAND U11135 ( .A(n10458), .B(n10457), .Z(n10462) );
  NAND U11136 ( .A(a[48]), .B(b[30]), .Z(n10461) );
  OR U11137 ( .A(n10462), .B(n10461), .Z(n10464) );
  XOR U11138 ( .A(n10460), .B(n10459), .Z(n10848) );
  XOR U11139 ( .A(n10462), .B(n10461), .Z(n10849) );
  NAND U11140 ( .A(n10848), .B(n10849), .Z(n10463) );
  NAND U11141 ( .A(n10464), .B(n10463), .Z(n10467) );
  AND U11142 ( .A(b[30]), .B(a[49]), .Z(n10468) );
  OR U11143 ( .A(n10467), .B(n10468), .Z(n10470) );
  XNOR U11144 ( .A(n10466), .B(n10465), .Z(n10855) );
  XOR U11145 ( .A(n10468), .B(n10467), .Z(n10854) );
  NANDN U11146 ( .A(n10855), .B(n10854), .Z(n10469) );
  NAND U11147 ( .A(n10470), .B(n10469), .Z(n10474) );
  NAND U11148 ( .A(a[50]), .B(b[30]), .Z(n10473) );
  OR U11149 ( .A(n10474), .B(n10473), .Z(n10476) );
  XOR U11150 ( .A(n10472), .B(n10471), .Z(n10860) );
  XOR U11151 ( .A(n10474), .B(n10473), .Z(n10861) );
  NAND U11152 ( .A(n10860), .B(n10861), .Z(n10475) );
  NAND U11153 ( .A(n10476), .B(n10475), .Z(n10479) );
  AND U11154 ( .A(b[30]), .B(a[51]), .Z(n10480) );
  OR U11155 ( .A(n10479), .B(n10480), .Z(n10482) );
  XNOR U11156 ( .A(n10478), .B(n10477), .Z(n10867) );
  XOR U11157 ( .A(n10480), .B(n10479), .Z(n10866) );
  NANDN U11158 ( .A(n10867), .B(n10866), .Z(n10481) );
  NAND U11159 ( .A(n10482), .B(n10481), .Z(n10486) );
  NAND U11160 ( .A(a[52]), .B(b[30]), .Z(n10485) );
  OR U11161 ( .A(n10486), .B(n10485), .Z(n10488) );
  XOR U11162 ( .A(n10484), .B(n10483), .Z(n10872) );
  XOR U11163 ( .A(n10486), .B(n10485), .Z(n10873) );
  NAND U11164 ( .A(n10872), .B(n10873), .Z(n10487) );
  NAND U11165 ( .A(n10488), .B(n10487), .Z(n10491) );
  AND U11166 ( .A(b[30]), .B(a[53]), .Z(n10492) );
  OR U11167 ( .A(n10491), .B(n10492), .Z(n10494) );
  XNOR U11168 ( .A(n10490), .B(n10489), .Z(n10879) );
  XOR U11169 ( .A(n10492), .B(n10491), .Z(n10878) );
  NANDN U11170 ( .A(n10879), .B(n10878), .Z(n10493) );
  NAND U11171 ( .A(n10494), .B(n10493), .Z(n10498) );
  NAND U11172 ( .A(a[54]), .B(b[30]), .Z(n10497) );
  OR U11173 ( .A(n10498), .B(n10497), .Z(n10500) );
  XOR U11174 ( .A(n10496), .B(n10495), .Z(n10884) );
  XOR U11175 ( .A(n10498), .B(n10497), .Z(n10885) );
  NAND U11176 ( .A(n10884), .B(n10885), .Z(n10499) );
  NAND U11177 ( .A(n10500), .B(n10499), .Z(n10503) );
  AND U11178 ( .A(b[30]), .B(a[55]), .Z(n10504) );
  OR U11179 ( .A(n10503), .B(n10504), .Z(n10506) );
  XNOR U11180 ( .A(n10502), .B(n10501), .Z(n10891) );
  XOR U11181 ( .A(n10504), .B(n10503), .Z(n10890) );
  NANDN U11182 ( .A(n10891), .B(n10890), .Z(n10505) );
  NAND U11183 ( .A(n10506), .B(n10505), .Z(n10510) );
  NAND U11184 ( .A(a[56]), .B(b[30]), .Z(n10509) );
  OR U11185 ( .A(n10510), .B(n10509), .Z(n10512) );
  XOR U11186 ( .A(n10508), .B(n10507), .Z(n10896) );
  XOR U11187 ( .A(n10510), .B(n10509), .Z(n10897) );
  NAND U11188 ( .A(n10896), .B(n10897), .Z(n10511) );
  NAND U11189 ( .A(n10512), .B(n10511), .Z(n10515) );
  AND U11190 ( .A(b[30]), .B(a[57]), .Z(n10516) );
  OR U11191 ( .A(n10515), .B(n10516), .Z(n10518) );
  XNOR U11192 ( .A(n10514), .B(n10513), .Z(n10903) );
  XOR U11193 ( .A(n10516), .B(n10515), .Z(n10902) );
  NANDN U11194 ( .A(n10903), .B(n10902), .Z(n10517) );
  NAND U11195 ( .A(n10518), .B(n10517), .Z(n10522) );
  NAND U11196 ( .A(a[58]), .B(b[30]), .Z(n10521) );
  OR U11197 ( .A(n10522), .B(n10521), .Z(n10524) );
  XOR U11198 ( .A(n10520), .B(n10519), .Z(n10908) );
  XOR U11199 ( .A(n10522), .B(n10521), .Z(n10909) );
  NAND U11200 ( .A(n10908), .B(n10909), .Z(n10523) );
  NAND U11201 ( .A(n10524), .B(n10523), .Z(n10527) );
  AND U11202 ( .A(b[30]), .B(a[59]), .Z(n10528) );
  OR U11203 ( .A(n10527), .B(n10528), .Z(n10530) );
  XNOR U11204 ( .A(n10526), .B(n10525), .Z(n10915) );
  XOR U11205 ( .A(n10528), .B(n10527), .Z(n10914) );
  NANDN U11206 ( .A(n10915), .B(n10914), .Z(n10529) );
  NAND U11207 ( .A(n10530), .B(n10529), .Z(n10534) );
  NAND U11208 ( .A(a[60]), .B(b[30]), .Z(n10533) );
  OR U11209 ( .A(n10534), .B(n10533), .Z(n10536) );
  XOR U11210 ( .A(n10532), .B(n10531), .Z(n10921) );
  XOR U11211 ( .A(n10534), .B(n10533), .Z(n10920) );
  NAND U11212 ( .A(n10921), .B(n10920), .Z(n10535) );
  NAND U11213 ( .A(n10536), .B(n10535), .Z(n10539) );
  AND U11214 ( .A(b[30]), .B(a[61]), .Z(n10540) );
  OR U11215 ( .A(n10539), .B(n10540), .Z(n10542) );
  XNOR U11216 ( .A(n10538), .B(n10537), .Z(n10927) );
  XOR U11217 ( .A(n10540), .B(n10539), .Z(n10926) );
  NANDN U11218 ( .A(n10927), .B(n10926), .Z(n10541) );
  NAND U11219 ( .A(n10542), .B(n10541), .Z(n10546) );
  NAND U11220 ( .A(a[62]), .B(b[30]), .Z(n10545) );
  OR U11221 ( .A(n10546), .B(n10545), .Z(n10548) );
  XOR U11222 ( .A(n10544), .B(n10543), .Z(n10932) );
  XOR U11223 ( .A(n10546), .B(n10545), .Z(n10933) );
  NAND U11224 ( .A(n10932), .B(n10933), .Z(n10547) );
  NAND U11225 ( .A(n10548), .B(n10547), .Z(n10551) );
  AND U11226 ( .A(b[30]), .B(a[63]), .Z(n10552) );
  OR U11227 ( .A(n10551), .B(n10552), .Z(n10554) );
  XNOR U11228 ( .A(n10550), .B(n10549), .Z(n10562) );
  XOR U11229 ( .A(n10552), .B(n10551), .Z(n10561) );
  NANDN U11230 ( .A(n10562), .B(n10561), .Z(n10553) );
  AND U11231 ( .A(n10554), .B(n10553), .Z(n10559) );
  NAND U11232 ( .A(n10560), .B(n10559), .Z(n10558) );
  XOR U11233 ( .A(n10556), .B(n10555), .Z(n10557) );
  NANDN U11234 ( .A(n10558), .B(n10557), .Z(n21987) );
  XOR U11235 ( .A(n10558), .B(n10557), .Z(n24198) );
  XOR U11236 ( .A(n10560), .B(n10559), .Z(n21982) );
  XNOR U11237 ( .A(n10562), .B(n10561), .Z(n21979) );
  NAND U11238 ( .A(a[62]), .B(b[29]), .Z(n10928) );
  NAND U11239 ( .A(a[60]), .B(b[29]), .Z(n10916) );
  NAND U11240 ( .A(a[58]), .B(b[29]), .Z(n10904) );
  NAND U11241 ( .A(a[56]), .B(b[29]), .Z(n10892) );
  NAND U11242 ( .A(a[54]), .B(b[29]), .Z(n10880) );
  NAND U11243 ( .A(a[52]), .B(b[29]), .Z(n10868) );
  NAND U11244 ( .A(a[50]), .B(b[29]), .Z(n10856) );
  NAND U11245 ( .A(a[48]), .B(b[29]), .Z(n10844) );
  NAND U11246 ( .A(a[46]), .B(b[29]), .Z(n10832) );
  NAND U11247 ( .A(a[44]), .B(b[29]), .Z(n10820) );
  NAND U11248 ( .A(a[42]), .B(b[29]), .Z(n10808) );
  NAND U11249 ( .A(a[40]), .B(b[29]), .Z(n10796) );
  NAND U11250 ( .A(a[38]), .B(b[29]), .Z(n10784) );
  ANDN U11251 ( .B(b[29]), .A(n21727), .Z(n10728) );
  ANDN U11252 ( .B(b[29]), .A(n166), .Z(n10596) );
  ANDN U11253 ( .B(b[29]), .A(n164), .Z(n10587) );
  ANDN U11254 ( .B(b[29]), .A(n21580), .Z(n10572) );
  NAND U11255 ( .A(b[30]), .B(a[1]), .Z(n10565) );
  AND U11256 ( .A(b[29]), .B(a[0]), .Z(n11323) );
  NANDN U11257 ( .A(n10565), .B(n11323), .Z(n10564) );
  NAND U11258 ( .A(a[2]), .B(b[29]), .Z(n10563) );
  AND U11259 ( .A(n10564), .B(n10563), .Z(n10571) );
  NANDN U11260 ( .A(n10565), .B(a[0]), .Z(n10566) );
  XNOR U11261 ( .A(a[2]), .B(n10566), .Z(n10567) );
  NAND U11262 ( .A(b[29]), .B(n10567), .Z(n10954) );
  AND U11263 ( .A(a[1]), .B(b[30]), .Z(n10568) );
  XNOR U11264 ( .A(n10569), .B(n10568), .Z(n10953) );
  NANDN U11265 ( .A(n10954), .B(n10953), .Z(n10570) );
  NANDN U11266 ( .A(n10571), .B(n10570), .Z(n10573) );
  NANDN U11267 ( .A(n10572), .B(n10573), .Z(n10577) );
  XOR U11268 ( .A(n10573), .B(n10572), .Z(n10958) );
  NANDN U11269 ( .A(n10958), .B(n10957), .Z(n10576) );
  NAND U11270 ( .A(n10577), .B(n10576), .Z(n10581) );
  XOR U11271 ( .A(n10579), .B(n10578), .Z(n10580) );
  NANDN U11272 ( .A(n10581), .B(n10580), .Z(n10583) );
  NAND U11273 ( .A(a[4]), .B(b[29]), .Z(n10963) );
  NANDN U11274 ( .A(n10963), .B(n10964), .Z(n10582) );
  NAND U11275 ( .A(n10583), .B(n10582), .Z(n10586) );
  OR U11276 ( .A(n10587), .B(n10586), .Z(n10589) );
  XOR U11277 ( .A(n10585), .B(n10584), .Z(n10941) );
  XOR U11278 ( .A(n10587), .B(n10586), .Z(n10940) );
  NAND U11279 ( .A(n10941), .B(n10940), .Z(n10588) );
  NAND U11280 ( .A(n10589), .B(n10588), .Z(n10593) );
  XOR U11281 ( .A(n10591), .B(n10590), .Z(n10592) );
  NAND U11282 ( .A(n10593), .B(n10592), .Z(n10595) );
  ANDN U11283 ( .B(b[29]), .A(n165), .Z(n10976) );
  XNOR U11284 ( .A(n10593), .B(n10592), .Z(n10975) );
  OR U11285 ( .A(n10976), .B(n10975), .Z(n10594) );
  AND U11286 ( .A(n10595), .B(n10594), .Z(n10597) );
  OR U11287 ( .A(n10596), .B(n10597), .Z(n10601) );
  XNOR U11288 ( .A(n10597), .B(n10596), .Z(n10980) );
  XNOR U11289 ( .A(n10599), .B(n10598), .Z(n10979) );
  OR U11290 ( .A(n10980), .B(n10979), .Z(n10600) );
  NAND U11291 ( .A(n10601), .B(n10600), .Z(n10604) );
  XOR U11292 ( .A(n10603), .B(n10602), .Z(n10605) );
  OR U11293 ( .A(n10604), .B(n10605), .Z(n10607) );
  NAND U11294 ( .A(a[8]), .B(b[29]), .Z(n10988) );
  XOR U11295 ( .A(n10605), .B(n10604), .Z(n10987) );
  NANDN U11296 ( .A(n10988), .B(n10987), .Z(n10606) );
  NAND U11297 ( .A(n10607), .B(n10606), .Z(n10608) );
  ANDN U11298 ( .B(b[29]), .A(n21615), .Z(n10609) );
  OR U11299 ( .A(n10608), .B(n10609), .Z(n10613) );
  XNOR U11300 ( .A(n10609), .B(n10608), .Z(n10991) );
  OR U11301 ( .A(n10991), .B(n10992), .Z(n10612) );
  NAND U11302 ( .A(n10613), .B(n10612), .Z(n10616) );
  XNOR U11303 ( .A(n10615), .B(n10614), .Z(n10617) );
  OR U11304 ( .A(n10616), .B(n10617), .Z(n10619) );
  XNOR U11305 ( .A(n10617), .B(n10616), .Z(n11000) );
  AND U11306 ( .A(b[29]), .B(a[10]), .Z(n10999) );
  NANDN U11307 ( .A(n11000), .B(n10999), .Z(n10618) );
  NAND U11308 ( .A(n10619), .B(n10618), .Z(n10622) );
  ANDN U11309 ( .B(b[29]), .A(n21164), .Z(n10623) );
  OR U11310 ( .A(n10622), .B(n10623), .Z(n10625) );
  XOR U11311 ( .A(n10621), .B(n10620), .Z(n11004) );
  XOR U11312 ( .A(n10623), .B(n10622), .Z(n11003) );
  NANDN U11313 ( .A(n11004), .B(n11003), .Z(n10624) );
  NAND U11314 ( .A(n10625), .B(n10624), .Z(n10628) );
  XNOR U11315 ( .A(n10627), .B(n10626), .Z(n10629) );
  OR U11316 ( .A(n10628), .B(n10629), .Z(n10631) );
  XNOR U11317 ( .A(n10629), .B(n10628), .Z(n11010) );
  NAND U11318 ( .A(a[12]), .B(b[29]), .Z(n11009) );
  OR U11319 ( .A(n11010), .B(n11009), .Z(n10630) );
  NAND U11320 ( .A(n10631), .B(n10630), .Z(n10634) );
  ANDN U11321 ( .B(b[29]), .A(n170), .Z(n10635) );
  OR U11322 ( .A(n10634), .B(n10635), .Z(n10637) );
  XOR U11323 ( .A(n10633), .B(n10632), .Z(n11016) );
  XOR U11324 ( .A(n10635), .B(n10634), .Z(n11015) );
  NANDN U11325 ( .A(n11016), .B(n11015), .Z(n10636) );
  NAND U11326 ( .A(n10637), .B(n10636), .Z(n10640) );
  XNOR U11327 ( .A(n10639), .B(n10638), .Z(n10641) );
  OR U11328 ( .A(n10640), .B(n10641), .Z(n10643) );
  XNOR U11329 ( .A(n10641), .B(n10640), .Z(n11022) );
  NAND U11330 ( .A(a[14]), .B(b[29]), .Z(n11021) );
  OR U11331 ( .A(n11022), .B(n11021), .Z(n10642) );
  NAND U11332 ( .A(n10643), .B(n10642), .Z(n10646) );
  ANDN U11333 ( .B(b[29]), .A(n172), .Z(n10647) );
  OR U11334 ( .A(n10646), .B(n10647), .Z(n10649) );
  XOR U11335 ( .A(n10645), .B(n10644), .Z(n11028) );
  XOR U11336 ( .A(n10647), .B(n10646), .Z(n11027) );
  NANDN U11337 ( .A(n11028), .B(n11027), .Z(n10648) );
  NAND U11338 ( .A(n10649), .B(n10648), .Z(n10652) );
  XNOR U11339 ( .A(n10651), .B(n10650), .Z(n10653) );
  OR U11340 ( .A(n10652), .B(n10653), .Z(n10655) );
  XNOR U11341 ( .A(n10653), .B(n10652), .Z(n11034) );
  NAND U11342 ( .A(a[16]), .B(b[29]), .Z(n11033) );
  OR U11343 ( .A(n11034), .B(n11033), .Z(n10654) );
  NAND U11344 ( .A(n10655), .B(n10654), .Z(n10658) );
  ANDN U11345 ( .B(b[29]), .A(n174), .Z(n10659) );
  OR U11346 ( .A(n10658), .B(n10659), .Z(n10661) );
  XOR U11347 ( .A(n10659), .B(n10658), .Z(n11039) );
  NANDN U11348 ( .A(n11040), .B(n11039), .Z(n10660) );
  NAND U11349 ( .A(n10661), .B(n10660), .Z(n10664) );
  XNOR U11350 ( .A(n10663), .B(n10662), .Z(n10665) );
  OR U11351 ( .A(n10664), .B(n10665), .Z(n10667) );
  XNOR U11352 ( .A(n10665), .B(n10664), .Z(n11046) );
  NAND U11353 ( .A(a[18]), .B(b[29]), .Z(n11045) );
  OR U11354 ( .A(n11046), .B(n11045), .Z(n10666) );
  NAND U11355 ( .A(n10667), .B(n10666), .Z(n10670) );
  ANDN U11356 ( .B(b[29]), .A(n21670), .Z(n10671) );
  OR U11357 ( .A(n10670), .B(n10671), .Z(n10673) );
  XOR U11358 ( .A(n10669), .B(n10668), .Z(n11052) );
  XOR U11359 ( .A(n10671), .B(n10670), .Z(n11051) );
  NANDN U11360 ( .A(n11052), .B(n11051), .Z(n10672) );
  NAND U11361 ( .A(n10673), .B(n10672), .Z(n10676) );
  XNOR U11362 ( .A(n10675), .B(n10674), .Z(n10677) );
  OR U11363 ( .A(n10676), .B(n10677), .Z(n10679) );
  XNOR U11364 ( .A(n10677), .B(n10676), .Z(n11058) );
  NAND U11365 ( .A(a[20]), .B(b[29]), .Z(n11057) );
  OR U11366 ( .A(n11058), .B(n11057), .Z(n10678) );
  NAND U11367 ( .A(n10679), .B(n10678), .Z(n10682) );
  ANDN U11368 ( .B(b[29]), .A(n21681), .Z(n10683) );
  OR U11369 ( .A(n10682), .B(n10683), .Z(n10685) );
  XOR U11370 ( .A(n10681), .B(n10680), .Z(n11064) );
  XOR U11371 ( .A(n10683), .B(n10682), .Z(n11063) );
  NANDN U11372 ( .A(n11064), .B(n11063), .Z(n10684) );
  NAND U11373 ( .A(n10685), .B(n10684), .Z(n10688) );
  XNOR U11374 ( .A(n10687), .B(n10686), .Z(n10689) );
  OR U11375 ( .A(n10688), .B(n10689), .Z(n10691) );
  XNOR U11376 ( .A(n10689), .B(n10688), .Z(n11070) );
  NAND U11377 ( .A(a[22]), .B(b[29]), .Z(n11069) );
  OR U11378 ( .A(n11070), .B(n11069), .Z(n10690) );
  NAND U11379 ( .A(n10691), .B(n10690), .Z(n10694) );
  ANDN U11380 ( .B(b[29]), .A(n21692), .Z(n10695) );
  OR U11381 ( .A(n10694), .B(n10695), .Z(n10697) );
  XOR U11382 ( .A(n10693), .B(n10692), .Z(n11076) );
  XOR U11383 ( .A(n10695), .B(n10694), .Z(n11075) );
  NANDN U11384 ( .A(n11076), .B(n11075), .Z(n10696) );
  NAND U11385 ( .A(n10697), .B(n10696), .Z(n10700) );
  XNOR U11386 ( .A(n10699), .B(n10698), .Z(n10701) );
  OR U11387 ( .A(n10700), .B(n10701), .Z(n10703) );
  XNOR U11388 ( .A(n10701), .B(n10700), .Z(n11082) );
  NAND U11389 ( .A(a[24]), .B(b[29]), .Z(n11081) );
  OR U11390 ( .A(n11082), .B(n11081), .Z(n10702) );
  NAND U11391 ( .A(n10703), .B(n10702), .Z(n10706) );
  ANDN U11392 ( .B(b[29]), .A(n21703), .Z(n10707) );
  OR U11393 ( .A(n10706), .B(n10707), .Z(n10709) );
  XOR U11394 ( .A(n10707), .B(n10706), .Z(n11087) );
  NANDN U11395 ( .A(n11088), .B(n11087), .Z(n10708) );
  NAND U11396 ( .A(n10709), .B(n10708), .Z(n10712) );
  XOR U11397 ( .A(n10711), .B(n10710), .Z(n10713) );
  OR U11398 ( .A(n10712), .B(n10713), .Z(n10715) );
  NAND U11399 ( .A(a[26]), .B(b[29]), .Z(n11094) );
  XOR U11400 ( .A(n10713), .B(n10712), .Z(n11093) );
  NANDN U11401 ( .A(n11094), .B(n11093), .Z(n10714) );
  NAND U11402 ( .A(n10715), .B(n10714), .Z(n10716) );
  ANDN U11403 ( .B(b[29]), .A(n21716), .Z(n10717) );
  OR U11404 ( .A(n10716), .B(n10717), .Z(n10721) );
  XNOR U11405 ( .A(n10717), .B(n10716), .Z(n11100) );
  XNOR U11406 ( .A(n10719), .B(n10718), .Z(n11099) );
  OR U11407 ( .A(n11100), .B(n11099), .Z(n10720) );
  AND U11408 ( .A(n10721), .B(n10720), .Z(n10724) );
  XOR U11409 ( .A(n10723), .B(n10722), .Z(n10725) );
  OR U11410 ( .A(n10724), .B(n10725), .Z(n10727) );
  ANDN U11411 ( .B(b[29]), .A(n180), .Z(n11108) );
  XOR U11412 ( .A(n10725), .B(n10724), .Z(n11107) );
  NANDN U11413 ( .A(n11108), .B(n11107), .Z(n10726) );
  AND U11414 ( .A(n10727), .B(n10726), .Z(n10729) );
  OR U11415 ( .A(n10728), .B(n10729), .Z(n10733) );
  XNOR U11416 ( .A(n10729), .B(n10728), .Z(n11112) );
  XNOR U11417 ( .A(n10731), .B(n10730), .Z(n11111) );
  OR U11418 ( .A(n11112), .B(n11111), .Z(n10732) );
  NAND U11419 ( .A(n10733), .B(n10732), .Z(n10736) );
  XNOR U11420 ( .A(n10735), .B(n10734), .Z(n10737) );
  OR U11421 ( .A(n10736), .B(n10737), .Z(n10739) );
  XNOR U11422 ( .A(n10737), .B(n10736), .Z(n11120) );
  NAND U11423 ( .A(a[30]), .B(b[29]), .Z(n11119) );
  OR U11424 ( .A(n11120), .B(n11119), .Z(n10738) );
  NAND U11425 ( .A(n10739), .B(n10738), .Z(n10742) );
  ANDN U11426 ( .B(b[29]), .A(n21740), .Z(n10743) );
  OR U11427 ( .A(n10742), .B(n10743), .Z(n10745) );
  XOR U11428 ( .A(n10741), .B(n10740), .Z(n11124) );
  XOR U11429 ( .A(n10743), .B(n10742), .Z(n11123) );
  NANDN U11430 ( .A(n11124), .B(n11123), .Z(n10744) );
  NAND U11431 ( .A(n10745), .B(n10744), .Z(n10748) );
  XNOR U11432 ( .A(n10747), .B(n10746), .Z(n10749) );
  OR U11433 ( .A(n10748), .B(n10749), .Z(n10751) );
  XNOR U11434 ( .A(n10749), .B(n10748), .Z(n11130) );
  NAND U11435 ( .A(a[32]), .B(b[29]), .Z(n11129) );
  OR U11436 ( .A(n11130), .B(n11129), .Z(n10750) );
  NAND U11437 ( .A(n10751), .B(n10750), .Z(n10754) );
  ANDN U11438 ( .B(b[29]), .A(n21751), .Z(n10755) );
  OR U11439 ( .A(n10754), .B(n10755), .Z(n10757) );
  XOR U11440 ( .A(n10753), .B(n10752), .Z(n11136) );
  XOR U11441 ( .A(n10755), .B(n10754), .Z(n11135) );
  NANDN U11442 ( .A(n11136), .B(n11135), .Z(n10756) );
  NAND U11443 ( .A(n10757), .B(n10756), .Z(n10760) );
  XNOR U11444 ( .A(n10759), .B(n10758), .Z(n10761) );
  OR U11445 ( .A(n10760), .B(n10761), .Z(n10763) );
  XNOR U11446 ( .A(n10761), .B(n10760), .Z(n11142) );
  NAND U11447 ( .A(a[34]), .B(b[29]), .Z(n11141) );
  OR U11448 ( .A(n11142), .B(n11141), .Z(n10762) );
  NAND U11449 ( .A(n10763), .B(n10762), .Z(n10764) );
  ANDN U11450 ( .B(b[29]), .A(n184), .Z(n10765) );
  OR U11451 ( .A(n10764), .B(n10765), .Z(n10769) );
  XOR U11452 ( .A(n10765), .B(n10764), .Z(n11147) );
  NAND U11453 ( .A(n11147), .B(n11148), .Z(n10768) );
  NAND U11454 ( .A(n10769), .B(n10768), .Z(n10773) );
  NAND U11455 ( .A(a[36]), .B(b[29]), .Z(n10772) );
  OR U11456 ( .A(n10773), .B(n10772), .Z(n10775) );
  XOR U11457 ( .A(n10771), .B(n10770), .Z(n11153) );
  XOR U11458 ( .A(n10773), .B(n10772), .Z(n11154) );
  NAND U11459 ( .A(n11153), .B(n11154), .Z(n10774) );
  NAND U11460 ( .A(n10775), .B(n10774), .Z(n10779) );
  XOR U11461 ( .A(n10777), .B(n10776), .Z(n10778) );
  NAND U11462 ( .A(n10779), .B(n10778), .Z(n10781) );
  XNOR U11463 ( .A(n10779), .B(n10778), .Z(n11160) );
  NAND U11464 ( .A(a[37]), .B(b[29]), .Z(n11159) );
  OR U11465 ( .A(n11160), .B(n11159), .Z(n10780) );
  NAND U11466 ( .A(n10781), .B(n10780), .Z(n10785) );
  NANDN U11467 ( .A(n10784), .B(n10785), .Z(n10787) );
  XNOR U11468 ( .A(n10783), .B(n10782), .Z(n11166) );
  XNOR U11469 ( .A(n10785), .B(n10784), .Z(n11165) );
  NANDN U11470 ( .A(n11166), .B(n11165), .Z(n10786) );
  NAND U11471 ( .A(n10787), .B(n10786), .Z(n10791) );
  XOR U11472 ( .A(n10789), .B(n10788), .Z(n10790) );
  NAND U11473 ( .A(n10791), .B(n10790), .Z(n10793) );
  XNOR U11474 ( .A(n10791), .B(n10790), .Z(n11172) );
  NAND U11475 ( .A(a[39]), .B(b[29]), .Z(n11171) );
  OR U11476 ( .A(n11172), .B(n11171), .Z(n10792) );
  NAND U11477 ( .A(n10793), .B(n10792), .Z(n10797) );
  NANDN U11478 ( .A(n10796), .B(n10797), .Z(n10799) );
  XNOR U11479 ( .A(n10795), .B(n10794), .Z(n11178) );
  XNOR U11480 ( .A(n10797), .B(n10796), .Z(n11177) );
  NANDN U11481 ( .A(n11178), .B(n11177), .Z(n10798) );
  NAND U11482 ( .A(n10799), .B(n10798), .Z(n10803) );
  XOR U11483 ( .A(n10801), .B(n10800), .Z(n10802) );
  NAND U11484 ( .A(n10803), .B(n10802), .Z(n10805) );
  XNOR U11485 ( .A(n10803), .B(n10802), .Z(n11184) );
  NAND U11486 ( .A(a[41]), .B(b[29]), .Z(n11183) );
  OR U11487 ( .A(n11184), .B(n11183), .Z(n10804) );
  NAND U11488 ( .A(n10805), .B(n10804), .Z(n10809) );
  NANDN U11489 ( .A(n10808), .B(n10809), .Z(n10811) );
  XNOR U11490 ( .A(n10807), .B(n10806), .Z(n11190) );
  XNOR U11491 ( .A(n10809), .B(n10808), .Z(n11189) );
  NANDN U11492 ( .A(n11190), .B(n11189), .Z(n10810) );
  NAND U11493 ( .A(n10811), .B(n10810), .Z(n10815) );
  XOR U11494 ( .A(n10813), .B(n10812), .Z(n10814) );
  NAND U11495 ( .A(n10815), .B(n10814), .Z(n10817) );
  XNOR U11496 ( .A(n10815), .B(n10814), .Z(n11196) );
  NAND U11497 ( .A(a[43]), .B(b[29]), .Z(n11195) );
  OR U11498 ( .A(n11196), .B(n11195), .Z(n10816) );
  NAND U11499 ( .A(n10817), .B(n10816), .Z(n10821) );
  NANDN U11500 ( .A(n10820), .B(n10821), .Z(n10823) );
  XNOR U11501 ( .A(n10819), .B(n10818), .Z(n11202) );
  XNOR U11502 ( .A(n10821), .B(n10820), .Z(n11201) );
  NANDN U11503 ( .A(n11202), .B(n11201), .Z(n10822) );
  NAND U11504 ( .A(n10823), .B(n10822), .Z(n10827) );
  XOR U11505 ( .A(n10825), .B(n10824), .Z(n10826) );
  NAND U11506 ( .A(n10827), .B(n10826), .Z(n10829) );
  XNOR U11507 ( .A(n10827), .B(n10826), .Z(n11208) );
  NAND U11508 ( .A(a[45]), .B(b[29]), .Z(n11207) );
  OR U11509 ( .A(n11208), .B(n11207), .Z(n10828) );
  NAND U11510 ( .A(n10829), .B(n10828), .Z(n10833) );
  NANDN U11511 ( .A(n10832), .B(n10833), .Z(n10835) );
  XNOR U11512 ( .A(n10831), .B(n10830), .Z(n11214) );
  XNOR U11513 ( .A(n10833), .B(n10832), .Z(n11213) );
  NANDN U11514 ( .A(n11214), .B(n11213), .Z(n10834) );
  NAND U11515 ( .A(n10835), .B(n10834), .Z(n10839) );
  XOR U11516 ( .A(n10837), .B(n10836), .Z(n10838) );
  NAND U11517 ( .A(n10839), .B(n10838), .Z(n10841) );
  XNOR U11518 ( .A(n10839), .B(n10838), .Z(n11220) );
  NAND U11519 ( .A(a[47]), .B(b[29]), .Z(n11219) );
  OR U11520 ( .A(n11220), .B(n11219), .Z(n10840) );
  NAND U11521 ( .A(n10841), .B(n10840), .Z(n10845) );
  NANDN U11522 ( .A(n10844), .B(n10845), .Z(n10847) );
  XNOR U11523 ( .A(n10843), .B(n10842), .Z(n11226) );
  XNOR U11524 ( .A(n10845), .B(n10844), .Z(n11225) );
  NANDN U11525 ( .A(n11226), .B(n11225), .Z(n10846) );
  NAND U11526 ( .A(n10847), .B(n10846), .Z(n10851) );
  XOR U11527 ( .A(n10849), .B(n10848), .Z(n10850) );
  NAND U11528 ( .A(n10851), .B(n10850), .Z(n10853) );
  XNOR U11529 ( .A(n10851), .B(n10850), .Z(n11232) );
  NAND U11530 ( .A(a[49]), .B(b[29]), .Z(n11231) );
  OR U11531 ( .A(n11232), .B(n11231), .Z(n10852) );
  NAND U11532 ( .A(n10853), .B(n10852), .Z(n10857) );
  NANDN U11533 ( .A(n10856), .B(n10857), .Z(n10859) );
  XNOR U11534 ( .A(n10855), .B(n10854), .Z(n11238) );
  XNOR U11535 ( .A(n10857), .B(n10856), .Z(n11237) );
  NANDN U11536 ( .A(n11238), .B(n11237), .Z(n10858) );
  NAND U11537 ( .A(n10859), .B(n10858), .Z(n10863) );
  XOR U11538 ( .A(n10861), .B(n10860), .Z(n10862) );
  NAND U11539 ( .A(n10863), .B(n10862), .Z(n10865) );
  XNOR U11540 ( .A(n10863), .B(n10862), .Z(n11244) );
  NAND U11541 ( .A(a[51]), .B(b[29]), .Z(n11243) );
  OR U11542 ( .A(n11244), .B(n11243), .Z(n10864) );
  NAND U11543 ( .A(n10865), .B(n10864), .Z(n10869) );
  NANDN U11544 ( .A(n10868), .B(n10869), .Z(n10871) );
  XNOR U11545 ( .A(n10867), .B(n10866), .Z(n11250) );
  XNOR U11546 ( .A(n10869), .B(n10868), .Z(n11249) );
  NANDN U11547 ( .A(n11250), .B(n11249), .Z(n10870) );
  NAND U11548 ( .A(n10871), .B(n10870), .Z(n10875) );
  XOR U11549 ( .A(n10873), .B(n10872), .Z(n10874) );
  NAND U11550 ( .A(n10875), .B(n10874), .Z(n10877) );
  XNOR U11551 ( .A(n10875), .B(n10874), .Z(n11256) );
  NAND U11552 ( .A(a[53]), .B(b[29]), .Z(n11255) );
  OR U11553 ( .A(n11256), .B(n11255), .Z(n10876) );
  NAND U11554 ( .A(n10877), .B(n10876), .Z(n10881) );
  NANDN U11555 ( .A(n10880), .B(n10881), .Z(n10883) );
  XNOR U11556 ( .A(n10879), .B(n10878), .Z(n11262) );
  XNOR U11557 ( .A(n10881), .B(n10880), .Z(n11261) );
  NANDN U11558 ( .A(n11262), .B(n11261), .Z(n10882) );
  NAND U11559 ( .A(n10883), .B(n10882), .Z(n10887) );
  XOR U11560 ( .A(n10885), .B(n10884), .Z(n10886) );
  NAND U11561 ( .A(n10887), .B(n10886), .Z(n10889) );
  XNOR U11562 ( .A(n10887), .B(n10886), .Z(n11268) );
  NAND U11563 ( .A(a[55]), .B(b[29]), .Z(n11267) );
  OR U11564 ( .A(n11268), .B(n11267), .Z(n10888) );
  NAND U11565 ( .A(n10889), .B(n10888), .Z(n10893) );
  NANDN U11566 ( .A(n10892), .B(n10893), .Z(n10895) );
  XNOR U11567 ( .A(n10891), .B(n10890), .Z(n11274) );
  XNOR U11568 ( .A(n10893), .B(n10892), .Z(n11273) );
  NANDN U11569 ( .A(n11274), .B(n11273), .Z(n10894) );
  NAND U11570 ( .A(n10895), .B(n10894), .Z(n10899) );
  XOR U11571 ( .A(n10897), .B(n10896), .Z(n10898) );
  NAND U11572 ( .A(n10899), .B(n10898), .Z(n10901) );
  XNOR U11573 ( .A(n10899), .B(n10898), .Z(n11280) );
  NAND U11574 ( .A(a[57]), .B(b[29]), .Z(n11279) );
  OR U11575 ( .A(n11280), .B(n11279), .Z(n10900) );
  NAND U11576 ( .A(n10901), .B(n10900), .Z(n10905) );
  NANDN U11577 ( .A(n10904), .B(n10905), .Z(n10907) );
  XNOR U11578 ( .A(n10903), .B(n10902), .Z(n11286) );
  XNOR U11579 ( .A(n10905), .B(n10904), .Z(n11285) );
  NANDN U11580 ( .A(n11286), .B(n11285), .Z(n10906) );
  NAND U11581 ( .A(n10907), .B(n10906), .Z(n10911) );
  XOR U11582 ( .A(n10909), .B(n10908), .Z(n10910) );
  NAND U11583 ( .A(n10911), .B(n10910), .Z(n10913) );
  XNOR U11584 ( .A(n10911), .B(n10910), .Z(n11292) );
  NAND U11585 ( .A(a[59]), .B(b[29]), .Z(n11291) );
  OR U11586 ( .A(n11292), .B(n11291), .Z(n10912) );
  NAND U11587 ( .A(n10913), .B(n10912), .Z(n10917) );
  NANDN U11588 ( .A(n10916), .B(n10917), .Z(n10919) );
  XNOR U11589 ( .A(n10915), .B(n10914), .Z(n11298) );
  XNOR U11590 ( .A(n10917), .B(n10916), .Z(n11297) );
  NANDN U11591 ( .A(n11298), .B(n11297), .Z(n10918) );
  NAND U11592 ( .A(n10919), .B(n10918), .Z(n10923) );
  XOR U11593 ( .A(n10921), .B(n10920), .Z(n10922) );
  NAND U11594 ( .A(n10923), .B(n10922), .Z(n10925) );
  XNOR U11595 ( .A(n10923), .B(n10922), .Z(n11304) );
  NAND U11596 ( .A(a[61]), .B(b[29]), .Z(n11303) );
  OR U11597 ( .A(n11304), .B(n11303), .Z(n10924) );
  NAND U11598 ( .A(n10925), .B(n10924), .Z(n10929) );
  NANDN U11599 ( .A(n10928), .B(n10929), .Z(n10931) );
  XNOR U11600 ( .A(n10927), .B(n10926), .Z(n10939) );
  XNOR U11601 ( .A(n10929), .B(n10928), .Z(n10938) );
  NANDN U11602 ( .A(n10939), .B(n10938), .Z(n10930) );
  NAND U11603 ( .A(n10931), .B(n10930), .Z(n10935) );
  XOR U11604 ( .A(n10933), .B(n10932), .Z(n10934) );
  NAND U11605 ( .A(n10935), .B(n10934), .Z(n10937) );
  XNOR U11606 ( .A(n10935), .B(n10934), .Z(n12064) );
  NAND U11607 ( .A(a[63]), .B(b[29]), .Z(n12063) );
  OR U11608 ( .A(n12064), .B(n12063), .Z(n10936) );
  AND U11609 ( .A(n10937), .B(n10936), .Z(n21978) );
  OR U11610 ( .A(n21979), .B(n21978), .Z(n21983) );
  NANDN U11611 ( .A(n21982), .B(n21983), .Z(n21985) );
  XNOR U11612 ( .A(n10939), .B(n10938), .Z(n12068) );
  AND U11613 ( .A(b[28]), .B(a[63]), .Z(n12065) );
  NAND U11614 ( .A(a[38]), .B(b[28]), .Z(n11161) );
  NAND U11615 ( .A(a[11]), .B(b[28]), .Z(n10998) );
  ANDN U11616 ( .B(b[28]), .A(n166), .Z(n10973) );
  XNOR U11617 ( .A(n10941), .B(n10940), .Z(n10970) );
  ANDN U11618 ( .B(b[28]), .A(n164), .Z(n10966) );
  ANDN U11619 ( .B(b[28]), .A(n21580), .Z(n10951) );
  NAND U11620 ( .A(b[29]), .B(a[1]), .Z(n10944) );
  AND U11621 ( .A(b[28]), .B(a[0]), .Z(n11694) );
  NANDN U11622 ( .A(n10944), .B(n11694), .Z(n10943) );
  NAND U11623 ( .A(a[2]), .B(b[28]), .Z(n10942) );
  AND U11624 ( .A(n10943), .B(n10942), .Z(n10950) );
  NANDN U11625 ( .A(n10944), .B(a[0]), .Z(n10945) );
  XNOR U11626 ( .A(a[2]), .B(n10945), .Z(n10946) );
  NAND U11627 ( .A(b[28]), .B(n10946), .Z(n11329) );
  AND U11628 ( .A(a[1]), .B(b[29]), .Z(n10947) );
  XNOR U11629 ( .A(n10948), .B(n10947), .Z(n11328) );
  NANDN U11630 ( .A(n11329), .B(n11328), .Z(n10949) );
  NANDN U11631 ( .A(n10950), .B(n10949), .Z(n10952) );
  NANDN U11632 ( .A(n10951), .B(n10952), .Z(n10956) );
  XOR U11633 ( .A(n10952), .B(n10951), .Z(n11333) );
  NANDN U11634 ( .A(n11333), .B(n11332), .Z(n10955) );
  NAND U11635 ( .A(n10956), .B(n10955), .Z(n10960) );
  XOR U11636 ( .A(n10958), .B(n10957), .Z(n10959) );
  NANDN U11637 ( .A(n10960), .B(n10959), .Z(n10962) );
  NAND U11638 ( .A(a[4]), .B(b[28]), .Z(n11338) );
  NANDN U11639 ( .A(n11338), .B(n11339), .Z(n10961) );
  NAND U11640 ( .A(n10962), .B(n10961), .Z(n10965) );
  OR U11641 ( .A(n10966), .B(n10965), .Z(n10968) );
  XOR U11642 ( .A(n10964), .B(n10963), .Z(n11316) );
  XOR U11643 ( .A(n10966), .B(n10965), .Z(n11315) );
  NAND U11644 ( .A(n11316), .B(n11315), .Z(n10967) );
  NAND U11645 ( .A(n10968), .B(n10967), .Z(n10969) );
  NANDN U11646 ( .A(n10970), .B(n10969), .Z(n10972) );
  ANDN U11647 ( .B(b[28]), .A(n165), .Z(n11351) );
  NANDN U11648 ( .A(n11351), .B(n11350), .Z(n10971) );
  NAND U11649 ( .A(n10972), .B(n10971), .Z(n10974) );
  NANDN U11650 ( .A(n10973), .B(n10974), .Z(n10978) );
  XOR U11651 ( .A(n10974), .B(n10973), .Z(n11355) );
  XOR U11652 ( .A(n10976), .B(n10975), .Z(n11354) );
  NANDN U11653 ( .A(n11355), .B(n11354), .Z(n10977) );
  NAND U11654 ( .A(n10978), .B(n10977), .Z(n10981) );
  XOR U11655 ( .A(n10980), .B(n10979), .Z(n10982) );
  OR U11656 ( .A(n10981), .B(n10982), .Z(n10984) );
  NAND U11657 ( .A(a[8]), .B(b[28]), .Z(n11363) );
  XOR U11658 ( .A(n10982), .B(n10981), .Z(n11362) );
  NANDN U11659 ( .A(n11363), .B(n11362), .Z(n10983) );
  NAND U11660 ( .A(n10984), .B(n10983), .Z(n10985) );
  ANDN U11661 ( .B(b[28]), .A(n21615), .Z(n10986) );
  OR U11662 ( .A(n10985), .B(n10986), .Z(n10990) );
  XNOR U11663 ( .A(n10986), .B(n10985), .Z(n11366) );
  OR U11664 ( .A(n11366), .B(n11367), .Z(n10989) );
  AND U11665 ( .A(n10990), .B(n10989), .Z(n10994) );
  XOR U11666 ( .A(n10992), .B(n10991), .Z(n10993) );
  NANDN U11667 ( .A(n10994), .B(n10993), .Z(n10996) );
  XOR U11668 ( .A(n10994), .B(n10993), .Z(n11374) );
  ANDN U11669 ( .B(b[28]), .A(n168), .Z(n11375) );
  OR U11670 ( .A(n11374), .B(n11375), .Z(n10995) );
  NAND U11671 ( .A(n10996), .B(n10995), .Z(n10997) );
  OR U11672 ( .A(n10998), .B(n10997), .Z(n11002) );
  XNOR U11673 ( .A(n10998), .B(n10997), .Z(n11379) );
  XNOR U11674 ( .A(n11000), .B(n10999), .Z(n11378) );
  NANDN U11675 ( .A(n11379), .B(n11378), .Z(n11001) );
  AND U11676 ( .A(n11002), .B(n11001), .Z(n11005) );
  XNOR U11677 ( .A(n11004), .B(n11003), .Z(n11006) );
  OR U11678 ( .A(n11005), .B(n11006), .Z(n11008) );
  XNOR U11679 ( .A(n11006), .B(n11005), .Z(n11387) );
  AND U11680 ( .A(b[28]), .B(a[12]), .Z(n11386) );
  NANDN U11681 ( .A(n11387), .B(n11386), .Z(n11007) );
  NAND U11682 ( .A(n11008), .B(n11007), .Z(n11011) );
  ANDN U11683 ( .B(b[28]), .A(n170), .Z(n11012) );
  OR U11684 ( .A(n11011), .B(n11012), .Z(n11014) );
  XOR U11685 ( .A(n11010), .B(n11009), .Z(n11391) );
  XOR U11686 ( .A(n11012), .B(n11011), .Z(n11390) );
  NANDN U11687 ( .A(n11391), .B(n11390), .Z(n11013) );
  NAND U11688 ( .A(n11014), .B(n11013), .Z(n11017) );
  XNOR U11689 ( .A(n11016), .B(n11015), .Z(n11018) );
  OR U11690 ( .A(n11017), .B(n11018), .Z(n11020) );
  XNOR U11691 ( .A(n11018), .B(n11017), .Z(n11397) );
  NAND U11692 ( .A(a[14]), .B(b[28]), .Z(n11396) );
  OR U11693 ( .A(n11397), .B(n11396), .Z(n11019) );
  NAND U11694 ( .A(n11020), .B(n11019), .Z(n11023) );
  ANDN U11695 ( .B(b[28]), .A(n172), .Z(n11024) );
  OR U11696 ( .A(n11023), .B(n11024), .Z(n11026) );
  XOR U11697 ( .A(n11022), .B(n11021), .Z(n11403) );
  XOR U11698 ( .A(n11024), .B(n11023), .Z(n11402) );
  NANDN U11699 ( .A(n11403), .B(n11402), .Z(n11025) );
  NAND U11700 ( .A(n11026), .B(n11025), .Z(n11029) );
  XNOR U11701 ( .A(n11028), .B(n11027), .Z(n11030) );
  OR U11702 ( .A(n11029), .B(n11030), .Z(n11032) );
  XNOR U11703 ( .A(n11030), .B(n11029), .Z(n11409) );
  NAND U11704 ( .A(a[16]), .B(b[28]), .Z(n11408) );
  OR U11705 ( .A(n11409), .B(n11408), .Z(n11031) );
  NAND U11706 ( .A(n11032), .B(n11031), .Z(n11035) );
  ANDN U11707 ( .B(b[28]), .A(n174), .Z(n11036) );
  OR U11708 ( .A(n11035), .B(n11036), .Z(n11038) );
  XOR U11709 ( .A(n11034), .B(n11033), .Z(n11415) );
  XOR U11710 ( .A(n11036), .B(n11035), .Z(n11414) );
  NANDN U11711 ( .A(n11415), .B(n11414), .Z(n11037) );
  NAND U11712 ( .A(n11038), .B(n11037), .Z(n11041) );
  XNOR U11713 ( .A(n11040), .B(n11039), .Z(n11042) );
  OR U11714 ( .A(n11041), .B(n11042), .Z(n11044) );
  XNOR U11715 ( .A(n11042), .B(n11041), .Z(n11421) );
  NAND U11716 ( .A(a[18]), .B(b[28]), .Z(n11420) );
  OR U11717 ( .A(n11421), .B(n11420), .Z(n11043) );
  NAND U11718 ( .A(n11044), .B(n11043), .Z(n11047) );
  ANDN U11719 ( .B(b[28]), .A(n21670), .Z(n11048) );
  OR U11720 ( .A(n11047), .B(n11048), .Z(n11050) );
  XOR U11721 ( .A(n11046), .B(n11045), .Z(n11427) );
  XOR U11722 ( .A(n11048), .B(n11047), .Z(n11426) );
  NANDN U11723 ( .A(n11427), .B(n11426), .Z(n11049) );
  NAND U11724 ( .A(n11050), .B(n11049), .Z(n11053) );
  XNOR U11725 ( .A(n11052), .B(n11051), .Z(n11054) );
  OR U11726 ( .A(n11053), .B(n11054), .Z(n11056) );
  XNOR U11727 ( .A(n11054), .B(n11053), .Z(n11433) );
  NAND U11728 ( .A(a[20]), .B(b[28]), .Z(n11432) );
  OR U11729 ( .A(n11433), .B(n11432), .Z(n11055) );
  NAND U11730 ( .A(n11056), .B(n11055), .Z(n11059) );
  ANDN U11731 ( .B(b[28]), .A(n21681), .Z(n11060) );
  OR U11732 ( .A(n11059), .B(n11060), .Z(n11062) );
  XOR U11733 ( .A(n11058), .B(n11057), .Z(n11439) );
  XOR U11734 ( .A(n11060), .B(n11059), .Z(n11438) );
  NANDN U11735 ( .A(n11439), .B(n11438), .Z(n11061) );
  NAND U11736 ( .A(n11062), .B(n11061), .Z(n11065) );
  XNOR U11737 ( .A(n11064), .B(n11063), .Z(n11066) );
  OR U11738 ( .A(n11065), .B(n11066), .Z(n11068) );
  XNOR U11739 ( .A(n11066), .B(n11065), .Z(n11445) );
  NAND U11740 ( .A(a[22]), .B(b[28]), .Z(n11444) );
  OR U11741 ( .A(n11445), .B(n11444), .Z(n11067) );
  NAND U11742 ( .A(n11068), .B(n11067), .Z(n11071) );
  ANDN U11743 ( .B(b[28]), .A(n21692), .Z(n11072) );
  OR U11744 ( .A(n11071), .B(n11072), .Z(n11074) );
  XOR U11745 ( .A(n11070), .B(n11069), .Z(n11451) );
  XOR U11746 ( .A(n11072), .B(n11071), .Z(n11450) );
  NANDN U11747 ( .A(n11451), .B(n11450), .Z(n11073) );
  NAND U11748 ( .A(n11074), .B(n11073), .Z(n11077) );
  XNOR U11749 ( .A(n11076), .B(n11075), .Z(n11078) );
  OR U11750 ( .A(n11077), .B(n11078), .Z(n11080) );
  XNOR U11751 ( .A(n11078), .B(n11077), .Z(n11457) );
  NAND U11752 ( .A(a[24]), .B(b[28]), .Z(n11456) );
  OR U11753 ( .A(n11457), .B(n11456), .Z(n11079) );
  NAND U11754 ( .A(n11080), .B(n11079), .Z(n11083) );
  ANDN U11755 ( .B(b[28]), .A(n21703), .Z(n11084) );
  OR U11756 ( .A(n11083), .B(n11084), .Z(n11086) );
  XOR U11757 ( .A(n11082), .B(n11081), .Z(n11463) );
  XOR U11758 ( .A(n11084), .B(n11083), .Z(n11462) );
  NANDN U11759 ( .A(n11463), .B(n11462), .Z(n11085) );
  NAND U11760 ( .A(n11086), .B(n11085), .Z(n11089) );
  XNOR U11761 ( .A(n11088), .B(n11087), .Z(n11090) );
  OR U11762 ( .A(n11089), .B(n11090), .Z(n11092) );
  XNOR U11763 ( .A(n11090), .B(n11089), .Z(n11469) );
  NAND U11764 ( .A(a[26]), .B(b[28]), .Z(n11468) );
  OR U11765 ( .A(n11469), .B(n11468), .Z(n11091) );
  NAND U11766 ( .A(n11092), .B(n11091), .Z(n11095) );
  ANDN U11767 ( .B(b[28]), .A(n21716), .Z(n11096) );
  OR U11768 ( .A(n11095), .B(n11096), .Z(n11098) );
  XOR U11769 ( .A(n11096), .B(n11095), .Z(n11474) );
  NANDN U11770 ( .A(n11475), .B(n11474), .Z(n11097) );
  NAND U11771 ( .A(n11098), .B(n11097), .Z(n11101) );
  XOR U11772 ( .A(n11100), .B(n11099), .Z(n11102) );
  OR U11773 ( .A(n11101), .B(n11102), .Z(n11104) );
  NAND U11774 ( .A(a[28]), .B(b[28]), .Z(n11481) );
  XOR U11775 ( .A(n11102), .B(n11101), .Z(n11480) );
  NANDN U11776 ( .A(n11481), .B(n11480), .Z(n11103) );
  NAND U11777 ( .A(n11104), .B(n11103), .Z(n11105) );
  ANDN U11778 ( .B(b[28]), .A(n21727), .Z(n11106) );
  OR U11779 ( .A(n11105), .B(n11106), .Z(n11110) );
  XNOR U11780 ( .A(n11106), .B(n11105), .Z(n11487) );
  XOR U11781 ( .A(n11108), .B(n11107), .Z(n11486) );
  OR U11782 ( .A(n11487), .B(n11486), .Z(n11109) );
  NAND U11783 ( .A(n11110), .B(n11109), .Z(n11113) );
  XOR U11784 ( .A(n11112), .B(n11111), .Z(n11114) );
  OR U11785 ( .A(n11113), .B(n11114), .Z(n11116) );
  NAND U11786 ( .A(a[30]), .B(b[28]), .Z(n11493) );
  XOR U11787 ( .A(n11114), .B(n11113), .Z(n11492) );
  NANDN U11788 ( .A(n11493), .B(n11492), .Z(n11115) );
  NAND U11789 ( .A(n11116), .B(n11115), .Z(n11117) );
  ANDN U11790 ( .B(b[28]), .A(n21740), .Z(n11118) );
  OR U11791 ( .A(n11117), .B(n11118), .Z(n11122) );
  XNOR U11792 ( .A(n11118), .B(n11117), .Z(n11498) );
  XOR U11793 ( .A(n11120), .B(n11119), .Z(n11499) );
  OR U11794 ( .A(n11498), .B(n11499), .Z(n11121) );
  NAND U11795 ( .A(n11122), .B(n11121), .Z(n11125) );
  XNOR U11796 ( .A(n11124), .B(n11123), .Z(n11126) );
  OR U11797 ( .A(n11125), .B(n11126), .Z(n11128) );
  XNOR U11798 ( .A(n11126), .B(n11125), .Z(n11507) );
  AND U11799 ( .A(b[28]), .B(a[32]), .Z(n11506) );
  NANDN U11800 ( .A(n11507), .B(n11506), .Z(n11127) );
  NAND U11801 ( .A(n11128), .B(n11127), .Z(n11131) );
  ANDN U11802 ( .B(b[28]), .A(n21751), .Z(n11132) );
  OR U11803 ( .A(n11131), .B(n11132), .Z(n11134) );
  XOR U11804 ( .A(n11130), .B(n11129), .Z(n11511) );
  XOR U11805 ( .A(n11132), .B(n11131), .Z(n11510) );
  NANDN U11806 ( .A(n11511), .B(n11510), .Z(n11133) );
  NAND U11807 ( .A(n11134), .B(n11133), .Z(n11137) );
  XNOR U11808 ( .A(n11136), .B(n11135), .Z(n11138) );
  OR U11809 ( .A(n11137), .B(n11138), .Z(n11140) );
  XNOR U11810 ( .A(n11138), .B(n11137), .Z(n11517) );
  NAND U11811 ( .A(a[34]), .B(b[28]), .Z(n11516) );
  OR U11812 ( .A(n11517), .B(n11516), .Z(n11139) );
  NAND U11813 ( .A(n11140), .B(n11139), .Z(n11143) );
  ANDN U11814 ( .B(b[28]), .A(n184), .Z(n11144) );
  OR U11815 ( .A(n11143), .B(n11144), .Z(n11146) );
  XOR U11816 ( .A(n11142), .B(n11141), .Z(n11523) );
  XOR U11817 ( .A(n11144), .B(n11143), .Z(n11522) );
  NANDN U11818 ( .A(n11523), .B(n11522), .Z(n11145) );
  NAND U11819 ( .A(n11146), .B(n11145), .Z(n11150) );
  AND U11820 ( .A(b[28]), .B(a[36]), .Z(n11149) );
  NANDN U11821 ( .A(n11150), .B(n11149), .Z(n11152) );
  XNOR U11822 ( .A(n11150), .B(n11149), .Z(n11530) );
  NANDN U11823 ( .A(n11531), .B(n11530), .Z(n11151) );
  NAND U11824 ( .A(n11152), .B(n11151), .Z(n11156) );
  XOR U11825 ( .A(n11154), .B(n11153), .Z(n11155) );
  NAND U11826 ( .A(n11156), .B(n11155), .Z(n11158) );
  XNOR U11827 ( .A(n11156), .B(n11155), .Z(n11537) );
  NAND U11828 ( .A(a[37]), .B(b[28]), .Z(n11536) );
  OR U11829 ( .A(n11537), .B(n11536), .Z(n11157) );
  NAND U11830 ( .A(n11158), .B(n11157), .Z(n11162) );
  NANDN U11831 ( .A(n11161), .B(n11162), .Z(n11164) );
  XOR U11832 ( .A(n11160), .B(n11159), .Z(n11540) );
  XNOR U11833 ( .A(n11162), .B(n11161), .Z(n11541) );
  NAND U11834 ( .A(n11540), .B(n11541), .Z(n11163) );
  NAND U11835 ( .A(n11164), .B(n11163), .Z(n11167) );
  AND U11836 ( .A(b[28]), .B(a[39]), .Z(n11168) );
  OR U11837 ( .A(n11167), .B(n11168), .Z(n11170) );
  XNOR U11838 ( .A(n11166), .B(n11165), .Z(n11547) );
  XOR U11839 ( .A(n11168), .B(n11167), .Z(n11546) );
  NANDN U11840 ( .A(n11547), .B(n11546), .Z(n11169) );
  NAND U11841 ( .A(n11170), .B(n11169), .Z(n11174) );
  NAND U11842 ( .A(a[40]), .B(b[28]), .Z(n11173) );
  OR U11843 ( .A(n11174), .B(n11173), .Z(n11176) );
  XOR U11844 ( .A(n11172), .B(n11171), .Z(n11552) );
  XOR U11845 ( .A(n11174), .B(n11173), .Z(n11553) );
  NAND U11846 ( .A(n11552), .B(n11553), .Z(n11175) );
  NAND U11847 ( .A(n11176), .B(n11175), .Z(n11179) );
  AND U11848 ( .A(b[28]), .B(a[41]), .Z(n11180) );
  OR U11849 ( .A(n11179), .B(n11180), .Z(n11182) );
  XNOR U11850 ( .A(n11178), .B(n11177), .Z(n11559) );
  XOR U11851 ( .A(n11180), .B(n11179), .Z(n11558) );
  NANDN U11852 ( .A(n11559), .B(n11558), .Z(n11181) );
  NAND U11853 ( .A(n11182), .B(n11181), .Z(n11186) );
  NAND U11854 ( .A(a[42]), .B(b[28]), .Z(n11185) );
  OR U11855 ( .A(n11186), .B(n11185), .Z(n11188) );
  XOR U11856 ( .A(n11184), .B(n11183), .Z(n11564) );
  XOR U11857 ( .A(n11186), .B(n11185), .Z(n11565) );
  NAND U11858 ( .A(n11564), .B(n11565), .Z(n11187) );
  NAND U11859 ( .A(n11188), .B(n11187), .Z(n11191) );
  AND U11860 ( .A(b[28]), .B(a[43]), .Z(n11192) );
  OR U11861 ( .A(n11191), .B(n11192), .Z(n11194) );
  XNOR U11862 ( .A(n11190), .B(n11189), .Z(n11571) );
  XOR U11863 ( .A(n11192), .B(n11191), .Z(n11570) );
  NANDN U11864 ( .A(n11571), .B(n11570), .Z(n11193) );
  NAND U11865 ( .A(n11194), .B(n11193), .Z(n11198) );
  NAND U11866 ( .A(a[44]), .B(b[28]), .Z(n11197) );
  OR U11867 ( .A(n11198), .B(n11197), .Z(n11200) );
  XOR U11868 ( .A(n11196), .B(n11195), .Z(n11576) );
  XOR U11869 ( .A(n11198), .B(n11197), .Z(n11577) );
  NAND U11870 ( .A(n11576), .B(n11577), .Z(n11199) );
  NAND U11871 ( .A(n11200), .B(n11199), .Z(n11203) );
  AND U11872 ( .A(b[28]), .B(a[45]), .Z(n11204) );
  OR U11873 ( .A(n11203), .B(n11204), .Z(n11206) );
  XNOR U11874 ( .A(n11202), .B(n11201), .Z(n11583) );
  XOR U11875 ( .A(n11204), .B(n11203), .Z(n11582) );
  NANDN U11876 ( .A(n11583), .B(n11582), .Z(n11205) );
  NAND U11877 ( .A(n11206), .B(n11205), .Z(n11210) );
  NAND U11878 ( .A(a[46]), .B(b[28]), .Z(n11209) );
  OR U11879 ( .A(n11210), .B(n11209), .Z(n11212) );
  XOR U11880 ( .A(n11208), .B(n11207), .Z(n11588) );
  XOR U11881 ( .A(n11210), .B(n11209), .Z(n11589) );
  NAND U11882 ( .A(n11588), .B(n11589), .Z(n11211) );
  NAND U11883 ( .A(n11212), .B(n11211), .Z(n11215) );
  AND U11884 ( .A(b[28]), .B(a[47]), .Z(n11216) );
  OR U11885 ( .A(n11215), .B(n11216), .Z(n11218) );
  XNOR U11886 ( .A(n11214), .B(n11213), .Z(n11595) );
  XOR U11887 ( .A(n11216), .B(n11215), .Z(n11594) );
  NANDN U11888 ( .A(n11595), .B(n11594), .Z(n11217) );
  NAND U11889 ( .A(n11218), .B(n11217), .Z(n11222) );
  NAND U11890 ( .A(a[48]), .B(b[28]), .Z(n11221) );
  OR U11891 ( .A(n11222), .B(n11221), .Z(n11224) );
  XOR U11892 ( .A(n11220), .B(n11219), .Z(n11600) );
  XOR U11893 ( .A(n11222), .B(n11221), .Z(n11601) );
  NAND U11894 ( .A(n11600), .B(n11601), .Z(n11223) );
  NAND U11895 ( .A(n11224), .B(n11223), .Z(n11227) );
  AND U11896 ( .A(b[28]), .B(a[49]), .Z(n11228) );
  OR U11897 ( .A(n11227), .B(n11228), .Z(n11230) );
  XNOR U11898 ( .A(n11226), .B(n11225), .Z(n11607) );
  XOR U11899 ( .A(n11228), .B(n11227), .Z(n11606) );
  NANDN U11900 ( .A(n11607), .B(n11606), .Z(n11229) );
  NAND U11901 ( .A(n11230), .B(n11229), .Z(n11234) );
  NAND U11902 ( .A(a[50]), .B(b[28]), .Z(n11233) );
  OR U11903 ( .A(n11234), .B(n11233), .Z(n11236) );
  XOR U11904 ( .A(n11232), .B(n11231), .Z(n11612) );
  XOR U11905 ( .A(n11234), .B(n11233), .Z(n11613) );
  NAND U11906 ( .A(n11612), .B(n11613), .Z(n11235) );
  NAND U11907 ( .A(n11236), .B(n11235), .Z(n11239) );
  AND U11908 ( .A(b[28]), .B(a[51]), .Z(n11240) );
  OR U11909 ( .A(n11239), .B(n11240), .Z(n11242) );
  XNOR U11910 ( .A(n11238), .B(n11237), .Z(n11619) );
  XOR U11911 ( .A(n11240), .B(n11239), .Z(n11618) );
  NANDN U11912 ( .A(n11619), .B(n11618), .Z(n11241) );
  NAND U11913 ( .A(n11242), .B(n11241), .Z(n11246) );
  NAND U11914 ( .A(a[52]), .B(b[28]), .Z(n11245) );
  OR U11915 ( .A(n11246), .B(n11245), .Z(n11248) );
  XOR U11916 ( .A(n11244), .B(n11243), .Z(n11624) );
  XOR U11917 ( .A(n11246), .B(n11245), .Z(n11625) );
  NAND U11918 ( .A(n11624), .B(n11625), .Z(n11247) );
  NAND U11919 ( .A(n11248), .B(n11247), .Z(n11251) );
  AND U11920 ( .A(b[28]), .B(a[53]), .Z(n11252) );
  OR U11921 ( .A(n11251), .B(n11252), .Z(n11254) );
  XNOR U11922 ( .A(n11250), .B(n11249), .Z(n11631) );
  XOR U11923 ( .A(n11252), .B(n11251), .Z(n11630) );
  NANDN U11924 ( .A(n11631), .B(n11630), .Z(n11253) );
  NAND U11925 ( .A(n11254), .B(n11253), .Z(n11258) );
  NAND U11926 ( .A(a[54]), .B(b[28]), .Z(n11257) );
  OR U11927 ( .A(n11258), .B(n11257), .Z(n11260) );
  XOR U11928 ( .A(n11256), .B(n11255), .Z(n11636) );
  XOR U11929 ( .A(n11258), .B(n11257), .Z(n11637) );
  NAND U11930 ( .A(n11636), .B(n11637), .Z(n11259) );
  NAND U11931 ( .A(n11260), .B(n11259), .Z(n11263) );
  AND U11932 ( .A(b[28]), .B(a[55]), .Z(n11264) );
  OR U11933 ( .A(n11263), .B(n11264), .Z(n11266) );
  XNOR U11934 ( .A(n11262), .B(n11261), .Z(n11643) );
  XOR U11935 ( .A(n11264), .B(n11263), .Z(n11642) );
  NANDN U11936 ( .A(n11643), .B(n11642), .Z(n11265) );
  NAND U11937 ( .A(n11266), .B(n11265), .Z(n11270) );
  NAND U11938 ( .A(a[56]), .B(b[28]), .Z(n11269) );
  OR U11939 ( .A(n11270), .B(n11269), .Z(n11272) );
  XOR U11940 ( .A(n11268), .B(n11267), .Z(n11648) );
  XOR U11941 ( .A(n11270), .B(n11269), .Z(n11649) );
  NAND U11942 ( .A(n11648), .B(n11649), .Z(n11271) );
  NAND U11943 ( .A(n11272), .B(n11271), .Z(n11275) );
  AND U11944 ( .A(b[28]), .B(a[57]), .Z(n11276) );
  OR U11945 ( .A(n11275), .B(n11276), .Z(n11278) );
  XNOR U11946 ( .A(n11274), .B(n11273), .Z(n11655) );
  XOR U11947 ( .A(n11276), .B(n11275), .Z(n11654) );
  NANDN U11948 ( .A(n11655), .B(n11654), .Z(n11277) );
  NAND U11949 ( .A(n11278), .B(n11277), .Z(n11282) );
  NAND U11950 ( .A(a[58]), .B(b[28]), .Z(n11281) );
  OR U11951 ( .A(n11282), .B(n11281), .Z(n11284) );
  XOR U11952 ( .A(n11280), .B(n11279), .Z(n11660) );
  XOR U11953 ( .A(n11282), .B(n11281), .Z(n11661) );
  NAND U11954 ( .A(n11660), .B(n11661), .Z(n11283) );
  NAND U11955 ( .A(n11284), .B(n11283), .Z(n11287) );
  AND U11956 ( .A(b[28]), .B(a[59]), .Z(n11288) );
  OR U11957 ( .A(n11287), .B(n11288), .Z(n11290) );
  XNOR U11958 ( .A(n11286), .B(n11285), .Z(n11667) );
  XOR U11959 ( .A(n11288), .B(n11287), .Z(n11666) );
  NANDN U11960 ( .A(n11667), .B(n11666), .Z(n11289) );
  NAND U11961 ( .A(n11290), .B(n11289), .Z(n11294) );
  NAND U11962 ( .A(a[60]), .B(b[28]), .Z(n11293) );
  OR U11963 ( .A(n11294), .B(n11293), .Z(n11296) );
  XOR U11964 ( .A(n11292), .B(n11291), .Z(n11313) );
  XOR U11965 ( .A(n11294), .B(n11293), .Z(n11314) );
  NAND U11966 ( .A(n11313), .B(n11314), .Z(n11295) );
  NAND U11967 ( .A(n11296), .B(n11295), .Z(n11299) );
  AND U11968 ( .A(b[28]), .B(a[61]), .Z(n11300) );
  OR U11969 ( .A(n11299), .B(n11300), .Z(n11302) );
  XNOR U11970 ( .A(n11298), .B(n11297), .Z(n11677) );
  XOR U11971 ( .A(n11300), .B(n11299), .Z(n11676) );
  NANDN U11972 ( .A(n11677), .B(n11676), .Z(n11301) );
  NAND U11973 ( .A(n11302), .B(n11301), .Z(n11306) );
  NAND U11974 ( .A(a[62]), .B(b[28]), .Z(n11305) );
  OR U11975 ( .A(n11306), .B(n11305), .Z(n11308) );
  XOR U11976 ( .A(n11304), .B(n11303), .Z(n11309) );
  XOR U11977 ( .A(n11306), .B(n11305), .Z(n11310) );
  NAND U11978 ( .A(n11309), .B(n11310), .Z(n11307) );
  NAND U11979 ( .A(n11308), .B(n11307), .Z(n12066) );
  XOR U11980 ( .A(n12065), .B(n12066), .Z(n12067) );
  XNOR U11981 ( .A(n12068), .B(n12067), .Z(n12062) );
  NAND U11982 ( .A(a[63]), .B(b[27]), .Z(n11311) );
  XOR U11983 ( .A(n11310), .B(n11309), .Z(n11312) );
  NANDN U11984 ( .A(n11311), .B(n11312), .Z(n11683) );
  XOR U11985 ( .A(n11312), .B(n11311), .Z(n11684) );
  XOR U11986 ( .A(n11314), .B(n11313), .Z(n11673) );
  NAND U11987 ( .A(a[60]), .B(b[27]), .Z(n11669) );
  NAND U11988 ( .A(a[58]), .B(b[27]), .Z(n11657) );
  NAND U11989 ( .A(a[56]), .B(b[27]), .Z(n11645) );
  NAND U11990 ( .A(a[54]), .B(b[27]), .Z(n11633) );
  NAND U11991 ( .A(a[52]), .B(b[27]), .Z(n11621) );
  NAND U11992 ( .A(a[50]), .B(b[27]), .Z(n11609) );
  NAND U11993 ( .A(a[48]), .B(b[27]), .Z(n11597) );
  NAND U11994 ( .A(a[46]), .B(b[27]), .Z(n11585) );
  NAND U11995 ( .A(a[44]), .B(b[27]), .Z(n11573) );
  NAND U11996 ( .A(a[42]), .B(b[27]), .Z(n11561) );
  NAND U11997 ( .A(a[40]), .B(b[27]), .Z(n11549) );
  NAND U11998 ( .A(a[33]), .B(b[27]), .Z(n11505) );
  NAND U11999 ( .A(a[13]), .B(b[27]), .Z(n11385) );
  ANDN U12000 ( .B(b[27]), .A(n21164), .Z(n11372) );
  ANDN U12001 ( .B(b[27]), .A(n166), .Z(n11348) );
  XNOR U12002 ( .A(n11316), .B(n11315), .Z(n11345) );
  ANDN U12003 ( .B(b[27]), .A(n164), .Z(n11341) );
  ANDN U12004 ( .B(b[27]), .A(n21580), .Z(n11326) );
  NAND U12005 ( .A(b[28]), .B(a[1]), .Z(n11319) );
  AND U12006 ( .A(b[27]), .B(a[0]), .Z(n12081) );
  NANDN U12007 ( .A(n11319), .B(n12081), .Z(n11318) );
  NAND U12008 ( .A(a[2]), .B(b[27]), .Z(n11317) );
  AND U12009 ( .A(n11318), .B(n11317), .Z(n11325) );
  NANDN U12010 ( .A(n11319), .B(a[0]), .Z(n11320) );
  XNOR U12011 ( .A(a[2]), .B(n11320), .Z(n11321) );
  NAND U12012 ( .A(b[27]), .B(n11321), .Z(n11700) );
  AND U12013 ( .A(a[1]), .B(b[28]), .Z(n11322) );
  XNOR U12014 ( .A(n11323), .B(n11322), .Z(n11699) );
  NANDN U12015 ( .A(n11700), .B(n11699), .Z(n11324) );
  NANDN U12016 ( .A(n11325), .B(n11324), .Z(n11327) );
  NANDN U12017 ( .A(n11326), .B(n11327), .Z(n11331) );
  XOR U12018 ( .A(n11327), .B(n11326), .Z(n11704) );
  NANDN U12019 ( .A(n11704), .B(n11703), .Z(n11330) );
  NAND U12020 ( .A(n11331), .B(n11330), .Z(n11335) );
  XOR U12021 ( .A(n11333), .B(n11332), .Z(n11334) );
  NANDN U12022 ( .A(n11335), .B(n11334), .Z(n11337) );
  NAND U12023 ( .A(a[4]), .B(b[27]), .Z(n11709) );
  NANDN U12024 ( .A(n11709), .B(n11710), .Z(n11336) );
  NAND U12025 ( .A(n11337), .B(n11336), .Z(n11340) );
  OR U12026 ( .A(n11341), .B(n11340), .Z(n11343) );
  XOR U12027 ( .A(n11339), .B(n11338), .Z(n11687) );
  XOR U12028 ( .A(n11341), .B(n11340), .Z(n11686) );
  NAND U12029 ( .A(n11687), .B(n11686), .Z(n11342) );
  NAND U12030 ( .A(n11343), .B(n11342), .Z(n11344) );
  NANDN U12031 ( .A(n11345), .B(n11344), .Z(n11347) );
  ANDN U12032 ( .B(b[27]), .A(n165), .Z(n11722) );
  NANDN U12033 ( .A(n11722), .B(n11721), .Z(n11346) );
  NAND U12034 ( .A(n11347), .B(n11346), .Z(n11349) );
  NANDN U12035 ( .A(n11348), .B(n11349), .Z(n11353) );
  XOR U12036 ( .A(n11349), .B(n11348), .Z(n11726) );
  XOR U12037 ( .A(n11351), .B(n11350), .Z(n11725) );
  OR U12038 ( .A(n11726), .B(n11725), .Z(n11352) );
  NAND U12039 ( .A(n11353), .B(n11352), .Z(n11357) );
  XOR U12040 ( .A(n11355), .B(n11354), .Z(n11356) );
  NANDN U12041 ( .A(n11357), .B(n11356), .Z(n11359) );
  NAND U12042 ( .A(a[8]), .B(b[27]), .Z(n11733) );
  NANDN U12043 ( .A(n11733), .B(n11734), .Z(n11358) );
  NAND U12044 ( .A(n11359), .B(n11358), .Z(n11360) );
  ANDN U12045 ( .B(b[27]), .A(n21615), .Z(n11361) );
  OR U12046 ( .A(n11360), .B(n11361), .Z(n11365) );
  XNOR U12047 ( .A(n11361), .B(n11360), .Z(n11737) );
  OR U12048 ( .A(n11737), .B(n11738), .Z(n11364) );
  AND U12049 ( .A(n11365), .B(n11364), .Z(n11369) );
  XOR U12050 ( .A(n11367), .B(n11366), .Z(n11368) );
  NANDN U12051 ( .A(n11369), .B(n11368), .Z(n11371) );
  XOR U12052 ( .A(n11369), .B(n11368), .Z(n11745) );
  ANDN U12053 ( .B(b[27]), .A(n168), .Z(n11746) );
  OR U12054 ( .A(n11745), .B(n11746), .Z(n11370) );
  AND U12055 ( .A(n11371), .B(n11370), .Z(n11373) );
  OR U12056 ( .A(n11372), .B(n11373), .Z(n11377) );
  XNOR U12057 ( .A(n11373), .B(n11372), .Z(n11750) );
  XNOR U12058 ( .A(n11375), .B(n11374), .Z(n11749) );
  OR U12059 ( .A(n11750), .B(n11749), .Z(n11376) );
  AND U12060 ( .A(n11377), .B(n11376), .Z(n11380) );
  OR U12061 ( .A(n11380), .B(n11381), .Z(n11383) );
  ANDN U12062 ( .B(b[27]), .A(n169), .Z(n11758) );
  XOR U12063 ( .A(n11381), .B(n11380), .Z(n11757) );
  NANDN U12064 ( .A(n11758), .B(n11757), .Z(n11382) );
  NAND U12065 ( .A(n11383), .B(n11382), .Z(n11384) );
  OR U12066 ( .A(n11385), .B(n11384), .Z(n11389) );
  XNOR U12067 ( .A(n11385), .B(n11384), .Z(n11762) );
  XNOR U12068 ( .A(n11387), .B(n11386), .Z(n11761) );
  NANDN U12069 ( .A(n11762), .B(n11761), .Z(n11388) );
  AND U12070 ( .A(n11389), .B(n11388), .Z(n11392) );
  XNOR U12071 ( .A(n11391), .B(n11390), .Z(n11393) );
  OR U12072 ( .A(n11392), .B(n11393), .Z(n11395) );
  XNOR U12073 ( .A(n11393), .B(n11392), .Z(n11770) );
  AND U12074 ( .A(b[27]), .B(a[14]), .Z(n11769) );
  NANDN U12075 ( .A(n11770), .B(n11769), .Z(n11394) );
  NAND U12076 ( .A(n11395), .B(n11394), .Z(n11398) );
  ANDN U12077 ( .B(b[27]), .A(n172), .Z(n11399) );
  OR U12078 ( .A(n11398), .B(n11399), .Z(n11401) );
  XOR U12079 ( .A(n11397), .B(n11396), .Z(n11774) );
  XOR U12080 ( .A(n11399), .B(n11398), .Z(n11773) );
  NANDN U12081 ( .A(n11774), .B(n11773), .Z(n11400) );
  NAND U12082 ( .A(n11401), .B(n11400), .Z(n11404) );
  XNOR U12083 ( .A(n11403), .B(n11402), .Z(n11405) );
  OR U12084 ( .A(n11404), .B(n11405), .Z(n11407) );
  XNOR U12085 ( .A(n11405), .B(n11404), .Z(n11780) );
  NAND U12086 ( .A(a[16]), .B(b[27]), .Z(n11779) );
  OR U12087 ( .A(n11780), .B(n11779), .Z(n11406) );
  NAND U12088 ( .A(n11407), .B(n11406), .Z(n11410) );
  ANDN U12089 ( .B(b[27]), .A(n174), .Z(n11411) );
  OR U12090 ( .A(n11410), .B(n11411), .Z(n11413) );
  XOR U12091 ( .A(n11409), .B(n11408), .Z(n11786) );
  XOR U12092 ( .A(n11411), .B(n11410), .Z(n11785) );
  NANDN U12093 ( .A(n11786), .B(n11785), .Z(n11412) );
  NAND U12094 ( .A(n11413), .B(n11412), .Z(n11416) );
  XNOR U12095 ( .A(n11415), .B(n11414), .Z(n11417) );
  OR U12096 ( .A(n11416), .B(n11417), .Z(n11419) );
  XNOR U12097 ( .A(n11417), .B(n11416), .Z(n11792) );
  NAND U12098 ( .A(a[18]), .B(b[27]), .Z(n11791) );
  OR U12099 ( .A(n11792), .B(n11791), .Z(n11418) );
  NAND U12100 ( .A(n11419), .B(n11418), .Z(n11422) );
  ANDN U12101 ( .B(b[27]), .A(n21670), .Z(n11423) );
  OR U12102 ( .A(n11422), .B(n11423), .Z(n11425) );
  XOR U12103 ( .A(n11421), .B(n11420), .Z(n11798) );
  XOR U12104 ( .A(n11423), .B(n11422), .Z(n11797) );
  NANDN U12105 ( .A(n11798), .B(n11797), .Z(n11424) );
  NAND U12106 ( .A(n11425), .B(n11424), .Z(n11428) );
  XNOR U12107 ( .A(n11427), .B(n11426), .Z(n11429) );
  OR U12108 ( .A(n11428), .B(n11429), .Z(n11431) );
  XNOR U12109 ( .A(n11429), .B(n11428), .Z(n11804) );
  NAND U12110 ( .A(a[20]), .B(b[27]), .Z(n11803) );
  OR U12111 ( .A(n11804), .B(n11803), .Z(n11430) );
  NAND U12112 ( .A(n11431), .B(n11430), .Z(n11434) );
  ANDN U12113 ( .B(b[27]), .A(n21681), .Z(n11435) );
  OR U12114 ( .A(n11434), .B(n11435), .Z(n11437) );
  XOR U12115 ( .A(n11433), .B(n11432), .Z(n11810) );
  XOR U12116 ( .A(n11435), .B(n11434), .Z(n11809) );
  NANDN U12117 ( .A(n11810), .B(n11809), .Z(n11436) );
  NAND U12118 ( .A(n11437), .B(n11436), .Z(n11440) );
  XNOR U12119 ( .A(n11439), .B(n11438), .Z(n11441) );
  OR U12120 ( .A(n11440), .B(n11441), .Z(n11443) );
  XNOR U12121 ( .A(n11441), .B(n11440), .Z(n11816) );
  NAND U12122 ( .A(a[22]), .B(b[27]), .Z(n11815) );
  OR U12123 ( .A(n11816), .B(n11815), .Z(n11442) );
  NAND U12124 ( .A(n11443), .B(n11442), .Z(n11446) );
  ANDN U12125 ( .B(b[27]), .A(n21692), .Z(n11447) );
  OR U12126 ( .A(n11446), .B(n11447), .Z(n11449) );
  XOR U12127 ( .A(n11445), .B(n11444), .Z(n11822) );
  XOR U12128 ( .A(n11447), .B(n11446), .Z(n11821) );
  NANDN U12129 ( .A(n11822), .B(n11821), .Z(n11448) );
  NAND U12130 ( .A(n11449), .B(n11448), .Z(n11452) );
  XNOR U12131 ( .A(n11451), .B(n11450), .Z(n11453) );
  OR U12132 ( .A(n11452), .B(n11453), .Z(n11455) );
  XNOR U12133 ( .A(n11453), .B(n11452), .Z(n11828) );
  NAND U12134 ( .A(a[24]), .B(b[27]), .Z(n11827) );
  OR U12135 ( .A(n11828), .B(n11827), .Z(n11454) );
  NAND U12136 ( .A(n11455), .B(n11454), .Z(n11458) );
  ANDN U12137 ( .B(b[27]), .A(n21703), .Z(n11459) );
  OR U12138 ( .A(n11458), .B(n11459), .Z(n11461) );
  XOR U12139 ( .A(n11457), .B(n11456), .Z(n11834) );
  XOR U12140 ( .A(n11459), .B(n11458), .Z(n11833) );
  NANDN U12141 ( .A(n11834), .B(n11833), .Z(n11460) );
  NAND U12142 ( .A(n11461), .B(n11460), .Z(n11464) );
  XNOR U12143 ( .A(n11463), .B(n11462), .Z(n11465) );
  OR U12144 ( .A(n11464), .B(n11465), .Z(n11467) );
  XNOR U12145 ( .A(n11465), .B(n11464), .Z(n11840) );
  NAND U12146 ( .A(a[26]), .B(b[27]), .Z(n11839) );
  OR U12147 ( .A(n11840), .B(n11839), .Z(n11466) );
  NAND U12148 ( .A(n11467), .B(n11466), .Z(n11470) );
  ANDN U12149 ( .B(b[27]), .A(n21716), .Z(n11471) );
  OR U12150 ( .A(n11470), .B(n11471), .Z(n11473) );
  XOR U12151 ( .A(n11469), .B(n11468), .Z(n11846) );
  XOR U12152 ( .A(n11471), .B(n11470), .Z(n11845) );
  NANDN U12153 ( .A(n11846), .B(n11845), .Z(n11472) );
  NAND U12154 ( .A(n11473), .B(n11472), .Z(n11476) );
  XNOR U12155 ( .A(n11475), .B(n11474), .Z(n11477) );
  OR U12156 ( .A(n11476), .B(n11477), .Z(n11479) );
  XNOR U12157 ( .A(n11477), .B(n11476), .Z(n11852) );
  NAND U12158 ( .A(a[28]), .B(b[27]), .Z(n11851) );
  OR U12159 ( .A(n11852), .B(n11851), .Z(n11478) );
  NAND U12160 ( .A(n11479), .B(n11478), .Z(n11482) );
  ANDN U12161 ( .B(b[27]), .A(n21727), .Z(n11483) );
  OR U12162 ( .A(n11482), .B(n11483), .Z(n11485) );
  XOR U12163 ( .A(n11483), .B(n11482), .Z(n11857) );
  NANDN U12164 ( .A(n11858), .B(n11857), .Z(n11484) );
  NAND U12165 ( .A(n11485), .B(n11484), .Z(n11488) );
  XOR U12166 ( .A(n11487), .B(n11486), .Z(n11489) );
  OR U12167 ( .A(n11488), .B(n11489), .Z(n11491) );
  NAND U12168 ( .A(a[30]), .B(b[27]), .Z(n11864) );
  XOR U12169 ( .A(n11489), .B(n11488), .Z(n11863) );
  NANDN U12170 ( .A(n11864), .B(n11863), .Z(n11490) );
  NAND U12171 ( .A(n11491), .B(n11490), .Z(n11494) );
  ANDN U12172 ( .B(b[27]), .A(n21740), .Z(n11495) );
  OR U12173 ( .A(n11494), .B(n11495), .Z(n11497) );
  XOR U12174 ( .A(n11495), .B(n11494), .Z(n11869) );
  NANDN U12175 ( .A(n11870), .B(n11869), .Z(n11496) );
  AND U12176 ( .A(n11497), .B(n11496), .Z(n11501) );
  XOR U12177 ( .A(n11499), .B(n11498), .Z(n11500) );
  NANDN U12178 ( .A(n11501), .B(n11500), .Z(n11503) );
  XOR U12179 ( .A(n11501), .B(n11500), .Z(n11877) );
  ANDN U12180 ( .B(b[27]), .A(n182), .Z(n11878) );
  OR U12181 ( .A(n11877), .B(n11878), .Z(n11502) );
  NAND U12182 ( .A(n11503), .B(n11502), .Z(n11504) );
  OR U12183 ( .A(n11505), .B(n11504), .Z(n11509) );
  XNOR U12184 ( .A(n11505), .B(n11504), .Z(n11882) );
  XNOR U12185 ( .A(n11507), .B(n11506), .Z(n11881) );
  NANDN U12186 ( .A(n11882), .B(n11881), .Z(n11508) );
  AND U12187 ( .A(n11509), .B(n11508), .Z(n11512) );
  XNOR U12188 ( .A(n11511), .B(n11510), .Z(n11513) );
  OR U12189 ( .A(n11512), .B(n11513), .Z(n11515) );
  XNOR U12190 ( .A(n11513), .B(n11512), .Z(n11890) );
  AND U12191 ( .A(b[27]), .B(a[34]), .Z(n11889) );
  NANDN U12192 ( .A(n11890), .B(n11889), .Z(n11514) );
  NAND U12193 ( .A(n11515), .B(n11514), .Z(n11518) );
  ANDN U12194 ( .B(b[27]), .A(n184), .Z(n11519) );
  OR U12195 ( .A(n11518), .B(n11519), .Z(n11521) );
  XOR U12196 ( .A(n11517), .B(n11516), .Z(n11894) );
  XOR U12197 ( .A(n11519), .B(n11518), .Z(n11893) );
  NANDN U12198 ( .A(n11894), .B(n11893), .Z(n11520) );
  NAND U12199 ( .A(n11521), .B(n11520), .Z(n11524) );
  XNOR U12200 ( .A(n11523), .B(n11522), .Z(n11525) );
  OR U12201 ( .A(n11524), .B(n11525), .Z(n11527) );
  XNOR U12202 ( .A(n11525), .B(n11524), .Z(n11900) );
  NAND U12203 ( .A(a[36]), .B(b[27]), .Z(n11899) );
  OR U12204 ( .A(n11900), .B(n11899), .Z(n11526) );
  NAND U12205 ( .A(n11527), .B(n11526), .Z(n11528) );
  ANDN U12206 ( .B(b[27]), .A(n21772), .Z(n11529) );
  OR U12207 ( .A(n11528), .B(n11529), .Z(n11533) );
  XOR U12208 ( .A(n11529), .B(n11528), .Z(n11905) );
  NAND U12209 ( .A(n11905), .B(n11906), .Z(n11532) );
  NAND U12210 ( .A(n11533), .B(n11532), .Z(n11535) );
  NAND U12211 ( .A(a[38]), .B(b[27]), .Z(n11534) );
  OR U12212 ( .A(n11535), .B(n11534), .Z(n11539) );
  XOR U12213 ( .A(n11535), .B(n11534), .Z(n11911) );
  XOR U12214 ( .A(n11537), .B(n11536), .Z(n11912) );
  NAND U12215 ( .A(n11911), .B(n11912), .Z(n11538) );
  NAND U12216 ( .A(n11539), .B(n11538), .Z(n11543) );
  XOR U12217 ( .A(n11541), .B(n11540), .Z(n11542) );
  NAND U12218 ( .A(n11543), .B(n11542), .Z(n11545) );
  XNOR U12219 ( .A(n11543), .B(n11542), .Z(n11920) );
  NAND U12220 ( .A(a[39]), .B(b[27]), .Z(n11919) );
  OR U12221 ( .A(n11920), .B(n11919), .Z(n11544) );
  NAND U12222 ( .A(n11545), .B(n11544), .Z(n11548) );
  NANDN U12223 ( .A(n11549), .B(n11548), .Z(n11551) );
  XNOR U12224 ( .A(n11547), .B(n11546), .Z(n11924) );
  NANDN U12225 ( .A(n11924), .B(n11923), .Z(n11550) );
  NAND U12226 ( .A(n11551), .B(n11550), .Z(n11555) );
  XOR U12227 ( .A(n11553), .B(n11552), .Z(n11554) );
  NAND U12228 ( .A(n11555), .B(n11554), .Z(n11557) );
  XNOR U12229 ( .A(n11555), .B(n11554), .Z(n11932) );
  NAND U12230 ( .A(a[41]), .B(b[27]), .Z(n11931) );
  OR U12231 ( .A(n11932), .B(n11931), .Z(n11556) );
  NAND U12232 ( .A(n11557), .B(n11556), .Z(n11560) );
  NANDN U12233 ( .A(n11561), .B(n11560), .Z(n11563) );
  XNOR U12234 ( .A(n11559), .B(n11558), .Z(n11936) );
  NANDN U12235 ( .A(n11936), .B(n11935), .Z(n11562) );
  NAND U12236 ( .A(n11563), .B(n11562), .Z(n11567) );
  XOR U12237 ( .A(n11565), .B(n11564), .Z(n11566) );
  NAND U12238 ( .A(n11567), .B(n11566), .Z(n11569) );
  XNOR U12239 ( .A(n11567), .B(n11566), .Z(n11944) );
  NAND U12240 ( .A(a[43]), .B(b[27]), .Z(n11943) );
  OR U12241 ( .A(n11944), .B(n11943), .Z(n11568) );
  NAND U12242 ( .A(n11569), .B(n11568), .Z(n11572) );
  NANDN U12243 ( .A(n11573), .B(n11572), .Z(n11575) );
  XNOR U12244 ( .A(n11571), .B(n11570), .Z(n11948) );
  NANDN U12245 ( .A(n11948), .B(n11947), .Z(n11574) );
  NAND U12246 ( .A(n11575), .B(n11574), .Z(n11579) );
  XOR U12247 ( .A(n11577), .B(n11576), .Z(n11578) );
  NAND U12248 ( .A(n11579), .B(n11578), .Z(n11581) );
  XNOR U12249 ( .A(n11579), .B(n11578), .Z(n11956) );
  NAND U12250 ( .A(a[45]), .B(b[27]), .Z(n11955) );
  OR U12251 ( .A(n11956), .B(n11955), .Z(n11580) );
  NAND U12252 ( .A(n11581), .B(n11580), .Z(n11584) );
  NANDN U12253 ( .A(n11585), .B(n11584), .Z(n11587) );
  XNOR U12254 ( .A(n11583), .B(n11582), .Z(n11960) );
  NANDN U12255 ( .A(n11960), .B(n11959), .Z(n11586) );
  NAND U12256 ( .A(n11587), .B(n11586), .Z(n11591) );
  XOR U12257 ( .A(n11589), .B(n11588), .Z(n11590) );
  NAND U12258 ( .A(n11591), .B(n11590), .Z(n11593) );
  XNOR U12259 ( .A(n11591), .B(n11590), .Z(n11968) );
  NAND U12260 ( .A(a[47]), .B(b[27]), .Z(n11967) );
  OR U12261 ( .A(n11968), .B(n11967), .Z(n11592) );
  NAND U12262 ( .A(n11593), .B(n11592), .Z(n11596) );
  NANDN U12263 ( .A(n11597), .B(n11596), .Z(n11599) );
  XNOR U12264 ( .A(n11595), .B(n11594), .Z(n11972) );
  NANDN U12265 ( .A(n11972), .B(n11971), .Z(n11598) );
  NAND U12266 ( .A(n11599), .B(n11598), .Z(n11603) );
  XOR U12267 ( .A(n11601), .B(n11600), .Z(n11602) );
  NAND U12268 ( .A(n11603), .B(n11602), .Z(n11605) );
  XNOR U12269 ( .A(n11603), .B(n11602), .Z(n11980) );
  NAND U12270 ( .A(a[49]), .B(b[27]), .Z(n11979) );
  OR U12271 ( .A(n11980), .B(n11979), .Z(n11604) );
  NAND U12272 ( .A(n11605), .B(n11604), .Z(n11608) );
  NANDN U12273 ( .A(n11609), .B(n11608), .Z(n11611) );
  XNOR U12274 ( .A(n11607), .B(n11606), .Z(n11984) );
  NANDN U12275 ( .A(n11984), .B(n11983), .Z(n11610) );
  NAND U12276 ( .A(n11611), .B(n11610), .Z(n11615) );
  XOR U12277 ( .A(n11613), .B(n11612), .Z(n11614) );
  NAND U12278 ( .A(n11615), .B(n11614), .Z(n11617) );
  XNOR U12279 ( .A(n11615), .B(n11614), .Z(n11992) );
  NAND U12280 ( .A(a[51]), .B(b[27]), .Z(n11991) );
  OR U12281 ( .A(n11992), .B(n11991), .Z(n11616) );
  NAND U12282 ( .A(n11617), .B(n11616), .Z(n11620) );
  NANDN U12283 ( .A(n11621), .B(n11620), .Z(n11623) );
  XNOR U12284 ( .A(n11619), .B(n11618), .Z(n11996) );
  NANDN U12285 ( .A(n11996), .B(n11995), .Z(n11622) );
  NAND U12286 ( .A(n11623), .B(n11622), .Z(n11627) );
  XOR U12287 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U12288 ( .A(n11627), .B(n11626), .Z(n11629) );
  XNOR U12289 ( .A(n11627), .B(n11626), .Z(n12004) );
  NAND U12290 ( .A(a[53]), .B(b[27]), .Z(n12003) );
  OR U12291 ( .A(n12004), .B(n12003), .Z(n11628) );
  NAND U12292 ( .A(n11629), .B(n11628), .Z(n11632) );
  NANDN U12293 ( .A(n11633), .B(n11632), .Z(n11635) );
  XNOR U12294 ( .A(n11631), .B(n11630), .Z(n12008) );
  NANDN U12295 ( .A(n12008), .B(n12007), .Z(n11634) );
  NAND U12296 ( .A(n11635), .B(n11634), .Z(n11639) );
  XOR U12297 ( .A(n11637), .B(n11636), .Z(n11638) );
  NAND U12298 ( .A(n11639), .B(n11638), .Z(n11641) );
  XNOR U12299 ( .A(n11639), .B(n11638), .Z(n12016) );
  NAND U12300 ( .A(a[55]), .B(b[27]), .Z(n12015) );
  OR U12301 ( .A(n12016), .B(n12015), .Z(n11640) );
  NAND U12302 ( .A(n11641), .B(n11640), .Z(n11644) );
  NANDN U12303 ( .A(n11645), .B(n11644), .Z(n11647) );
  XNOR U12304 ( .A(n11643), .B(n11642), .Z(n12020) );
  NANDN U12305 ( .A(n12020), .B(n12019), .Z(n11646) );
  NAND U12306 ( .A(n11647), .B(n11646), .Z(n11651) );
  XOR U12307 ( .A(n11649), .B(n11648), .Z(n11650) );
  NAND U12308 ( .A(n11651), .B(n11650), .Z(n11653) );
  XNOR U12309 ( .A(n11651), .B(n11650), .Z(n12028) );
  NAND U12310 ( .A(a[57]), .B(b[27]), .Z(n12027) );
  OR U12311 ( .A(n12028), .B(n12027), .Z(n11652) );
  NAND U12312 ( .A(n11653), .B(n11652), .Z(n11656) );
  NANDN U12313 ( .A(n11657), .B(n11656), .Z(n11659) );
  XNOR U12314 ( .A(n11655), .B(n11654), .Z(n12032) );
  NANDN U12315 ( .A(n12032), .B(n12031), .Z(n11658) );
  NAND U12316 ( .A(n11659), .B(n11658), .Z(n11663) );
  XOR U12317 ( .A(n11661), .B(n11660), .Z(n11662) );
  NAND U12318 ( .A(n11663), .B(n11662), .Z(n11665) );
  XNOR U12319 ( .A(n11663), .B(n11662), .Z(n12040) );
  NAND U12320 ( .A(a[59]), .B(b[27]), .Z(n12039) );
  OR U12321 ( .A(n12040), .B(n12039), .Z(n11664) );
  NAND U12322 ( .A(n11665), .B(n11664), .Z(n11668) );
  NANDN U12323 ( .A(n11669), .B(n11668), .Z(n11671) );
  XNOR U12324 ( .A(n11667), .B(n11666), .Z(n12046) );
  NANDN U12325 ( .A(n12046), .B(n12045), .Z(n11670) );
  NAND U12326 ( .A(n11671), .B(n11670), .Z(n11672) );
  OR U12327 ( .A(n11673), .B(n11672), .Z(n11675) );
  ANDN U12328 ( .B(b[27]), .A(n209), .Z(n12050) );
  XOR U12329 ( .A(n11673), .B(n11672), .Z(n12049) );
  NANDN U12330 ( .A(n12050), .B(n12049), .Z(n11674) );
  NAND U12331 ( .A(n11675), .B(n11674), .Z(n11679) );
  NAND U12332 ( .A(a[62]), .B(b[27]), .Z(n11678) );
  OR U12333 ( .A(n11679), .B(n11678), .Z(n11681) );
  XNOR U12334 ( .A(n11677), .B(n11676), .Z(n12058) );
  XOR U12335 ( .A(n11679), .B(n11678), .Z(n12057) );
  NANDN U12336 ( .A(n12058), .B(n12057), .Z(n11680) );
  NAND U12337 ( .A(n11681), .B(n11680), .Z(n11685) );
  NANDN U12338 ( .A(n11684), .B(n11685), .Z(n11682) );
  AND U12339 ( .A(n11683), .B(n11682), .Z(n12061) );
  XNOR U12340 ( .A(n12062), .B(n12061), .Z(n21974) );
  XOR U12341 ( .A(n11685), .B(n11684), .Z(n12449) );
  ANDN U12342 ( .B(b[26]), .A(n210), .Z(n12056) );
  ANDN U12343 ( .B(b[26]), .A(n209), .Z(n12044) );
  ANDN U12344 ( .B(b[26]), .A(n207), .Z(n12034) );
  ANDN U12345 ( .B(b[26]), .A(n205), .Z(n12022) );
  ANDN U12346 ( .B(b[26]), .A(n203), .Z(n12010) );
  ANDN U12347 ( .B(b[26]), .A(n201), .Z(n11998) );
  ANDN U12348 ( .B(b[26]), .A(n199), .Z(n11986) );
  ANDN U12349 ( .B(b[26]), .A(n197), .Z(n11974) );
  ANDN U12350 ( .B(b[26]), .A(n195), .Z(n11962) );
  ANDN U12351 ( .B(b[26]), .A(n193), .Z(n11950) );
  ANDN U12352 ( .B(b[26]), .A(n191), .Z(n11938) );
  ANDN U12353 ( .B(b[26]), .A(n189), .Z(n11926) );
  NAND U12354 ( .A(a[40]), .B(b[26]), .Z(n11918) );
  NAND U12355 ( .A(a[35]), .B(b[26]), .Z(n11888) );
  NAND U12356 ( .A(a[15]), .B(b[26]), .Z(n11768) );
  ANDN U12357 ( .B(b[26]), .A(n21164), .Z(n11743) );
  ANDN U12358 ( .B(b[26]), .A(n21615), .Z(n11732) );
  ANDN U12359 ( .B(b[26]), .A(n166), .Z(n11719) );
  XNOR U12360 ( .A(n11687), .B(n11686), .Z(n11716) );
  ANDN U12361 ( .B(b[26]), .A(n164), .Z(n11712) );
  ANDN U12362 ( .B(b[26]), .A(n21580), .Z(n11697) );
  NAND U12363 ( .A(b[27]), .B(a[1]), .Z(n11690) );
  AND U12364 ( .A(b[26]), .B(a[0]), .Z(n12460) );
  NANDN U12365 ( .A(n11690), .B(n12460), .Z(n11689) );
  NAND U12366 ( .A(a[2]), .B(b[26]), .Z(n11688) );
  AND U12367 ( .A(n11689), .B(n11688), .Z(n11696) );
  NANDN U12368 ( .A(n11690), .B(a[0]), .Z(n11691) );
  XNOR U12369 ( .A(a[2]), .B(n11691), .Z(n11692) );
  NAND U12370 ( .A(b[26]), .B(n11692), .Z(n12087) );
  AND U12371 ( .A(a[1]), .B(b[27]), .Z(n11693) );
  XNOR U12372 ( .A(n11694), .B(n11693), .Z(n12086) );
  NANDN U12373 ( .A(n12087), .B(n12086), .Z(n11695) );
  NANDN U12374 ( .A(n11696), .B(n11695), .Z(n11698) );
  NANDN U12375 ( .A(n11697), .B(n11698), .Z(n11702) );
  XOR U12376 ( .A(n11698), .B(n11697), .Z(n12091) );
  NANDN U12377 ( .A(n12091), .B(n12090), .Z(n11701) );
  NAND U12378 ( .A(n11702), .B(n11701), .Z(n11706) );
  XOR U12379 ( .A(n11704), .B(n11703), .Z(n11705) );
  NANDN U12380 ( .A(n11706), .B(n11705), .Z(n11708) );
  NAND U12381 ( .A(a[4]), .B(b[26]), .Z(n12096) );
  NANDN U12382 ( .A(n12096), .B(n12097), .Z(n11707) );
  NAND U12383 ( .A(n11708), .B(n11707), .Z(n11711) );
  OR U12384 ( .A(n11712), .B(n11711), .Z(n11714) );
  XOR U12385 ( .A(n11710), .B(n11709), .Z(n12074) );
  XOR U12386 ( .A(n11712), .B(n11711), .Z(n12073) );
  NAND U12387 ( .A(n12074), .B(n12073), .Z(n11713) );
  NAND U12388 ( .A(n11714), .B(n11713), .Z(n11715) );
  NANDN U12389 ( .A(n11716), .B(n11715), .Z(n11718) );
  ANDN U12390 ( .B(b[26]), .A(n165), .Z(n12109) );
  NANDN U12391 ( .A(n12109), .B(n12108), .Z(n11717) );
  NAND U12392 ( .A(n11718), .B(n11717), .Z(n11720) );
  NANDN U12393 ( .A(n11719), .B(n11720), .Z(n11724) );
  XOR U12394 ( .A(n11720), .B(n11719), .Z(n12113) );
  XOR U12395 ( .A(n11722), .B(n11721), .Z(n12112) );
  OR U12396 ( .A(n12113), .B(n12112), .Z(n11723) );
  NAND U12397 ( .A(n11724), .B(n11723), .Z(n11728) );
  XNOR U12398 ( .A(n11726), .B(n11725), .Z(n11727) );
  NANDN U12399 ( .A(n11728), .B(n11727), .Z(n11730) );
  NAND U12400 ( .A(a[8]), .B(b[26]), .Z(n12120) );
  NANDN U12401 ( .A(n12120), .B(n12121), .Z(n11729) );
  NAND U12402 ( .A(n11730), .B(n11729), .Z(n11731) );
  OR U12403 ( .A(n11732), .B(n11731), .Z(n11736) );
  XNOR U12404 ( .A(n11732), .B(n11731), .Z(n12124) );
  XOR U12405 ( .A(n11734), .B(n11733), .Z(n12125) );
  NANDN U12406 ( .A(n12124), .B(n12125), .Z(n11735) );
  NAND U12407 ( .A(n11736), .B(n11735), .Z(n11740) );
  XOR U12408 ( .A(n11738), .B(n11737), .Z(n11739) );
  NAND U12409 ( .A(n11740), .B(n11739), .Z(n11742) );
  ANDN U12410 ( .B(b[26]), .A(n168), .Z(n12133) );
  XNOR U12411 ( .A(n11740), .B(n11739), .Z(n12132) );
  OR U12412 ( .A(n12133), .B(n12132), .Z(n11741) );
  NAND U12413 ( .A(n11742), .B(n11741), .Z(n11744) );
  NANDN U12414 ( .A(n11743), .B(n11744), .Z(n11748) );
  XOR U12415 ( .A(n11744), .B(n11743), .Z(n12137) );
  XNOR U12416 ( .A(n11746), .B(n11745), .Z(n12136) );
  OR U12417 ( .A(n12137), .B(n12136), .Z(n11747) );
  NAND U12418 ( .A(n11748), .B(n11747), .Z(n11751) );
  XNOR U12419 ( .A(n11750), .B(n11749), .Z(n11752) );
  NANDN U12420 ( .A(n11751), .B(n11752), .Z(n11754) );
  NAND U12421 ( .A(a[12]), .B(b[26]), .Z(n12144) );
  XNOR U12422 ( .A(n11752), .B(n11751), .Z(n12145) );
  NANDN U12423 ( .A(n12144), .B(n12145), .Z(n11753) );
  NAND U12424 ( .A(n11754), .B(n11753), .Z(n11755) );
  ANDN U12425 ( .B(b[26]), .A(n170), .Z(n11756) );
  OR U12426 ( .A(n11755), .B(n11756), .Z(n11760) );
  XNOR U12427 ( .A(n11756), .B(n11755), .Z(n12149) );
  OR U12428 ( .A(n12149), .B(n12148), .Z(n11759) );
  AND U12429 ( .A(n11760), .B(n11759), .Z(n11763) );
  OR U12430 ( .A(n11763), .B(n11764), .Z(n11766) );
  ANDN U12431 ( .B(b[26]), .A(n171), .Z(n12157) );
  XOR U12432 ( .A(n11764), .B(n11763), .Z(n12156) );
  NANDN U12433 ( .A(n12157), .B(n12156), .Z(n11765) );
  NAND U12434 ( .A(n11766), .B(n11765), .Z(n11767) );
  OR U12435 ( .A(n11768), .B(n11767), .Z(n11772) );
  XNOR U12436 ( .A(n11768), .B(n11767), .Z(n12161) );
  XNOR U12437 ( .A(n11770), .B(n11769), .Z(n12160) );
  NANDN U12438 ( .A(n12161), .B(n12160), .Z(n11771) );
  AND U12439 ( .A(n11772), .B(n11771), .Z(n11775) );
  XNOR U12440 ( .A(n11774), .B(n11773), .Z(n11776) );
  OR U12441 ( .A(n11775), .B(n11776), .Z(n11778) );
  XNOR U12442 ( .A(n11776), .B(n11775), .Z(n12169) );
  AND U12443 ( .A(b[26]), .B(a[16]), .Z(n12168) );
  NANDN U12444 ( .A(n12169), .B(n12168), .Z(n11777) );
  NAND U12445 ( .A(n11778), .B(n11777), .Z(n11781) );
  ANDN U12446 ( .B(b[26]), .A(n174), .Z(n11782) );
  OR U12447 ( .A(n11781), .B(n11782), .Z(n11784) );
  XOR U12448 ( .A(n11780), .B(n11779), .Z(n12173) );
  XOR U12449 ( .A(n11782), .B(n11781), .Z(n12172) );
  NANDN U12450 ( .A(n12173), .B(n12172), .Z(n11783) );
  NAND U12451 ( .A(n11784), .B(n11783), .Z(n11787) );
  XNOR U12452 ( .A(n11786), .B(n11785), .Z(n11788) );
  OR U12453 ( .A(n11787), .B(n11788), .Z(n11790) );
  XNOR U12454 ( .A(n11788), .B(n11787), .Z(n12179) );
  NAND U12455 ( .A(a[18]), .B(b[26]), .Z(n12178) );
  OR U12456 ( .A(n12179), .B(n12178), .Z(n11789) );
  NAND U12457 ( .A(n11790), .B(n11789), .Z(n11793) );
  ANDN U12458 ( .B(b[26]), .A(n21670), .Z(n11794) );
  OR U12459 ( .A(n11793), .B(n11794), .Z(n11796) );
  XOR U12460 ( .A(n11792), .B(n11791), .Z(n12185) );
  XOR U12461 ( .A(n11794), .B(n11793), .Z(n12184) );
  NANDN U12462 ( .A(n12185), .B(n12184), .Z(n11795) );
  NAND U12463 ( .A(n11796), .B(n11795), .Z(n11799) );
  XNOR U12464 ( .A(n11798), .B(n11797), .Z(n11800) );
  OR U12465 ( .A(n11799), .B(n11800), .Z(n11802) );
  XNOR U12466 ( .A(n11800), .B(n11799), .Z(n12191) );
  NAND U12467 ( .A(a[20]), .B(b[26]), .Z(n12190) );
  OR U12468 ( .A(n12191), .B(n12190), .Z(n11801) );
  NAND U12469 ( .A(n11802), .B(n11801), .Z(n11805) );
  ANDN U12470 ( .B(b[26]), .A(n21681), .Z(n11806) );
  OR U12471 ( .A(n11805), .B(n11806), .Z(n11808) );
  XOR U12472 ( .A(n11804), .B(n11803), .Z(n12197) );
  XOR U12473 ( .A(n11806), .B(n11805), .Z(n12196) );
  NANDN U12474 ( .A(n12197), .B(n12196), .Z(n11807) );
  NAND U12475 ( .A(n11808), .B(n11807), .Z(n11811) );
  XNOR U12476 ( .A(n11810), .B(n11809), .Z(n11812) );
  OR U12477 ( .A(n11811), .B(n11812), .Z(n11814) );
  XNOR U12478 ( .A(n11812), .B(n11811), .Z(n12203) );
  NAND U12479 ( .A(a[22]), .B(b[26]), .Z(n12202) );
  OR U12480 ( .A(n12203), .B(n12202), .Z(n11813) );
  NAND U12481 ( .A(n11814), .B(n11813), .Z(n11817) );
  ANDN U12482 ( .B(b[26]), .A(n21692), .Z(n11818) );
  OR U12483 ( .A(n11817), .B(n11818), .Z(n11820) );
  XOR U12484 ( .A(n11816), .B(n11815), .Z(n12209) );
  XOR U12485 ( .A(n11818), .B(n11817), .Z(n12208) );
  NANDN U12486 ( .A(n12209), .B(n12208), .Z(n11819) );
  NAND U12487 ( .A(n11820), .B(n11819), .Z(n11823) );
  XNOR U12488 ( .A(n11822), .B(n11821), .Z(n11824) );
  OR U12489 ( .A(n11823), .B(n11824), .Z(n11826) );
  XNOR U12490 ( .A(n11824), .B(n11823), .Z(n12215) );
  NAND U12491 ( .A(a[24]), .B(b[26]), .Z(n12214) );
  OR U12492 ( .A(n12215), .B(n12214), .Z(n11825) );
  NAND U12493 ( .A(n11826), .B(n11825), .Z(n11829) );
  ANDN U12494 ( .B(b[26]), .A(n21703), .Z(n11830) );
  OR U12495 ( .A(n11829), .B(n11830), .Z(n11832) );
  XOR U12496 ( .A(n11828), .B(n11827), .Z(n12221) );
  XOR U12497 ( .A(n11830), .B(n11829), .Z(n12220) );
  NANDN U12498 ( .A(n12221), .B(n12220), .Z(n11831) );
  NAND U12499 ( .A(n11832), .B(n11831), .Z(n11835) );
  XNOR U12500 ( .A(n11834), .B(n11833), .Z(n11836) );
  OR U12501 ( .A(n11835), .B(n11836), .Z(n11838) );
  XNOR U12502 ( .A(n11836), .B(n11835), .Z(n12227) );
  NAND U12503 ( .A(a[26]), .B(b[26]), .Z(n12226) );
  OR U12504 ( .A(n12227), .B(n12226), .Z(n11837) );
  NAND U12505 ( .A(n11838), .B(n11837), .Z(n11841) );
  ANDN U12506 ( .B(b[26]), .A(n21716), .Z(n11842) );
  OR U12507 ( .A(n11841), .B(n11842), .Z(n11844) );
  XOR U12508 ( .A(n11840), .B(n11839), .Z(n12233) );
  XOR U12509 ( .A(n11842), .B(n11841), .Z(n12232) );
  NANDN U12510 ( .A(n12233), .B(n12232), .Z(n11843) );
  NAND U12511 ( .A(n11844), .B(n11843), .Z(n11847) );
  XNOR U12512 ( .A(n11846), .B(n11845), .Z(n11848) );
  OR U12513 ( .A(n11847), .B(n11848), .Z(n11850) );
  XNOR U12514 ( .A(n11848), .B(n11847), .Z(n12239) );
  NAND U12515 ( .A(a[28]), .B(b[26]), .Z(n12238) );
  OR U12516 ( .A(n12239), .B(n12238), .Z(n11849) );
  NAND U12517 ( .A(n11850), .B(n11849), .Z(n11853) );
  ANDN U12518 ( .B(b[26]), .A(n21727), .Z(n11854) );
  OR U12519 ( .A(n11853), .B(n11854), .Z(n11856) );
  XOR U12520 ( .A(n11852), .B(n11851), .Z(n12245) );
  XOR U12521 ( .A(n11854), .B(n11853), .Z(n12244) );
  NANDN U12522 ( .A(n12245), .B(n12244), .Z(n11855) );
  NAND U12523 ( .A(n11856), .B(n11855), .Z(n11859) );
  XNOR U12524 ( .A(n11858), .B(n11857), .Z(n11860) );
  OR U12525 ( .A(n11859), .B(n11860), .Z(n11862) );
  XNOR U12526 ( .A(n11860), .B(n11859), .Z(n12251) );
  NAND U12527 ( .A(a[30]), .B(b[26]), .Z(n12250) );
  OR U12528 ( .A(n12251), .B(n12250), .Z(n11861) );
  NAND U12529 ( .A(n11862), .B(n11861), .Z(n11865) );
  ANDN U12530 ( .B(b[26]), .A(n21740), .Z(n11866) );
  OR U12531 ( .A(n11865), .B(n11866), .Z(n11868) );
  XOR U12532 ( .A(n11866), .B(n11865), .Z(n12256) );
  NANDN U12533 ( .A(n12257), .B(n12256), .Z(n11867) );
  NAND U12534 ( .A(n11868), .B(n11867), .Z(n11871) );
  XNOR U12535 ( .A(n11870), .B(n11869), .Z(n11872) );
  OR U12536 ( .A(n11871), .B(n11872), .Z(n11874) );
  XNOR U12537 ( .A(n11872), .B(n11871), .Z(n12263) );
  NAND U12538 ( .A(a[32]), .B(b[26]), .Z(n12262) );
  OR U12539 ( .A(n12263), .B(n12262), .Z(n11873) );
  NAND U12540 ( .A(n11874), .B(n11873), .Z(n11875) );
  ANDN U12541 ( .B(b[26]), .A(n21751), .Z(n11876) );
  OR U12542 ( .A(n11875), .B(n11876), .Z(n11880) );
  XNOR U12543 ( .A(n11876), .B(n11875), .Z(n12269) );
  XNOR U12544 ( .A(n11878), .B(n11877), .Z(n12268) );
  OR U12545 ( .A(n12269), .B(n12268), .Z(n11879) );
  AND U12546 ( .A(n11880), .B(n11879), .Z(n11883) );
  OR U12547 ( .A(n11883), .B(n11884), .Z(n11886) );
  ANDN U12548 ( .B(b[26]), .A(n183), .Z(n12277) );
  XOR U12549 ( .A(n11884), .B(n11883), .Z(n12276) );
  NANDN U12550 ( .A(n12277), .B(n12276), .Z(n11885) );
  NAND U12551 ( .A(n11886), .B(n11885), .Z(n11887) );
  OR U12552 ( .A(n11888), .B(n11887), .Z(n11892) );
  XNOR U12553 ( .A(n11888), .B(n11887), .Z(n12281) );
  XNOR U12554 ( .A(n11890), .B(n11889), .Z(n12280) );
  NANDN U12555 ( .A(n12281), .B(n12280), .Z(n11891) );
  AND U12556 ( .A(n11892), .B(n11891), .Z(n11895) );
  XNOR U12557 ( .A(n11894), .B(n11893), .Z(n11896) );
  OR U12558 ( .A(n11895), .B(n11896), .Z(n11898) );
  XNOR U12559 ( .A(n11896), .B(n11895), .Z(n12289) );
  AND U12560 ( .A(b[26]), .B(a[36]), .Z(n12288) );
  NANDN U12561 ( .A(n12289), .B(n12288), .Z(n11897) );
  NAND U12562 ( .A(n11898), .B(n11897), .Z(n11901) );
  ANDN U12563 ( .B(b[26]), .A(n21772), .Z(n11902) );
  OR U12564 ( .A(n11901), .B(n11902), .Z(n11904) );
  XOR U12565 ( .A(n11900), .B(n11899), .Z(n12293) );
  XOR U12566 ( .A(n11902), .B(n11901), .Z(n12292) );
  NANDN U12567 ( .A(n12293), .B(n12292), .Z(n11903) );
  NAND U12568 ( .A(n11904), .B(n11903), .Z(n11908) );
  AND U12569 ( .A(b[26]), .B(a[38]), .Z(n11907) );
  NANDN U12570 ( .A(n11908), .B(n11907), .Z(n11910) );
  XNOR U12571 ( .A(n11908), .B(n11907), .Z(n12300) );
  NANDN U12572 ( .A(n12301), .B(n12300), .Z(n11909) );
  NAND U12573 ( .A(n11910), .B(n11909), .Z(n11914) );
  NAND U12574 ( .A(n11914), .B(n11913), .Z(n11916) );
  XNOR U12575 ( .A(n11914), .B(n11913), .Z(n12305) );
  NAND U12576 ( .A(a[39]), .B(b[26]), .Z(n12304) );
  OR U12577 ( .A(n12305), .B(n12304), .Z(n11915) );
  NAND U12578 ( .A(n11916), .B(n11915), .Z(n11917) );
  NANDN U12579 ( .A(n11918), .B(n11917), .Z(n11922) );
  XOR U12580 ( .A(n11920), .B(n11919), .Z(n12311) );
  NAND U12581 ( .A(n12310), .B(n12311), .Z(n11921) );
  NAND U12582 ( .A(n11922), .B(n11921), .Z(n11925) );
  OR U12583 ( .A(n11926), .B(n11925), .Z(n11928) );
  XNOR U12584 ( .A(n11924), .B(n11923), .Z(n12317) );
  XOR U12585 ( .A(n11926), .B(n11925), .Z(n12316) );
  NANDN U12586 ( .A(n12317), .B(n12316), .Z(n11927) );
  NAND U12587 ( .A(n11928), .B(n11927), .Z(n11930) );
  NAND U12588 ( .A(a[42]), .B(b[26]), .Z(n11929) );
  OR U12589 ( .A(n11930), .B(n11929), .Z(n11934) );
  XOR U12590 ( .A(n11930), .B(n11929), .Z(n12322) );
  XOR U12591 ( .A(n11932), .B(n11931), .Z(n12323) );
  NAND U12592 ( .A(n12322), .B(n12323), .Z(n11933) );
  NAND U12593 ( .A(n11934), .B(n11933), .Z(n11937) );
  OR U12594 ( .A(n11938), .B(n11937), .Z(n11940) );
  XNOR U12595 ( .A(n11936), .B(n11935), .Z(n12329) );
  XOR U12596 ( .A(n11938), .B(n11937), .Z(n12328) );
  NANDN U12597 ( .A(n12329), .B(n12328), .Z(n11939) );
  NAND U12598 ( .A(n11940), .B(n11939), .Z(n11942) );
  NAND U12599 ( .A(a[44]), .B(b[26]), .Z(n11941) );
  OR U12600 ( .A(n11942), .B(n11941), .Z(n11946) );
  XOR U12601 ( .A(n11942), .B(n11941), .Z(n12334) );
  XOR U12602 ( .A(n11944), .B(n11943), .Z(n12335) );
  NAND U12603 ( .A(n12334), .B(n12335), .Z(n11945) );
  NAND U12604 ( .A(n11946), .B(n11945), .Z(n11949) );
  OR U12605 ( .A(n11950), .B(n11949), .Z(n11952) );
  XNOR U12606 ( .A(n11948), .B(n11947), .Z(n12341) );
  XOR U12607 ( .A(n11950), .B(n11949), .Z(n12340) );
  NANDN U12608 ( .A(n12341), .B(n12340), .Z(n11951) );
  NAND U12609 ( .A(n11952), .B(n11951), .Z(n11954) );
  NAND U12610 ( .A(a[46]), .B(b[26]), .Z(n11953) );
  OR U12611 ( .A(n11954), .B(n11953), .Z(n11958) );
  XOR U12612 ( .A(n11954), .B(n11953), .Z(n12346) );
  XOR U12613 ( .A(n11956), .B(n11955), .Z(n12347) );
  NAND U12614 ( .A(n12346), .B(n12347), .Z(n11957) );
  NAND U12615 ( .A(n11958), .B(n11957), .Z(n11961) );
  OR U12616 ( .A(n11962), .B(n11961), .Z(n11964) );
  XNOR U12617 ( .A(n11960), .B(n11959), .Z(n12353) );
  XOR U12618 ( .A(n11962), .B(n11961), .Z(n12352) );
  NANDN U12619 ( .A(n12353), .B(n12352), .Z(n11963) );
  NAND U12620 ( .A(n11964), .B(n11963), .Z(n11966) );
  NAND U12621 ( .A(a[48]), .B(b[26]), .Z(n11965) );
  OR U12622 ( .A(n11966), .B(n11965), .Z(n11970) );
  XOR U12623 ( .A(n11966), .B(n11965), .Z(n12358) );
  XOR U12624 ( .A(n11968), .B(n11967), .Z(n12359) );
  NAND U12625 ( .A(n12358), .B(n12359), .Z(n11969) );
  NAND U12626 ( .A(n11970), .B(n11969), .Z(n11973) );
  OR U12627 ( .A(n11974), .B(n11973), .Z(n11976) );
  XNOR U12628 ( .A(n11972), .B(n11971), .Z(n12365) );
  XOR U12629 ( .A(n11974), .B(n11973), .Z(n12364) );
  NANDN U12630 ( .A(n12365), .B(n12364), .Z(n11975) );
  NAND U12631 ( .A(n11976), .B(n11975), .Z(n11978) );
  NAND U12632 ( .A(a[50]), .B(b[26]), .Z(n11977) );
  OR U12633 ( .A(n11978), .B(n11977), .Z(n11982) );
  XOR U12634 ( .A(n11978), .B(n11977), .Z(n12370) );
  XOR U12635 ( .A(n11980), .B(n11979), .Z(n12371) );
  NAND U12636 ( .A(n12370), .B(n12371), .Z(n11981) );
  NAND U12637 ( .A(n11982), .B(n11981), .Z(n11985) );
  OR U12638 ( .A(n11986), .B(n11985), .Z(n11988) );
  XNOR U12639 ( .A(n11984), .B(n11983), .Z(n12377) );
  XOR U12640 ( .A(n11986), .B(n11985), .Z(n12376) );
  NANDN U12641 ( .A(n12377), .B(n12376), .Z(n11987) );
  NAND U12642 ( .A(n11988), .B(n11987), .Z(n11990) );
  NAND U12643 ( .A(a[52]), .B(b[26]), .Z(n11989) );
  OR U12644 ( .A(n11990), .B(n11989), .Z(n11994) );
  XOR U12645 ( .A(n11990), .B(n11989), .Z(n12382) );
  XOR U12646 ( .A(n11992), .B(n11991), .Z(n12383) );
  NAND U12647 ( .A(n12382), .B(n12383), .Z(n11993) );
  NAND U12648 ( .A(n11994), .B(n11993), .Z(n11997) );
  OR U12649 ( .A(n11998), .B(n11997), .Z(n12000) );
  XNOR U12650 ( .A(n11996), .B(n11995), .Z(n12389) );
  XOR U12651 ( .A(n11998), .B(n11997), .Z(n12388) );
  NANDN U12652 ( .A(n12389), .B(n12388), .Z(n11999) );
  NAND U12653 ( .A(n12000), .B(n11999), .Z(n12002) );
  NAND U12654 ( .A(a[54]), .B(b[26]), .Z(n12001) );
  OR U12655 ( .A(n12002), .B(n12001), .Z(n12006) );
  XOR U12656 ( .A(n12002), .B(n12001), .Z(n12394) );
  XOR U12657 ( .A(n12004), .B(n12003), .Z(n12395) );
  NAND U12658 ( .A(n12394), .B(n12395), .Z(n12005) );
  NAND U12659 ( .A(n12006), .B(n12005), .Z(n12009) );
  OR U12660 ( .A(n12010), .B(n12009), .Z(n12012) );
  XNOR U12661 ( .A(n12008), .B(n12007), .Z(n12401) );
  XOR U12662 ( .A(n12010), .B(n12009), .Z(n12400) );
  NANDN U12663 ( .A(n12401), .B(n12400), .Z(n12011) );
  NAND U12664 ( .A(n12012), .B(n12011), .Z(n12014) );
  NAND U12665 ( .A(a[56]), .B(b[26]), .Z(n12013) );
  OR U12666 ( .A(n12014), .B(n12013), .Z(n12018) );
  XOR U12667 ( .A(n12014), .B(n12013), .Z(n12406) );
  XOR U12668 ( .A(n12016), .B(n12015), .Z(n12407) );
  NAND U12669 ( .A(n12406), .B(n12407), .Z(n12017) );
  NAND U12670 ( .A(n12018), .B(n12017), .Z(n12021) );
  OR U12671 ( .A(n12022), .B(n12021), .Z(n12024) );
  XNOR U12672 ( .A(n12020), .B(n12019), .Z(n12413) );
  XOR U12673 ( .A(n12022), .B(n12021), .Z(n12412) );
  NANDN U12674 ( .A(n12413), .B(n12412), .Z(n12023) );
  NAND U12675 ( .A(n12024), .B(n12023), .Z(n12026) );
  NAND U12676 ( .A(a[58]), .B(b[26]), .Z(n12025) );
  OR U12677 ( .A(n12026), .B(n12025), .Z(n12030) );
  XOR U12678 ( .A(n12026), .B(n12025), .Z(n12418) );
  XOR U12679 ( .A(n12028), .B(n12027), .Z(n12419) );
  NAND U12680 ( .A(n12418), .B(n12419), .Z(n12029) );
  NAND U12681 ( .A(n12030), .B(n12029), .Z(n12033) );
  OR U12682 ( .A(n12034), .B(n12033), .Z(n12036) );
  XNOR U12683 ( .A(n12032), .B(n12031), .Z(n12425) );
  XOR U12684 ( .A(n12034), .B(n12033), .Z(n12424) );
  NANDN U12685 ( .A(n12425), .B(n12424), .Z(n12035) );
  NAND U12686 ( .A(n12036), .B(n12035), .Z(n12038) );
  NAND U12687 ( .A(a[60]), .B(b[26]), .Z(n12037) );
  OR U12688 ( .A(n12038), .B(n12037), .Z(n12042) );
  XOR U12689 ( .A(n12038), .B(n12037), .Z(n12430) );
  XOR U12690 ( .A(n12040), .B(n12039), .Z(n12431) );
  NAND U12691 ( .A(n12430), .B(n12431), .Z(n12041) );
  AND U12692 ( .A(n12042), .B(n12041), .Z(n12043) );
  NANDN U12693 ( .A(n12044), .B(n12043), .Z(n12048) );
  XOR U12694 ( .A(n12046), .B(n12045), .Z(n12436) );
  NANDN U12695 ( .A(n12437), .B(n12436), .Z(n12047) );
  NAND U12696 ( .A(n12048), .B(n12047), .Z(n12052) );
  NAND U12697 ( .A(a[62]), .B(b[26]), .Z(n12051) );
  OR U12698 ( .A(n12052), .B(n12051), .Z(n12054) );
  XOR U12699 ( .A(n12052), .B(n12051), .Z(n12071) );
  NAND U12700 ( .A(n12072), .B(n12071), .Z(n12053) );
  NAND U12701 ( .A(n12054), .B(n12053), .Z(n12055) );
  OR U12702 ( .A(n12056), .B(n12055), .Z(n12060) );
  XNOR U12703 ( .A(n12056), .B(n12055), .Z(n12446) );
  XOR U12704 ( .A(n12058), .B(n12057), .Z(n12447) );
  NANDN U12705 ( .A(n12446), .B(n12447), .Z(n12059) );
  NAND U12706 ( .A(n12060), .B(n12059), .Z(n12448) );
  OR U12707 ( .A(n12449), .B(n12448), .Z(n24181) );
  IV U12708 ( .A(n24181), .Z(n21975) );
  ANDN U12709 ( .B(n21974), .A(n21975), .Z(n24187) );
  OR U12710 ( .A(n12062), .B(n12061), .Z(n24183) );
  IV U12711 ( .A(n24183), .Z(n21977) );
  XOR U12712 ( .A(n12064), .B(n12063), .Z(n21980) );
  OR U12713 ( .A(n12066), .B(n12065), .Z(n12070) );
  NANDN U12714 ( .A(n12068), .B(n12067), .Z(n12069) );
  AND U12715 ( .A(n12070), .B(n12069), .Z(n21981) );
  XNOR U12716 ( .A(n21980), .B(n21981), .Z(n24182) );
  NANDN U12717 ( .A(n21977), .B(n24182), .Z(n24190) );
  XNOR U12718 ( .A(n12072), .B(n12071), .Z(n12442) );
  NAND U12719 ( .A(a[62]), .B(b[25]), .Z(n12438) );
  NAND U12720 ( .A(a[60]), .B(b[25]), .Z(n12426) );
  NAND U12721 ( .A(a[58]), .B(b[25]), .Z(n12414) );
  NAND U12722 ( .A(a[56]), .B(b[25]), .Z(n12402) );
  NAND U12723 ( .A(a[54]), .B(b[25]), .Z(n12390) );
  NAND U12724 ( .A(a[52]), .B(b[25]), .Z(n12378) );
  NAND U12725 ( .A(a[50]), .B(b[25]), .Z(n12366) );
  NAND U12726 ( .A(a[48]), .B(b[25]), .Z(n12354) );
  NAND U12727 ( .A(a[46]), .B(b[25]), .Z(n12342) );
  NAND U12728 ( .A(a[44]), .B(b[25]), .Z(n12330) );
  NAND U12729 ( .A(a[42]), .B(b[25]), .Z(n12318) );
  NAND U12730 ( .A(a[37]), .B(b[25]), .Z(n12287) );
  NAND U12731 ( .A(a[17]), .B(b[25]), .Z(n12167) );
  ANDN U12732 ( .B(b[25]), .A(n172), .Z(n12154) );
  ANDN U12733 ( .B(b[25]), .A(n170), .Z(n12143) );
  ANDN U12734 ( .B(b[25]), .A(n21164), .Z(n12131) );
  ANDN U12735 ( .B(b[25]), .A(n21615), .Z(n12119) );
  ANDN U12736 ( .B(b[25]), .A(n166), .Z(n12106) );
  XNOR U12737 ( .A(n12074), .B(n12073), .Z(n12103) );
  ANDN U12738 ( .B(b[25]), .A(n164), .Z(n12099) );
  ANDN U12739 ( .B(b[25]), .A(n21580), .Z(n12084) );
  NAND U12740 ( .A(b[26]), .B(a[1]), .Z(n12077) );
  AND U12741 ( .A(b[25]), .B(a[0]), .Z(n12843) );
  NANDN U12742 ( .A(n12077), .B(n12843), .Z(n12076) );
  NAND U12743 ( .A(a[2]), .B(b[25]), .Z(n12075) );
  AND U12744 ( .A(n12076), .B(n12075), .Z(n12083) );
  NANDN U12745 ( .A(n12077), .B(a[0]), .Z(n12078) );
  XNOR U12746 ( .A(a[2]), .B(n12078), .Z(n12079) );
  NAND U12747 ( .A(b[25]), .B(n12079), .Z(n12466) );
  AND U12748 ( .A(a[1]), .B(b[26]), .Z(n12080) );
  XNOR U12749 ( .A(n12081), .B(n12080), .Z(n12465) );
  NANDN U12750 ( .A(n12466), .B(n12465), .Z(n12082) );
  NANDN U12751 ( .A(n12083), .B(n12082), .Z(n12085) );
  NANDN U12752 ( .A(n12084), .B(n12085), .Z(n12089) );
  XOR U12753 ( .A(n12085), .B(n12084), .Z(n12470) );
  NANDN U12754 ( .A(n12470), .B(n12469), .Z(n12088) );
  NAND U12755 ( .A(n12089), .B(n12088), .Z(n12093) );
  XOR U12756 ( .A(n12091), .B(n12090), .Z(n12092) );
  NANDN U12757 ( .A(n12093), .B(n12092), .Z(n12095) );
  NAND U12758 ( .A(a[4]), .B(b[25]), .Z(n12475) );
  NANDN U12759 ( .A(n12475), .B(n12476), .Z(n12094) );
  NAND U12760 ( .A(n12095), .B(n12094), .Z(n12098) );
  OR U12761 ( .A(n12099), .B(n12098), .Z(n12101) );
  XOR U12762 ( .A(n12097), .B(n12096), .Z(n12453) );
  XOR U12763 ( .A(n12099), .B(n12098), .Z(n12452) );
  NAND U12764 ( .A(n12453), .B(n12452), .Z(n12100) );
  NAND U12765 ( .A(n12101), .B(n12100), .Z(n12102) );
  NANDN U12766 ( .A(n12103), .B(n12102), .Z(n12105) );
  ANDN U12767 ( .B(b[25]), .A(n165), .Z(n12488) );
  NANDN U12768 ( .A(n12488), .B(n12487), .Z(n12104) );
  NAND U12769 ( .A(n12105), .B(n12104), .Z(n12107) );
  NANDN U12770 ( .A(n12106), .B(n12107), .Z(n12111) );
  XOR U12771 ( .A(n12107), .B(n12106), .Z(n12492) );
  XOR U12772 ( .A(n12109), .B(n12108), .Z(n12491) );
  OR U12773 ( .A(n12492), .B(n12491), .Z(n12110) );
  NAND U12774 ( .A(n12111), .B(n12110), .Z(n12115) );
  XNOR U12775 ( .A(n12113), .B(n12112), .Z(n12114) );
  NANDN U12776 ( .A(n12115), .B(n12114), .Z(n12117) );
  NAND U12777 ( .A(a[8]), .B(b[25]), .Z(n12499) );
  NANDN U12778 ( .A(n12499), .B(n12500), .Z(n12116) );
  NAND U12779 ( .A(n12117), .B(n12116), .Z(n12118) );
  OR U12780 ( .A(n12119), .B(n12118), .Z(n12123) );
  XNOR U12781 ( .A(n12119), .B(n12118), .Z(n12503) );
  XOR U12782 ( .A(n12121), .B(n12120), .Z(n12504) );
  NANDN U12783 ( .A(n12503), .B(n12504), .Z(n12122) );
  NAND U12784 ( .A(n12123), .B(n12122), .Z(n12126) );
  XOR U12785 ( .A(n12125), .B(n12124), .Z(n12127) );
  NANDN U12786 ( .A(n12126), .B(n12127), .Z(n12129) );
  NAND U12787 ( .A(a[10]), .B(b[25]), .Z(n12511) );
  XNOR U12788 ( .A(n12127), .B(n12126), .Z(n12512) );
  NANDN U12789 ( .A(n12511), .B(n12512), .Z(n12128) );
  NAND U12790 ( .A(n12129), .B(n12128), .Z(n12130) );
  OR U12791 ( .A(n12131), .B(n12130), .Z(n12135) );
  XOR U12792 ( .A(n12131), .B(n12130), .Z(n12515) );
  XOR U12793 ( .A(n12133), .B(n12132), .Z(n12516) );
  NAND U12794 ( .A(n12515), .B(n12516), .Z(n12134) );
  NAND U12795 ( .A(n12135), .B(n12134), .Z(n12139) );
  XNOR U12796 ( .A(n12137), .B(n12136), .Z(n12138) );
  NANDN U12797 ( .A(n12139), .B(n12138), .Z(n12141) );
  NAND U12798 ( .A(a[12]), .B(b[25]), .Z(n12523) );
  NANDN U12799 ( .A(n12523), .B(n12524), .Z(n12140) );
  NAND U12800 ( .A(n12141), .B(n12140), .Z(n12142) );
  OR U12801 ( .A(n12143), .B(n12142), .Z(n12147) );
  XNOR U12802 ( .A(n12143), .B(n12142), .Z(n12527) );
  XOR U12803 ( .A(n12145), .B(n12144), .Z(n12528) );
  NANDN U12804 ( .A(n12527), .B(n12528), .Z(n12146) );
  NAND U12805 ( .A(n12147), .B(n12146), .Z(n12151) );
  XOR U12806 ( .A(n12149), .B(n12148), .Z(n12150) );
  NAND U12807 ( .A(n12151), .B(n12150), .Z(n12153) );
  ANDN U12808 ( .B(b[25]), .A(n171), .Z(n12534) );
  XNOR U12809 ( .A(n12151), .B(n12150), .Z(n12533) );
  OR U12810 ( .A(n12534), .B(n12533), .Z(n12152) );
  AND U12811 ( .A(n12153), .B(n12152), .Z(n12155) );
  OR U12812 ( .A(n12154), .B(n12155), .Z(n12159) );
  XNOR U12813 ( .A(n12155), .B(n12154), .Z(n12540) );
  OR U12814 ( .A(n12540), .B(n12539), .Z(n12158) );
  AND U12815 ( .A(n12159), .B(n12158), .Z(n12162) );
  OR U12816 ( .A(n12162), .B(n12163), .Z(n12165) );
  ANDN U12817 ( .B(b[25]), .A(n173), .Z(n12548) );
  XOR U12818 ( .A(n12163), .B(n12162), .Z(n12547) );
  NANDN U12819 ( .A(n12548), .B(n12547), .Z(n12164) );
  NAND U12820 ( .A(n12165), .B(n12164), .Z(n12166) );
  OR U12821 ( .A(n12167), .B(n12166), .Z(n12171) );
  XNOR U12822 ( .A(n12167), .B(n12166), .Z(n12552) );
  XNOR U12823 ( .A(n12169), .B(n12168), .Z(n12551) );
  NANDN U12824 ( .A(n12552), .B(n12551), .Z(n12170) );
  AND U12825 ( .A(n12171), .B(n12170), .Z(n12174) );
  XNOR U12826 ( .A(n12173), .B(n12172), .Z(n12175) );
  OR U12827 ( .A(n12174), .B(n12175), .Z(n12177) );
  XNOR U12828 ( .A(n12175), .B(n12174), .Z(n12558) );
  NAND U12829 ( .A(a[18]), .B(b[25]), .Z(n12557) );
  OR U12830 ( .A(n12558), .B(n12557), .Z(n12176) );
  NAND U12831 ( .A(n12177), .B(n12176), .Z(n12180) );
  ANDN U12832 ( .B(b[25]), .A(n21670), .Z(n12181) );
  OR U12833 ( .A(n12180), .B(n12181), .Z(n12183) );
  XOR U12834 ( .A(n12179), .B(n12178), .Z(n12564) );
  XOR U12835 ( .A(n12181), .B(n12180), .Z(n12563) );
  NANDN U12836 ( .A(n12564), .B(n12563), .Z(n12182) );
  NAND U12837 ( .A(n12183), .B(n12182), .Z(n12186) );
  XNOR U12838 ( .A(n12185), .B(n12184), .Z(n12187) );
  OR U12839 ( .A(n12186), .B(n12187), .Z(n12189) );
  XNOR U12840 ( .A(n12187), .B(n12186), .Z(n12570) );
  NAND U12841 ( .A(a[20]), .B(b[25]), .Z(n12569) );
  OR U12842 ( .A(n12570), .B(n12569), .Z(n12188) );
  NAND U12843 ( .A(n12189), .B(n12188), .Z(n12192) );
  ANDN U12844 ( .B(b[25]), .A(n21681), .Z(n12193) );
  OR U12845 ( .A(n12192), .B(n12193), .Z(n12195) );
  XOR U12846 ( .A(n12191), .B(n12190), .Z(n12576) );
  XOR U12847 ( .A(n12193), .B(n12192), .Z(n12575) );
  NANDN U12848 ( .A(n12576), .B(n12575), .Z(n12194) );
  NAND U12849 ( .A(n12195), .B(n12194), .Z(n12198) );
  XNOR U12850 ( .A(n12197), .B(n12196), .Z(n12199) );
  OR U12851 ( .A(n12198), .B(n12199), .Z(n12201) );
  XNOR U12852 ( .A(n12199), .B(n12198), .Z(n12582) );
  NAND U12853 ( .A(a[22]), .B(b[25]), .Z(n12581) );
  OR U12854 ( .A(n12582), .B(n12581), .Z(n12200) );
  NAND U12855 ( .A(n12201), .B(n12200), .Z(n12204) );
  ANDN U12856 ( .B(b[25]), .A(n21692), .Z(n12205) );
  OR U12857 ( .A(n12204), .B(n12205), .Z(n12207) );
  XOR U12858 ( .A(n12203), .B(n12202), .Z(n12588) );
  XOR U12859 ( .A(n12205), .B(n12204), .Z(n12587) );
  NANDN U12860 ( .A(n12588), .B(n12587), .Z(n12206) );
  NAND U12861 ( .A(n12207), .B(n12206), .Z(n12210) );
  XNOR U12862 ( .A(n12209), .B(n12208), .Z(n12211) );
  OR U12863 ( .A(n12210), .B(n12211), .Z(n12213) );
  XNOR U12864 ( .A(n12211), .B(n12210), .Z(n12594) );
  NAND U12865 ( .A(a[24]), .B(b[25]), .Z(n12593) );
  OR U12866 ( .A(n12594), .B(n12593), .Z(n12212) );
  NAND U12867 ( .A(n12213), .B(n12212), .Z(n12216) );
  ANDN U12868 ( .B(b[25]), .A(n21703), .Z(n12217) );
  OR U12869 ( .A(n12216), .B(n12217), .Z(n12219) );
  XOR U12870 ( .A(n12215), .B(n12214), .Z(n12600) );
  XOR U12871 ( .A(n12217), .B(n12216), .Z(n12599) );
  NANDN U12872 ( .A(n12600), .B(n12599), .Z(n12218) );
  NAND U12873 ( .A(n12219), .B(n12218), .Z(n12222) );
  XNOR U12874 ( .A(n12221), .B(n12220), .Z(n12223) );
  OR U12875 ( .A(n12222), .B(n12223), .Z(n12225) );
  XNOR U12876 ( .A(n12223), .B(n12222), .Z(n12606) );
  NAND U12877 ( .A(a[26]), .B(b[25]), .Z(n12605) );
  OR U12878 ( .A(n12606), .B(n12605), .Z(n12224) );
  NAND U12879 ( .A(n12225), .B(n12224), .Z(n12228) );
  ANDN U12880 ( .B(b[25]), .A(n21716), .Z(n12229) );
  OR U12881 ( .A(n12228), .B(n12229), .Z(n12231) );
  XOR U12882 ( .A(n12227), .B(n12226), .Z(n12612) );
  XOR U12883 ( .A(n12229), .B(n12228), .Z(n12611) );
  NANDN U12884 ( .A(n12612), .B(n12611), .Z(n12230) );
  NAND U12885 ( .A(n12231), .B(n12230), .Z(n12234) );
  XNOR U12886 ( .A(n12233), .B(n12232), .Z(n12235) );
  OR U12887 ( .A(n12234), .B(n12235), .Z(n12237) );
  XNOR U12888 ( .A(n12235), .B(n12234), .Z(n12618) );
  NAND U12889 ( .A(a[28]), .B(b[25]), .Z(n12617) );
  OR U12890 ( .A(n12618), .B(n12617), .Z(n12236) );
  NAND U12891 ( .A(n12237), .B(n12236), .Z(n12240) );
  ANDN U12892 ( .B(b[25]), .A(n21727), .Z(n12241) );
  OR U12893 ( .A(n12240), .B(n12241), .Z(n12243) );
  XOR U12894 ( .A(n12239), .B(n12238), .Z(n12624) );
  XOR U12895 ( .A(n12241), .B(n12240), .Z(n12623) );
  NANDN U12896 ( .A(n12624), .B(n12623), .Z(n12242) );
  NAND U12897 ( .A(n12243), .B(n12242), .Z(n12246) );
  XNOR U12898 ( .A(n12245), .B(n12244), .Z(n12247) );
  OR U12899 ( .A(n12246), .B(n12247), .Z(n12249) );
  XNOR U12900 ( .A(n12247), .B(n12246), .Z(n12630) );
  NAND U12901 ( .A(a[30]), .B(b[25]), .Z(n12629) );
  OR U12902 ( .A(n12630), .B(n12629), .Z(n12248) );
  NAND U12903 ( .A(n12249), .B(n12248), .Z(n12252) );
  ANDN U12904 ( .B(b[25]), .A(n21740), .Z(n12253) );
  OR U12905 ( .A(n12252), .B(n12253), .Z(n12255) );
  XOR U12906 ( .A(n12251), .B(n12250), .Z(n12636) );
  XOR U12907 ( .A(n12253), .B(n12252), .Z(n12635) );
  NANDN U12908 ( .A(n12636), .B(n12635), .Z(n12254) );
  NAND U12909 ( .A(n12255), .B(n12254), .Z(n12258) );
  XNOR U12910 ( .A(n12257), .B(n12256), .Z(n12259) );
  OR U12911 ( .A(n12258), .B(n12259), .Z(n12261) );
  XNOR U12912 ( .A(n12259), .B(n12258), .Z(n12642) );
  NAND U12913 ( .A(a[32]), .B(b[25]), .Z(n12641) );
  OR U12914 ( .A(n12642), .B(n12641), .Z(n12260) );
  NAND U12915 ( .A(n12261), .B(n12260), .Z(n12264) );
  ANDN U12916 ( .B(b[25]), .A(n21751), .Z(n12265) );
  OR U12917 ( .A(n12264), .B(n12265), .Z(n12267) );
  XOR U12918 ( .A(n12263), .B(n12262), .Z(n12648) );
  XOR U12919 ( .A(n12265), .B(n12264), .Z(n12647) );
  NANDN U12920 ( .A(n12648), .B(n12647), .Z(n12266) );
  NAND U12921 ( .A(n12267), .B(n12266), .Z(n12270) );
  XOR U12922 ( .A(n12269), .B(n12268), .Z(n12271) );
  OR U12923 ( .A(n12270), .B(n12271), .Z(n12273) );
  NAND U12924 ( .A(a[34]), .B(b[25]), .Z(n12654) );
  XOR U12925 ( .A(n12271), .B(n12270), .Z(n12653) );
  NANDN U12926 ( .A(n12654), .B(n12653), .Z(n12272) );
  NAND U12927 ( .A(n12273), .B(n12272), .Z(n12274) );
  ANDN U12928 ( .B(b[25]), .A(n184), .Z(n12275) );
  OR U12929 ( .A(n12274), .B(n12275), .Z(n12279) );
  XNOR U12930 ( .A(n12275), .B(n12274), .Z(n12660) );
  XOR U12931 ( .A(n12277), .B(n12276), .Z(n12659) );
  OR U12932 ( .A(n12660), .B(n12659), .Z(n12278) );
  AND U12933 ( .A(n12279), .B(n12278), .Z(n12282) );
  OR U12934 ( .A(n12282), .B(n12283), .Z(n12285) );
  ANDN U12935 ( .B(b[25]), .A(n185), .Z(n12668) );
  XOR U12936 ( .A(n12283), .B(n12282), .Z(n12667) );
  NANDN U12937 ( .A(n12668), .B(n12667), .Z(n12284) );
  NAND U12938 ( .A(n12285), .B(n12284), .Z(n12286) );
  OR U12939 ( .A(n12287), .B(n12286), .Z(n12291) );
  XNOR U12940 ( .A(n12287), .B(n12286), .Z(n12672) );
  XNOR U12941 ( .A(n12289), .B(n12288), .Z(n12671) );
  NANDN U12942 ( .A(n12672), .B(n12671), .Z(n12290) );
  AND U12943 ( .A(n12291), .B(n12290), .Z(n12294) );
  XNOR U12944 ( .A(n12293), .B(n12292), .Z(n12295) );
  OR U12945 ( .A(n12294), .B(n12295), .Z(n12297) );
  XNOR U12946 ( .A(n12295), .B(n12294), .Z(n12678) );
  NAND U12947 ( .A(a[38]), .B(b[25]), .Z(n12677) );
  OR U12948 ( .A(n12678), .B(n12677), .Z(n12296) );
  NAND U12949 ( .A(n12297), .B(n12296), .Z(n12298) );
  ANDN U12950 ( .B(b[25]), .A(n187), .Z(n12299) );
  OR U12951 ( .A(n12298), .B(n12299), .Z(n12303) );
  XOR U12952 ( .A(n12299), .B(n12298), .Z(n12683) );
  NAND U12953 ( .A(n12683), .B(n12684), .Z(n12302) );
  NAND U12954 ( .A(n12303), .B(n12302), .Z(n12307) );
  NAND U12955 ( .A(a[40]), .B(b[25]), .Z(n12306) );
  OR U12956 ( .A(n12307), .B(n12306), .Z(n12309) );
  XOR U12957 ( .A(n12305), .B(n12304), .Z(n12689) );
  XOR U12958 ( .A(n12307), .B(n12306), .Z(n12690) );
  NAND U12959 ( .A(n12689), .B(n12690), .Z(n12308) );
  NAND U12960 ( .A(n12309), .B(n12308), .Z(n12313) );
  NAND U12961 ( .A(n12313), .B(n12312), .Z(n12315) );
  XNOR U12962 ( .A(n12313), .B(n12312), .Z(n12696) );
  NAND U12963 ( .A(a[41]), .B(b[25]), .Z(n12695) );
  OR U12964 ( .A(n12696), .B(n12695), .Z(n12314) );
  NAND U12965 ( .A(n12315), .B(n12314), .Z(n12319) );
  NANDN U12966 ( .A(n12318), .B(n12319), .Z(n12321) );
  XNOR U12967 ( .A(n12317), .B(n12316), .Z(n12702) );
  XNOR U12968 ( .A(n12319), .B(n12318), .Z(n12701) );
  NANDN U12969 ( .A(n12702), .B(n12701), .Z(n12320) );
  NAND U12970 ( .A(n12321), .B(n12320), .Z(n12325) );
  NAND U12971 ( .A(n12325), .B(n12324), .Z(n12327) );
  XNOR U12972 ( .A(n12325), .B(n12324), .Z(n12708) );
  NAND U12973 ( .A(a[43]), .B(b[25]), .Z(n12707) );
  OR U12974 ( .A(n12708), .B(n12707), .Z(n12326) );
  NAND U12975 ( .A(n12327), .B(n12326), .Z(n12331) );
  NANDN U12976 ( .A(n12330), .B(n12331), .Z(n12333) );
  XNOR U12977 ( .A(n12329), .B(n12328), .Z(n12714) );
  XNOR U12978 ( .A(n12331), .B(n12330), .Z(n12713) );
  NANDN U12979 ( .A(n12714), .B(n12713), .Z(n12332) );
  NAND U12980 ( .A(n12333), .B(n12332), .Z(n12337) );
  NAND U12981 ( .A(n12337), .B(n12336), .Z(n12339) );
  XNOR U12982 ( .A(n12337), .B(n12336), .Z(n12720) );
  NAND U12983 ( .A(a[45]), .B(b[25]), .Z(n12719) );
  OR U12984 ( .A(n12720), .B(n12719), .Z(n12338) );
  NAND U12985 ( .A(n12339), .B(n12338), .Z(n12343) );
  NANDN U12986 ( .A(n12342), .B(n12343), .Z(n12345) );
  XNOR U12987 ( .A(n12341), .B(n12340), .Z(n12726) );
  XNOR U12988 ( .A(n12343), .B(n12342), .Z(n12725) );
  NANDN U12989 ( .A(n12726), .B(n12725), .Z(n12344) );
  NAND U12990 ( .A(n12345), .B(n12344), .Z(n12349) );
  NAND U12991 ( .A(n12349), .B(n12348), .Z(n12351) );
  XNOR U12992 ( .A(n12349), .B(n12348), .Z(n12732) );
  NAND U12993 ( .A(a[47]), .B(b[25]), .Z(n12731) );
  OR U12994 ( .A(n12732), .B(n12731), .Z(n12350) );
  NAND U12995 ( .A(n12351), .B(n12350), .Z(n12355) );
  NANDN U12996 ( .A(n12354), .B(n12355), .Z(n12357) );
  XNOR U12997 ( .A(n12353), .B(n12352), .Z(n12738) );
  XNOR U12998 ( .A(n12355), .B(n12354), .Z(n12737) );
  NANDN U12999 ( .A(n12738), .B(n12737), .Z(n12356) );
  NAND U13000 ( .A(n12357), .B(n12356), .Z(n12361) );
  NAND U13001 ( .A(n12361), .B(n12360), .Z(n12363) );
  XNOR U13002 ( .A(n12361), .B(n12360), .Z(n12744) );
  NAND U13003 ( .A(a[49]), .B(b[25]), .Z(n12743) );
  OR U13004 ( .A(n12744), .B(n12743), .Z(n12362) );
  NAND U13005 ( .A(n12363), .B(n12362), .Z(n12367) );
  NANDN U13006 ( .A(n12366), .B(n12367), .Z(n12369) );
  XNOR U13007 ( .A(n12365), .B(n12364), .Z(n12750) );
  XNOR U13008 ( .A(n12367), .B(n12366), .Z(n12749) );
  NANDN U13009 ( .A(n12750), .B(n12749), .Z(n12368) );
  NAND U13010 ( .A(n12369), .B(n12368), .Z(n12373) );
  NAND U13011 ( .A(n12373), .B(n12372), .Z(n12375) );
  XNOR U13012 ( .A(n12373), .B(n12372), .Z(n12756) );
  NAND U13013 ( .A(a[51]), .B(b[25]), .Z(n12755) );
  OR U13014 ( .A(n12756), .B(n12755), .Z(n12374) );
  NAND U13015 ( .A(n12375), .B(n12374), .Z(n12379) );
  NANDN U13016 ( .A(n12378), .B(n12379), .Z(n12381) );
  XNOR U13017 ( .A(n12377), .B(n12376), .Z(n12762) );
  XNOR U13018 ( .A(n12379), .B(n12378), .Z(n12761) );
  NANDN U13019 ( .A(n12762), .B(n12761), .Z(n12380) );
  NAND U13020 ( .A(n12381), .B(n12380), .Z(n12385) );
  NAND U13021 ( .A(n12385), .B(n12384), .Z(n12387) );
  XNOR U13022 ( .A(n12385), .B(n12384), .Z(n12768) );
  NAND U13023 ( .A(a[53]), .B(b[25]), .Z(n12767) );
  OR U13024 ( .A(n12768), .B(n12767), .Z(n12386) );
  NAND U13025 ( .A(n12387), .B(n12386), .Z(n12391) );
  NANDN U13026 ( .A(n12390), .B(n12391), .Z(n12393) );
  XNOR U13027 ( .A(n12389), .B(n12388), .Z(n12774) );
  XNOR U13028 ( .A(n12391), .B(n12390), .Z(n12773) );
  NANDN U13029 ( .A(n12774), .B(n12773), .Z(n12392) );
  NAND U13030 ( .A(n12393), .B(n12392), .Z(n12397) );
  NAND U13031 ( .A(n12397), .B(n12396), .Z(n12399) );
  XNOR U13032 ( .A(n12397), .B(n12396), .Z(n12780) );
  NAND U13033 ( .A(a[55]), .B(b[25]), .Z(n12779) );
  OR U13034 ( .A(n12780), .B(n12779), .Z(n12398) );
  NAND U13035 ( .A(n12399), .B(n12398), .Z(n12403) );
  NANDN U13036 ( .A(n12402), .B(n12403), .Z(n12405) );
  XNOR U13037 ( .A(n12401), .B(n12400), .Z(n12786) );
  XNOR U13038 ( .A(n12403), .B(n12402), .Z(n12785) );
  NANDN U13039 ( .A(n12786), .B(n12785), .Z(n12404) );
  NAND U13040 ( .A(n12405), .B(n12404), .Z(n12409) );
  NAND U13041 ( .A(n12409), .B(n12408), .Z(n12411) );
  XNOR U13042 ( .A(n12409), .B(n12408), .Z(n12792) );
  NAND U13043 ( .A(a[57]), .B(b[25]), .Z(n12791) );
  OR U13044 ( .A(n12792), .B(n12791), .Z(n12410) );
  NAND U13045 ( .A(n12411), .B(n12410), .Z(n12415) );
  NANDN U13046 ( .A(n12414), .B(n12415), .Z(n12417) );
  XNOR U13047 ( .A(n12413), .B(n12412), .Z(n12798) );
  XNOR U13048 ( .A(n12415), .B(n12414), .Z(n12797) );
  NANDN U13049 ( .A(n12798), .B(n12797), .Z(n12416) );
  NAND U13050 ( .A(n12417), .B(n12416), .Z(n12421) );
  NAND U13051 ( .A(n12421), .B(n12420), .Z(n12423) );
  XNOR U13052 ( .A(n12421), .B(n12420), .Z(n12804) );
  NAND U13053 ( .A(a[59]), .B(b[25]), .Z(n12803) );
  OR U13054 ( .A(n12804), .B(n12803), .Z(n12422) );
  NAND U13055 ( .A(n12423), .B(n12422), .Z(n12427) );
  NANDN U13056 ( .A(n12426), .B(n12427), .Z(n12429) );
  XNOR U13057 ( .A(n12425), .B(n12424), .Z(n12810) );
  XNOR U13058 ( .A(n12427), .B(n12426), .Z(n12809) );
  NANDN U13059 ( .A(n12810), .B(n12809), .Z(n12428) );
  NAND U13060 ( .A(n12429), .B(n12428), .Z(n12433) );
  NAND U13061 ( .A(n12433), .B(n12432), .Z(n12435) );
  XNOR U13062 ( .A(n12433), .B(n12432), .Z(n12816) );
  NAND U13063 ( .A(a[61]), .B(b[25]), .Z(n12815) );
  OR U13064 ( .A(n12816), .B(n12815), .Z(n12434) );
  NAND U13065 ( .A(n12435), .B(n12434), .Z(n12439) );
  NANDN U13066 ( .A(n12438), .B(n12439), .Z(n12441) );
  XNOR U13067 ( .A(n12439), .B(n12438), .Z(n12821) );
  NAND U13068 ( .A(n12822), .B(n12821), .Z(n12440) );
  AND U13069 ( .A(n12441), .B(n12440), .Z(n12443) );
  OR U13070 ( .A(n12442), .B(n12443), .Z(n12445) );
  XNOR U13071 ( .A(n12443), .B(n12442), .Z(n12451) );
  AND U13072 ( .A(b[25]), .B(a[63]), .Z(n12450) );
  NANDN U13073 ( .A(n12451), .B(n12450), .Z(n12444) );
  AND U13074 ( .A(n12445), .B(n12444), .Z(n12827) );
  XOR U13075 ( .A(n12447), .B(n12446), .Z(n12828) );
  NANDN U13076 ( .A(n12827), .B(n12828), .Z(n24175) );
  XOR U13077 ( .A(n12449), .B(n12448), .Z(n24174) );
  IV U13078 ( .A(n24174), .Z(n21976) );
  XOR U13079 ( .A(n12451), .B(n12450), .Z(n12832) );
  NAND U13080 ( .A(a[42]), .B(b[24]), .Z(n12697) );
  ANDN U13081 ( .B(b[24]), .A(n187), .Z(n12679) );
  ANDN U13082 ( .B(b[24]), .A(n21670), .Z(n12559) );
  ANDN U13083 ( .B(b[24]), .A(n174), .Z(n12545) );
  ANDN U13084 ( .B(b[24]), .A(n172), .Z(n12536) );
  ANDN U13085 ( .B(b[24]), .A(n170), .Z(n12522) );
  ANDN U13086 ( .B(b[24]), .A(n21164), .Z(n12510) );
  ANDN U13087 ( .B(b[24]), .A(n21615), .Z(n12498) );
  ANDN U13088 ( .B(b[24]), .A(n166), .Z(n12485) );
  XNOR U13089 ( .A(n12453), .B(n12452), .Z(n12482) );
  ANDN U13090 ( .B(b[24]), .A(n164), .Z(n12478) );
  ANDN U13091 ( .B(b[24]), .A(n21580), .Z(n12463) );
  NAND U13092 ( .A(b[25]), .B(a[1]), .Z(n12456) );
  AND U13093 ( .A(b[24]), .B(a[0]), .Z(n13224) );
  NANDN U13094 ( .A(n12456), .B(n13224), .Z(n12455) );
  NAND U13095 ( .A(a[2]), .B(b[24]), .Z(n12454) );
  AND U13096 ( .A(n12455), .B(n12454), .Z(n12462) );
  NANDN U13097 ( .A(n12456), .B(a[0]), .Z(n12457) );
  XNOR U13098 ( .A(a[2]), .B(n12457), .Z(n12458) );
  NAND U13099 ( .A(b[24]), .B(n12458), .Z(n12849) );
  AND U13100 ( .A(a[1]), .B(b[25]), .Z(n12459) );
  XNOR U13101 ( .A(n12460), .B(n12459), .Z(n12848) );
  NANDN U13102 ( .A(n12849), .B(n12848), .Z(n12461) );
  NANDN U13103 ( .A(n12462), .B(n12461), .Z(n12464) );
  NANDN U13104 ( .A(n12463), .B(n12464), .Z(n12468) );
  XOR U13105 ( .A(n12464), .B(n12463), .Z(n12853) );
  NANDN U13106 ( .A(n12853), .B(n12852), .Z(n12467) );
  NAND U13107 ( .A(n12468), .B(n12467), .Z(n12472) );
  XOR U13108 ( .A(n12470), .B(n12469), .Z(n12471) );
  NANDN U13109 ( .A(n12472), .B(n12471), .Z(n12474) );
  NAND U13110 ( .A(a[4]), .B(b[24]), .Z(n12858) );
  NANDN U13111 ( .A(n12858), .B(n12859), .Z(n12473) );
  NAND U13112 ( .A(n12474), .B(n12473), .Z(n12477) );
  OR U13113 ( .A(n12478), .B(n12477), .Z(n12480) );
  XOR U13114 ( .A(n12476), .B(n12475), .Z(n12836) );
  XOR U13115 ( .A(n12478), .B(n12477), .Z(n12835) );
  NAND U13116 ( .A(n12836), .B(n12835), .Z(n12479) );
  NAND U13117 ( .A(n12480), .B(n12479), .Z(n12481) );
  NANDN U13118 ( .A(n12482), .B(n12481), .Z(n12484) );
  ANDN U13119 ( .B(b[24]), .A(n165), .Z(n12871) );
  NANDN U13120 ( .A(n12871), .B(n12870), .Z(n12483) );
  NAND U13121 ( .A(n12484), .B(n12483), .Z(n12486) );
  NANDN U13122 ( .A(n12485), .B(n12486), .Z(n12490) );
  XOR U13123 ( .A(n12486), .B(n12485), .Z(n12875) );
  XOR U13124 ( .A(n12488), .B(n12487), .Z(n12874) );
  OR U13125 ( .A(n12875), .B(n12874), .Z(n12489) );
  NAND U13126 ( .A(n12490), .B(n12489), .Z(n12494) );
  XNOR U13127 ( .A(n12492), .B(n12491), .Z(n12493) );
  NANDN U13128 ( .A(n12494), .B(n12493), .Z(n12496) );
  NAND U13129 ( .A(a[8]), .B(b[24]), .Z(n12882) );
  NANDN U13130 ( .A(n12882), .B(n12883), .Z(n12495) );
  NAND U13131 ( .A(n12496), .B(n12495), .Z(n12497) );
  OR U13132 ( .A(n12498), .B(n12497), .Z(n12502) );
  XNOR U13133 ( .A(n12498), .B(n12497), .Z(n12886) );
  XOR U13134 ( .A(n12500), .B(n12499), .Z(n12887) );
  NANDN U13135 ( .A(n12886), .B(n12887), .Z(n12501) );
  NAND U13136 ( .A(n12502), .B(n12501), .Z(n12505) );
  XOR U13137 ( .A(n12504), .B(n12503), .Z(n12506) );
  NANDN U13138 ( .A(n12505), .B(n12506), .Z(n12508) );
  NAND U13139 ( .A(a[10]), .B(b[24]), .Z(n12894) );
  XNOR U13140 ( .A(n12506), .B(n12505), .Z(n12895) );
  NANDN U13141 ( .A(n12894), .B(n12895), .Z(n12507) );
  NAND U13142 ( .A(n12508), .B(n12507), .Z(n12509) );
  OR U13143 ( .A(n12510), .B(n12509), .Z(n12514) );
  XNOR U13144 ( .A(n12510), .B(n12509), .Z(n12898) );
  XOR U13145 ( .A(n12512), .B(n12511), .Z(n12899) );
  NANDN U13146 ( .A(n12898), .B(n12899), .Z(n12513) );
  NAND U13147 ( .A(n12514), .B(n12513), .Z(n12518) );
  NAND U13148 ( .A(n12518), .B(n12517), .Z(n12520) );
  ANDN U13149 ( .B(b[24]), .A(n169), .Z(n12905) );
  XNOR U13150 ( .A(n12518), .B(n12517), .Z(n12904) );
  OR U13151 ( .A(n12905), .B(n12904), .Z(n12519) );
  NAND U13152 ( .A(n12520), .B(n12519), .Z(n12521) );
  NANDN U13153 ( .A(n12522), .B(n12521), .Z(n12526) );
  XOR U13154 ( .A(n12524), .B(n12523), .Z(n12910) );
  NANDN U13155 ( .A(n12911), .B(n12910), .Z(n12525) );
  NAND U13156 ( .A(n12526), .B(n12525), .Z(n12529) );
  XOR U13157 ( .A(n12528), .B(n12527), .Z(n12530) );
  NANDN U13158 ( .A(n12529), .B(n12530), .Z(n12532) );
  NAND U13159 ( .A(a[14]), .B(b[24]), .Z(n12918) );
  XNOR U13160 ( .A(n12530), .B(n12529), .Z(n12919) );
  NANDN U13161 ( .A(n12918), .B(n12919), .Z(n12531) );
  NAND U13162 ( .A(n12532), .B(n12531), .Z(n12535) );
  OR U13163 ( .A(n12536), .B(n12535), .Z(n12538) );
  XOR U13164 ( .A(n12534), .B(n12533), .Z(n12833) );
  XOR U13165 ( .A(n12536), .B(n12535), .Z(n12834) );
  NAND U13166 ( .A(n12833), .B(n12834), .Z(n12537) );
  NAND U13167 ( .A(n12538), .B(n12537), .Z(n12542) );
  XOR U13168 ( .A(n12540), .B(n12539), .Z(n12541) );
  NAND U13169 ( .A(n12542), .B(n12541), .Z(n12544) );
  ANDN U13170 ( .B(b[24]), .A(n173), .Z(n12927) );
  XNOR U13171 ( .A(n12542), .B(n12541), .Z(n12926) );
  OR U13172 ( .A(n12927), .B(n12926), .Z(n12543) );
  AND U13173 ( .A(n12544), .B(n12543), .Z(n12546) );
  OR U13174 ( .A(n12545), .B(n12546), .Z(n12550) );
  XNOR U13175 ( .A(n12546), .B(n12545), .Z(n12933) );
  OR U13176 ( .A(n12933), .B(n12932), .Z(n12549) );
  AND U13177 ( .A(n12550), .B(n12549), .Z(n12553) );
  OR U13178 ( .A(n12553), .B(n12554), .Z(n12556) );
  ANDN U13179 ( .B(b[24]), .A(n175), .Z(n12941) );
  XOR U13180 ( .A(n12554), .B(n12553), .Z(n12940) );
  NANDN U13181 ( .A(n12941), .B(n12940), .Z(n12555) );
  AND U13182 ( .A(n12556), .B(n12555), .Z(n12560) );
  OR U13183 ( .A(n12559), .B(n12560), .Z(n12562) );
  XOR U13184 ( .A(n12558), .B(n12557), .Z(n12945) );
  XOR U13185 ( .A(n12560), .B(n12559), .Z(n12944) );
  NANDN U13186 ( .A(n12945), .B(n12944), .Z(n12561) );
  NAND U13187 ( .A(n12562), .B(n12561), .Z(n12565) );
  XNOR U13188 ( .A(n12564), .B(n12563), .Z(n12566) );
  OR U13189 ( .A(n12565), .B(n12566), .Z(n12568) );
  XNOR U13190 ( .A(n12566), .B(n12565), .Z(n12951) );
  NAND U13191 ( .A(a[20]), .B(b[24]), .Z(n12950) );
  OR U13192 ( .A(n12951), .B(n12950), .Z(n12567) );
  NAND U13193 ( .A(n12568), .B(n12567), .Z(n12571) );
  ANDN U13194 ( .B(b[24]), .A(n21681), .Z(n12572) );
  OR U13195 ( .A(n12571), .B(n12572), .Z(n12574) );
  XOR U13196 ( .A(n12570), .B(n12569), .Z(n12957) );
  XOR U13197 ( .A(n12572), .B(n12571), .Z(n12956) );
  NANDN U13198 ( .A(n12957), .B(n12956), .Z(n12573) );
  NAND U13199 ( .A(n12574), .B(n12573), .Z(n12577) );
  XNOR U13200 ( .A(n12576), .B(n12575), .Z(n12578) );
  OR U13201 ( .A(n12577), .B(n12578), .Z(n12580) );
  XNOR U13202 ( .A(n12578), .B(n12577), .Z(n12963) );
  NAND U13203 ( .A(a[22]), .B(b[24]), .Z(n12962) );
  OR U13204 ( .A(n12963), .B(n12962), .Z(n12579) );
  NAND U13205 ( .A(n12580), .B(n12579), .Z(n12583) );
  ANDN U13206 ( .B(b[24]), .A(n21692), .Z(n12584) );
  OR U13207 ( .A(n12583), .B(n12584), .Z(n12586) );
  XOR U13208 ( .A(n12582), .B(n12581), .Z(n12969) );
  XOR U13209 ( .A(n12584), .B(n12583), .Z(n12968) );
  NANDN U13210 ( .A(n12969), .B(n12968), .Z(n12585) );
  NAND U13211 ( .A(n12586), .B(n12585), .Z(n12589) );
  XNOR U13212 ( .A(n12588), .B(n12587), .Z(n12590) );
  OR U13213 ( .A(n12589), .B(n12590), .Z(n12592) );
  XNOR U13214 ( .A(n12590), .B(n12589), .Z(n12975) );
  NAND U13215 ( .A(a[24]), .B(b[24]), .Z(n12974) );
  OR U13216 ( .A(n12975), .B(n12974), .Z(n12591) );
  NAND U13217 ( .A(n12592), .B(n12591), .Z(n12595) );
  ANDN U13218 ( .B(b[24]), .A(n21703), .Z(n12596) );
  OR U13219 ( .A(n12595), .B(n12596), .Z(n12598) );
  XOR U13220 ( .A(n12594), .B(n12593), .Z(n12981) );
  XOR U13221 ( .A(n12596), .B(n12595), .Z(n12980) );
  NANDN U13222 ( .A(n12981), .B(n12980), .Z(n12597) );
  NAND U13223 ( .A(n12598), .B(n12597), .Z(n12601) );
  XNOR U13224 ( .A(n12600), .B(n12599), .Z(n12602) );
  OR U13225 ( .A(n12601), .B(n12602), .Z(n12604) );
  XNOR U13226 ( .A(n12602), .B(n12601), .Z(n12987) );
  NAND U13227 ( .A(a[26]), .B(b[24]), .Z(n12986) );
  OR U13228 ( .A(n12987), .B(n12986), .Z(n12603) );
  NAND U13229 ( .A(n12604), .B(n12603), .Z(n12607) );
  ANDN U13230 ( .B(b[24]), .A(n21716), .Z(n12608) );
  OR U13231 ( .A(n12607), .B(n12608), .Z(n12610) );
  XOR U13232 ( .A(n12606), .B(n12605), .Z(n12993) );
  XOR U13233 ( .A(n12608), .B(n12607), .Z(n12992) );
  NANDN U13234 ( .A(n12993), .B(n12992), .Z(n12609) );
  NAND U13235 ( .A(n12610), .B(n12609), .Z(n12613) );
  XNOR U13236 ( .A(n12612), .B(n12611), .Z(n12614) );
  OR U13237 ( .A(n12613), .B(n12614), .Z(n12616) );
  XNOR U13238 ( .A(n12614), .B(n12613), .Z(n12999) );
  NAND U13239 ( .A(a[28]), .B(b[24]), .Z(n12998) );
  OR U13240 ( .A(n12999), .B(n12998), .Z(n12615) );
  NAND U13241 ( .A(n12616), .B(n12615), .Z(n12619) );
  ANDN U13242 ( .B(b[24]), .A(n21727), .Z(n12620) );
  OR U13243 ( .A(n12619), .B(n12620), .Z(n12622) );
  XOR U13244 ( .A(n12618), .B(n12617), .Z(n13005) );
  XOR U13245 ( .A(n12620), .B(n12619), .Z(n13004) );
  NANDN U13246 ( .A(n13005), .B(n13004), .Z(n12621) );
  NAND U13247 ( .A(n12622), .B(n12621), .Z(n12625) );
  XNOR U13248 ( .A(n12624), .B(n12623), .Z(n12626) );
  OR U13249 ( .A(n12625), .B(n12626), .Z(n12628) );
  XNOR U13250 ( .A(n12626), .B(n12625), .Z(n13011) );
  NAND U13251 ( .A(a[30]), .B(b[24]), .Z(n13010) );
  OR U13252 ( .A(n13011), .B(n13010), .Z(n12627) );
  NAND U13253 ( .A(n12628), .B(n12627), .Z(n12631) );
  ANDN U13254 ( .B(b[24]), .A(n21740), .Z(n12632) );
  OR U13255 ( .A(n12631), .B(n12632), .Z(n12634) );
  XOR U13256 ( .A(n12630), .B(n12629), .Z(n13017) );
  XOR U13257 ( .A(n12632), .B(n12631), .Z(n13016) );
  NANDN U13258 ( .A(n13017), .B(n13016), .Z(n12633) );
  NAND U13259 ( .A(n12634), .B(n12633), .Z(n12637) );
  XNOR U13260 ( .A(n12636), .B(n12635), .Z(n12638) );
  OR U13261 ( .A(n12637), .B(n12638), .Z(n12640) );
  XNOR U13262 ( .A(n12638), .B(n12637), .Z(n13023) );
  NAND U13263 ( .A(a[32]), .B(b[24]), .Z(n13022) );
  OR U13264 ( .A(n13023), .B(n13022), .Z(n12639) );
  NAND U13265 ( .A(n12640), .B(n12639), .Z(n12643) );
  ANDN U13266 ( .B(b[24]), .A(n21751), .Z(n12644) );
  OR U13267 ( .A(n12643), .B(n12644), .Z(n12646) );
  XOR U13268 ( .A(n12642), .B(n12641), .Z(n13029) );
  XOR U13269 ( .A(n12644), .B(n12643), .Z(n13028) );
  NANDN U13270 ( .A(n13029), .B(n13028), .Z(n12645) );
  NAND U13271 ( .A(n12646), .B(n12645), .Z(n12649) );
  XNOR U13272 ( .A(n12648), .B(n12647), .Z(n12650) );
  OR U13273 ( .A(n12649), .B(n12650), .Z(n12652) );
  XNOR U13274 ( .A(n12650), .B(n12649), .Z(n13035) );
  NAND U13275 ( .A(a[34]), .B(b[24]), .Z(n13034) );
  OR U13276 ( .A(n13035), .B(n13034), .Z(n12651) );
  NAND U13277 ( .A(n12652), .B(n12651), .Z(n12655) );
  ANDN U13278 ( .B(b[24]), .A(n184), .Z(n12656) );
  OR U13279 ( .A(n12655), .B(n12656), .Z(n12658) );
  XOR U13280 ( .A(n12656), .B(n12655), .Z(n13040) );
  NANDN U13281 ( .A(n13041), .B(n13040), .Z(n12657) );
  NAND U13282 ( .A(n12658), .B(n12657), .Z(n12661) );
  XOR U13283 ( .A(n12660), .B(n12659), .Z(n12662) );
  OR U13284 ( .A(n12661), .B(n12662), .Z(n12664) );
  NAND U13285 ( .A(a[36]), .B(b[24]), .Z(n13046) );
  XOR U13286 ( .A(n12662), .B(n12661), .Z(n13047) );
  NANDN U13287 ( .A(n13046), .B(n13047), .Z(n12663) );
  NAND U13288 ( .A(n12664), .B(n12663), .Z(n12665) );
  ANDN U13289 ( .B(b[24]), .A(n21772), .Z(n12666) );
  OR U13290 ( .A(n12665), .B(n12666), .Z(n12670) );
  XNOR U13291 ( .A(n12666), .B(n12665), .Z(n13053) );
  XOR U13292 ( .A(n12668), .B(n12667), .Z(n13052) );
  OR U13293 ( .A(n13053), .B(n13052), .Z(n12669) );
  AND U13294 ( .A(n12670), .B(n12669), .Z(n12673) );
  OR U13295 ( .A(n12673), .B(n12674), .Z(n12676) );
  ANDN U13296 ( .B(b[24]), .A(n186), .Z(n13061) );
  XOR U13297 ( .A(n12674), .B(n12673), .Z(n13060) );
  NANDN U13298 ( .A(n13061), .B(n13060), .Z(n12675) );
  AND U13299 ( .A(n12676), .B(n12675), .Z(n12680) );
  OR U13300 ( .A(n12679), .B(n12680), .Z(n12682) );
  XOR U13301 ( .A(n12678), .B(n12677), .Z(n13065) );
  XOR U13302 ( .A(n12680), .B(n12679), .Z(n13064) );
  NANDN U13303 ( .A(n13065), .B(n13064), .Z(n12681) );
  NAND U13304 ( .A(n12682), .B(n12681), .Z(n12686) );
  AND U13305 ( .A(b[24]), .B(a[40]), .Z(n12685) );
  NANDN U13306 ( .A(n12686), .B(n12685), .Z(n12688) );
  XNOR U13307 ( .A(n12686), .B(n12685), .Z(n13072) );
  NANDN U13308 ( .A(n13073), .B(n13072), .Z(n12687) );
  NAND U13309 ( .A(n12688), .B(n12687), .Z(n12692) );
  XOR U13310 ( .A(n12690), .B(n12689), .Z(n12691) );
  NAND U13311 ( .A(n12692), .B(n12691), .Z(n12694) );
  XNOR U13312 ( .A(n12692), .B(n12691), .Z(n13077) );
  NAND U13313 ( .A(a[41]), .B(b[24]), .Z(n13076) );
  OR U13314 ( .A(n13077), .B(n13076), .Z(n12693) );
  NAND U13315 ( .A(n12694), .B(n12693), .Z(n12698) );
  NANDN U13316 ( .A(n12697), .B(n12698), .Z(n12700) );
  XOR U13317 ( .A(n12696), .B(n12695), .Z(n13082) );
  XNOR U13318 ( .A(n12698), .B(n12697), .Z(n13083) );
  NAND U13319 ( .A(n13082), .B(n13083), .Z(n12699) );
  NAND U13320 ( .A(n12700), .B(n12699), .Z(n12703) );
  AND U13321 ( .A(b[24]), .B(a[43]), .Z(n12704) );
  OR U13322 ( .A(n12703), .B(n12704), .Z(n12706) );
  XNOR U13323 ( .A(n12702), .B(n12701), .Z(n13089) );
  XOR U13324 ( .A(n12704), .B(n12703), .Z(n13088) );
  NANDN U13325 ( .A(n13089), .B(n13088), .Z(n12705) );
  NAND U13326 ( .A(n12706), .B(n12705), .Z(n12710) );
  NAND U13327 ( .A(a[44]), .B(b[24]), .Z(n12709) );
  OR U13328 ( .A(n12710), .B(n12709), .Z(n12712) );
  XOR U13329 ( .A(n12708), .B(n12707), .Z(n13094) );
  XOR U13330 ( .A(n12710), .B(n12709), .Z(n13095) );
  NAND U13331 ( .A(n13094), .B(n13095), .Z(n12711) );
  NAND U13332 ( .A(n12712), .B(n12711), .Z(n12715) );
  AND U13333 ( .A(b[24]), .B(a[45]), .Z(n12716) );
  OR U13334 ( .A(n12715), .B(n12716), .Z(n12718) );
  XNOR U13335 ( .A(n12714), .B(n12713), .Z(n13101) );
  XOR U13336 ( .A(n12716), .B(n12715), .Z(n13100) );
  NANDN U13337 ( .A(n13101), .B(n13100), .Z(n12717) );
  NAND U13338 ( .A(n12718), .B(n12717), .Z(n12722) );
  NAND U13339 ( .A(a[46]), .B(b[24]), .Z(n12721) );
  OR U13340 ( .A(n12722), .B(n12721), .Z(n12724) );
  XOR U13341 ( .A(n12720), .B(n12719), .Z(n13106) );
  XOR U13342 ( .A(n12722), .B(n12721), .Z(n13107) );
  NAND U13343 ( .A(n13106), .B(n13107), .Z(n12723) );
  NAND U13344 ( .A(n12724), .B(n12723), .Z(n12727) );
  AND U13345 ( .A(b[24]), .B(a[47]), .Z(n12728) );
  OR U13346 ( .A(n12727), .B(n12728), .Z(n12730) );
  XNOR U13347 ( .A(n12726), .B(n12725), .Z(n13113) );
  XOR U13348 ( .A(n12728), .B(n12727), .Z(n13112) );
  NANDN U13349 ( .A(n13113), .B(n13112), .Z(n12729) );
  NAND U13350 ( .A(n12730), .B(n12729), .Z(n12734) );
  NAND U13351 ( .A(a[48]), .B(b[24]), .Z(n12733) );
  OR U13352 ( .A(n12734), .B(n12733), .Z(n12736) );
  XOR U13353 ( .A(n12732), .B(n12731), .Z(n13118) );
  XOR U13354 ( .A(n12734), .B(n12733), .Z(n13119) );
  NAND U13355 ( .A(n13118), .B(n13119), .Z(n12735) );
  NAND U13356 ( .A(n12736), .B(n12735), .Z(n12739) );
  AND U13357 ( .A(b[24]), .B(a[49]), .Z(n12740) );
  OR U13358 ( .A(n12739), .B(n12740), .Z(n12742) );
  XNOR U13359 ( .A(n12738), .B(n12737), .Z(n13125) );
  XOR U13360 ( .A(n12740), .B(n12739), .Z(n13124) );
  NANDN U13361 ( .A(n13125), .B(n13124), .Z(n12741) );
  NAND U13362 ( .A(n12742), .B(n12741), .Z(n12746) );
  NAND U13363 ( .A(a[50]), .B(b[24]), .Z(n12745) );
  OR U13364 ( .A(n12746), .B(n12745), .Z(n12748) );
  XOR U13365 ( .A(n12744), .B(n12743), .Z(n13130) );
  XOR U13366 ( .A(n12746), .B(n12745), .Z(n13131) );
  NAND U13367 ( .A(n13130), .B(n13131), .Z(n12747) );
  NAND U13368 ( .A(n12748), .B(n12747), .Z(n12751) );
  AND U13369 ( .A(b[24]), .B(a[51]), .Z(n12752) );
  OR U13370 ( .A(n12751), .B(n12752), .Z(n12754) );
  XNOR U13371 ( .A(n12750), .B(n12749), .Z(n13137) );
  XOR U13372 ( .A(n12752), .B(n12751), .Z(n13136) );
  NANDN U13373 ( .A(n13137), .B(n13136), .Z(n12753) );
  NAND U13374 ( .A(n12754), .B(n12753), .Z(n12758) );
  NAND U13375 ( .A(a[52]), .B(b[24]), .Z(n12757) );
  OR U13376 ( .A(n12758), .B(n12757), .Z(n12760) );
  XOR U13377 ( .A(n12756), .B(n12755), .Z(n13142) );
  XOR U13378 ( .A(n12758), .B(n12757), .Z(n13143) );
  NAND U13379 ( .A(n13142), .B(n13143), .Z(n12759) );
  NAND U13380 ( .A(n12760), .B(n12759), .Z(n12763) );
  AND U13381 ( .A(b[24]), .B(a[53]), .Z(n12764) );
  OR U13382 ( .A(n12763), .B(n12764), .Z(n12766) );
  XNOR U13383 ( .A(n12762), .B(n12761), .Z(n13149) );
  XOR U13384 ( .A(n12764), .B(n12763), .Z(n13148) );
  NANDN U13385 ( .A(n13149), .B(n13148), .Z(n12765) );
  NAND U13386 ( .A(n12766), .B(n12765), .Z(n12770) );
  NAND U13387 ( .A(a[54]), .B(b[24]), .Z(n12769) );
  OR U13388 ( .A(n12770), .B(n12769), .Z(n12772) );
  XOR U13389 ( .A(n12768), .B(n12767), .Z(n13154) );
  XOR U13390 ( .A(n12770), .B(n12769), .Z(n13155) );
  NAND U13391 ( .A(n13154), .B(n13155), .Z(n12771) );
  NAND U13392 ( .A(n12772), .B(n12771), .Z(n12775) );
  AND U13393 ( .A(b[24]), .B(a[55]), .Z(n12776) );
  OR U13394 ( .A(n12775), .B(n12776), .Z(n12778) );
  XNOR U13395 ( .A(n12774), .B(n12773), .Z(n13161) );
  XOR U13396 ( .A(n12776), .B(n12775), .Z(n13160) );
  NANDN U13397 ( .A(n13161), .B(n13160), .Z(n12777) );
  NAND U13398 ( .A(n12778), .B(n12777), .Z(n12782) );
  NAND U13399 ( .A(a[56]), .B(b[24]), .Z(n12781) );
  OR U13400 ( .A(n12782), .B(n12781), .Z(n12784) );
  XOR U13401 ( .A(n12780), .B(n12779), .Z(n13166) );
  XOR U13402 ( .A(n12782), .B(n12781), .Z(n13167) );
  NAND U13403 ( .A(n13166), .B(n13167), .Z(n12783) );
  NAND U13404 ( .A(n12784), .B(n12783), .Z(n12787) );
  AND U13405 ( .A(b[24]), .B(a[57]), .Z(n12788) );
  OR U13406 ( .A(n12787), .B(n12788), .Z(n12790) );
  XNOR U13407 ( .A(n12786), .B(n12785), .Z(n13173) );
  XOR U13408 ( .A(n12788), .B(n12787), .Z(n13172) );
  NANDN U13409 ( .A(n13173), .B(n13172), .Z(n12789) );
  NAND U13410 ( .A(n12790), .B(n12789), .Z(n12794) );
  NAND U13411 ( .A(a[58]), .B(b[24]), .Z(n12793) );
  OR U13412 ( .A(n12794), .B(n12793), .Z(n12796) );
  XOR U13413 ( .A(n12792), .B(n12791), .Z(n13178) );
  XOR U13414 ( .A(n12794), .B(n12793), .Z(n13179) );
  NAND U13415 ( .A(n13178), .B(n13179), .Z(n12795) );
  NAND U13416 ( .A(n12796), .B(n12795), .Z(n12799) );
  AND U13417 ( .A(b[24]), .B(a[59]), .Z(n12800) );
  OR U13418 ( .A(n12799), .B(n12800), .Z(n12802) );
  XNOR U13419 ( .A(n12798), .B(n12797), .Z(n13185) );
  XOR U13420 ( .A(n12800), .B(n12799), .Z(n13184) );
  NANDN U13421 ( .A(n13185), .B(n13184), .Z(n12801) );
  NAND U13422 ( .A(n12802), .B(n12801), .Z(n12806) );
  NAND U13423 ( .A(a[60]), .B(b[24]), .Z(n12805) );
  OR U13424 ( .A(n12806), .B(n12805), .Z(n12808) );
  XOR U13425 ( .A(n12804), .B(n12803), .Z(n13190) );
  XOR U13426 ( .A(n12806), .B(n12805), .Z(n13191) );
  NAND U13427 ( .A(n13190), .B(n13191), .Z(n12807) );
  NAND U13428 ( .A(n12808), .B(n12807), .Z(n12811) );
  AND U13429 ( .A(b[24]), .B(a[61]), .Z(n12812) );
  OR U13430 ( .A(n12811), .B(n12812), .Z(n12814) );
  XNOR U13431 ( .A(n12810), .B(n12809), .Z(n13195) );
  XOR U13432 ( .A(n12812), .B(n12811), .Z(n13194) );
  NANDN U13433 ( .A(n13195), .B(n13194), .Z(n12813) );
  NAND U13434 ( .A(n12814), .B(n12813), .Z(n12818) );
  NAND U13435 ( .A(a[62]), .B(b[24]), .Z(n12817) );
  OR U13436 ( .A(n12818), .B(n12817), .Z(n12820) );
  XOR U13437 ( .A(n12816), .B(n12815), .Z(n13200) );
  XOR U13438 ( .A(n12818), .B(n12817), .Z(n13201) );
  NAND U13439 ( .A(n13200), .B(n13201), .Z(n12819) );
  NAND U13440 ( .A(n12820), .B(n12819), .Z(n12823) );
  AND U13441 ( .A(b[24]), .B(a[63]), .Z(n12824) );
  OR U13442 ( .A(n12823), .B(n12824), .Z(n12826) );
  XOR U13443 ( .A(n12822), .B(n12821), .Z(n13207) );
  XOR U13444 ( .A(n12824), .B(n12823), .Z(n13206) );
  NANDN U13445 ( .A(n13207), .B(n13206), .Z(n12825) );
  NAND U13446 ( .A(n12826), .B(n12825), .Z(n12831) );
  OR U13447 ( .A(n12832), .B(n12831), .Z(n12830) );
  XOR U13448 ( .A(n12828), .B(n12827), .Z(n12829) );
  NAND U13449 ( .A(n12830), .B(n12829), .Z(n21973) );
  XNOR U13450 ( .A(n12830), .B(n12829), .Z(n24173) );
  XOR U13451 ( .A(n12832), .B(n12831), .Z(n21970) );
  NAND U13452 ( .A(a[60]), .B(b[23]), .Z(n13186) );
  NAND U13453 ( .A(a[58]), .B(b[23]), .Z(n13174) );
  NAND U13454 ( .A(a[56]), .B(b[23]), .Z(n13162) );
  NAND U13455 ( .A(a[54]), .B(b[23]), .Z(n13150) );
  NAND U13456 ( .A(a[52]), .B(b[23]), .Z(n13138) );
  NAND U13457 ( .A(a[50]), .B(b[23]), .Z(n13126) );
  NAND U13458 ( .A(a[48]), .B(b[23]), .Z(n13114) );
  NAND U13459 ( .A(a[46]), .B(b[23]), .Z(n13102) );
  NAND U13460 ( .A(a[44]), .B(b[23]), .Z(n13090) );
  ANDN U13461 ( .B(b[23]), .A(n21772), .Z(n13049) );
  ANDN U13462 ( .B(b[23]), .A(n184), .Z(n13037) );
  ANDN U13463 ( .B(b[23]), .A(n21751), .Z(n13025) );
  ANDN U13464 ( .B(b[23]), .A(n21740), .Z(n13013) );
  ANDN U13465 ( .B(b[23]), .A(n21727), .Z(n13001) );
  ANDN U13466 ( .B(b[23]), .A(n21716), .Z(n12989) );
  ANDN U13467 ( .B(b[23]), .A(n21703), .Z(n12977) );
  ANDN U13468 ( .B(b[23]), .A(n21692), .Z(n12965) );
  ANDN U13469 ( .B(b[23]), .A(n21681), .Z(n12953) );
  ANDN U13470 ( .B(b[23]), .A(n21670), .Z(n12938) );
  ANDN U13471 ( .B(b[23]), .A(n174), .Z(n12929) );
  ANDN U13472 ( .B(b[23]), .A(n172), .Z(n12917) );
  ANDN U13473 ( .B(b[23]), .A(n170), .Z(n12907) );
  ANDN U13474 ( .B(b[23]), .A(n21164), .Z(n12893) );
  ANDN U13475 ( .B(b[23]), .A(n21615), .Z(n12881) );
  ANDN U13476 ( .B(b[23]), .A(n166), .Z(n12868) );
  XNOR U13477 ( .A(n12836), .B(n12835), .Z(n12865) );
  ANDN U13478 ( .B(b[23]), .A(n164), .Z(n12861) );
  ANDN U13479 ( .B(b[23]), .A(n21580), .Z(n12846) );
  NAND U13480 ( .A(b[24]), .B(a[1]), .Z(n12839) );
  AND U13481 ( .A(b[23]), .B(a[0]), .Z(n13603) );
  NANDN U13482 ( .A(n12839), .B(n13603), .Z(n12838) );
  NAND U13483 ( .A(a[2]), .B(b[23]), .Z(n12837) );
  AND U13484 ( .A(n12838), .B(n12837), .Z(n12845) );
  NANDN U13485 ( .A(n12839), .B(a[0]), .Z(n12840) );
  XNOR U13486 ( .A(a[2]), .B(n12840), .Z(n12841) );
  NAND U13487 ( .A(b[23]), .B(n12841), .Z(n13230) );
  AND U13488 ( .A(a[1]), .B(b[24]), .Z(n12842) );
  XNOR U13489 ( .A(n12843), .B(n12842), .Z(n13229) );
  NANDN U13490 ( .A(n13230), .B(n13229), .Z(n12844) );
  NANDN U13491 ( .A(n12845), .B(n12844), .Z(n12847) );
  NANDN U13492 ( .A(n12846), .B(n12847), .Z(n12851) );
  XOR U13493 ( .A(n12847), .B(n12846), .Z(n13234) );
  NANDN U13494 ( .A(n13234), .B(n13233), .Z(n12850) );
  NAND U13495 ( .A(n12851), .B(n12850), .Z(n12855) );
  XOR U13496 ( .A(n12853), .B(n12852), .Z(n12854) );
  NANDN U13497 ( .A(n12855), .B(n12854), .Z(n12857) );
  NAND U13498 ( .A(a[4]), .B(b[23]), .Z(n13241) );
  NANDN U13499 ( .A(n13241), .B(n13242), .Z(n12856) );
  NAND U13500 ( .A(n12857), .B(n12856), .Z(n12860) );
  OR U13501 ( .A(n12861), .B(n12860), .Z(n12863) );
  XOR U13502 ( .A(n12859), .B(n12858), .Z(n13217) );
  XOR U13503 ( .A(n12861), .B(n12860), .Z(n13216) );
  NAND U13504 ( .A(n13217), .B(n13216), .Z(n12862) );
  NAND U13505 ( .A(n12863), .B(n12862), .Z(n12864) );
  NANDN U13506 ( .A(n12865), .B(n12864), .Z(n12867) );
  ANDN U13507 ( .B(b[23]), .A(n165), .Z(n13252) );
  NANDN U13508 ( .A(n13252), .B(n13251), .Z(n12866) );
  NAND U13509 ( .A(n12867), .B(n12866), .Z(n12869) );
  NANDN U13510 ( .A(n12868), .B(n12869), .Z(n12873) );
  XOR U13511 ( .A(n12869), .B(n12868), .Z(n13256) );
  XOR U13512 ( .A(n12871), .B(n12870), .Z(n13255) );
  OR U13513 ( .A(n13256), .B(n13255), .Z(n12872) );
  NAND U13514 ( .A(n12873), .B(n12872), .Z(n12877) );
  XNOR U13515 ( .A(n12875), .B(n12874), .Z(n12876) );
  NANDN U13516 ( .A(n12877), .B(n12876), .Z(n12879) );
  NAND U13517 ( .A(a[8]), .B(b[23]), .Z(n13261) );
  NANDN U13518 ( .A(n13261), .B(n13262), .Z(n12878) );
  NAND U13519 ( .A(n12879), .B(n12878), .Z(n12880) );
  OR U13520 ( .A(n12881), .B(n12880), .Z(n12885) );
  XNOR U13521 ( .A(n12881), .B(n12880), .Z(n13267) );
  XOR U13522 ( .A(n12883), .B(n12882), .Z(n13268) );
  NANDN U13523 ( .A(n13267), .B(n13268), .Z(n12884) );
  NAND U13524 ( .A(n12885), .B(n12884), .Z(n12888) );
  XOR U13525 ( .A(n12887), .B(n12886), .Z(n12889) );
  NANDN U13526 ( .A(n12888), .B(n12889), .Z(n12891) );
  NAND U13527 ( .A(a[10]), .B(b[23]), .Z(n13275) );
  XNOR U13528 ( .A(n12889), .B(n12888), .Z(n13276) );
  NANDN U13529 ( .A(n13275), .B(n13276), .Z(n12890) );
  NAND U13530 ( .A(n12891), .B(n12890), .Z(n12892) );
  OR U13531 ( .A(n12893), .B(n12892), .Z(n12897) );
  XNOR U13532 ( .A(n12893), .B(n12892), .Z(n13279) );
  XOR U13533 ( .A(n12895), .B(n12894), .Z(n13280) );
  NANDN U13534 ( .A(n13279), .B(n13280), .Z(n12896) );
  NAND U13535 ( .A(n12897), .B(n12896), .Z(n12900) );
  XOR U13536 ( .A(n12899), .B(n12898), .Z(n12901) );
  NANDN U13537 ( .A(n12900), .B(n12901), .Z(n12903) );
  NAND U13538 ( .A(a[12]), .B(b[23]), .Z(n13287) );
  XNOR U13539 ( .A(n12901), .B(n12900), .Z(n13288) );
  NANDN U13540 ( .A(n13287), .B(n13288), .Z(n12902) );
  NAND U13541 ( .A(n12903), .B(n12902), .Z(n12906) );
  OR U13542 ( .A(n12907), .B(n12906), .Z(n12909) );
  XOR U13543 ( .A(n12905), .B(n12904), .Z(n13214) );
  XOR U13544 ( .A(n12907), .B(n12906), .Z(n13215) );
  NAND U13545 ( .A(n13214), .B(n13215), .Z(n12908) );
  NAND U13546 ( .A(n12909), .B(n12908), .Z(n12912) );
  NANDN U13547 ( .A(n12912), .B(n12913), .Z(n12915) );
  NAND U13548 ( .A(a[14]), .B(b[23]), .Z(n13297) );
  XNOR U13549 ( .A(n12913), .B(n12912), .Z(n13298) );
  NANDN U13550 ( .A(n13297), .B(n13298), .Z(n12914) );
  NAND U13551 ( .A(n12915), .B(n12914), .Z(n12916) );
  OR U13552 ( .A(n12917), .B(n12916), .Z(n12921) );
  XNOR U13553 ( .A(n12917), .B(n12916), .Z(n13301) );
  XOR U13554 ( .A(n12919), .B(n12918), .Z(n13302) );
  NANDN U13555 ( .A(n13301), .B(n13302), .Z(n12920) );
  NAND U13556 ( .A(n12921), .B(n12920), .Z(n12922) );
  OR U13557 ( .A(n12923), .B(n12922), .Z(n12925) );
  NAND U13558 ( .A(a[16]), .B(b[23]), .Z(n13309) );
  XOR U13559 ( .A(n12923), .B(n12922), .Z(n13310) );
  NANDN U13560 ( .A(n13309), .B(n13310), .Z(n12924) );
  NAND U13561 ( .A(n12925), .B(n12924), .Z(n12928) );
  OR U13562 ( .A(n12929), .B(n12928), .Z(n12931) );
  XOR U13563 ( .A(n12927), .B(n12926), .Z(n13212) );
  XOR U13564 ( .A(n12929), .B(n12928), .Z(n13213) );
  NAND U13565 ( .A(n13212), .B(n13213), .Z(n12930) );
  NAND U13566 ( .A(n12931), .B(n12930), .Z(n12935) );
  XOR U13567 ( .A(n12933), .B(n12932), .Z(n12934) );
  NAND U13568 ( .A(n12935), .B(n12934), .Z(n12937) );
  ANDN U13569 ( .B(b[23]), .A(n175), .Z(n13318) );
  XNOR U13570 ( .A(n12935), .B(n12934), .Z(n13317) );
  OR U13571 ( .A(n13318), .B(n13317), .Z(n12936) );
  NAND U13572 ( .A(n12937), .B(n12936), .Z(n12939) );
  NANDN U13573 ( .A(n12938), .B(n12939), .Z(n12943) );
  XOR U13574 ( .A(n12939), .B(n12938), .Z(n13324) );
  XOR U13575 ( .A(n12941), .B(n12940), .Z(n13323) );
  OR U13576 ( .A(n13324), .B(n13323), .Z(n12942) );
  NAND U13577 ( .A(n12943), .B(n12942), .Z(n12946) );
  NANDN U13578 ( .A(n12946), .B(n12947), .Z(n12949) );
  NAND U13579 ( .A(a[20]), .B(b[23]), .Z(n13331) );
  XNOR U13580 ( .A(n12947), .B(n12946), .Z(n13332) );
  NANDN U13581 ( .A(n13331), .B(n13332), .Z(n12948) );
  NAND U13582 ( .A(n12949), .B(n12948), .Z(n12952) );
  OR U13583 ( .A(n12953), .B(n12952), .Z(n12955) );
  XNOR U13584 ( .A(n12951), .B(n12950), .Z(n13336) );
  XOR U13585 ( .A(n12953), .B(n12952), .Z(n13335) );
  NAND U13586 ( .A(n13336), .B(n13335), .Z(n12954) );
  NAND U13587 ( .A(n12955), .B(n12954), .Z(n12958) );
  NANDN U13588 ( .A(n12958), .B(n12959), .Z(n12961) );
  NAND U13589 ( .A(a[22]), .B(b[23]), .Z(n13343) );
  XNOR U13590 ( .A(n12959), .B(n12958), .Z(n13344) );
  NANDN U13591 ( .A(n13343), .B(n13344), .Z(n12960) );
  NAND U13592 ( .A(n12961), .B(n12960), .Z(n12964) );
  OR U13593 ( .A(n12965), .B(n12964), .Z(n12967) );
  XNOR U13594 ( .A(n12963), .B(n12962), .Z(n13348) );
  XOR U13595 ( .A(n12965), .B(n12964), .Z(n13347) );
  NAND U13596 ( .A(n13348), .B(n13347), .Z(n12966) );
  NAND U13597 ( .A(n12967), .B(n12966), .Z(n12970) );
  NANDN U13598 ( .A(n12970), .B(n12971), .Z(n12973) );
  NAND U13599 ( .A(a[24]), .B(b[23]), .Z(n13355) );
  XNOR U13600 ( .A(n12971), .B(n12970), .Z(n13356) );
  NANDN U13601 ( .A(n13355), .B(n13356), .Z(n12972) );
  NAND U13602 ( .A(n12973), .B(n12972), .Z(n12976) );
  OR U13603 ( .A(n12977), .B(n12976), .Z(n12979) );
  XNOR U13604 ( .A(n12975), .B(n12974), .Z(n13360) );
  XOR U13605 ( .A(n12977), .B(n12976), .Z(n13359) );
  NAND U13606 ( .A(n13360), .B(n13359), .Z(n12978) );
  NAND U13607 ( .A(n12979), .B(n12978), .Z(n12982) );
  NANDN U13608 ( .A(n12982), .B(n12983), .Z(n12985) );
  NAND U13609 ( .A(a[26]), .B(b[23]), .Z(n13367) );
  XNOR U13610 ( .A(n12983), .B(n12982), .Z(n13368) );
  NANDN U13611 ( .A(n13367), .B(n13368), .Z(n12984) );
  NAND U13612 ( .A(n12985), .B(n12984), .Z(n12988) );
  OR U13613 ( .A(n12989), .B(n12988), .Z(n12991) );
  XNOR U13614 ( .A(n12987), .B(n12986), .Z(n13372) );
  XOR U13615 ( .A(n12989), .B(n12988), .Z(n13371) );
  NAND U13616 ( .A(n13372), .B(n13371), .Z(n12990) );
  NAND U13617 ( .A(n12991), .B(n12990), .Z(n12994) );
  NANDN U13618 ( .A(n12994), .B(n12995), .Z(n12997) );
  NAND U13619 ( .A(a[28]), .B(b[23]), .Z(n13379) );
  XNOR U13620 ( .A(n12995), .B(n12994), .Z(n13380) );
  NANDN U13621 ( .A(n13379), .B(n13380), .Z(n12996) );
  NAND U13622 ( .A(n12997), .B(n12996), .Z(n13000) );
  OR U13623 ( .A(n13001), .B(n13000), .Z(n13003) );
  XNOR U13624 ( .A(n12999), .B(n12998), .Z(n13384) );
  XOR U13625 ( .A(n13001), .B(n13000), .Z(n13383) );
  NAND U13626 ( .A(n13384), .B(n13383), .Z(n13002) );
  NAND U13627 ( .A(n13003), .B(n13002), .Z(n13006) );
  NANDN U13628 ( .A(n13006), .B(n13007), .Z(n13009) );
  NAND U13629 ( .A(a[30]), .B(b[23]), .Z(n13391) );
  XNOR U13630 ( .A(n13007), .B(n13006), .Z(n13392) );
  NANDN U13631 ( .A(n13391), .B(n13392), .Z(n13008) );
  NAND U13632 ( .A(n13009), .B(n13008), .Z(n13012) );
  OR U13633 ( .A(n13013), .B(n13012), .Z(n13015) );
  XNOR U13634 ( .A(n13011), .B(n13010), .Z(n13396) );
  XOR U13635 ( .A(n13013), .B(n13012), .Z(n13395) );
  NAND U13636 ( .A(n13396), .B(n13395), .Z(n13014) );
  NAND U13637 ( .A(n13015), .B(n13014), .Z(n13018) );
  NANDN U13638 ( .A(n13018), .B(n13019), .Z(n13021) );
  NAND U13639 ( .A(a[32]), .B(b[23]), .Z(n13403) );
  XNOR U13640 ( .A(n13019), .B(n13018), .Z(n13404) );
  NANDN U13641 ( .A(n13403), .B(n13404), .Z(n13020) );
  NAND U13642 ( .A(n13021), .B(n13020), .Z(n13024) );
  OR U13643 ( .A(n13025), .B(n13024), .Z(n13027) );
  XNOR U13644 ( .A(n13023), .B(n13022), .Z(n13408) );
  XOR U13645 ( .A(n13025), .B(n13024), .Z(n13407) );
  NAND U13646 ( .A(n13408), .B(n13407), .Z(n13026) );
  NAND U13647 ( .A(n13027), .B(n13026), .Z(n13030) );
  NANDN U13648 ( .A(n13030), .B(n13031), .Z(n13033) );
  NAND U13649 ( .A(a[34]), .B(b[23]), .Z(n13415) );
  XNOR U13650 ( .A(n13031), .B(n13030), .Z(n13416) );
  NANDN U13651 ( .A(n13415), .B(n13416), .Z(n13032) );
  NAND U13652 ( .A(n13033), .B(n13032), .Z(n13036) );
  OR U13653 ( .A(n13037), .B(n13036), .Z(n13039) );
  XNOR U13654 ( .A(n13035), .B(n13034), .Z(n13420) );
  XOR U13655 ( .A(n13037), .B(n13036), .Z(n13419) );
  NAND U13656 ( .A(n13420), .B(n13419), .Z(n13038) );
  NAND U13657 ( .A(n13039), .B(n13038), .Z(n13042) );
  NANDN U13658 ( .A(n13042), .B(n13043), .Z(n13045) );
  NAND U13659 ( .A(a[36]), .B(b[23]), .Z(n13427) );
  XNOR U13660 ( .A(n13043), .B(n13042), .Z(n13428) );
  NANDN U13661 ( .A(n13427), .B(n13428), .Z(n13044) );
  NAND U13662 ( .A(n13045), .B(n13044), .Z(n13048) );
  OR U13663 ( .A(n13049), .B(n13048), .Z(n13051) );
  XNOR U13664 ( .A(n13047), .B(n13046), .Z(n13432) );
  XOR U13665 ( .A(n13049), .B(n13048), .Z(n13431) );
  NANDN U13666 ( .A(n13432), .B(n13431), .Z(n13050) );
  NAND U13667 ( .A(n13051), .B(n13050), .Z(n13054) );
  XNOR U13668 ( .A(n13053), .B(n13052), .Z(n13055) );
  NANDN U13669 ( .A(n13054), .B(n13055), .Z(n13057) );
  NAND U13670 ( .A(a[38]), .B(b[23]), .Z(n13439) );
  XNOR U13671 ( .A(n13055), .B(n13054), .Z(n13440) );
  NANDN U13672 ( .A(n13439), .B(n13440), .Z(n13056) );
  NAND U13673 ( .A(n13057), .B(n13056), .Z(n13058) );
  ANDN U13674 ( .B(b[23]), .A(n187), .Z(n13059) );
  OR U13675 ( .A(n13058), .B(n13059), .Z(n13063) );
  XNOR U13676 ( .A(n13059), .B(n13058), .Z(n13444) );
  XOR U13677 ( .A(n13061), .B(n13060), .Z(n13443) );
  OR U13678 ( .A(n13444), .B(n13443), .Z(n13062) );
  NAND U13679 ( .A(n13063), .B(n13062), .Z(n13066) );
  XNOR U13680 ( .A(n13065), .B(n13064), .Z(n13067) );
  OR U13681 ( .A(n13066), .B(n13067), .Z(n13069) );
  XNOR U13682 ( .A(n13067), .B(n13066), .Z(n13450) );
  NAND U13683 ( .A(a[40]), .B(b[23]), .Z(n13449) );
  OR U13684 ( .A(n13450), .B(n13449), .Z(n13068) );
  NAND U13685 ( .A(n13069), .B(n13068), .Z(n13070) );
  ANDN U13686 ( .B(b[23]), .A(n189), .Z(n13071) );
  OR U13687 ( .A(n13070), .B(n13071), .Z(n13075) );
  XOR U13688 ( .A(n13071), .B(n13070), .Z(n13455) );
  NAND U13689 ( .A(n13455), .B(n13456), .Z(n13074) );
  NAND U13690 ( .A(n13075), .B(n13074), .Z(n13079) );
  NAND U13691 ( .A(a[42]), .B(b[23]), .Z(n13078) );
  OR U13692 ( .A(n13079), .B(n13078), .Z(n13081) );
  XOR U13693 ( .A(n13077), .B(n13076), .Z(n13461) );
  XOR U13694 ( .A(n13079), .B(n13078), .Z(n13462) );
  NAND U13695 ( .A(n13461), .B(n13462), .Z(n13080) );
  NAND U13696 ( .A(n13081), .B(n13080), .Z(n13085) );
  XOR U13697 ( .A(n13083), .B(n13082), .Z(n13084) );
  NAND U13698 ( .A(n13085), .B(n13084), .Z(n13087) );
  XNOR U13699 ( .A(n13085), .B(n13084), .Z(n13468) );
  NAND U13700 ( .A(a[43]), .B(b[23]), .Z(n13467) );
  OR U13701 ( .A(n13468), .B(n13467), .Z(n13086) );
  NAND U13702 ( .A(n13087), .B(n13086), .Z(n13091) );
  NANDN U13703 ( .A(n13090), .B(n13091), .Z(n13093) );
  XNOR U13704 ( .A(n13089), .B(n13088), .Z(n13474) );
  XNOR U13705 ( .A(n13091), .B(n13090), .Z(n13473) );
  NANDN U13706 ( .A(n13474), .B(n13473), .Z(n13092) );
  NAND U13707 ( .A(n13093), .B(n13092), .Z(n13097) );
  XOR U13708 ( .A(n13095), .B(n13094), .Z(n13096) );
  NAND U13709 ( .A(n13097), .B(n13096), .Z(n13099) );
  XNOR U13710 ( .A(n13097), .B(n13096), .Z(n13480) );
  NAND U13711 ( .A(a[45]), .B(b[23]), .Z(n13479) );
  OR U13712 ( .A(n13480), .B(n13479), .Z(n13098) );
  NAND U13713 ( .A(n13099), .B(n13098), .Z(n13103) );
  NANDN U13714 ( .A(n13102), .B(n13103), .Z(n13105) );
  XNOR U13715 ( .A(n13101), .B(n13100), .Z(n13486) );
  XNOR U13716 ( .A(n13103), .B(n13102), .Z(n13485) );
  NANDN U13717 ( .A(n13486), .B(n13485), .Z(n13104) );
  NAND U13718 ( .A(n13105), .B(n13104), .Z(n13109) );
  XOR U13719 ( .A(n13107), .B(n13106), .Z(n13108) );
  NAND U13720 ( .A(n13109), .B(n13108), .Z(n13111) );
  XNOR U13721 ( .A(n13109), .B(n13108), .Z(n13492) );
  NAND U13722 ( .A(a[47]), .B(b[23]), .Z(n13491) );
  OR U13723 ( .A(n13492), .B(n13491), .Z(n13110) );
  NAND U13724 ( .A(n13111), .B(n13110), .Z(n13115) );
  NANDN U13725 ( .A(n13114), .B(n13115), .Z(n13117) );
  XNOR U13726 ( .A(n13113), .B(n13112), .Z(n13498) );
  XNOR U13727 ( .A(n13115), .B(n13114), .Z(n13497) );
  NANDN U13728 ( .A(n13498), .B(n13497), .Z(n13116) );
  NAND U13729 ( .A(n13117), .B(n13116), .Z(n13121) );
  XOR U13730 ( .A(n13119), .B(n13118), .Z(n13120) );
  NAND U13731 ( .A(n13121), .B(n13120), .Z(n13123) );
  XNOR U13732 ( .A(n13121), .B(n13120), .Z(n13504) );
  NAND U13733 ( .A(a[49]), .B(b[23]), .Z(n13503) );
  OR U13734 ( .A(n13504), .B(n13503), .Z(n13122) );
  NAND U13735 ( .A(n13123), .B(n13122), .Z(n13127) );
  NANDN U13736 ( .A(n13126), .B(n13127), .Z(n13129) );
  XNOR U13737 ( .A(n13125), .B(n13124), .Z(n13510) );
  XNOR U13738 ( .A(n13127), .B(n13126), .Z(n13509) );
  NANDN U13739 ( .A(n13510), .B(n13509), .Z(n13128) );
  NAND U13740 ( .A(n13129), .B(n13128), .Z(n13133) );
  XOR U13741 ( .A(n13131), .B(n13130), .Z(n13132) );
  NAND U13742 ( .A(n13133), .B(n13132), .Z(n13135) );
  XNOR U13743 ( .A(n13133), .B(n13132), .Z(n13516) );
  NAND U13744 ( .A(a[51]), .B(b[23]), .Z(n13515) );
  OR U13745 ( .A(n13516), .B(n13515), .Z(n13134) );
  NAND U13746 ( .A(n13135), .B(n13134), .Z(n13139) );
  NANDN U13747 ( .A(n13138), .B(n13139), .Z(n13141) );
  XNOR U13748 ( .A(n13137), .B(n13136), .Z(n13522) );
  XNOR U13749 ( .A(n13139), .B(n13138), .Z(n13521) );
  NANDN U13750 ( .A(n13522), .B(n13521), .Z(n13140) );
  NAND U13751 ( .A(n13141), .B(n13140), .Z(n13145) );
  XOR U13752 ( .A(n13143), .B(n13142), .Z(n13144) );
  NAND U13753 ( .A(n13145), .B(n13144), .Z(n13147) );
  XNOR U13754 ( .A(n13145), .B(n13144), .Z(n13528) );
  NAND U13755 ( .A(a[53]), .B(b[23]), .Z(n13527) );
  OR U13756 ( .A(n13528), .B(n13527), .Z(n13146) );
  NAND U13757 ( .A(n13147), .B(n13146), .Z(n13151) );
  NANDN U13758 ( .A(n13150), .B(n13151), .Z(n13153) );
  XNOR U13759 ( .A(n13149), .B(n13148), .Z(n13534) );
  XNOR U13760 ( .A(n13151), .B(n13150), .Z(n13533) );
  NANDN U13761 ( .A(n13534), .B(n13533), .Z(n13152) );
  NAND U13762 ( .A(n13153), .B(n13152), .Z(n13157) );
  XOR U13763 ( .A(n13155), .B(n13154), .Z(n13156) );
  NAND U13764 ( .A(n13157), .B(n13156), .Z(n13159) );
  XNOR U13765 ( .A(n13157), .B(n13156), .Z(n13540) );
  NAND U13766 ( .A(a[55]), .B(b[23]), .Z(n13539) );
  OR U13767 ( .A(n13540), .B(n13539), .Z(n13158) );
  NAND U13768 ( .A(n13159), .B(n13158), .Z(n13163) );
  NANDN U13769 ( .A(n13162), .B(n13163), .Z(n13165) );
  XNOR U13770 ( .A(n13161), .B(n13160), .Z(n13546) );
  XNOR U13771 ( .A(n13163), .B(n13162), .Z(n13545) );
  NANDN U13772 ( .A(n13546), .B(n13545), .Z(n13164) );
  NAND U13773 ( .A(n13165), .B(n13164), .Z(n13169) );
  XOR U13774 ( .A(n13167), .B(n13166), .Z(n13168) );
  NAND U13775 ( .A(n13169), .B(n13168), .Z(n13171) );
  XNOR U13776 ( .A(n13169), .B(n13168), .Z(n13552) );
  NAND U13777 ( .A(a[57]), .B(b[23]), .Z(n13551) );
  OR U13778 ( .A(n13552), .B(n13551), .Z(n13170) );
  NAND U13779 ( .A(n13171), .B(n13170), .Z(n13175) );
  NANDN U13780 ( .A(n13174), .B(n13175), .Z(n13177) );
  XNOR U13781 ( .A(n13173), .B(n13172), .Z(n13558) );
  XNOR U13782 ( .A(n13175), .B(n13174), .Z(n13557) );
  NANDN U13783 ( .A(n13558), .B(n13557), .Z(n13176) );
  NAND U13784 ( .A(n13177), .B(n13176), .Z(n13181) );
  XOR U13785 ( .A(n13179), .B(n13178), .Z(n13180) );
  NAND U13786 ( .A(n13181), .B(n13180), .Z(n13183) );
  XNOR U13787 ( .A(n13181), .B(n13180), .Z(n13564) );
  NAND U13788 ( .A(a[59]), .B(b[23]), .Z(n13563) );
  OR U13789 ( .A(n13564), .B(n13563), .Z(n13182) );
  NAND U13790 ( .A(n13183), .B(n13182), .Z(n13187) );
  NANDN U13791 ( .A(n13186), .B(n13187), .Z(n13189) );
  XNOR U13792 ( .A(n13185), .B(n13184), .Z(n13570) );
  XNOR U13793 ( .A(n13187), .B(n13186), .Z(n13569) );
  NANDN U13794 ( .A(n13570), .B(n13569), .Z(n13188) );
  NAND U13795 ( .A(n13189), .B(n13188), .Z(n13192) );
  XOR U13796 ( .A(n13191), .B(n13190), .Z(n13193) );
  AND U13797 ( .A(b[23]), .B(a[61]), .Z(n13576) );
  XOR U13798 ( .A(n13193), .B(n13192), .Z(n13575) );
  NAND U13799 ( .A(a[62]), .B(b[23]), .Z(n13196) );
  OR U13800 ( .A(n13197), .B(n13196), .Z(n13199) );
  XNOR U13801 ( .A(n13195), .B(n13194), .Z(n13582) );
  XOR U13802 ( .A(n13197), .B(n13196), .Z(n13581) );
  NANDN U13803 ( .A(n13582), .B(n13581), .Z(n13198) );
  NAND U13804 ( .A(n13199), .B(n13198), .Z(n13203) );
  XOR U13805 ( .A(n13201), .B(n13200), .Z(n13202) );
  NAND U13806 ( .A(n13203), .B(n13202), .Z(n13205) );
  XNOR U13807 ( .A(n13203), .B(n13202), .Z(n13211) );
  NAND U13808 ( .A(a[63]), .B(b[23]), .Z(n13210) );
  OR U13809 ( .A(n13211), .B(n13210), .Z(n13204) );
  NAND U13810 ( .A(n13205), .B(n13204), .Z(n13208) );
  XNOR U13811 ( .A(n13207), .B(n13206), .Z(n13209) );
  ANDN U13812 ( .B(n13208), .A(n13209), .Z(n21971) );
  XNOR U13813 ( .A(n13209), .B(n13208), .Z(n21968) );
  XNOR U13814 ( .A(n13211), .B(n13210), .Z(n13588) );
  NAND U13815 ( .A(a[44]), .B(b[22]), .Z(n13469) );
  ANDN U13816 ( .B(b[22]), .A(n187), .Z(n13438) );
  ANDN U13817 ( .B(b[22]), .A(n21772), .Z(n13426) );
  ANDN U13818 ( .B(b[22]), .A(n184), .Z(n13414) );
  ANDN U13819 ( .B(b[22]), .A(n21751), .Z(n13402) );
  ANDN U13820 ( .B(b[22]), .A(n21740), .Z(n13390) );
  ANDN U13821 ( .B(b[22]), .A(n21727), .Z(n13378) );
  ANDN U13822 ( .B(b[22]), .A(n21716), .Z(n13366) );
  ANDN U13823 ( .B(b[22]), .A(n21703), .Z(n13354) );
  ANDN U13824 ( .B(b[22]), .A(n21692), .Z(n13342) );
  ANDN U13825 ( .B(b[22]), .A(n21681), .Z(n13330) );
  ANDN U13826 ( .B(b[22]), .A(n21670), .Z(n13320) );
  ANDN U13827 ( .B(b[22]), .A(n174), .Z(n13308) );
  ANDN U13828 ( .B(b[22]), .A(n172), .Z(n13296) );
  ANDN U13829 ( .B(b[22]), .A(n170), .Z(n13286) );
  ANDN U13830 ( .B(b[22]), .A(n21164), .Z(n13274) );
  ANDN U13831 ( .B(b[22]), .A(n21615), .Z(n13264) );
  ANDN U13832 ( .B(b[22]), .A(n166), .Z(n13249) );
  XNOR U13833 ( .A(n13217), .B(n13216), .Z(n13246) );
  ANDN U13834 ( .B(b[22]), .A(n164), .Z(n13240) );
  ANDN U13835 ( .B(b[22]), .A(n21580), .Z(n13227) );
  NAND U13836 ( .A(b[23]), .B(a[1]), .Z(n13220) );
  AND U13837 ( .A(b[22]), .B(a[0]), .Z(n13984) );
  NANDN U13838 ( .A(n13220), .B(n13984), .Z(n13219) );
  NAND U13839 ( .A(a[2]), .B(b[22]), .Z(n13218) );
  AND U13840 ( .A(n13219), .B(n13218), .Z(n13226) );
  NANDN U13841 ( .A(n13220), .B(a[0]), .Z(n13221) );
  XNOR U13842 ( .A(a[2]), .B(n13221), .Z(n13222) );
  NAND U13843 ( .A(b[22]), .B(n13222), .Z(n13609) );
  AND U13844 ( .A(a[1]), .B(b[23]), .Z(n13223) );
  XNOR U13845 ( .A(n13224), .B(n13223), .Z(n13608) );
  NANDN U13846 ( .A(n13609), .B(n13608), .Z(n13225) );
  NANDN U13847 ( .A(n13226), .B(n13225), .Z(n13228) );
  NANDN U13848 ( .A(n13227), .B(n13228), .Z(n13232) );
  XOR U13849 ( .A(n13228), .B(n13227), .Z(n13613) );
  NANDN U13850 ( .A(n13613), .B(n13612), .Z(n13231) );
  NAND U13851 ( .A(n13232), .B(n13231), .Z(n13236) );
  XOR U13852 ( .A(n13234), .B(n13233), .Z(n13235) );
  NANDN U13853 ( .A(n13236), .B(n13235), .Z(n13238) );
  NAND U13854 ( .A(a[4]), .B(b[22]), .Z(n13620) );
  NANDN U13855 ( .A(n13620), .B(n13621), .Z(n13237) );
  NAND U13856 ( .A(n13238), .B(n13237), .Z(n13239) );
  OR U13857 ( .A(n13240), .B(n13239), .Z(n13244) );
  XNOR U13858 ( .A(n13240), .B(n13239), .Z(n13624) );
  XOR U13859 ( .A(n13242), .B(n13241), .Z(n13625) );
  NANDN U13860 ( .A(n13624), .B(n13625), .Z(n13243) );
  NAND U13861 ( .A(n13244), .B(n13243), .Z(n13245) );
  NANDN U13862 ( .A(n13246), .B(n13245), .Z(n13248) );
  ANDN U13863 ( .B(b[22]), .A(n165), .Z(n13631) );
  NANDN U13864 ( .A(n13631), .B(n13630), .Z(n13247) );
  NAND U13865 ( .A(n13248), .B(n13247), .Z(n13250) );
  NANDN U13866 ( .A(n13249), .B(n13250), .Z(n13254) );
  XOR U13867 ( .A(n13250), .B(n13249), .Z(n13637) );
  XOR U13868 ( .A(n13252), .B(n13251), .Z(n13636) );
  OR U13869 ( .A(n13637), .B(n13636), .Z(n13253) );
  NAND U13870 ( .A(n13254), .B(n13253), .Z(n13258) );
  XNOR U13871 ( .A(n13256), .B(n13255), .Z(n13257) );
  NANDN U13872 ( .A(n13258), .B(n13257), .Z(n13260) );
  NAND U13873 ( .A(a[8]), .B(b[22]), .Z(n13642) );
  NANDN U13874 ( .A(n13642), .B(n13643), .Z(n13259) );
  NAND U13875 ( .A(n13260), .B(n13259), .Z(n13263) );
  OR U13876 ( .A(n13264), .B(n13263), .Z(n13266) );
  XOR U13877 ( .A(n13262), .B(n13261), .Z(n13596) );
  XOR U13878 ( .A(n13264), .B(n13263), .Z(n13595) );
  NAND U13879 ( .A(n13596), .B(n13595), .Z(n13265) );
  NAND U13880 ( .A(n13266), .B(n13265), .Z(n13269) );
  XOR U13881 ( .A(n13268), .B(n13267), .Z(n13270) );
  NANDN U13882 ( .A(n13269), .B(n13270), .Z(n13272) );
  NAND U13883 ( .A(a[10]), .B(b[22]), .Z(n13654) );
  XNOR U13884 ( .A(n13270), .B(n13269), .Z(n13655) );
  NANDN U13885 ( .A(n13654), .B(n13655), .Z(n13271) );
  NAND U13886 ( .A(n13272), .B(n13271), .Z(n13273) );
  OR U13887 ( .A(n13274), .B(n13273), .Z(n13278) );
  XNOR U13888 ( .A(n13274), .B(n13273), .Z(n13658) );
  XOR U13889 ( .A(n13276), .B(n13275), .Z(n13659) );
  NANDN U13890 ( .A(n13658), .B(n13659), .Z(n13277) );
  NAND U13891 ( .A(n13278), .B(n13277), .Z(n13281) );
  XOR U13892 ( .A(n13280), .B(n13279), .Z(n13282) );
  NANDN U13893 ( .A(n13281), .B(n13282), .Z(n13284) );
  NAND U13894 ( .A(a[12]), .B(b[22]), .Z(n13666) );
  XNOR U13895 ( .A(n13282), .B(n13281), .Z(n13667) );
  NANDN U13896 ( .A(n13666), .B(n13667), .Z(n13283) );
  NAND U13897 ( .A(n13284), .B(n13283), .Z(n13285) );
  OR U13898 ( .A(n13286), .B(n13285), .Z(n13290) );
  XNOR U13899 ( .A(n13286), .B(n13285), .Z(n13670) );
  XOR U13900 ( .A(n13288), .B(n13287), .Z(n13671) );
  NANDN U13901 ( .A(n13670), .B(n13671), .Z(n13289) );
  NAND U13902 ( .A(n13290), .B(n13289), .Z(n13291) );
  OR U13903 ( .A(n13292), .B(n13291), .Z(n13294) );
  NAND U13904 ( .A(a[14]), .B(b[22]), .Z(n13678) );
  XOR U13905 ( .A(n13292), .B(n13291), .Z(n13679) );
  NANDN U13906 ( .A(n13678), .B(n13679), .Z(n13293) );
  NAND U13907 ( .A(n13294), .B(n13293), .Z(n13295) );
  OR U13908 ( .A(n13296), .B(n13295), .Z(n13300) );
  XNOR U13909 ( .A(n13296), .B(n13295), .Z(n13682) );
  XOR U13910 ( .A(n13298), .B(n13297), .Z(n13683) );
  NANDN U13911 ( .A(n13682), .B(n13683), .Z(n13299) );
  NAND U13912 ( .A(n13300), .B(n13299), .Z(n13303) );
  XOR U13913 ( .A(n13302), .B(n13301), .Z(n13304) );
  NANDN U13914 ( .A(n13303), .B(n13304), .Z(n13306) );
  NAND U13915 ( .A(a[16]), .B(b[22]), .Z(n13690) );
  XNOR U13916 ( .A(n13304), .B(n13303), .Z(n13691) );
  NANDN U13917 ( .A(n13690), .B(n13691), .Z(n13305) );
  NAND U13918 ( .A(n13306), .B(n13305), .Z(n13307) );
  OR U13919 ( .A(n13308), .B(n13307), .Z(n13312) );
  XNOR U13920 ( .A(n13308), .B(n13307), .Z(n13694) );
  XOR U13921 ( .A(n13310), .B(n13309), .Z(n13695) );
  NANDN U13922 ( .A(n13694), .B(n13695), .Z(n13311) );
  NAND U13923 ( .A(n13312), .B(n13311), .Z(n13313) );
  OR U13924 ( .A(n13314), .B(n13313), .Z(n13316) );
  NAND U13925 ( .A(a[18]), .B(b[22]), .Z(n13702) );
  XOR U13926 ( .A(n13314), .B(n13313), .Z(n13703) );
  NANDN U13927 ( .A(n13702), .B(n13703), .Z(n13315) );
  NAND U13928 ( .A(n13316), .B(n13315), .Z(n13319) );
  OR U13929 ( .A(n13320), .B(n13319), .Z(n13322) );
  XOR U13930 ( .A(n13318), .B(n13317), .Z(n13593) );
  XOR U13931 ( .A(n13320), .B(n13319), .Z(n13594) );
  NAND U13932 ( .A(n13593), .B(n13594), .Z(n13321) );
  NAND U13933 ( .A(n13322), .B(n13321), .Z(n13326) );
  XOR U13934 ( .A(n13324), .B(n13323), .Z(n13325) );
  NAND U13935 ( .A(n13326), .B(n13325), .Z(n13328) );
  ANDN U13936 ( .B(b[22]), .A(n176), .Z(n13711) );
  XNOR U13937 ( .A(n13326), .B(n13325), .Z(n13710) );
  OR U13938 ( .A(n13711), .B(n13710), .Z(n13327) );
  NAND U13939 ( .A(n13328), .B(n13327), .Z(n13329) );
  NANDN U13940 ( .A(n13330), .B(n13329), .Z(n13334) );
  XOR U13941 ( .A(n13332), .B(n13331), .Z(n13716) );
  NANDN U13942 ( .A(n13717), .B(n13716), .Z(n13333) );
  NAND U13943 ( .A(n13334), .B(n13333), .Z(n13337) );
  XOR U13944 ( .A(n13336), .B(n13335), .Z(n13338) );
  OR U13945 ( .A(n13337), .B(n13338), .Z(n13340) );
  NAND U13946 ( .A(a[22]), .B(b[22]), .Z(n13724) );
  XOR U13947 ( .A(n13338), .B(n13337), .Z(n13725) );
  NANDN U13948 ( .A(n13724), .B(n13725), .Z(n13339) );
  NAND U13949 ( .A(n13340), .B(n13339), .Z(n13341) );
  OR U13950 ( .A(n13342), .B(n13341), .Z(n13346) );
  XNOR U13951 ( .A(n13342), .B(n13341), .Z(n13728) );
  XOR U13952 ( .A(n13344), .B(n13343), .Z(n13729) );
  NANDN U13953 ( .A(n13728), .B(n13729), .Z(n13345) );
  NAND U13954 ( .A(n13346), .B(n13345), .Z(n13349) );
  XOR U13955 ( .A(n13348), .B(n13347), .Z(n13350) );
  OR U13956 ( .A(n13349), .B(n13350), .Z(n13352) );
  NAND U13957 ( .A(a[24]), .B(b[22]), .Z(n13736) );
  XOR U13958 ( .A(n13350), .B(n13349), .Z(n13737) );
  NANDN U13959 ( .A(n13736), .B(n13737), .Z(n13351) );
  NAND U13960 ( .A(n13352), .B(n13351), .Z(n13353) );
  OR U13961 ( .A(n13354), .B(n13353), .Z(n13358) );
  XNOR U13962 ( .A(n13354), .B(n13353), .Z(n13740) );
  XOR U13963 ( .A(n13356), .B(n13355), .Z(n13741) );
  NANDN U13964 ( .A(n13740), .B(n13741), .Z(n13357) );
  NAND U13965 ( .A(n13358), .B(n13357), .Z(n13361) );
  XOR U13966 ( .A(n13360), .B(n13359), .Z(n13362) );
  OR U13967 ( .A(n13361), .B(n13362), .Z(n13364) );
  NAND U13968 ( .A(a[26]), .B(b[22]), .Z(n13748) );
  XOR U13969 ( .A(n13362), .B(n13361), .Z(n13749) );
  NANDN U13970 ( .A(n13748), .B(n13749), .Z(n13363) );
  NAND U13971 ( .A(n13364), .B(n13363), .Z(n13365) );
  OR U13972 ( .A(n13366), .B(n13365), .Z(n13370) );
  XNOR U13973 ( .A(n13366), .B(n13365), .Z(n13752) );
  XOR U13974 ( .A(n13368), .B(n13367), .Z(n13753) );
  NANDN U13975 ( .A(n13752), .B(n13753), .Z(n13369) );
  NAND U13976 ( .A(n13370), .B(n13369), .Z(n13373) );
  XOR U13977 ( .A(n13372), .B(n13371), .Z(n13374) );
  OR U13978 ( .A(n13373), .B(n13374), .Z(n13376) );
  NAND U13979 ( .A(a[28]), .B(b[22]), .Z(n13760) );
  XOR U13980 ( .A(n13374), .B(n13373), .Z(n13761) );
  NANDN U13981 ( .A(n13760), .B(n13761), .Z(n13375) );
  NAND U13982 ( .A(n13376), .B(n13375), .Z(n13377) );
  OR U13983 ( .A(n13378), .B(n13377), .Z(n13382) );
  XNOR U13984 ( .A(n13378), .B(n13377), .Z(n13764) );
  XOR U13985 ( .A(n13380), .B(n13379), .Z(n13765) );
  NANDN U13986 ( .A(n13764), .B(n13765), .Z(n13381) );
  NAND U13987 ( .A(n13382), .B(n13381), .Z(n13385) );
  XOR U13988 ( .A(n13384), .B(n13383), .Z(n13386) );
  OR U13989 ( .A(n13385), .B(n13386), .Z(n13388) );
  NAND U13990 ( .A(a[30]), .B(b[22]), .Z(n13772) );
  XOR U13991 ( .A(n13386), .B(n13385), .Z(n13773) );
  NANDN U13992 ( .A(n13772), .B(n13773), .Z(n13387) );
  NAND U13993 ( .A(n13388), .B(n13387), .Z(n13389) );
  OR U13994 ( .A(n13390), .B(n13389), .Z(n13394) );
  XNOR U13995 ( .A(n13390), .B(n13389), .Z(n13776) );
  XOR U13996 ( .A(n13392), .B(n13391), .Z(n13777) );
  NANDN U13997 ( .A(n13776), .B(n13777), .Z(n13393) );
  NAND U13998 ( .A(n13394), .B(n13393), .Z(n13397) );
  XOR U13999 ( .A(n13396), .B(n13395), .Z(n13398) );
  OR U14000 ( .A(n13397), .B(n13398), .Z(n13400) );
  NAND U14001 ( .A(a[32]), .B(b[22]), .Z(n13784) );
  XOR U14002 ( .A(n13398), .B(n13397), .Z(n13785) );
  NANDN U14003 ( .A(n13784), .B(n13785), .Z(n13399) );
  NAND U14004 ( .A(n13400), .B(n13399), .Z(n13401) );
  OR U14005 ( .A(n13402), .B(n13401), .Z(n13406) );
  XNOR U14006 ( .A(n13402), .B(n13401), .Z(n13788) );
  XOR U14007 ( .A(n13404), .B(n13403), .Z(n13789) );
  NANDN U14008 ( .A(n13788), .B(n13789), .Z(n13405) );
  NAND U14009 ( .A(n13406), .B(n13405), .Z(n13409) );
  XOR U14010 ( .A(n13408), .B(n13407), .Z(n13410) );
  OR U14011 ( .A(n13409), .B(n13410), .Z(n13412) );
  NAND U14012 ( .A(a[34]), .B(b[22]), .Z(n13796) );
  XOR U14013 ( .A(n13410), .B(n13409), .Z(n13797) );
  NANDN U14014 ( .A(n13796), .B(n13797), .Z(n13411) );
  NAND U14015 ( .A(n13412), .B(n13411), .Z(n13413) );
  OR U14016 ( .A(n13414), .B(n13413), .Z(n13418) );
  XNOR U14017 ( .A(n13414), .B(n13413), .Z(n13800) );
  XOR U14018 ( .A(n13416), .B(n13415), .Z(n13801) );
  NANDN U14019 ( .A(n13800), .B(n13801), .Z(n13417) );
  NAND U14020 ( .A(n13418), .B(n13417), .Z(n13421) );
  XOR U14021 ( .A(n13420), .B(n13419), .Z(n13422) );
  OR U14022 ( .A(n13421), .B(n13422), .Z(n13424) );
  NAND U14023 ( .A(a[36]), .B(b[22]), .Z(n13808) );
  XOR U14024 ( .A(n13422), .B(n13421), .Z(n13809) );
  NANDN U14025 ( .A(n13808), .B(n13809), .Z(n13423) );
  NAND U14026 ( .A(n13424), .B(n13423), .Z(n13425) );
  OR U14027 ( .A(n13426), .B(n13425), .Z(n13430) );
  XNOR U14028 ( .A(n13426), .B(n13425), .Z(n13812) );
  XOR U14029 ( .A(n13428), .B(n13427), .Z(n13813) );
  NANDN U14030 ( .A(n13812), .B(n13813), .Z(n13429) );
  NAND U14031 ( .A(n13430), .B(n13429), .Z(n13433) );
  XNOR U14032 ( .A(n13432), .B(n13431), .Z(n13434) );
  OR U14033 ( .A(n13433), .B(n13434), .Z(n13436) );
  NAND U14034 ( .A(a[38]), .B(b[22]), .Z(n13820) );
  XOR U14035 ( .A(n13434), .B(n13433), .Z(n13821) );
  NANDN U14036 ( .A(n13820), .B(n13821), .Z(n13435) );
  NAND U14037 ( .A(n13436), .B(n13435), .Z(n13437) );
  OR U14038 ( .A(n13438), .B(n13437), .Z(n13442) );
  XNOR U14039 ( .A(n13438), .B(n13437), .Z(n13824) );
  XOR U14040 ( .A(n13440), .B(n13439), .Z(n13825) );
  NANDN U14041 ( .A(n13824), .B(n13825), .Z(n13441) );
  NAND U14042 ( .A(n13442), .B(n13441), .Z(n13445) );
  XOR U14043 ( .A(n13444), .B(n13443), .Z(n13446) );
  OR U14044 ( .A(n13445), .B(n13446), .Z(n13448) );
  NAND U14045 ( .A(a[40]), .B(b[22]), .Z(n13831) );
  XOR U14046 ( .A(n13446), .B(n13445), .Z(n13830) );
  NANDN U14047 ( .A(n13831), .B(n13830), .Z(n13447) );
  NAND U14048 ( .A(n13448), .B(n13447), .Z(n13451) );
  ANDN U14049 ( .B(b[22]), .A(n189), .Z(n13452) );
  OR U14050 ( .A(n13451), .B(n13452), .Z(n13454) );
  XOR U14051 ( .A(n13450), .B(n13449), .Z(n13837) );
  XOR U14052 ( .A(n13452), .B(n13451), .Z(n13836) );
  NANDN U14053 ( .A(n13837), .B(n13836), .Z(n13453) );
  NAND U14054 ( .A(n13454), .B(n13453), .Z(n13458) );
  AND U14055 ( .A(b[22]), .B(a[42]), .Z(n13457) );
  NANDN U14056 ( .A(n13458), .B(n13457), .Z(n13460) );
  XNOR U14057 ( .A(n13458), .B(n13457), .Z(n13844) );
  NANDN U14058 ( .A(n13845), .B(n13844), .Z(n13459) );
  NAND U14059 ( .A(n13460), .B(n13459), .Z(n13464) );
  XOR U14060 ( .A(n13462), .B(n13461), .Z(n13463) );
  NAND U14061 ( .A(n13464), .B(n13463), .Z(n13466) );
  XNOR U14062 ( .A(n13464), .B(n13463), .Z(n13849) );
  NAND U14063 ( .A(a[43]), .B(b[22]), .Z(n13848) );
  OR U14064 ( .A(n13849), .B(n13848), .Z(n13465) );
  NAND U14065 ( .A(n13466), .B(n13465), .Z(n13470) );
  NANDN U14066 ( .A(n13469), .B(n13470), .Z(n13472) );
  XOR U14067 ( .A(n13468), .B(n13467), .Z(n13854) );
  XNOR U14068 ( .A(n13470), .B(n13469), .Z(n13855) );
  NAND U14069 ( .A(n13854), .B(n13855), .Z(n13471) );
  NAND U14070 ( .A(n13472), .B(n13471), .Z(n13475) );
  AND U14071 ( .A(b[22]), .B(a[45]), .Z(n13476) );
  OR U14072 ( .A(n13475), .B(n13476), .Z(n13478) );
  XNOR U14073 ( .A(n13474), .B(n13473), .Z(n13861) );
  XOR U14074 ( .A(n13476), .B(n13475), .Z(n13860) );
  NANDN U14075 ( .A(n13861), .B(n13860), .Z(n13477) );
  NAND U14076 ( .A(n13478), .B(n13477), .Z(n13482) );
  NAND U14077 ( .A(a[46]), .B(b[22]), .Z(n13481) );
  OR U14078 ( .A(n13482), .B(n13481), .Z(n13484) );
  XOR U14079 ( .A(n13480), .B(n13479), .Z(n13866) );
  XOR U14080 ( .A(n13482), .B(n13481), .Z(n13867) );
  NAND U14081 ( .A(n13866), .B(n13867), .Z(n13483) );
  NAND U14082 ( .A(n13484), .B(n13483), .Z(n13487) );
  AND U14083 ( .A(b[22]), .B(a[47]), .Z(n13488) );
  OR U14084 ( .A(n13487), .B(n13488), .Z(n13490) );
  XNOR U14085 ( .A(n13486), .B(n13485), .Z(n13873) );
  XOR U14086 ( .A(n13488), .B(n13487), .Z(n13872) );
  NANDN U14087 ( .A(n13873), .B(n13872), .Z(n13489) );
  NAND U14088 ( .A(n13490), .B(n13489), .Z(n13494) );
  NAND U14089 ( .A(a[48]), .B(b[22]), .Z(n13493) );
  OR U14090 ( .A(n13494), .B(n13493), .Z(n13496) );
  XOR U14091 ( .A(n13492), .B(n13491), .Z(n13878) );
  XOR U14092 ( .A(n13494), .B(n13493), .Z(n13879) );
  NAND U14093 ( .A(n13878), .B(n13879), .Z(n13495) );
  NAND U14094 ( .A(n13496), .B(n13495), .Z(n13499) );
  AND U14095 ( .A(b[22]), .B(a[49]), .Z(n13500) );
  OR U14096 ( .A(n13499), .B(n13500), .Z(n13502) );
  XNOR U14097 ( .A(n13498), .B(n13497), .Z(n13885) );
  XOR U14098 ( .A(n13500), .B(n13499), .Z(n13884) );
  NANDN U14099 ( .A(n13885), .B(n13884), .Z(n13501) );
  NAND U14100 ( .A(n13502), .B(n13501), .Z(n13506) );
  NAND U14101 ( .A(a[50]), .B(b[22]), .Z(n13505) );
  OR U14102 ( .A(n13506), .B(n13505), .Z(n13508) );
  XOR U14103 ( .A(n13504), .B(n13503), .Z(n13890) );
  XOR U14104 ( .A(n13506), .B(n13505), .Z(n13891) );
  NAND U14105 ( .A(n13890), .B(n13891), .Z(n13507) );
  NAND U14106 ( .A(n13508), .B(n13507), .Z(n13511) );
  AND U14107 ( .A(b[22]), .B(a[51]), .Z(n13512) );
  OR U14108 ( .A(n13511), .B(n13512), .Z(n13514) );
  XNOR U14109 ( .A(n13510), .B(n13509), .Z(n13897) );
  XOR U14110 ( .A(n13512), .B(n13511), .Z(n13896) );
  NANDN U14111 ( .A(n13897), .B(n13896), .Z(n13513) );
  NAND U14112 ( .A(n13514), .B(n13513), .Z(n13518) );
  NAND U14113 ( .A(a[52]), .B(b[22]), .Z(n13517) );
  OR U14114 ( .A(n13518), .B(n13517), .Z(n13520) );
  XOR U14115 ( .A(n13516), .B(n13515), .Z(n13902) );
  XOR U14116 ( .A(n13518), .B(n13517), .Z(n13903) );
  NAND U14117 ( .A(n13902), .B(n13903), .Z(n13519) );
  NAND U14118 ( .A(n13520), .B(n13519), .Z(n13523) );
  AND U14119 ( .A(b[22]), .B(a[53]), .Z(n13524) );
  OR U14120 ( .A(n13523), .B(n13524), .Z(n13526) );
  XNOR U14121 ( .A(n13522), .B(n13521), .Z(n13909) );
  XOR U14122 ( .A(n13524), .B(n13523), .Z(n13908) );
  NANDN U14123 ( .A(n13909), .B(n13908), .Z(n13525) );
  NAND U14124 ( .A(n13526), .B(n13525), .Z(n13530) );
  NAND U14125 ( .A(a[54]), .B(b[22]), .Z(n13529) );
  OR U14126 ( .A(n13530), .B(n13529), .Z(n13532) );
  XOR U14127 ( .A(n13528), .B(n13527), .Z(n13914) );
  XOR U14128 ( .A(n13530), .B(n13529), .Z(n13915) );
  NAND U14129 ( .A(n13914), .B(n13915), .Z(n13531) );
  NAND U14130 ( .A(n13532), .B(n13531), .Z(n13535) );
  AND U14131 ( .A(b[22]), .B(a[55]), .Z(n13536) );
  OR U14132 ( .A(n13535), .B(n13536), .Z(n13538) );
  XNOR U14133 ( .A(n13534), .B(n13533), .Z(n13921) );
  XOR U14134 ( .A(n13536), .B(n13535), .Z(n13920) );
  NANDN U14135 ( .A(n13921), .B(n13920), .Z(n13537) );
  NAND U14136 ( .A(n13538), .B(n13537), .Z(n13542) );
  NAND U14137 ( .A(a[56]), .B(b[22]), .Z(n13541) );
  OR U14138 ( .A(n13542), .B(n13541), .Z(n13544) );
  XOR U14139 ( .A(n13540), .B(n13539), .Z(n13926) );
  XOR U14140 ( .A(n13542), .B(n13541), .Z(n13927) );
  NAND U14141 ( .A(n13926), .B(n13927), .Z(n13543) );
  NAND U14142 ( .A(n13544), .B(n13543), .Z(n13547) );
  AND U14143 ( .A(b[22]), .B(a[57]), .Z(n13548) );
  OR U14144 ( .A(n13547), .B(n13548), .Z(n13550) );
  XNOR U14145 ( .A(n13546), .B(n13545), .Z(n13931) );
  XOR U14146 ( .A(n13548), .B(n13547), .Z(n13930) );
  NANDN U14147 ( .A(n13931), .B(n13930), .Z(n13549) );
  NAND U14148 ( .A(n13550), .B(n13549), .Z(n13554) );
  NAND U14149 ( .A(a[58]), .B(b[22]), .Z(n13553) );
  OR U14150 ( .A(n13554), .B(n13553), .Z(n13556) );
  XOR U14151 ( .A(n13552), .B(n13551), .Z(n13936) );
  XOR U14152 ( .A(n13554), .B(n13553), .Z(n13937) );
  NAND U14153 ( .A(n13936), .B(n13937), .Z(n13555) );
  NAND U14154 ( .A(n13556), .B(n13555), .Z(n13559) );
  AND U14155 ( .A(b[22]), .B(a[59]), .Z(n13560) );
  OR U14156 ( .A(n13559), .B(n13560), .Z(n13562) );
  XNOR U14157 ( .A(n13558), .B(n13557), .Z(n13943) );
  XOR U14158 ( .A(n13560), .B(n13559), .Z(n13942) );
  NANDN U14159 ( .A(n13943), .B(n13942), .Z(n13561) );
  NAND U14160 ( .A(n13562), .B(n13561), .Z(n13566) );
  NAND U14161 ( .A(a[60]), .B(b[22]), .Z(n13565) );
  OR U14162 ( .A(n13566), .B(n13565), .Z(n13568) );
  XOR U14163 ( .A(n13564), .B(n13563), .Z(n13589) );
  XOR U14164 ( .A(n13566), .B(n13565), .Z(n13590) );
  NAND U14165 ( .A(n13589), .B(n13590), .Z(n13567) );
  NAND U14166 ( .A(n13568), .B(n13567), .Z(n13571) );
  AND U14167 ( .A(b[22]), .B(a[61]), .Z(n13572) );
  OR U14168 ( .A(n13571), .B(n13572), .Z(n13574) );
  XNOR U14169 ( .A(n13570), .B(n13569), .Z(n13951) );
  XOR U14170 ( .A(n13572), .B(n13571), .Z(n13950) );
  NANDN U14171 ( .A(n13951), .B(n13950), .Z(n13573) );
  NAND U14172 ( .A(n13574), .B(n13573), .Z(n13578) );
  NAND U14173 ( .A(a[62]), .B(b[22]), .Z(n13577) );
  OR U14174 ( .A(n13578), .B(n13577), .Z(n13580) );
  XOR U14175 ( .A(n13576), .B(n13575), .Z(n13957) );
  XOR U14176 ( .A(n13578), .B(n13577), .Z(n13956) );
  NAND U14177 ( .A(n13957), .B(n13956), .Z(n13579) );
  NAND U14178 ( .A(n13580), .B(n13579), .Z(n13583) );
  AND U14179 ( .A(b[22]), .B(a[63]), .Z(n13584) );
  OR U14180 ( .A(n13583), .B(n13584), .Z(n13586) );
  XNOR U14181 ( .A(n13582), .B(n13581), .Z(n13963) );
  XOR U14182 ( .A(n13584), .B(n13583), .Z(n13962) );
  NANDN U14183 ( .A(n13963), .B(n13962), .Z(n13585) );
  NAND U14184 ( .A(n13586), .B(n13585), .Z(n13587) );
  NOR U14185 ( .A(n13588), .B(n13587), .Z(n21969) );
  XOR U14186 ( .A(n13588), .B(n13587), .Z(n13964) );
  NAND U14187 ( .A(a[62]), .B(b[21]), .Z(n13952) );
  NAND U14188 ( .A(a[61]), .B(b[21]), .Z(n13592) );
  XOR U14189 ( .A(n13590), .B(n13589), .Z(n13591) );
  NANDN U14190 ( .A(n13592), .B(n13591), .Z(n13949) );
  XOR U14191 ( .A(n13592), .B(n13591), .Z(n14331) );
  NAND U14192 ( .A(a[60]), .B(b[21]), .Z(n13944) );
  NAND U14193 ( .A(a[56]), .B(b[21]), .Z(n13922) );
  NAND U14194 ( .A(a[54]), .B(b[21]), .Z(n13910) );
  NAND U14195 ( .A(a[52]), .B(b[21]), .Z(n13898) );
  NAND U14196 ( .A(a[50]), .B(b[21]), .Z(n13886) );
  NAND U14197 ( .A(a[48]), .B(b[21]), .Z(n13874) );
  NAND U14198 ( .A(a[46]), .B(b[21]), .Z(n13862) );
  ANDN U14199 ( .B(b[21]), .A(n187), .Z(n13819) );
  ANDN U14200 ( .B(b[21]), .A(n21772), .Z(n13807) );
  ANDN U14201 ( .B(b[21]), .A(n184), .Z(n13795) );
  ANDN U14202 ( .B(b[21]), .A(n21751), .Z(n13783) );
  ANDN U14203 ( .B(b[21]), .A(n21740), .Z(n13771) );
  ANDN U14204 ( .B(b[21]), .A(n21727), .Z(n13759) );
  ANDN U14205 ( .B(b[21]), .A(n21716), .Z(n13747) );
  ANDN U14206 ( .B(b[21]), .A(n21703), .Z(n13735) );
  ANDN U14207 ( .B(b[21]), .A(n21692), .Z(n13723) );
  ANDN U14208 ( .B(b[21]), .A(n21681), .Z(n13713) );
  ANDN U14209 ( .B(b[21]), .A(n21670), .Z(n13701) );
  ANDN U14210 ( .B(b[21]), .A(n174), .Z(n13689) );
  ANDN U14211 ( .B(b[21]), .A(n172), .Z(n13677) );
  ANDN U14212 ( .B(b[21]), .A(n170), .Z(n13665) );
  NAND U14213 ( .A(a[11]), .B(b[21]), .Z(n13653) );
  XNOR U14214 ( .A(n13596), .B(n13595), .Z(n13649) );
  ANDN U14215 ( .B(b[21]), .A(n21615), .Z(n13645) );
  ANDN U14216 ( .B(b[21]), .A(n166), .Z(n13633) );
  ANDN U14217 ( .B(b[21]), .A(n164), .Z(n13619) );
  ANDN U14218 ( .B(b[21]), .A(n21580), .Z(n13606) );
  NAND U14219 ( .A(b[22]), .B(a[1]), .Z(n13599) );
  AND U14220 ( .A(b[21]), .B(a[0]), .Z(n14357) );
  NANDN U14221 ( .A(n13599), .B(n14357), .Z(n13598) );
  NAND U14222 ( .A(a[2]), .B(b[21]), .Z(n13597) );
  AND U14223 ( .A(n13598), .B(n13597), .Z(n13605) );
  NANDN U14224 ( .A(n13599), .B(a[0]), .Z(n13600) );
  XNOR U14225 ( .A(a[2]), .B(n13600), .Z(n13601) );
  NAND U14226 ( .A(b[21]), .B(n13601), .Z(n13990) );
  AND U14227 ( .A(a[1]), .B(b[22]), .Z(n13602) );
  XNOR U14228 ( .A(n13603), .B(n13602), .Z(n13989) );
  NANDN U14229 ( .A(n13990), .B(n13989), .Z(n13604) );
  NANDN U14230 ( .A(n13605), .B(n13604), .Z(n13607) );
  NANDN U14231 ( .A(n13606), .B(n13607), .Z(n13611) );
  XOR U14232 ( .A(n13607), .B(n13606), .Z(n13994) );
  NANDN U14233 ( .A(n13994), .B(n13993), .Z(n13610) );
  NAND U14234 ( .A(n13611), .B(n13610), .Z(n13615) );
  XOR U14235 ( .A(n13613), .B(n13612), .Z(n13614) );
  NANDN U14236 ( .A(n13615), .B(n13614), .Z(n13617) );
  NAND U14237 ( .A(a[4]), .B(b[21]), .Z(n14001) );
  NANDN U14238 ( .A(n14001), .B(n14002), .Z(n13616) );
  NAND U14239 ( .A(n13617), .B(n13616), .Z(n13618) );
  OR U14240 ( .A(n13619), .B(n13618), .Z(n13623) );
  XNOR U14241 ( .A(n13619), .B(n13618), .Z(n13976) );
  XOR U14242 ( .A(n13621), .B(n13620), .Z(n13977) );
  NANDN U14243 ( .A(n13976), .B(n13977), .Z(n13622) );
  NAND U14244 ( .A(n13623), .B(n13622), .Z(n13626) );
  XOR U14245 ( .A(n13625), .B(n13624), .Z(n13627) );
  NANDN U14246 ( .A(n13626), .B(n13627), .Z(n13629) );
  NAND U14247 ( .A(a[6]), .B(b[21]), .Z(n14011) );
  XNOR U14248 ( .A(n13627), .B(n13626), .Z(n14012) );
  NANDN U14249 ( .A(n14011), .B(n14012), .Z(n13628) );
  NAND U14250 ( .A(n13629), .B(n13628), .Z(n13632) );
  OR U14251 ( .A(n13633), .B(n13632), .Z(n13635) );
  XOR U14252 ( .A(n13631), .B(n13630), .Z(n14015) );
  XOR U14253 ( .A(n13633), .B(n13632), .Z(n14016) );
  NANDN U14254 ( .A(n14015), .B(n14016), .Z(n13634) );
  NAND U14255 ( .A(n13635), .B(n13634), .Z(n13639) );
  XNOR U14256 ( .A(n13637), .B(n13636), .Z(n13638) );
  NANDN U14257 ( .A(n13639), .B(n13638), .Z(n13641) );
  NAND U14258 ( .A(a[8]), .B(b[21]), .Z(n14023) );
  NANDN U14259 ( .A(n14023), .B(n14024), .Z(n13640) );
  NAND U14260 ( .A(n13641), .B(n13640), .Z(n13644) );
  OR U14261 ( .A(n13645), .B(n13644), .Z(n13647) );
  XOR U14262 ( .A(n13643), .B(n13642), .Z(n13975) );
  XOR U14263 ( .A(n13645), .B(n13644), .Z(n13974) );
  NAND U14264 ( .A(n13975), .B(n13974), .Z(n13646) );
  NAND U14265 ( .A(n13647), .B(n13646), .Z(n13648) );
  NANDN U14266 ( .A(n13649), .B(n13648), .Z(n13651) );
  ANDN U14267 ( .B(b[21]), .A(n168), .Z(n14034) );
  NANDN U14268 ( .A(n14034), .B(n14033), .Z(n13650) );
  AND U14269 ( .A(n13651), .B(n13650), .Z(n13652) );
  NANDN U14270 ( .A(n13653), .B(n13652), .Z(n13657) );
  XNOR U14271 ( .A(n13655), .B(n13654), .Z(n13973) );
  NAND U14272 ( .A(n13972), .B(n13973), .Z(n13656) );
  AND U14273 ( .A(n13657), .B(n13656), .Z(n13660) );
  XOR U14274 ( .A(n13659), .B(n13658), .Z(n13661) );
  NANDN U14275 ( .A(n13660), .B(n13661), .Z(n13663) );
  NAND U14276 ( .A(a[12]), .B(b[21]), .Z(n14043) );
  XNOR U14277 ( .A(n13661), .B(n13660), .Z(n14044) );
  NANDN U14278 ( .A(n14043), .B(n14044), .Z(n13662) );
  NAND U14279 ( .A(n13663), .B(n13662), .Z(n13664) );
  OR U14280 ( .A(n13665), .B(n13664), .Z(n13669) );
  XNOR U14281 ( .A(n13665), .B(n13664), .Z(n14047) );
  XOR U14282 ( .A(n13667), .B(n13666), .Z(n14048) );
  NANDN U14283 ( .A(n14047), .B(n14048), .Z(n13668) );
  NAND U14284 ( .A(n13669), .B(n13668), .Z(n13672) );
  XOR U14285 ( .A(n13671), .B(n13670), .Z(n13673) );
  NANDN U14286 ( .A(n13672), .B(n13673), .Z(n13675) );
  NAND U14287 ( .A(a[14]), .B(b[21]), .Z(n14055) );
  XNOR U14288 ( .A(n13673), .B(n13672), .Z(n14056) );
  NANDN U14289 ( .A(n14055), .B(n14056), .Z(n13674) );
  NAND U14290 ( .A(n13675), .B(n13674), .Z(n13676) );
  OR U14291 ( .A(n13677), .B(n13676), .Z(n13681) );
  XNOR U14292 ( .A(n13677), .B(n13676), .Z(n14059) );
  XOR U14293 ( .A(n13679), .B(n13678), .Z(n14060) );
  NANDN U14294 ( .A(n14059), .B(n14060), .Z(n13680) );
  NAND U14295 ( .A(n13681), .B(n13680), .Z(n13684) );
  XOR U14296 ( .A(n13683), .B(n13682), .Z(n13685) );
  NANDN U14297 ( .A(n13684), .B(n13685), .Z(n13687) );
  NAND U14298 ( .A(a[16]), .B(b[21]), .Z(n14067) );
  XNOR U14299 ( .A(n13685), .B(n13684), .Z(n14068) );
  NANDN U14300 ( .A(n14067), .B(n14068), .Z(n13686) );
  NAND U14301 ( .A(n13687), .B(n13686), .Z(n13688) );
  OR U14302 ( .A(n13689), .B(n13688), .Z(n13693) );
  XNOR U14303 ( .A(n13689), .B(n13688), .Z(n14071) );
  XOR U14304 ( .A(n13691), .B(n13690), .Z(n14072) );
  NANDN U14305 ( .A(n14071), .B(n14072), .Z(n13692) );
  NAND U14306 ( .A(n13693), .B(n13692), .Z(n13696) );
  XOR U14307 ( .A(n13695), .B(n13694), .Z(n13697) );
  NANDN U14308 ( .A(n13696), .B(n13697), .Z(n13699) );
  NAND U14309 ( .A(a[18]), .B(b[21]), .Z(n14079) );
  XNOR U14310 ( .A(n13697), .B(n13696), .Z(n14080) );
  NANDN U14311 ( .A(n14079), .B(n14080), .Z(n13698) );
  NAND U14312 ( .A(n13699), .B(n13698), .Z(n13700) );
  OR U14313 ( .A(n13701), .B(n13700), .Z(n13705) );
  XNOR U14314 ( .A(n13701), .B(n13700), .Z(n14083) );
  XOR U14315 ( .A(n13703), .B(n13702), .Z(n14084) );
  NANDN U14316 ( .A(n14083), .B(n14084), .Z(n13704) );
  NAND U14317 ( .A(n13705), .B(n13704), .Z(n13706) );
  OR U14318 ( .A(n13707), .B(n13706), .Z(n13709) );
  NAND U14319 ( .A(a[20]), .B(b[21]), .Z(n14091) );
  XOR U14320 ( .A(n13707), .B(n13706), .Z(n14092) );
  NANDN U14321 ( .A(n14091), .B(n14092), .Z(n13708) );
  NAND U14322 ( .A(n13709), .B(n13708), .Z(n13712) );
  OR U14323 ( .A(n13713), .B(n13712), .Z(n13715) );
  XOR U14324 ( .A(n13711), .B(n13710), .Z(n13970) );
  XOR U14325 ( .A(n13713), .B(n13712), .Z(n13971) );
  NAND U14326 ( .A(n13970), .B(n13971), .Z(n13714) );
  NAND U14327 ( .A(n13715), .B(n13714), .Z(n13718) );
  NANDN U14328 ( .A(n13718), .B(n13719), .Z(n13721) );
  NAND U14329 ( .A(a[22]), .B(b[21]), .Z(n14101) );
  XNOR U14330 ( .A(n13719), .B(n13718), .Z(n14102) );
  NANDN U14331 ( .A(n14101), .B(n14102), .Z(n13720) );
  NAND U14332 ( .A(n13721), .B(n13720), .Z(n13722) );
  OR U14333 ( .A(n13723), .B(n13722), .Z(n13727) );
  XNOR U14334 ( .A(n13723), .B(n13722), .Z(n14105) );
  XOR U14335 ( .A(n13725), .B(n13724), .Z(n14106) );
  NANDN U14336 ( .A(n14105), .B(n14106), .Z(n13726) );
  NAND U14337 ( .A(n13727), .B(n13726), .Z(n13730) );
  XOR U14338 ( .A(n13729), .B(n13728), .Z(n13731) );
  NANDN U14339 ( .A(n13730), .B(n13731), .Z(n13733) );
  NAND U14340 ( .A(a[24]), .B(b[21]), .Z(n14113) );
  XNOR U14341 ( .A(n13731), .B(n13730), .Z(n14114) );
  NANDN U14342 ( .A(n14113), .B(n14114), .Z(n13732) );
  NAND U14343 ( .A(n13733), .B(n13732), .Z(n13734) );
  OR U14344 ( .A(n13735), .B(n13734), .Z(n13739) );
  XNOR U14345 ( .A(n13735), .B(n13734), .Z(n14117) );
  XOR U14346 ( .A(n13737), .B(n13736), .Z(n14118) );
  NANDN U14347 ( .A(n14117), .B(n14118), .Z(n13738) );
  NAND U14348 ( .A(n13739), .B(n13738), .Z(n13742) );
  XOR U14349 ( .A(n13741), .B(n13740), .Z(n13743) );
  NANDN U14350 ( .A(n13742), .B(n13743), .Z(n13745) );
  NAND U14351 ( .A(a[26]), .B(b[21]), .Z(n14125) );
  XNOR U14352 ( .A(n13743), .B(n13742), .Z(n14126) );
  NANDN U14353 ( .A(n14125), .B(n14126), .Z(n13744) );
  NAND U14354 ( .A(n13745), .B(n13744), .Z(n13746) );
  OR U14355 ( .A(n13747), .B(n13746), .Z(n13751) );
  XNOR U14356 ( .A(n13747), .B(n13746), .Z(n14129) );
  XOR U14357 ( .A(n13749), .B(n13748), .Z(n14130) );
  NANDN U14358 ( .A(n14129), .B(n14130), .Z(n13750) );
  NAND U14359 ( .A(n13751), .B(n13750), .Z(n13754) );
  XOR U14360 ( .A(n13753), .B(n13752), .Z(n13755) );
  NANDN U14361 ( .A(n13754), .B(n13755), .Z(n13757) );
  NAND U14362 ( .A(a[28]), .B(b[21]), .Z(n14137) );
  XNOR U14363 ( .A(n13755), .B(n13754), .Z(n14138) );
  NANDN U14364 ( .A(n14137), .B(n14138), .Z(n13756) );
  NAND U14365 ( .A(n13757), .B(n13756), .Z(n13758) );
  OR U14366 ( .A(n13759), .B(n13758), .Z(n13763) );
  XNOR U14367 ( .A(n13759), .B(n13758), .Z(n14141) );
  XOR U14368 ( .A(n13761), .B(n13760), .Z(n14142) );
  NANDN U14369 ( .A(n14141), .B(n14142), .Z(n13762) );
  NAND U14370 ( .A(n13763), .B(n13762), .Z(n13766) );
  XOR U14371 ( .A(n13765), .B(n13764), .Z(n13767) );
  NANDN U14372 ( .A(n13766), .B(n13767), .Z(n13769) );
  NAND U14373 ( .A(a[30]), .B(b[21]), .Z(n14149) );
  XNOR U14374 ( .A(n13767), .B(n13766), .Z(n14150) );
  NANDN U14375 ( .A(n14149), .B(n14150), .Z(n13768) );
  NAND U14376 ( .A(n13769), .B(n13768), .Z(n13770) );
  OR U14377 ( .A(n13771), .B(n13770), .Z(n13775) );
  XNOR U14378 ( .A(n13771), .B(n13770), .Z(n14153) );
  XOR U14379 ( .A(n13773), .B(n13772), .Z(n14154) );
  NANDN U14380 ( .A(n14153), .B(n14154), .Z(n13774) );
  NAND U14381 ( .A(n13775), .B(n13774), .Z(n13778) );
  XOR U14382 ( .A(n13777), .B(n13776), .Z(n13779) );
  NANDN U14383 ( .A(n13778), .B(n13779), .Z(n13781) );
  NAND U14384 ( .A(a[32]), .B(b[21]), .Z(n14161) );
  XNOR U14385 ( .A(n13779), .B(n13778), .Z(n14162) );
  NANDN U14386 ( .A(n14161), .B(n14162), .Z(n13780) );
  NAND U14387 ( .A(n13781), .B(n13780), .Z(n13782) );
  OR U14388 ( .A(n13783), .B(n13782), .Z(n13787) );
  XNOR U14389 ( .A(n13783), .B(n13782), .Z(n14165) );
  XOR U14390 ( .A(n13785), .B(n13784), .Z(n14166) );
  NANDN U14391 ( .A(n14165), .B(n14166), .Z(n13786) );
  NAND U14392 ( .A(n13787), .B(n13786), .Z(n13790) );
  XOR U14393 ( .A(n13789), .B(n13788), .Z(n13791) );
  NANDN U14394 ( .A(n13790), .B(n13791), .Z(n13793) );
  NAND U14395 ( .A(a[34]), .B(b[21]), .Z(n14173) );
  XNOR U14396 ( .A(n13791), .B(n13790), .Z(n14174) );
  NANDN U14397 ( .A(n14173), .B(n14174), .Z(n13792) );
  NAND U14398 ( .A(n13793), .B(n13792), .Z(n13794) );
  OR U14399 ( .A(n13795), .B(n13794), .Z(n13799) );
  XNOR U14400 ( .A(n13795), .B(n13794), .Z(n14177) );
  XOR U14401 ( .A(n13797), .B(n13796), .Z(n14178) );
  NANDN U14402 ( .A(n14177), .B(n14178), .Z(n13798) );
  NAND U14403 ( .A(n13799), .B(n13798), .Z(n13802) );
  XOR U14404 ( .A(n13801), .B(n13800), .Z(n13803) );
  NANDN U14405 ( .A(n13802), .B(n13803), .Z(n13805) );
  NAND U14406 ( .A(a[36]), .B(b[21]), .Z(n14185) );
  XNOR U14407 ( .A(n13803), .B(n13802), .Z(n14186) );
  NANDN U14408 ( .A(n14185), .B(n14186), .Z(n13804) );
  NAND U14409 ( .A(n13805), .B(n13804), .Z(n13806) );
  OR U14410 ( .A(n13807), .B(n13806), .Z(n13811) );
  XNOR U14411 ( .A(n13807), .B(n13806), .Z(n14189) );
  XOR U14412 ( .A(n13809), .B(n13808), .Z(n14190) );
  NANDN U14413 ( .A(n14189), .B(n14190), .Z(n13810) );
  NAND U14414 ( .A(n13811), .B(n13810), .Z(n13814) );
  XOR U14415 ( .A(n13813), .B(n13812), .Z(n13815) );
  NANDN U14416 ( .A(n13814), .B(n13815), .Z(n13817) );
  NAND U14417 ( .A(a[38]), .B(b[21]), .Z(n14197) );
  XNOR U14418 ( .A(n13815), .B(n13814), .Z(n14198) );
  NANDN U14419 ( .A(n14197), .B(n14198), .Z(n13816) );
  NAND U14420 ( .A(n13817), .B(n13816), .Z(n13818) );
  OR U14421 ( .A(n13819), .B(n13818), .Z(n13823) );
  XNOR U14422 ( .A(n13819), .B(n13818), .Z(n14201) );
  XOR U14423 ( .A(n13821), .B(n13820), .Z(n14202) );
  NANDN U14424 ( .A(n14201), .B(n14202), .Z(n13822) );
  NAND U14425 ( .A(n13823), .B(n13822), .Z(n13826) );
  XOR U14426 ( .A(n13825), .B(n13824), .Z(n13827) );
  NANDN U14427 ( .A(n13826), .B(n13827), .Z(n13829) );
  NAND U14428 ( .A(a[40]), .B(b[21]), .Z(n14209) );
  XNOR U14429 ( .A(n13827), .B(n13826), .Z(n14210) );
  NANDN U14430 ( .A(n14209), .B(n14210), .Z(n13828) );
  NAND U14431 ( .A(n13829), .B(n13828), .Z(n13832) );
  ANDN U14432 ( .B(b[21]), .A(n189), .Z(n13833) );
  OR U14433 ( .A(n13832), .B(n13833), .Z(n13835) );
  XOR U14434 ( .A(n13833), .B(n13832), .Z(n14213) );
  NANDN U14435 ( .A(n14214), .B(n14213), .Z(n13834) );
  NAND U14436 ( .A(n13835), .B(n13834), .Z(n13838) );
  XNOR U14437 ( .A(n13837), .B(n13836), .Z(n13839) );
  OR U14438 ( .A(n13838), .B(n13839), .Z(n13841) );
  XNOR U14439 ( .A(n13839), .B(n13838), .Z(n14220) );
  NAND U14440 ( .A(a[42]), .B(b[21]), .Z(n14219) );
  OR U14441 ( .A(n14220), .B(n14219), .Z(n13840) );
  NAND U14442 ( .A(n13841), .B(n13840), .Z(n13842) );
  ANDN U14443 ( .B(b[21]), .A(n191), .Z(n13843) );
  OR U14444 ( .A(n13842), .B(n13843), .Z(n13847) );
  XOR U14445 ( .A(n13843), .B(n13842), .Z(n14225) );
  NAND U14446 ( .A(n14225), .B(n14226), .Z(n13846) );
  NAND U14447 ( .A(n13847), .B(n13846), .Z(n13851) );
  NAND U14448 ( .A(a[44]), .B(b[21]), .Z(n13850) );
  OR U14449 ( .A(n13851), .B(n13850), .Z(n13853) );
  XOR U14450 ( .A(n13849), .B(n13848), .Z(n14231) );
  XOR U14451 ( .A(n13851), .B(n13850), .Z(n14232) );
  NAND U14452 ( .A(n14231), .B(n14232), .Z(n13852) );
  NAND U14453 ( .A(n13853), .B(n13852), .Z(n13857) );
  XOR U14454 ( .A(n13855), .B(n13854), .Z(n13856) );
  NAND U14455 ( .A(n13857), .B(n13856), .Z(n13859) );
  XNOR U14456 ( .A(n13857), .B(n13856), .Z(n14238) );
  NAND U14457 ( .A(a[45]), .B(b[21]), .Z(n14237) );
  OR U14458 ( .A(n14238), .B(n14237), .Z(n13858) );
  NAND U14459 ( .A(n13859), .B(n13858), .Z(n13863) );
  NANDN U14460 ( .A(n13862), .B(n13863), .Z(n13865) );
  XNOR U14461 ( .A(n13861), .B(n13860), .Z(n14244) );
  XNOR U14462 ( .A(n13863), .B(n13862), .Z(n14243) );
  NANDN U14463 ( .A(n14244), .B(n14243), .Z(n13864) );
  NAND U14464 ( .A(n13865), .B(n13864), .Z(n13869) );
  XOR U14465 ( .A(n13867), .B(n13866), .Z(n13868) );
  NAND U14466 ( .A(n13869), .B(n13868), .Z(n13871) );
  XNOR U14467 ( .A(n13869), .B(n13868), .Z(n14250) );
  NAND U14468 ( .A(a[47]), .B(b[21]), .Z(n14249) );
  OR U14469 ( .A(n14250), .B(n14249), .Z(n13870) );
  NAND U14470 ( .A(n13871), .B(n13870), .Z(n13875) );
  NANDN U14471 ( .A(n13874), .B(n13875), .Z(n13877) );
  XNOR U14472 ( .A(n13873), .B(n13872), .Z(n14256) );
  XNOR U14473 ( .A(n13875), .B(n13874), .Z(n14255) );
  NANDN U14474 ( .A(n14256), .B(n14255), .Z(n13876) );
  NAND U14475 ( .A(n13877), .B(n13876), .Z(n13881) );
  XOR U14476 ( .A(n13879), .B(n13878), .Z(n13880) );
  NAND U14477 ( .A(n13881), .B(n13880), .Z(n13883) );
  XNOR U14478 ( .A(n13881), .B(n13880), .Z(n14262) );
  NAND U14479 ( .A(a[49]), .B(b[21]), .Z(n14261) );
  OR U14480 ( .A(n14262), .B(n14261), .Z(n13882) );
  NAND U14481 ( .A(n13883), .B(n13882), .Z(n13887) );
  NANDN U14482 ( .A(n13886), .B(n13887), .Z(n13889) );
  XNOR U14483 ( .A(n13885), .B(n13884), .Z(n14268) );
  XNOR U14484 ( .A(n13887), .B(n13886), .Z(n14267) );
  NANDN U14485 ( .A(n14268), .B(n14267), .Z(n13888) );
  NAND U14486 ( .A(n13889), .B(n13888), .Z(n13893) );
  XOR U14487 ( .A(n13891), .B(n13890), .Z(n13892) );
  NAND U14488 ( .A(n13893), .B(n13892), .Z(n13895) );
  XNOR U14489 ( .A(n13893), .B(n13892), .Z(n14274) );
  NAND U14490 ( .A(a[51]), .B(b[21]), .Z(n14273) );
  OR U14491 ( .A(n14274), .B(n14273), .Z(n13894) );
  NAND U14492 ( .A(n13895), .B(n13894), .Z(n13899) );
  NANDN U14493 ( .A(n13898), .B(n13899), .Z(n13901) );
  XNOR U14494 ( .A(n13897), .B(n13896), .Z(n14280) );
  XNOR U14495 ( .A(n13899), .B(n13898), .Z(n14279) );
  NANDN U14496 ( .A(n14280), .B(n14279), .Z(n13900) );
  NAND U14497 ( .A(n13901), .B(n13900), .Z(n13905) );
  XOR U14498 ( .A(n13903), .B(n13902), .Z(n13904) );
  NAND U14499 ( .A(n13905), .B(n13904), .Z(n13907) );
  XNOR U14500 ( .A(n13905), .B(n13904), .Z(n14286) );
  NAND U14501 ( .A(a[53]), .B(b[21]), .Z(n14285) );
  OR U14502 ( .A(n14286), .B(n14285), .Z(n13906) );
  NAND U14503 ( .A(n13907), .B(n13906), .Z(n13911) );
  NANDN U14504 ( .A(n13910), .B(n13911), .Z(n13913) );
  XNOR U14505 ( .A(n13909), .B(n13908), .Z(n14292) );
  XNOR U14506 ( .A(n13911), .B(n13910), .Z(n14291) );
  NANDN U14507 ( .A(n14292), .B(n14291), .Z(n13912) );
  NAND U14508 ( .A(n13913), .B(n13912), .Z(n13917) );
  XOR U14509 ( .A(n13915), .B(n13914), .Z(n13916) );
  NAND U14510 ( .A(n13917), .B(n13916), .Z(n13919) );
  XNOR U14511 ( .A(n13917), .B(n13916), .Z(n14298) );
  NAND U14512 ( .A(a[55]), .B(b[21]), .Z(n14297) );
  OR U14513 ( .A(n14298), .B(n14297), .Z(n13918) );
  NAND U14514 ( .A(n13919), .B(n13918), .Z(n13923) );
  NANDN U14515 ( .A(n13922), .B(n13923), .Z(n13925) );
  XNOR U14516 ( .A(n13921), .B(n13920), .Z(n14304) );
  XNOR U14517 ( .A(n13923), .B(n13922), .Z(n14303) );
  NANDN U14518 ( .A(n14304), .B(n14303), .Z(n13924) );
  NAND U14519 ( .A(n13925), .B(n13924), .Z(n13928) );
  XOR U14520 ( .A(n13927), .B(n13926), .Z(n13929) );
  AND U14521 ( .A(b[21]), .B(a[57]), .Z(n14310) );
  XOR U14522 ( .A(n13929), .B(n13928), .Z(n14309) );
  NAND U14523 ( .A(a[58]), .B(b[21]), .Z(n13932) );
  OR U14524 ( .A(n13933), .B(n13932), .Z(n13935) );
  XNOR U14525 ( .A(n13931), .B(n13930), .Z(n14316) );
  XOR U14526 ( .A(n13933), .B(n13932), .Z(n14315) );
  NANDN U14527 ( .A(n14316), .B(n14315), .Z(n13934) );
  NAND U14528 ( .A(n13935), .B(n13934), .Z(n13939) );
  XOR U14529 ( .A(n13937), .B(n13936), .Z(n13938) );
  NAND U14530 ( .A(n13939), .B(n13938), .Z(n13941) );
  XNOR U14531 ( .A(n13939), .B(n13938), .Z(n14322) );
  NAND U14532 ( .A(a[59]), .B(b[21]), .Z(n14321) );
  OR U14533 ( .A(n14322), .B(n14321), .Z(n13940) );
  NAND U14534 ( .A(n13941), .B(n13940), .Z(n13945) );
  NANDN U14535 ( .A(n13944), .B(n13945), .Z(n13947) );
  XNOR U14536 ( .A(n13943), .B(n13942), .Z(n14330) );
  XNOR U14537 ( .A(n13945), .B(n13944), .Z(n14329) );
  NANDN U14538 ( .A(n14330), .B(n14329), .Z(n13946) );
  NAND U14539 ( .A(n13947), .B(n13946), .Z(n14332) );
  NANDN U14540 ( .A(n14331), .B(n14332), .Z(n13948) );
  NAND U14541 ( .A(n13949), .B(n13948), .Z(n13953) );
  NANDN U14542 ( .A(n13952), .B(n13953), .Z(n13955) );
  XNOR U14543 ( .A(n13951), .B(n13950), .Z(n14338) );
  XNOR U14544 ( .A(n13953), .B(n13952), .Z(n14337) );
  NANDN U14545 ( .A(n14338), .B(n14337), .Z(n13954) );
  NAND U14546 ( .A(n13955), .B(n13954), .Z(n13958) );
  XOR U14547 ( .A(n13957), .B(n13956), .Z(n13959) );
  OR U14548 ( .A(n13958), .B(n13959), .Z(n13961) );
  AND U14549 ( .A(b[21]), .B(a[63]), .Z(n13969) );
  XOR U14550 ( .A(n13959), .B(n13958), .Z(n13968) );
  NANDN U14551 ( .A(n13969), .B(n13968), .Z(n13960) );
  NAND U14552 ( .A(n13961), .B(n13960), .Z(n13966) );
  XNOR U14553 ( .A(n13963), .B(n13962), .Z(n13967) );
  OR U14554 ( .A(n13966), .B(n13967), .Z(n13965) );
  NANDN U14555 ( .A(n13964), .B(n13965), .Z(n21967) );
  XNOR U14556 ( .A(n13965), .B(n13964), .Z(n24166) );
  XOR U14557 ( .A(n13967), .B(n13966), .Z(n24162) );
  XOR U14558 ( .A(n13969), .B(n13968), .Z(n14721) );
  AND U14559 ( .A(b[20]), .B(a[61]), .Z(n14328) );
  NAND U14560 ( .A(a[46]), .B(b[20]), .Z(n14239) );
  ANDN U14561 ( .B(b[20]), .A(n189), .Z(n14208) );
  ANDN U14562 ( .B(b[20]), .A(n187), .Z(n14196) );
  ANDN U14563 ( .B(b[20]), .A(n21772), .Z(n14184) );
  ANDN U14564 ( .B(b[20]), .A(n184), .Z(n14172) );
  ANDN U14565 ( .B(b[20]), .A(n21751), .Z(n14160) );
  ANDN U14566 ( .B(b[20]), .A(n21740), .Z(n14148) );
  ANDN U14567 ( .B(b[20]), .A(n21727), .Z(n14136) );
  ANDN U14568 ( .B(b[20]), .A(n21716), .Z(n14124) );
  ANDN U14569 ( .B(b[20]), .A(n21703), .Z(n14112) );
  ANDN U14570 ( .B(b[20]), .A(n21692), .Z(n14100) );
  ANDN U14571 ( .B(b[20]), .A(n21681), .Z(n14090) );
  ANDN U14572 ( .B(b[20]), .A(n21670), .Z(n14078) );
  ANDN U14573 ( .B(b[20]), .A(n174), .Z(n14066) );
  ANDN U14574 ( .B(b[20]), .A(n172), .Z(n14054) );
  NAND U14575 ( .A(a[13]), .B(b[20]), .Z(n14042) );
  ANDN U14576 ( .B(b[20]), .A(n21164), .Z(n14031) );
  XNOR U14577 ( .A(n13975), .B(n13974), .Z(n14028) );
  ANDN U14578 ( .B(b[20]), .A(n21615), .Z(n14022) );
  NAND U14579 ( .A(a[7]), .B(b[20]), .Z(n14010) );
  NAND U14580 ( .A(a[6]), .B(b[20]), .Z(n14005) );
  XOR U14581 ( .A(n13977), .B(n13976), .Z(n14006) );
  NANDN U14582 ( .A(n14005), .B(n14006), .Z(n14008) );
  ANDN U14583 ( .B(b[20]), .A(n164), .Z(n14000) );
  ANDN U14584 ( .B(b[20]), .A(n21580), .Z(n13987) );
  NAND U14585 ( .A(b[21]), .B(a[1]), .Z(n13980) );
  AND U14586 ( .A(b[20]), .B(a[0]), .Z(n14736) );
  NANDN U14587 ( .A(n13980), .B(n14736), .Z(n13979) );
  NAND U14588 ( .A(a[2]), .B(b[20]), .Z(n13978) );
  AND U14589 ( .A(n13979), .B(n13978), .Z(n13986) );
  NANDN U14590 ( .A(n13980), .B(a[0]), .Z(n13981) );
  XNOR U14591 ( .A(a[2]), .B(n13981), .Z(n13982) );
  NAND U14592 ( .A(b[20]), .B(n13982), .Z(n14363) );
  AND U14593 ( .A(a[1]), .B(b[21]), .Z(n13983) );
  XNOR U14594 ( .A(n13984), .B(n13983), .Z(n14362) );
  NANDN U14595 ( .A(n14363), .B(n14362), .Z(n13985) );
  NANDN U14596 ( .A(n13986), .B(n13985), .Z(n13988) );
  NANDN U14597 ( .A(n13987), .B(n13988), .Z(n13992) );
  XOR U14598 ( .A(n13988), .B(n13987), .Z(n14367) );
  NANDN U14599 ( .A(n14367), .B(n14366), .Z(n13991) );
  NAND U14600 ( .A(n13992), .B(n13991), .Z(n13996) );
  XOR U14601 ( .A(n13994), .B(n13993), .Z(n13995) );
  NANDN U14602 ( .A(n13996), .B(n13995), .Z(n13998) );
  NAND U14603 ( .A(a[4]), .B(b[20]), .Z(n14374) );
  NANDN U14604 ( .A(n14374), .B(n14375), .Z(n13997) );
  NAND U14605 ( .A(n13998), .B(n13997), .Z(n13999) );
  OR U14606 ( .A(n14000), .B(n13999), .Z(n14004) );
  XNOR U14607 ( .A(n14000), .B(n13999), .Z(n14349) );
  XOR U14608 ( .A(n14002), .B(n14001), .Z(n14350) );
  NANDN U14609 ( .A(n14349), .B(n14350), .Z(n14003) );
  NAND U14610 ( .A(n14004), .B(n14003), .Z(n14384) );
  XNOR U14611 ( .A(n14006), .B(n14005), .Z(n14385) );
  NANDN U14612 ( .A(n14384), .B(n14385), .Z(n14007) );
  NAND U14613 ( .A(n14008), .B(n14007), .Z(n14009) );
  NANDN U14614 ( .A(n14010), .B(n14009), .Z(n14014) );
  XNOR U14615 ( .A(n14012), .B(n14011), .Z(n14348) );
  NAND U14616 ( .A(n14347), .B(n14348), .Z(n14013) );
  AND U14617 ( .A(n14014), .B(n14013), .Z(n14018) );
  XOR U14618 ( .A(n14016), .B(n14015), .Z(n14017) );
  NANDN U14619 ( .A(n14018), .B(n14017), .Z(n14020) );
  NAND U14620 ( .A(a[8]), .B(b[20]), .Z(n14394) );
  NANDN U14621 ( .A(n14394), .B(n14395), .Z(n14019) );
  NAND U14622 ( .A(n14020), .B(n14019), .Z(n14021) );
  OR U14623 ( .A(n14022), .B(n14021), .Z(n14026) );
  XNOR U14624 ( .A(n14022), .B(n14021), .Z(n14398) );
  XOR U14625 ( .A(n14024), .B(n14023), .Z(n14399) );
  NANDN U14626 ( .A(n14398), .B(n14399), .Z(n14025) );
  NAND U14627 ( .A(n14026), .B(n14025), .Z(n14027) );
  NANDN U14628 ( .A(n14028), .B(n14027), .Z(n14030) );
  ANDN U14629 ( .B(b[20]), .A(n168), .Z(n14405) );
  NANDN U14630 ( .A(n14405), .B(n14404), .Z(n14029) );
  NAND U14631 ( .A(n14030), .B(n14029), .Z(n14032) );
  NANDN U14632 ( .A(n14031), .B(n14032), .Z(n14036) );
  XOR U14633 ( .A(n14032), .B(n14031), .Z(n14411) );
  XOR U14634 ( .A(n14034), .B(n14033), .Z(n14410) );
  OR U14635 ( .A(n14411), .B(n14410), .Z(n14035) );
  AND U14636 ( .A(n14036), .B(n14035), .Z(n14037) );
  OR U14637 ( .A(n14038), .B(n14037), .Z(n14040) );
  ANDN U14638 ( .B(b[20]), .A(n169), .Z(n14419) );
  XNOR U14639 ( .A(n14038), .B(n14037), .Z(n14418) );
  OR U14640 ( .A(n14419), .B(n14418), .Z(n14039) );
  AND U14641 ( .A(n14040), .B(n14039), .Z(n14041) );
  NANDN U14642 ( .A(n14042), .B(n14041), .Z(n14046) );
  XNOR U14643 ( .A(n14044), .B(n14043), .Z(n14346) );
  NAND U14644 ( .A(n14345), .B(n14346), .Z(n14045) );
  AND U14645 ( .A(n14046), .B(n14045), .Z(n14049) );
  XOR U14646 ( .A(n14048), .B(n14047), .Z(n14050) );
  NANDN U14647 ( .A(n14049), .B(n14050), .Z(n14052) );
  NAND U14648 ( .A(a[14]), .B(b[20]), .Z(n14428) );
  XNOR U14649 ( .A(n14050), .B(n14049), .Z(n14429) );
  NANDN U14650 ( .A(n14428), .B(n14429), .Z(n14051) );
  NAND U14651 ( .A(n14052), .B(n14051), .Z(n14053) );
  OR U14652 ( .A(n14054), .B(n14053), .Z(n14058) );
  XNOR U14653 ( .A(n14054), .B(n14053), .Z(n14432) );
  XOR U14654 ( .A(n14056), .B(n14055), .Z(n14433) );
  NANDN U14655 ( .A(n14432), .B(n14433), .Z(n14057) );
  NAND U14656 ( .A(n14058), .B(n14057), .Z(n14061) );
  XOR U14657 ( .A(n14060), .B(n14059), .Z(n14062) );
  NANDN U14658 ( .A(n14061), .B(n14062), .Z(n14064) );
  NAND U14659 ( .A(a[16]), .B(b[20]), .Z(n14440) );
  XNOR U14660 ( .A(n14062), .B(n14061), .Z(n14441) );
  NANDN U14661 ( .A(n14440), .B(n14441), .Z(n14063) );
  NAND U14662 ( .A(n14064), .B(n14063), .Z(n14065) );
  OR U14663 ( .A(n14066), .B(n14065), .Z(n14070) );
  XNOR U14664 ( .A(n14066), .B(n14065), .Z(n14444) );
  XOR U14665 ( .A(n14068), .B(n14067), .Z(n14445) );
  NANDN U14666 ( .A(n14444), .B(n14445), .Z(n14069) );
  NAND U14667 ( .A(n14070), .B(n14069), .Z(n14073) );
  XOR U14668 ( .A(n14072), .B(n14071), .Z(n14074) );
  NANDN U14669 ( .A(n14073), .B(n14074), .Z(n14076) );
  NAND U14670 ( .A(a[18]), .B(b[20]), .Z(n14452) );
  XNOR U14671 ( .A(n14074), .B(n14073), .Z(n14453) );
  NANDN U14672 ( .A(n14452), .B(n14453), .Z(n14075) );
  NAND U14673 ( .A(n14076), .B(n14075), .Z(n14077) );
  OR U14674 ( .A(n14078), .B(n14077), .Z(n14082) );
  XNOR U14675 ( .A(n14078), .B(n14077), .Z(n14456) );
  XOR U14676 ( .A(n14080), .B(n14079), .Z(n14457) );
  NANDN U14677 ( .A(n14456), .B(n14457), .Z(n14081) );
  NAND U14678 ( .A(n14082), .B(n14081), .Z(n14085) );
  XOR U14679 ( .A(n14084), .B(n14083), .Z(n14086) );
  NANDN U14680 ( .A(n14085), .B(n14086), .Z(n14088) );
  NAND U14681 ( .A(a[20]), .B(b[20]), .Z(n14464) );
  XNOR U14682 ( .A(n14086), .B(n14085), .Z(n14465) );
  NANDN U14683 ( .A(n14464), .B(n14465), .Z(n14087) );
  NAND U14684 ( .A(n14088), .B(n14087), .Z(n14089) );
  OR U14685 ( .A(n14090), .B(n14089), .Z(n14094) );
  XNOR U14686 ( .A(n14090), .B(n14089), .Z(n14468) );
  XOR U14687 ( .A(n14092), .B(n14091), .Z(n14469) );
  NANDN U14688 ( .A(n14468), .B(n14469), .Z(n14093) );
  NAND U14689 ( .A(n14094), .B(n14093), .Z(n14095) );
  OR U14690 ( .A(n14096), .B(n14095), .Z(n14098) );
  NAND U14691 ( .A(a[22]), .B(b[20]), .Z(n14476) );
  XOR U14692 ( .A(n14096), .B(n14095), .Z(n14477) );
  NANDN U14693 ( .A(n14476), .B(n14477), .Z(n14097) );
  NAND U14694 ( .A(n14098), .B(n14097), .Z(n14099) );
  OR U14695 ( .A(n14100), .B(n14099), .Z(n14104) );
  XNOR U14696 ( .A(n14100), .B(n14099), .Z(n14480) );
  XOR U14697 ( .A(n14102), .B(n14101), .Z(n14481) );
  NANDN U14698 ( .A(n14480), .B(n14481), .Z(n14103) );
  NAND U14699 ( .A(n14104), .B(n14103), .Z(n14107) );
  XOR U14700 ( .A(n14106), .B(n14105), .Z(n14108) );
  NANDN U14701 ( .A(n14107), .B(n14108), .Z(n14110) );
  NAND U14702 ( .A(a[24]), .B(b[20]), .Z(n14488) );
  XNOR U14703 ( .A(n14108), .B(n14107), .Z(n14489) );
  NANDN U14704 ( .A(n14488), .B(n14489), .Z(n14109) );
  NAND U14705 ( .A(n14110), .B(n14109), .Z(n14111) );
  OR U14706 ( .A(n14112), .B(n14111), .Z(n14116) );
  XNOR U14707 ( .A(n14112), .B(n14111), .Z(n14492) );
  XOR U14708 ( .A(n14114), .B(n14113), .Z(n14493) );
  NANDN U14709 ( .A(n14492), .B(n14493), .Z(n14115) );
  NAND U14710 ( .A(n14116), .B(n14115), .Z(n14119) );
  XOR U14711 ( .A(n14118), .B(n14117), .Z(n14120) );
  NANDN U14712 ( .A(n14119), .B(n14120), .Z(n14122) );
  NAND U14713 ( .A(a[26]), .B(b[20]), .Z(n14500) );
  XNOR U14714 ( .A(n14120), .B(n14119), .Z(n14501) );
  NANDN U14715 ( .A(n14500), .B(n14501), .Z(n14121) );
  NAND U14716 ( .A(n14122), .B(n14121), .Z(n14123) );
  OR U14717 ( .A(n14124), .B(n14123), .Z(n14128) );
  XNOR U14718 ( .A(n14124), .B(n14123), .Z(n14504) );
  XOR U14719 ( .A(n14126), .B(n14125), .Z(n14505) );
  NANDN U14720 ( .A(n14504), .B(n14505), .Z(n14127) );
  NAND U14721 ( .A(n14128), .B(n14127), .Z(n14131) );
  XOR U14722 ( .A(n14130), .B(n14129), .Z(n14132) );
  NANDN U14723 ( .A(n14131), .B(n14132), .Z(n14134) );
  NAND U14724 ( .A(a[28]), .B(b[20]), .Z(n14512) );
  XNOR U14725 ( .A(n14132), .B(n14131), .Z(n14513) );
  NANDN U14726 ( .A(n14512), .B(n14513), .Z(n14133) );
  NAND U14727 ( .A(n14134), .B(n14133), .Z(n14135) );
  OR U14728 ( .A(n14136), .B(n14135), .Z(n14140) );
  XNOR U14729 ( .A(n14136), .B(n14135), .Z(n14516) );
  XOR U14730 ( .A(n14138), .B(n14137), .Z(n14517) );
  NANDN U14731 ( .A(n14516), .B(n14517), .Z(n14139) );
  NAND U14732 ( .A(n14140), .B(n14139), .Z(n14143) );
  XOR U14733 ( .A(n14142), .B(n14141), .Z(n14144) );
  NANDN U14734 ( .A(n14143), .B(n14144), .Z(n14146) );
  NAND U14735 ( .A(a[30]), .B(b[20]), .Z(n14524) );
  XNOR U14736 ( .A(n14144), .B(n14143), .Z(n14525) );
  NANDN U14737 ( .A(n14524), .B(n14525), .Z(n14145) );
  NAND U14738 ( .A(n14146), .B(n14145), .Z(n14147) );
  OR U14739 ( .A(n14148), .B(n14147), .Z(n14152) );
  XNOR U14740 ( .A(n14148), .B(n14147), .Z(n14528) );
  XOR U14741 ( .A(n14150), .B(n14149), .Z(n14529) );
  NANDN U14742 ( .A(n14528), .B(n14529), .Z(n14151) );
  NAND U14743 ( .A(n14152), .B(n14151), .Z(n14155) );
  XOR U14744 ( .A(n14154), .B(n14153), .Z(n14156) );
  NANDN U14745 ( .A(n14155), .B(n14156), .Z(n14158) );
  NAND U14746 ( .A(a[32]), .B(b[20]), .Z(n14536) );
  XNOR U14747 ( .A(n14156), .B(n14155), .Z(n14537) );
  NANDN U14748 ( .A(n14536), .B(n14537), .Z(n14157) );
  NAND U14749 ( .A(n14158), .B(n14157), .Z(n14159) );
  OR U14750 ( .A(n14160), .B(n14159), .Z(n14164) );
  XNOR U14751 ( .A(n14160), .B(n14159), .Z(n14540) );
  XOR U14752 ( .A(n14162), .B(n14161), .Z(n14541) );
  NANDN U14753 ( .A(n14540), .B(n14541), .Z(n14163) );
  NAND U14754 ( .A(n14164), .B(n14163), .Z(n14167) );
  XOR U14755 ( .A(n14166), .B(n14165), .Z(n14168) );
  NANDN U14756 ( .A(n14167), .B(n14168), .Z(n14170) );
  NAND U14757 ( .A(a[34]), .B(b[20]), .Z(n14548) );
  XNOR U14758 ( .A(n14168), .B(n14167), .Z(n14549) );
  NANDN U14759 ( .A(n14548), .B(n14549), .Z(n14169) );
  NAND U14760 ( .A(n14170), .B(n14169), .Z(n14171) );
  OR U14761 ( .A(n14172), .B(n14171), .Z(n14176) );
  XNOR U14762 ( .A(n14172), .B(n14171), .Z(n14552) );
  XOR U14763 ( .A(n14174), .B(n14173), .Z(n14553) );
  NANDN U14764 ( .A(n14552), .B(n14553), .Z(n14175) );
  NAND U14765 ( .A(n14176), .B(n14175), .Z(n14179) );
  XOR U14766 ( .A(n14178), .B(n14177), .Z(n14180) );
  NANDN U14767 ( .A(n14179), .B(n14180), .Z(n14182) );
  NAND U14768 ( .A(a[36]), .B(b[20]), .Z(n14560) );
  XNOR U14769 ( .A(n14180), .B(n14179), .Z(n14561) );
  NANDN U14770 ( .A(n14560), .B(n14561), .Z(n14181) );
  NAND U14771 ( .A(n14182), .B(n14181), .Z(n14183) );
  OR U14772 ( .A(n14184), .B(n14183), .Z(n14188) );
  XNOR U14773 ( .A(n14184), .B(n14183), .Z(n14564) );
  XOR U14774 ( .A(n14186), .B(n14185), .Z(n14565) );
  NANDN U14775 ( .A(n14564), .B(n14565), .Z(n14187) );
  NAND U14776 ( .A(n14188), .B(n14187), .Z(n14191) );
  XOR U14777 ( .A(n14190), .B(n14189), .Z(n14192) );
  NANDN U14778 ( .A(n14191), .B(n14192), .Z(n14194) );
  NAND U14779 ( .A(a[38]), .B(b[20]), .Z(n14572) );
  XNOR U14780 ( .A(n14192), .B(n14191), .Z(n14573) );
  NANDN U14781 ( .A(n14572), .B(n14573), .Z(n14193) );
  NAND U14782 ( .A(n14194), .B(n14193), .Z(n14195) );
  OR U14783 ( .A(n14196), .B(n14195), .Z(n14200) );
  XNOR U14784 ( .A(n14196), .B(n14195), .Z(n14576) );
  XOR U14785 ( .A(n14198), .B(n14197), .Z(n14577) );
  NANDN U14786 ( .A(n14576), .B(n14577), .Z(n14199) );
  NAND U14787 ( .A(n14200), .B(n14199), .Z(n14203) );
  XOR U14788 ( .A(n14202), .B(n14201), .Z(n14204) );
  NANDN U14789 ( .A(n14203), .B(n14204), .Z(n14206) );
  NAND U14790 ( .A(a[40]), .B(b[20]), .Z(n14584) );
  XNOR U14791 ( .A(n14204), .B(n14203), .Z(n14585) );
  NANDN U14792 ( .A(n14584), .B(n14585), .Z(n14205) );
  NAND U14793 ( .A(n14206), .B(n14205), .Z(n14207) );
  OR U14794 ( .A(n14208), .B(n14207), .Z(n14212) );
  XNOR U14795 ( .A(n14208), .B(n14207), .Z(n14588) );
  XOR U14796 ( .A(n14210), .B(n14209), .Z(n14589) );
  NANDN U14797 ( .A(n14588), .B(n14589), .Z(n14211) );
  NAND U14798 ( .A(n14212), .B(n14211), .Z(n14215) );
  XNOR U14799 ( .A(n14214), .B(n14213), .Z(n14216) );
  OR U14800 ( .A(n14215), .B(n14216), .Z(n14218) );
  XNOR U14801 ( .A(n14216), .B(n14215), .Z(n14595) );
  NAND U14802 ( .A(a[42]), .B(b[20]), .Z(n14594) );
  OR U14803 ( .A(n14595), .B(n14594), .Z(n14217) );
  NAND U14804 ( .A(n14218), .B(n14217), .Z(n14221) );
  ANDN U14805 ( .B(b[20]), .A(n191), .Z(n14222) );
  OR U14806 ( .A(n14221), .B(n14222), .Z(n14224) );
  XOR U14807 ( .A(n14220), .B(n14219), .Z(n14601) );
  XOR U14808 ( .A(n14222), .B(n14221), .Z(n14600) );
  NANDN U14809 ( .A(n14601), .B(n14600), .Z(n14223) );
  NAND U14810 ( .A(n14224), .B(n14223), .Z(n14228) );
  AND U14811 ( .A(b[20]), .B(a[44]), .Z(n14227) );
  NANDN U14812 ( .A(n14228), .B(n14227), .Z(n14230) );
  XNOR U14813 ( .A(n14228), .B(n14227), .Z(n14608) );
  NANDN U14814 ( .A(n14609), .B(n14608), .Z(n14229) );
  NAND U14815 ( .A(n14230), .B(n14229), .Z(n14234) );
  XOR U14816 ( .A(n14232), .B(n14231), .Z(n14233) );
  NAND U14817 ( .A(n14234), .B(n14233), .Z(n14236) );
  XNOR U14818 ( .A(n14234), .B(n14233), .Z(n14613) );
  NAND U14819 ( .A(a[45]), .B(b[20]), .Z(n14612) );
  OR U14820 ( .A(n14613), .B(n14612), .Z(n14235) );
  NAND U14821 ( .A(n14236), .B(n14235), .Z(n14240) );
  NANDN U14822 ( .A(n14239), .B(n14240), .Z(n14242) );
  XOR U14823 ( .A(n14238), .B(n14237), .Z(n14618) );
  XNOR U14824 ( .A(n14240), .B(n14239), .Z(n14619) );
  NAND U14825 ( .A(n14618), .B(n14619), .Z(n14241) );
  NAND U14826 ( .A(n14242), .B(n14241), .Z(n14245) );
  AND U14827 ( .A(b[20]), .B(a[47]), .Z(n14246) );
  OR U14828 ( .A(n14245), .B(n14246), .Z(n14248) );
  XNOR U14829 ( .A(n14244), .B(n14243), .Z(n14625) );
  XOR U14830 ( .A(n14246), .B(n14245), .Z(n14624) );
  NANDN U14831 ( .A(n14625), .B(n14624), .Z(n14247) );
  NAND U14832 ( .A(n14248), .B(n14247), .Z(n14252) );
  NAND U14833 ( .A(a[48]), .B(b[20]), .Z(n14251) );
  OR U14834 ( .A(n14252), .B(n14251), .Z(n14254) );
  XOR U14835 ( .A(n14250), .B(n14249), .Z(n14630) );
  XOR U14836 ( .A(n14252), .B(n14251), .Z(n14631) );
  NAND U14837 ( .A(n14630), .B(n14631), .Z(n14253) );
  NAND U14838 ( .A(n14254), .B(n14253), .Z(n14257) );
  AND U14839 ( .A(b[20]), .B(a[49]), .Z(n14258) );
  OR U14840 ( .A(n14257), .B(n14258), .Z(n14260) );
  XNOR U14841 ( .A(n14256), .B(n14255), .Z(n14637) );
  XOR U14842 ( .A(n14258), .B(n14257), .Z(n14636) );
  NANDN U14843 ( .A(n14637), .B(n14636), .Z(n14259) );
  NAND U14844 ( .A(n14260), .B(n14259), .Z(n14264) );
  NAND U14845 ( .A(a[50]), .B(b[20]), .Z(n14263) );
  OR U14846 ( .A(n14264), .B(n14263), .Z(n14266) );
  XOR U14847 ( .A(n14262), .B(n14261), .Z(n14642) );
  XOR U14848 ( .A(n14264), .B(n14263), .Z(n14643) );
  NAND U14849 ( .A(n14642), .B(n14643), .Z(n14265) );
  NAND U14850 ( .A(n14266), .B(n14265), .Z(n14269) );
  AND U14851 ( .A(b[20]), .B(a[51]), .Z(n14270) );
  OR U14852 ( .A(n14269), .B(n14270), .Z(n14272) );
  XNOR U14853 ( .A(n14268), .B(n14267), .Z(n14649) );
  XOR U14854 ( .A(n14270), .B(n14269), .Z(n14648) );
  NANDN U14855 ( .A(n14649), .B(n14648), .Z(n14271) );
  NAND U14856 ( .A(n14272), .B(n14271), .Z(n14276) );
  NAND U14857 ( .A(a[52]), .B(b[20]), .Z(n14275) );
  OR U14858 ( .A(n14276), .B(n14275), .Z(n14278) );
  XOR U14859 ( .A(n14274), .B(n14273), .Z(n14654) );
  XOR U14860 ( .A(n14276), .B(n14275), .Z(n14655) );
  NAND U14861 ( .A(n14654), .B(n14655), .Z(n14277) );
  NAND U14862 ( .A(n14278), .B(n14277), .Z(n14281) );
  AND U14863 ( .A(b[20]), .B(a[53]), .Z(n14282) );
  OR U14864 ( .A(n14281), .B(n14282), .Z(n14284) );
  XNOR U14865 ( .A(n14280), .B(n14279), .Z(n14661) );
  XOR U14866 ( .A(n14282), .B(n14281), .Z(n14660) );
  NANDN U14867 ( .A(n14661), .B(n14660), .Z(n14283) );
  NAND U14868 ( .A(n14284), .B(n14283), .Z(n14288) );
  NAND U14869 ( .A(a[54]), .B(b[20]), .Z(n14287) );
  OR U14870 ( .A(n14288), .B(n14287), .Z(n14290) );
  XOR U14871 ( .A(n14286), .B(n14285), .Z(n14666) );
  XOR U14872 ( .A(n14288), .B(n14287), .Z(n14667) );
  NAND U14873 ( .A(n14666), .B(n14667), .Z(n14289) );
  NAND U14874 ( .A(n14290), .B(n14289), .Z(n14293) );
  AND U14875 ( .A(b[20]), .B(a[55]), .Z(n14294) );
  OR U14876 ( .A(n14293), .B(n14294), .Z(n14296) );
  XNOR U14877 ( .A(n14292), .B(n14291), .Z(n14673) );
  XOR U14878 ( .A(n14294), .B(n14293), .Z(n14672) );
  NANDN U14879 ( .A(n14673), .B(n14672), .Z(n14295) );
  NAND U14880 ( .A(n14296), .B(n14295), .Z(n14300) );
  NAND U14881 ( .A(a[56]), .B(b[20]), .Z(n14299) );
  OR U14882 ( .A(n14300), .B(n14299), .Z(n14302) );
  XOR U14883 ( .A(n14298), .B(n14297), .Z(n14678) );
  XOR U14884 ( .A(n14300), .B(n14299), .Z(n14679) );
  NAND U14885 ( .A(n14678), .B(n14679), .Z(n14301) );
  NAND U14886 ( .A(n14302), .B(n14301), .Z(n14305) );
  AND U14887 ( .A(b[20]), .B(a[57]), .Z(n14306) );
  OR U14888 ( .A(n14305), .B(n14306), .Z(n14308) );
  XNOR U14889 ( .A(n14304), .B(n14303), .Z(n14685) );
  XOR U14890 ( .A(n14306), .B(n14305), .Z(n14684) );
  NANDN U14891 ( .A(n14685), .B(n14684), .Z(n14307) );
  NAND U14892 ( .A(n14308), .B(n14307), .Z(n14312) );
  NAND U14893 ( .A(a[58]), .B(b[20]), .Z(n14311) );
  OR U14894 ( .A(n14312), .B(n14311), .Z(n14314) );
  XOR U14895 ( .A(n14310), .B(n14309), .Z(n14691) );
  XOR U14896 ( .A(n14312), .B(n14311), .Z(n14690) );
  NAND U14897 ( .A(n14691), .B(n14690), .Z(n14313) );
  NAND U14898 ( .A(n14314), .B(n14313), .Z(n14317) );
  AND U14899 ( .A(b[20]), .B(a[59]), .Z(n14318) );
  OR U14900 ( .A(n14317), .B(n14318), .Z(n14320) );
  XNOR U14901 ( .A(n14316), .B(n14315), .Z(n14697) );
  XOR U14902 ( .A(n14318), .B(n14317), .Z(n14696) );
  NANDN U14903 ( .A(n14697), .B(n14696), .Z(n14319) );
  NAND U14904 ( .A(n14320), .B(n14319), .Z(n14324) );
  NAND U14905 ( .A(a[60]), .B(b[20]), .Z(n14323) );
  OR U14906 ( .A(n14324), .B(n14323), .Z(n14326) );
  XOR U14907 ( .A(n14322), .B(n14321), .Z(n14702) );
  XOR U14908 ( .A(n14324), .B(n14323), .Z(n14703) );
  NAND U14909 ( .A(n14702), .B(n14703), .Z(n14325) );
  AND U14910 ( .A(n14326), .B(n14325), .Z(n14327) );
  XOR U14911 ( .A(n14328), .B(n14327), .Z(n14708) );
  XOR U14912 ( .A(n14330), .B(n14329), .Z(n14709) );
  NAND U14913 ( .A(a[62]), .B(b[20]), .Z(n14333) );
  OR U14914 ( .A(n14334), .B(n14333), .Z(n14336) );
  XNOR U14915 ( .A(n14332), .B(n14331), .Z(n14343) );
  XOR U14916 ( .A(n14334), .B(n14333), .Z(n14344) );
  NAND U14917 ( .A(n14343), .B(n14344), .Z(n14335) );
  NAND U14918 ( .A(n14336), .B(n14335), .Z(n14339) );
  AND U14919 ( .A(b[20]), .B(a[63]), .Z(n14340) );
  OR U14920 ( .A(n14339), .B(n14340), .Z(n14342) );
  XOR U14921 ( .A(n14338), .B(n14337), .Z(n14719) );
  XOR U14922 ( .A(n14340), .B(n14339), .Z(n14718) );
  NAND U14923 ( .A(n14719), .B(n14718), .Z(n14341) );
  AND U14924 ( .A(n14342), .B(n14341), .Z(n14720) );
  NAND U14925 ( .A(n14721), .B(n14720), .Z(n24163) );
  XNOR U14926 ( .A(n14344), .B(n14343), .Z(n14715) );
  NAND U14927 ( .A(a[63]), .B(b[19]), .Z(n14714) );
  OR U14928 ( .A(n14715), .B(n14714), .Z(n14717) );
  NAND U14929 ( .A(a[62]), .B(b[19]), .Z(n14710) );
  NAND U14930 ( .A(a[58]), .B(b[19]), .Z(n14686) );
  NAND U14931 ( .A(a[56]), .B(b[19]), .Z(n14674) );
  NAND U14932 ( .A(a[54]), .B(b[19]), .Z(n14662) );
  NAND U14933 ( .A(a[52]), .B(b[19]), .Z(n14650) );
  NAND U14934 ( .A(a[50]), .B(b[19]), .Z(n14638) );
  NAND U14935 ( .A(a[48]), .B(b[19]), .Z(n14626) );
  ANDN U14936 ( .B(b[19]), .A(n189), .Z(n14583) );
  ANDN U14937 ( .B(b[19]), .A(n187), .Z(n14571) );
  ANDN U14938 ( .B(b[19]), .A(n21772), .Z(n14559) );
  ANDN U14939 ( .B(b[19]), .A(n184), .Z(n14547) );
  ANDN U14940 ( .B(b[19]), .A(n21751), .Z(n14535) );
  ANDN U14941 ( .B(b[19]), .A(n21740), .Z(n14523) );
  ANDN U14942 ( .B(b[19]), .A(n21727), .Z(n14511) );
  ANDN U14943 ( .B(b[19]), .A(n21716), .Z(n14499) );
  ANDN U14944 ( .B(b[19]), .A(n21703), .Z(n14487) );
  ANDN U14945 ( .B(b[19]), .A(n21692), .Z(n14475) );
  ANDN U14946 ( .B(b[19]), .A(n21681), .Z(n14463) );
  ANDN U14947 ( .B(b[19]), .A(n21670), .Z(n14451) );
  ANDN U14948 ( .B(b[19]), .A(n174), .Z(n14439) );
  NAND U14949 ( .A(a[15]), .B(b[19]), .Z(n14427) );
  ANDN U14950 ( .B(b[19]), .A(n170), .Z(n14417) );
  ANDN U14951 ( .B(b[19]), .A(n21164), .Z(n14407) );
  ANDN U14952 ( .B(b[19]), .A(n21615), .Z(n14393) );
  ANDN U14953 ( .B(b[19]), .A(n166), .Z(n14383) );
  NAND U14954 ( .A(a[6]), .B(b[19]), .Z(n14378) );
  XOR U14955 ( .A(n14350), .B(n14349), .Z(n14379) );
  NANDN U14956 ( .A(n14378), .B(n14379), .Z(n14381) );
  ANDN U14957 ( .B(b[19]), .A(n164), .Z(n14373) );
  ANDN U14958 ( .B(b[19]), .A(n21580), .Z(n14360) );
  NAND U14959 ( .A(b[20]), .B(a[1]), .Z(n14353) );
  AND U14960 ( .A(b[19]), .B(a[0]), .Z(n15117) );
  NANDN U14961 ( .A(n14353), .B(n15117), .Z(n14352) );
  NAND U14962 ( .A(a[2]), .B(b[19]), .Z(n14351) );
  AND U14963 ( .A(n14352), .B(n14351), .Z(n14359) );
  NANDN U14964 ( .A(n14353), .B(a[0]), .Z(n14354) );
  XNOR U14965 ( .A(a[2]), .B(n14354), .Z(n14355) );
  NAND U14966 ( .A(b[19]), .B(n14355), .Z(n14742) );
  AND U14967 ( .A(a[1]), .B(b[20]), .Z(n14356) );
  XNOR U14968 ( .A(n14357), .B(n14356), .Z(n14741) );
  NANDN U14969 ( .A(n14742), .B(n14741), .Z(n14358) );
  NANDN U14970 ( .A(n14359), .B(n14358), .Z(n14361) );
  NANDN U14971 ( .A(n14360), .B(n14361), .Z(n14365) );
  XOR U14972 ( .A(n14361), .B(n14360), .Z(n14746) );
  NANDN U14973 ( .A(n14746), .B(n14745), .Z(n14364) );
  NAND U14974 ( .A(n14365), .B(n14364), .Z(n14369) );
  XOR U14975 ( .A(n14367), .B(n14366), .Z(n14368) );
  NANDN U14976 ( .A(n14369), .B(n14368), .Z(n14371) );
  NAND U14977 ( .A(a[4]), .B(b[19]), .Z(n14753) );
  NANDN U14978 ( .A(n14753), .B(n14754), .Z(n14370) );
  NAND U14979 ( .A(n14371), .B(n14370), .Z(n14372) );
  OR U14980 ( .A(n14373), .B(n14372), .Z(n14377) );
  XNOR U14981 ( .A(n14373), .B(n14372), .Z(n14728) );
  XOR U14982 ( .A(n14375), .B(n14374), .Z(n14729) );
  NANDN U14983 ( .A(n14728), .B(n14729), .Z(n14376) );
  NAND U14984 ( .A(n14377), .B(n14376), .Z(n14763) );
  XNOR U14985 ( .A(n14379), .B(n14378), .Z(n14764) );
  NANDN U14986 ( .A(n14763), .B(n14764), .Z(n14380) );
  NAND U14987 ( .A(n14381), .B(n14380), .Z(n14382) );
  OR U14988 ( .A(n14383), .B(n14382), .Z(n14387) );
  XNOR U14989 ( .A(n14383), .B(n14382), .Z(n14767) );
  XOR U14990 ( .A(n14385), .B(n14384), .Z(n14768) );
  NANDN U14991 ( .A(n14767), .B(n14768), .Z(n14386) );
  AND U14992 ( .A(n14387), .B(n14386), .Z(n14388) );
  OR U14993 ( .A(n14389), .B(n14388), .Z(n14391) );
  ANDN U14994 ( .B(b[19]), .A(n167), .Z(n14776) );
  XNOR U14995 ( .A(n14389), .B(n14388), .Z(n14775) );
  OR U14996 ( .A(n14776), .B(n14775), .Z(n14390) );
  NAND U14997 ( .A(n14391), .B(n14390), .Z(n14392) );
  NANDN U14998 ( .A(n14393), .B(n14392), .Z(n14397) );
  XOR U14999 ( .A(n14395), .B(n14394), .Z(n14779) );
  NANDN U15000 ( .A(n14780), .B(n14779), .Z(n14396) );
  NAND U15001 ( .A(n14397), .B(n14396), .Z(n14400) );
  XOR U15002 ( .A(n14399), .B(n14398), .Z(n14401) );
  NANDN U15003 ( .A(n14400), .B(n14401), .Z(n14403) );
  NAND U15004 ( .A(a[10]), .B(b[19]), .Z(n14787) );
  XNOR U15005 ( .A(n14401), .B(n14400), .Z(n14788) );
  NANDN U15006 ( .A(n14787), .B(n14788), .Z(n14402) );
  NAND U15007 ( .A(n14403), .B(n14402), .Z(n14406) );
  OR U15008 ( .A(n14407), .B(n14406), .Z(n14409) );
  XOR U15009 ( .A(n14405), .B(n14404), .Z(n14791) );
  XOR U15010 ( .A(n14407), .B(n14406), .Z(n14792) );
  NANDN U15011 ( .A(n14791), .B(n14792), .Z(n14408) );
  NAND U15012 ( .A(n14409), .B(n14408), .Z(n14413) );
  XNOR U15013 ( .A(n14411), .B(n14410), .Z(n14412) );
  NANDN U15014 ( .A(n14413), .B(n14412), .Z(n14415) );
  NAND U15015 ( .A(a[12]), .B(b[19]), .Z(n14799) );
  NANDN U15016 ( .A(n14799), .B(n14800), .Z(n14414) );
  NAND U15017 ( .A(n14415), .B(n14414), .Z(n14416) );
  OR U15018 ( .A(n14417), .B(n14416), .Z(n14421) );
  XOR U15019 ( .A(n14417), .B(n14416), .Z(n14803) );
  XOR U15020 ( .A(n14419), .B(n14418), .Z(n14804) );
  NAND U15021 ( .A(n14803), .B(n14804), .Z(n14420) );
  AND U15022 ( .A(n14421), .B(n14420), .Z(n14422) );
  OR U15023 ( .A(n14423), .B(n14422), .Z(n14425) );
  ANDN U15024 ( .B(b[19]), .A(n171), .Z(n14812) );
  XNOR U15025 ( .A(n14423), .B(n14422), .Z(n14811) );
  OR U15026 ( .A(n14812), .B(n14811), .Z(n14424) );
  AND U15027 ( .A(n14425), .B(n14424), .Z(n14426) );
  NANDN U15028 ( .A(n14427), .B(n14426), .Z(n14431) );
  XNOR U15029 ( .A(n14429), .B(n14428), .Z(n14727) );
  NAND U15030 ( .A(n14726), .B(n14727), .Z(n14430) );
  AND U15031 ( .A(n14431), .B(n14430), .Z(n14434) );
  XOR U15032 ( .A(n14433), .B(n14432), .Z(n14435) );
  NANDN U15033 ( .A(n14434), .B(n14435), .Z(n14437) );
  NAND U15034 ( .A(a[16]), .B(b[19]), .Z(n14821) );
  XNOR U15035 ( .A(n14435), .B(n14434), .Z(n14822) );
  NANDN U15036 ( .A(n14821), .B(n14822), .Z(n14436) );
  NAND U15037 ( .A(n14437), .B(n14436), .Z(n14438) );
  OR U15038 ( .A(n14439), .B(n14438), .Z(n14443) );
  XNOR U15039 ( .A(n14439), .B(n14438), .Z(n14825) );
  XOR U15040 ( .A(n14441), .B(n14440), .Z(n14826) );
  NANDN U15041 ( .A(n14825), .B(n14826), .Z(n14442) );
  NAND U15042 ( .A(n14443), .B(n14442), .Z(n14446) );
  XOR U15043 ( .A(n14445), .B(n14444), .Z(n14447) );
  NANDN U15044 ( .A(n14446), .B(n14447), .Z(n14449) );
  NAND U15045 ( .A(a[18]), .B(b[19]), .Z(n14833) );
  XNOR U15046 ( .A(n14447), .B(n14446), .Z(n14834) );
  NANDN U15047 ( .A(n14833), .B(n14834), .Z(n14448) );
  NAND U15048 ( .A(n14449), .B(n14448), .Z(n14450) );
  OR U15049 ( .A(n14451), .B(n14450), .Z(n14455) );
  XNOR U15050 ( .A(n14451), .B(n14450), .Z(n14837) );
  XOR U15051 ( .A(n14453), .B(n14452), .Z(n14838) );
  NANDN U15052 ( .A(n14837), .B(n14838), .Z(n14454) );
  NAND U15053 ( .A(n14455), .B(n14454), .Z(n14458) );
  XOR U15054 ( .A(n14457), .B(n14456), .Z(n14459) );
  NANDN U15055 ( .A(n14458), .B(n14459), .Z(n14461) );
  NAND U15056 ( .A(a[20]), .B(b[19]), .Z(n14845) );
  XNOR U15057 ( .A(n14459), .B(n14458), .Z(n14846) );
  NANDN U15058 ( .A(n14845), .B(n14846), .Z(n14460) );
  NAND U15059 ( .A(n14461), .B(n14460), .Z(n14462) );
  OR U15060 ( .A(n14463), .B(n14462), .Z(n14467) );
  XNOR U15061 ( .A(n14463), .B(n14462), .Z(n14849) );
  XOR U15062 ( .A(n14465), .B(n14464), .Z(n14850) );
  NANDN U15063 ( .A(n14849), .B(n14850), .Z(n14466) );
  NAND U15064 ( .A(n14467), .B(n14466), .Z(n14470) );
  XOR U15065 ( .A(n14469), .B(n14468), .Z(n14471) );
  NANDN U15066 ( .A(n14470), .B(n14471), .Z(n14473) );
  NAND U15067 ( .A(a[22]), .B(b[19]), .Z(n14857) );
  XNOR U15068 ( .A(n14471), .B(n14470), .Z(n14858) );
  NANDN U15069 ( .A(n14857), .B(n14858), .Z(n14472) );
  NAND U15070 ( .A(n14473), .B(n14472), .Z(n14474) );
  OR U15071 ( .A(n14475), .B(n14474), .Z(n14479) );
  XNOR U15072 ( .A(n14475), .B(n14474), .Z(n14861) );
  XOR U15073 ( .A(n14477), .B(n14476), .Z(n14862) );
  NANDN U15074 ( .A(n14861), .B(n14862), .Z(n14478) );
  NAND U15075 ( .A(n14479), .B(n14478), .Z(n14482) );
  XOR U15076 ( .A(n14481), .B(n14480), .Z(n14483) );
  NANDN U15077 ( .A(n14482), .B(n14483), .Z(n14485) );
  NAND U15078 ( .A(a[24]), .B(b[19]), .Z(n14869) );
  XNOR U15079 ( .A(n14483), .B(n14482), .Z(n14870) );
  NANDN U15080 ( .A(n14869), .B(n14870), .Z(n14484) );
  NAND U15081 ( .A(n14485), .B(n14484), .Z(n14486) );
  OR U15082 ( .A(n14487), .B(n14486), .Z(n14491) );
  XNOR U15083 ( .A(n14487), .B(n14486), .Z(n14873) );
  XOR U15084 ( .A(n14489), .B(n14488), .Z(n14874) );
  NANDN U15085 ( .A(n14873), .B(n14874), .Z(n14490) );
  NAND U15086 ( .A(n14491), .B(n14490), .Z(n14494) );
  XOR U15087 ( .A(n14493), .B(n14492), .Z(n14495) );
  NANDN U15088 ( .A(n14494), .B(n14495), .Z(n14497) );
  NAND U15089 ( .A(a[26]), .B(b[19]), .Z(n14881) );
  XNOR U15090 ( .A(n14495), .B(n14494), .Z(n14882) );
  NANDN U15091 ( .A(n14881), .B(n14882), .Z(n14496) );
  NAND U15092 ( .A(n14497), .B(n14496), .Z(n14498) );
  OR U15093 ( .A(n14499), .B(n14498), .Z(n14503) );
  XNOR U15094 ( .A(n14499), .B(n14498), .Z(n14885) );
  XOR U15095 ( .A(n14501), .B(n14500), .Z(n14886) );
  NANDN U15096 ( .A(n14885), .B(n14886), .Z(n14502) );
  NAND U15097 ( .A(n14503), .B(n14502), .Z(n14506) );
  XOR U15098 ( .A(n14505), .B(n14504), .Z(n14507) );
  NANDN U15099 ( .A(n14506), .B(n14507), .Z(n14509) );
  NAND U15100 ( .A(a[28]), .B(b[19]), .Z(n14893) );
  XNOR U15101 ( .A(n14507), .B(n14506), .Z(n14894) );
  NANDN U15102 ( .A(n14893), .B(n14894), .Z(n14508) );
  NAND U15103 ( .A(n14509), .B(n14508), .Z(n14510) );
  OR U15104 ( .A(n14511), .B(n14510), .Z(n14515) );
  XNOR U15105 ( .A(n14511), .B(n14510), .Z(n14897) );
  XOR U15106 ( .A(n14513), .B(n14512), .Z(n14898) );
  NANDN U15107 ( .A(n14897), .B(n14898), .Z(n14514) );
  NAND U15108 ( .A(n14515), .B(n14514), .Z(n14518) );
  XOR U15109 ( .A(n14517), .B(n14516), .Z(n14519) );
  NANDN U15110 ( .A(n14518), .B(n14519), .Z(n14521) );
  NAND U15111 ( .A(a[30]), .B(b[19]), .Z(n14905) );
  XNOR U15112 ( .A(n14519), .B(n14518), .Z(n14906) );
  NANDN U15113 ( .A(n14905), .B(n14906), .Z(n14520) );
  NAND U15114 ( .A(n14521), .B(n14520), .Z(n14522) );
  OR U15115 ( .A(n14523), .B(n14522), .Z(n14527) );
  XNOR U15116 ( .A(n14523), .B(n14522), .Z(n14909) );
  XOR U15117 ( .A(n14525), .B(n14524), .Z(n14910) );
  NANDN U15118 ( .A(n14909), .B(n14910), .Z(n14526) );
  NAND U15119 ( .A(n14527), .B(n14526), .Z(n14530) );
  XOR U15120 ( .A(n14529), .B(n14528), .Z(n14531) );
  NANDN U15121 ( .A(n14530), .B(n14531), .Z(n14533) );
  NAND U15122 ( .A(a[32]), .B(b[19]), .Z(n14917) );
  XNOR U15123 ( .A(n14531), .B(n14530), .Z(n14918) );
  NANDN U15124 ( .A(n14917), .B(n14918), .Z(n14532) );
  NAND U15125 ( .A(n14533), .B(n14532), .Z(n14534) );
  OR U15126 ( .A(n14535), .B(n14534), .Z(n14539) );
  XNOR U15127 ( .A(n14535), .B(n14534), .Z(n14921) );
  XOR U15128 ( .A(n14537), .B(n14536), .Z(n14922) );
  NANDN U15129 ( .A(n14921), .B(n14922), .Z(n14538) );
  NAND U15130 ( .A(n14539), .B(n14538), .Z(n14542) );
  XOR U15131 ( .A(n14541), .B(n14540), .Z(n14543) );
  NANDN U15132 ( .A(n14542), .B(n14543), .Z(n14545) );
  NAND U15133 ( .A(a[34]), .B(b[19]), .Z(n14929) );
  XNOR U15134 ( .A(n14543), .B(n14542), .Z(n14930) );
  NANDN U15135 ( .A(n14929), .B(n14930), .Z(n14544) );
  NAND U15136 ( .A(n14545), .B(n14544), .Z(n14546) );
  OR U15137 ( .A(n14547), .B(n14546), .Z(n14551) );
  XNOR U15138 ( .A(n14547), .B(n14546), .Z(n14933) );
  XOR U15139 ( .A(n14549), .B(n14548), .Z(n14934) );
  NANDN U15140 ( .A(n14933), .B(n14934), .Z(n14550) );
  NAND U15141 ( .A(n14551), .B(n14550), .Z(n14554) );
  XOR U15142 ( .A(n14553), .B(n14552), .Z(n14555) );
  NANDN U15143 ( .A(n14554), .B(n14555), .Z(n14557) );
  NAND U15144 ( .A(a[36]), .B(b[19]), .Z(n14941) );
  XNOR U15145 ( .A(n14555), .B(n14554), .Z(n14942) );
  NANDN U15146 ( .A(n14941), .B(n14942), .Z(n14556) );
  NAND U15147 ( .A(n14557), .B(n14556), .Z(n14558) );
  OR U15148 ( .A(n14559), .B(n14558), .Z(n14563) );
  XNOR U15149 ( .A(n14559), .B(n14558), .Z(n14945) );
  XOR U15150 ( .A(n14561), .B(n14560), .Z(n14946) );
  NANDN U15151 ( .A(n14945), .B(n14946), .Z(n14562) );
  NAND U15152 ( .A(n14563), .B(n14562), .Z(n14566) );
  XOR U15153 ( .A(n14565), .B(n14564), .Z(n14567) );
  NANDN U15154 ( .A(n14566), .B(n14567), .Z(n14569) );
  NAND U15155 ( .A(a[38]), .B(b[19]), .Z(n14953) );
  XNOR U15156 ( .A(n14567), .B(n14566), .Z(n14954) );
  NANDN U15157 ( .A(n14953), .B(n14954), .Z(n14568) );
  NAND U15158 ( .A(n14569), .B(n14568), .Z(n14570) );
  OR U15159 ( .A(n14571), .B(n14570), .Z(n14575) );
  XNOR U15160 ( .A(n14571), .B(n14570), .Z(n14957) );
  XOR U15161 ( .A(n14573), .B(n14572), .Z(n14958) );
  NANDN U15162 ( .A(n14957), .B(n14958), .Z(n14574) );
  NAND U15163 ( .A(n14575), .B(n14574), .Z(n14578) );
  XOR U15164 ( .A(n14577), .B(n14576), .Z(n14579) );
  NANDN U15165 ( .A(n14578), .B(n14579), .Z(n14581) );
  NAND U15166 ( .A(a[40]), .B(b[19]), .Z(n14965) );
  XNOR U15167 ( .A(n14579), .B(n14578), .Z(n14966) );
  NANDN U15168 ( .A(n14965), .B(n14966), .Z(n14580) );
  NAND U15169 ( .A(n14581), .B(n14580), .Z(n14582) );
  OR U15170 ( .A(n14583), .B(n14582), .Z(n14587) );
  XNOR U15171 ( .A(n14583), .B(n14582), .Z(n14969) );
  XOR U15172 ( .A(n14585), .B(n14584), .Z(n14970) );
  NANDN U15173 ( .A(n14969), .B(n14970), .Z(n14586) );
  NAND U15174 ( .A(n14587), .B(n14586), .Z(n14590) );
  XOR U15175 ( .A(n14589), .B(n14588), .Z(n14591) );
  NANDN U15176 ( .A(n14590), .B(n14591), .Z(n14593) );
  NAND U15177 ( .A(a[42]), .B(b[19]), .Z(n14977) );
  XNOR U15178 ( .A(n14591), .B(n14590), .Z(n14978) );
  NANDN U15179 ( .A(n14977), .B(n14978), .Z(n14592) );
  NAND U15180 ( .A(n14593), .B(n14592), .Z(n14596) );
  ANDN U15181 ( .B(b[19]), .A(n191), .Z(n14597) );
  OR U15182 ( .A(n14596), .B(n14597), .Z(n14599) );
  XOR U15183 ( .A(n14595), .B(n14594), .Z(n14982) );
  XOR U15184 ( .A(n14597), .B(n14596), .Z(n14981) );
  NANDN U15185 ( .A(n14982), .B(n14981), .Z(n14598) );
  NAND U15186 ( .A(n14599), .B(n14598), .Z(n14602) );
  XNOR U15187 ( .A(n14601), .B(n14600), .Z(n14603) );
  OR U15188 ( .A(n14602), .B(n14603), .Z(n14605) );
  XNOR U15189 ( .A(n14603), .B(n14602), .Z(n14988) );
  NAND U15190 ( .A(a[44]), .B(b[19]), .Z(n14987) );
  OR U15191 ( .A(n14988), .B(n14987), .Z(n14604) );
  NAND U15192 ( .A(n14605), .B(n14604), .Z(n14606) );
  ANDN U15193 ( .B(b[19]), .A(n193), .Z(n14607) );
  OR U15194 ( .A(n14606), .B(n14607), .Z(n14611) );
  XOR U15195 ( .A(n14607), .B(n14606), .Z(n14993) );
  NAND U15196 ( .A(n14993), .B(n14994), .Z(n14610) );
  NAND U15197 ( .A(n14611), .B(n14610), .Z(n14615) );
  NAND U15198 ( .A(a[46]), .B(b[19]), .Z(n14614) );
  OR U15199 ( .A(n14615), .B(n14614), .Z(n14617) );
  XOR U15200 ( .A(n14613), .B(n14612), .Z(n14999) );
  XOR U15201 ( .A(n14615), .B(n14614), .Z(n15000) );
  NAND U15202 ( .A(n14999), .B(n15000), .Z(n14616) );
  NAND U15203 ( .A(n14617), .B(n14616), .Z(n14621) );
  XOR U15204 ( .A(n14619), .B(n14618), .Z(n14620) );
  NAND U15205 ( .A(n14621), .B(n14620), .Z(n14623) );
  XNOR U15206 ( .A(n14621), .B(n14620), .Z(n15006) );
  NAND U15207 ( .A(a[47]), .B(b[19]), .Z(n15005) );
  OR U15208 ( .A(n15006), .B(n15005), .Z(n14622) );
  NAND U15209 ( .A(n14623), .B(n14622), .Z(n14627) );
  NANDN U15210 ( .A(n14626), .B(n14627), .Z(n14629) );
  XNOR U15211 ( .A(n14625), .B(n14624), .Z(n15012) );
  XNOR U15212 ( .A(n14627), .B(n14626), .Z(n15011) );
  NANDN U15213 ( .A(n15012), .B(n15011), .Z(n14628) );
  NAND U15214 ( .A(n14629), .B(n14628), .Z(n14633) );
  XOR U15215 ( .A(n14631), .B(n14630), .Z(n14632) );
  NAND U15216 ( .A(n14633), .B(n14632), .Z(n14635) );
  XNOR U15217 ( .A(n14633), .B(n14632), .Z(n15018) );
  NAND U15218 ( .A(a[49]), .B(b[19]), .Z(n15017) );
  OR U15219 ( .A(n15018), .B(n15017), .Z(n14634) );
  NAND U15220 ( .A(n14635), .B(n14634), .Z(n14639) );
  NANDN U15221 ( .A(n14638), .B(n14639), .Z(n14641) );
  XNOR U15222 ( .A(n14637), .B(n14636), .Z(n15024) );
  XNOR U15223 ( .A(n14639), .B(n14638), .Z(n15023) );
  NANDN U15224 ( .A(n15024), .B(n15023), .Z(n14640) );
  NAND U15225 ( .A(n14641), .B(n14640), .Z(n14645) );
  XOR U15226 ( .A(n14643), .B(n14642), .Z(n14644) );
  NAND U15227 ( .A(n14645), .B(n14644), .Z(n14647) );
  XNOR U15228 ( .A(n14645), .B(n14644), .Z(n15030) );
  NAND U15229 ( .A(a[51]), .B(b[19]), .Z(n15029) );
  OR U15230 ( .A(n15030), .B(n15029), .Z(n14646) );
  NAND U15231 ( .A(n14647), .B(n14646), .Z(n14651) );
  NANDN U15232 ( .A(n14650), .B(n14651), .Z(n14653) );
  XNOR U15233 ( .A(n14649), .B(n14648), .Z(n15036) );
  XNOR U15234 ( .A(n14651), .B(n14650), .Z(n15035) );
  NANDN U15235 ( .A(n15036), .B(n15035), .Z(n14652) );
  NAND U15236 ( .A(n14653), .B(n14652), .Z(n14657) );
  XOR U15237 ( .A(n14655), .B(n14654), .Z(n14656) );
  NAND U15238 ( .A(n14657), .B(n14656), .Z(n14659) );
  XNOR U15239 ( .A(n14657), .B(n14656), .Z(n15042) );
  NAND U15240 ( .A(a[53]), .B(b[19]), .Z(n15041) );
  OR U15241 ( .A(n15042), .B(n15041), .Z(n14658) );
  NAND U15242 ( .A(n14659), .B(n14658), .Z(n14663) );
  NANDN U15243 ( .A(n14662), .B(n14663), .Z(n14665) );
  XNOR U15244 ( .A(n14661), .B(n14660), .Z(n15048) );
  XNOR U15245 ( .A(n14663), .B(n14662), .Z(n15047) );
  NANDN U15246 ( .A(n15048), .B(n15047), .Z(n14664) );
  NAND U15247 ( .A(n14665), .B(n14664), .Z(n14669) );
  XOR U15248 ( .A(n14667), .B(n14666), .Z(n14668) );
  NAND U15249 ( .A(n14669), .B(n14668), .Z(n14671) );
  XNOR U15250 ( .A(n14669), .B(n14668), .Z(n15054) );
  NAND U15251 ( .A(a[55]), .B(b[19]), .Z(n15053) );
  OR U15252 ( .A(n15054), .B(n15053), .Z(n14670) );
  NAND U15253 ( .A(n14671), .B(n14670), .Z(n14675) );
  NANDN U15254 ( .A(n14674), .B(n14675), .Z(n14677) );
  XNOR U15255 ( .A(n14673), .B(n14672), .Z(n15060) );
  XNOR U15256 ( .A(n14675), .B(n14674), .Z(n15059) );
  NANDN U15257 ( .A(n15060), .B(n15059), .Z(n14676) );
  NAND U15258 ( .A(n14677), .B(n14676), .Z(n14681) );
  XOR U15259 ( .A(n14679), .B(n14678), .Z(n14680) );
  NAND U15260 ( .A(n14681), .B(n14680), .Z(n14683) );
  XNOR U15261 ( .A(n14681), .B(n14680), .Z(n15066) );
  NAND U15262 ( .A(a[57]), .B(b[19]), .Z(n15065) );
  OR U15263 ( .A(n15066), .B(n15065), .Z(n14682) );
  NAND U15264 ( .A(n14683), .B(n14682), .Z(n14687) );
  NANDN U15265 ( .A(n14686), .B(n14687), .Z(n14689) );
  XNOR U15266 ( .A(n14685), .B(n14684), .Z(n15072) );
  XNOR U15267 ( .A(n14687), .B(n14686), .Z(n15071) );
  NANDN U15268 ( .A(n15072), .B(n15071), .Z(n14688) );
  NAND U15269 ( .A(n14689), .B(n14688), .Z(n14692) );
  XOR U15270 ( .A(n14691), .B(n14690), .Z(n14693) );
  OR U15271 ( .A(n14692), .B(n14693), .Z(n14695) );
  AND U15272 ( .A(b[19]), .B(a[59]), .Z(n15078) );
  XOR U15273 ( .A(n14693), .B(n14692), .Z(n15077) );
  NANDN U15274 ( .A(n15078), .B(n15077), .Z(n14694) );
  NAND U15275 ( .A(n14695), .B(n14694), .Z(n14699) );
  NAND U15276 ( .A(a[60]), .B(b[19]), .Z(n14698) );
  OR U15277 ( .A(n14699), .B(n14698), .Z(n14701) );
  XNOR U15278 ( .A(n14697), .B(n14696), .Z(n15084) );
  XOR U15279 ( .A(n14699), .B(n14698), .Z(n15083) );
  NANDN U15280 ( .A(n15084), .B(n15083), .Z(n14700) );
  NAND U15281 ( .A(n14701), .B(n14700), .Z(n14705) );
  XOR U15282 ( .A(n14703), .B(n14702), .Z(n14704) );
  NAND U15283 ( .A(n14705), .B(n14704), .Z(n14707) );
  XNOR U15284 ( .A(n14705), .B(n14704), .Z(n15090) );
  NAND U15285 ( .A(a[61]), .B(b[19]), .Z(n15089) );
  OR U15286 ( .A(n15090), .B(n15089), .Z(n14706) );
  NAND U15287 ( .A(n14707), .B(n14706), .Z(n14711) );
  NANDN U15288 ( .A(n14710), .B(n14711), .Z(n14713) );
  XOR U15289 ( .A(n14709), .B(n14708), .Z(n15096) );
  XNOR U15290 ( .A(n14711), .B(n14710), .Z(n15095) );
  NAND U15291 ( .A(n15096), .B(n15095), .Z(n14712) );
  NAND U15292 ( .A(n14713), .B(n14712), .Z(n14725) );
  XOR U15293 ( .A(n14715), .B(n14714), .Z(n14724) );
  NAND U15294 ( .A(n14725), .B(n14724), .Z(n14716) );
  AND U15295 ( .A(n14717), .B(n14716), .Z(n14722) );
  XNOR U15296 ( .A(n14719), .B(n14718), .Z(n14723) );
  NANDN U15297 ( .A(n14722), .B(n14723), .Z(n24161) );
  XOR U15298 ( .A(n14721), .B(n14720), .Z(n24158) );
  XNOR U15299 ( .A(n14723), .B(n14722), .Z(n24154) );
  XOR U15300 ( .A(n14725), .B(n14724), .Z(n15102) );
  NAND U15301 ( .A(a[48]), .B(b[18]), .Z(n15007) );
  ANDN U15302 ( .B(b[18]), .A(n191), .Z(n14976) );
  ANDN U15303 ( .B(b[18]), .A(n189), .Z(n14964) );
  ANDN U15304 ( .B(b[18]), .A(n187), .Z(n14952) );
  ANDN U15305 ( .B(b[18]), .A(n21772), .Z(n14940) );
  ANDN U15306 ( .B(b[18]), .A(n184), .Z(n14928) );
  ANDN U15307 ( .B(b[18]), .A(n21751), .Z(n14916) );
  ANDN U15308 ( .B(b[18]), .A(n21740), .Z(n14904) );
  ANDN U15309 ( .B(b[18]), .A(n21727), .Z(n14892) );
  ANDN U15310 ( .B(b[18]), .A(n21716), .Z(n14880) );
  ANDN U15311 ( .B(b[18]), .A(n21703), .Z(n14868) );
  ANDN U15312 ( .B(b[18]), .A(n21692), .Z(n14856) );
  ANDN U15313 ( .B(b[18]), .A(n21681), .Z(n14844) );
  ANDN U15314 ( .B(b[18]), .A(n21670), .Z(n14832) );
  NAND U15315 ( .A(a[17]), .B(b[18]), .Z(n14820) );
  ANDN U15316 ( .B(b[18]), .A(n172), .Z(n14809) );
  ANDN U15317 ( .B(b[18]), .A(n170), .Z(n14798) );
  ANDN U15318 ( .B(b[18]), .A(n21164), .Z(n14786) );
  ANDN U15319 ( .B(b[18]), .A(n21615), .Z(n14774) );
  ANDN U15320 ( .B(b[18]), .A(n166), .Z(n14762) );
  NAND U15321 ( .A(a[6]), .B(b[18]), .Z(n14757) );
  XOR U15322 ( .A(n14729), .B(n14728), .Z(n14758) );
  NANDN U15323 ( .A(n14757), .B(n14758), .Z(n14760) );
  ANDN U15324 ( .B(b[18]), .A(n164), .Z(n14752) );
  ANDN U15325 ( .B(b[18]), .A(n21580), .Z(n14739) );
  NAND U15326 ( .A(b[19]), .B(a[1]), .Z(n14732) );
  AND U15327 ( .A(b[18]), .B(a[0]), .Z(n15496) );
  NANDN U15328 ( .A(n14732), .B(n15496), .Z(n14731) );
  NAND U15329 ( .A(a[2]), .B(b[18]), .Z(n14730) );
  AND U15330 ( .A(n14731), .B(n14730), .Z(n14738) );
  NANDN U15331 ( .A(n14732), .B(a[0]), .Z(n14733) );
  XNOR U15332 ( .A(a[2]), .B(n14733), .Z(n14734) );
  NAND U15333 ( .A(b[18]), .B(n14734), .Z(n15123) );
  AND U15334 ( .A(a[1]), .B(b[19]), .Z(n14735) );
  XNOR U15335 ( .A(n14736), .B(n14735), .Z(n15122) );
  NANDN U15336 ( .A(n15123), .B(n15122), .Z(n14737) );
  NANDN U15337 ( .A(n14738), .B(n14737), .Z(n14740) );
  NANDN U15338 ( .A(n14739), .B(n14740), .Z(n14744) );
  XOR U15339 ( .A(n14740), .B(n14739), .Z(n15127) );
  NANDN U15340 ( .A(n15127), .B(n15126), .Z(n14743) );
  NAND U15341 ( .A(n14744), .B(n14743), .Z(n14748) );
  XOR U15342 ( .A(n14746), .B(n14745), .Z(n14747) );
  NANDN U15343 ( .A(n14748), .B(n14747), .Z(n14750) );
  NAND U15344 ( .A(a[4]), .B(b[18]), .Z(n15134) );
  NANDN U15345 ( .A(n15134), .B(n15135), .Z(n14749) );
  NAND U15346 ( .A(n14750), .B(n14749), .Z(n14751) );
  OR U15347 ( .A(n14752), .B(n14751), .Z(n14756) );
  XNOR U15348 ( .A(n14752), .B(n14751), .Z(n15109) );
  XOR U15349 ( .A(n14754), .B(n14753), .Z(n15110) );
  NANDN U15350 ( .A(n15109), .B(n15110), .Z(n14755) );
  NAND U15351 ( .A(n14756), .B(n14755), .Z(n15144) );
  XNOR U15352 ( .A(n14758), .B(n14757), .Z(n15145) );
  NANDN U15353 ( .A(n15144), .B(n15145), .Z(n14759) );
  NAND U15354 ( .A(n14760), .B(n14759), .Z(n14761) );
  OR U15355 ( .A(n14762), .B(n14761), .Z(n14766) );
  XNOR U15356 ( .A(n14762), .B(n14761), .Z(n15148) );
  XOR U15357 ( .A(n14764), .B(n14763), .Z(n15149) );
  NANDN U15358 ( .A(n15148), .B(n15149), .Z(n14765) );
  NAND U15359 ( .A(n14766), .B(n14765), .Z(n14769) );
  XOR U15360 ( .A(n14768), .B(n14767), .Z(n14770) );
  NANDN U15361 ( .A(n14769), .B(n14770), .Z(n14772) );
  NAND U15362 ( .A(a[8]), .B(b[18]), .Z(n15156) );
  XNOR U15363 ( .A(n14770), .B(n14769), .Z(n15157) );
  NANDN U15364 ( .A(n15156), .B(n15157), .Z(n14771) );
  NAND U15365 ( .A(n14772), .B(n14771), .Z(n14773) );
  OR U15366 ( .A(n14774), .B(n14773), .Z(n14778) );
  XOR U15367 ( .A(n14774), .B(n14773), .Z(n15160) );
  XOR U15368 ( .A(n14776), .B(n14775), .Z(n15161) );
  NAND U15369 ( .A(n15160), .B(n15161), .Z(n14777) );
  NAND U15370 ( .A(n14778), .B(n14777), .Z(n14781) );
  NANDN U15371 ( .A(n14781), .B(n14782), .Z(n14784) );
  NAND U15372 ( .A(a[10]), .B(b[18]), .Z(n15168) );
  XNOR U15373 ( .A(n14782), .B(n14781), .Z(n15169) );
  NANDN U15374 ( .A(n15168), .B(n15169), .Z(n14783) );
  NAND U15375 ( .A(n14784), .B(n14783), .Z(n14785) );
  OR U15376 ( .A(n14786), .B(n14785), .Z(n14790) );
  XNOR U15377 ( .A(n14786), .B(n14785), .Z(n15172) );
  XOR U15378 ( .A(n14788), .B(n14787), .Z(n15173) );
  NANDN U15379 ( .A(n15172), .B(n15173), .Z(n14789) );
  NAND U15380 ( .A(n14790), .B(n14789), .Z(n14794) );
  XOR U15381 ( .A(n14792), .B(n14791), .Z(n14793) );
  NANDN U15382 ( .A(n14794), .B(n14793), .Z(n14796) );
  NAND U15383 ( .A(a[12]), .B(b[18]), .Z(n15180) );
  NANDN U15384 ( .A(n15180), .B(n15181), .Z(n14795) );
  NAND U15385 ( .A(n14796), .B(n14795), .Z(n14797) );
  OR U15386 ( .A(n14798), .B(n14797), .Z(n14802) );
  XNOR U15387 ( .A(n14798), .B(n14797), .Z(n15184) );
  XOR U15388 ( .A(n14800), .B(n14799), .Z(n15185) );
  NANDN U15389 ( .A(n15184), .B(n15185), .Z(n14801) );
  NAND U15390 ( .A(n14802), .B(n14801), .Z(n14806) );
  NAND U15391 ( .A(n14806), .B(n14805), .Z(n14808) );
  ANDN U15392 ( .B(b[18]), .A(n171), .Z(n15191) );
  XNOR U15393 ( .A(n14806), .B(n14805), .Z(n15190) );
  OR U15394 ( .A(n15191), .B(n15190), .Z(n14807) );
  NAND U15395 ( .A(n14808), .B(n14807), .Z(n14810) );
  NANDN U15396 ( .A(n14809), .B(n14810), .Z(n14814) );
  XOR U15397 ( .A(n14810), .B(n14809), .Z(n15108) );
  XOR U15398 ( .A(n14812), .B(n14811), .Z(n15107) );
  NANDN U15399 ( .A(n15108), .B(n15107), .Z(n14813) );
  AND U15400 ( .A(n14814), .B(n14813), .Z(n14815) );
  OR U15401 ( .A(n14816), .B(n14815), .Z(n14818) );
  ANDN U15402 ( .B(b[18]), .A(n173), .Z(n15203) );
  XNOR U15403 ( .A(n14816), .B(n14815), .Z(n15202) );
  OR U15404 ( .A(n15203), .B(n15202), .Z(n14817) );
  AND U15405 ( .A(n14818), .B(n14817), .Z(n14819) );
  NANDN U15406 ( .A(n14820), .B(n14819), .Z(n14824) );
  XNOR U15407 ( .A(n14822), .B(n14821), .Z(n15106) );
  NAND U15408 ( .A(n15105), .B(n15106), .Z(n14823) );
  AND U15409 ( .A(n14824), .B(n14823), .Z(n14827) );
  XOR U15410 ( .A(n14826), .B(n14825), .Z(n14828) );
  NANDN U15411 ( .A(n14827), .B(n14828), .Z(n14830) );
  NAND U15412 ( .A(a[18]), .B(b[18]), .Z(n15212) );
  XNOR U15413 ( .A(n14828), .B(n14827), .Z(n15213) );
  NANDN U15414 ( .A(n15212), .B(n15213), .Z(n14829) );
  NAND U15415 ( .A(n14830), .B(n14829), .Z(n14831) );
  OR U15416 ( .A(n14832), .B(n14831), .Z(n14836) );
  XNOR U15417 ( .A(n14832), .B(n14831), .Z(n15216) );
  XOR U15418 ( .A(n14834), .B(n14833), .Z(n15217) );
  NANDN U15419 ( .A(n15216), .B(n15217), .Z(n14835) );
  NAND U15420 ( .A(n14836), .B(n14835), .Z(n14839) );
  XOR U15421 ( .A(n14838), .B(n14837), .Z(n14840) );
  NANDN U15422 ( .A(n14839), .B(n14840), .Z(n14842) );
  NAND U15423 ( .A(a[20]), .B(b[18]), .Z(n15224) );
  XNOR U15424 ( .A(n14840), .B(n14839), .Z(n15225) );
  NANDN U15425 ( .A(n15224), .B(n15225), .Z(n14841) );
  NAND U15426 ( .A(n14842), .B(n14841), .Z(n14843) );
  OR U15427 ( .A(n14844), .B(n14843), .Z(n14848) );
  XNOR U15428 ( .A(n14844), .B(n14843), .Z(n15228) );
  XOR U15429 ( .A(n14846), .B(n14845), .Z(n15229) );
  NANDN U15430 ( .A(n15228), .B(n15229), .Z(n14847) );
  NAND U15431 ( .A(n14848), .B(n14847), .Z(n14851) );
  XOR U15432 ( .A(n14850), .B(n14849), .Z(n14852) );
  NANDN U15433 ( .A(n14851), .B(n14852), .Z(n14854) );
  NAND U15434 ( .A(a[22]), .B(b[18]), .Z(n15236) );
  XNOR U15435 ( .A(n14852), .B(n14851), .Z(n15237) );
  NANDN U15436 ( .A(n15236), .B(n15237), .Z(n14853) );
  NAND U15437 ( .A(n14854), .B(n14853), .Z(n14855) );
  OR U15438 ( .A(n14856), .B(n14855), .Z(n14860) );
  XNOR U15439 ( .A(n14856), .B(n14855), .Z(n15240) );
  XOR U15440 ( .A(n14858), .B(n14857), .Z(n15241) );
  NANDN U15441 ( .A(n15240), .B(n15241), .Z(n14859) );
  NAND U15442 ( .A(n14860), .B(n14859), .Z(n14863) );
  XOR U15443 ( .A(n14862), .B(n14861), .Z(n14864) );
  NANDN U15444 ( .A(n14863), .B(n14864), .Z(n14866) );
  NAND U15445 ( .A(a[24]), .B(b[18]), .Z(n15248) );
  XNOR U15446 ( .A(n14864), .B(n14863), .Z(n15249) );
  NANDN U15447 ( .A(n15248), .B(n15249), .Z(n14865) );
  NAND U15448 ( .A(n14866), .B(n14865), .Z(n14867) );
  OR U15449 ( .A(n14868), .B(n14867), .Z(n14872) );
  XNOR U15450 ( .A(n14868), .B(n14867), .Z(n15252) );
  XOR U15451 ( .A(n14870), .B(n14869), .Z(n15253) );
  NANDN U15452 ( .A(n15252), .B(n15253), .Z(n14871) );
  NAND U15453 ( .A(n14872), .B(n14871), .Z(n14875) );
  XOR U15454 ( .A(n14874), .B(n14873), .Z(n14876) );
  NANDN U15455 ( .A(n14875), .B(n14876), .Z(n14878) );
  NAND U15456 ( .A(a[26]), .B(b[18]), .Z(n15260) );
  XNOR U15457 ( .A(n14876), .B(n14875), .Z(n15261) );
  NANDN U15458 ( .A(n15260), .B(n15261), .Z(n14877) );
  NAND U15459 ( .A(n14878), .B(n14877), .Z(n14879) );
  OR U15460 ( .A(n14880), .B(n14879), .Z(n14884) );
  XNOR U15461 ( .A(n14880), .B(n14879), .Z(n15264) );
  XOR U15462 ( .A(n14882), .B(n14881), .Z(n15265) );
  NANDN U15463 ( .A(n15264), .B(n15265), .Z(n14883) );
  NAND U15464 ( .A(n14884), .B(n14883), .Z(n14887) );
  XOR U15465 ( .A(n14886), .B(n14885), .Z(n14888) );
  NANDN U15466 ( .A(n14887), .B(n14888), .Z(n14890) );
  NAND U15467 ( .A(a[28]), .B(b[18]), .Z(n15272) );
  XNOR U15468 ( .A(n14888), .B(n14887), .Z(n15273) );
  NANDN U15469 ( .A(n15272), .B(n15273), .Z(n14889) );
  NAND U15470 ( .A(n14890), .B(n14889), .Z(n14891) );
  OR U15471 ( .A(n14892), .B(n14891), .Z(n14896) );
  XNOR U15472 ( .A(n14892), .B(n14891), .Z(n15276) );
  XOR U15473 ( .A(n14894), .B(n14893), .Z(n15277) );
  NANDN U15474 ( .A(n15276), .B(n15277), .Z(n14895) );
  NAND U15475 ( .A(n14896), .B(n14895), .Z(n14899) );
  XOR U15476 ( .A(n14898), .B(n14897), .Z(n14900) );
  NANDN U15477 ( .A(n14899), .B(n14900), .Z(n14902) );
  NAND U15478 ( .A(a[30]), .B(b[18]), .Z(n15284) );
  XNOR U15479 ( .A(n14900), .B(n14899), .Z(n15285) );
  NANDN U15480 ( .A(n15284), .B(n15285), .Z(n14901) );
  NAND U15481 ( .A(n14902), .B(n14901), .Z(n14903) );
  OR U15482 ( .A(n14904), .B(n14903), .Z(n14908) );
  XNOR U15483 ( .A(n14904), .B(n14903), .Z(n15288) );
  XOR U15484 ( .A(n14906), .B(n14905), .Z(n15289) );
  NANDN U15485 ( .A(n15288), .B(n15289), .Z(n14907) );
  NAND U15486 ( .A(n14908), .B(n14907), .Z(n14911) );
  XOR U15487 ( .A(n14910), .B(n14909), .Z(n14912) );
  NANDN U15488 ( .A(n14911), .B(n14912), .Z(n14914) );
  NAND U15489 ( .A(a[32]), .B(b[18]), .Z(n15296) );
  XNOR U15490 ( .A(n14912), .B(n14911), .Z(n15297) );
  NANDN U15491 ( .A(n15296), .B(n15297), .Z(n14913) );
  NAND U15492 ( .A(n14914), .B(n14913), .Z(n14915) );
  OR U15493 ( .A(n14916), .B(n14915), .Z(n14920) );
  XNOR U15494 ( .A(n14916), .B(n14915), .Z(n15300) );
  XOR U15495 ( .A(n14918), .B(n14917), .Z(n15301) );
  NANDN U15496 ( .A(n15300), .B(n15301), .Z(n14919) );
  NAND U15497 ( .A(n14920), .B(n14919), .Z(n14923) );
  XOR U15498 ( .A(n14922), .B(n14921), .Z(n14924) );
  NANDN U15499 ( .A(n14923), .B(n14924), .Z(n14926) );
  NAND U15500 ( .A(a[34]), .B(b[18]), .Z(n15308) );
  XNOR U15501 ( .A(n14924), .B(n14923), .Z(n15309) );
  NANDN U15502 ( .A(n15308), .B(n15309), .Z(n14925) );
  NAND U15503 ( .A(n14926), .B(n14925), .Z(n14927) );
  OR U15504 ( .A(n14928), .B(n14927), .Z(n14932) );
  XNOR U15505 ( .A(n14928), .B(n14927), .Z(n15312) );
  XOR U15506 ( .A(n14930), .B(n14929), .Z(n15313) );
  NANDN U15507 ( .A(n15312), .B(n15313), .Z(n14931) );
  NAND U15508 ( .A(n14932), .B(n14931), .Z(n14935) );
  XOR U15509 ( .A(n14934), .B(n14933), .Z(n14936) );
  NANDN U15510 ( .A(n14935), .B(n14936), .Z(n14938) );
  NAND U15511 ( .A(a[36]), .B(b[18]), .Z(n15320) );
  XNOR U15512 ( .A(n14936), .B(n14935), .Z(n15321) );
  NANDN U15513 ( .A(n15320), .B(n15321), .Z(n14937) );
  NAND U15514 ( .A(n14938), .B(n14937), .Z(n14939) );
  OR U15515 ( .A(n14940), .B(n14939), .Z(n14944) );
  XNOR U15516 ( .A(n14940), .B(n14939), .Z(n15324) );
  XOR U15517 ( .A(n14942), .B(n14941), .Z(n15325) );
  NANDN U15518 ( .A(n15324), .B(n15325), .Z(n14943) );
  NAND U15519 ( .A(n14944), .B(n14943), .Z(n14947) );
  XOR U15520 ( .A(n14946), .B(n14945), .Z(n14948) );
  NANDN U15521 ( .A(n14947), .B(n14948), .Z(n14950) );
  NAND U15522 ( .A(a[38]), .B(b[18]), .Z(n15332) );
  XNOR U15523 ( .A(n14948), .B(n14947), .Z(n15333) );
  NANDN U15524 ( .A(n15332), .B(n15333), .Z(n14949) );
  NAND U15525 ( .A(n14950), .B(n14949), .Z(n14951) );
  OR U15526 ( .A(n14952), .B(n14951), .Z(n14956) );
  XNOR U15527 ( .A(n14952), .B(n14951), .Z(n15336) );
  XOR U15528 ( .A(n14954), .B(n14953), .Z(n15337) );
  NANDN U15529 ( .A(n15336), .B(n15337), .Z(n14955) );
  NAND U15530 ( .A(n14956), .B(n14955), .Z(n14959) );
  XOR U15531 ( .A(n14958), .B(n14957), .Z(n14960) );
  NANDN U15532 ( .A(n14959), .B(n14960), .Z(n14962) );
  NAND U15533 ( .A(a[40]), .B(b[18]), .Z(n15344) );
  XNOR U15534 ( .A(n14960), .B(n14959), .Z(n15345) );
  NANDN U15535 ( .A(n15344), .B(n15345), .Z(n14961) );
  NAND U15536 ( .A(n14962), .B(n14961), .Z(n14963) );
  OR U15537 ( .A(n14964), .B(n14963), .Z(n14968) );
  XNOR U15538 ( .A(n14964), .B(n14963), .Z(n15348) );
  XOR U15539 ( .A(n14966), .B(n14965), .Z(n15349) );
  NANDN U15540 ( .A(n15348), .B(n15349), .Z(n14967) );
  NAND U15541 ( .A(n14968), .B(n14967), .Z(n14971) );
  XOR U15542 ( .A(n14970), .B(n14969), .Z(n14972) );
  NANDN U15543 ( .A(n14971), .B(n14972), .Z(n14974) );
  NAND U15544 ( .A(a[42]), .B(b[18]), .Z(n15356) );
  XNOR U15545 ( .A(n14972), .B(n14971), .Z(n15357) );
  NANDN U15546 ( .A(n15356), .B(n15357), .Z(n14973) );
  NAND U15547 ( .A(n14974), .B(n14973), .Z(n14975) );
  OR U15548 ( .A(n14976), .B(n14975), .Z(n14980) );
  XNOR U15549 ( .A(n14976), .B(n14975), .Z(n15360) );
  XOR U15550 ( .A(n14978), .B(n14977), .Z(n15361) );
  NANDN U15551 ( .A(n15360), .B(n15361), .Z(n14979) );
  NAND U15552 ( .A(n14980), .B(n14979), .Z(n14983) );
  XNOR U15553 ( .A(n14982), .B(n14981), .Z(n14984) );
  OR U15554 ( .A(n14983), .B(n14984), .Z(n14986) );
  XNOR U15555 ( .A(n14984), .B(n14983), .Z(n15367) );
  NAND U15556 ( .A(a[44]), .B(b[18]), .Z(n15366) );
  OR U15557 ( .A(n15367), .B(n15366), .Z(n14985) );
  NAND U15558 ( .A(n14986), .B(n14985), .Z(n14989) );
  ANDN U15559 ( .B(b[18]), .A(n193), .Z(n14990) );
  OR U15560 ( .A(n14989), .B(n14990), .Z(n14992) );
  XOR U15561 ( .A(n14988), .B(n14987), .Z(n15373) );
  XOR U15562 ( .A(n14990), .B(n14989), .Z(n15372) );
  NANDN U15563 ( .A(n15373), .B(n15372), .Z(n14991) );
  NAND U15564 ( .A(n14992), .B(n14991), .Z(n14996) );
  AND U15565 ( .A(b[18]), .B(a[46]), .Z(n14995) );
  NANDN U15566 ( .A(n14996), .B(n14995), .Z(n14998) );
  XNOR U15567 ( .A(n14996), .B(n14995), .Z(n15380) );
  NANDN U15568 ( .A(n15381), .B(n15380), .Z(n14997) );
  NAND U15569 ( .A(n14998), .B(n14997), .Z(n15002) );
  XOR U15570 ( .A(n15000), .B(n14999), .Z(n15001) );
  NAND U15571 ( .A(n15002), .B(n15001), .Z(n15004) );
  XNOR U15572 ( .A(n15002), .B(n15001), .Z(n15385) );
  NAND U15573 ( .A(a[47]), .B(b[18]), .Z(n15384) );
  OR U15574 ( .A(n15385), .B(n15384), .Z(n15003) );
  NAND U15575 ( .A(n15004), .B(n15003), .Z(n15008) );
  NANDN U15576 ( .A(n15007), .B(n15008), .Z(n15010) );
  XOR U15577 ( .A(n15006), .B(n15005), .Z(n15390) );
  XNOR U15578 ( .A(n15008), .B(n15007), .Z(n15391) );
  NAND U15579 ( .A(n15390), .B(n15391), .Z(n15009) );
  NAND U15580 ( .A(n15010), .B(n15009), .Z(n15013) );
  AND U15581 ( .A(b[18]), .B(a[49]), .Z(n15014) );
  OR U15582 ( .A(n15013), .B(n15014), .Z(n15016) );
  XNOR U15583 ( .A(n15012), .B(n15011), .Z(n15397) );
  XOR U15584 ( .A(n15014), .B(n15013), .Z(n15396) );
  NANDN U15585 ( .A(n15397), .B(n15396), .Z(n15015) );
  NAND U15586 ( .A(n15016), .B(n15015), .Z(n15020) );
  NAND U15587 ( .A(a[50]), .B(b[18]), .Z(n15019) );
  OR U15588 ( .A(n15020), .B(n15019), .Z(n15022) );
  XOR U15589 ( .A(n15018), .B(n15017), .Z(n15402) );
  XOR U15590 ( .A(n15020), .B(n15019), .Z(n15403) );
  NAND U15591 ( .A(n15402), .B(n15403), .Z(n15021) );
  NAND U15592 ( .A(n15022), .B(n15021), .Z(n15025) );
  AND U15593 ( .A(b[18]), .B(a[51]), .Z(n15026) );
  OR U15594 ( .A(n15025), .B(n15026), .Z(n15028) );
  XNOR U15595 ( .A(n15024), .B(n15023), .Z(n15409) );
  XOR U15596 ( .A(n15026), .B(n15025), .Z(n15408) );
  NANDN U15597 ( .A(n15409), .B(n15408), .Z(n15027) );
  NAND U15598 ( .A(n15028), .B(n15027), .Z(n15032) );
  NAND U15599 ( .A(a[52]), .B(b[18]), .Z(n15031) );
  OR U15600 ( .A(n15032), .B(n15031), .Z(n15034) );
  XOR U15601 ( .A(n15030), .B(n15029), .Z(n15414) );
  XOR U15602 ( .A(n15032), .B(n15031), .Z(n15415) );
  NAND U15603 ( .A(n15414), .B(n15415), .Z(n15033) );
  NAND U15604 ( .A(n15034), .B(n15033), .Z(n15037) );
  AND U15605 ( .A(b[18]), .B(a[53]), .Z(n15038) );
  OR U15606 ( .A(n15037), .B(n15038), .Z(n15040) );
  XNOR U15607 ( .A(n15036), .B(n15035), .Z(n15421) );
  XOR U15608 ( .A(n15038), .B(n15037), .Z(n15420) );
  NANDN U15609 ( .A(n15421), .B(n15420), .Z(n15039) );
  NAND U15610 ( .A(n15040), .B(n15039), .Z(n15044) );
  NAND U15611 ( .A(a[54]), .B(b[18]), .Z(n15043) );
  OR U15612 ( .A(n15044), .B(n15043), .Z(n15046) );
  XOR U15613 ( .A(n15042), .B(n15041), .Z(n15426) );
  XOR U15614 ( .A(n15044), .B(n15043), .Z(n15427) );
  NAND U15615 ( .A(n15426), .B(n15427), .Z(n15045) );
  NAND U15616 ( .A(n15046), .B(n15045), .Z(n15049) );
  AND U15617 ( .A(b[18]), .B(a[55]), .Z(n15050) );
  OR U15618 ( .A(n15049), .B(n15050), .Z(n15052) );
  XNOR U15619 ( .A(n15048), .B(n15047), .Z(n15433) );
  XOR U15620 ( .A(n15050), .B(n15049), .Z(n15432) );
  NANDN U15621 ( .A(n15433), .B(n15432), .Z(n15051) );
  NAND U15622 ( .A(n15052), .B(n15051), .Z(n15056) );
  NAND U15623 ( .A(a[56]), .B(b[18]), .Z(n15055) );
  OR U15624 ( .A(n15056), .B(n15055), .Z(n15058) );
  XOR U15625 ( .A(n15054), .B(n15053), .Z(n15438) );
  XOR U15626 ( .A(n15056), .B(n15055), .Z(n15439) );
  NAND U15627 ( .A(n15438), .B(n15439), .Z(n15057) );
  NAND U15628 ( .A(n15058), .B(n15057), .Z(n15061) );
  AND U15629 ( .A(b[18]), .B(a[57]), .Z(n15062) );
  OR U15630 ( .A(n15061), .B(n15062), .Z(n15064) );
  XNOR U15631 ( .A(n15060), .B(n15059), .Z(n15445) );
  XOR U15632 ( .A(n15062), .B(n15061), .Z(n15444) );
  NANDN U15633 ( .A(n15445), .B(n15444), .Z(n15063) );
  NAND U15634 ( .A(n15064), .B(n15063), .Z(n15068) );
  NAND U15635 ( .A(a[58]), .B(b[18]), .Z(n15067) );
  OR U15636 ( .A(n15068), .B(n15067), .Z(n15070) );
  XOR U15637 ( .A(n15066), .B(n15065), .Z(n15450) );
  XOR U15638 ( .A(n15068), .B(n15067), .Z(n15451) );
  NAND U15639 ( .A(n15450), .B(n15451), .Z(n15069) );
  NAND U15640 ( .A(n15070), .B(n15069), .Z(n15073) );
  AND U15641 ( .A(b[18]), .B(a[59]), .Z(n15074) );
  OR U15642 ( .A(n15073), .B(n15074), .Z(n15076) );
  XNOR U15643 ( .A(n15072), .B(n15071), .Z(n15457) );
  XOR U15644 ( .A(n15074), .B(n15073), .Z(n15456) );
  NANDN U15645 ( .A(n15457), .B(n15456), .Z(n15075) );
  NAND U15646 ( .A(n15076), .B(n15075), .Z(n15080) );
  NAND U15647 ( .A(a[60]), .B(b[18]), .Z(n15079) );
  OR U15648 ( .A(n15080), .B(n15079), .Z(n15082) );
  XOR U15649 ( .A(n15078), .B(n15077), .Z(n15463) );
  XOR U15650 ( .A(n15080), .B(n15079), .Z(n15462) );
  NAND U15651 ( .A(n15463), .B(n15462), .Z(n15081) );
  NAND U15652 ( .A(n15082), .B(n15081), .Z(n15085) );
  AND U15653 ( .A(b[18]), .B(a[61]), .Z(n15086) );
  OR U15654 ( .A(n15085), .B(n15086), .Z(n15088) );
  XNOR U15655 ( .A(n15084), .B(n15083), .Z(n15469) );
  XOR U15656 ( .A(n15086), .B(n15085), .Z(n15468) );
  NANDN U15657 ( .A(n15469), .B(n15468), .Z(n15087) );
  NAND U15658 ( .A(n15088), .B(n15087), .Z(n15092) );
  NAND U15659 ( .A(a[62]), .B(b[18]), .Z(n15091) );
  OR U15660 ( .A(n15092), .B(n15091), .Z(n15094) );
  XOR U15661 ( .A(n15090), .B(n15089), .Z(n15474) );
  XOR U15662 ( .A(n15092), .B(n15091), .Z(n15475) );
  NAND U15663 ( .A(n15474), .B(n15475), .Z(n15093) );
  NAND U15664 ( .A(n15094), .B(n15093), .Z(n15097) );
  AND U15665 ( .A(b[18]), .B(a[63]), .Z(n15098) );
  OR U15666 ( .A(n15097), .B(n15098), .Z(n15100) );
  XOR U15667 ( .A(n15096), .B(n15095), .Z(n15104) );
  XOR U15668 ( .A(n15098), .B(n15097), .Z(n15103) );
  NANDN U15669 ( .A(n15104), .B(n15103), .Z(n15099) );
  NAND U15670 ( .A(n15100), .B(n15099), .Z(n15101) );
  XOR U15671 ( .A(n15102), .B(n15101), .Z(n24151) );
  XNOR U15672 ( .A(n15104), .B(n15103), .Z(n15479) );
  NAND U15673 ( .A(a[62]), .B(b[17]), .Z(n15470) );
  NAND U15674 ( .A(a[60]), .B(b[17]), .Z(n15458) );
  NAND U15675 ( .A(a[58]), .B(b[17]), .Z(n15446) );
  NAND U15676 ( .A(a[56]), .B(b[17]), .Z(n15434) );
  NAND U15677 ( .A(a[54]), .B(b[17]), .Z(n15422) );
  NAND U15678 ( .A(a[52]), .B(b[17]), .Z(n15410) );
  NAND U15679 ( .A(a[50]), .B(b[17]), .Z(n15398) );
  ANDN U15680 ( .B(b[17]), .A(n191), .Z(n15355) );
  ANDN U15681 ( .B(b[17]), .A(n189), .Z(n15343) );
  ANDN U15682 ( .B(b[17]), .A(n187), .Z(n15331) );
  ANDN U15683 ( .B(b[17]), .A(n21772), .Z(n15319) );
  ANDN U15684 ( .B(b[17]), .A(n184), .Z(n15307) );
  ANDN U15685 ( .B(b[17]), .A(n21751), .Z(n15295) );
  ANDN U15686 ( .B(b[17]), .A(n21740), .Z(n15283) );
  ANDN U15687 ( .B(b[17]), .A(n21727), .Z(n15271) );
  ANDN U15688 ( .B(b[17]), .A(n21716), .Z(n15259) );
  ANDN U15689 ( .B(b[17]), .A(n21703), .Z(n15247) );
  ANDN U15690 ( .B(b[17]), .A(n21692), .Z(n15235) );
  ANDN U15691 ( .B(b[17]), .A(n21681), .Z(n15223) );
  NAND U15692 ( .A(a[19]), .B(b[17]), .Z(n15211) );
  ANDN U15693 ( .B(b[17]), .A(n174), .Z(n15200) );
  XOR U15694 ( .A(n15108), .B(n15107), .Z(n15196) );
  ANDN U15695 ( .B(b[17]), .A(n172), .Z(n15193) );
  ANDN U15696 ( .B(b[17]), .A(n170), .Z(n15179) );
  ANDN U15697 ( .B(b[17]), .A(n21164), .Z(n15167) );
  ANDN U15698 ( .B(b[17]), .A(n21615), .Z(n15155) );
  ANDN U15699 ( .B(b[17]), .A(n166), .Z(n15143) );
  NAND U15700 ( .A(a[6]), .B(b[17]), .Z(n15138) );
  XOR U15701 ( .A(n15110), .B(n15109), .Z(n15139) );
  NANDN U15702 ( .A(n15138), .B(n15139), .Z(n15141) );
  ANDN U15703 ( .B(b[17]), .A(n164), .Z(n15133) );
  ANDN U15704 ( .B(b[17]), .A(n21580), .Z(n15120) );
  NAND U15705 ( .A(b[18]), .B(a[1]), .Z(n15113) );
  AND U15706 ( .A(b[17]), .B(a[0]), .Z(n15871) );
  NANDN U15707 ( .A(n15113), .B(n15871), .Z(n15112) );
  NAND U15708 ( .A(a[2]), .B(b[17]), .Z(n15111) );
  AND U15709 ( .A(n15112), .B(n15111), .Z(n15119) );
  NANDN U15710 ( .A(n15113), .B(a[0]), .Z(n15114) );
  XNOR U15711 ( .A(a[2]), .B(n15114), .Z(n15115) );
  NAND U15712 ( .A(b[17]), .B(n15115), .Z(n15502) );
  AND U15713 ( .A(a[1]), .B(b[18]), .Z(n15116) );
  XNOR U15714 ( .A(n15117), .B(n15116), .Z(n15501) );
  NANDN U15715 ( .A(n15502), .B(n15501), .Z(n15118) );
  NANDN U15716 ( .A(n15119), .B(n15118), .Z(n15121) );
  NANDN U15717 ( .A(n15120), .B(n15121), .Z(n15125) );
  XOR U15718 ( .A(n15121), .B(n15120), .Z(n15506) );
  NANDN U15719 ( .A(n15506), .B(n15505), .Z(n15124) );
  NAND U15720 ( .A(n15125), .B(n15124), .Z(n15129) );
  XOR U15721 ( .A(n15127), .B(n15126), .Z(n15128) );
  NANDN U15722 ( .A(n15129), .B(n15128), .Z(n15131) );
  NAND U15723 ( .A(a[4]), .B(b[17]), .Z(n15513) );
  NANDN U15724 ( .A(n15513), .B(n15514), .Z(n15130) );
  NAND U15725 ( .A(n15131), .B(n15130), .Z(n15132) );
  OR U15726 ( .A(n15133), .B(n15132), .Z(n15137) );
  XNOR U15727 ( .A(n15133), .B(n15132), .Z(n15488) );
  XOR U15728 ( .A(n15135), .B(n15134), .Z(n15489) );
  NANDN U15729 ( .A(n15488), .B(n15489), .Z(n15136) );
  NAND U15730 ( .A(n15137), .B(n15136), .Z(n15523) );
  XNOR U15731 ( .A(n15139), .B(n15138), .Z(n15524) );
  NANDN U15732 ( .A(n15523), .B(n15524), .Z(n15140) );
  NAND U15733 ( .A(n15141), .B(n15140), .Z(n15142) );
  OR U15734 ( .A(n15143), .B(n15142), .Z(n15147) );
  XNOR U15735 ( .A(n15143), .B(n15142), .Z(n15527) );
  XOR U15736 ( .A(n15145), .B(n15144), .Z(n15528) );
  NANDN U15737 ( .A(n15527), .B(n15528), .Z(n15146) );
  NAND U15738 ( .A(n15147), .B(n15146), .Z(n15150) );
  XOR U15739 ( .A(n15149), .B(n15148), .Z(n15151) );
  NANDN U15740 ( .A(n15150), .B(n15151), .Z(n15153) );
  NAND U15741 ( .A(a[8]), .B(b[17]), .Z(n15535) );
  XNOR U15742 ( .A(n15151), .B(n15150), .Z(n15536) );
  NANDN U15743 ( .A(n15535), .B(n15536), .Z(n15152) );
  NAND U15744 ( .A(n15153), .B(n15152), .Z(n15154) );
  OR U15745 ( .A(n15155), .B(n15154), .Z(n15159) );
  XNOR U15746 ( .A(n15155), .B(n15154), .Z(n15539) );
  XOR U15747 ( .A(n15157), .B(n15156), .Z(n15540) );
  NANDN U15748 ( .A(n15539), .B(n15540), .Z(n15158) );
  NAND U15749 ( .A(n15159), .B(n15158), .Z(n15163) );
  NAND U15750 ( .A(n15163), .B(n15162), .Z(n15165) );
  ANDN U15751 ( .B(b[17]), .A(n168), .Z(n15546) );
  XNOR U15752 ( .A(n15163), .B(n15162), .Z(n15545) );
  OR U15753 ( .A(n15546), .B(n15545), .Z(n15164) );
  NAND U15754 ( .A(n15165), .B(n15164), .Z(n15166) );
  NANDN U15755 ( .A(n15167), .B(n15166), .Z(n15171) );
  XOR U15756 ( .A(n15169), .B(n15168), .Z(n15551) );
  NANDN U15757 ( .A(n15552), .B(n15551), .Z(n15170) );
  NAND U15758 ( .A(n15171), .B(n15170), .Z(n15174) );
  XOR U15759 ( .A(n15173), .B(n15172), .Z(n15175) );
  NANDN U15760 ( .A(n15174), .B(n15175), .Z(n15177) );
  NAND U15761 ( .A(a[12]), .B(b[17]), .Z(n15559) );
  XNOR U15762 ( .A(n15175), .B(n15174), .Z(n15560) );
  NANDN U15763 ( .A(n15559), .B(n15560), .Z(n15176) );
  NAND U15764 ( .A(n15177), .B(n15176), .Z(n15178) );
  OR U15765 ( .A(n15179), .B(n15178), .Z(n15183) );
  XNOR U15766 ( .A(n15179), .B(n15178), .Z(n15563) );
  XOR U15767 ( .A(n15181), .B(n15180), .Z(n15564) );
  NANDN U15768 ( .A(n15563), .B(n15564), .Z(n15182) );
  NAND U15769 ( .A(n15183), .B(n15182), .Z(n15186) );
  XOR U15770 ( .A(n15185), .B(n15184), .Z(n15187) );
  NANDN U15771 ( .A(n15186), .B(n15187), .Z(n15189) );
  NAND U15772 ( .A(a[14]), .B(b[17]), .Z(n15571) );
  XNOR U15773 ( .A(n15187), .B(n15186), .Z(n15572) );
  NANDN U15774 ( .A(n15571), .B(n15572), .Z(n15188) );
  NAND U15775 ( .A(n15189), .B(n15188), .Z(n15192) );
  OR U15776 ( .A(n15193), .B(n15192), .Z(n15195) );
  XOR U15777 ( .A(n15191), .B(n15190), .Z(n15486) );
  XOR U15778 ( .A(n15193), .B(n15192), .Z(n15487) );
  NAND U15779 ( .A(n15486), .B(n15487), .Z(n15194) );
  NAND U15780 ( .A(n15195), .B(n15194), .Z(n15197) );
  NANDN U15781 ( .A(n15196), .B(n15197), .Z(n15199) );
  ANDN U15782 ( .B(b[17]), .A(n173), .Z(n15580) );
  XOR U15783 ( .A(n15197), .B(n15196), .Z(n15579) );
  OR U15784 ( .A(n15580), .B(n15579), .Z(n15198) );
  NAND U15785 ( .A(n15199), .B(n15198), .Z(n15201) );
  NANDN U15786 ( .A(n15200), .B(n15201), .Z(n15205) );
  XOR U15787 ( .A(n15201), .B(n15200), .Z(n15485) );
  XOR U15788 ( .A(n15203), .B(n15202), .Z(n15484) );
  NANDN U15789 ( .A(n15485), .B(n15484), .Z(n15204) );
  AND U15790 ( .A(n15205), .B(n15204), .Z(n15206) );
  OR U15791 ( .A(n15207), .B(n15206), .Z(n15209) );
  ANDN U15792 ( .B(b[17]), .A(n175), .Z(n15592) );
  XNOR U15793 ( .A(n15207), .B(n15206), .Z(n15591) );
  OR U15794 ( .A(n15592), .B(n15591), .Z(n15208) );
  AND U15795 ( .A(n15209), .B(n15208), .Z(n15210) );
  NANDN U15796 ( .A(n15211), .B(n15210), .Z(n15215) );
  XNOR U15797 ( .A(n15213), .B(n15212), .Z(n15483) );
  NAND U15798 ( .A(n15482), .B(n15483), .Z(n15214) );
  AND U15799 ( .A(n15215), .B(n15214), .Z(n15218) );
  XOR U15800 ( .A(n15217), .B(n15216), .Z(n15219) );
  NANDN U15801 ( .A(n15218), .B(n15219), .Z(n15221) );
  NAND U15802 ( .A(a[20]), .B(b[17]), .Z(n15601) );
  XNOR U15803 ( .A(n15219), .B(n15218), .Z(n15602) );
  NANDN U15804 ( .A(n15601), .B(n15602), .Z(n15220) );
  NAND U15805 ( .A(n15221), .B(n15220), .Z(n15222) );
  OR U15806 ( .A(n15223), .B(n15222), .Z(n15227) );
  XNOR U15807 ( .A(n15223), .B(n15222), .Z(n15605) );
  XOR U15808 ( .A(n15225), .B(n15224), .Z(n15606) );
  NANDN U15809 ( .A(n15605), .B(n15606), .Z(n15226) );
  NAND U15810 ( .A(n15227), .B(n15226), .Z(n15230) );
  XOR U15811 ( .A(n15229), .B(n15228), .Z(n15231) );
  NANDN U15812 ( .A(n15230), .B(n15231), .Z(n15233) );
  NAND U15813 ( .A(a[22]), .B(b[17]), .Z(n15613) );
  XNOR U15814 ( .A(n15231), .B(n15230), .Z(n15614) );
  NANDN U15815 ( .A(n15613), .B(n15614), .Z(n15232) );
  NAND U15816 ( .A(n15233), .B(n15232), .Z(n15234) );
  OR U15817 ( .A(n15235), .B(n15234), .Z(n15239) );
  XNOR U15818 ( .A(n15235), .B(n15234), .Z(n15617) );
  XOR U15819 ( .A(n15237), .B(n15236), .Z(n15618) );
  NANDN U15820 ( .A(n15617), .B(n15618), .Z(n15238) );
  NAND U15821 ( .A(n15239), .B(n15238), .Z(n15242) );
  XOR U15822 ( .A(n15241), .B(n15240), .Z(n15243) );
  NANDN U15823 ( .A(n15242), .B(n15243), .Z(n15245) );
  NAND U15824 ( .A(a[24]), .B(b[17]), .Z(n15625) );
  XNOR U15825 ( .A(n15243), .B(n15242), .Z(n15626) );
  NANDN U15826 ( .A(n15625), .B(n15626), .Z(n15244) );
  NAND U15827 ( .A(n15245), .B(n15244), .Z(n15246) );
  OR U15828 ( .A(n15247), .B(n15246), .Z(n15251) );
  XNOR U15829 ( .A(n15247), .B(n15246), .Z(n15629) );
  XOR U15830 ( .A(n15249), .B(n15248), .Z(n15630) );
  NANDN U15831 ( .A(n15629), .B(n15630), .Z(n15250) );
  NAND U15832 ( .A(n15251), .B(n15250), .Z(n15254) );
  XOR U15833 ( .A(n15253), .B(n15252), .Z(n15255) );
  NANDN U15834 ( .A(n15254), .B(n15255), .Z(n15257) );
  NAND U15835 ( .A(a[26]), .B(b[17]), .Z(n15637) );
  XNOR U15836 ( .A(n15255), .B(n15254), .Z(n15638) );
  NANDN U15837 ( .A(n15637), .B(n15638), .Z(n15256) );
  NAND U15838 ( .A(n15257), .B(n15256), .Z(n15258) );
  OR U15839 ( .A(n15259), .B(n15258), .Z(n15263) );
  XNOR U15840 ( .A(n15259), .B(n15258), .Z(n15641) );
  XOR U15841 ( .A(n15261), .B(n15260), .Z(n15642) );
  NANDN U15842 ( .A(n15641), .B(n15642), .Z(n15262) );
  NAND U15843 ( .A(n15263), .B(n15262), .Z(n15266) );
  XOR U15844 ( .A(n15265), .B(n15264), .Z(n15267) );
  NANDN U15845 ( .A(n15266), .B(n15267), .Z(n15269) );
  NAND U15846 ( .A(a[28]), .B(b[17]), .Z(n15649) );
  XNOR U15847 ( .A(n15267), .B(n15266), .Z(n15650) );
  NANDN U15848 ( .A(n15649), .B(n15650), .Z(n15268) );
  NAND U15849 ( .A(n15269), .B(n15268), .Z(n15270) );
  OR U15850 ( .A(n15271), .B(n15270), .Z(n15275) );
  XNOR U15851 ( .A(n15271), .B(n15270), .Z(n15653) );
  XOR U15852 ( .A(n15273), .B(n15272), .Z(n15654) );
  NANDN U15853 ( .A(n15653), .B(n15654), .Z(n15274) );
  NAND U15854 ( .A(n15275), .B(n15274), .Z(n15278) );
  XOR U15855 ( .A(n15277), .B(n15276), .Z(n15279) );
  NANDN U15856 ( .A(n15278), .B(n15279), .Z(n15281) );
  NAND U15857 ( .A(a[30]), .B(b[17]), .Z(n15661) );
  XNOR U15858 ( .A(n15279), .B(n15278), .Z(n15662) );
  NANDN U15859 ( .A(n15661), .B(n15662), .Z(n15280) );
  NAND U15860 ( .A(n15281), .B(n15280), .Z(n15282) );
  OR U15861 ( .A(n15283), .B(n15282), .Z(n15287) );
  XNOR U15862 ( .A(n15283), .B(n15282), .Z(n15665) );
  XOR U15863 ( .A(n15285), .B(n15284), .Z(n15666) );
  NANDN U15864 ( .A(n15665), .B(n15666), .Z(n15286) );
  NAND U15865 ( .A(n15287), .B(n15286), .Z(n15290) );
  XOR U15866 ( .A(n15289), .B(n15288), .Z(n15291) );
  NANDN U15867 ( .A(n15290), .B(n15291), .Z(n15293) );
  NAND U15868 ( .A(a[32]), .B(b[17]), .Z(n15673) );
  XNOR U15869 ( .A(n15291), .B(n15290), .Z(n15674) );
  NANDN U15870 ( .A(n15673), .B(n15674), .Z(n15292) );
  NAND U15871 ( .A(n15293), .B(n15292), .Z(n15294) );
  OR U15872 ( .A(n15295), .B(n15294), .Z(n15299) );
  XNOR U15873 ( .A(n15295), .B(n15294), .Z(n15677) );
  XOR U15874 ( .A(n15297), .B(n15296), .Z(n15678) );
  NANDN U15875 ( .A(n15677), .B(n15678), .Z(n15298) );
  NAND U15876 ( .A(n15299), .B(n15298), .Z(n15302) );
  XOR U15877 ( .A(n15301), .B(n15300), .Z(n15303) );
  NANDN U15878 ( .A(n15302), .B(n15303), .Z(n15305) );
  NAND U15879 ( .A(a[34]), .B(b[17]), .Z(n15685) );
  XNOR U15880 ( .A(n15303), .B(n15302), .Z(n15686) );
  NANDN U15881 ( .A(n15685), .B(n15686), .Z(n15304) );
  NAND U15882 ( .A(n15305), .B(n15304), .Z(n15306) );
  OR U15883 ( .A(n15307), .B(n15306), .Z(n15311) );
  XNOR U15884 ( .A(n15307), .B(n15306), .Z(n15689) );
  XOR U15885 ( .A(n15309), .B(n15308), .Z(n15690) );
  NANDN U15886 ( .A(n15689), .B(n15690), .Z(n15310) );
  NAND U15887 ( .A(n15311), .B(n15310), .Z(n15314) );
  XOR U15888 ( .A(n15313), .B(n15312), .Z(n15315) );
  NANDN U15889 ( .A(n15314), .B(n15315), .Z(n15317) );
  NAND U15890 ( .A(a[36]), .B(b[17]), .Z(n15697) );
  XNOR U15891 ( .A(n15315), .B(n15314), .Z(n15698) );
  NANDN U15892 ( .A(n15697), .B(n15698), .Z(n15316) );
  NAND U15893 ( .A(n15317), .B(n15316), .Z(n15318) );
  OR U15894 ( .A(n15319), .B(n15318), .Z(n15323) );
  XNOR U15895 ( .A(n15319), .B(n15318), .Z(n15701) );
  XOR U15896 ( .A(n15321), .B(n15320), .Z(n15702) );
  NANDN U15897 ( .A(n15701), .B(n15702), .Z(n15322) );
  NAND U15898 ( .A(n15323), .B(n15322), .Z(n15326) );
  XOR U15899 ( .A(n15325), .B(n15324), .Z(n15327) );
  NANDN U15900 ( .A(n15326), .B(n15327), .Z(n15329) );
  NAND U15901 ( .A(a[38]), .B(b[17]), .Z(n15709) );
  XNOR U15902 ( .A(n15327), .B(n15326), .Z(n15710) );
  NANDN U15903 ( .A(n15709), .B(n15710), .Z(n15328) );
  NAND U15904 ( .A(n15329), .B(n15328), .Z(n15330) );
  OR U15905 ( .A(n15331), .B(n15330), .Z(n15335) );
  XNOR U15906 ( .A(n15331), .B(n15330), .Z(n15713) );
  XOR U15907 ( .A(n15333), .B(n15332), .Z(n15714) );
  NANDN U15908 ( .A(n15713), .B(n15714), .Z(n15334) );
  NAND U15909 ( .A(n15335), .B(n15334), .Z(n15338) );
  XOR U15910 ( .A(n15337), .B(n15336), .Z(n15339) );
  NANDN U15911 ( .A(n15338), .B(n15339), .Z(n15341) );
  NAND U15912 ( .A(a[40]), .B(b[17]), .Z(n15721) );
  XNOR U15913 ( .A(n15339), .B(n15338), .Z(n15722) );
  NANDN U15914 ( .A(n15721), .B(n15722), .Z(n15340) );
  NAND U15915 ( .A(n15341), .B(n15340), .Z(n15342) );
  OR U15916 ( .A(n15343), .B(n15342), .Z(n15347) );
  XNOR U15917 ( .A(n15343), .B(n15342), .Z(n15725) );
  XOR U15918 ( .A(n15345), .B(n15344), .Z(n15726) );
  NANDN U15919 ( .A(n15725), .B(n15726), .Z(n15346) );
  NAND U15920 ( .A(n15347), .B(n15346), .Z(n15350) );
  XOR U15921 ( .A(n15349), .B(n15348), .Z(n15351) );
  NANDN U15922 ( .A(n15350), .B(n15351), .Z(n15353) );
  NAND U15923 ( .A(a[42]), .B(b[17]), .Z(n15733) );
  XNOR U15924 ( .A(n15351), .B(n15350), .Z(n15734) );
  NANDN U15925 ( .A(n15733), .B(n15734), .Z(n15352) );
  NAND U15926 ( .A(n15353), .B(n15352), .Z(n15354) );
  OR U15927 ( .A(n15355), .B(n15354), .Z(n15359) );
  XNOR U15928 ( .A(n15355), .B(n15354), .Z(n15737) );
  XOR U15929 ( .A(n15357), .B(n15356), .Z(n15738) );
  NANDN U15930 ( .A(n15737), .B(n15738), .Z(n15358) );
  NAND U15931 ( .A(n15359), .B(n15358), .Z(n15362) );
  XOR U15932 ( .A(n15361), .B(n15360), .Z(n15363) );
  NANDN U15933 ( .A(n15362), .B(n15363), .Z(n15365) );
  NAND U15934 ( .A(a[44]), .B(b[17]), .Z(n15745) );
  XNOR U15935 ( .A(n15363), .B(n15362), .Z(n15746) );
  NANDN U15936 ( .A(n15745), .B(n15746), .Z(n15364) );
  NAND U15937 ( .A(n15365), .B(n15364), .Z(n15368) );
  ANDN U15938 ( .B(b[17]), .A(n193), .Z(n15369) );
  OR U15939 ( .A(n15368), .B(n15369), .Z(n15371) );
  XOR U15940 ( .A(n15367), .B(n15366), .Z(n15750) );
  XOR U15941 ( .A(n15369), .B(n15368), .Z(n15749) );
  NANDN U15942 ( .A(n15750), .B(n15749), .Z(n15370) );
  NAND U15943 ( .A(n15371), .B(n15370), .Z(n15374) );
  XNOR U15944 ( .A(n15373), .B(n15372), .Z(n15375) );
  OR U15945 ( .A(n15374), .B(n15375), .Z(n15377) );
  XNOR U15946 ( .A(n15375), .B(n15374), .Z(n15756) );
  NAND U15947 ( .A(a[46]), .B(b[17]), .Z(n15755) );
  OR U15948 ( .A(n15756), .B(n15755), .Z(n15376) );
  NAND U15949 ( .A(n15377), .B(n15376), .Z(n15378) );
  ANDN U15950 ( .B(b[17]), .A(n195), .Z(n15379) );
  OR U15951 ( .A(n15378), .B(n15379), .Z(n15383) );
  XOR U15952 ( .A(n15379), .B(n15378), .Z(n15761) );
  NAND U15953 ( .A(n15761), .B(n15762), .Z(n15382) );
  NAND U15954 ( .A(n15383), .B(n15382), .Z(n15387) );
  NAND U15955 ( .A(a[48]), .B(b[17]), .Z(n15386) );
  OR U15956 ( .A(n15387), .B(n15386), .Z(n15389) );
  XOR U15957 ( .A(n15385), .B(n15384), .Z(n15767) );
  XOR U15958 ( .A(n15387), .B(n15386), .Z(n15768) );
  NAND U15959 ( .A(n15767), .B(n15768), .Z(n15388) );
  NAND U15960 ( .A(n15389), .B(n15388), .Z(n15393) );
  XOR U15961 ( .A(n15391), .B(n15390), .Z(n15392) );
  NAND U15962 ( .A(n15393), .B(n15392), .Z(n15395) );
  XNOR U15963 ( .A(n15393), .B(n15392), .Z(n15774) );
  NAND U15964 ( .A(a[49]), .B(b[17]), .Z(n15773) );
  OR U15965 ( .A(n15774), .B(n15773), .Z(n15394) );
  NAND U15966 ( .A(n15395), .B(n15394), .Z(n15399) );
  NANDN U15967 ( .A(n15398), .B(n15399), .Z(n15401) );
  XNOR U15968 ( .A(n15397), .B(n15396), .Z(n15780) );
  XNOR U15969 ( .A(n15399), .B(n15398), .Z(n15779) );
  NANDN U15970 ( .A(n15780), .B(n15779), .Z(n15400) );
  NAND U15971 ( .A(n15401), .B(n15400), .Z(n15405) );
  XOR U15972 ( .A(n15403), .B(n15402), .Z(n15404) );
  NAND U15973 ( .A(n15405), .B(n15404), .Z(n15407) );
  XNOR U15974 ( .A(n15405), .B(n15404), .Z(n15786) );
  NAND U15975 ( .A(a[51]), .B(b[17]), .Z(n15785) );
  OR U15976 ( .A(n15786), .B(n15785), .Z(n15406) );
  NAND U15977 ( .A(n15407), .B(n15406), .Z(n15411) );
  NANDN U15978 ( .A(n15410), .B(n15411), .Z(n15413) );
  XNOR U15979 ( .A(n15409), .B(n15408), .Z(n15792) );
  XNOR U15980 ( .A(n15411), .B(n15410), .Z(n15791) );
  NANDN U15981 ( .A(n15792), .B(n15791), .Z(n15412) );
  NAND U15982 ( .A(n15413), .B(n15412), .Z(n15417) );
  XOR U15983 ( .A(n15415), .B(n15414), .Z(n15416) );
  NAND U15984 ( .A(n15417), .B(n15416), .Z(n15419) );
  XNOR U15985 ( .A(n15417), .B(n15416), .Z(n15798) );
  NAND U15986 ( .A(a[53]), .B(b[17]), .Z(n15797) );
  OR U15987 ( .A(n15798), .B(n15797), .Z(n15418) );
  NAND U15988 ( .A(n15419), .B(n15418), .Z(n15423) );
  NANDN U15989 ( .A(n15422), .B(n15423), .Z(n15425) );
  XNOR U15990 ( .A(n15421), .B(n15420), .Z(n15804) );
  XNOR U15991 ( .A(n15423), .B(n15422), .Z(n15803) );
  NANDN U15992 ( .A(n15804), .B(n15803), .Z(n15424) );
  NAND U15993 ( .A(n15425), .B(n15424), .Z(n15429) );
  XOR U15994 ( .A(n15427), .B(n15426), .Z(n15428) );
  NAND U15995 ( .A(n15429), .B(n15428), .Z(n15431) );
  XNOR U15996 ( .A(n15429), .B(n15428), .Z(n15810) );
  NAND U15997 ( .A(a[55]), .B(b[17]), .Z(n15809) );
  OR U15998 ( .A(n15810), .B(n15809), .Z(n15430) );
  NAND U15999 ( .A(n15431), .B(n15430), .Z(n15435) );
  NANDN U16000 ( .A(n15434), .B(n15435), .Z(n15437) );
  XNOR U16001 ( .A(n15433), .B(n15432), .Z(n15816) );
  XNOR U16002 ( .A(n15435), .B(n15434), .Z(n15815) );
  NANDN U16003 ( .A(n15816), .B(n15815), .Z(n15436) );
  NAND U16004 ( .A(n15437), .B(n15436), .Z(n15441) );
  XOR U16005 ( .A(n15439), .B(n15438), .Z(n15440) );
  NAND U16006 ( .A(n15441), .B(n15440), .Z(n15443) );
  XNOR U16007 ( .A(n15441), .B(n15440), .Z(n15822) );
  NAND U16008 ( .A(a[57]), .B(b[17]), .Z(n15821) );
  OR U16009 ( .A(n15822), .B(n15821), .Z(n15442) );
  NAND U16010 ( .A(n15443), .B(n15442), .Z(n15447) );
  NANDN U16011 ( .A(n15446), .B(n15447), .Z(n15449) );
  XNOR U16012 ( .A(n15445), .B(n15444), .Z(n15828) );
  XNOR U16013 ( .A(n15447), .B(n15446), .Z(n15827) );
  NANDN U16014 ( .A(n15828), .B(n15827), .Z(n15448) );
  NAND U16015 ( .A(n15449), .B(n15448), .Z(n15453) );
  XOR U16016 ( .A(n15451), .B(n15450), .Z(n15452) );
  NAND U16017 ( .A(n15453), .B(n15452), .Z(n15455) );
  XNOR U16018 ( .A(n15453), .B(n15452), .Z(n15834) );
  NAND U16019 ( .A(a[59]), .B(b[17]), .Z(n15833) );
  OR U16020 ( .A(n15834), .B(n15833), .Z(n15454) );
  NAND U16021 ( .A(n15455), .B(n15454), .Z(n15459) );
  NANDN U16022 ( .A(n15458), .B(n15459), .Z(n15461) );
  XNOR U16023 ( .A(n15457), .B(n15456), .Z(n15840) );
  XNOR U16024 ( .A(n15459), .B(n15458), .Z(n15839) );
  NANDN U16025 ( .A(n15840), .B(n15839), .Z(n15460) );
  NAND U16026 ( .A(n15461), .B(n15460), .Z(n15465) );
  XOR U16027 ( .A(n15463), .B(n15462), .Z(n15464) );
  NAND U16028 ( .A(n15465), .B(n15464), .Z(n15467) );
  XNOR U16029 ( .A(n15465), .B(n15464), .Z(n15846) );
  NAND U16030 ( .A(a[61]), .B(b[17]), .Z(n15845) );
  OR U16031 ( .A(n15846), .B(n15845), .Z(n15466) );
  NAND U16032 ( .A(n15467), .B(n15466), .Z(n15471) );
  NANDN U16033 ( .A(n15470), .B(n15471), .Z(n15473) );
  XNOR U16034 ( .A(n15469), .B(n15468), .Z(n15852) );
  XNOR U16035 ( .A(n15471), .B(n15470), .Z(n15851) );
  NANDN U16036 ( .A(n15852), .B(n15851), .Z(n15472) );
  NAND U16037 ( .A(n15473), .B(n15472), .Z(n15476) );
  XOR U16038 ( .A(n15475), .B(n15474), .Z(n15477) );
  AND U16039 ( .A(b[17]), .B(a[63]), .Z(n15481) );
  XOR U16040 ( .A(n15477), .B(n15476), .Z(n15480) );
  NANDN U16041 ( .A(n15479), .B(n15478), .Z(n24150) );
  XNOR U16042 ( .A(n15479), .B(n15478), .Z(n21962) );
  XOR U16043 ( .A(n15481), .B(n15480), .Z(n15858) );
  NAND U16044 ( .A(a[50]), .B(b[16]), .Z(n15775) );
  ANDN U16045 ( .B(b[16]), .A(n193), .Z(n15744) );
  ANDN U16046 ( .B(b[16]), .A(n191), .Z(n15732) );
  ANDN U16047 ( .B(b[16]), .A(n189), .Z(n15720) );
  ANDN U16048 ( .B(b[16]), .A(n187), .Z(n15708) );
  ANDN U16049 ( .B(b[16]), .A(n21772), .Z(n15696) );
  ANDN U16050 ( .B(b[16]), .A(n184), .Z(n15684) );
  ANDN U16051 ( .B(b[16]), .A(n21751), .Z(n15672) );
  ANDN U16052 ( .B(b[16]), .A(n21740), .Z(n15660) );
  ANDN U16053 ( .B(b[16]), .A(n21727), .Z(n15648) );
  ANDN U16054 ( .B(b[16]), .A(n21716), .Z(n15636) );
  ANDN U16055 ( .B(b[16]), .A(n21703), .Z(n15624) );
  ANDN U16056 ( .B(b[16]), .A(n21692), .Z(n15612) );
  NAND U16057 ( .A(a[21]), .B(b[16]), .Z(n15600) );
  ANDN U16058 ( .B(b[16]), .A(n21670), .Z(n15589) );
  XOR U16059 ( .A(n15485), .B(n15484), .Z(n15585) );
  ANDN U16060 ( .B(b[16]), .A(n174), .Z(n15582) );
  ANDN U16061 ( .B(b[16]), .A(n172), .Z(n15570) );
  ANDN U16062 ( .B(b[16]), .A(n170), .Z(n15558) );
  ANDN U16063 ( .B(b[16]), .A(n21164), .Z(n15548) );
  ANDN U16064 ( .B(b[16]), .A(n21615), .Z(n15534) );
  ANDN U16065 ( .B(b[16]), .A(n166), .Z(n15522) );
  NAND U16066 ( .A(a[6]), .B(b[16]), .Z(n15517) );
  XOR U16067 ( .A(n15489), .B(n15488), .Z(n15518) );
  NANDN U16068 ( .A(n15517), .B(n15518), .Z(n15520) );
  ANDN U16069 ( .B(b[16]), .A(n164), .Z(n15512) );
  ANDN U16070 ( .B(b[16]), .A(n21580), .Z(n15499) );
  NAND U16071 ( .A(b[17]), .B(a[1]), .Z(n15492) );
  AND U16072 ( .A(b[16]), .B(a[0]), .Z(n16246) );
  NANDN U16073 ( .A(n15492), .B(n16246), .Z(n15491) );
  NAND U16074 ( .A(a[2]), .B(b[16]), .Z(n15490) );
  AND U16075 ( .A(n15491), .B(n15490), .Z(n15498) );
  NANDN U16076 ( .A(n15492), .B(a[0]), .Z(n15493) );
  XNOR U16077 ( .A(a[2]), .B(n15493), .Z(n15494) );
  NAND U16078 ( .A(b[16]), .B(n15494), .Z(n15877) );
  AND U16079 ( .A(a[1]), .B(b[17]), .Z(n15495) );
  XNOR U16080 ( .A(n15496), .B(n15495), .Z(n15876) );
  NANDN U16081 ( .A(n15877), .B(n15876), .Z(n15497) );
  NANDN U16082 ( .A(n15498), .B(n15497), .Z(n15500) );
  NANDN U16083 ( .A(n15499), .B(n15500), .Z(n15504) );
  XOR U16084 ( .A(n15500), .B(n15499), .Z(n15881) );
  NANDN U16085 ( .A(n15881), .B(n15880), .Z(n15503) );
  NAND U16086 ( .A(n15504), .B(n15503), .Z(n15508) );
  XOR U16087 ( .A(n15506), .B(n15505), .Z(n15507) );
  NANDN U16088 ( .A(n15508), .B(n15507), .Z(n15510) );
  NAND U16089 ( .A(a[4]), .B(b[16]), .Z(n15888) );
  NANDN U16090 ( .A(n15888), .B(n15889), .Z(n15509) );
  NAND U16091 ( .A(n15510), .B(n15509), .Z(n15511) );
  OR U16092 ( .A(n15512), .B(n15511), .Z(n15516) );
  XNOR U16093 ( .A(n15512), .B(n15511), .Z(n15892) );
  XOR U16094 ( .A(n15514), .B(n15513), .Z(n15893) );
  NANDN U16095 ( .A(n15892), .B(n15893), .Z(n15515) );
  NAND U16096 ( .A(n15516), .B(n15515), .Z(n15900) );
  XNOR U16097 ( .A(n15518), .B(n15517), .Z(n15901) );
  NANDN U16098 ( .A(n15900), .B(n15901), .Z(n15519) );
  NAND U16099 ( .A(n15520), .B(n15519), .Z(n15521) );
  OR U16100 ( .A(n15522), .B(n15521), .Z(n15526) );
  XNOR U16101 ( .A(n15522), .B(n15521), .Z(n15904) );
  XOR U16102 ( .A(n15524), .B(n15523), .Z(n15905) );
  NANDN U16103 ( .A(n15904), .B(n15905), .Z(n15525) );
  NAND U16104 ( .A(n15526), .B(n15525), .Z(n15529) );
  XOR U16105 ( .A(n15528), .B(n15527), .Z(n15530) );
  NANDN U16106 ( .A(n15529), .B(n15530), .Z(n15532) );
  NAND U16107 ( .A(a[8]), .B(b[16]), .Z(n15912) );
  XNOR U16108 ( .A(n15530), .B(n15529), .Z(n15913) );
  NANDN U16109 ( .A(n15912), .B(n15913), .Z(n15531) );
  NAND U16110 ( .A(n15532), .B(n15531), .Z(n15533) );
  OR U16111 ( .A(n15534), .B(n15533), .Z(n15538) );
  XNOR U16112 ( .A(n15534), .B(n15533), .Z(n15916) );
  XOR U16113 ( .A(n15536), .B(n15535), .Z(n15917) );
  NANDN U16114 ( .A(n15916), .B(n15917), .Z(n15537) );
  NAND U16115 ( .A(n15538), .B(n15537), .Z(n15541) );
  XOR U16116 ( .A(n15540), .B(n15539), .Z(n15542) );
  NANDN U16117 ( .A(n15541), .B(n15542), .Z(n15544) );
  NAND U16118 ( .A(a[10]), .B(b[16]), .Z(n15924) );
  XNOR U16119 ( .A(n15542), .B(n15541), .Z(n15925) );
  NANDN U16120 ( .A(n15924), .B(n15925), .Z(n15543) );
  NAND U16121 ( .A(n15544), .B(n15543), .Z(n15547) );
  OR U16122 ( .A(n15548), .B(n15547), .Z(n15550) );
  XOR U16123 ( .A(n15546), .B(n15545), .Z(n15928) );
  XOR U16124 ( .A(n15548), .B(n15547), .Z(n15929) );
  NAND U16125 ( .A(n15928), .B(n15929), .Z(n15549) );
  NAND U16126 ( .A(n15550), .B(n15549), .Z(n15553) );
  NANDN U16127 ( .A(n15553), .B(n15554), .Z(n15556) );
  NAND U16128 ( .A(a[12]), .B(b[16]), .Z(n15936) );
  XNOR U16129 ( .A(n15554), .B(n15553), .Z(n15937) );
  NANDN U16130 ( .A(n15936), .B(n15937), .Z(n15555) );
  NAND U16131 ( .A(n15556), .B(n15555), .Z(n15557) );
  OR U16132 ( .A(n15558), .B(n15557), .Z(n15562) );
  XNOR U16133 ( .A(n15558), .B(n15557), .Z(n15940) );
  XOR U16134 ( .A(n15560), .B(n15559), .Z(n15941) );
  NANDN U16135 ( .A(n15940), .B(n15941), .Z(n15561) );
  NAND U16136 ( .A(n15562), .B(n15561), .Z(n15565) );
  XOR U16137 ( .A(n15564), .B(n15563), .Z(n15566) );
  NANDN U16138 ( .A(n15565), .B(n15566), .Z(n15568) );
  NAND U16139 ( .A(a[14]), .B(b[16]), .Z(n15948) );
  XNOR U16140 ( .A(n15566), .B(n15565), .Z(n15949) );
  NANDN U16141 ( .A(n15948), .B(n15949), .Z(n15567) );
  NAND U16142 ( .A(n15568), .B(n15567), .Z(n15569) );
  OR U16143 ( .A(n15570), .B(n15569), .Z(n15574) );
  XNOR U16144 ( .A(n15570), .B(n15569), .Z(n15952) );
  XOR U16145 ( .A(n15572), .B(n15571), .Z(n15953) );
  NANDN U16146 ( .A(n15952), .B(n15953), .Z(n15573) );
  NAND U16147 ( .A(n15574), .B(n15573), .Z(n15575) );
  OR U16148 ( .A(n15576), .B(n15575), .Z(n15578) );
  NAND U16149 ( .A(a[16]), .B(b[16]), .Z(n15960) );
  XOR U16150 ( .A(n15576), .B(n15575), .Z(n15961) );
  NANDN U16151 ( .A(n15960), .B(n15961), .Z(n15577) );
  NAND U16152 ( .A(n15578), .B(n15577), .Z(n15581) );
  OR U16153 ( .A(n15582), .B(n15581), .Z(n15584) );
  XOR U16154 ( .A(n15580), .B(n15579), .Z(n15863) );
  XOR U16155 ( .A(n15582), .B(n15581), .Z(n15864) );
  NAND U16156 ( .A(n15863), .B(n15864), .Z(n15583) );
  NAND U16157 ( .A(n15584), .B(n15583), .Z(n15586) );
  NANDN U16158 ( .A(n15585), .B(n15586), .Z(n15588) );
  ANDN U16159 ( .B(b[16]), .A(n175), .Z(n15969) );
  XOR U16160 ( .A(n15586), .B(n15585), .Z(n15968) );
  OR U16161 ( .A(n15969), .B(n15968), .Z(n15587) );
  NAND U16162 ( .A(n15588), .B(n15587), .Z(n15590) );
  NANDN U16163 ( .A(n15589), .B(n15590), .Z(n15594) );
  XOR U16164 ( .A(n15590), .B(n15589), .Z(n15862) );
  XOR U16165 ( .A(n15592), .B(n15591), .Z(n15861) );
  NANDN U16166 ( .A(n15862), .B(n15861), .Z(n15593) );
  AND U16167 ( .A(n15594), .B(n15593), .Z(n15595) );
  OR U16168 ( .A(n15596), .B(n15595), .Z(n15598) );
  ANDN U16169 ( .B(b[16]), .A(n176), .Z(n15981) );
  XNOR U16170 ( .A(n15596), .B(n15595), .Z(n15980) );
  OR U16171 ( .A(n15981), .B(n15980), .Z(n15597) );
  AND U16172 ( .A(n15598), .B(n15597), .Z(n15599) );
  NANDN U16173 ( .A(n15600), .B(n15599), .Z(n15604) );
  XNOR U16174 ( .A(n15602), .B(n15601), .Z(n15860) );
  NAND U16175 ( .A(n15859), .B(n15860), .Z(n15603) );
  AND U16176 ( .A(n15604), .B(n15603), .Z(n15607) );
  XOR U16177 ( .A(n15606), .B(n15605), .Z(n15608) );
  NANDN U16178 ( .A(n15607), .B(n15608), .Z(n15610) );
  NAND U16179 ( .A(a[22]), .B(b[16]), .Z(n15990) );
  XNOR U16180 ( .A(n15608), .B(n15607), .Z(n15991) );
  NANDN U16181 ( .A(n15990), .B(n15991), .Z(n15609) );
  NAND U16182 ( .A(n15610), .B(n15609), .Z(n15611) );
  OR U16183 ( .A(n15612), .B(n15611), .Z(n15616) );
  XNOR U16184 ( .A(n15612), .B(n15611), .Z(n15994) );
  XOR U16185 ( .A(n15614), .B(n15613), .Z(n15995) );
  NANDN U16186 ( .A(n15994), .B(n15995), .Z(n15615) );
  NAND U16187 ( .A(n15616), .B(n15615), .Z(n15619) );
  XOR U16188 ( .A(n15618), .B(n15617), .Z(n15620) );
  NANDN U16189 ( .A(n15619), .B(n15620), .Z(n15622) );
  NAND U16190 ( .A(a[24]), .B(b[16]), .Z(n16002) );
  XNOR U16191 ( .A(n15620), .B(n15619), .Z(n16003) );
  NANDN U16192 ( .A(n16002), .B(n16003), .Z(n15621) );
  NAND U16193 ( .A(n15622), .B(n15621), .Z(n15623) );
  OR U16194 ( .A(n15624), .B(n15623), .Z(n15628) );
  XNOR U16195 ( .A(n15624), .B(n15623), .Z(n16006) );
  XOR U16196 ( .A(n15626), .B(n15625), .Z(n16007) );
  NANDN U16197 ( .A(n16006), .B(n16007), .Z(n15627) );
  NAND U16198 ( .A(n15628), .B(n15627), .Z(n15631) );
  XOR U16199 ( .A(n15630), .B(n15629), .Z(n15632) );
  NANDN U16200 ( .A(n15631), .B(n15632), .Z(n15634) );
  NAND U16201 ( .A(a[26]), .B(b[16]), .Z(n16014) );
  XNOR U16202 ( .A(n15632), .B(n15631), .Z(n16015) );
  NANDN U16203 ( .A(n16014), .B(n16015), .Z(n15633) );
  NAND U16204 ( .A(n15634), .B(n15633), .Z(n15635) );
  OR U16205 ( .A(n15636), .B(n15635), .Z(n15640) );
  XNOR U16206 ( .A(n15636), .B(n15635), .Z(n16018) );
  XOR U16207 ( .A(n15638), .B(n15637), .Z(n16019) );
  NANDN U16208 ( .A(n16018), .B(n16019), .Z(n15639) );
  NAND U16209 ( .A(n15640), .B(n15639), .Z(n15643) );
  XOR U16210 ( .A(n15642), .B(n15641), .Z(n15644) );
  NANDN U16211 ( .A(n15643), .B(n15644), .Z(n15646) );
  NAND U16212 ( .A(a[28]), .B(b[16]), .Z(n16026) );
  XNOR U16213 ( .A(n15644), .B(n15643), .Z(n16027) );
  NANDN U16214 ( .A(n16026), .B(n16027), .Z(n15645) );
  NAND U16215 ( .A(n15646), .B(n15645), .Z(n15647) );
  OR U16216 ( .A(n15648), .B(n15647), .Z(n15652) );
  XNOR U16217 ( .A(n15648), .B(n15647), .Z(n16030) );
  XOR U16218 ( .A(n15650), .B(n15649), .Z(n16031) );
  NANDN U16219 ( .A(n16030), .B(n16031), .Z(n15651) );
  NAND U16220 ( .A(n15652), .B(n15651), .Z(n15655) );
  XOR U16221 ( .A(n15654), .B(n15653), .Z(n15656) );
  NANDN U16222 ( .A(n15655), .B(n15656), .Z(n15658) );
  NAND U16223 ( .A(a[30]), .B(b[16]), .Z(n16038) );
  XNOR U16224 ( .A(n15656), .B(n15655), .Z(n16039) );
  NANDN U16225 ( .A(n16038), .B(n16039), .Z(n15657) );
  NAND U16226 ( .A(n15658), .B(n15657), .Z(n15659) );
  OR U16227 ( .A(n15660), .B(n15659), .Z(n15664) );
  XNOR U16228 ( .A(n15660), .B(n15659), .Z(n16042) );
  XOR U16229 ( .A(n15662), .B(n15661), .Z(n16043) );
  NANDN U16230 ( .A(n16042), .B(n16043), .Z(n15663) );
  NAND U16231 ( .A(n15664), .B(n15663), .Z(n15667) );
  XOR U16232 ( .A(n15666), .B(n15665), .Z(n15668) );
  NANDN U16233 ( .A(n15667), .B(n15668), .Z(n15670) );
  NAND U16234 ( .A(a[32]), .B(b[16]), .Z(n16050) );
  XNOR U16235 ( .A(n15668), .B(n15667), .Z(n16051) );
  NANDN U16236 ( .A(n16050), .B(n16051), .Z(n15669) );
  NAND U16237 ( .A(n15670), .B(n15669), .Z(n15671) );
  OR U16238 ( .A(n15672), .B(n15671), .Z(n15676) );
  XNOR U16239 ( .A(n15672), .B(n15671), .Z(n16054) );
  XOR U16240 ( .A(n15674), .B(n15673), .Z(n16055) );
  NANDN U16241 ( .A(n16054), .B(n16055), .Z(n15675) );
  NAND U16242 ( .A(n15676), .B(n15675), .Z(n15679) );
  XOR U16243 ( .A(n15678), .B(n15677), .Z(n15680) );
  NANDN U16244 ( .A(n15679), .B(n15680), .Z(n15682) );
  NAND U16245 ( .A(a[34]), .B(b[16]), .Z(n16062) );
  XNOR U16246 ( .A(n15680), .B(n15679), .Z(n16063) );
  NANDN U16247 ( .A(n16062), .B(n16063), .Z(n15681) );
  NAND U16248 ( .A(n15682), .B(n15681), .Z(n15683) );
  OR U16249 ( .A(n15684), .B(n15683), .Z(n15688) );
  XNOR U16250 ( .A(n15684), .B(n15683), .Z(n16066) );
  XOR U16251 ( .A(n15686), .B(n15685), .Z(n16067) );
  NANDN U16252 ( .A(n16066), .B(n16067), .Z(n15687) );
  NAND U16253 ( .A(n15688), .B(n15687), .Z(n15691) );
  XOR U16254 ( .A(n15690), .B(n15689), .Z(n15692) );
  NANDN U16255 ( .A(n15691), .B(n15692), .Z(n15694) );
  NAND U16256 ( .A(a[36]), .B(b[16]), .Z(n16074) );
  XNOR U16257 ( .A(n15692), .B(n15691), .Z(n16075) );
  NANDN U16258 ( .A(n16074), .B(n16075), .Z(n15693) );
  NAND U16259 ( .A(n15694), .B(n15693), .Z(n15695) );
  OR U16260 ( .A(n15696), .B(n15695), .Z(n15700) );
  XNOR U16261 ( .A(n15696), .B(n15695), .Z(n16078) );
  XOR U16262 ( .A(n15698), .B(n15697), .Z(n16079) );
  NANDN U16263 ( .A(n16078), .B(n16079), .Z(n15699) );
  NAND U16264 ( .A(n15700), .B(n15699), .Z(n15703) );
  XOR U16265 ( .A(n15702), .B(n15701), .Z(n15704) );
  NANDN U16266 ( .A(n15703), .B(n15704), .Z(n15706) );
  NAND U16267 ( .A(a[38]), .B(b[16]), .Z(n16086) );
  XNOR U16268 ( .A(n15704), .B(n15703), .Z(n16087) );
  NANDN U16269 ( .A(n16086), .B(n16087), .Z(n15705) );
  NAND U16270 ( .A(n15706), .B(n15705), .Z(n15707) );
  OR U16271 ( .A(n15708), .B(n15707), .Z(n15712) );
  XNOR U16272 ( .A(n15708), .B(n15707), .Z(n16090) );
  XOR U16273 ( .A(n15710), .B(n15709), .Z(n16091) );
  NANDN U16274 ( .A(n16090), .B(n16091), .Z(n15711) );
  NAND U16275 ( .A(n15712), .B(n15711), .Z(n15715) );
  XOR U16276 ( .A(n15714), .B(n15713), .Z(n15716) );
  NANDN U16277 ( .A(n15715), .B(n15716), .Z(n15718) );
  NAND U16278 ( .A(a[40]), .B(b[16]), .Z(n16098) );
  XNOR U16279 ( .A(n15716), .B(n15715), .Z(n16099) );
  NANDN U16280 ( .A(n16098), .B(n16099), .Z(n15717) );
  NAND U16281 ( .A(n15718), .B(n15717), .Z(n15719) );
  OR U16282 ( .A(n15720), .B(n15719), .Z(n15724) );
  XNOR U16283 ( .A(n15720), .B(n15719), .Z(n16102) );
  XOR U16284 ( .A(n15722), .B(n15721), .Z(n16103) );
  NANDN U16285 ( .A(n16102), .B(n16103), .Z(n15723) );
  NAND U16286 ( .A(n15724), .B(n15723), .Z(n15727) );
  XOR U16287 ( .A(n15726), .B(n15725), .Z(n15728) );
  NANDN U16288 ( .A(n15727), .B(n15728), .Z(n15730) );
  NAND U16289 ( .A(a[42]), .B(b[16]), .Z(n16110) );
  XNOR U16290 ( .A(n15728), .B(n15727), .Z(n16111) );
  NANDN U16291 ( .A(n16110), .B(n16111), .Z(n15729) );
  NAND U16292 ( .A(n15730), .B(n15729), .Z(n15731) );
  OR U16293 ( .A(n15732), .B(n15731), .Z(n15736) );
  XNOR U16294 ( .A(n15732), .B(n15731), .Z(n16114) );
  XOR U16295 ( .A(n15734), .B(n15733), .Z(n16115) );
  NANDN U16296 ( .A(n16114), .B(n16115), .Z(n15735) );
  NAND U16297 ( .A(n15736), .B(n15735), .Z(n15739) );
  XOR U16298 ( .A(n15738), .B(n15737), .Z(n15740) );
  NANDN U16299 ( .A(n15739), .B(n15740), .Z(n15742) );
  NAND U16300 ( .A(a[44]), .B(b[16]), .Z(n16122) );
  XNOR U16301 ( .A(n15740), .B(n15739), .Z(n16123) );
  NANDN U16302 ( .A(n16122), .B(n16123), .Z(n15741) );
  NAND U16303 ( .A(n15742), .B(n15741), .Z(n15743) );
  OR U16304 ( .A(n15744), .B(n15743), .Z(n15748) );
  XNOR U16305 ( .A(n15744), .B(n15743), .Z(n16126) );
  XOR U16306 ( .A(n15746), .B(n15745), .Z(n16127) );
  NANDN U16307 ( .A(n16126), .B(n16127), .Z(n15747) );
  NAND U16308 ( .A(n15748), .B(n15747), .Z(n15751) );
  XNOR U16309 ( .A(n15750), .B(n15749), .Z(n15752) );
  OR U16310 ( .A(n15751), .B(n15752), .Z(n15754) );
  XNOR U16311 ( .A(n15752), .B(n15751), .Z(n16133) );
  NAND U16312 ( .A(a[46]), .B(b[16]), .Z(n16132) );
  OR U16313 ( .A(n16133), .B(n16132), .Z(n15753) );
  NAND U16314 ( .A(n15754), .B(n15753), .Z(n15757) );
  ANDN U16315 ( .B(b[16]), .A(n195), .Z(n15758) );
  OR U16316 ( .A(n15757), .B(n15758), .Z(n15760) );
  XOR U16317 ( .A(n15756), .B(n15755), .Z(n16139) );
  XOR U16318 ( .A(n15758), .B(n15757), .Z(n16138) );
  NANDN U16319 ( .A(n16139), .B(n16138), .Z(n15759) );
  NAND U16320 ( .A(n15760), .B(n15759), .Z(n15764) );
  AND U16321 ( .A(b[16]), .B(a[48]), .Z(n15763) );
  NANDN U16322 ( .A(n15764), .B(n15763), .Z(n15766) );
  XNOR U16323 ( .A(n15764), .B(n15763), .Z(n16146) );
  NANDN U16324 ( .A(n16147), .B(n16146), .Z(n15765) );
  NAND U16325 ( .A(n15766), .B(n15765), .Z(n15770) );
  XOR U16326 ( .A(n15768), .B(n15767), .Z(n15769) );
  NAND U16327 ( .A(n15770), .B(n15769), .Z(n15772) );
  XNOR U16328 ( .A(n15770), .B(n15769), .Z(n16151) );
  NAND U16329 ( .A(a[49]), .B(b[16]), .Z(n16150) );
  OR U16330 ( .A(n16151), .B(n16150), .Z(n15771) );
  NAND U16331 ( .A(n15772), .B(n15771), .Z(n15776) );
  NANDN U16332 ( .A(n15775), .B(n15776), .Z(n15778) );
  XOR U16333 ( .A(n15774), .B(n15773), .Z(n16156) );
  XNOR U16334 ( .A(n15776), .B(n15775), .Z(n16157) );
  NAND U16335 ( .A(n16156), .B(n16157), .Z(n15777) );
  NAND U16336 ( .A(n15778), .B(n15777), .Z(n15781) );
  AND U16337 ( .A(b[16]), .B(a[51]), .Z(n15782) );
  OR U16338 ( .A(n15781), .B(n15782), .Z(n15784) );
  XNOR U16339 ( .A(n15780), .B(n15779), .Z(n16163) );
  XOR U16340 ( .A(n15782), .B(n15781), .Z(n16162) );
  NANDN U16341 ( .A(n16163), .B(n16162), .Z(n15783) );
  NAND U16342 ( .A(n15784), .B(n15783), .Z(n15788) );
  NAND U16343 ( .A(a[52]), .B(b[16]), .Z(n15787) );
  OR U16344 ( .A(n15788), .B(n15787), .Z(n15790) );
  XOR U16345 ( .A(n15786), .B(n15785), .Z(n16168) );
  XOR U16346 ( .A(n15788), .B(n15787), .Z(n16169) );
  NAND U16347 ( .A(n16168), .B(n16169), .Z(n15789) );
  NAND U16348 ( .A(n15790), .B(n15789), .Z(n15793) );
  AND U16349 ( .A(b[16]), .B(a[53]), .Z(n15794) );
  OR U16350 ( .A(n15793), .B(n15794), .Z(n15796) );
  XNOR U16351 ( .A(n15792), .B(n15791), .Z(n16175) );
  XOR U16352 ( .A(n15794), .B(n15793), .Z(n16174) );
  NANDN U16353 ( .A(n16175), .B(n16174), .Z(n15795) );
  NAND U16354 ( .A(n15796), .B(n15795), .Z(n15800) );
  NAND U16355 ( .A(a[54]), .B(b[16]), .Z(n15799) );
  OR U16356 ( .A(n15800), .B(n15799), .Z(n15802) );
  XOR U16357 ( .A(n15798), .B(n15797), .Z(n16180) );
  XOR U16358 ( .A(n15800), .B(n15799), .Z(n16181) );
  NAND U16359 ( .A(n16180), .B(n16181), .Z(n15801) );
  NAND U16360 ( .A(n15802), .B(n15801), .Z(n15805) );
  AND U16361 ( .A(b[16]), .B(a[55]), .Z(n15806) );
  OR U16362 ( .A(n15805), .B(n15806), .Z(n15808) );
  XNOR U16363 ( .A(n15804), .B(n15803), .Z(n16187) );
  XOR U16364 ( .A(n15806), .B(n15805), .Z(n16186) );
  NANDN U16365 ( .A(n16187), .B(n16186), .Z(n15807) );
  NAND U16366 ( .A(n15808), .B(n15807), .Z(n15812) );
  NAND U16367 ( .A(a[56]), .B(b[16]), .Z(n15811) );
  OR U16368 ( .A(n15812), .B(n15811), .Z(n15814) );
  XOR U16369 ( .A(n15810), .B(n15809), .Z(n16192) );
  XOR U16370 ( .A(n15812), .B(n15811), .Z(n16193) );
  NAND U16371 ( .A(n16192), .B(n16193), .Z(n15813) );
  NAND U16372 ( .A(n15814), .B(n15813), .Z(n15817) );
  AND U16373 ( .A(b[16]), .B(a[57]), .Z(n15818) );
  OR U16374 ( .A(n15817), .B(n15818), .Z(n15820) );
  XNOR U16375 ( .A(n15816), .B(n15815), .Z(n16199) );
  XOR U16376 ( .A(n15818), .B(n15817), .Z(n16198) );
  NANDN U16377 ( .A(n16199), .B(n16198), .Z(n15819) );
  NAND U16378 ( .A(n15820), .B(n15819), .Z(n15824) );
  NAND U16379 ( .A(a[58]), .B(b[16]), .Z(n15823) );
  OR U16380 ( .A(n15824), .B(n15823), .Z(n15826) );
  XOR U16381 ( .A(n15822), .B(n15821), .Z(n16204) );
  XOR U16382 ( .A(n15824), .B(n15823), .Z(n16205) );
  NAND U16383 ( .A(n16204), .B(n16205), .Z(n15825) );
  NAND U16384 ( .A(n15826), .B(n15825), .Z(n15829) );
  AND U16385 ( .A(b[16]), .B(a[59]), .Z(n15830) );
  OR U16386 ( .A(n15829), .B(n15830), .Z(n15832) );
  XNOR U16387 ( .A(n15828), .B(n15827), .Z(n16211) );
  XOR U16388 ( .A(n15830), .B(n15829), .Z(n16210) );
  NANDN U16389 ( .A(n16211), .B(n16210), .Z(n15831) );
  NAND U16390 ( .A(n15832), .B(n15831), .Z(n15836) );
  NAND U16391 ( .A(a[60]), .B(b[16]), .Z(n15835) );
  OR U16392 ( .A(n15836), .B(n15835), .Z(n15838) );
  XOR U16393 ( .A(n15834), .B(n15833), .Z(n16216) );
  XOR U16394 ( .A(n15836), .B(n15835), .Z(n16217) );
  NAND U16395 ( .A(n16216), .B(n16217), .Z(n15837) );
  NAND U16396 ( .A(n15838), .B(n15837), .Z(n15841) );
  AND U16397 ( .A(b[16]), .B(a[61]), .Z(n15842) );
  OR U16398 ( .A(n15841), .B(n15842), .Z(n15844) );
  XNOR U16399 ( .A(n15840), .B(n15839), .Z(n16223) );
  XOR U16400 ( .A(n15842), .B(n15841), .Z(n16222) );
  NANDN U16401 ( .A(n16223), .B(n16222), .Z(n15843) );
  NAND U16402 ( .A(n15844), .B(n15843), .Z(n15848) );
  NAND U16403 ( .A(a[62]), .B(b[16]), .Z(n15847) );
  OR U16404 ( .A(n15848), .B(n15847), .Z(n15850) );
  XOR U16405 ( .A(n15846), .B(n15845), .Z(n16228) );
  XOR U16406 ( .A(n15848), .B(n15847), .Z(n16229) );
  NAND U16407 ( .A(n16228), .B(n16229), .Z(n15849) );
  NAND U16408 ( .A(n15850), .B(n15849), .Z(n15853) );
  AND U16409 ( .A(b[16]), .B(a[63]), .Z(n15854) );
  OR U16410 ( .A(n15853), .B(n15854), .Z(n15856) );
  XNOR U16411 ( .A(n15852), .B(n15851), .Z(n16233) );
  XOR U16412 ( .A(n15854), .B(n15853), .Z(n16232) );
  NANDN U16413 ( .A(n16233), .B(n16232), .Z(n15855) );
  NAND U16414 ( .A(n15856), .B(n15855), .Z(n15857) );
  OR U16415 ( .A(n21962), .B(n21963), .Z(n21965) );
  XOR U16416 ( .A(n15858), .B(n15857), .Z(n21961) );
  NAND U16417 ( .A(a[62]), .B(b[15]), .Z(n16224) );
  NAND U16418 ( .A(a[60]), .B(b[15]), .Z(n16212) );
  NAND U16419 ( .A(a[58]), .B(b[15]), .Z(n16200) );
  NAND U16420 ( .A(a[56]), .B(b[15]), .Z(n16188) );
  NAND U16421 ( .A(a[54]), .B(b[15]), .Z(n16176) );
  NAND U16422 ( .A(a[52]), .B(b[15]), .Z(n16164) );
  ANDN U16423 ( .B(b[15]), .A(n193), .Z(n16121) );
  ANDN U16424 ( .B(b[15]), .A(n191), .Z(n16109) );
  ANDN U16425 ( .B(b[15]), .A(n189), .Z(n16097) );
  ANDN U16426 ( .B(b[15]), .A(n187), .Z(n16085) );
  ANDN U16427 ( .B(b[15]), .A(n21772), .Z(n16073) );
  ANDN U16428 ( .B(b[15]), .A(n184), .Z(n16061) );
  ANDN U16429 ( .B(b[15]), .A(n21751), .Z(n16049) );
  ANDN U16430 ( .B(b[15]), .A(n21740), .Z(n16037) );
  ANDN U16431 ( .B(b[15]), .A(n21727), .Z(n16025) );
  ANDN U16432 ( .B(b[15]), .A(n21716), .Z(n16013) );
  ANDN U16433 ( .B(b[15]), .A(n21703), .Z(n16001) );
  ANDN U16434 ( .B(b[15]), .A(n21692), .Z(n15989) );
  ANDN U16435 ( .B(b[15]), .A(n21681), .Z(n15978) );
  XOR U16436 ( .A(n15862), .B(n15861), .Z(n15974) );
  ANDN U16437 ( .B(b[15]), .A(n21670), .Z(n15971) );
  ANDN U16438 ( .B(b[15]), .A(n174), .Z(n15959) );
  ANDN U16439 ( .B(b[15]), .A(n172), .Z(n15947) );
  NAND U16440 ( .A(a[13]), .B(b[15]), .Z(n15935) );
  ANDN U16441 ( .B(b[15]), .A(n21164), .Z(n15923) );
  ANDN U16442 ( .B(b[15]), .A(n21615), .Z(n15911) );
  ANDN U16443 ( .B(b[15]), .A(n166), .Z(n15899) );
  ANDN U16444 ( .B(b[15]), .A(n164), .Z(n15887) );
  ANDN U16445 ( .B(b[15]), .A(n21580), .Z(n15874) );
  NAND U16446 ( .A(b[16]), .B(a[1]), .Z(n15867) );
  AND U16447 ( .A(b[15]), .B(a[0]), .Z(n16639) );
  NANDN U16448 ( .A(n15867), .B(n16639), .Z(n15866) );
  NAND U16449 ( .A(a[2]), .B(b[15]), .Z(n15865) );
  AND U16450 ( .A(n15866), .B(n15865), .Z(n15873) );
  NANDN U16451 ( .A(n15867), .B(a[0]), .Z(n15868) );
  XNOR U16452 ( .A(a[2]), .B(n15868), .Z(n15869) );
  NAND U16453 ( .A(b[15]), .B(n15869), .Z(n16252) );
  AND U16454 ( .A(a[1]), .B(b[16]), .Z(n15870) );
  XNOR U16455 ( .A(n15871), .B(n15870), .Z(n16251) );
  NANDN U16456 ( .A(n16252), .B(n16251), .Z(n15872) );
  NANDN U16457 ( .A(n15873), .B(n15872), .Z(n15875) );
  NANDN U16458 ( .A(n15874), .B(n15875), .Z(n15879) );
  XOR U16459 ( .A(n15875), .B(n15874), .Z(n16256) );
  NANDN U16460 ( .A(n16256), .B(n16255), .Z(n15878) );
  NAND U16461 ( .A(n15879), .B(n15878), .Z(n15883) );
  XOR U16462 ( .A(n15881), .B(n15880), .Z(n15882) );
  NANDN U16463 ( .A(n15883), .B(n15882), .Z(n15885) );
  NAND U16464 ( .A(a[4]), .B(b[15]), .Z(n16263) );
  NANDN U16465 ( .A(n16263), .B(n16264), .Z(n15884) );
  NAND U16466 ( .A(n15885), .B(n15884), .Z(n15886) );
  OR U16467 ( .A(n15887), .B(n15886), .Z(n15891) );
  XNOR U16468 ( .A(n15887), .B(n15886), .Z(n16267) );
  XOR U16469 ( .A(n15889), .B(n15888), .Z(n16268) );
  NANDN U16470 ( .A(n16267), .B(n16268), .Z(n15890) );
  NAND U16471 ( .A(n15891), .B(n15890), .Z(n15894) );
  XOR U16472 ( .A(n15893), .B(n15892), .Z(n15895) );
  NANDN U16473 ( .A(n15894), .B(n15895), .Z(n15897) );
  NAND U16474 ( .A(a[6]), .B(b[15]), .Z(n16275) );
  XNOR U16475 ( .A(n15895), .B(n15894), .Z(n16276) );
  NANDN U16476 ( .A(n16275), .B(n16276), .Z(n15896) );
  NAND U16477 ( .A(n15897), .B(n15896), .Z(n15898) );
  OR U16478 ( .A(n15899), .B(n15898), .Z(n15903) );
  XNOR U16479 ( .A(n15899), .B(n15898), .Z(n16279) );
  XOR U16480 ( .A(n15901), .B(n15900), .Z(n16280) );
  NANDN U16481 ( .A(n16279), .B(n16280), .Z(n15902) );
  NAND U16482 ( .A(n15903), .B(n15902), .Z(n15906) );
  XOR U16483 ( .A(n15905), .B(n15904), .Z(n15907) );
  NANDN U16484 ( .A(n15906), .B(n15907), .Z(n15909) );
  NAND U16485 ( .A(a[8]), .B(b[15]), .Z(n16285) );
  XNOR U16486 ( .A(n15907), .B(n15906), .Z(n16286) );
  NANDN U16487 ( .A(n16285), .B(n16286), .Z(n15908) );
  NAND U16488 ( .A(n15909), .B(n15908), .Z(n15910) );
  OR U16489 ( .A(n15911), .B(n15910), .Z(n15915) );
  XNOR U16490 ( .A(n15911), .B(n15910), .Z(n16291) );
  XOR U16491 ( .A(n15913), .B(n15912), .Z(n16292) );
  NANDN U16492 ( .A(n16291), .B(n16292), .Z(n15914) );
  NAND U16493 ( .A(n15915), .B(n15914), .Z(n15918) );
  XOR U16494 ( .A(n15917), .B(n15916), .Z(n15919) );
  NANDN U16495 ( .A(n15918), .B(n15919), .Z(n15921) );
  NAND U16496 ( .A(a[10]), .B(b[15]), .Z(n16299) );
  XNOR U16497 ( .A(n15919), .B(n15918), .Z(n16300) );
  NANDN U16498 ( .A(n16299), .B(n16300), .Z(n15920) );
  NAND U16499 ( .A(n15921), .B(n15920), .Z(n15922) );
  OR U16500 ( .A(n15923), .B(n15922), .Z(n15927) );
  XNOR U16501 ( .A(n15923), .B(n15922), .Z(n16303) );
  XOR U16502 ( .A(n15925), .B(n15924), .Z(n16304) );
  NANDN U16503 ( .A(n16303), .B(n16304), .Z(n15926) );
  NAND U16504 ( .A(n15927), .B(n15926), .Z(n15931) );
  NAND U16505 ( .A(n15931), .B(n15930), .Z(n15933) );
  ANDN U16506 ( .B(b[15]), .A(n169), .Z(n16312) );
  XNOR U16507 ( .A(n15931), .B(n15930), .Z(n16311) );
  OR U16508 ( .A(n16312), .B(n16311), .Z(n15932) );
  AND U16509 ( .A(n15933), .B(n15932), .Z(n15934) );
  NANDN U16510 ( .A(n15935), .B(n15934), .Z(n15939) );
  XNOR U16511 ( .A(n15937), .B(n15936), .Z(n16239) );
  NAND U16512 ( .A(n16238), .B(n16239), .Z(n15938) );
  AND U16513 ( .A(n15939), .B(n15938), .Z(n15942) );
  XOR U16514 ( .A(n15941), .B(n15940), .Z(n15943) );
  NANDN U16515 ( .A(n15942), .B(n15943), .Z(n15945) );
  NAND U16516 ( .A(a[14]), .B(b[15]), .Z(n16321) );
  XNOR U16517 ( .A(n15943), .B(n15942), .Z(n16322) );
  NANDN U16518 ( .A(n16321), .B(n16322), .Z(n15944) );
  NAND U16519 ( .A(n15945), .B(n15944), .Z(n15946) );
  OR U16520 ( .A(n15947), .B(n15946), .Z(n15951) );
  XNOR U16521 ( .A(n15947), .B(n15946), .Z(n16325) );
  XOR U16522 ( .A(n15949), .B(n15948), .Z(n16326) );
  NANDN U16523 ( .A(n16325), .B(n16326), .Z(n15950) );
  NAND U16524 ( .A(n15951), .B(n15950), .Z(n15954) );
  XOR U16525 ( .A(n15953), .B(n15952), .Z(n15955) );
  NANDN U16526 ( .A(n15954), .B(n15955), .Z(n15957) );
  NAND U16527 ( .A(a[16]), .B(b[15]), .Z(n16331) );
  XNOR U16528 ( .A(n15955), .B(n15954), .Z(n16332) );
  NANDN U16529 ( .A(n16331), .B(n16332), .Z(n15956) );
  NAND U16530 ( .A(n15957), .B(n15956), .Z(n15958) );
  OR U16531 ( .A(n15959), .B(n15958), .Z(n15963) );
  XNOR U16532 ( .A(n15959), .B(n15958), .Z(n16337) );
  XOR U16533 ( .A(n15961), .B(n15960), .Z(n16338) );
  NANDN U16534 ( .A(n16337), .B(n16338), .Z(n15962) );
  NAND U16535 ( .A(n15963), .B(n15962), .Z(n15964) );
  OR U16536 ( .A(n15965), .B(n15964), .Z(n15967) );
  NAND U16537 ( .A(a[18]), .B(b[15]), .Z(n16343) );
  XOR U16538 ( .A(n15965), .B(n15964), .Z(n16344) );
  NANDN U16539 ( .A(n16343), .B(n16344), .Z(n15966) );
  NAND U16540 ( .A(n15967), .B(n15966), .Z(n15970) );
  OR U16541 ( .A(n15971), .B(n15970), .Z(n15973) );
  XOR U16542 ( .A(n15969), .B(n15968), .Z(n16236) );
  XOR U16543 ( .A(n15971), .B(n15970), .Z(n16237) );
  NAND U16544 ( .A(n16236), .B(n16237), .Z(n15972) );
  NAND U16545 ( .A(n15973), .B(n15972), .Z(n15975) );
  NANDN U16546 ( .A(n15974), .B(n15975), .Z(n15977) );
  ANDN U16547 ( .B(b[15]), .A(n176), .Z(n16354) );
  XOR U16548 ( .A(n15975), .B(n15974), .Z(n16353) );
  OR U16549 ( .A(n16354), .B(n16353), .Z(n15976) );
  NAND U16550 ( .A(n15977), .B(n15976), .Z(n15979) );
  NANDN U16551 ( .A(n15978), .B(n15979), .Z(n15983) );
  XOR U16552 ( .A(n15979), .B(n15978), .Z(n16235) );
  XOR U16553 ( .A(n15981), .B(n15980), .Z(n16234) );
  NANDN U16554 ( .A(n16235), .B(n16234), .Z(n15982) );
  AND U16555 ( .A(n15983), .B(n15982), .Z(n15984) );
  OR U16556 ( .A(n15985), .B(n15984), .Z(n15987) );
  ANDN U16557 ( .B(b[15]), .A(n177), .Z(n16366) );
  XNOR U16558 ( .A(n15985), .B(n15984), .Z(n16365) );
  OR U16559 ( .A(n16366), .B(n16365), .Z(n15986) );
  NAND U16560 ( .A(n15987), .B(n15986), .Z(n15988) );
  NANDN U16561 ( .A(n15989), .B(n15988), .Z(n15993) );
  XOR U16562 ( .A(n15991), .B(n15990), .Z(n16369) );
  NANDN U16563 ( .A(n16370), .B(n16369), .Z(n15992) );
  NAND U16564 ( .A(n15993), .B(n15992), .Z(n15996) );
  XOR U16565 ( .A(n15995), .B(n15994), .Z(n15997) );
  NANDN U16566 ( .A(n15996), .B(n15997), .Z(n15999) );
  NAND U16567 ( .A(a[24]), .B(b[15]), .Z(n16375) );
  XNOR U16568 ( .A(n15997), .B(n15996), .Z(n16376) );
  NANDN U16569 ( .A(n16375), .B(n16376), .Z(n15998) );
  NAND U16570 ( .A(n15999), .B(n15998), .Z(n16000) );
  OR U16571 ( .A(n16001), .B(n16000), .Z(n16005) );
  XNOR U16572 ( .A(n16001), .B(n16000), .Z(n16381) );
  XOR U16573 ( .A(n16003), .B(n16002), .Z(n16382) );
  NANDN U16574 ( .A(n16381), .B(n16382), .Z(n16004) );
  NAND U16575 ( .A(n16005), .B(n16004), .Z(n16008) );
  XOR U16576 ( .A(n16007), .B(n16006), .Z(n16009) );
  NANDN U16577 ( .A(n16008), .B(n16009), .Z(n16011) );
  NAND U16578 ( .A(a[26]), .B(b[15]), .Z(n16387) );
  XNOR U16579 ( .A(n16009), .B(n16008), .Z(n16388) );
  NANDN U16580 ( .A(n16387), .B(n16388), .Z(n16010) );
  NAND U16581 ( .A(n16011), .B(n16010), .Z(n16012) );
  OR U16582 ( .A(n16013), .B(n16012), .Z(n16017) );
  XNOR U16583 ( .A(n16013), .B(n16012), .Z(n16393) );
  XOR U16584 ( .A(n16015), .B(n16014), .Z(n16394) );
  NANDN U16585 ( .A(n16393), .B(n16394), .Z(n16016) );
  NAND U16586 ( .A(n16017), .B(n16016), .Z(n16020) );
  XOR U16587 ( .A(n16019), .B(n16018), .Z(n16021) );
  NANDN U16588 ( .A(n16020), .B(n16021), .Z(n16023) );
  NAND U16589 ( .A(a[28]), .B(b[15]), .Z(n16399) );
  XNOR U16590 ( .A(n16021), .B(n16020), .Z(n16400) );
  NANDN U16591 ( .A(n16399), .B(n16400), .Z(n16022) );
  NAND U16592 ( .A(n16023), .B(n16022), .Z(n16024) );
  OR U16593 ( .A(n16025), .B(n16024), .Z(n16029) );
  XNOR U16594 ( .A(n16025), .B(n16024), .Z(n16405) );
  XOR U16595 ( .A(n16027), .B(n16026), .Z(n16406) );
  NANDN U16596 ( .A(n16405), .B(n16406), .Z(n16028) );
  NAND U16597 ( .A(n16029), .B(n16028), .Z(n16032) );
  XOR U16598 ( .A(n16031), .B(n16030), .Z(n16033) );
  NANDN U16599 ( .A(n16032), .B(n16033), .Z(n16035) );
  NAND U16600 ( .A(a[30]), .B(b[15]), .Z(n16411) );
  XNOR U16601 ( .A(n16033), .B(n16032), .Z(n16412) );
  NANDN U16602 ( .A(n16411), .B(n16412), .Z(n16034) );
  NAND U16603 ( .A(n16035), .B(n16034), .Z(n16036) );
  OR U16604 ( .A(n16037), .B(n16036), .Z(n16041) );
  XNOR U16605 ( .A(n16037), .B(n16036), .Z(n16417) );
  XOR U16606 ( .A(n16039), .B(n16038), .Z(n16418) );
  NANDN U16607 ( .A(n16417), .B(n16418), .Z(n16040) );
  NAND U16608 ( .A(n16041), .B(n16040), .Z(n16044) );
  XOR U16609 ( .A(n16043), .B(n16042), .Z(n16045) );
  NANDN U16610 ( .A(n16044), .B(n16045), .Z(n16047) );
  NAND U16611 ( .A(a[32]), .B(b[15]), .Z(n16423) );
  XNOR U16612 ( .A(n16045), .B(n16044), .Z(n16424) );
  NANDN U16613 ( .A(n16423), .B(n16424), .Z(n16046) );
  NAND U16614 ( .A(n16047), .B(n16046), .Z(n16048) );
  OR U16615 ( .A(n16049), .B(n16048), .Z(n16053) );
  XNOR U16616 ( .A(n16049), .B(n16048), .Z(n16429) );
  XOR U16617 ( .A(n16051), .B(n16050), .Z(n16430) );
  NANDN U16618 ( .A(n16429), .B(n16430), .Z(n16052) );
  NAND U16619 ( .A(n16053), .B(n16052), .Z(n16056) );
  XOR U16620 ( .A(n16055), .B(n16054), .Z(n16057) );
  NANDN U16621 ( .A(n16056), .B(n16057), .Z(n16059) );
  NAND U16622 ( .A(a[34]), .B(b[15]), .Z(n16435) );
  XNOR U16623 ( .A(n16057), .B(n16056), .Z(n16436) );
  NANDN U16624 ( .A(n16435), .B(n16436), .Z(n16058) );
  NAND U16625 ( .A(n16059), .B(n16058), .Z(n16060) );
  OR U16626 ( .A(n16061), .B(n16060), .Z(n16065) );
  XNOR U16627 ( .A(n16061), .B(n16060), .Z(n16441) );
  XOR U16628 ( .A(n16063), .B(n16062), .Z(n16442) );
  NANDN U16629 ( .A(n16441), .B(n16442), .Z(n16064) );
  NAND U16630 ( .A(n16065), .B(n16064), .Z(n16068) );
  XOR U16631 ( .A(n16067), .B(n16066), .Z(n16069) );
  NANDN U16632 ( .A(n16068), .B(n16069), .Z(n16071) );
  NAND U16633 ( .A(a[36]), .B(b[15]), .Z(n16447) );
  XNOR U16634 ( .A(n16069), .B(n16068), .Z(n16448) );
  NANDN U16635 ( .A(n16447), .B(n16448), .Z(n16070) );
  NAND U16636 ( .A(n16071), .B(n16070), .Z(n16072) );
  OR U16637 ( .A(n16073), .B(n16072), .Z(n16077) );
  XNOR U16638 ( .A(n16073), .B(n16072), .Z(n16453) );
  XOR U16639 ( .A(n16075), .B(n16074), .Z(n16454) );
  NANDN U16640 ( .A(n16453), .B(n16454), .Z(n16076) );
  NAND U16641 ( .A(n16077), .B(n16076), .Z(n16080) );
  XOR U16642 ( .A(n16079), .B(n16078), .Z(n16081) );
  NANDN U16643 ( .A(n16080), .B(n16081), .Z(n16083) );
  NAND U16644 ( .A(a[38]), .B(b[15]), .Z(n16459) );
  XNOR U16645 ( .A(n16081), .B(n16080), .Z(n16460) );
  NANDN U16646 ( .A(n16459), .B(n16460), .Z(n16082) );
  NAND U16647 ( .A(n16083), .B(n16082), .Z(n16084) );
  OR U16648 ( .A(n16085), .B(n16084), .Z(n16089) );
  XNOR U16649 ( .A(n16085), .B(n16084), .Z(n16465) );
  XOR U16650 ( .A(n16087), .B(n16086), .Z(n16466) );
  NANDN U16651 ( .A(n16465), .B(n16466), .Z(n16088) );
  NAND U16652 ( .A(n16089), .B(n16088), .Z(n16092) );
  XOR U16653 ( .A(n16091), .B(n16090), .Z(n16093) );
  NANDN U16654 ( .A(n16092), .B(n16093), .Z(n16095) );
  NAND U16655 ( .A(a[40]), .B(b[15]), .Z(n16471) );
  XNOR U16656 ( .A(n16093), .B(n16092), .Z(n16472) );
  NANDN U16657 ( .A(n16471), .B(n16472), .Z(n16094) );
  NAND U16658 ( .A(n16095), .B(n16094), .Z(n16096) );
  OR U16659 ( .A(n16097), .B(n16096), .Z(n16101) );
  XNOR U16660 ( .A(n16097), .B(n16096), .Z(n16477) );
  XOR U16661 ( .A(n16099), .B(n16098), .Z(n16478) );
  NANDN U16662 ( .A(n16477), .B(n16478), .Z(n16100) );
  NAND U16663 ( .A(n16101), .B(n16100), .Z(n16104) );
  XOR U16664 ( .A(n16103), .B(n16102), .Z(n16105) );
  NANDN U16665 ( .A(n16104), .B(n16105), .Z(n16107) );
  NAND U16666 ( .A(a[42]), .B(b[15]), .Z(n16483) );
  XNOR U16667 ( .A(n16105), .B(n16104), .Z(n16484) );
  NANDN U16668 ( .A(n16483), .B(n16484), .Z(n16106) );
  NAND U16669 ( .A(n16107), .B(n16106), .Z(n16108) );
  OR U16670 ( .A(n16109), .B(n16108), .Z(n16113) );
  XNOR U16671 ( .A(n16109), .B(n16108), .Z(n16489) );
  XOR U16672 ( .A(n16111), .B(n16110), .Z(n16490) );
  NANDN U16673 ( .A(n16489), .B(n16490), .Z(n16112) );
  NAND U16674 ( .A(n16113), .B(n16112), .Z(n16116) );
  XOR U16675 ( .A(n16115), .B(n16114), .Z(n16117) );
  NANDN U16676 ( .A(n16116), .B(n16117), .Z(n16119) );
  NAND U16677 ( .A(a[44]), .B(b[15]), .Z(n16495) );
  XNOR U16678 ( .A(n16117), .B(n16116), .Z(n16496) );
  NANDN U16679 ( .A(n16495), .B(n16496), .Z(n16118) );
  NAND U16680 ( .A(n16119), .B(n16118), .Z(n16120) );
  OR U16681 ( .A(n16121), .B(n16120), .Z(n16125) );
  XNOR U16682 ( .A(n16121), .B(n16120), .Z(n16501) );
  XOR U16683 ( .A(n16123), .B(n16122), .Z(n16502) );
  NANDN U16684 ( .A(n16501), .B(n16502), .Z(n16124) );
  NAND U16685 ( .A(n16125), .B(n16124), .Z(n16128) );
  XOR U16686 ( .A(n16127), .B(n16126), .Z(n16129) );
  NANDN U16687 ( .A(n16128), .B(n16129), .Z(n16131) );
  NAND U16688 ( .A(a[46]), .B(b[15]), .Z(n16507) );
  XNOR U16689 ( .A(n16129), .B(n16128), .Z(n16508) );
  NANDN U16690 ( .A(n16507), .B(n16508), .Z(n16130) );
  NAND U16691 ( .A(n16131), .B(n16130), .Z(n16134) );
  ANDN U16692 ( .B(b[15]), .A(n195), .Z(n16135) );
  OR U16693 ( .A(n16134), .B(n16135), .Z(n16137) );
  XOR U16694 ( .A(n16133), .B(n16132), .Z(n16514) );
  XOR U16695 ( .A(n16135), .B(n16134), .Z(n16513) );
  NANDN U16696 ( .A(n16514), .B(n16513), .Z(n16136) );
  NAND U16697 ( .A(n16137), .B(n16136), .Z(n16140) );
  XNOR U16698 ( .A(n16139), .B(n16138), .Z(n16141) );
  OR U16699 ( .A(n16140), .B(n16141), .Z(n16143) );
  XNOR U16700 ( .A(n16141), .B(n16140), .Z(n16522) );
  NAND U16701 ( .A(a[48]), .B(b[15]), .Z(n16521) );
  OR U16702 ( .A(n16522), .B(n16521), .Z(n16142) );
  NAND U16703 ( .A(n16143), .B(n16142), .Z(n16144) );
  ANDN U16704 ( .B(b[15]), .A(n197), .Z(n16145) );
  OR U16705 ( .A(n16144), .B(n16145), .Z(n16149) );
  XOR U16706 ( .A(n16145), .B(n16144), .Z(n16525) );
  NAND U16707 ( .A(n16525), .B(n16526), .Z(n16148) );
  NAND U16708 ( .A(n16149), .B(n16148), .Z(n16153) );
  NAND U16709 ( .A(a[50]), .B(b[15]), .Z(n16152) );
  OR U16710 ( .A(n16153), .B(n16152), .Z(n16155) );
  XOR U16711 ( .A(n16151), .B(n16150), .Z(n16531) );
  XOR U16712 ( .A(n16153), .B(n16152), .Z(n16532) );
  NAND U16713 ( .A(n16531), .B(n16532), .Z(n16154) );
  NAND U16714 ( .A(n16155), .B(n16154), .Z(n16159) );
  XOR U16715 ( .A(n16157), .B(n16156), .Z(n16158) );
  NAND U16716 ( .A(n16159), .B(n16158), .Z(n16161) );
  XNOR U16717 ( .A(n16159), .B(n16158), .Z(n16538) );
  NAND U16718 ( .A(a[51]), .B(b[15]), .Z(n16537) );
  OR U16719 ( .A(n16538), .B(n16537), .Z(n16160) );
  NAND U16720 ( .A(n16161), .B(n16160), .Z(n16165) );
  NANDN U16721 ( .A(n16164), .B(n16165), .Z(n16167) );
  XNOR U16722 ( .A(n16163), .B(n16162), .Z(n16544) );
  XNOR U16723 ( .A(n16165), .B(n16164), .Z(n16543) );
  NANDN U16724 ( .A(n16544), .B(n16543), .Z(n16166) );
  NAND U16725 ( .A(n16167), .B(n16166), .Z(n16171) );
  XOR U16726 ( .A(n16169), .B(n16168), .Z(n16170) );
  NAND U16727 ( .A(n16171), .B(n16170), .Z(n16173) );
  XNOR U16728 ( .A(n16171), .B(n16170), .Z(n16550) );
  NAND U16729 ( .A(a[53]), .B(b[15]), .Z(n16549) );
  OR U16730 ( .A(n16550), .B(n16549), .Z(n16172) );
  NAND U16731 ( .A(n16173), .B(n16172), .Z(n16177) );
  NANDN U16732 ( .A(n16176), .B(n16177), .Z(n16179) );
  XNOR U16733 ( .A(n16175), .B(n16174), .Z(n16556) );
  XNOR U16734 ( .A(n16177), .B(n16176), .Z(n16555) );
  NANDN U16735 ( .A(n16556), .B(n16555), .Z(n16178) );
  NAND U16736 ( .A(n16179), .B(n16178), .Z(n16183) );
  XOR U16737 ( .A(n16181), .B(n16180), .Z(n16182) );
  NAND U16738 ( .A(n16183), .B(n16182), .Z(n16185) );
  XNOR U16739 ( .A(n16183), .B(n16182), .Z(n16562) );
  NAND U16740 ( .A(a[55]), .B(b[15]), .Z(n16561) );
  OR U16741 ( .A(n16562), .B(n16561), .Z(n16184) );
  NAND U16742 ( .A(n16185), .B(n16184), .Z(n16189) );
  NANDN U16743 ( .A(n16188), .B(n16189), .Z(n16191) );
  XNOR U16744 ( .A(n16187), .B(n16186), .Z(n16568) );
  XNOR U16745 ( .A(n16189), .B(n16188), .Z(n16567) );
  NANDN U16746 ( .A(n16568), .B(n16567), .Z(n16190) );
  NAND U16747 ( .A(n16191), .B(n16190), .Z(n16195) );
  XOR U16748 ( .A(n16193), .B(n16192), .Z(n16194) );
  NAND U16749 ( .A(n16195), .B(n16194), .Z(n16197) );
  XNOR U16750 ( .A(n16195), .B(n16194), .Z(n16574) );
  NAND U16751 ( .A(a[57]), .B(b[15]), .Z(n16573) );
  OR U16752 ( .A(n16574), .B(n16573), .Z(n16196) );
  NAND U16753 ( .A(n16197), .B(n16196), .Z(n16201) );
  NANDN U16754 ( .A(n16200), .B(n16201), .Z(n16203) );
  XNOR U16755 ( .A(n16199), .B(n16198), .Z(n16580) );
  XNOR U16756 ( .A(n16201), .B(n16200), .Z(n16579) );
  NANDN U16757 ( .A(n16580), .B(n16579), .Z(n16202) );
  NAND U16758 ( .A(n16203), .B(n16202), .Z(n16207) );
  XOR U16759 ( .A(n16205), .B(n16204), .Z(n16206) );
  NAND U16760 ( .A(n16207), .B(n16206), .Z(n16209) );
  XNOR U16761 ( .A(n16207), .B(n16206), .Z(n16586) );
  NAND U16762 ( .A(a[59]), .B(b[15]), .Z(n16585) );
  OR U16763 ( .A(n16586), .B(n16585), .Z(n16208) );
  NAND U16764 ( .A(n16209), .B(n16208), .Z(n16213) );
  NANDN U16765 ( .A(n16212), .B(n16213), .Z(n16215) );
  XNOR U16766 ( .A(n16211), .B(n16210), .Z(n16592) );
  XNOR U16767 ( .A(n16213), .B(n16212), .Z(n16591) );
  NANDN U16768 ( .A(n16592), .B(n16591), .Z(n16214) );
  NAND U16769 ( .A(n16215), .B(n16214), .Z(n16219) );
  XOR U16770 ( .A(n16217), .B(n16216), .Z(n16218) );
  NAND U16771 ( .A(n16219), .B(n16218), .Z(n16221) );
  XNOR U16772 ( .A(n16219), .B(n16218), .Z(n16598) );
  NAND U16773 ( .A(a[61]), .B(b[15]), .Z(n16597) );
  OR U16774 ( .A(n16598), .B(n16597), .Z(n16220) );
  NAND U16775 ( .A(n16221), .B(n16220), .Z(n16225) );
  NANDN U16776 ( .A(n16224), .B(n16225), .Z(n16227) );
  XNOR U16777 ( .A(n16223), .B(n16222), .Z(n16604) );
  XNOR U16778 ( .A(n16225), .B(n16224), .Z(n16603) );
  NANDN U16779 ( .A(n16604), .B(n16603), .Z(n16226) );
  NAND U16780 ( .A(n16227), .B(n16226), .Z(n16230) );
  XOR U16781 ( .A(n16229), .B(n16228), .Z(n16231) );
  AND U16782 ( .A(b[15]), .B(a[63]), .Z(n16610) );
  XOR U16783 ( .A(n16231), .B(n16230), .Z(n16609) );
  XNOR U16784 ( .A(n16233), .B(n16232), .Z(n16612) );
  NOR U16785 ( .A(n16611), .B(n16612), .Z(n21960) );
  NAND U16786 ( .A(a[52]), .B(b[14]), .Z(n16539) );
  ANDN U16787 ( .B(b[14]), .A(n195), .Z(n16510) );
  ANDN U16788 ( .B(b[14]), .A(n193), .Z(n16498) );
  ANDN U16789 ( .B(b[14]), .A(n191), .Z(n16486) );
  ANDN U16790 ( .B(b[14]), .A(n189), .Z(n16474) );
  ANDN U16791 ( .B(b[14]), .A(n187), .Z(n16462) );
  ANDN U16792 ( .B(b[14]), .A(n21772), .Z(n16450) );
  ANDN U16793 ( .B(b[14]), .A(n184), .Z(n16438) );
  ANDN U16794 ( .B(b[14]), .A(n21751), .Z(n16426) );
  ANDN U16795 ( .B(b[14]), .A(n21740), .Z(n16414) );
  ANDN U16796 ( .B(b[14]), .A(n21727), .Z(n16402) );
  ANDN U16797 ( .B(b[14]), .A(n21716), .Z(n16390) );
  ANDN U16798 ( .B(b[14]), .A(n21703), .Z(n16378) );
  ANDN U16799 ( .B(b[14]), .A(n21692), .Z(n16363) );
  XOR U16800 ( .A(n16235), .B(n16234), .Z(n16359) );
  ANDN U16801 ( .B(b[14]), .A(n21681), .Z(n16356) );
  ANDN U16802 ( .B(b[14]), .A(n21670), .Z(n16346) );
  ANDN U16803 ( .B(b[14]), .A(n174), .Z(n16334) );
  NAND U16804 ( .A(a[15]), .B(b[14]), .Z(n16320) );
  ANDN U16805 ( .B(b[14]), .A(n170), .Z(n16310) );
  NAND U16806 ( .A(a[12]), .B(b[14]), .Z(n16306) );
  NAND U16807 ( .A(a[11]), .B(b[14]), .Z(n16298) );
  NAND U16808 ( .A(a[9]), .B(b[14]), .Z(n16288) );
  ANDN U16809 ( .B(b[14]), .A(n166), .Z(n16274) );
  ANDN U16810 ( .B(b[14]), .A(n164), .Z(n16262) );
  ANDN U16811 ( .B(b[14]), .A(n21580), .Z(n16249) );
  NAND U16812 ( .A(b[15]), .B(a[1]), .Z(n16242) );
  AND U16813 ( .A(b[14]), .B(a[0]), .Z(n16994) );
  NANDN U16814 ( .A(n16242), .B(n16994), .Z(n16241) );
  NAND U16815 ( .A(a[2]), .B(b[14]), .Z(n16240) );
  AND U16816 ( .A(n16241), .B(n16240), .Z(n16248) );
  NANDN U16817 ( .A(n16242), .B(a[0]), .Z(n16243) );
  XNOR U16818 ( .A(a[2]), .B(n16243), .Z(n16244) );
  NAND U16819 ( .A(b[14]), .B(n16244), .Z(n16645) );
  AND U16820 ( .A(a[1]), .B(b[15]), .Z(n16245) );
  XNOR U16821 ( .A(n16246), .B(n16245), .Z(n16644) );
  NANDN U16822 ( .A(n16645), .B(n16644), .Z(n16247) );
  NANDN U16823 ( .A(n16248), .B(n16247), .Z(n16250) );
  NANDN U16824 ( .A(n16249), .B(n16250), .Z(n16254) );
  XOR U16825 ( .A(n16250), .B(n16249), .Z(n16649) );
  NANDN U16826 ( .A(n16649), .B(n16648), .Z(n16253) );
  NAND U16827 ( .A(n16254), .B(n16253), .Z(n16258) );
  XOR U16828 ( .A(n16256), .B(n16255), .Z(n16257) );
  NANDN U16829 ( .A(n16258), .B(n16257), .Z(n16260) );
  NAND U16830 ( .A(a[4]), .B(b[14]), .Z(n16656) );
  NANDN U16831 ( .A(n16656), .B(n16657), .Z(n16259) );
  NAND U16832 ( .A(n16260), .B(n16259), .Z(n16261) );
  OR U16833 ( .A(n16262), .B(n16261), .Z(n16266) );
  XNOR U16834 ( .A(n16262), .B(n16261), .Z(n16631) );
  XOR U16835 ( .A(n16264), .B(n16263), .Z(n16632) );
  NANDN U16836 ( .A(n16631), .B(n16632), .Z(n16265) );
  NAND U16837 ( .A(n16266), .B(n16265), .Z(n16269) );
  XOR U16838 ( .A(n16268), .B(n16267), .Z(n16270) );
  NANDN U16839 ( .A(n16269), .B(n16270), .Z(n16272) );
  NAND U16840 ( .A(a[6]), .B(b[14]), .Z(n16666) );
  XNOR U16841 ( .A(n16270), .B(n16269), .Z(n16667) );
  NANDN U16842 ( .A(n16666), .B(n16667), .Z(n16271) );
  NAND U16843 ( .A(n16272), .B(n16271), .Z(n16273) );
  OR U16844 ( .A(n16274), .B(n16273), .Z(n16278) );
  XNOR U16845 ( .A(n16274), .B(n16273), .Z(n16670) );
  XOR U16846 ( .A(n16276), .B(n16275), .Z(n16671) );
  NANDN U16847 ( .A(n16670), .B(n16671), .Z(n16277) );
  NAND U16848 ( .A(n16278), .B(n16277), .Z(n16281) );
  XOR U16849 ( .A(n16280), .B(n16279), .Z(n16282) );
  NANDN U16850 ( .A(n16281), .B(n16282), .Z(n16284) );
  NAND U16851 ( .A(a[8]), .B(b[14]), .Z(n16678) );
  XNOR U16852 ( .A(n16282), .B(n16281), .Z(n16679) );
  NANDN U16853 ( .A(n16678), .B(n16679), .Z(n16283) );
  NAND U16854 ( .A(n16284), .B(n16283), .Z(n16287) );
  NANDN U16855 ( .A(n16288), .B(n16287), .Z(n16290) );
  XOR U16856 ( .A(n16286), .B(n16285), .Z(n16685) );
  NANDN U16857 ( .A(n16685), .B(n16684), .Z(n16289) );
  AND U16858 ( .A(n16290), .B(n16289), .Z(n16293) );
  XOR U16859 ( .A(n16292), .B(n16291), .Z(n16294) );
  NANDN U16860 ( .A(n16293), .B(n16294), .Z(n16296) );
  NAND U16861 ( .A(a[10]), .B(b[14]), .Z(n16688) );
  XNOR U16862 ( .A(n16294), .B(n16293), .Z(n16689) );
  NANDN U16863 ( .A(n16688), .B(n16689), .Z(n16295) );
  NAND U16864 ( .A(n16296), .B(n16295), .Z(n16297) );
  NANDN U16865 ( .A(n16298), .B(n16297), .Z(n16302) );
  XNOR U16866 ( .A(n16300), .B(n16299), .Z(n16695) );
  NAND U16867 ( .A(n16694), .B(n16695), .Z(n16301) );
  NAND U16868 ( .A(n16302), .B(n16301), .Z(n16305) );
  NANDN U16869 ( .A(n16306), .B(n16305), .Z(n16308) );
  XOR U16870 ( .A(n16304), .B(n16303), .Z(n16701) );
  NAND U16871 ( .A(n16701), .B(n16700), .Z(n16307) );
  NAND U16872 ( .A(n16308), .B(n16307), .Z(n16309) );
  OR U16873 ( .A(n16310), .B(n16309), .Z(n16314) );
  XOR U16874 ( .A(n16310), .B(n16309), .Z(n16629) );
  XOR U16875 ( .A(n16312), .B(n16311), .Z(n16630) );
  NAND U16876 ( .A(n16629), .B(n16630), .Z(n16313) );
  AND U16877 ( .A(n16314), .B(n16313), .Z(n16315) );
  OR U16878 ( .A(n16316), .B(n16315), .Z(n16318) );
  ANDN U16879 ( .B(b[14]), .A(n171), .Z(n16711) );
  XOR U16880 ( .A(n16316), .B(n16315), .Z(n16710) );
  NANDN U16881 ( .A(n16711), .B(n16710), .Z(n16317) );
  AND U16882 ( .A(n16318), .B(n16317), .Z(n16319) );
  NANDN U16883 ( .A(n16320), .B(n16319), .Z(n16324) );
  XNOR U16884 ( .A(n16322), .B(n16321), .Z(n16628) );
  NAND U16885 ( .A(n16627), .B(n16628), .Z(n16323) );
  AND U16886 ( .A(n16324), .B(n16323), .Z(n16327) );
  XOR U16887 ( .A(n16326), .B(n16325), .Z(n16328) );
  NANDN U16888 ( .A(n16327), .B(n16328), .Z(n16330) );
  NAND U16889 ( .A(a[16]), .B(b[14]), .Z(n16720) );
  XNOR U16890 ( .A(n16328), .B(n16327), .Z(n16721) );
  NANDN U16891 ( .A(n16720), .B(n16721), .Z(n16329) );
  NAND U16892 ( .A(n16330), .B(n16329), .Z(n16333) );
  OR U16893 ( .A(n16334), .B(n16333), .Z(n16336) );
  XOR U16894 ( .A(n16332), .B(n16331), .Z(n16726) );
  XOR U16895 ( .A(n16334), .B(n16333), .Z(n16727) );
  NAND U16896 ( .A(n16726), .B(n16727), .Z(n16335) );
  NAND U16897 ( .A(n16336), .B(n16335), .Z(n16339) );
  XOR U16898 ( .A(n16338), .B(n16337), .Z(n16340) );
  NANDN U16899 ( .A(n16339), .B(n16340), .Z(n16342) );
  NAND U16900 ( .A(a[18]), .B(b[14]), .Z(n16732) );
  XNOR U16901 ( .A(n16340), .B(n16339), .Z(n16733) );
  NANDN U16902 ( .A(n16732), .B(n16733), .Z(n16341) );
  NAND U16903 ( .A(n16342), .B(n16341), .Z(n16345) );
  OR U16904 ( .A(n16346), .B(n16345), .Z(n16348) );
  XOR U16905 ( .A(n16344), .B(n16343), .Z(n16738) );
  XOR U16906 ( .A(n16346), .B(n16345), .Z(n16739) );
  NAND U16907 ( .A(n16738), .B(n16739), .Z(n16347) );
  NAND U16908 ( .A(n16348), .B(n16347), .Z(n16349) );
  OR U16909 ( .A(n16350), .B(n16349), .Z(n16352) );
  NAND U16910 ( .A(a[20]), .B(b[14]), .Z(n16744) );
  XOR U16911 ( .A(n16350), .B(n16349), .Z(n16745) );
  NANDN U16912 ( .A(n16744), .B(n16745), .Z(n16351) );
  NAND U16913 ( .A(n16352), .B(n16351), .Z(n16355) );
  OR U16914 ( .A(n16356), .B(n16355), .Z(n16358) );
  XOR U16915 ( .A(n16354), .B(n16353), .Z(n16625) );
  XOR U16916 ( .A(n16356), .B(n16355), .Z(n16626) );
  NAND U16917 ( .A(n16625), .B(n16626), .Z(n16357) );
  NAND U16918 ( .A(n16358), .B(n16357), .Z(n16360) );
  NANDN U16919 ( .A(n16359), .B(n16360), .Z(n16362) );
  ANDN U16920 ( .B(b[14]), .A(n177), .Z(n16757) );
  XOR U16921 ( .A(n16360), .B(n16359), .Z(n16756) );
  OR U16922 ( .A(n16757), .B(n16756), .Z(n16361) );
  NAND U16923 ( .A(n16362), .B(n16361), .Z(n16364) );
  NANDN U16924 ( .A(n16363), .B(n16364), .Z(n16368) );
  XOR U16925 ( .A(n16364), .B(n16363), .Z(n16624) );
  XOR U16926 ( .A(n16366), .B(n16365), .Z(n16623) );
  NANDN U16927 ( .A(n16624), .B(n16623), .Z(n16367) );
  NAND U16928 ( .A(n16368), .B(n16367), .Z(n16371) );
  NANDN U16929 ( .A(n16371), .B(n16372), .Z(n16374) );
  NAND U16930 ( .A(a[24]), .B(b[14]), .Z(n16764) );
  XNOR U16931 ( .A(n16372), .B(n16371), .Z(n16765) );
  NANDN U16932 ( .A(n16764), .B(n16765), .Z(n16373) );
  NAND U16933 ( .A(n16374), .B(n16373), .Z(n16377) );
  OR U16934 ( .A(n16378), .B(n16377), .Z(n16380) );
  XOR U16935 ( .A(n16376), .B(n16375), .Z(n16770) );
  XOR U16936 ( .A(n16378), .B(n16377), .Z(n16771) );
  NAND U16937 ( .A(n16770), .B(n16771), .Z(n16379) );
  NAND U16938 ( .A(n16380), .B(n16379), .Z(n16383) );
  XOR U16939 ( .A(n16382), .B(n16381), .Z(n16384) );
  NANDN U16940 ( .A(n16383), .B(n16384), .Z(n16386) );
  NAND U16941 ( .A(a[26]), .B(b[14]), .Z(n16776) );
  XNOR U16942 ( .A(n16384), .B(n16383), .Z(n16777) );
  NANDN U16943 ( .A(n16776), .B(n16777), .Z(n16385) );
  NAND U16944 ( .A(n16386), .B(n16385), .Z(n16389) );
  OR U16945 ( .A(n16390), .B(n16389), .Z(n16392) );
  XOR U16946 ( .A(n16388), .B(n16387), .Z(n16782) );
  XOR U16947 ( .A(n16390), .B(n16389), .Z(n16783) );
  NAND U16948 ( .A(n16782), .B(n16783), .Z(n16391) );
  NAND U16949 ( .A(n16392), .B(n16391), .Z(n16395) );
  XOR U16950 ( .A(n16394), .B(n16393), .Z(n16396) );
  NANDN U16951 ( .A(n16395), .B(n16396), .Z(n16398) );
  NAND U16952 ( .A(a[28]), .B(b[14]), .Z(n16788) );
  XNOR U16953 ( .A(n16396), .B(n16395), .Z(n16789) );
  NANDN U16954 ( .A(n16788), .B(n16789), .Z(n16397) );
  NAND U16955 ( .A(n16398), .B(n16397), .Z(n16401) );
  OR U16956 ( .A(n16402), .B(n16401), .Z(n16404) );
  XOR U16957 ( .A(n16400), .B(n16399), .Z(n16794) );
  XOR U16958 ( .A(n16402), .B(n16401), .Z(n16795) );
  NAND U16959 ( .A(n16794), .B(n16795), .Z(n16403) );
  NAND U16960 ( .A(n16404), .B(n16403), .Z(n16407) );
  XOR U16961 ( .A(n16406), .B(n16405), .Z(n16408) );
  NANDN U16962 ( .A(n16407), .B(n16408), .Z(n16410) );
  NAND U16963 ( .A(a[30]), .B(b[14]), .Z(n16800) );
  XNOR U16964 ( .A(n16408), .B(n16407), .Z(n16801) );
  NANDN U16965 ( .A(n16800), .B(n16801), .Z(n16409) );
  NAND U16966 ( .A(n16410), .B(n16409), .Z(n16413) );
  OR U16967 ( .A(n16414), .B(n16413), .Z(n16416) );
  XOR U16968 ( .A(n16412), .B(n16411), .Z(n16806) );
  XOR U16969 ( .A(n16414), .B(n16413), .Z(n16807) );
  NAND U16970 ( .A(n16806), .B(n16807), .Z(n16415) );
  NAND U16971 ( .A(n16416), .B(n16415), .Z(n16419) );
  XOR U16972 ( .A(n16418), .B(n16417), .Z(n16420) );
  NANDN U16973 ( .A(n16419), .B(n16420), .Z(n16422) );
  NAND U16974 ( .A(a[32]), .B(b[14]), .Z(n16812) );
  XNOR U16975 ( .A(n16420), .B(n16419), .Z(n16813) );
  NANDN U16976 ( .A(n16812), .B(n16813), .Z(n16421) );
  NAND U16977 ( .A(n16422), .B(n16421), .Z(n16425) );
  OR U16978 ( .A(n16426), .B(n16425), .Z(n16428) );
  XOR U16979 ( .A(n16424), .B(n16423), .Z(n16818) );
  XOR U16980 ( .A(n16426), .B(n16425), .Z(n16819) );
  NAND U16981 ( .A(n16818), .B(n16819), .Z(n16427) );
  NAND U16982 ( .A(n16428), .B(n16427), .Z(n16431) );
  XOR U16983 ( .A(n16430), .B(n16429), .Z(n16432) );
  NANDN U16984 ( .A(n16431), .B(n16432), .Z(n16434) );
  NAND U16985 ( .A(a[34]), .B(b[14]), .Z(n16824) );
  XNOR U16986 ( .A(n16432), .B(n16431), .Z(n16825) );
  NANDN U16987 ( .A(n16824), .B(n16825), .Z(n16433) );
  NAND U16988 ( .A(n16434), .B(n16433), .Z(n16437) );
  OR U16989 ( .A(n16438), .B(n16437), .Z(n16440) );
  XOR U16990 ( .A(n16436), .B(n16435), .Z(n16830) );
  XOR U16991 ( .A(n16438), .B(n16437), .Z(n16831) );
  NAND U16992 ( .A(n16830), .B(n16831), .Z(n16439) );
  NAND U16993 ( .A(n16440), .B(n16439), .Z(n16443) );
  XOR U16994 ( .A(n16442), .B(n16441), .Z(n16444) );
  NANDN U16995 ( .A(n16443), .B(n16444), .Z(n16446) );
  NAND U16996 ( .A(a[36]), .B(b[14]), .Z(n16836) );
  XNOR U16997 ( .A(n16444), .B(n16443), .Z(n16837) );
  NANDN U16998 ( .A(n16836), .B(n16837), .Z(n16445) );
  NAND U16999 ( .A(n16446), .B(n16445), .Z(n16449) );
  OR U17000 ( .A(n16450), .B(n16449), .Z(n16452) );
  XOR U17001 ( .A(n16448), .B(n16447), .Z(n16842) );
  XOR U17002 ( .A(n16450), .B(n16449), .Z(n16843) );
  NAND U17003 ( .A(n16842), .B(n16843), .Z(n16451) );
  NAND U17004 ( .A(n16452), .B(n16451), .Z(n16455) );
  XOR U17005 ( .A(n16454), .B(n16453), .Z(n16456) );
  NANDN U17006 ( .A(n16455), .B(n16456), .Z(n16458) );
  NAND U17007 ( .A(a[38]), .B(b[14]), .Z(n16848) );
  XNOR U17008 ( .A(n16456), .B(n16455), .Z(n16849) );
  NANDN U17009 ( .A(n16848), .B(n16849), .Z(n16457) );
  NAND U17010 ( .A(n16458), .B(n16457), .Z(n16461) );
  OR U17011 ( .A(n16462), .B(n16461), .Z(n16464) );
  XOR U17012 ( .A(n16460), .B(n16459), .Z(n16854) );
  XOR U17013 ( .A(n16462), .B(n16461), .Z(n16855) );
  NAND U17014 ( .A(n16854), .B(n16855), .Z(n16463) );
  NAND U17015 ( .A(n16464), .B(n16463), .Z(n16467) );
  XOR U17016 ( .A(n16466), .B(n16465), .Z(n16468) );
  NANDN U17017 ( .A(n16467), .B(n16468), .Z(n16470) );
  NAND U17018 ( .A(a[40]), .B(b[14]), .Z(n16860) );
  XNOR U17019 ( .A(n16468), .B(n16467), .Z(n16861) );
  NANDN U17020 ( .A(n16860), .B(n16861), .Z(n16469) );
  NAND U17021 ( .A(n16470), .B(n16469), .Z(n16473) );
  OR U17022 ( .A(n16474), .B(n16473), .Z(n16476) );
  XOR U17023 ( .A(n16472), .B(n16471), .Z(n16866) );
  XOR U17024 ( .A(n16474), .B(n16473), .Z(n16867) );
  NAND U17025 ( .A(n16866), .B(n16867), .Z(n16475) );
  NAND U17026 ( .A(n16476), .B(n16475), .Z(n16479) );
  XOR U17027 ( .A(n16478), .B(n16477), .Z(n16480) );
  NANDN U17028 ( .A(n16479), .B(n16480), .Z(n16482) );
  NAND U17029 ( .A(a[42]), .B(b[14]), .Z(n16872) );
  XNOR U17030 ( .A(n16480), .B(n16479), .Z(n16873) );
  NANDN U17031 ( .A(n16872), .B(n16873), .Z(n16481) );
  NAND U17032 ( .A(n16482), .B(n16481), .Z(n16485) );
  OR U17033 ( .A(n16486), .B(n16485), .Z(n16488) );
  XOR U17034 ( .A(n16484), .B(n16483), .Z(n16878) );
  XOR U17035 ( .A(n16486), .B(n16485), .Z(n16879) );
  NAND U17036 ( .A(n16878), .B(n16879), .Z(n16487) );
  NAND U17037 ( .A(n16488), .B(n16487), .Z(n16491) );
  XOR U17038 ( .A(n16490), .B(n16489), .Z(n16492) );
  NANDN U17039 ( .A(n16491), .B(n16492), .Z(n16494) );
  NAND U17040 ( .A(a[44]), .B(b[14]), .Z(n16884) );
  XNOR U17041 ( .A(n16492), .B(n16491), .Z(n16885) );
  NANDN U17042 ( .A(n16884), .B(n16885), .Z(n16493) );
  NAND U17043 ( .A(n16494), .B(n16493), .Z(n16497) );
  OR U17044 ( .A(n16498), .B(n16497), .Z(n16500) );
  XOR U17045 ( .A(n16496), .B(n16495), .Z(n16890) );
  XOR U17046 ( .A(n16498), .B(n16497), .Z(n16891) );
  NAND U17047 ( .A(n16890), .B(n16891), .Z(n16499) );
  NAND U17048 ( .A(n16500), .B(n16499), .Z(n16503) );
  XOR U17049 ( .A(n16502), .B(n16501), .Z(n16504) );
  NANDN U17050 ( .A(n16503), .B(n16504), .Z(n16506) );
  NAND U17051 ( .A(a[46]), .B(b[14]), .Z(n16896) );
  XNOR U17052 ( .A(n16504), .B(n16503), .Z(n16897) );
  NANDN U17053 ( .A(n16896), .B(n16897), .Z(n16505) );
  NAND U17054 ( .A(n16506), .B(n16505), .Z(n16509) );
  OR U17055 ( .A(n16510), .B(n16509), .Z(n16512) );
  XOR U17056 ( .A(n16508), .B(n16507), .Z(n16902) );
  XOR U17057 ( .A(n16510), .B(n16509), .Z(n16903) );
  NAND U17058 ( .A(n16902), .B(n16903), .Z(n16511) );
  NAND U17059 ( .A(n16512), .B(n16511), .Z(n16515) );
  XNOR U17060 ( .A(n16514), .B(n16513), .Z(n16516) );
  OR U17061 ( .A(n16515), .B(n16516), .Z(n16518) );
  XNOR U17062 ( .A(n16516), .B(n16515), .Z(n16911) );
  ANDN U17063 ( .B(b[14]), .A(n196), .Z(n16910) );
  NANDN U17064 ( .A(n16911), .B(n16910), .Z(n16517) );
  NAND U17065 ( .A(n16518), .B(n16517), .Z(n16519) );
  ANDN U17066 ( .B(b[14]), .A(n197), .Z(n16520) );
  OR U17067 ( .A(n16519), .B(n16520), .Z(n16524) );
  XNOR U17068 ( .A(n16520), .B(n16519), .Z(n16914) );
  XOR U17069 ( .A(n16522), .B(n16521), .Z(n16915) );
  OR U17070 ( .A(n16914), .B(n16915), .Z(n16523) );
  NAND U17071 ( .A(n16524), .B(n16523), .Z(n16528) );
  AND U17072 ( .A(b[14]), .B(a[50]), .Z(n16527) );
  NANDN U17073 ( .A(n16528), .B(n16527), .Z(n16530) );
  XNOR U17074 ( .A(n16528), .B(n16527), .Z(n16922) );
  NANDN U17075 ( .A(n16923), .B(n16922), .Z(n16529) );
  NAND U17076 ( .A(n16530), .B(n16529), .Z(n16534) );
  XOR U17077 ( .A(n16532), .B(n16531), .Z(n16533) );
  NAND U17078 ( .A(n16534), .B(n16533), .Z(n16536) );
  XNOR U17079 ( .A(n16534), .B(n16533), .Z(n16929) );
  NAND U17080 ( .A(a[51]), .B(b[14]), .Z(n16928) );
  OR U17081 ( .A(n16929), .B(n16928), .Z(n16535) );
  NAND U17082 ( .A(n16536), .B(n16535), .Z(n16540) );
  NANDN U17083 ( .A(n16539), .B(n16540), .Z(n16542) );
  XOR U17084 ( .A(n16538), .B(n16537), .Z(n16621) );
  XNOR U17085 ( .A(n16540), .B(n16539), .Z(n16622) );
  NAND U17086 ( .A(n16621), .B(n16622), .Z(n16541) );
  NAND U17087 ( .A(n16542), .B(n16541), .Z(n16545) );
  AND U17088 ( .A(b[14]), .B(a[53]), .Z(n16546) );
  OR U17089 ( .A(n16545), .B(n16546), .Z(n16548) );
  XNOR U17090 ( .A(n16544), .B(n16543), .Z(n16939) );
  XOR U17091 ( .A(n16546), .B(n16545), .Z(n16938) );
  NANDN U17092 ( .A(n16939), .B(n16938), .Z(n16547) );
  NAND U17093 ( .A(n16548), .B(n16547), .Z(n16552) );
  NAND U17094 ( .A(a[54]), .B(b[14]), .Z(n16551) );
  OR U17095 ( .A(n16552), .B(n16551), .Z(n16554) );
  XOR U17096 ( .A(n16550), .B(n16549), .Z(n16619) );
  XOR U17097 ( .A(n16552), .B(n16551), .Z(n16620) );
  NAND U17098 ( .A(n16619), .B(n16620), .Z(n16553) );
  NAND U17099 ( .A(n16554), .B(n16553), .Z(n16557) );
  AND U17100 ( .A(b[14]), .B(a[55]), .Z(n16558) );
  OR U17101 ( .A(n16557), .B(n16558), .Z(n16560) );
  XNOR U17102 ( .A(n16556), .B(n16555), .Z(n16949) );
  XOR U17103 ( .A(n16558), .B(n16557), .Z(n16948) );
  NANDN U17104 ( .A(n16949), .B(n16948), .Z(n16559) );
  NAND U17105 ( .A(n16560), .B(n16559), .Z(n16564) );
  NAND U17106 ( .A(a[56]), .B(b[14]), .Z(n16563) );
  OR U17107 ( .A(n16564), .B(n16563), .Z(n16566) );
  XOR U17108 ( .A(n16562), .B(n16561), .Z(n16617) );
  XOR U17109 ( .A(n16564), .B(n16563), .Z(n16618) );
  NAND U17110 ( .A(n16617), .B(n16618), .Z(n16565) );
  NAND U17111 ( .A(n16566), .B(n16565), .Z(n16569) );
  AND U17112 ( .A(b[14]), .B(a[57]), .Z(n16570) );
  OR U17113 ( .A(n16569), .B(n16570), .Z(n16572) );
  XNOR U17114 ( .A(n16568), .B(n16567), .Z(n16959) );
  XOR U17115 ( .A(n16570), .B(n16569), .Z(n16958) );
  NANDN U17116 ( .A(n16959), .B(n16958), .Z(n16571) );
  NAND U17117 ( .A(n16572), .B(n16571), .Z(n16576) );
  NAND U17118 ( .A(a[58]), .B(b[14]), .Z(n16575) );
  OR U17119 ( .A(n16576), .B(n16575), .Z(n16578) );
  XOR U17120 ( .A(n16574), .B(n16573), .Z(n16615) );
  XOR U17121 ( .A(n16576), .B(n16575), .Z(n16616) );
  NAND U17122 ( .A(n16615), .B(n16616), .Z(n16577) );
  NAND U17123 ( .A(n16578), .B(n16577), .Z(n16581) );
  AND U17124 ( .A(b[14]), .B(a[59]), .Z(n16582) );
  OR U17125 ( .A(n16581), .B(n16582), .Z(n16584) );
  XNOR U17126 ( .A(n16580), .B(n16579), .Z(n16969) );
  XOR U17127 ( .A(n16582), .B(n16581), .Z(n16968) );
  NANDN U17128 ( .A(n16969), .B(n16968), .Z(n16583) );
  NAND U17129 ( .A(n16584), .B(n16583), .Z(n16588) );
  NAND U17130 ( .A(a[60]), .B(b[14]), .Z(n16587) );
  OR U17131 ( .A(n16588), .B(n16587), .Z(n16590) );
  XOR U17132 ( .A(n16586), .B(n16585), .Z(n16972) );
  XOR U17133 ( .A(n16588), .B(n16587), .Z(n16973) );
  NAND U17134 ( .A(n16972), .B(n16973), .Z(n16589) );
  NAND U17135 ( .A(n16590), .B(n16589), .Z(n16593) );
  AND U17136 ( .A(b[14]), .B(a[61]), .Z(n16594) );
  OR U17137 ( .A(n16593), .B(n16594), .Z(n16596) );
  XNOR U17138 ( .A(n16592), .B(n16591), .Z(n16981) );
  XOR U17139 ( .A(n16594), .B(n16593), .Z(n16980) );
  NANDN U17140 ( .A(n16981), .B(n16980), .Z(n16595) );
  NAND U17141 ( .A(n16596), .B(n16595), .Z(n16600) );
  NAND U17142 ( .A(a[62]), .B(b[14]), .Z(n16599) );
  OR U17143 ( .A(n16600), .B(n16599), .Z(n16602) );
  XOR U17144 ( .A(n16598), .B(n16597), .Z(n16982) );
  XOR U17145 ( .A(n16600), .B(n16599), .Z(n16983) );
  NAND U17146 ( .A(n16982), .B(n16983), .Z(n16601) );
  NAND U17147 ( .A(n16602), .B(n16601), .Z(n16605) );
  AND U17148 ( .A(b[14]), .B(a[63]), .Z(n16606) );
  OR U17149 ( .A(n16605), .B(n16606), .Z(n16608) );
  XNOR U17150 ( .A(n16604), .B(n16603), .Z(n17360) );
  XOR U17151 ( .A(n16606), .B(n16605), .Z(n17359) );
  NANDN U17152 ( .A(n17360), .B(n17359), .Z(n16607) );
  NAND U17153 ( .A(n16608), .B(n16607), .Z(n21956) );
  XOR U17154 ( .A(n16610), .B(n16609), .Z(n21957) );
  NANDN U17155 ( .A(n21956), .B(n21957), .Z(n16614) );
  XOR U17156 ( .A(n16612), .B(n16611), .Z(n16613) );
  NANDN U17157 ( .A(n16614), .B(n16613), .Z(n21959) );
  XOR U17158 ( .A(n16614), .B(n16613), .Z(n24144) );
  NAND U17159 ( .A(a[62]), .B(b[13]), .Z(n16978) );
  NAND U17160 ( .A(a[60]), .B(b[13]), .Z(n16966) );
  XOR U17161 ( .A(n16616), .B(n16615), .Z(n16962) );
  NAND U17162 ( .A(a[58]), .B(b[13]), .Z(n16956) );
  XOR U17163 ( .A(n16618), .B(n16617), .Z(n16952) );
  NAND U17164 ( .A(a[56]), .B(b[13]), .Z(n16946) );
  XOR U17165 ( .A(n16620), .B(n16619), .Z(n16942) );
  NAND U17166 ( .A(a[54]), .B(b[13]), .Z(n16936) );
  XOR U17167 ( .A(n16622), .B(n16621), .Z(n16932) );
  ANDN U17168 ( .B(b[13]), .A(n195), .Z(n16899) );
  ANDN U17169 ( .B(b[13]), .A(n193), .Z(n16887) );
  ANDN U17170 ( .B(b[13]), .A(n191), .Z(n16875) );
  ANDN U17171 ( .B(b[13]), .A(n189), .Z(n16863) );
  ANDN U17172 ( .B(b[13]), .A(n187), .Z(n16851) );
  ANDN U17173 ( .B(b[13]), .A(n21772), .Z(n16839) );
  ANDN U17174 ( .B(b[13]), .A(n184), .Z(n16827) );
  ANDN U17175 ( .B(b[13]), .A(n21751), .Z(n16815) );
  ANDN U17176 ( .B(b[13]), .A(n21740), .Z(n16803) );
  ANDN U17177 ( .B(b[13]), .A(n21727), .Z(n16791) );
  ANDN U17178 ( .B(b[13]), .A(n21716), .Z(n16779) );
  XOR U17179 ( .A(n16624), .B(n16623), .Z(n16760) );
  ANDN U17180 ( .B(b[13]), .A(n21692), .Z(n16755) );
  ANDN U17181 ( .B(b[13]), .A(n21681), .Z(n16747) );
  ANDN U17182 ( .B(b[13]), .A(n21670), .Z(n16735) );
  ANDN U17183 ( .B(b[13]), .A(n172), .Z(n16713) );
  ANDN U17184 ( .B(b[13]), .A(n170), .Z(n16703) );
  NAND U17185 ( .A(a[11]), .B(b[13]), .Z(n16691) );
  ANDN U17186 ( .B(b[13]), .A(n21615), .Z(n16677) );
  ANDN U17187 ( .B(b[13]), .A(n166), .Z(n16665) );
  NAND U17188 ( .A(a[6]), .B(b[13]), .Z(n16660) );
  XOR U17189 ( .A(n16632), .B(n16631), .Z(n16661) );
  NANDN U17190 ( .A(n16660), .B(n16661), .Z(n16663) );
  ANDN U17191 ( .B(b[13]), .A(n164), .Z(n16655) );
  ANDN U17192 ( .B(b[13]), .A(n21580), .Z(n16642) );
  NAND U17193 ( .A(b[14]), .B(a[1]), .Z(n16635) );
  AND U17194 ( .A(b[13]), .B(a[0]), .Z(n17379) );
  NANDN U17195 ( .A(n16635), .B(n17379), .Z(n16634) );
  NAND U17196 ( .A(b[13]), .B(a[2]), .Z(n16633) );
  AND U17197 ( .A(n16634), .B(n16633), .Z(n16641) );
  NANDN U17198 ( .A(n16635), .B(a[0]), .Z(n16636) );
  XNOR U17199 ( .A(a[2]), .B(n16636), .Z(n16637) );
  NAND U17200 ( .A(b[13]), .B(n16637), .Z(n17000) );
  AND U17201 ( .A(a[1]), .B(b[14]), .Z(n16638) );
  XNOR U17202 ( .A(n16639), .B(n16638), .Z(n16999) );
  NANDN U17203 ( .A(n17000), .B(n16999), .Z(n16640) );
  NANDN U17204 ( .A(n16641), .B(n16640), .Z(n16643) );
  NANDN U17205 ( .A(n16642), .B(n16643), .Z(n16647) );
  XOR U17206 ( .A(n16643), .B(n16642), .Z(n17004) );
  NANDN U17207 ( .A(n17004), .B(n17003), .Z(n16646) );
  NAND U17208 ( .A(n16647), .B(n16646), .Z(n16651) );
  XOR U17209 ( .A(n16649), .B(n16648), .Z(n16650) );
  NANDN U17210 ( .A(n16651), .B(n16650), .Z(n16653) );
  NAND U17211 ( .A(a[4]), .B(b[13]), .Z(n17011) );
  NANDN U17212 ( .A(n17011), .B(n17012), .Z(n16652) );
  NAND U17213 ( .A(n16653), .B(n16652), .Z(n16654) );
  OR U17214 ( .A(n16655), .B(n16654), .Z(n16659) );
  XNOR U17215 ( .A(n16655), .B(n16654), .Z(n16986) );
  XOR U17216 ( .A(n16657), .B(n16656), .Z(n16987) );
  NANDN U17217 ( .A(n16986), .B(n16987), .Z(n16658) );
  NAND U17218 ( .A(n16659), .B(n16658), .Z(n17021) );
  XNOR U17219 ( .A(n16661), .B(n16660), .Z(n17022) );
  NANDN U17220 ( .A(n17021), .B(n17022), .Z(n16662) );
  NAND U17221 ( .A(n16663), .B(n16662), .Z(n16664) );
  OR U17222 ( .A(n16665), .B(n16664), .Z(n16669) );
  XNOR U17223 ( .A(n16665), .B(n16664), .Z(n17025) );
  XOR U17224 ( .A(n16667), .B(n16666), .Z(n17026) );
  NANDN U17225 ( .A(n17025), .B(n17026), .Z(n16668) );
  NAND U17226 ( .A(n16669), .B(n16668), .Z(n16672) );
  XOR U17227 ( .A(n16671), .B(n16670), .Z(n16673) );
  NANDN U17228 ( .A(n16672), .B(n16673), .Z(n16675) );
  NAND U17229 ( .A(a[8]), .B(b[13]), .Z(n17033) );
  XNOR U17230 ( .A(n16673), .B(n16672), .Z(n17034) );
  NANDN U17231 ( .A(n17033), .B(n17034), .Z(n16674) );
  NAND U17232 ( .A(n16675), .B(n16674), .Z(n16676) );
  OR U17233 ( .A(n16677), .B(n16676), .Z(n16681) );
  XNOR U17234 ( .A(n16677), .B(n16676), .Z(n17037) );
  XOR U17235 ( .A(n16679), .B(n16678), .Z(n17038) );
  NANDN U17236 ( .A(n17037), .B(n17038), .Z(n16680) );
  NAND U17237 ( .A(n16681), .B(n16680), .Z(n16683) );
  NAND U17238 ( .A(b[13]), .B(a[10]), .Z(n16682) );
  OR U17239 ( .A(n16683), .B(n16682), .Z(n16687) );
  XOR U17240 ( .A(n16683), .B(n16682), .Z(n17043) );
  XNOR U17241 ( .A(n16685), .B(n16684), .Z(n17044) );
  NAND U17242 ( .A(n17043), .B(n17044), .Z(n16686) );
  NAND U17243 ( .A(n16687), .B(n16686), .Z(n16690) );
  NANDN U17244 ( .A(n16691), .B(n16690), .Z(n16693) );
  XOR U17245 ( .A(n16689), .B(n16688), .Z(n17052) );
  NANDN U17246 ( .A(n17052), .B(n17051), .Z(n16692) );
  NAND U17247 ( .A(n16693), .B(n16692), .Z(n16697) );
  NAND U17248 ( .A(n16697), .B(n16696), .Z(n16699) );
  XNOR U17249 ( .A(n16697), .B(n16696), .Z(n17058) );
  NAND U17250 ( .A(a[12]), .B(b[13]), .Z(n17057) );
  OR U17251 ( .A(n17058), .B(n17057), .Z(n16698) );
  NAND U17252 ( .A(n16699), .B(n16698), .Z(n16702) );
  OR U17253 ( .A(n16703), .B(n16702), .Z(n16705) );
  XOR U17254 ( .A(n16701), .B(n16700), .Z(n17062) );
  XOR U17255 ( .A(n16703), .B(n16702), .Z(n17061) );
  NANDN U17256 ( .A(n17062), .B(n17061), .Z(n16704) );
  NAND U17257 ( .A(n16705), .B(n16704), .Z(n16706) );
  OR U17258 ( .A(n16707), .B(n16706), .Z(n16709) );
  NAND U17259 ( .A(b[13]), .B(a[14]), .Z(n17067) );
  XOR U17260 ( .A(n16707), .B(n16706), .Z(n17068) );
  NANDN U17261 ( .A(n17067), .B(n17068), .Z(n16708) );
  NAND U17262 ( .A(n16709), .B(n16708), .Z(n16712) );
  OR U17263 ( .A(n16713), .B(n16712), .Z(n16715) );
  XOR U17264 ( .A(n16713), .B(n16712), .Z(n16985) );
  NANDN U17265 ( .A(n16984), .B(n16985), .Z(n16714) );
  AND U17266 ( .A(n16715), .B(n16714), .Z(n16716) );
  OR U17267 ( .A(n16717), .B(n16716), .Z(n16719) );
  ANDN U17268 ( .B(b[13]), .A(n173), .Z(n17078) );
  XOR U17269 ( .A(n16717), .B(n16716), .Z(n17077) );
  NANDN U17270 ( .A(n17078), .B(n17077), .Z(n16718) );
  NAND U17271 ( .A(n16719), .B(n16718), .Z(n16722) );
  NANDN U17272 ( .A(n153), .B(a[17]), .Z(n16723) );
  NAND U17273 ( .A(n16722), .B(n16723), .Z(n16725) );
  XOR U17274 ( .A(n16721), .B(n16720), .Z(n17083) );
  NAND U17275 ( .A(n17083), .B(n17084), .Z(n16724) );
  NAND U17276 ( .A(n16725), .B(n16724), .Z(n16728) );
  NANDN U17277 ( .A(n16728), .B(n16729), .Z(n16731) );
  NAND U17278 ( .A(b[13]), .B(a[18]), .Z(n17091) );
  XNOR U17279 ( .A(n16729), .B(n16728), .Z(n17092) );
  NANDN U17280 ( .A(n17091), .B(n17092), .Z(n16730) );
  NAND U17281 ( .A(n16731), .B(n16730), .Z(n16734) );
  OR U17282 ( .A(n16735), .B(n16734), .Z(n16737) );
  XOR U17283 ( .A(n16733), .B(n16732), .Z(n17095) );
  XOR U17284 ( .A(n16735), .B(n16734), .Z(n17096) );
  NAND U17285 ( .A(n17095), .B(n17096), .Z(n16736) );
  NAND U17286 ( .A(n16737), .B(n16736), .Z(n16740) );
  NANDN U17287 ( .A(n16740), .B(n16741), .Z(n16743) );
  NAND U17288 ( .A(b[13]), .B(a[20]), .Z(n17103) );
  XNOR U17289 ( .A(n16741), .B(n16740), .Z(n17104) );
  NANDN U17290 ( .A(n17103), .B(n17104), .Z(n16742) );
  NAND U17291 ( .A(n16743), .B(n16742), .Z(n16746) );
  OR U17292 ( .A(n16747), .B(n16746), .Z(n16749) );
  XOR U17293 ( .A(n16745), .B(n16744), .Z(n17107) );
  XOR U17294 ( .A(n16747), .B(n16746), .Z(n17108) );
  NAND U17295 ( .A(n17107), .B(n17108), .Z(n16748) );
  NAND U17296 ( .A(n16749), .B(n16748), .Z(n16750) );
  OR U17297 ( .A(n16751), .B(n16750), .Z(n16753) );
  NAND U17298 ( .A(b[13]), .B(a[22]), .Z(n17115) );
  XOR U17299 ( .A(n16751), .B(n16750), .Z(n17116) );
  NANDN U17300 ( .A(n17115), .B(n17116), .Z(n16752) );
  AND U17301 ( .A(n16753), .B(n16752), .Z(n16754) );
  NANDN U17302 ( .A(n16755), .B(n16754), .Z(n16759) );
  XOR U17303 ( .A(n16757), .B(n16756), .Z(n17119) );
  NANDN U17304 ( .A(n17120), .B(n17119), .Z(n16758) );
  NAND U17305 ( .A(n16759), .B(n16758), .Z(n16761) );
  NANDN U17306 ( .A(n16760), .B(n16761), .Z(n16763) );
  ANDN U17307 ( .B(b[13]), .A(n178), .Z(n17126) );
  XNOR U17308 ( .A(n16761), .B(n16760), .Z(n17125) );
  NANDN U17309 ( .A(n17126), .B(n17125), .Z(n16762) );
  NAND U17310 ( .A(n16763), .B(n16762), .Z(n16766) );
  NANDN U17311 ( .A(n153), .B(a[25]), .Z(n16767) );
  NAND U17312 ( .A(n16766), .B(n16767), .Z(n16769) );
  XOR U17313 ( .A(n16765), .B(n16764), .Z(n17131) );
  NAND U17314 ( .A(n17131), .B(n17132), .Z(n16768) );
  NAND U17315 ( .A(n16769), .B(n16768), .Z(n16772) );
  NANDN U17316 ( .A(n16772), .B(n16773), .Z(n16775) );
  NAND U17317 ( .A(b[13]), .B(a[26]), .Z(n17139) );
  XNOR U17318 ( .A(n16773), .B(n16772), .Z(n17140) );
  NANDN U17319 ( .A(n17139), .B(n17140), .Z(n16774) );
  NAND U17320 ( .A(n16775), .B(n16774), .Z(n16778) );
  OR U17321 ( .A(n16779), .B(n16778), .Z(n16781) );
  XOR U17322 ( .A(n16777), .B(n16776), .Z(n17143) );
  XOR U17323 ( .A(n16779), .B(n16778), .Z(n17144) );
  NAND U17324 ( .A(n17143), .B(n17144), .Z(n16780) );
  NAND U17325 ( .A(n16781), .B(n16780), .Z(n16784) );
  NANDN U17326 ( .A(n16784), .B(n16785), .Z(n16787) );
  NAND U17327 ( .A(b[13]), .B(a[28]), .Z(n17151) );
  XNOR U17328 ( .A(n16785), .B(n16784), .Z(n17152) );
  NANDN U17329 ( .A(n17151), .B(n17152), .Z(n16786) );
  NAND U17330 ( .A(n16787), .B(n16786), .Z(n16790) );
  OR U17331 ( .A(n16791), .B(n16790), .Z(n16793) );
  XOR U17332 ( .A(n16789), .B(n16788), .Z(n17155) );
  XOR U17333 ( .A(n16791), .B(n16790), .Z(n17156) );
  NAND U17334 ( .A(n17155), .B(n17156), .Z(n16792) );
  NAND U17335 ( .A(n16793), .B(n16792), .Z(n16796) );
  NANDN U17336 ( .A(n16796), .B(n16797), .Z(n16799) );
  NAND U17337 ( .A(b[13]), .B(a[30]), .Z(n17163) );
  XNOR U17338 ( .A(n16797), .B(n16796), .Z(n17164) );
  NANDN U17339 ( .A(n17163), .B(n17164), .Z(n16798) );
  NAND U17340 ( .A(n16799), .B(n16798), .Z(n16802) );
  OR U17341 ( .A(n16803), .B(n16802), .Z(n16805) );
  XOR U17342 ( .A(n16801), .B(n16800), .Z(n17167) );
  XOR U17343 ( .A(n16803), .B(n16802), .Z(n17168) );
  NAND U17344 ( .A(n17167), .B(n17168), .Z(n16804) );
  NAND U17345 ( .A(n16805), .B(n16804), .Z(n16808) );
  NANDN U17346 ( .A(n16808), .B(n16809), .Z(n16811) );
  NAND U17347 ( .A(b[13]), .B(a[32]), .Z(n17175) );
  XNOR U17348 ( .A(n16809), .B(n16808), .Z(n17176) );
  NANDN U17349 ( .A(n17175), .B(n17176), .Z(n16810) );
  NAND U17350 ( .A(n16811), .B(n16810), .Z(n16814) );
  OR U17351 ( .A(n16815), .B(n16814), .Z(n16817) );
  XOR U17352 ( .A(n16813), .B(n16812), .Z(n17179) );
  XOR U17353 ( .A(n16815), .B(n16814), .Z(n17180) );
  NAND U17354 ( .A(n17179), .B(n17180), .Z(n16816) );
  NAND U17355 ( .A(n16817), .B(n16816), .Z(n16820) );
  NANDN U17356 ( .A(n16820), .B(n16821), .Z(n16823) );
  NAND U17357 ( .A(b[13]), .B(a[34]), .Z(n17187) );
  XNOR U17358 ( .A(n16821), .B(n16820), .Z(n17188) );
  NANDN U17359 ( .A(n17187), .B(n17188), .Z(n16822) );
  NAND U17360 ( .A(n16823), .B(n16822), .Z(n16826) );
  OR U17361 ( .A(n16827), .B(n16826), .Z(n16829) );
  XOR U17362 ( .A(n16825), .B(n16824), .Z(n17191) );
  XOR U17363 ( .A(n16827), .B(n16826), .Z(n17192) );
  NAND U17364 ( .A(n17191), .B(n17192), .Z(n16828) );
  NAND U17365 ( .A(n16829), .B(n16828), .Z(n16832) );
  NANDN U17366 ( .A(n16832), .B(n16833), .Z(n16835) );
  NAND U17367 ( .A(b[13]), .B(a[36]), .Z(n17199) );
  XNOR U17368 ( .A(n16833), .B(n16832), .Z(n17200) );
  NANDN U17369 ( .A(n17199), .B(n17200), .Z(n16834) );
  NAND U17370 ( .A(n16835), .B(n16834), .Z(n16838) );
  OR U17371 ( .A(n16839), .B(n16838), .Z(n16841) );
  XOR U17372 ( .A(n16837), .B(n16836), .Z(n17203) );
  XOR U17373 ( .A(n16839), .B(n16838), .Z(n17204) );
  NAND U17374 ( .A(n17203), .B(n17204), .Z(n16840) );
  NAND U17375 ( .A(n16841), .B(n16840), .Z(n16844) );
  NANDN U17376 ( .A(n16844), .B(n16845), .Z(n16847) );
  NAND U17377 ( .A(b[13]), .B(a[38]), .Z(n17211) );
  XNOR U17378 ( .A(n16845), .B(n16844), .Z(n17212) );
  NANDN U17379 ( .A(n17211), .B(n17212), .Z(n16846) );
  NAND U17380 ( .A(n16847), .B(n16846), .Z(n16850) );
  OR U17381 ( .A(n16851), .B(n16850), .Z(n16853) );
  XOR U17382 ( .A(n16849), .B(n16848), .Z(n17215) );
  XOR U17383 ( .A(n16851), .B(n16850), .Z(n17216) );
  NAND U17384 ( .A(n17215), .B(n17216), .Z(n16852) );
  NAND U17385 ( .A(n16853), .B(n16852), .Z(n16856) );
  NANDN U17386 ( .A(n16856), .B(n16857), .Z(n16859) );
  NAND U17387 ( .A(b[13]), .B(a[40]), .Z(n17223) );
  XNOR U17388 ( .A(n16857), .B(n16856), .Z(n17224) );
  NANDN U17389 ( .A(n17223), .B(n17224), .Z(n16858) );
  NAND U17390 ( .A(n16859), .B(n16858), .Z(n16862) );
  OR U17391 ( .A(n16863), .B(n16862), .Z(n16865) );
  XOR U17392 ( .A(n16861), .B(n16860), .Z(n17227) );
  XOR U17393 ( .A(n16863), .B(n16862), .Z(n17228) );
  NAND U17394 ( .A(n17227), .B(n17228), .Z(n16864) );
  NAND U17395 ( .A(n16865), .B(n16864), .Z(n16868) );
  NANDN U17396 ( .A(n16868), .B(n16869), .Z(n16871) );
  NAND U17397 ( .A(b[13]), .B(a[42]), .Z(n17235) );
  XNOR U17398 ( .A(n16869), .B(n16868), .Z(n17236) );
  NANDN U17399 ( .A(n17235), .B(n17236), .Z(n16870) );
  NAND U17400 ( .A(n16871), .B(n16870), .Z(n16874) );
  OR U17401 ( .A(n16875), .B(n16874), .Z(n16877) );
  XOR U17402 ( .A(n16873), .B(n16872), .Z(n17239) );
  XOR U17403 ( .A(n16875), .B(n16874), .Z(n17240) );
  NAND U17404 ( .A(n17239), .B(n17240), .Z(n16876) );
  NAND U17405 ( .A(n16877), .B(n16876), .Z(n16880) );
  NANDN U17406 ( .A(n16880), .B(n16881), .Z(n16883) );
  NAND U17407 ( .A(b[13]), .B(a[44]), .Z(n17247) );
  XNOR U17408 ( .A(n16881), .B(n16880), .Z(n17248) );
  NANDN U17409 ( .A(n17247), .B(n17248), .Z(n16882) );
  NAND U17410 ( .A(n16883), .B(n16882), .Z(n16886) );
  OR U17411 ( .A(n16887), .B(n16886), .Z(n16889) );
  XOR U17412 ( .A(n16885), .B(n16884), .Z(n17251) );
  XOR U17413 ( .A(n16887), .B(n16886), .Z(n17252) );
  NAND U17414 ( .A(n17251), .B(n17252), .Z(n16888) );
  NAND U17415 ( .A(n16889), .B(n16888), .Z(n16892) );
  NANDN U17416 ( .A(n16892), .B(n16893), .Z(n16895) );
  NAND U17417 ( .A(b[13]), .B(a[46]), .Z(n17259) );
  XNOR U17418 ( .A(n16893), .B(n16892), .Z(n17260) );
  NANDN U17419 ( .A(n17259), .B(n17260), .Z(n16894) );
  NAND U17420 ( .A(n16895), .B(n16894), .Z(n16898) );
  OR U17421 ( .A(n16899), .B(n16898), .Z(n16901) );
  XOR U17422 ( .A(n16897), .B(n16896), .Z(n17263) );
  XOR U17423 ( .A(n16899), .B(n16898), .Z(n17264) );
  NAND U17424 ( .A(n17263), .B(n17264), .Z(n16900) );
  NAND U17425 ( .A(n16901), .B(n16900), .Z(n16904) );
  NANDN U17426 ( .A(n16904), .B(n16905), .Z(n16907) );
  NAND U17427 ( .A(b[13]), .B(a[48]), .Z(n17271) );
  XNOR U17428 ( .A(n16905), .B(n16904), .Z(n17272) );
  NANDN U17429 ( .A(n17271), .B(n17272), .Z(n16906) );
  NAND U17430 ( .A(n16907), .B(n16906), .Z(n16908) );
  ANDN U17431 ( .B(b[13]), .A(n197), .Z(n16909) );
  OR U17432 ( .A(n16908), .B(n16909), .Z(n16913) );
  XNOR U17433 ( .A(n16909), .B(n16908), .Z(n17275) );
  XNOR U17434 ( .A(n16911), .B(n16910), .Z(n17276) );
  OR U17435 ( .A(n17275), .B(n17276), .Z(n16912) );
  NAND U17436 ( .A(n16913), .B(n16912), .Z(n16916) );
  XOR U17437 ( .A(n16915), .B(n16914), .Z(n16917) );
  OR U17438 ( .A(n16916), .B(n16917), .Z(n16919) );
  XNOR U17439 ( .A(n16917), .B(n16916), .Z(n17284) );
  AND U17440 ( .A(a[50]), .B(b[13]), .Z(n17283) );
  NANDN U17441 ( .A(n17284), .B(n17283), .Z(n16918) );
  NAND U17442 ( .A(n16919), .B(n16918), .Z(n16920) );
  ANDN U17443 ( .B(b[13]), .A(n199), .Z(n16921) );
  OR U17444 ( .A(n16920), .B(n16921), .Z(n16925) );
  XNOR U17445 ( .A(n16921), .B(n16920), .Z(n17289) );
  XNOR U17446 ( .A(n16923), .B(n16922), .Z(n17290) );
  OR U17447 ( .A(n17289), .B(n17290), .Z(n16924) );
  NAND U17448 ( .A(n16925), .B(n16924), .Z(n16927) );
  NAND U17449 ( .A(b[13]), .B(a[52]), .Z(n16926) );
  OR U17450 ( .A(n16927), .B(n16926), .Z(n16931) );
  XOR U17451 ( .A(n16927), .B(n16926), .Z(n17295) );
  XOR U17452 ( .A(n16929), .B(n16928), .Z(n17296) );
  NAND U17453 ( .A(n17295), .B(n17296), .Z(n16930) );
  NAND U17454 ( .A(n16931), .B(n16930), .Z(n16933) );
  NAND U17455 ( .A(n16932), .B(n16933), .Z(n16935) );
  NAND U17456 ( .A(a[53]), .B(b[13]), .Z(n17301) );
  NANDN U17457 ( .A(n17301), .B(n17302), .Z(n16934) );
  NAND U17458 ( .A(n16935), .B(n16934), .Z(n16937) );
  NANDN U17459 ( .A(n16936), .B(n16937), .Z(n16941) );
  XOR U17460 ( .A(n16937), .B(n16936), .Z(n17308) );
  XOR U17461 ( .A(n16939), .B(n16938), .Z(n17307) );
  NANDN U17462 ( .A(n17308), .B(n17307), .Z(n16940) );
  NAND U17463 ( .A(n16941), .B(n16940), .Z(n16943) );
  NAND U17464 ( .A(n16942), .B(n16943), .Z(n16945) );
  NAND U17465 ( .A(a[55]), .B(b[13]), .Z(n17313) );
  NANDN U17466 ( .A(n17313), .B(n17314), .Z(n16944) );
  NAND U17467 ( .A(n16945), .B(n16944), .Z(n16947) );
  NANDN U17468 ( .A(n16946), .B(n16947), .Z(n16951) );
  XOR U17469 ( .A(n16947), .B(n16946), .Z(n17320) );
  XOR U17470 ( .A(n16949), .B(n16948), .Z(n17319) );
  NANDN U17471 ( .A(n17320), .B(n17319), .Z(n16950) );
  NAND U17472 ( .A(n16951), .B(n16950), .Z(n16953) );
  NAND U17473 ( .A(n16952), .B(n16953), .Z(n16955) );
  NAND U17474 ( .A(a[57]), .B(b[13]), .Z(n17325) );
  NANDN U17475 ( .A(n17325), .B(n17326), .Z(n16954) );
  NAND U17476 ( .A(n16955), .B(n16954), .Z(n16957) );
  NANDN U17477 ( .A(n16956), .B(n16957), .Z(n16961) );
  XOR U17478 ( .A(n16957), .B(n16956), .Z(n17330) );
  XOR U17479 ( .A(n16959), .B(n16958), .Z(n17329) );
  NANDN U17480 ( .A(n17330), .B(n17329), .Z(n16960) );
  NAND U17481 ( .A(n16961), .B(n16960), .Z(n16963) );
  NAND U17482 ( .A(n16962), .B(n16963), .Z(n16965) );
  NAND U17483 ( .A(a[59]), .B(b[13]), .Z(n17337) );
  NANDN U17484 ( .A(n17337), .B(n17338), .Z(n16964) );
  NAND U17485 ( .A(n16965), .B(n16964), .Z(n16967) );
  NANDN U17486 ( .A(n16966), .B(n16967), .Z(n16971) );
  XOR U17487 ( .A(n16967), .B(n16966), .Z(n17342) );
  XOR U17488 ( .A(n16969), .B(n16968), .Z(n17341) );
  NANDN U17489 ( .A(n17342), .B(n17341), .Z(n16970) );
  NAND U17490 ( .A(n16971), .B(n16970), .Z(n16975) );
  XOR U17491 ( .A(n16973), .B(n16972), .Z(n16974) );
  NAND U17492 ( .A(n16975), .B(n16974), .Z(n16977) );
  NAND U17493 ( .A(a[61]), .B(b[13]), .Z(n17347) );
  XOR U17494 ( .A(n16975), .B(n16974), .Z(n17348) );
  NANDN U17495 ( .A(n17347), .B(n17348), .Z(n16976) );
  NAND U17496 ( .A(n16977), .B(n16976), .Z(n16979) );
  XOR U17497 ( .A(n16979), .B(n16978), .Z(n17353) );
  XOR U17498 ( .A(n16981), .B(n16980), .Z(n17354) );
  XOR U17499 ( .A(n16983), .B(n16982), .Z(n17361) );
  AND U17500 ( .A(a[63]), .B(b[13]), .Z(n17363) );
  XOR U17501 ( .A(n17364), .B(n17363), .Z(n18500) );
  ANDN U17502 ( .B(b[12]), .A(n209), .Z(n17344) );
  ANDN U17503 ( .B(b[12]), .A(n207), .Z(n17332) );
  ANDN U17504 ( .B(b[12]), .A(n205), .Z(n17318) );
  ANDN U17505 ( .B(b[12]), .A(n203), .Z(n17306) );
  NAND U17506 ( .A(a[54]), .B(b[12]), .Z(n17299) );
  NAND U17507 ( .A(a[53]), .B(b[12]), .Z(n17293) );
  ANDN U17508 ( .B(b[12]), .A(n197), .Z(n17270) );
  ANDN U17509 ( .B(b[12]), .A(n195), .Z(n17258) );
  ANDN U17510 ( .B(b[12]), .A(n193), .Z(n17246) );
  ANDN U17511 ( .B(b[12]), .A(n191), .Z(n17234) );
  ANDN U17512 ( .B(b[12]), .A(n189), .Z(n17222) );
  ANDN U17513 ( .B(b[12]), .A(n187), .Z(n17210) );
  ANDN U17514 ( .B(b[12]), .A(n21772), .Z(n17198) );
  ANDN U17515 ( .B(b[12]), .A(n184), .Z(n17186) );
  ANDN U17516 ( .B(b[12]), .A(n21751), .Z(n17174) );
  ANDN U17517 ( .B(b[12]), .A(n21740), .Z(n17162) );
  ANDN U17518 ( .B(b[12]), .A(n21727), .Z(n17150) );
  ANDN U17519 ( .B(b[12]), .A(n21716), .Z(n17138) );
  ANDN U17520 ( .B(b[12]), .A(n21703), .Z(n17128) );
  ANDN U17521 ( .B(b[12]), .A(n21692), .Z(n17114) );
  ANDN U17522 ( .B(b[12]), .A(n21681), .Z(n17102) );
  ANDN U17523 ( .B(b[12]), .A(n21670), .Z(n17090) );
  XOR U17524 ( .A(n16985), .B(n16984), .Z(n17073) );
  ANDN U17525 ( .B(b[12]), .A(n172), .Z(n17070) );
  ANDN U17526 ( .B(b[12]), .A(n170), .Z(n17056) );
  ANDN U17527 ( .B(b[12]), .A(n21164), .Z(n17046) );
  ANDN U17528 ( .B(b[12]), .A(n21615), .Z(n17032) );
  ANDN U17529 ( .B(b[12]), .A(n166), .Z(n17020) );
  NAND U17530 ( .A(a[6]), .B(b[12]), .Z(n17015) );
  XOR U17531 ( .A(n16987), .B(n16986), .Z(n17016) );
  NANDN U17532 ( .A(n17015), .B(n17016), .Z(n17018) );
  ANDN U17533 ( .B(b[12]), .A(n164), .Z(n17010) );
  ANDN U17534 ( .B(b[12]), .A(n21580), .Z(n16997) );
  NAND U17535 ( .A(b[13]), .B(a[1]), .Z(n16990) );
  AND U17536 ( .A(b[12]), .B(a[0]), .Z(n17754) );
  NANDN U17537 ( .A(n16990), .B(n17754), .Z(n16989) );
  NAND U17538 ( .A(b[12]), .B(a[2]), .Z(n16988) );
  AND U17539 ( .A(n16989), .B(n16988), .Z(n16996) );
  NANDN U17540 ( .A(n16990), .B(a[0]), .Z(n16991) );
  XNOR U17541 ( .A(a[2]), .B(n16991), .Z(n16992) );
  NAND U17542 ( .A(b[12]), .B(n16992), .Z(n17385) );
  AND U17543 ( .A(a[1]), .B(b[13]), .Z(n16993) );
  XNOR U17544 ( .A(n16994), .B(n16993), .Z(n17384) );
  NANDN U17545 ( .A(n17385), .B(n17384), .Z(n16995) );
  NANDN U17546 ( .A(n16996), .B(n16995), .Z(n16998) );
  NANDN U17547 ( .A(n16997), .B(n16998), .Z(n17002) );
  XOR U17548 ( .A(n16998), .B(n16997), .Z(n17389) );
  NANDN U17549 ( .A(n17389), .B(n17388), .Z(n17001) );
  NAND U17550 ( .A(n17002), .B(n17001), .Z(n17006) );
  XOR U17551 ( .A(n17004), .B(n17003), .Z(n17005) );
  NANDN U17552 ( .A(n17006), .B(n17005), .Z(n17008) );
  NAND U17553 ( .A(a[4]), .B(b[12]), .Z(n17396) );
  NANDN U17554 ( .A(n17396), .B(n17397), .Z(n17007) );
  NAND U17555 ( .A(n17008), .B(n17007), .Z(n17009) );
  OR U17556 ( .A(n17010), .B(n17009), .Z(n17014) );
  XNOR U17557 ( .A(n17010), .B(n17009), .Z(n17400) );
  XOR U17558 ( .A(n17012), .B(n17011), .Z(n17401) );
  NANDN U17559 ( .A(n17400), .B(n17401), .Z(n17013) );
  NAND U17560 ( .A(n17014), .B(n17013), .Z(n17408) );
  XNOR U17561 ( .A(n17016), .B(n17015), .Z(n17409) );
  NANDN U17562 ( .A(n17408), .B(n17409), .Z(n17017) );
  NAND U17563 ( .A(n17018), .B(n17017), .Z(n17019) );
  OR U17564 ( .A(n17020), .B(n17019), .Z(n17024) );
  XNOR U17565 ( .A(n17020), .B(n17019), .Z(n17412) );
  XOR U17566 ( .A(n17022), .B(n17021), .Z(n17413) );
  NANDN U17567 ( .A(n17412), .B(n17413), .Z(n17023) );
  NAND U17568 ( .A(n17024), .B(n17023), .Z(n17027) );
  XOR U17569 ( .A(n17026), .B(n17025), .Z(n17028) );
  NANDN U17570 ( .A(n17027), .B(n17028), .Z(n17030) );
  NAND U17571 ( .A(a[8]), .B(b[12]), .Z(n17420) );
  XNOR U17572 ( .A(n17028), .B(n17027), .Z(n17421) );
  NANDN U17573 ( .A(n17420), .B(n17421), .Z(n17029) );
  NAND U17574 ( .A(n17030), .B(n17029), .Z(n17031) );
  OR U17575 ( .A(n17032), .B(n17031), .Z(n17036) );
  XNOR U17576 ( .A(n17032), .B(n17031), .Z(n17424) );
  XOR U17577 ( .A(n17034), .B(n17033), .Z(n17425) );
  NANDN U17578 ( .A(n17424), .B(n17425), .Z(n17035) );
  NAND U17579 ( .A(n17036), .B(n17035), .Z(n17039) );
  XOR U17580 ( .A(n17038), .B(n17037), .Z(n17040) );
  NANDN U17581 ( .A(n17039), .B(n17040), .Z(n17042) );
  NAND U17582 ( .A(a[10]), .B(b[12]), .Z(n17432) );
  XNOR U17583 ( .A(n17040), .B(n17039), .Z(n17433) );
  NANDN U17584 ( .A(n17432), .B(n17433), .Z(n17041) );
  NAND U17585 ( .A(n17042), .B(n17041), .Z(n17045) );
  OR U17586 ( .A(n17046), .B(n17045), .Z(n17048) );
  XOR U17587 ( .A(n17046), .B(n17045), .Z(n17436) );
  NANDN U17588 ( .A(n17437), .B(n17436), .Z(n17047) );
  NAND U17589 ( .A(n17048), .B(n17047), .Z(n17050) );
  NAND U17590 ( .A(b[12]), .B(a[12]), .Z(n17049) );
  OR U17591 ( .A(n17050), .B(n17049), .Z(n17054) );
  XOR U17592 ( .A(n17050), .B(n17049), .Z(n17442) );
  XNOR U17593 ( .A(n17052), .B(n17051), .Z(n17443) );
  NAND U17594 ( .A(n17442), .B(n17443), .Z(n17053) );
  NAND U17595 ( .A(n17054), .B(n17053), .Z(n17055) );
  OR U17596 ( .A(n17056), .B(n17055), .Z(n17060) );
  XNOR U17597 ( .A(n17056), .B(n17055), .Z(n17448) );
  XNOR U17598 ( .A(n17058), .B(n17057), .Z(n17449) );
  NANDN U17599 ( .A(n17448), .B(n17449), .Z(n17059) );
  NAND U17600 ( .A(n17060), .B(n17059), .Z(n17063) );
  XNOR U17601 ( .A(n17062), .B(n17061), .Z(n17064) );
  OR U17602 ( .A(n17063), .B(n17064), .Z(n17066) );
  NAND U17603 ( .A(b[12]), .B(a[14]), .Z(n17456) );
  XOR U17604 ( .A(n17064), .B(n17063), .Z(n17457) );
  NANDN U17605 ( .A(n17456), .B(n17457), .Z(n17065) );
  NAND U17606 ( .A(n17066), .B(n17065), .Z(n17069) );
  OR U17607 ( .A(n17070), .B(n17069), .Z(n17072) );
  XOR U17608 ( .A(n17068), .B(n17067), .Z(n17372) );
  XOR U17609 ( .A(n17070), .B(n17069), .Z(n17371) );
  NAND U17610 ( .A(n17372), .B(n17371), .Z(n17071) );
  NAND U17611 ( .A(n17072), .B(n17071), .Z(n17074) );
  NANDN U17612 ( .A(n17073), .B(n17074), .Z(n17076) );
  ANDN U17613 ( .B(b[12]), .A(n173), .Z(n17465) );
  XOR U17614 ( .A(n17074), .B(n17073), .Z(n17464) );
  OR U17615 ( .A(n17465), .B(n17464), .Z(n17075) );
  NAND U17616 ( .A(n17076), .B(n17075), .Z(n17079) );
  NAND U17617 ( .A(n17079), .B(n17080), .Z(n17082) );
  XOR U17618 ( .A(n17078), .B(n17077), .Z(n17470) );
  NANDN U17619 ( .A(n17470), .B(n17471), .Z(n17081) );
  NAND U17620 ( .A(n17082), .B(n17081), .Z(n17085) );
  NANDN U17621 ( .A(n17085), .B(n17086), .Z(n17088) );
  NAND U17622 ( .A(a[18]), .B(b[12]), .Z(n17478) );
  XNOR U17623 ( .A(n17086), .B(n17085), .Z(n17479) );
  NANDN U17624 ( .A(n17478), .B(n17479), .Z(n17087) );
  AND U17625 ( .A(n17088), .B(n17087), .Z(n17089) );
  NANDN U17626 ( .A(n17090), .B(n17089), .Z(n17094) );
  XOR U17627 ( .A(n17092), .B(n17091), .Z(n17482) );
  NANDN U17628 ( .A(n17483), .B(n17482), .Z(n17093) );
  NAND U17629 ( .A(n17094), .B(n17093), .Z(n17097) );
  NANDN U17630 ( .A(n17097), .B(n17098), .Z(n17100) );
  NAND U17631 ( .A(a[20]), .B(b[12]), .Z(n17490) );
  XNOR U17632 ( .A(n17098), .B(n17097), .Z(n17491) );
  NANDN U17633 ( .A(n17490), .B(n17491), .Z(n17099) );
  AND U17634 ( .A(n17100), .B(n17099), .Z(n17101) );
  NANDN U17635 ( .A(n17102), .B(n17101), .Z(n17106) );
  XOR U17636 ( .A(n17104), .B(n17103), .Z(n17494) );
  NANDN U17637 ( .A(n17495), .B(n17494), .Z(n17105) );
  NAND U17638 ( .A(n17106), .B(n17105), .Z(n17109) );
  NANDN U17639 ( .A(n17109), .B(n17110), .Z(n17112) );
  NAND U17640 ( .A(a[22]), .B(b[12]), .Z(n17502) );
  XNOR U17641 ( .A(n17110), .B(n17109), .Z(n17503) );
  NANDN U17642 ( .A(n17502), .B(n17503), .Z(n17111) );
  AND U17643 ( .A(n17112), .B(n17111), .Z(n17113) );
  NANDN U17644 ( .A(n17114), .B(n17113), .Z(n17118) );
  XOR U17645 ( .A(n17116), .B(n17115), .Z(n17506) );
  NANDN U17646 ( .A(n17507), .B(n17506), .Z(n17117) );
  NAND U17647 ( .A(n17118), .B(n17117), .Z(n17121) );
  NANDN U17648 ( .A(n17121), .B(n17122), .Z(n17124) );
  NAND U17649 ( .A(a[24]), .B(b[12]), .Z(n17514) );
  XNOR U17650 ( .A(n17122), .B(n17121), .Z(n17515) );
  NANDN U17651 ( .A(n17514), .B(n17515), .Z(n17123) );
  NAND U17652 ( .A(n17124), .B(n17123), .Z(n17127) );
  OR U17653 ( .A(n17128), .B(n17127), .Z(n17130) );
  XOR U17654 ( .A(n17126), .B(n17125), .Z(n17519) );
  XOR U17655 ( .A(n17128), .B(n17127), .Z(n17518) );
  NANDN U17656 ( .A(n17519), .B(n17518), .Z(n17129) );
  NAND U17657 ( .A(n17130), .B(n17129), .Z(n17133) );
  NANDN U17658 ( .A(n17133), .B(n17134), .Z(n17136) );
  NAND U17659 ( .A(a[26]), .B(b[12]), .Z(n17526) );
  XNOR U17660 ( .A(n17134), .B(n17133), .Z(n17527) );
  NANDN U17661 ( .A(n17526), .B(n17527), .Z(n17135) );
  AND U17662 ( .A(n17136), .B(n17135), .Z(n17137) );
  NANDN U17663 ( .A(n17138), .B(n17137), .Z(n17142) );
  XOR U17664 ( .A(n17140), .B(n17139), .Z(n17530) );
  NANDN U17665 ( .A(n17531), .B(n17530), .Z(n17141) );
  NAND U17666 ( .A(n17142), .B(n17141), .Z(n17145) );
  NANDN U17667 ( .A(n17145), .B(n17146), .Z(n17148) );
  NAND U17668 ( .A(a[28]), .B(b[12]), .Z(n17538) );
  XNOR U17669 ( .A(n17146), .B(n17145), .Z(n17539) );
  NANDN U17670 ( .A(n17538), .B(n17539), .Z(n17147) );
  AND U17671 ( .A(n17148), .B(n17147), .Z(n17149) );
  NANDN U17672 ( .A(n17150), .B(n17149), .Z(n17154) );
  XOR U17673 ( .A(n17152), .B(n17151), .Z(n17542) );
  NANDN U17674 ( .A(n17543), .B(n17542), .Z(n17153) );
  NAND U17675 ( .A(n17154), .B(n17153), .Z(n17157) );
  NANDN U17676 ( .A(n17157), .B(n17158), .Z(n17160) );
  NAND U17677 ( .A(a[30]), .B(b[12]), .Z(n17550) );
  XNOR U17678 ( .A(n17158), .B(n17157), .Z(n17551) );
  NANDN U17679 ( .A(n17550), .B(n17551), .Z(n17159) );
  AND U17680 ( .A(n17160), .B(n17159), .Z(n17161) );
  NANDN U17681 ( .A(n17162), .B(n17161), .Z(n17166) );
  XOR U17682 ( .A(n17164), .B(n17163), .Z(n17554) );
  NANDN U17683 ( .A(n17555), .B(n17554), .Z(n17165) );
  NAND U17684 ( .A(n17166), .B(n17165), .Z(n17169) );
  NANDN U17685 ( .A(n17169), .B(n17170), .Z(n17172) );
  NAND U17686 ( .A(a[32]), .B(b[12]), .Z(n17562) );
  XNOR U17687 ( .A(n17170), .B(n17169), .Z(n17563) );
  NANDN U17688 ( .A(n17562), .B(n17563), .Z(n17171) );
  AND U17689 ( .A(n17172), .B(n17171), .Z(n17173) );
  NANDN U17690 ( .A(n17174), .B(n17173), .Z(n17178) );
  XOR U17691 ( .A(n17176), .B(n17175), .Z(n17566) );
  NANDN U17692 ( .A(n17567), .B(n17566), .Z(n17177) );
  NAND U17693 ( .A(n17178), .B(n17177), .Z(n17181) );
  NANDN U17694 ( .A(n17181), .B(n17182), .Z(n17184) );
  NAND U17695 ( .A(a[34]), .B(b[12]), .Z(n17574) );
  XNOR U17696 ( .A(n17182), .B(n17181), .Z(n17575) );
  NANDN U17697 ( .A(n17574), .B(n17575), .Z(n17183) );
  AND U17698 ( .A(n17184), .B(n17183), .Z(n17185) );
  NANDN U17699 ( .A(n17186), .B(n17185), .Z(n17190) );
  XOR U17700 ( .A(n17188), .B(n17187), .Z(n17578) );
  NANDN U17701 ( .A(n17579), .B(n17578), .Z(n17189) );
  NAND U17702 ( .A(n17190), .B(n17189), .Z(n17193) );
  NANDN U17703 ( .A(n17193), .B(n17194), .Z(n17196) );
  NAND U17704 ( .A(a[36]), .B(b[12]), .Z(n17586) );
  XNOR U17705 ( .A(n17194), .B(n17193), .Z(n17587) );
  NANDN U17706 ( .A(n17586), .B(n17587), .Z(n17195) );
  AND U17707 ( .A(n17196), .B(n17195), .Z(n17197) );
  NANDN U17708 ( .A(n17198), .B(n17197), .Z(n17202) );
  XOR U17709 ( .A(n17200), .B(n17199), .Z(n17590) );
  NANDN U17710 ( .A(n17591), .B(n17590), .Z(n17201) );
  NAND U17711 ( .A(n17202), .B(n17201), .Z(n17205) );
  NANDN U17712 ( .A(n17205), .B(n17206), .Z(n17208) );
  NAND U17713 ( .A(a[38]), .B(b[12]), .Z(n17598) );
  XNOR U17714 ( .A(n17206), .B(n17205), .Z(n17599) );
  NANDN U17715 ( .A(n17598), .B(n17599), .Z(n17207) );
  AND U17716 ( .A(n17208), .B(n17207), .Z(n17209) );
  NANDN U17717 ( .A(n17210), .B(n17209), .Z(n17214) );
  XOR U17718 ( .A(n17212), .B(n17211), .Z(n17602) );
  NANDN U17719 ( .A(n17603), .B(n17602), .Z(n17213) );
  NAND U17720 ( .A(n17214), .B(n17213), .Z(n17217) );
  NANDN U17721 ( .A(n17217), .B(n17218), .Z(n17220) );
  NAND U17722 ( .A(a[40]), .B(b[12]), .Z(n17610) );
  XNOR U17723 ( .A(n17218), .B(n17217), .Z(n17611) );
  NANDN U17724 ( .A(n17610), .B(n17611), .Z(n17219) );
  AND U17725 ( .A(n17220), .B(n17219), .Z(n17221) );
  NANDN U17726 ( .A(n17222), .B(n17221), .Z(n17226) );
  XOR U17727 ( .A(n17224), .B(n17223), .Z(n17614) );
  NANDN U17728 ( .A(n17615), .B(n17614), .Z(n17225) );
  NAND U17729 ( .A(n17226), .B(n17225), .Z(n17229) );
  NANDN U17730 ( .A(n17229), .B(n17230), .Z(n17232) );
  NAND U17731 ( .A(a[42]), .B(b[12]), .Z(n17622) );
  XNOR U17732 ( .A(n17230), .B(n17229), .Z(n17623) );
  NANDN U17733 ( .A(n17622), .B(n17623), .Z(n17231) );
  AND U17734 ( .A(n17232), .B(n17231), .Z(n17233) );
  NANDN U17735 ( .A(n17234), .B(n17233), .Z(n17238) );
  XOR U17736 ( .A(n17236), .B(n17235), .Z(n17626) );
  NANDN U17737 ( .A(n17627), .B(n17626), .Z(n17237) );
  NAND U17738 ( .A(n17238), .B(n17237), .Z(n17241) );
  NANDN U17739 ( .A(n17241), .B(n17242), .Z(n17244) );
  NAND U17740 ( .A(a[44]), .B(b[12]), .Z(n17634) );
  XNOR U17741 ( .A(n17242), .B(n17241), .Z(n17635) );
  NANDN U17742 ( .A(n17634), .B(n17635), .Z(n17243) );
  AND U17743 ( .A(n17244), .B(n17243), .Z(n17245) );
  NANDN U17744 ( .A(n17246), .B(n17245), .Z(n17250) );
  XOR U17745 ( .A(n17248), .B(n17247), .Z(n17638) );
  NANDN U17746 ( .A(n17639), .B(n17638), .Z(n17249) );
  NAND U17747 ( .A(n17250), .B(n17249), .Z(n17253) );
  NANDN U17748 ( .A(n17253), .B(n17254), .Z(n17256) );
  NAND U17749 ( .A(a[46]), .B(b[12]), .Z(n17646) );
  XNOR U17750 ( .A(n17254), .B(n17253), .Z(n17647) );
  NANDN U17751 ( .A(n17646), .B(n17647), .Z(n17255) );
  AND U17752 ( .A(n17256), .B(n17255), .Z(n17257) );
  NANDN U17753 ( .A(n17258), .B(n17257), .Z(n17262) );
  XOR U17754 ( .A(n17260), .B(n17259), .Z(n17650) );
  NANDN U17755 ( .A(n17651), .B(n17650), .Z(n17261) );
  NAND U17756 ( .A(n17262), .B(n17261), .Z(n17265) );
  NANDN U17757 ( .A(n17265), .B(n17266), .Z(n17268) );
  NAND U17758 ( .A(a[48]), .B(b[12]), .Z(n17658) );
  XNOR U17759 ( .A(n17266), .B(n17265), .Z(n17659) );
  NANDN U17760 ( .A(n17658), .B(n17659), .Z(n17267) );
  AND U17761 ( .A(n17268), .B(n17267), .Z(n17269) );
  NANDN U17762 ( .A(n17270), .B(n17269), .Z(n17274) );
  XOR U17763 ( .A(n17272), .B(n17271), .Z(n17662) );
  NANDN U17764 ( .A(n17663), .B(n17662), .Z(n17273) );
  NAND U17765 ( .A(n17274), .B(n17273), .Z(n17277) );
  XNOR U17766 ( .A(n17276), .B(n17275), .Z(n17278) );
  NANDN U17767 ( .A(n17277), .B(n17278), .Z(n17280) );
  XOR U17768 ( .A(n17278), .B(n17277), .Z(n17669) );
  NAND U17769 ( .A(a[50]), .B(b[12]), .Z(n17668) );
  OR U17770 ( .A(n17669), .B(n17668), .Z(n17279) );
  NAND U17771 ( .A(n17280), .B(n17279), .Z(n17281) );
  NAND U17772 ( .A(b[12]), .B(a[51]), .Z(n17282) );
  NANDN U17773 ( .A(n17281), .B(n17282), .Z(n17286) );
  XOR U17774 ( .A(n17282), .B(n17281), .Z(n17674) );
  XOR U17775 ( .A(n17284), .B(n17283), .Z(n17675) );
  NANDN U17776 ( .A(n17674), .B(n17675), .Z(n17285) );
  NAND U17777 ( .A(n17286), .B(n17285), .Z(n17288) );
  NAND U17778 ( .A(a[52]), .B(b[12]), .Z(n17287) );
  OR U17779 ( .A(n17288), .B(n17287), .Z(n17292) );
  XNOR U17780 ( .A(n17288), .B(n17287), .Z(n17680) );
  XNOR U17781 ( .A(n17290), .B(n17289), .Z(n17681) );
  NANDN U17782 ( .A(n17680), .B(n17681), .Z(n17291) );
  NAND U17783 ( .A(n17292), .B(n17291), .Z(n17294) );
  NANDN U17784 ( .A(n17293), .B(n17294), .Z(n17298) );
  XOR U17785 ( .A(n17294), .B(n17293), .Z(n17687) );
  NANDN U17786 ( .A(n17687), .B(n17686), .Z(n17297) );
  NAND U17787 ( .A(n17298), .B(n17297), .Z(n17300) );
  NANDN U17788 ( .A(n17299), .B(n17300), .Z(n17304) );
  XOR U17789 ( .A(n17300), .B(n17299), .Z(n17693) );
  XNOR U17790 ( .A(n17302), .B(n17301), .Z(n17692) );
  NANDN U17791 ( .A(n17693), .B(n17692), .Z(n17303) );
  NAND U17792 ( .A(n17304), .B(n17303), .Z(n17305) );
  OR U17793 ( .A(n17306), .B(n17305), .Z(n17310) );
  XNOR U17794 ( .A(n17306), .B(n17305), .Z(n17700) );
  NANDN U17795 ( .A(n17700), .B(n17701), .Z(n17309) );
  NAND U17796 ( .A(n17310), .B(n17309), .Z(n17312) );
  NAND U17797 ( .A(b[12]), .B(a[56]), .Z(n17311) );
  OR U17798 ( .A(n17312), .B(n17311), .Z(n17316) );
  XOR U17799 ( .A(n17312), .B(n17311), .Z(n17704) );
  XNOR U17800 ( .A(n17314), .B(n17313), .Z(n17705) );
  NAND U17801 ( .A(n17704), .B(n17705), .Z(n17315) );
  NAND U17802 ( .A(n17316), .B(n17315), .Z(n17317) );
  OR U17803 ( .A(n17318), .B(n17317), .Z(n17322) );
  XNOR U17804 ( .A(n17318), .B(n17317), .Z(n17712) );
  NANDN U17805 ( .A(n17712), .B(n17713), .Z(n17321) );
  NAND U17806 ( .A(n17322), .B(n17321), .Z(n17324) );
  NAND U17807 ( .A(b[12]), .B(a[58]), .Z(n17323) );
  OR U17808 ( .A(n17324), .B(n17323), .Z(n17328) );
  XOR U17809 ( .A(n17324), .B(n17323), .Z(n17716) );
  XNOR U17810 ( .A(n17326), .B(n17325), .Z(n17717) );
  NAND U17811 ( .A(n17716), .B(n17717), .Z(n17327) );
  NAND U17812 ( .A(n17328), .B(n17327), .Z(n17331) );
  OR U17813 ( .A(n17332), .B(n17331), .Z(n17334) );
  XOR U17814 ( .A(n17332), .B(n17331), .Z(n17722) );
  NAND U17815 ( .A(n17723), .B(n17722), .Z(n17333) );
  NAND U17816 ( .A(n17334), .B(n17333), .Z(n17336) );
  NAND U17817 ( .A(b[12]), .B(a[60]), .Z(n17335) );
  OR U17818 ( .A(n17336), .B(n17335), .Z(n17340) );
  XOR U17819 ( .A(n17336), .B(n17335), .Z(n17728) );
  XNOR U17820 ( .A(n17338), .B(n17337), .Z(n17729) );
  NAND U17821 ( .A(n17728), .B(n17729), .Z(n17339) );
  NAND U17822 ( .A(n17340), .B(n17339), .Z(n17343) );
  OR U17823 ( .A(n17344), .B(n17343), .Z(n17346) );
  XOR U17824 ( .A(n17344), .B(n17343), .Z(n17734) );
  NAND U17825 ( .A(n17735), .B(n17734), .Z(n17345) );
  NAND U17826 ( .A(n17346), .B(n17345), .Z(n17350) );
  NAND U17827 ( .A(b[12]), .B(a[62]), .Z(n17349) );
  OR U17828 ( .A(n17350), .B(n17349), .Z(n17352) );
  XOR U17829 ( .A(n17348), .B(n17347), .Z(n17369) );
  XOR U17830 ( .A(n17350), .B(n17349), .Z(n17370) );
  NANDN U17831 ( .A(n17369), .B(n17370), .Z(n17351) );
  NAND U17832 ( .A(n17352), .B(n17351), .Z(n17355) );
  AND U17833 ( .A(a[63]), .B(b[12]), .Z(n17356) );
  OR U17834 ( .A(n17355), .B(n17356), .Z(n17358) );
  XOR U17835 ( .A(n17354), .B(n17353), .Z(n17368) );
  XOR U17836 ( .A(n17356), .B(n17355), .Z(n17367) );
  NAND U17837 ( .A(n17368), .B(n17367), .Z(n17357) );
  NAND U17838 ( .A(n17358), .B(n17357), .Z(n18499) );
  OR U17839 ( .A(n18500), .B(n18499), .Z(n24139) );
  XNOR U17840 ( .A(n17360), .B(n17359), .Z(n21952) );
  NANDN U17841 ( .A(n17362), .B(n17361), .Z(n17366) );
  NANDN U17842 ( .A(n17364), .B(n17363), .Z(n17365) );
  AND U17843 ( .A(n17366), .B(n17365), .Z(n21953) );
  XOR U17844 ( .A(n21952), .B(n21953), .Z(n24138) );
  ANDN U17845 ( .B(n24139), .A(n24138), .Z(n21951) );
  XOR U17846 ( .A(n17368), .B(n17367), .Z(n21941) );
  XNOR U17847 ( .A(n17370), .B(n17369), .Z(n17741) );
  ANDN U17848 ( .B(b[11]), .A(n210), .Z(n17740) );
  NAND U17849 ( .A(a[62]), .B(b[11]), .Z(n17736) );
  NAND U17850 ( .A(a[60]), .B(b[11]), .Z(n17724) );
  ANDN U17851 ( .B(b[11]), .A(n197), .Z(n17657) );
  ANDN U17852 ( .B(b[11]), .A(n195), .Z(n17645) );
  ANDN U17853 ( .B(b[11]), .A(n193), .Z(n17633) );
  ANDN U17854 ( .B(b[11]), .A(n191), .Z(n17621) );
  ANDN U17855 ( .B(b[11]), .A(n189), .Z(n17609) );
  ANDN U17856 ( .B(b[11]), .A(n187), .Z(n17597) );
  ANDN U17857 ( .B(b[11]), .A(n21772), .Z(n17585) );
  ANDN U17858 ( .B(b[11]), .A(n184), .Z(n17573) );
  ANDN U17859 ( .B(b[11]), .A(n21751), .Z(n17561) );
  ANDN U17860 ( .B(b[11]), .A(n21740), .Z(n17549) );
  ANDN U17861 ( .B(b[11]), .A(n21727), .Z(n17537) );
  ANDN U17862 ( .B(b[11]), .A(n21716), .Z(n17525) );
  ANDN U17863 ( .B(b[11]), .A(n21703), .Z(n17513) );
  ANDN U17864 ( .B(b[11]), .A(n21692), .Z(n17501) );
  ANDN U17865 ( .B(b[11]), .A(n21681), .Z(n17489) );
  ANDN U17866 ( .B(b[11]), .A(n21670), .Z(n17477) );
  ANDN U17867 ( .B(b[11]), .A(n174), .Z(n17466) );
  XNOR U17868 ( .A(n17372), .B(n17371), .Z(n17461) );
  NAND U17869 ( .A(a[15]), .B(b[11]), .Z(n17455) );
  ANDN U17870 ( .B(b[11]), .A(n170), .Z(n17445) );
  ANDN U17871 ( .B(b[11]), .A(n21164), .Z(n17431) );
  ANDN U17872 ( .B(b[11]), .A(n21615), .Z(n17419) );
  ANDN U17873 ( .B(b[11]), .A(n166), .Z(n17407) );
  ANDN U17874 ( .B(b[11]), .A(n164), .Z(n17395) );
  ANDN U17875 ( .B(b[11]), .A(n21580), .Z(n17382) );
  NAND U17876 ( .A(b[12]), .B(a[1]), .Z(n17375) );
  AND U17877 ( .A(b[11]), .B(a[0]), .Z(n18133) );
  NANDN U17878 ( .A(n17375), .B(n18133), .Z(n17374) );
  NAND U17879 ( .A(a[2]), .B(b[11]), .Z(n17373) );
  AND U17880 ( .A(n17374), .B(n17373), .Z(n17381) );
  NANDN U17881 ( .A(n17375), .B(a[0]), .Z(n17376) );
  XNOR U17882 ( .A(a[2]), .B(n17376), .Z(n17377) );
  NAND U17883 ( .A(b[11]), .B(n17377), .Z(n17760) );
  AND U17884 ( .A(a[1]), .B(b[12]), .Z(n17378) );
  XNOR U17885 ( .A(n17379), .B(n17378), .Z(n17759) );
  NANDN U17886 ( .A(n17760), .B(n17759), .Z(n17380) );
  NANDN U17887 ( .A(n17381), .B(n17380), .Z(n17383) );
  NANDN U17888 ( .A(n17382), .B(n17383), .Z(n17387) );
  XOR U17889 ( .A(n17383), .B(n17382), .Z(n17764) );
  NANDN U17890 ( .A(n17764), .B(n17763), .Z(n17386) );
  NAND U17891 ( .A(n17387), .B(n17386), .Z(n17391) );
  XOR U17892 ( .A(n17389), .B(n17388), .Z(n17390) );
  NANDN U17893 ( .A(n17391), .B(n17390), .Z(n17393) );
  NAND U17894 ( .A(a[4]), .B(b[11]), .Z(n17771) );
  NANDN U17895 ( .A(n17771), .B(n17772), .Z(n17392) );
  NAND U17896 ( .A(n17393), .B(n17392), .Z(n17394) );
  OR U17897 ( .A(n17395), .B(n17394), .Z(n17399) );
  XNOR U17898 ( .A(n17395), .B(n17394), .Z(n17775) );
  XOR U17899 ( .A(n17397), .B(n17396), .Z(n17776) );
  NANDN U17900 ( .A(n17775), .B(n17776), .Z(n17398) );
  NAND U17901 ( .A(n17399), .B(n17398), .Z(n17402) );
  XOR U17902 ( .A(n17401), .B(n17400), .Z(n17403) );
  NANDN U17903 ( .A(n17402), .B(n17403), .Z(n17405) );
  NAND U17904 ( .A(a[6]), .B(b[11]), .Z(n17783) );
  XNOR U17905 ( .A(n17403), .B(n17402), .Z(n17784) );
  NANDN U17906 ( .A(n17783), .B(n17784), .Z(n17404) );
  NAND U17907 ( .A(n17405), .B(n17404), .Z(n17406) );
  OR U17908 ( .A(n17407), .B(n17406), .Z(n17411) );
  XNOR U17909 ( .A(n17407), .B(n17406), .Z(n17787) );
  XOR U17910 ( .A(n17409), .B(n17408), .Z(n17788) );
  NANDN U17911 ( .A(n17787), .B(n17788), .Z(n17410) );
  NAND U17912 ( .A(n17411), .B(n17410), .Z(n17414) );
  XOR U17913 ( .A(n17413), .B(n17412), .Z(n17415) );
  NANDN U17914 ( .A(n17414), .B(n17415), .Z(n17417) );
  NAND U17915 ( .A(a[8]), .B(b[11]), .Z(n17795) );
  XNOR U17916 ( .A(n17415), .B(n17414), .Z(n17796) );
  NANDN U17917 ( .A(n17795), .B(n17796), .Z(n17416) );
  NAND U17918 ( .A(n17417), .B(n17416), .Z(n17418) );
  OR U17919 ( .A(n17419), .B(n17418), .Z(n17423) );
  XNOR U17920 ( .A(n17419), .B(n17418), .Z(n17799) );
  XOR U17921 ( .A(n17421), .B(n17420), .Z(n17800) );
  NANDN U17922 ( .A(n17799), .B(n17800), .Z(n17422) );
  NAND U17923 ( .A(n17423), .B(n17422), .Z(n17426) );
  XOR U17924 ( .A(n17425), .B(n17424), .Z(n17427) );
  NANDN U17925 ( .A(n17426), .B(n17427), .Z(n17429) );
  NAND U17926 ( .A(a[10]), .B(b[11]), .Z(n17807) );
  XNOR U17927 ( .A(n17427), .B(n17426), .Z(n17808) );
  NANDN U17928 ( .A(n17807), .B(n17808), .Z(n17428) );
  NAND U17929 ( .A(n17429), .B(n17428), .Z(n17430) );
  OR U17930 ( .A(n17431), .B(n17430), .Z(n17435) );
  XNOR U17931 ( .A(n17431), .B(n17430), .Z(n17811) );
  XOR U17932 ( .A(n17433), .B(n17432), .Z(n17812) );
  NANDN U17933 ( .A(n17811), .B(n17812), .Z(n17434) );
  NAND U17934 ( .A(n17435), .B(n17434), .Z(n17438) );
  NANDN U17935 ( .A(n17438), .B(n17439), .Z(n17441) );
  NAND U17936 ( .A(a[12]), .B(b[11]), .Z(n17819) );
  XNOR U17937 ( .A(n17439), .B(n17438), .Z(n17820) );
  NANDN U17938 ( .A(n17819), .B(n17820), .Z(n17440) );
  NAND U17939 ( .A(n17441), .B(n17440), .Z(n17444) );
  OR U17940 ( .A(n17445), .B(n17444), .Z(n17447) );
  XOR U17941 ( .A(n17445), .B(n17444), .Z(n17823) );
  NANDN U17942 ( .A(n17824), .B(n17823), .Z(n17446) );
  NAND U17943 ( .A(n17447), .B(n17446), .Z(n17450) );
  XOR U17944 ( .A(n17449), .B(n17448), .Z(n17451) );
  NANDN U17945 ( .A(n17450), .B(n17451), .Z(n17453) );
  NAND U17946 ( .A(a[14]), .B(b[11]), .Z(n17831) );
  XNOR U17947 ( .A(n17451), .B(n17450), .Z(n17832) );
  NANDN U17948 ( .A(n17831), .B(n17832), .Z(n17452) );
  NAND U17949 ( .A(n17453), .B(n17452), .Z(n17454) );
  NANDN U17950 ( .A(n17455), .B(n17454), .Z(n17459) );
  XNOR U17951 ( .A(n17457), .B(n17456), .Z(n17747) );
  NAND U17952 ( .A(n17746), .B(n17747), .Z(n17458) );
  AND U17953 ( .A(n17459), .B(n17458), .Z(n17460) );
  NANDN U17954 ( .A(n17461), .B(n17460), .Z(n17463) );
  ANDN U17955 ( .B(b[11]), .A(n173), .Z(n17840) );
  NANDN U17956 ( .A(n17840), .B(n17839), .Z(n17462) );
  NAND U17957 ( .A(n17463), .B(n17462), .Z(n17467) );
  NANDN U17958 ( .A(n17466), .B(n17467), .Z(n17469) );
  XNOR U17959 ( .A(n17465), .B(n17464), .Z(n17846) );
  XOR U17960 ( .A(n17467), .B(n17466), .Z(n17845) );
  OR U17961 ( .A(n17846), .B(n17845), .Z(n17468) );
  NAND U17962 ( .A(n17469), .B(n17468), .Z(n17473) );
  XOR U17963 ( .A(n17471), .B(n17470), .Z(n17472) );
  NANDN U17964 ( .A(n17473), .B(n17472), .Z(n17475) );
  NAND U17965 ( .A(a[18]), .B(b[11]), .Z(n17853) );
  NANDN U17966 ( .A(n17853), .B(n17854), .Z(n17474) );
  NAND U17967 ( .A(n17475), .B(n17474), .Z(n17476) );
  OR U17968 ( .A(n17477), .B(n17476), .Z(n17481) );
  XNOR U17969 ( .A(n17477), .B(n17476), .Z(n17857) );
  XOR U17970 ( .A(n17479), .B(n17478), .Z(n17858) );
  NANDN U17971 ( .A(n17857), .B(n17858), .Z(n17480) );
  NAND U17972 ( .A(n17481), .B(n17480), .Z(n17484) );
  NANDN U17973 ( .A(n17484), .B(n17485), .Z(n17487) );
  NAND U17974 ( .A(a[20]), .B(b[11]), .Z(n17865) );
  XNOR U17975 ( .A(n17485), .B(n17484), .Z(n17866) );
  NANDN U17976 ( .A(n17865), .B(n17866), .Z(n17486) );
  NAND U17977 ( .A(n17487), .B(n17486), .Z(n17488) );
  OR U17978 ( .A(n17489), .B(n17488), .Z(n17493) );
  XNOR U17979 ( .A(n17489), .B(n17488), .Z(n17869) );
  XOR U17980 ( .A(n17491), .B(n17490), .Z(n17870) );
  NANDN U17981 ( .A(n17869), .B(n17870), .Z(n17492) );
  NAND U17982 ( .A(n17493), .B(n17492), .Z(n17496) );
  NANDN U17983 ( .A(n17496), .B(n17497), .Z(n17499) );
  NAND U17984 ( .A(a[22]), .B(b[11]), .Z(n17877) );
  XNOR U17985 ( .A(n17497), .B(n17496), .Z(n17878) );
  NANDN U17986 ( .A(n17877), .B(n17878), .Z(n17498) );
  NAND U17987 ( .A(n17499), .B(n17498), .Z(n17500) );
  OR U17988 ( .A(n17501), .B(n17500), .Z(n17505) );
  XNOR U17989 ( .A(n17501), .B(n17500), .Z(n17881) );
  XOR U17990 ( .A(n17503), .B(n17502), .Z(n17882) );
  NANDN U17991 ( .A(n17881), .B(n17882), .Z(n17504) );
  NAND U17992 ( .A(n17505), .B(n17504), .Z(n17508) );
  NANDN U17993 ( .A(n17508), .B(n17509), .Z(n17511) );
  NAND U17994 ( .A(a[24]), .B(b[11]), .Z(n17889) );
  XNOR U17995 ( .A(n17509), .B(n17508), .Z(n17890) );
  NANDN U17996 ( .A(n17889), .B(n17890), .Z(n17510) );
  NAND U17997 ( .A(n17511), .B(n17510), .Z(n17512) );
  OR U17998 ( .A(n17513), .B(n17512), .Z(n17517) );
  XNOR U17999 ( .A(n17513), .B(n17512), .Z(n17893) );
  XOR U18000 ( .A(n17515), .B(n17514), .Z(n17894) );
  NANDN U18001 ( .A(n17893), .B(n17894), .Z(n17516) );
  NAND U18002 ( .A(n17517), .B(n17516), .Z(n17521) );
  XOR U18003 ( .A(n17519), .B(n17518), .Z(n17520) );
  NANDN U18004 ( .A(n17521), .B(n17520), .Z(n17523) );
  NAND U18005 ( .A(a[26]), .B(b[11]), .Z(n17901) );
  NANDN U18006 ( .A(n17901), .B(n17902), .Z(n17522) );
  NAND U18007 ( .A(n17523), .B(n17522), .Z(n17524) );
  OR U18008 ( .A(n17525), .B(n17524), .Z(n17529) );
  XNOR U18009 ( .A(n17525), .B(n17524), .Z(n17905) );
  XOR U18010 ( .A(n17527), .B(n17526), .Z(n17906) );
  NANDN U18011 ( .A(n17905), .B(n17906), .Z(n17528) );
  NAND U18012 ( .A(n17529), .B(n17528), .Z(n17532) );
  NANDN U18013 ( .A(n17532), .B(n17533), .Z(n17535) );
  NAND U18014 ( .A(a[28]), .B(b[11]), .Z(n17913) );
  XNOR U18015 ( .A(n17533), .B(n17532), .Z(n17914) );
  NANDN U18016 ( .A(n17913), .B(n17914), .Z(n17534) );
  NAND U18017 ( .A(n17535), .B(n17534), .Z(n17536) );
  OR U18018 ( .A(n17537), .B(n17536), .Z(n17541) );
  XNOR U18019 ( .A(n17537), .B(n17536), .Z(n17917) );
  XOR U18020 ( .A(n17539), .B(n17538), .Z(n17918) );
  NANDN U18021 ( .A(n17917), .B(n17918), .Z(n17540) );
  NAND U18022 ( .A(n17541), .B(n17540), .Z(n17544) );
  NANDN U18023 ( .A(n17544), .B(n17545), .Z(n17547) );
  NAND U18024 ( .A(a[30]), .B(b[11]), .Z(n17925) );
  XNOR U18025 ( .A(n17545), .B(n17544), .Z(n17926) );
  NANDN U18026 ( .A(n17925), .B(n17926), .Z(n17546) );
  NAND U18027 ( .A(n17547), .B(n17546), .Z(n17548) );
  OR U18028 ( .A(n17549), .B(n17548), .Z(n17553) );
  XNOR U18029 ( .A(n17549), .B(n17548), .Z(n17929) );
  XOR U18030 ( .A(n17551), .B(n17550), .Z(n17930) );
  NANDN U18031 ( .A(n17929), .B(n17930), .Z(n17552) );
  NAND U18032 ( .A(n17553), .B(n17552), .Z(n17556) );
  NANDN U18033 ( .A(n17556), .B(n17557), .Z(n17559) );
  NAND U18034 ( .A(a[32]), .B(b[11]), .Z(n17937) );
  XNOR U18035 ( .A(n17557), .B(n17556), .Z(n17938) );
  NANDN U18036 ( .A(n17937), .B(n17938), .Z(n17558) );
  NAND U18037 ( .A(n17559), .B(n17558), .Z(n17560) );
  OR U18038 ( .A(n17561), .B(n17560), .Z(n17565) );
  XNOR U18039 ( .A(n17561), .B(n17560), .Z(n17941) );
  XOR U18040 ( .A(n17563), .B(n17562), .Z(n17942) );
  NANDN U18041 ( .A(n17941), .B(n17942), .Z(n17564) );
  NAND U18042 ( .A(n17565), .B(n17564), .Z(n17568) );
  NANDN U18043 ( .A(n17568), .B(n17569), .Z(n17571) );
  NAND U18044 ( .A(a[34]), .B(b[11]), .Z(n17949) );
  XNOR U18045 ( .A(n17569), .B(n17568), .Z(n17950) );
  NANDN U18046 ( .A(n17949), .B(n17950), .Z(n17570) );
  NAND U18047 ( .A(n17571), .B(n17570), .Z(n17572) );
  OR U18048 ( .A(n17573), .B(n17572), .Z(n17577) );
  XNOR U18049 ( .A(n17573), .B(n17572), .Z(n17953) );
  XOR U18050 ( .A(n17575), .B(n17574), .Z(n17954) );
  NANDN U18051 ( .A(n17953), .B(n17954), .Z(n17576) );
  NAND U18052 ( .A(n17577), .B(n17576), .Z(n17580) );
  NANDN U18053 ( .A(n17580), .B(n17581), .Z(n17583) );
  NAND U18054 ( .A(a[36]), .B(b[11]), .Z(n17961) );
  XNOR U18055 ( .A(n17581), .B(n17580), .Z(n17962) );
  NANDN U18056 ( .A(n17961), .B(n17962), .Z(n17582) );
  NAND U18057 ( .A(n17583), .B(n17582), .Z(n17584) );
  OR U18058 ( .A(n17585), .B(n17584), .Z(n17589) );
  XNOR U18059 ( .A(n17585), .B(n17584), .Z(n17965) );
  XOR U18060 ( .A(n17587), .B(n17586), .Z(n17966) );
  NANDN U18061 ( .A(n17965), .B(n17966), .Z(n17588) );
  NAND U18062 ( .A(n17589), .B(n17588), .Z(n17592) );
  NANDN U18063 ( .A(n17592), .B(n17593), .Z(n17595) );
  NAND U18064 ( .A(a[38]), .B(b[11]), .Z(n17973) );
  XNOR U18065 ( .A(n17593), .B(n17592), .Z(n17974) );
  NANDN U18066 ( .A(n17973), .B(n17974), .Z(n17594) );
  NAND U18067 ( .A(n17595), .B(n17594), .Z(n17596) );
  OR U18068 ( .A(n17597), .B(n17596), .Z(n17601) );
  XNOR U18069 ( .A(n17597), .B(n17596), .Z(n17977) );
  XOR U18070 ( .A(n17599), .B(n17598), .Z(n17978) );
  NANDN U18071 ( .A(n17977), .B(n17978), .Z(n17600) );
  NAND U18072 ( .A(n17601), .B(n17600), .Z(n17604) );
  NANDN U18073 ( .A(n17604), .B(n17605), .Z(n17607) );
  NAND U18074 ( .A(a[40]), .B(b[11]), .Z(n17985) );
  XNOR U18075 ( .A(n17605), .B(n17604), .Z(n17986) );
  NANDN U18076 ( .A(n17985), .B(n17986), .Z(n17606) );
  NAND U18077 ( .A(n17607), .B(n17606), .Z(n17608) );
  OR U18078 ( .A(n17609), .B(n17608), .Z(n17613) );
  XNOR U18079 ( .A(n17609), .B(n17608), .Z(n17989) );
  XOR U18080 ( .A(n17611), .B(n17610), .Z(n17990) );
  NANDN U18081 ( .A(n17989), .B(n17990), .Z(n17612) );
  NAND U18082 ( .A(n17613), .B(n17612), .Z(n17616) );
  NANDN U18083 ( .A(n17616), .B(n17617), .Z(n17619) );
  NAND U18084 ( .A(a[42]), .B(b[11]), .Z(n17997) );
  XNOR U18085 ( .A(n17617), .B(n17616), .Z(n17998) );
  NANDN U18086 ( .A(n17997), .B(n17998), .Z(n17618) );
  NAND U18087 ( .A(n17619), .B(n17618), .Z(n17620) );
  OR U18088 ( .A(n17621), .B(n17620), .Z(n17625) );
  XNOR U18089 ( .A(n17621), .B(n17620), .Z(n18001) );
  XOR U18090 ( .A(n17623), .B(n17622), .Z(n18002) );
  NANDN U18091 ( .A(n18001), .B(n18002), .Z(n17624) );
  NAND U18092 ( .A(n17625), .B(n17624), .Z(n17628) );
  NANDN U18093 ( .A(n17628), .B(n17629), .Z(n17631) );
  NAND U18094 ( .A(a[44]), .B(b[11]), .Z(n18009) );
  XNOR U18095 ( .A(n17629), .B(n17628), .Z(n18010) );
  NANDN U18096 ( .A(n18009), .B(n18010), .Z(n17630) );
  NAND U18097 ( .A(n17631), .B(n17630), .Z(n17632) );
  OR U18098 ( .A(n17633), .B(n17632), .Z(n17637) );
  XNOR U18099 ( .A(n17633), .B(n17632), .Z(n18013) );
  XOR U18100 ( .A(n17635), .B(n17634), .Z(n18014) );
  NANDN U18101 ( .A(n18013), .B(n18014), .Z(n17636) );
  NAND U18102 ( .A(n17637), .B(n17636), .Z(n17640) );
  NANDN U18103 ( .A(n17640), .B(n17641), .Z(n17643) );
  NAND U18104 ( .A(a[46]), .B(b[11]), .Z(n18021) );
  XNOR U18105 ( .A(n17641), .B(n17640), .Z(n18022) );
  NANDN U18106 ( .A(n18021), .B(n18022), .Z(n17642) );
  NAND U18107 ( .A(n17643), .B(n17642), .Z(n17644) );
  OR U18108 ( .A(n17645), .B(n17644), .Z(n17649) );
  XNOR U18109 ( .A(n17645), .B(n17644), .Z(n18025) );
  XOR U18110 ( .A(n17647), .B(n17646), .Z(n18026) );
  NANDN U18111 ( .A(n18025), .B(n18026), .Z(n17648) );
  NAND U18112 ( .A(n17649), .B(n17648), .Z(n17652) );
  NANDN U18113 ( .A(n17652), .B(n17653), .Z(n17655) );
  NAND U18114 ( .A(a[48]), .B(b[11]), .Z(n18033) );
  XNOR U18115 ( .A(n17653), .B(n17652), .Z(n18034) );
  NANDN U18116 ( .A(n18033), .B(n18034), .Z(n17654) );
  NAND U18117 ( .A(n17655), .B(n17654), .Z(n17656) );
  OR U18118 ( .A(n17657), .B(n17656), .Z(n17661) );
  XNOR U18119 ( .A(n17657), .B(n17656), .Z(n18037) );
  XOR U18120 ( .A(n17659), .B(n17658), .Z(n18038) );
  NANDN U18121 ( .A(n18037), .B(n18038), .Z(n17660) );
  NAND U18122 ( .A(n17661), .B(n17660), .Z(n17664) );
  NANDN U18123 ( .A(n17664), .B(n17665), .Z(n17667) );
  NAND U18124 ( .A(a[50]), .B(b[11]), .Z(n18045) );
  XNOR U18125 ( .A(n17665), .B(n17664), .Z(n18046) );
  NANDN U18126 ( .A(n18045), .B(n18046), .Z(n17666) );
  NAND U18127 ( .A(n17667), .B(n17666), .Z(n17670) );
  ANDN U18128 ( .B(b[11]), .A(n199), .Z(n17671) );
  OR U18129 ( .A(n17670), .B(n17671), .Z(n17673) );
  XOR U18130 ( .A(n17669), .B(n17668), .Z(n18050) );
  XOR U18131 ( .A(n17671), .B(n17670), .Z(n18049) );
  NANDN U18132 ( .A(n18050), .B(n18049), .Z(n17672) );
  NAND U18133 ( .A(n17673), .B(n17672), .Z(n17677) );
  XOR U18134 ( .A(n17675), .B(n17674), .Z(n17676) );
  NANDN U18135 ( .A(n17677), .B(n17676), .Z(n17679) );
  NAND U18136 ( .A(a[52]), .B(b[11]), .Z(n18056) );
  NANDN U18137 ( .A(n18056), .B(n18055), .Z(n17678) );
  NAND U18138 ( .A(n17679), .B(n17678), .Z(n17682) );
  ANDN U18139 ( .B(b[11]), .A(n201), .Z(n17683) );
  OR U18140 ( .A(n17682), .B(n17683), .Z(n17685) );
  XNOR U18141 ( .A(n17681), .B(n17680), .Z(n18064) );
  XOR U18142 ( .A(n17683), .B(n17682), .Z(n18063) );
  NANDN U18143 ( .A(n18064), .B(n18063), .Z(n17684) );
  NAND U18144 ( .A(n17685), .B(n17684), .Z(n17689) );
  AND U18145 ( .A(b[11]), .B(a[54]), .Z(n17688) );
  NANDN U18146 ( .A(n17689), .B(n17688), .Z(n17691) );
  XOR U18147 ( .A(n17687), .B(n17686), .Z(n17744) );
  XNOR U18148 ( .A(n17689), .B(n17688), .Z(n17745) );
  NANDN U18149 ( .A(n17744), .B(n17745), .Z(n17690) );
  AND U18150 ( .A(n17691), .B(n17690), .Z(n17695) );
  XNOR U18151 ( .A(n17693), .B(n17692), .Z(n17694) );
  NANDN U18152 ( .A(n17695), .B(n17694), .Z(n17697) );
  AND U18153 ( .A(b[11]), .B(a[55]), .Z(n18073) );
  NANDN U18154 ( .A(n18074), .B(n18073), .Z(n17696) );
  AND U18155 ( .A(n17697), .B(n17696), .Z(n17699) );
  AND U18156 ( .A(b[11]), .B(a[56]), .Z(n17698) );
  NANDN U18157 ( .A(n17699), .B(n17698), .Z(n17703) );
  XOR U18158 ( .A(n17699), .B(n17698), .Z(n18077) );
  XOR U18159 ( .A(n17701), .B(n17700), .Z(n18078) );
  NANDN U18160 ( .A(n18077), .B(n18078), .Z(n17702) );
  AND U18161 ( .A(n17703), .B(n17702), .Z(n17707) );
  NANDN U18162 ( .A(n17707), .B(n17706), .Z(n17709) );
  XOR U18163 ( .A(n17707), .B(n17706), .Z(n18086) );
  AND U18164 ( .A(b[11]), .B(a[57]), .Z(n18085) );
  NANDN U18165 ( .A(n18086), .B(n18085), .Z(n17708) );
  AND U18166 ( .A(n17709), .B(n17708), .Z(n17711) );
  AND U18167 ( .A(b[11]), .B(a[58]), .Z(n17710) );
  NANDN U18168 ( .A(n17711), .B(n17710), .Z(n17715) );
  XOR U18169 ( .A(n17711), .B(n17710), .Z(n18089) );
  XOR U18170 ( .A(n17713), .B(n17712), .Z(n18090) );
  NANDN U18171 ( .A(n18089), .B(n18090), .Z(n17714) );
  AND U18172 ( .A(n17715), .B(n17714), .Z(n17719) );
  NANDN U18173 ( .A(n17719), .B(n17718), .Z(n17721) );
  XOR U18174 ( .A(n17719), .B(n17718), .Z(n18098) );
  NAND U18175 ( .A(a[59]), .B(b[11]), .Z(n18097) );
  OR U18176 ( .A(n18098), .B(n18097), .Z(n17720) );
  AND U18177 ( .A(n17721), .B(n17720), .Z(n17725) );
  OR U18178 ( .A(n17724), .B(n17725), .Z(n17727) );
  XOR U18179 ( .A(n17723), .B(n17722), .Z(n18104) );
  XOR U18180 ( .A(n17725), .B(n17724), .Z(n18103) );
  NANDN U18181 ( .A(n18104), .B(n18103), .Z(n17726) );
  AND U18182 ( .A(n17727), .B(n17726), .Z(n17731) );
  NANDN U18183 ( .A(n17731), .B(n17730), .Z(n17733) );
  XOR U18184 ( .A(n17731), .B(n17730), .Z(n18110) );
  NAND U18185 ( .A(a[61]), .B(b[11]), .Z(n18109) );
  OR U18186 ( .A(n18110), .B(n18109), .Z(n17732) );
  AND U18187 ( .A(n17733), .B(n17732), .Z(n17737) );
  OR U18188 ( .A(n17736), .B(n17737), .Z(n17739) );
  XOR U18189 ( .A(n17735), .B(n17734), .Z(n18116) );
  XOR U18190 ( .A(n17737), .B(n17736), .Z(n18115) );
  NANDN U18191 ( .A(n18116), .B(n18115), .Z(n17738) );
  AND U18192 ( .A(n17739), .B(n17738), .Z(n17743) );
  XOR U18193 ( .A(n17741), .B(n17740), .Z(n17742) );
  XOR U18194 ( .A(n21941), .B(n21942), .Z(n24126) );
  XOR U18195 ( .A(n17743), .B(n17742), .Z(n18497) );
  ANDN U18196 ( .B(b[10]), .A(n207), .Z(n18092) );
  ANDN U18197 ( .B(b[10]), .A(n205), .Z(n18080) );
  NAND U18198 ( .A(a[56]), .B(b[10]), .Z(n18072) );
  XOR U18199 ( .A(n17745), .B(n17744), .Z(n18067) );
  ANDN U18200 ( .B(b[10]), .A(n199), .Z(n18044) );
  ANDN U18201 ( .B(b[10]), .A(n197), .Z(n18032) );
  ANDN U18202 ( .B(b[10]), .A(n195), .Z(n18020) );
  ANDN U18203 ( .B(b[10]), .A(n193), .Z(n18008) );
  ANDN U18204 ( .B(b[10]), .A(n191), .Z(n17996) );
  ANDN U18205 ( .B(b[10]), .A(n189), .Z(n17984) );
  ANDN U18206 ( .B(b[10]), .A(n187), .Z(n17972) );
  ANDN U18207 ( .B(b[10]), .A(n21772), .Z(n17960) );
  ANDN U18208 ( .B(b[10]), .A(n184), .Z(n17948) );
  ANDN U18209 ( .B(b[10]), .A(n21751), .Z(n17936) );
  ANDN U18210 ( .B(b[10]), .A(n21740), .Z(n17924) );
  ANDN U18211 ( .B(b[10]), .A(n21727), .Z(n17912) );
  ANDN U18212 ( .B(b[10]), .A(n21716), .Z(n17900) );
  ANDN U18213 ( .B(b[10]), .A(n21703), .Z(n17888) );
  ANDN U18214 ( .B(b[10]), .A(n21692), .Z(n17876) );
  ANDN U18215 ( .B(b[10]), .A(n21681), .Z(n17864) );
  ANDN U18216 ( .B(b[10]), .A(n21670), .Z(n17852) );
  ANDN U18217 ( .B(b[10]), .A(n174), .Z(n17842) );
  NAND U18218 ( .A(a[16]), .B(b[10]), .Z(n17836) );
  NANDN U18219 ( .A(n17836), .B(n17835), .Z(n17838) );
  ANDN U18220 ( .B(b[10]), .A(n172), .Z(n17830) );
  ANDN U18221 ( .B(b[10]), .A(n170), .Z(n17818) );
  ANDN U18222 ( .B(b[10]), .A(n21164), .Z(n17806) );
  ANDN U18223 ( .B(b[10]), .A(n21615), .Z(n17794) );
  ANDN U18224 ( .B(b[10]), .A(n166), .Z(n17782) );
  ANDN U18225 ( .B(b[10]), .A(n164), .Z(n17770) );
  ANDN U18226 ( .B(b[10]), .A(n21580), .Z(n17757) );
  NAND U18227 ( .A(b[11]), .B(a[1]), .Z(n17750) );
  AND U18228 ( .A(b[10]), .B(a[0]), .Z(n18513) );
  NANDN U18229 ( .A(n17750), .B(n18513), .Z(n17749) );
  NAND U18230 ( .A(a[2]), .B(b[10]), .Z(n17748) );
  AND U18231 ( .A(n17749), .B(n17748), .Z(n17756) );
  NANDN U18232 ( .A(n17750), .B(a[0]), .Z(n17751) );
  XNOR U18233 ( .A(a[2]), .B(n17751), .Z(n17752) );
  NAND U18234 ( .A(b[10]), .B(n17752), .Z(n18139) );
  AND U18235 ( .A(a[1]), .B(b[11]), .Z(n17753) );
  XNOR U18236 ( .A(n17754), .B(n17753), .Z(n18138) );
  NANDN U18237 ( .A(n18139), .B(n18138), .Z(n17755) );
  NANDN U18238 ( .A(n17756), .B(n17755), .Z(n17758) );
  NANDN U18239 ( .A(n17757), .B(n17758), .Z(n17762) );
  XOR U18240 ( .A(n17758), .B(n17757), .Z(n18143) );
  NANDN U18241 ( .A(n18143), .B(n18142), .Z(n17761) );
  NAND U18242 ( .A(n17762), .B(n17761), .Z(n17766) );
  XOR U18243 ( .A(n17764), .B(n17763), .Z(n17765) );
  NANDN U18244 ( .A(n17766), .B(n17765), .Z(n17768) );
  NAND U18245 ( .A(a[4]), .B(b[10]), .Z(n18150) );
  NANDN U18246 ( .A(n18150), .B(n18151), .Z(n17767) );
  NAND U18247 ( .A(n17768), .B(n17767), .Z(n17769) );
  OR U18248 ( .A(n17770), .B(n17769), .Z(n17774) );
  XNOR U18249 ( .A(n17770), .B(n17769), .Z(n18125) );
  XOR U18250 ( .A(n17772), .B(n17771), .Z(n18126) );
  NANDN U18251 ( .A(n18125), .B(n18126), .Z(n17773) );
  NAND U18252 ( .A(n17774), .B(n17773), .Z(n17777) );
  XOR U18253 ( .A(n17776), .B(n17775), .Z(n17778) );
  NANDN U18254 ( .A(n17777), .B(n17778), .Z(n17780) );
  NAND U18255 ( .A(a[6]), .B(b[10]), .Z(n18160) );
  XNOR U18256 ( .A(n17778), .B(n17777), .Z(n18161) );
  NANDN U18257 ( .A(n18160), .B(n18161), .Z(n17779) );
  NAND U18258 ( .A(n17780), .B(n17779), .Z(n17781) );
  OR U18259 ( .A(n17782), .B(n17781), .Z(n17786) );
  XNOR U18260 ( .A(n17782), .B(n17781), .Z(n18164) );
  XOR U18261 ( .A(n17784), .B(n17783), .Z(n18165) );
  NANDN U18262 ( .A(n18164), .B(n18165), .Z(n17785) );
  NAND U18263 ( .A(n17786), .B(n17785), .Z(n17789) );
  XOR U18264 ( .A(n17788), .B(n17787), .Z(n17790) );
  NANDN U18265 ( .A(n17789), .B(n17790), .Z(n17792) );
  NAND U18266 ( .A(a[8]), .B(b[10]), .Z(n18172) );
  XNOR U18267 ( .A(n17790), .B(n17789), .Z(n18173) );
  NANDN U18268 ( .A(n18172), .B(n18173), .Z(n17791) );
  NAND U18269 ( .A(n17792), .B(n17791), .Z(n17793) );
  OR U18270 ( .A(n17794), .B(n17793), .Z(n17798) );
  XNOR U18271 ( .A(n17794), .B(n17793), .Z(n18176) );
  XOR U18272 ( .A(n17796), .B(n17795), .Z(n18177) );
  NANDN U18273 ( .A(n18176), .B(n18177), .Z(n17797) );
  NAND U18274 ( .A(n17798), .B(n17797), .Z(n17802) );
  NAND U18275 ( .A(a[10]), .B(b[10]), .Z(n17801) );
  OR U18276 ( .A(n17802), .B(n17801), .Z(n17804) );
  XOR U18277 ( .A(n17800), .B(n17799), .Z(n18183) );
  XOR U18278 ( .A(n17802), .B(n17801), .Z(n18182) );
  NAND U18279 ( .A(n18183), .B(n18182), .Z(n17803) );
  NAND U18280 ( .A(n17804), .B(n17803), .Z(n17805) );
  OR U18281 ( .A(n17806), .B(n17805), .Z(n17810) );
  XNOR U18282 ( .A(n17806), .B(n17805), .Z(n18188) );
  XOR U18283 ( .A(n17808), .B(n17807), .Z(n18189) );
  NANDN U18284 ( .A(n18188), .B(n18189), .Z(n17809) );
  NAND U18285 ( .A(n17810), .B(n17809), .Z(n17814) );
  NAND U18286 ( .A(a[12]), .B(b[10]), .Z(n17813) );
  OR U18287 ( .A(n17814), .B(n17813), .Z(n17816) );
  XOR U18288 ( .A(n17812), .B(n17811), .Z(n18195) );
  XOR U18289 ( .A(n17814), .B(n17813), .Z(n18194) );
  NAND U18290 ( .A(n18195), .B(n18194), .Z(n17815) );
  NAND U18291 ( .A(n17816), .B(n17815), .Z(n17817) );
  OR U18292 ( .A(n17818), .B(n17817), .Z(n17822) );
  XNOR U18293 ( .A(n17818), .B(n17817), .Z(n18200) );
  XOR U18294 ( .A(n17820), .B(n17819), .Z(n18201) );
  NANDN U18295 ( .A(n18200), .B(n18201), .Z(n17821) );
  NAND U18296 ( .A(n17822), .B(n17821), .Z(n17825) );
  NANDN U18297 ( .A(n17825), .B(n17826), .Z(n17828) );
  NAND U18298 ( .A(a[14]), .B(b[10]), .Z(n18206) );
  XNOR U18299 ( .A(n17826), .B(n17825), .Z(n18207) );
  NANDN U18300 ( .A(n18206), .B(n18207), .Z(n17827) );
  NAND U18301 ( .A(n17828), .B(n17827), .Z(n17829) );
  OR U18302 ( .A(n17830), .B(n17829), .Z(n17834) );
  XNOR U18303 ( .A(n17830), .B(n17829), .Z(n18123) );
  XOR U18304 ( .A(n17832), .B(n17831), .Z(n18124) );
  NANDN U18305 ( .A(n18123), .B(n18124), .Z(n17833) );
  NAND U18306 ( .A(n17834), .B(n17833), .Z(n18219) );
  XNOR U18307 ( .A(n17836), .B(n17835), .Z(n18218) );
  NANDN U18308 ( .A(n18219), .B(n18218), .Z(n17837) );
  NAND U18309 ( .A(n17838), .B(n17837), .Z(n17841) );
  OR U18310 ( .A(n17842), .B(n17841), .Z(n17844) );
  XOR U18311 ( .A(n17840), .B(n17839), .Z(n18222) );
  XOR U18312 ( .A(n17842), .B(n17841), .Z(n18223) );
  NANDN U18313 ( .A(n18222), .B(n18223), .Z(n17843) );
  NAND U18314 ( .A(n17844), .B(n17843), .Z(n17848) );
  XNOR U18315 ( .A(n17846), .B(n17845), .Z(n17847) );
  NANDN U18316 ( .A(n17848), .B(n17847), .Z(n17850) );
  NAND U18317 ( .A(a[18]), .B(b[10]), .Z(n18230) );
  NANDN U18318 ( .A(n18230), .B(n18231), .Z(n17849) );
  NAND U18319 ( .A(n17850), .B(n17849), .Z(n17851) );
  OR U18320 ( .A(n17852), .B(n17851), .Z(n17856) );
  XNOR U18321 ( .A(n17852), .B(n17851), .Z(n18234) );
  XOR U18322 ( .A(n17854), .B(n17853), .Z(n18235) );
  NANDN U18323 ( .A(n18234), .B(n18235), .Z(n17855) );
  NAND U18324 ( .A(n17856), .B(n17855), .Z(n17859) );
  XOR U18325 ( .A(n17858), .B(n17857), .Z(n17860) );
  NANDN U18326 ( .A(n17859), .B(n17860), .Z(n17862) );
  NAND U18327 ( .A(a[20]), .B(b[10]), .Z(n18242) );
  XNOR U18328 ( .A(n17860), .B(n17859), .Z(n18243) );
  NANDN U18329 ( .A(n18242), .B(n18243), .Z(n17861) );
  NAND U18330 ( .A(n17862), .B(n17861), .Z(n17863) );
  OR U18331 ( .A(n17864), .B(n17863), .Z(n17868) );
  XNOR U18332 ( .A(n17864), .B(n17863), .Z(n18246) );
  XOR U18333 ( .A(n17866), .B(n17865), .Z(n18247) );
  NANDN U18334 ( .A(n18246), .B(n18247), .Z(n17867) );
  NAND U18335 ( .A(n17868), .B(n17867), .Z(n17871) );
  XOR U18336 ( .A(n17870), .B(n17869), .Z(n17872) );
  NANDN U18337 ( .A(n17871), .B(n17872), .Z(n17874) );
  NAND U18338 ( .A(a[22]), .B(b[10]), .Z(n18254) );
  XNOR U18339 ( .A(n17872), .B(n17871), .Z(n18255) );
  NANDN U18340 ( .A(n18254), .B(n18255), .Z(n17873) );
  NAND U18341 ( .A(n17874), .B(n17873), .Z(n17875) );
  OR U18342 ( .A(n17876), .B(n17875), .Z(n17880) );
  XNOR U18343 ( .A(n17876), .B(n17875), .Z(n18258) );
  XOR U18344 ( .A(n17878), .B(n17877), .Z(n18259) );
  NANDN U18345 ( .A(n18258), .B(n18259), .Z(n17879) );
  NAND U18346 ( .A(n17880), .B(n17879), .Z(n17883) );
  XOR U18347 ( .A(n17882), .B(n17881), .Z(n17884) );
  NANDN U18348 ( .A(n17883), .B(n17884), .Z(n17886) );
  NAND U18349 ( .A(a[24]), .B(b[10]), .Z(n18266) );
  XNOR U18350 ( .A(n17884), .B(n17883), .Z(n18267) );
  NANDN U18351 ( .A(n18266), .B(n18267), .Z(n17885) );
  NAND U18352 ( .A(n17886), .B(n17885), .Z(n17887) );
  OR U18353 ( .A(n17888), .B(n17887), .Z(n17892) );
  XNOR U18354 ( .A(n17888), .B(n17887), .Z(n18270) );
  XOR U18355 ( .A(n17890), .B(n17889), .Z(n18271) );
  NANDN U18356 ( .A(n18270), .B(n18271), .Z(n17891) );
  NAND U18357 ( .A(n17892), .B(n17891), .Z(n17895) );
  XOR U18358 ( .A(n17894), .B(n17893), .Z(n17896) );
  NANDN U18359 ( .A(n17895), .B(n17896), .Z(n17898) );
  NAND U18360 ( .A(a[26]), .B(b[10]), .Z(n18278) );
  XNOR U18361 ( .A(n17896), .B(n17895), .Z(n18279) );
  NANDN U18362 ( .A(n18278), .B(n18279), .Z(n17897) );
  NAND U18363 ( .A(n17898), .B(n17897), .Z(n17899) );
  OR U18364 ( .A(n17900), .B(n17899), .Z(n17904) );
  XNOR U18365 ( .A(n17900), .B(n17899), .Z(n18282) );
  XOR U18366 ( .A(n17902), .B(n17901), .Z(n18283) );
  NANDN U18367 ( .A(n18282), .B(n18283), .Z(n17903) );
  NAND U18368 ( .A(n17904), .B(n17903), .Z(n17907) );
  XOR U18369 ( .A(n17906), .B(n17905), .Z(n17908) );
  NANDN U18370 ( .A(n17907), .B(n17908), .Z(n17910) );
  NAND U18371 ( .A(a[28]), .B(b[10]), .Z(n18290) );
  XNOR U18372 ( .A(n17908), .B(n17907), .Z(n18291) );
  NANDN U18373 ( .A(n18290), .B(n18291), .Z(n17909) );
  NAND U18374 ( .A(n17910), .B(n17909), .Z(n17911) );
  OR U18375 ( .A(n17912), .B(n17911), .Z(n17916) );
  XNOR U18376 ( .A(n17912), .B(n17911), .Z(n18294) );
  XOR U18377 ( .A(n17914), .B(n17913), .Z(n18295) );
  NANDN U18378 ( .A(n18294), .B(n18295), .Z(n17915) );
  NAND U18379 ( .A(n17916), .B(n17915), .Z(n17919) );
  XOR U18380 ( .A(n17918), .B(n17917), .Z(n17920) );
  NANDN U18381 ( .A(n17919), .B(n17920), .Z(n17922) );
  NAND U18382 ( .A(a[30]), .B(b[10]), .Z(n18302) );
  XNOR U18383 ( .A(n17920), .B(n17919), .Z(n18303) );
  NANDN U18384 ( .A(n18302), .B(n18303), .Z(n17921) );
  NAND U18385 ( .A(n17922), .B(n17921), .Z(n17923) );
  OR U18386 ( .A(n17924), .B(n17923), .Z(n17928) );
  XNOR U18387 ( .A(n17924), .B(n17923), .Z(n18306) );
  XOR U18388 ( .A(n17926), .B(n17925), .Z(n18307) );
  NANDN U18389 ( .A(n18306), .B(n18307), .Z(n17927) );
  NAND U18390 ( .A(n17928), .B(n17927), .Z(n17931) );
  XOR U18391 ( .A(n17930), .B(n17929), .Z(n17932) );
  NANDN U18392 ( .A(n17931), .B(n17932), .Z(n17934) );
  NAND U18393 ( .A(a[32]), .B(b[10]), .Z(n18314) );
  XNOR U18394 ( .A(n17932), .B(n17931), .Z(n18315) );
  NANDN U18395 ( .A(n18314), .B(n18315), .Z(n17933) );
  NAND U18396 ( .A(n17934), .B(n17933), .Z(n17935) );
  OR U18397 ( .A(n17936), .B(n17935), .Z(n17940) );
  XNOR U18398 ( .A(n17936), .B(n17935), .Z(n18318) );
  XOR U18399 ( .A(n17938), .B(n17937), .Z(n18319) );
  NANDN U18400 ( .A(n18318), .B(n18319), .Z(n17939) );
  NAND U18401 ( .A(n17940), .B(n17939), .Z(n17943) );
  XOR U18402 ( .A(n17942), .B(n17941), .Z(n17944) );
  NANDN U18403 ( .A(n17943), .B(n17944), .Z(n17946) );
  NAND U18404 ( .A(a[34]), .B(b[10]), .Z(n18326) );
  XNOR U18405 ( .A(n17944), .B(n17943), .Z(n18327) );
  NANDN U18406 ( .A(n18326), .B(n18327), .Z(n17945) );
  NAND U18407 ( .A(n17946), .B(n17945), .Z(n17947) );
  OR U18408 ( .A(n17948), .B(n17947), .Z(n17952) );
  XNOR U18409 ( .A(n17948), .B(n17947), .Z(n18330) );
  XOR U18410 ( .A(n17950), .B(n17949), .Z(n18331) );
  NANDN U18411 ( .A(n18330), .B(n18331), .Z(n17951) );
  NAND U18412 ( .A(n17952), .B(n17951), .Z(n17955) );
  XOR U18413 ( .A(n17954), .B(n17953), .Z(n17956) );
  NANDN U18414 ( .A(n17955), .B(n17956), .Z(n17958) );
  NAND U18415 ( .A(a[36]), .B(b[10]), .Z(n18338) );
  XNOR U18416 ( .A(n17956), .B(n17955), .Z(n18339) );
  NANDN U18417 ( .A(n18338), .B(n18339), .Z(n17957) );
  NAND U18418 ( .A(n17958), .B(n17957), .Z(n17959) );
  OR U18419 ( .A(n17960), .B(n17959), .Z(n17964) );
  XNOR U18420 ( .A(n17960), .B(n17959), .Z(n18342) );
  XOR U18421 ( .A(n17962), .B(n17961), .Z(n18343) );
  NANDN U18422 ( .A(n18342), .B(n18343), .Z(n17963) );
  NAND U18423 ( .A(n17964), .B(n17963), .Z(n17967) );
  XOR U18424 ( .A(n17966), .B(n17965), .Z(n17968) );
  NANDN U18425 ( .A(n17967), .B(n17968), .Z(n17970) );
  NAND U18426 ( .A(a[38]), .B(b[10]), .Z(n18350) );
  XNOR U18427 ( .A(n17968), .B(n17967), .Z(n18351) );
  NANDN U18428 ( .A(n18350), .B(n18351), .Z(n17969) );
  NAND U18429 ( .A(n17970), .B(n17969), .Z(n17971) );
  OR U18430 ( .A(n17972), .B(n17971), .Z(n17976) );
  XNOR U18431 ( .A(n17972), .B(n17971), .Z(n18354) );
  XOR U18432 ( .A(n17974), .B(n17973), .Z(n18355) );
  NANDN U18433 ( .A(n18354), .B(n18355), .Z(n17975) );
  NAND U18434 ( .A(n17976), .B(n17975), .Z(n17979) );
  XOR U18435 ( .A(n17978), .B(n17977), .Z(n17980) );
  NANDN U18436 ( .A(n17979), .B(n17980), .Z(n17982) );
  NAND U18437 ( .A(a[40]), .B(b[10]), .Z(n18362) );
  XNOR U18438 ( .A(n17980), .B(n17979), .Z(n18363) );
  NANDN U18439 ( .A(n18362), .B(n18363), .Z(n17981) );
  NAND U18440 ( .A(n17982), .B(n17981), .Z(n17983) );
  OR U18441 ( .A(n17984), .B(n17983), .Z(n17988) );
  XNOR U18442 ( .A(n17984), .B(n17983), .Z(n18366) );
  XOR U18443 ( .A(n17986), .B(n17985), .Z(n18367) );
  NANDN U18444 ( .A(n18366), .B(n18367), .Z(n17987) );
  NAND U18445 ( .A(n17988), .B(n17987), .Z(n17991) );
  XOR U18446 ( .A(n17990), .B(n17989), .Z(n17992) );
  NANDN U18447 ( .A(n17991), .B(n17992), .Z(n17994) );
  NAND U18448 ( .A(a[42]), .B(b[10]), .Z(n18374) );
  XNOR U18449 ( .A(n17992), .B(n17991), .Z(n18375) );
  NANDN U18450 ( .A(n18374), .B(n18375), .Z(n17993) );
  NAND U18451 ( .A(n17994), .B(n17993), .Z(n17995) );
  OR U18452 ( .A(n17996), .B(n17995), .Z(n18000) );
  XNOR U18453 ( .A(n17996), .B(n17995), .Z(n18378) );
  XOR U18454 ( .A(n17998), .B(n17997), .Z(n18379) );
  NANDN U18455 ( .A(n18378), .B(n18379), .Z(n17999) );
  NAND U18456 ( .A(n18000), .B(n17999), .Z(n18003) );
  XOR U18457 ( .A(n18002), .B(n18001), .Z(n18004) );
  NANDN U18458 ( .A(n18003), .B(n18004), .Z(n18006) );
  NAND U18459 ( .A(a[44]), .B(b[10]), .Z(n18386) );
  XNOR U18460 ( .A(n18004), .B(n18003), .Z(n18387) );
  NANDN U18461 ( .A(n18386), .B(n18387), .Z(n18005) );
  NAND U18462 ( .A(n18006), .B(n18005), .Z(n18007) );
  OR U18463 ( .A(n18008), .B(n18007), .Z(n18012) );
  XNOR U18464 ( .A(n18008), .B(n18007), .Z(n18390) );
  XOR U18465 ( .A(n18010), .B(n18009), .Z(n18391) );
  NANDN U18466 ( .A(n18390), .B(n18391), .Z(n18011) );
  NAND U18467 ( .A(n18012), .B(n18011), .Z(n18015) );
  XOR U18468 ( .A(n18014), .B(n18013), .Z(n18016) );
  NANDN U18469 ( .A(n18015), .B(n18016), .Z(n18018) );
  NAND U18470 ( .A(a[46]), .B(b[10]), .Z(n18398) );
  XNOR U18471 ( .A(n18016), .B(n18015), .Z(n18399) );
  NANDN U18472 ( .A(n18398), .B(n18399), .Z(n18017) );
  NAND U18473 ( .A(n18018), .B(n18017), .Z(n18019) );
  OR U18474 ( .A(n18020), .B(n18019), .Z(n18024) );
  XNOR U18475 ( .A(n18020), .B(n18019), .Z(n18402) );
  XOR U18476 ( .A(n18022), .B(n18021), .Z(n18403) );
  NANDN U18477 ( .A(n18402), .B(n18403), .Z(n18023) );
  NAND U18478 ( .A(n18024), .B(n18023), .Z(n18027) );
  XOR U18479 ( .A(n18026), .B(n18025), .Z(n18028) );
  NANDN U18480 ( .A(n18027), .B(n18028), .Z(n18030) );
  NAND U18481 ( .A(a[48]), .B(b[10]), .Z(n18410) );
  XNOR U18482 ( .A(n18028), .B(n18027), .Z(n18411) );
  NANDN U18483 ( .A(n18410), .B(n18411), .Z(n18029) );
  NAND U18484 ( .A(n18030), .B(n18029), .Z(n18031) );
  OR U18485 ( .A(n18032), .B(n18031), .Z(n18036) );
  XNOR U18486 ( .A(n18032), .B(n18031), .Z(n18414) );
  XOR U18487 ( .A(n18034), .B(n18033), .Z(n18415) );
  NANDN U18488 ( .A(n18414), .B(n18415), .Z(n18035) );
  NAND U18489 ( .A(n18036), .B(n18035), .Z(n18039) );
  XOR U18490 ( .A(n18038), .B(n18037), .Z(n18040) );
  NANDN U18491 ( .A(n18039), .B(n18040), .Z(n18042) );
  NAND U18492 ( .A(a[50]), .B(b[10]), .Z(n18422) );
  XNOR U18493 ( .A(n18040), .B(n18039), .Z(n18423) );
  NANDN U18494 ( .A(n18422), .B(n18423), .Z(n18041) );
  NAND U18495 ( .A(n18042), .B(n18041), .Z(n18043) );
  OR U18496 ( .A(n18044), .B(n18043), .Z(n18048) );
  XNOR U18497 ( .A(n18044), .B(n18043), .Z(n18426) );
  XOR U18498 ( .A(n18046), .B(n18045), .Z(n18427) );
  NANDN U18499 ( .A(n18426), .B(n18427), .Z(n18047) );
  NAND U18500 ( .A(n18048), .B(n18047), .Z(n18051) );
  XNOR U18501 ( .A(n18050), .B(n18049), .Z(n18052) );
  OR U18502 ( .A(n18051), .B(n18052), .Z(n18054) );
  XNOR U18503 ( .A(n18052), .B(n18051), .Z(n18433) );
  NAND U18504 ( .A(a[52]), .B(b[10]), .Z(n18432) );
  OR U18505 ( .A(n18433), .B(n18432), .Z(n18053) );
  NAND U18506 ( .A(n18054), .B(n18053), .Z(n18057) );
  ANDN U18507 ( .B(b[10]), .A(n201), .Z(n18058) );
  OR U18508 ( .A(n18057), .B(n18058), .Z(n18060) );
  XOR U18509 ( .A(n18058), .B(n18057), .Z(n18438) );
  NANDN U18510 ( .A(n18439), .B(n18438), .Z(n18059) );
  NAND U18511 ( .A(n18060), .B(n18059), .Z(n18062) );
  AND U18512 ( .A(b[10]), .B(a[54]), .Z(n18061) );
  NANDN U18513 ( .A(n18062), .B(n18061), .Z(n18066) );
  XNOR U18514 ( .A(n18062), .B(n18061), .Z(n18444) );
  NAND U18515 ( .A(n18444), .B(n18445), .Z(n18065) );
  NAND U18516 ( .A(n18066), .B(n18065), .Z(n18068) );
  NANDN U18517 ( .A(n18067), .B(n18068), .Z(n18070) );
  XOR U18518 ( .A(n18068), .B(n18067), .Z(n18451) );
  NAND U18519 ( .A(a[55]), .B(b[10]), .Z(n18450) );
  OR U18520 ( .A(n18451), .B(n18450), .Z(n18069) );
  NAND U18521 ( .A(n18070), .B(n18069), .Z(n18071) );
  NANDN U18522 ( .A(n18072), .B(n18071), .Z(n18076) );
  XNOR U18523 ( .A(n18074), .B(n18073), .Z(n18457) );
  NAND U18524 ( .A(n18456), .B(n18457), .Z(n18075) );
  NAND U18525 ( .A(n18076), .B(n18075), .Z(n18079) );
  OR U18526 ( .A(n18080), .B(n18079), .Z(n18082) );
  XNOR U18527 ( .A(n18078), .B(n18077), .Z(n18463) );
  XOR U18528 ( .A(n18080), .B(n18079), .Z(n18462) );
  NANDN U18529 ( .A(n18463), .B(n18462), .Z(n18081) );
  NAND U18530 ( .A(n18082), .B(n18081), .Z(n18084) );
  NAND U18531 ( .A(a[58]), .B(b[10]), .Z(n18083) );
  OR U18532 ( .A(n18084), .B(n18083), .Z(n18088) );
  XOR U18533 ( .A(n18084), .B(n18083), .Z(n18468) );
  XNOR U18534 ( .A(n18086), .B(n18085), .Z(n18469) );
  NAND U18535 ( .A(n18468), .B(n18469), .Z(n18087) );
  NAND U18536 ( .A(n18088), .B(n18087), .Z(n18091) );
  OR U18537 ( .A(n18092), .B(n18091), .Z(n18094) );
  XNOR U18538 ( .A(n18090), .B(n18089), .Z(n18475) );
  XOR U18539 ( .A(n18092), .B(n18091), .Z(n18474) );
  NANDN U18540 ( .A(n18475), .B(n18474), .Z(n18093) );
  NAND U18541 ( .A(n18094), .B(n18093), .Z(n18096) );
  AND U18542 ( .A(b[10]), .B(a[60]), .Z(n18095) );
  NANDN U18543 ( .A(n18096), .B(n18095), .Z(n18100) );
  XNOR U18544 ( .A(n18096), .B(n18095), .Z(n18122) );
  XOR U18545 ( .A(n18098), .B(n18097), .Z(n18121) );
  NAND U18546 ( .A(n18122), .B(n18121), .Z(n18099) );
  NAND U18547 ( .A(n18100), .B(n18099), .Z(n18101) );
  NAND U18548 ( .A(a[61]), .B(b[10]), .Z(n18102) );
  NANDN U18549 ( .A(n18101), .B(n18102), .Z(n18106) );
  XOR U18550 ( .A(n18102), .B(n18101), .Z(n18484) );
  XOR U18551 ( .A(n18104), .B(n18103), .Z(n18485) );
  NANDN U18552 ( .A(n18484), .B(n18485), .Z(n18105) );
  NAND U18553 ( .A(n18106), .B(n18105), .Z(n18108) );
  AND U18554 ( .A(b[10]), .B(a[62]), .Z(n18107) );
  NANDN U18555 ( .A(n18108), .B(n18107), .Z(n18112) );
  XNOR U18556 ( .A(n18108), .B(n18107), .Z(n18120) );
  XOR U18557 ( .A(n18110), .B(n18109), .Z(n18119) );
  NAND U18558 ( .A(n18120), .B(n18119), .Z(n18111) );
  NAND U18559 ( .A(n18112), .B(n18111), .Z(n18113) );
  ANDN U18560 ( .B(b[10]), .A(n210), .Z(n18114) );
  OR U18561 ( .A(n18113), .B(n18114), .Z(n18118) );
  XNOR U18562 ( .A(n18114), .B(n18113), .Z(n18494) );
  OR U18563 ( .A(n18494), .B(n18495), .Z(n18117) );
  NAND U18564 ( .A(n18118), .B(n18117), .Z(n18496) );
  IV U18565 ( .A(n24127), .Z(n24123) );
  NANDN U18566 ( .A(n24126), .B(n24123), .Z(n18498) );
  XNOR U18567 ( .A(n18120), .B(n18119), .Z(n18490) );
  NAND U18568 ( .A(a[62]), .B(b[9]), .Z(n18486) );
  XNOR U18569 ( .A(n18122), .B(n18121), .Z(n18480) );
  NAND U18570 ( .A(a[60]), .B(b[9]), .Z(n18476) );
  NAND U18571 ( .A(a[58]), .B(b[9]), .Z(n18464) );
  ANDN U18572 ( .B(b[9]), .A(n199), .Z(n18421) );
  ANDN U18573 ( .B(b[9]), .A(n197), .Z(n18409) );
  ANDN U18574 ( .B(b[9]), .A(n195), .Z(n18397) );
  ANDN U18575 ( .B(b[9]), .A(n193), .Z(n18385) );
  ANDN U18576 ( .B(b[9]), .A(n191), .Z(n18373) );
  ANDN U18577 ( .B(b[9]), .A(n189), .Z(n18361) );
  ANDN U18578 ( .B(b[9]), .A(n187), .Z(n18349) );
  ANDN U18579 ( .B(b[9]), .A(n21772), .Z(n18337) );
  ANDN U18580 ( .B(b[9]), .A(n184), .Z(n18325) );
  ANDN U18581 ( .B(b[9]), .A(n21751), .Z(n18313) );
  ANDN U18582 ( .B(b[9]), .A(n21740), .Z(n18301) );
  ANDN U18583 ( .B(b[9]), .A(n21727), .Z(n18289) );
  ANDN U18584 ( .B(b[9]), .A(n21716), .Z(n18277) );
  ANDN U18585 ( .B(b[9]), .A(n21703), .Z(n18265) );
  ANDN U18586 ( .B(b[9]), .A(n21692), .Z(n18253) );
  ANDN U18587 ( .B(b[9]), .A(n21681), .Z(n18241) );
  ANDN U18588 ( .B(b[9]), .A(n21670), .Z(n18229) );
  ANDN U18589 ( .B(b[9]), .A(n174), .Z(n18217) );
  NAND U18590 ( .A(a[16]), .B(b[9]), .Z(n18212) );
  XOR U18591 ( .A(n18124), .B(n18123), .Z(n18213) );
  NANDN U18592 ( .A(n18212), .B(n18213), .Z(n18215) );
  ANDN U18593 ( .B(b[9]), .A(n172), .Z(n18209) );
  ANDN U18594 ( .B(b[9]), .A(n170), .Z(n18197) );
  ANDN U18595 ( .B(b[9]), .A(n21164), .Z(n18185) );
  ANDN U18596 ( .B(b[9]), .A(n21615), .Z(n18171) );
  ANDN U18597 ( .B(b[9]), .A(n166), .Z(n18159) );
  NAND U18598 ( .A(a[6]), .B(b[9]), .Z(n18154) );
  XOR U18599 ( .A(n18126), .B(n18125), .Z(n18155) );
  NANDN U18600 ( .A(n18154), .B(n18155), .Z(n18157) );
  ANDN U18601 ( .B(b[9]), .A(n164), .Z(n18149) );
  ANDN U18602 ( .B(b[9]), .A(n21580), .Z(n18136) );
  NAND U18603 ( .A(b[10]), .B(a[1]), .Z(n18129) );
  AND U18604 ( .A(b[9]), .B(a[0]), .Z(n18894) );
  NANDN U18605 ( .A(n18129), .B(n18894), .Z(n18128) );
  NAND U18606 ( .A(a[2]), .B(b[9]), .Z(n18127) );
  AND U18607 ( .A(n18128), .B(n18127), .Z(n18135) );
  NANDN U18608 ( .A(n18129), .B(a[0]), .Z(n18130) );
  XNOR U18609 ( .A(a[2]), .B(n18130), .Z(n18131) );
  NAND U18610 ( .A(b[9]), .B(n18131), .Z(n18521) );
  AND U18611 ( .A(a[1]), .B(b[10]), .Z(n18132) );
  XOR U18612 ( .A(n18133), .B(n18132), .Z(n18522) );
  OR U18613 ( .A(n18521), .B(n18522), .Z(n18134) );
  NANDN U18614 ( .A(n18135), .B(n18134), .Z(n18137) );
  NANDN U18615 ( .A(n18136), .B(n18137), .Z(n18141) );
  XOR U18616 ( .A(n18137), .B(n18136), .Z(n18526) );
  NANDN U18617 ( .A(n18526), .B(n18525), .Z(n18140) );
  NAND U18618 ( .A(n18141), .B(n18140), .Z(n18145) );
  XOR U18619 ( .A(n18143), .B(n18142), .Z(n18144) );
  NANDN U18620 ( .A(n18145), .B(n18144), .Z(n18147) );
  NAND U18621 ( .A(a[4]), .B(b[9]), .Z(n18533) );
  NANDN U18622 ( .A(n18533), .B(n18534), .Z(n18146) );
  NAND U18623 ( .A(n18147), .B(n18146), .Z(n18148) );
  OR U18624 ( .A(n18149), .B(n18148), .Z(n18153) );
  XNOR U18625 ( .A(n18149), .B(n18148), .Z(n18508) );
  XOR U18626 ( .A(n18151), .B(n18150), .Z(n18509) );
  NANDN U18627 ( .A(n18508), .B(n18509), .Z(n18152) );
  NAND U18628 ( .A(n18153), .B(n18152), .Z(n18543) );
  XNOR U18629 ( .A(n18155), .B(n18154), .Z(n18544) );
  NANDN U18630 ( .A(n18543), .B(n18544), .Z(n18156) );
  NAND U18631 ( .A(n18157), .B(n18156), .Z(n18158) );
  OR U18632 ( .A(n18159), .B(n18158), .Z(n18163) );
  XNOR U18633 ( .A(n18159), .B(n18158), .Z(n18547) );
  XOR U18634 ( .A(n18161), .B(n18160), .Z(n18548) );
  NANDN U18635 ( .A(n18547), .B(n18548), .Z(n18162) );
  NAND U18636 ( .A(n18163), .B(n18162), .Z(n18166) );
  XOR U18637 ( .A(n18165), .B(n18164), .Z(n18167) );
  NANDN U18638 ( .A(n18166), .B(n18167), .Z(n18169) );
  NAND U18639 ( .A(a[8]), .B(b[9]), .Z(n18555) );
  XNOR U18640 ( .A(n18167), .B(n18166), .Z(n18556) );
  NANDN U18641 ( .A(n18555), .B(n18556), .Z(n18168) );
  NAND U18642 ( .A(n18169), .B(n18168), .Z(n18170) );
  OR U18643 ( .A(n18171), .B(n18170), .Z(n18175) );
  XNOR U18644 ( .A(n18171), .B(n18170), .Z(n18559) );
  XOR U18645 ( .A(n18173), .B(n18172), .Z(n18560) );
  NANDN U18646 ( .A(n18559), .B(n18560), .Z(n18174) );
  NAND U18647 ( .A(n18175), .B(n18174), .Z(n18178) );
  XOR U18648 ( .A(n18177), .B(n18176), .Z(n18179) );
  NANDN U18649 ( .A(n18178), .B(n18179), .Z(n18181) );
  NAND U18650 ( .A(a[10]), .B(b[9]), .Z(n18567) );
  XNOR U18651 ( .A(n18179), .B(n18178), .Z(n18568) );
  NANDN U18652 ( .A(n18567), .B(n18568), .Z(n18180) );
  NAND U18653 ( .A(n18181), .B(n18180), .Z(n18184) );
  OR U18654 ( .A(n18185), .B(n18184), .Z(n18187) );
  XOR U18655 ( .A(n18183), .B(n18182), .Z(n18572) );
  XOR U18656 ( .A(n18185), .B(n18184), .Z(n18571) );
  NANDN U18657 ( .A(n18572), .B(n18571), .Z(n18186) );
  NAND U18658 ( .A(n18187), .B(n18186), .Z(n18190) );
  XOR U18659 ( .A(n18189), .B(n18188), .Z(n18191) );
  NANDN U18660 ( .A(n18190), .B(n18191), .Z(n18193) );
  NAND U18661 ( .A(a[12]), .B(b[9]), .Z(n18579) );
  XNOR U18662 ( .A(n18191), .B(n18190), .Z(n18580) );
  NANDN U18663 ( .A(n18579), .B(n18580), .Z(n18192) );
  NAND U18664 ( .A(n18193), .B(n18192), .Z(n18196) );
  OR U18665 ( .A(n18197), .B(n18196), .Z(n18199) );
  XOR U18666 ( .A(n18195), .B(n18194), .Z(n18507) );
  XOR U18667 ( .A(n18197), .B(n18196), .Z(n18506) );
  NANDN U18668 ( .A(n18507), .B(n18506), .Z(n18198) );
  NAND U18669 ( .A(n18199), .B(n18198), .Z(n18202) );
  XOR U18670 ( .A(n18201), .B(n18200), .Z(n18203) );
  NANDN U18671 ( .A(n18202), .B(n18203), .Z(n18205) );
  NAND U18672 ( .A(a[14]), .B(b[9]), .Z(n18589) );
  XNOR U18673 ( .A(n18203), .B(n18202), .Z(n18590) );
  NANDN U18674 ( .A(n18589), .B(n18590), .Z(n18204) );
  NAND U18675 ( .A(n18205), .B(n18204), .Z(n18208) );
  OR U18676 ( .A(n18209), .B(n18208), .Z(n18211) );
  XOR U18677 ( .A(n18207), .B(n18206), .Z(n18505) );
  XOR U18678 ( .A(n18209), .B(n18208), .Z(n18504) );
  NAND U18679 ( .A(n18505), .B(n18504), .Z(n18210) );
  NAND U18680 ( .A(n18211), .B(n18210), .Z(n18597) );
  XNOR U18681 ( .A(n18213), .B(n18212), .Z(n18598) );
  NANDN U18682 ( .A(n18597), .B(n18598), .Z(n18214) );
  NAND U18683 ( .A(n18215), .B(n18214), .Z(n18216) );
  OR U18684 ( .A(n18217), .B(n18216), .Z(n18221) );
  XNOR U18685 ( .A(n18217), .B(n18216), .Z(n18603) );
  XOR U18686 ( .A(n18219), .B(n18218), .Z(n18604) );
  NANDN U18687 ( .A(n18603), .B(n18604), .Z(n18220) );
  NAND U18688 ( .A(n18221), .B(n18220), .Z(n18225) );
  XOR U18689 ( .A(n18223), .B(n18222), .Z(n18224) );
  NANDN U18690 ( .A(n18225), .B(n18224), .Z(n18227) );
  NAND U18691 ( .A(a[18]), .B(b[9]), .Z(n18609) );
  NANDN U18692 ( .A(n18609), .B(n18610), .Z(n18226) );
  NAND U18693 ( .A(n18227), .B(n18226), .Z(n18228) );
  OR U18694 ( .A(n18229), .B(n18228), .Z(n18233) );
  XNOR U18695 ( .A(n18229), .B(n18228), .Z(n18615) );
  XOR U18696 ( .A(n18231), .B(n18230), .Z(n18616) );
  NANDN U18697 ( .A(n18615), .B(n18616), .Z(n18232) );
  NAND U18698 ( .A(n18233), .B(n18232), .Z(n18236) );
  XOR U18699 ( .A(n18235), .B(n18234), .Z(n18237) );
  NANDN U18700 ( .A(n18236), .B(n18237), .Z(n18239) );
  NAND U18701 ( .A(a[20]), .B(b[9]), .Z(n18623) );
  XNOR U18702 ( .A(n18237), .B(n18236), .Z(n18624) );
  NANDN U18703 ( .A(n18623), .B(n18624), .Z(n18238) );
  NAND U18704 ( .A(n18239), .B(n18238), .Z(n18240) );
  OR U18705 ( .A(n18241), .B(n18240), .Z(n18245) );
  XNOR U18706 ( .A(n18241), .B(n18240), .Z(n18627) );
  XOR U18707 ( .A(n18243), .B(n18242), .Z(n18628) );
  NANDN U18708 ( .A(n18627), .B(n18628), .Z(n18244) );
  NAND U18709 ( .A(n18245), .B(n18244), .Z(n18248) );
  XOR U18710 ( .A(n18247), .B(n18246), .Z(n18249) );
  NANDN U18711 ( .A(n18248), .B(n18249), .Z(n18251) );
  NAND U18712 ( .A(a[22]), .B(b[9]), .Z(n18635) );
  XNOR U18713 ( .A(n18249), .B(n18248), .Z(n18636) );
  NANDN U18714 ( .A(n18635), .B(n18636), .Z(n18250) );
  NAND U18715 ( .A(n18251), .B(n18250), .Z(n18252) );
  OR U18716 ( .A(n18253), .B(n18252), .Z(n18257) );
  XNOR U18717 ( .A(n18253), .B(n18252), .Z(n18639) );
  XOR U18718 ( .A(n18255), .B(n18254), .Z(n18640) );
  NANDN U18719 ( .A(n18639), .B(n18640), .Z(n18256) );
  NAND U18720 ( .A(n18257), .B(n18256), .Z(n18260) );
  XOR U18721 ( .A(n18259), .B(n18258), .Z(n18261) );
  NANDN U18722 ( .A(n18260), .B(n18261), .Z(n18263) );
  NAND U18723 ( .A(a[24]), .B(b[9]), .Z(n18647) );
  XNOR U18724 ( .A(n18261), .B(n18260), .Z(n18648) );
  NANDN U18725 ( .A(n18647), .B(n18648), .Z(n18262) );
  NAND U18726 ( .A(n18263), .B(n18262), .Z(n18264) );
  OR U18727 ( .A(n18265), .B(n18264), .Z(n18269) );
  XNOR U18728 ( .A(n18265), .B(n18264), .Z(n18651) );
  XOR U18729 ( .A(n18267), .B(n18266), .Z(n18652) );
  NANDN U18730 ( .A(n18651), .B(n18652), .Z(n18268) );
  NAND U18731 ( .A(n18269), .B(n18268), .Z(n18272) );
  XOR U18732 ( .A(n18271), .B(n18270), .Z(n18273) );
  NANDN U18733 ( .A(n18272), .B(n18273), .Z(n18275) );
  NAND U18734 ( .A(a[26]), .B(b[9]), .Z(n18659) );
  XNOR U18735 ( .A(n18273), .B(n18272), .Z(n18660) );
  NANDN U18736 ( .A(n18659), .B(n18660), .Z(n18274) );
  NAND U18737 ( .A(n18275), .B(n18274), .Z(n18276) );
  OR U18738 ( .A(n18277), .B(n18276), .Z(n18281) );
  XNOR U18739 ( .A(n18277), .B(n18276), .Z(n18663) );
  XOR U18740 ( .A(n18279), .B(n18278), .Z(n18664) );
  NANDN U18741 ( .A(n18663), .B(n18664), .Z(n18280) );
  NAND U18742 ( .A(n18281), .B(n18280), .Z(n18284) );
  XOR U18743 ( .A(n18283), .B(n18282), .Z(n18285) );
  NANDN U18744 ( .A(n18284), .B(n18285), .Z(n18287) );
  NAND U18745 ( .A(a[28]), .B(b[9]), .Z(n18671) );
  XNOR U18746 ( .A(n18285), .B(n18284), .Z(n18672) );
  NANDN U18747 ( .A(n18671), .B(n18672), .Z(n18286) );
  NAND U18748 ( .A(n18287), .B(n18286), .Z(n18288) );
  OR U18749 ( .A(n18289), .B(n18288), .Z(n18293) );
  XNOR U18750 ( .A(n18289), .B(n18288), .Z(n18675) );
  XOR U18751 ( .A(n18291), .B(n18290), .Z(n18676) );
  NANDN U18752 ( .A(n18675), .B(n18676), .Z(n18292) );
  NAND U18753 ( .A(n18293), .B(n18292), .Z(n18296) );
  XOR U18754 ( .A(n18295), .B(n18294), .Z(n18297) );
  NANDN U18755 ( .A(n18296), .B(n18297), .Z(n18299) );
  NAND U18756 ( .A(a[30]), .B(b[9]), .Z(n18683) );
  XNOR U18757 ( .A(n18297), .B(n18296), .Z(n18684) );
  NANDN U18758 ( .A(n18683), .B(n18684), .Z(n18298) );
  NAND U18759 ( .A(n18299), .B(n18298), .Z(n18300) );
  OR U18760 ( .A(n18301), .B(n18300), .Z(n18305) );
  XNOR U18761 ( .A(n18301), .B(n18300), .Z(n18687) );
  XOR U18762 ( .A(n18303), .B(n18302), .Z(n18688) );
  NANDN U18763 ( .A(n18687), .B(n18688), .Z(n18304) );
  NAND U18764 ( .A(n18305), .B(n18304), .Z(n18308) );
  XOR U18765 ( .A(n18307), .B(n18306), .Z(n18309) );
  NANDN U18766 ( .A(n18308), .B(n18309), .Z(n18311) );
  NAND U18767 ( .A(a[32]), .B(b[9]), .Z(n18695) );
  XNOR U18768 ( .A(n18309), .B(n18308), .Z(n18696) );
  NANDN U18769 ( .A(n18695), .B(n18696), .Z(n18310) );
  NAND U18770 ( .A(n18311), .B(n18310), .Z(n18312) );
  OR U18771 ( .A(n18313), .B(n18312), .Z(n18317) );
  XNOR U18772 ( .A(n18313), .B(n18312), .Z(n18699) );
  XOR U18773 ( .A(n18315), .B(n18314), .Z(n18700) );
  NANDN U18774 ( .A(n18699), .B(n18700), .Z(n18316) );
  NAND U18775 ( .A(n18317), .B(n18316), .Z(n18320) );
  XOR U18776 ( .A(n18319), .B(n18318), .Z(n18321) );
  NANDN U18777 ( .A(n18320), .B(n18321), .Z(n18323) );
  NAND U18778 ( .A(a[34]), .B(b[9]), .Z(n18707) );
  XNOR U18779 ( .A(n18321), .B(n18320), .Z(n18708) );
  NANDN U18780 ( .A(n18707), .B(n18708), .Z(n18322) );
  NAND U18781 ( .A(n18323), .B(n18322), .Z(n18324) );
  OR U18782 ( .A(n18325), .B(n18324), .Z(n18329) );
  XNOR U18783 ( .A(n18325), .B(n18324), .Z(n18711) );
  XOR U18784 ( .A(n18327), .B(n18326), .Z(n18712) );
  NANDN U18785 ( .A(n18711), .B(n18712), .Z(n18328) );
  NAND U18786 ( .A(n18329), .B(n18328), .Z(n18332) );
  XOR U18787 ( .A(n18331), .B(n18330), .Z(n18333) );
  NANDN U18788 ( .A(n18332), .B(n18333), .Z(n18335) );
  NAND U18789 ( .A(a[36]), .B(b[9]), .Z(n18719) );
  XNOR U18790 ( .A(n18333), .B(n18332), .Z(n18720) );
  NANDN U18791 ( .A(n18719), .B(n18720), .Z(n18334) );
  NAND U18792 ( .A(n18335), .B(n18334), .Z(n18336) );
  OR U18793 ( .A(n18337), .B(n18336), .Z(n18341) );
  XNOR U18794 ( .A(n18337), .B(n18336), .Z(n18723) );
  XOR U18795 ( .A(n18339), .B(n18338), .Z(n18724) );
  NANDN U18796 ( .A(n18723), .B(n18724), .Z(n18340) );
  NAND U18797 ( .A(n18341), .B(n18340), .Z(n18344) );
  XOR U18798 ( .A(n18343), .B(n18342), .Z(n18345) );
  NANDN U18799 ( .A(n18344), .B(n18345), .Z(n18347) );
  NAND U18800 ( .A(a[38]), .B(b[9]), .Z(n18731) );
  XNOR U18801 ( .A(n18345), .B(n18344), .Z(n18732) );
  NANDN U18802 ( .A(n18731), .B(n18732), .Z(n18346) );
  NAND U18803 ( .A(n18347), .B(n18346), .Z(n18348) );
  OR U18804 ( .A(n18349), .B(n18348), .Z(n18353) );
  XNOR U18805 ( .A(n18349), .B(n18348), .Z(n18735) );
  XOR U18806 ( .A(n18351), .B(n18350), .Z(n18736) );
  NANDN U18807 ( .A(n18735), .B(n18736), .Z(n18352) );
  NAND U18808 ( .A(n18353), .B(n18352), .Z(n18356) );
  XOR U18809 ( .A(n18355), .B(n18354), .Z(n18357) );
  NANDN U18810 ( .A(n18356), .B(n18357), .Z(n18359) );
  NAND U18811 ( .A(a[40]), .B(b[9]), .Z(n18743) );
  XNOR U18812 ( .A(n18357), .B(n18356), .Z(n18744) );
  NANDN U18813 ( .A(n18743), .B(n18744), .Z(n18358) );
  NAND U18814 ( .A(n18359), .B(n18358), .Z(n18360) );
  OR U18815 ( .A(n18361), .B(n18360), .Z(n18365) );
  XNOR U18816 ( .A(n18361), .B(n18360), .Z(n18747) );
  XOR U18817 ( .A(n18363), .B(n18362), .Z(n18748) );
  NANDN U18818 ( .A(n18747), .B(n18748), .Z(n18364) );
  NAND U18819 ( .A(n18365), .B(n18364), .Z(n18368) );
  XOR U18820 ( .A(n18367), .B(n18366), .Z(n18369) );
  NANDN U18821 ( .A(n18368), .B(n18369), .Z(n18371) );
  NAND U18822 ( .A(a[42]), .B(b[9]), .Z(n18755) );
  XNOR U18823 ( .A(n18369), .B(n18368), .Z(n18756) );
  NANDN U18824 ( .A(n18755), .B(n18756), .Z(n18370) );
  NAND U18825 ( .A(n18371), .B(n18370), .Z(n18372) );
  OR U18826 ( .A(n18373), .B(n18372), .Z(n18377) );
  XNOR U18827 ( .A(n18373), .B(n18372), .Z(n18759) );
  XOR U18828 ( .A(n18375), .B(n18374), .Z(n18760) );
  NANDN U18829 ( .A(n18759), .B(n18760), .Z(n18376) );
  NAND U18830 ( .A(n18377), .B(n18376), .Z(n18380) );
  XOR U18831 ( .A(n18379), .B(n18378), .Z(n18381) );
  NANDN U18832 ( .A(n18380), .B(n18381), .Z(n18383) );
  NAND U18833 ( .A(a[44]), .B(b[9]), .Z(n18767) );
  XNOR U18834 ( .A(n18381), .B(n18380), .Z(n18768) );
  NANDN U18835 ( .A(n18767), .B(n18768), .Z(n18382) );
  NAND U18836 ( .A(n18383), .B(n18382), .Z(n18384) );
  OR U18837 ( .A(n18385), .B(n18384), .Z(n18389) );
  XNOR U18838 ( .A(n18385), .B(n18384), .Z(n18771) );
  XOR U18839 ( .A(n18387), .B(n18386), .Z(n18772) );
  NANDN U18840 ( .A(n18771), .B(n18772), .Z(n18388) );
  NAND U18841 ( .A(n18389), .B(n18388), .Z(n18392) );
  XOR U18842 ( .A(n18391), .B(n18390), .Z(n18393) );
  NANDN U18843 ( .A(n18392), .B(n18393), .Z(n18395) );
  NAND U18844 ( .A(a[46]), .B(b[9]), .Z(n18779) );
  XNOR U18845 ( .A(n18393), .B(n18392), .Z(n18780) );
  NANDN U18846 ( .A(n18779), .B(n18780), .Z(n18394) );
  NAND U18847 ( .A(n18395), .B(n18394), .Z(n18396) );
  OR U18848 ( .A(n18397), .B(n18396), .Z(n18401) );
  XNOR U18849 ( .A(n18397), .B(n18396), .Z(n18783) );
  XOR U18850 ( .A(n18399), .B(n18398), .Z(n18784) );
  NANDN U18851 ( .A(n18783), .B(n18784), .Z(n18400) );
  NAND U18852 ( .A(n18401), .B(n18400), .Z(n18404) );
  XOR U18853 ( .A(n18403), .B(n18402), .Z(n18405) );
  NANDN U18854 ( .A(n18404), .B(n18405), .Z(n18407) );
  NAND U18855 ( .A(a[48]), .B(b[9]), .Z(n18791) );
  XNOR U18856 ( .A(n18405), .B(n18404), .Z(n18792) );
  NANDN U18857 ( .A(n18791), .B(n18792), .Z(n18406) );
  NAND U18858 ( .A(n18407), .B(n18406), .Z(n18408) );
  OR U18859 ( .A(n18409), .B(n18408), .Z(n18413) );
  XNOR U18860 ( .A(n18409), .B(n18408), .Z(n18795) );
  XOR U18861 ( .A(n18411), .B(n18410), .Z(n18796) );
  NANDN U18862 ( .A(n18795), .B(n18796), .Z(n18412) );
  NAND U18863 ( .A(n18413), .B(n18412), .Z(n18416) );
  XOR U18864 ( .A(n18415), .B(n18414), .Z(n18417) );
  NANDN U18865 ( .A(n18416), .B(n18417), .Z(n18419) );
  NAND U18866 ( .A(a[50]), .B(b[9]), .Z(n18803) );
  XNOR U18867 ( .A(n18417), .B(n18416), .Z(n18804) );
  NANDN U18868 ( .A(n18803), .B(n18804), .Z(n18418) );
  NAND U18869 ( .A(n18419), .B(n18418), .Z(n18420) );
  OR U18870 ( .A(n18421), .B(n18420), .Z(n18425) );
  XNOR U18871 ( .A(n18421), .B(n18420), .Z(n18807) );
  XOR U18872 ( .A(n18423), .B(n18422), .Z(n18808) );
  NANDN U18873 ( .A(n18807), .B(n18808), .Z(n18424) );
  NAND U18874 ( .A(n18425), .B(n18424), .Z(n18428) );
  XOR U18875 ( .A(n18427), .B(n18426), .Z(n18429) );
  NANDN U18876 ( .A(n18428), .B(n18429), .Z(n18431) );
  NAND U18877 ( .A(a[52]), .B(b[9]), .Z(n18815) );
  XNOR U18878 ( .A(n18429), .B(n18428), .Z(n18816) );
  NANDN U18879 ( .A(n18815), .B(n18816), .Z(n18430) );
  NAND U18880 ( .A(n18431), .B(n18430), .Z(n18434) );
  ANDN U18881 ( .B(b[9]), .A(n201), .Z(n18435) );
  OR U18882 ( .A(n18434), .B(n18435), .Z(n18437) );
  XOR U18883 ( .A(n18433), .B(n18432), .Z(n18820) );
  XOR U18884 ( .A(n18435), .B(n18434), .Z(n18819) );
  NANDN U18885 ( .A(n18820), .B(n18819), .Z(n18436) );
  NAND U18886 ( .A(n18437), .B(n18436), .Z(n18440) );
  XNOR U18887 ( .A(n18439), .B(n18438), .Z(n18441) );
  OR U18888 ( .A(n18440), .B(n18441), .Z(n18443) );
  XNOR U18889 ( .A(n18441), .B(n18440), .Z(n18826) );
  NAND U18890 ( .A(a[54]), .B(b[9]), .Z(n18825) );
  OR U18891 ( .A(n18826), .B(n18825), .Z(n18442) );
  NAND U18892 ( .A(n18443), .B(n18442), .Z(n18446) );
  ANDN U18893 ( .B(b[9]), .A(n203), .Z(n18447) );
  OR U18894 ( .A(n18446), .B(n18447), .Z(n18449) );
  XOR U18895 ( .A(n18447), .B(n18446), .Z(n18833) );
  NANDN U18896 ( .A(n18834), .B(n18833), .Z(n18448) );
  NAND U18897 ( .A(n18449), .B(n18448), .Z(n18453) );
  NAND U18898 ( .A(a[56]), .B(b[9]), .Z(n18452) );
  OR U18899 ( .A(n18453), .B(n18452), .Z(n18455) );
  XOR U18900 ( .A(n18451), .B(n18450), .Z(n18837) );
  XOR U18901 ( .A(n18453), .B(n18452), .Z(n18838) );
  NAND U18902 ( .A(n18837), .B(n18838), .Z(n18454) );
  NAND U18903 ( .A(n18455), .B(n18454), .Z(n18459) );
  NAND U18904 ( .A(n18459), .B(n18458), .Z(n18461) );
  XNOR U18905 ( .A(n18459), .B(n18458), .Z(n18844) );
  NAND U18906 ( .A(a[57]), .B(b[9]), .Z(n18843) );
  OR U18907 ( .A(n18844), .B(n18843), .Z(n18460) );
  NAND U18908 ( .A(n18461), .B(n18460), .Z(n18465) );
  NANDN U18909 ( .A(n18464), .B(n18465), .Z(n18467) );
  XNOR U18910 ( .A(n18463), .B(n18462), .Z(n18850) );
  XNOR U18911 ( .A(n18465), .B(n18464), .Z(n18849) );
  NANDN U18912 ( .A(n18850), .B(n18849), .Z(n18466) );
  NAND U18913 ( .A(n18467), .B(n18466), .Z(n18471) );
  NAND U18914 ( .A(n18471), .B(n18470), .Z(n18473) );
  XNOR U18915 ( .A(n18471), .B(n18470), .Z(n18856) );
  NAND U18916 ( .A(a[59]), .B(b[9]), .Z(n18855) );
  OR U18917 ( .A(n18856), .B(n18855), .Z(n18472) );
  NAND U18918 ( .A(n18473), .B(n18472), .Z(n18477) );
  NANDN U18919 ( .A(n18476), .B(n18477), .Z(n18479) );
  XNOR U18920 ( .A(n18475), .B(n18474), .Z(n18862) );
  XNOR U18921 ( .A(n18477), .B(n18476), .Z(n18861) );
  NANDN U18922 ( .A(n18862), .B(n18861), .Z(n18478) );
  NAND U18923 ( .A(n18479), .B(n18478), .Z(n18481) );
  NANDN U18924 ( .A(n18480), .B(n18481), .Z(n18483) );
  NAND U18925 ( .A(a[61]), .B(b[9]), .Z(n18867) );
  XNOR U18926 ( .A(n18481), .B(n18480), .Z(n18868) );
  NANDN U18927 ( .A(n18867), .B(n18868), .Z(n18482) );
  NAND U18928 ( .A(n18483), .B(n18482), .Z(n18487) );
  NANDN U18929 ( .A(n18486), .B(n18487), .Z(n18489) );
  XNOR U18930 ( .A(n18485), .B(n18484), .Z(n18874) );
  XNOR U18931 ( .A(n18487), .B(n18486), .Z(n18873) );
  NANDN U18932 ( .A(n18874), .B(n18873), .Z(n18488) );
  AND U18933 ( .A(n18489), .B(n18488), .Z(n18491) );
  OR U18934 ( .A(n18490), .B(n18491), .Z(n18493) );
  XNOR U18935 ( .A(n18491), .B(n18490), .Z(n18503) );
  AND U18936 ( .A(b[9]), .B(a[63]), .Z(n18502) );
  NANDN U18937 ( .A(n18503), .B(n18502), .Z(n18492) );
  AND U18938 ( .A(n18493), .B(n18492), .Z(n18879) );
  XNOR U18939 ( .A(n18495), .B(n18494), .Z(n18880) );
  NANDN U18940 ( .A(n18879), .B(n18880), .Z(n24117) );
  XNOR U18941 ( .A(n18497), .B(n18496), .Z(n24119) );
  NAND U18942 ( .A(n18498), .B(n24122), .Z(n24129) );
  NOR U18943 ( .A(n21942), .B(n21941), .Z(n24133) );
  IV U18944 ( .A(n24133), .Z(n21939) );
  XNOR U18945 ( .A(n18500), .B(n18499), .Z(n24132) );
  NAND U18946 ( .A(n21939), .B(n24132), .Z(n18501) );
  NANDN U18947 ( .A(n24129), .B(n18501), .Z(n21938) );
  XOR U18948 ( .A(n18503), .B(n18502), .Z(n18884) );
  NAND U18949 ( .A(a[58]), .B(b[8]), .Z(n18845) );
  ANDN U18950 ( .B(b[8]), .A(n201), .Z(n18814) );
  ANDN U18951 ( .B(b[8]), .A(n199), .Z(n18802) );
  ANDN U18952 ( .B(b[8]), .A(n197), .Z(n18790) );
  ANDN U18953 ( .B(b[8]), .A(n195), .Z(n18778) );
  ANDN U18954 ( .B(b[8]), .A(n193), .Z(n18766) );
  ANDN U18955 ( .B(b[8]), .A(n191), .Z(n18754) );
  ANDN U18956 ( .B(b[8]), .A(n189), .Z(n18742) );
  ANDN U18957 ( .B(b[8]), .A(n187), .Z(n18730) );
  ANDN U18958 ( .B(b[8]), .A(n21772), .Z(n18718) );
  ANDN U18959 ( .B(b[8]), .A(n184), .Z(n18706) );
  ANDN U18960 ( .B(b[8]), .A(n21751), .Z(n18694) );
  ANDN U18961 ( .B(b[8]), .A(n21740), .Z(n18682) );
  ANDN U18962 ( .B(b[8]), .A(n21727), .Z(n18670) );
  ANDN U18963 ( .B(b[8]), .A(n21716), .Z(n18658) );
  ANDN U18964 ( .B(b[8]), .A(n21703), .Z(n18646) );
  ANDN U18965 ( .B(b[8]), .A(n21692), .Z(n18634) );
  ANDN U18966 ( .B(b[8]), .A(n21681), .Z(n18622) );
  ANDN U18967 ( .B(b[8]), .A(n21670), .Z(n18612) );
  ANDN U18968 ( .B(b[8]), .A(n174), .Z(n18600) );
  XNOR U18969 ( .A(n18505), .B(n18504), .Z(n18594) );
  ANDN U18970 ( .B(b[8]), .A(n172), .Z(n18588) );
  XNOR U18971 ( .A(n18507), .B(n18506), .Z(n18584) );
  NAND U18972 ( .A(a[13]), .B(b[8]), .Z(n18578) );
  ANDN U18973 ( .B(b[8]), .A(n21164), .Z(n18566) );
  ANDN U18974 ( .B(b[8]), .A(n21615), .Z(n18554) );
  ANDN U18975 ( .B(b[8]), .A(n166), .Z(n18542) );
  NAND U18976 ( .A(a[6]), .B(b[8]), .Z(n18537) );
  XOR U18977 ( .A(n18509), .B(n18508), .Z(n18538) );
  NANDN U18978 ( .A(n18537), .B(n18538), .Z(n18540) );
  ANDN U18979 ( .B(b[8]), .A(n164), .Z(n18532) );
  ANDN U18980 ( .B(b[8]), .A(n21580), .Z(n18519) );
  NAND U18981 ( .A(b[9]), .B(a[1]), .Z(n18514) );
  NANDN U18982 ( .A(n18514), .B(a[0]), .Z(n18510) );
  XNOR U18983 ( .A(a[2]), .B(n18510), .Z(n18511) );
  NAND U18984 ( .A(b[8]), .B(n18511), .Z(n18902) );
  AND U18985 ( .A(a[1]), .B(b[9]), .Z(n18512) );
  XOR U18986 ( .A(n18513), .B(n18512), .Z(n18903) );
  OR U18987 ( .A(n18902), .B(n18903), .Z(n18518) );
  AND U18988 ( .A(b[8]), .B(a[0]), .Z(n19269) );
  NANDN U18989 ( .A(n18514), .B(n19269), .Z(n18516) );
  NAND U18990 ( .A(a[2]), .B(b[8]), .Z(n18515) );
  AND U18991 ( .A(n18516), .B(n18515), .Z(n18517) );
  ANDN U18992 ( .B(n18518), .A(n18517), .Z(n18520) );
  OR U18993 ( .A(n18519), .B(n18520), .Z(n18524) );
  XNOR U18994 ( .A(n18520), .B(n18519), .Z(n18907) );
  XNOR U18995 ( .A(n18522), .B(n18521), .Z(n18906) );
  OR U18996 ( .A(n18907), .B(n18906), .Z(n18523) );
  NAND U18997 ( .A(n18524), .B(n18523), .Z(n18528) );
  XOR U18998 ( .A(n18526), .B(n18525), .Z(n18527) );
  NANDN U18999 ( .A(n18528), .B(n18527), .Z(n18530) );
  NAND U19000 ( .A(a[4]), .B(b[8]), .Z(n18914) );
  NANDN U19001 ( .A(n18914), .B(n18915), .Z(n18529) );
  NAND U19002 ( .A(n18530), .B(n18529), .Z(n18531) );
  OR U19003 ( .A(n18532), .B(n18531), .Z(n18536) );
  XNOR U19004 ( .A(n18532), .B(n18531), .Z(n18889) );
  XOR U19005 ( .A(n18534), .B(n18533), .Z(n18890) );
  NANDN U19006 ( .A(n18889), .B(n18890), .Z(n18535) );
  NAND U19007 ( .A(n18536), .B(n18535), .Z(n18924) );
  XNOR U19008 ( .A(n18538), .B(n18537), .Z(n18925) );
  NANDN U19009 ( .A(n18924), .B(n18925), .Z(n18539) );
  NAND U19010 ( .A(n18540), .B(n18539), .Z(n18541) );
  OR U19011 ( .A(n18542), .B(n18541), .Z(n18546) );
  XNOR U19012 ( .A(n18542), .B(n18541), .Z(n18928) );
  XOR U19013 ( .A(n18544), .B(n18543), .Z(n18929) );
  NANDN U19014 ( .A(n18928), .B(n18929), .Z(n18545) );
  NAND U19015 ( .A(n18546), .B(n18545), .Z(n18549) );
  XOR U19016 ( .A(n18548), .B(n18547), .Z(n18550) );
  NANDN U19017 ( .A(n18549), .B(n18550), .Z(n18552) );
  NAND U19018 ( .A(a[8]), .B(b[8]), .Z(n18936) );
  XNOR U19019 ( .A(n18550), .B(n18549), .Z(n18937) );
  NANDN U19020 ( .A(n18936), .B(n18937), .Z(n18551) );
  NAND U19021 ( .A(n18552), .B(n18551), .Z(n18553) );
  OR U19022 ( .A(n18554), .B(n18553), .Z(n18558) );
  XNOR U19023 ( .A(n18554), .B(n18553), .Z(n18940) );
  XOR U19024 ( .A(n18556), .B(n18555), .Z(n18941) );
  NANDN U19025 ( .A(n18940), .B(n18941), .Z(n18557) );
  NAND U19026 ( .A(n18558), .B(n18557), .Z(n18561) );
  XOR U19027 ( .A(n18560), .B(n18559), .Z(n18562) );
  NANDN U19028 ( .A(n18561), .B(n18562), .Z(n18564) );
  NAND U19029 ( .A(a[10]), .B(b[8]), .Z(n18948) );
  XNOR U19030 ( .A(n18562), .B(n18561), .Z(n18949) );
  NANDN U19031 ( .A(n18948), .B(n18949), .Z(n18563) );
  NAND U19032 ( .A(n18564), .B(n18563), .Z(n18565) );
  OR U19033 ( .A(n18566), .B(n18565), .Z(n18570) );
  XNOR U19034 ( .A(n18566), .B(n18565), .Z(n18952) );
  XOR U19035 ( .A(n18568), .B(n18567), .Z(n18953) );
  NANDN U19036 ( .A(n18952), .B(n18953), .Z(n18569) );
  NAND U19037 ( .A(n18570), .B(n18569), .Z(n18573) );
  XNOR U19038 ( .A(n18572), .B(n18571), .Z(n18574) );
  OR U19039 ( .A(n18573), .B(n18574), .Z(n18576) );
  NAND U19040 ( .A(a[12]), .B(b[8]), .Z(n18960) );
  XOR U19041 ( .A(n18574), .B(n18573), .Z(n18961) );
  NANDN U19042 ( .A(n18960), .B(n18961), .Z(n18575) );
  NAND U19043 ( .A(n18576), .B(n18575), .Z(n18577) );
  NANDN U19044 ( .A(n18578), .B(n18577), .Z(n18582) );
  XNOR U19045 ( .A(n18580), .B(n18579), .Z(n18967) );
  NAND U19046 ( .A(n18966), .B(n18967), .Z(n18581) );
  AND U19047 ( .A(n18582), .B(n18581), .Z(n18583) );
  OR U19048 ( .A(n18584), .B(n18583), .Z(n18586) );
  NAND U19049 ( .A(a[14]), .B(b[8]), .Z(n18972) );
  XOR U19050 ( .A(n18584), .B(n18583), .Z(n18973) );
  NANDN U19051 ( .A(n18972), .B(n18973), .Z(n18585) );
  NAND U19052 ( .A(n18586), .B(n18585), .Z(n18587) );
  OR U19053 ( .A(n18588), .B(n18587), .Z(n18592) );
  XNOR U19054 ( .A(n18588), .B(n18587), .Z(n18976) );
  XOR U19055 ( .A(n18590), .B(n18589), .Z(n18977) );
  NANDN U19056 ( .A(n18976), .B(n18977), .Z(n18591) );
  NAND U19057 ( .A(n18592), .B(n18591), .Z(n18593) );
  NANDN U19058 ( .A(n18594), .B(n18593), .Z(n18596) );
  ANDN U19059 ( .B(b[8]), .A(n173), .Z(n18985) );
  NANDN U19060 ( .A(n18985), .B(n18984), .Z(n18595) );
  AND U19061 ( .A(n18596), .B(n18595), .Z(n18599) );
  OR U19062 ( .A(n18600), .B(n18599), .Z(n18602) );
  XNOR U19063 ( .A(n18598), .B(n18597), .Z(n18989) );
  XNOR U19064 ( .A(n18600), .B(n18599), .Z(n18988) );
  OR U19065 ( .A(n18989), .B(n18988), .Z(n18601) );
  NAND U19066 ( .A(n18602), .B(n18601), .Z(n18605) );
  XOR U19067 ( .A(n18604), .B(n18603), .Z(n18606) );
  NANDN U19068 ( .A(n18605), .B(n18606), .Z(n18608) );
  NAND U19069 ( .A(a[18]), .B(b[8]), .Z(n18996) );
  XNOR U19070 ( .A(n18606), .B(n18605), .Z(n18997) );
  NANDN U19071 ( .A(n18996), .B(n18997), .Z(n18607) );
  NAND U19072 ( .A(n18608), .B(n18607), .Z(n18611) );
  OR U19073 ( .A(n18612), .B(n18611), .Z(n18614) );
  XOR U19074 ( .A(n18610), .B(n18609), .Z(n18888) );
  XOR U19075 ( .A(n18612), .B(n18611), .Z(n18887) );
  NAND U19076 ( .A(n18888), .B(n18887), .Z(n18613) );
  NAND U19077 ( .A(n18614), .B(n18613), .Z(n18617) );
  XOR U19078 ( .A(n18616), .B(n18615), .Z(n18618) );
  NANDN U19079 ( .A(n18617), .B(n18618), .Z(n18620) );
  NAND U19080 ( .A(a[20]), .B(b[8]), .Z(n19006) );
  XNOR U19081 ( .A(n18618), .B(n18617), .Z(n19007) );
  NANDN U19082 ( .A(n19006), .B(n19007), .Z(n18619) );
  NAND U19083 ( .A(n18620), .B(n18619), .Z(n18621) );
  OR U19084 ( .A(n18622), .B(n18621), .Z(n18626) );
  XNOR U19085 ( .A(n18622), .B(n18621), .Z(n19010) );
  XOR U19086 ( .A(n18624), .B(n18623), .Z(n19011) );
  NANDN U19087 ( .A(n19010), .B(n19011), .Z(n18625) );
  NAND U19088 ( .A(n18626), .B(n18625), .Z(n18629) );
  XOR U19089 ( .A(n18628), .B(n18627), .Z(n18630) );
  NANDN U19090 ( .A(n18629), .B(n18630), .Z(n18632) );
  NAND U19091 ( .A(a[22]), .B(b[8]), .Z(n19018) );
  XNOR U19092 ( .A(n18630), .B(n18629), .Z(n19019) );
  NANDN U19093 ( .A(n19018), .B(n19019), .Z(n18631) );
  NAND U19094 ( .A(n18632), .B(n18631), .Z(n18633) );
  OR U19095 ( .A(n18634), .B(n18633), .Z(n18638) );
  XNOR U19096 ( .A(n18634), .B(n18633), .Z(n19022) );
  XOR U19097 ( .A(n18636), .B(n18635), .Z(n19023) );
  NANDN U19098 ( .A(n19022), .B(n19023), .Z(n18637) );
  NAND U19099 ( .A(n18638), .B(n18637), .Z(n18641) );
  XOR U19100 ( .A(n18640), .B(n18639), .Z(n18642) );
  NANDN U19101 ( .A(n18641), .B(n18642), .Z(n18644) );
  NAND U19102 ( .A(a[24]), .B(b[8]), .Z(n19030) );
  XNOR U19103 ( .A(n18642), .B(n18641), .Z(n19031) );
  NANDN U19104 ( .A(n19030), .B(n19031), .Z(n18643) );
  NAND U19105 ( .A(n18644), .B(n18643), .Z(n18645) );
  OR U19106 ( .A(n18646), .B(n18645), .Z(n18650) );
  XNOR U19107 ( .A(n18646), .B(n18645), .Z(n19034) );
  XOR U19108 ( .A(n18648), .B(n18647), .Z(n19035) );
  NANDN U19109 ( .A(n19034), .B(n19035), .Z(n18649) );
  NAND U19110 ( .A(n18650), .B(n18649), .Z(n18653) );
  XOR U19111 ( .A(n18652), .B(n18651), .Z(n18654) );
  NANDN U19112 ( .A(n18653), .B(n18654), .Z(n18656) );
  NAND U19113 ( .A(a[26]), .B(b[8]), .Z(n19042) );
  XNOR U19114 ( .A(n18654), .B(n18653), .Z(n19043) );
  NANDN U19115 ( .A(n19042), .B(n19043), .Z(n18655) );
  NAND U19116 ( .A(n18656), .B(n18655), .Z(n18657) );
  OR U19117 ( .A(n18658), .B(n18657), .Z(n18662) );
  XNOR U19118 ( .A(n18658), .B(n18657), .Z(n19046) );
  XOR U19119 ( .A(n18660), .B(n18659), .Z(n19047) );
  NANDN U19120 ( .A(n19046), .B(n19047), .Z(n18661) );
  NAND U19121 ( .A(n18662), .B(n18661), .Z(n18665) );
  XOR U19122 ( .A(n18664), .B(n18663), .Z(n18666) );
  NANDN U19123 ( .A(n18665), .B(n18666), .Z(n18668) );
  NAND U19124 ( .A(a[28]), .B(b[8]), .Z(n19054) );
  XNOR U19125 ( .A(n18666), .B(n18665), .Z(n19055) );
  NANDN U19126 ( .A(n19054), .B(n19055), .Z(n18667) );
  NAND U19127 ( .A(n18668), .B(n18667), .Z(n18669) );
  OR U19128 ( .A(n18670), .B(n18669), .Z(n18674) );
  XNOR U19129 ( .A(n18670), .B(n18669), .Z(n19058) );
  XOR U19130 ( .A(n18672), .B(n18671), .Z(n19059) );
  NANDN U19131 ( .A(n19058), .B(n19059), .Z(n18673) );
  NAND U19132 ( .A(n18674), .B(n18673), .Z(n18677) );
  XOR U19133 ( .A(n18676), .B(n18675), .Z(n18678) );
  NANDN U19134 ( .A(n18677), .B(n18678), .Z(n18680) );
  NAND U19135 ( .A(a[30]), .B(b[8]), .Z(n19066) );
  XNOR U19136 ( .A(n18678), .B(n18677), .Z(n19067) );
  NANDN U19137 ( .A(n19066), .B(n19067), .Z(n18679) );
  NAND U19138 ( .A(n18680), .B(n18679), .Z(n18681) );
  OR U19139 ( .A(n18682), .B(n18681), .Z(n18686) );
  XNOR U19140 ( .A(n18682), .B(n18681), .Z(n19070) );
  XOR U19141 ( .A(n18684), .B(n18683), .Z(n19071) );
  NANDN U19142 ( .A(n19070), .B(n19071), .Z(n18685) );
  NAND U19143 ( .A(n18686), .B(n18685), .Z(n18689) );
  XOR U19144 ( .A(n18688), .B(n18687), .Z(n18690) );
  NANDN U19145 ( .A(n18689), .B(n18690), .Z(n18692) );
  NAND U19146 ( .A(a[32]), .B(b[8]), .Z(n19078) );
  XNOR U19147 ( .A(n18690), .B(n18689), .Z(n19079) );
  NANDN U19148 ( .A(n19078), .B(n19079), .Z(n18691) );
  NAND U19149 ( .A(n18692), .B(n18691), .Z(n18693) );
  OR U19150 ( .A(n18694), .B(n18693), .Z(n18698) );
  XNOR U19151 ( .A(n18694), .B(n18693), .Z(n19082) );
  XOR U19152 ( .A(n18696), .B(n18695), .Z(n19083) );
  NANDN U19153 ( .A(n19082), .B(n19083), .Z(n18697) );
  NAND U19154 ( .A(n18698), .B(n18697), .Z(n18701) );
  XOR U19155 ( .A(n18700), .B(n18699), .Z(n18702) );
  NANDN U19156 ( .A(n18701), .B(n18702), .Z(n18704) );
  NAND U19157 ( .A(a[34]), .B(b[8]), .Z(n19090) );
  XNOR U19158 ( .A(n18702), .B(n18701), .Z(n19091) );
  NANDN U19159 ( .A(n19090), .B(n19091), .Z(n18703) );
  NAND U19160 ( .A(n18704), .B(n18703), .Z(n18705) );
  OR U19161 ( .A(n18706), .B(n18705), .Z(n18710) );
  XNOR U19162 ( .A(n18706), .B(n18705), .Z(n19094) );
  XOR U19163 ( .A(n18708), .B(n18707), .Z(n19095) );
  NANDN U19164 ( .A(n19094), .B(n19095), .Z(n18709) );
  NAND U19165 ( .A(n18710), .B(n18709), .Z(n18713) );
  XOR U19166 ( .A(n18712), .B(n18711), .Z(n18714) );
  NANDN U19167 ( .A(n18713), .B(n18714), .Z(n18716) );
  NAND U19168 ( .A(a[36]), .B(b[8]), .Z(n19102) );
  XNOR U19169 ( .A(n18714), .B(n18713), .Z(n19103) );
  NANDN U19170 ( .A(n19102), .B(n19103), .Z(n18715) );
  NAND U19171 ( .A(n18716), .B(n18715), .Z(n18717) );
  OR U19172 ( .A(n18718), .B(n18717), .Z(n18722) );
  XNOR U19173 ( .A(n18718), .B(n18717), .Z(n19106) );
  XOR U19174 ( .A(n18720), .B(n18719), .Z(n19107) );
  NANDN U19175 ( .A(n19106), .B(n19107), .Z(n18721) );
  NAND U19176 ( .A(n18722), .B(n18721), .Z(n18725) );
  XOR U19177 ( .A(n18724), .B(n18723), .Z(n18726) );
  NANDN U19178 ( .A(n18725), .B(n18726), .Z(n18728) );
  NAND U19179 ( .A(a[38]), .B(b[8]), .Z(n19114) );
  XNOR U19180 ( .A(n18726), .B(n18725), .Z(n19115) );
  NANDN U19181 ( .A(n19114), .B(n19115), .Z(n18727) );
  NAND U19182 ( .A(n18728), .B(n18727), .Z(n18729) );
  OR U19183 ( .A(n18730), .B(n18729), .Z(n18734) );
  XNOR U19184 ( .A(n18730), .B(n18729), .Z(n19118) );
  XOR U19185 ( .A(n18732), .B(n18731), .Z(n19119) );
  NANDN U19186 ( .A(n19118), .B(n19119), .Z(n18733) );
  NAND U19187 ( .A(n18734), .B(n18733), .Z(n18737) );
  XOR U19188 ( .A(n18736), .B(n18735), .Z(n18738) );
  NANDN U19189 ( .A(n18737), .B(n18738), .Z(n18740) );
  NAND U19190 ( .A(a[40]), .B(b[8]), .Z(n19126) );
  XNOR U19191 ( .A(n18738), .B(n18737), .Z(n19127) );
  NANDN U19192 ( .A(n19126), .B(n19127), .Z(n18739) );
  NAND U19193 ( .A(n18740), .B(n18739), .Z(n18741) );
  OR U19194 ( .A(n18742), .B(n18741), .Z(n18746) );
  XNOR U19195 ( .A(n18742), .B(n18741), .Z(n19130) );
  XOR U19196 ( .A(n18744), .B(n18743), .Z(n19131) );
  NANDN U19197 ( .A(n19130), .B(n19131), .Z(n18745) );
  NAND U19198 ( .A(n18746), .B(n18745), .Z(n18749) );
  XOR U19199 ( .A(n18748), .B(n18747), .Z(n18750) );
  NANDN U19200 ( .A(n18749), .B(n18750), .Z(n18752) );
  NAND U19201 ( .A(a[42]), .B(b[8]), .Z(n19138) );
  XNOR U19202 ( .A(n18750), .B(n18749), .Z(n19139) );
  NANDN U19203 ( .A(n19138), .B(n19139), .Z(n18751) );
  NAND U19204 ( .A(n18752), .B(n18751), .Z(n18753) );
  OR U19205 ( .A(n18754), .B(n18753), .Z(n18758) );
  XNOR U19206 ( .A(n18754), .B(n18753), .Z(n19142) );
  XOR U19207 ( .A(n18756), .B(n18755), .Z(n19143) );
  NANDN U19208 ( .A(n19142), .B(n19143), .Z(n18757) );
  NAND U19209 ( .A(n18758), .B(n18757), .Z(n18761) );
  XOR U19210 ( .A(n18760), .B(n18759), .Z(n18762) );
  NANDN U19211 ( .A(n18761), .B(n18762), .Z(n18764) );
  NAND U19212 ( .A(a[44]), .B(b[8]), .Z(n19150) );
  XNOR U19213 ( .A(n18762), .B(n18761), .Z(n19151) );
  NANDN U19214 ( .A(n19150), .B(n19151), .Z(n18763) );
  NAND U19215 ( .A(n18764), .B(n18763), .Z(n18765) );
  OR U19216 ( .A(n18766), .B(n18765), .Z(n18770) );
  XNOR U19217 ( .A(n18766), .B(n18765), .Z(n19154) );
  XOR U19218 ( .A(n18768), .B(n18767), .Z(n19155) );
  NANDN U19219 ( .A(n19154), .B(n19155), .Z(n18769) );
  NAND U19220 ( .A(n18770), .B(n18769), .Z(n18773) );
  XOR U19221 ( .A(n18772), .B(n18771), .Z(n18774) );
  NANDN U19222 ( .A(n18773), .B(n18774), .Z(n18776) );
  NAND U19223 ( .A(a[46]), .B(b[8]), .Z(n19162) );
  XNOR U19224 ( .A(n18774), .B(n18773), .Z(n19163) );
  NANDN U19225 ( .A(n19162), .B(n19163), .Z(n18775) );
  NAND U19226 ( .A(n18776), .B(n18775), .Z(n18777) );
  OR U19227 ( .A(n18778), .B(n18777), .Z(n18782) );
  XNOR U19228 ( .A(n18778), .B(n18777), .Z(n19166) );
  XOR U19229 ( .A(n18780), .B(n18779), .Z(n19167) );
  NANDN U19230 ( .A(n19166), .B(n19167), .Z(n18781) );
  NAND U19231 ( .A(n18782), .B(n18781), .Z(n18785) );
  XOR U19232 ( .A(n18784), .B(n18783), .Z(n18786) );
  NANDN U19233 ( .A(n18785), .B(n18786), .Z(n18788) );
  NAND U19234 ( .A(a[48]), .B(b[8]), .Z(n19174) );
  XNOR U19235 ( .A(n18786), .B(n18785), .Z(n19175) );
  NANDN U19236 ( .A(n19174), .B(n19175), .Z(n18787) );
  NAND U19237 ( .A(n18788), .B(n18787), .Z(n18789) );
  OR U19238 ( .A(n18790), .B(n18789), .Z(n18794) );
  XNOR U19239 ( .A(n18790), .B(n18789), .Z(n19178) );
  XOR U19240 ( .A(n18792), .B(n18791), .Z(n19179) );
  NANDN U19241 ( .A(n19178), .B(n19179), .Z(n18793) );
  NAND U19242 ( .A(n18794), .B(n18793), .Z(n18797) );
  XOR U19243 ( .A(n18796), .B(n18795), .Z(n18798) );
  NANDN U19244 ( .A(n18797), .B(n18798), .Z(n18800) );
  NAND U19245 ( .A(a[50]), .B(b[8]), .Z(n19186) );
  XNOR U19246 ( .A(n18798), .B(n18797), .Z(n19187) );
  NANDN U19247 ( .A(n19186), .B(n19187), .Z(n18799) );
  NAND U19248 ( .A(n18800), .B(n18799), .Z(n18801) );
  OR U19249 ( .A(n18802), .B(n18801), .Z(n18806) );
  XNOR U19250 ( .A(n18802), .B(n18801), .Z(n19190) );
  XOR U19251 ( .A(n18804), .B(n18803), .Z(n19191) );
  NANDN U19252 ( .A(n19190), .B(n19191), .Z(n18805) );
  NAND U19253 ( .A(n18806), .B(n18805), .Z(n18809) );
  XOR U19254 ( .A(n18808), .B(n18807), .Z(n18810) );
  NANDN U19255 ( .A(n18809), .B(n18810), .Z(n18812) );
  NAND U19256 ( .A(a[52]), .B(b[8]), .Z(n19198) );
  XNOR U19257 ( .A(n18810), .B(n18809), .Z(n19199) );
  NANDN U19258 ( .A(n19198), .B(n19199), .Z(n18811) );
  NAND U19259 ( .A(n18812), .B(n18811), .Z(n18813) );
  OR U19260 ( .A(n18814), .B(n18813), .Z(n18818) );
  XNOR U19261 ( .A(n18814), .B(n18813), .Z(n19202) );
  XOR U19262 ( .A(n18816), .B(n18815), .Z(n19203) );
  NANDN U19263 ( .A(n19202), .B(n19203), .Z(n18817) );
  NAND U19264 ( .A(n18818), .B(n18817), .Z(n18821) );
  XNOR U19265 ( .A(n18820), .B(n18819), .Z(n18822) );
  OR U19266 ( .A(n18821), .B(n18822), .Z(n18824) );
  XNOR U19267 ( .A(n18822), .B(n18821), .Z(n19209) );
  NAND U19268 ( .A(a[54]), .B(b[8]), .Z(n19208) );
  OR U19269 ( .A(n19209), .B(n19208), .Z(n18823) );
  NAND U19270 ( .A(n18824), .B(n18823), .Z(n18827) );
  ANDN U19271 ( .B(b[8]), .A(n203), .Z(n18828) );
  OR U19272 ( .A(n18827), .B(n18828), .Z(n18830) );
  XOR U19273 ( .A(n18826), .B(n18825), .Z(n19215) );
  XOR U19274 ( .A(n18828), .B(n18827), .Z(n19214) );
  NANDN U19275 ( .A(n19215), .B(n19214), .Z(n18829) );
  NAND U19276 ( .A(n18830), .B(n18829), .Z(n18832) );
  AND U19277 ( .A(b[8]), .B(a[56]), .Z(n18831) );
  NANDN U19278 ( .A(n18832), .B(n18831), .Z(n18836) );
  XNOR U19279 ( .A(n18832), .B(n18831), .Z(n19220) );
  NAND U19280 ( .A(n19220), .B(n19221), .Z(n18835) );
  NAND U19281 ( .A(n18836), .B(n18835), .Z(n18840) );
  XOR U19282 ( .A(n18838), .B(n18837), .Z(n18839) );
  NAND U19283 ( .A(n18840), .B(n18839), .Z(n18842) );
  XNOR U19284 ( .A(n18840), .B(n18839), .Z(n19227) );
  NAND U19285 ( .A(a[57]), .B(b[8]), .Z(n19226) );
  OR U19286 ( .A(n19227), .B(n19226), .Z(n18841) );
  NAND U19287 ( .A(n18842), .B(n18841), .Z(n18846) );
  NANDN U19288 ( .A(n18845), .B(n18846), .Z(n18848) );
  XOR U19289 ( .A(n18844), .B(n18843), .Z(n19232) );
  XNOR U19290 ( .A(n18846), .B(n18845), .Z(n19233) );
  NAND U19291 ( .A(n19232), .B(n19233), .Z(n18847) );
  NAND U19292 ( .A(n18848), .B(n18847), .Z(n18851) );
  AND U19293 ( .A(b[8]), .B(a[59]), .Z(n18852) );
  OR U19294 ( .A(n18851), .B(n18852), .Z(n18854) );
  XNOR U19295 ( .A(n18850), .B(n18849), .Z(n19239) );
  XOR U19296 ( .A(n18852), .B(n18851), .Z(n19238) );
  NANDN U19297 ( .A(n19239), .B(n19238), .Z(n18853) );
  NAND U19298 ( .A(n18854), .B(n18853), .Z(n18858) );
  NAND U19299 ( .A(a[60]), .B(b[8]), .Z(n18857) );
  OR U19300 ( .A(n18858), .B(n18857), .Z(n18860) );
  XOR U19301 ( .A(n18856), .B(n18855), .Z(n19244) );
  XOR U19302 ( .A(n18858), .B(n18857), .Z(n19245) );
  NAND U19303 ( .A(n19244), .B(n19245), .Z(n18859) );
  NAND U19304 ( .A(n18860), .B(n18859), .Z(n18863) );
  AND U19305 ( .A(b[8]), .B(a[61]), .Z(n18864) );
  OR U19306 ( .A(n18863), .B(n18864), .Z(n18866) );
  XNOR U19307 ( .A(n18862), .B(n18861), .Z(n19249) );
  XOR U19308 ( .A(n18864), .B(n18863), .Z(n19248) );
  NANDN U19309 ( .A(n19249), .B(n19248), .Z(n18865) );
  NAND U19310 ( .A(n18866), .B(n18865), .Z(n18870) );
  NAND U19311 ( .A(a[62]), .B(b[8]), .Z(n18869) );
  OR U19312 ( .A(n18870), .B(n18869), .Z(n18872) );
  XOR U19313 ( .A(n18868), .B(n18867), .Z(n19254) );
  XOR U19314 ( .A(n18870), .B(n18869), .Z(n19255) );
  NANDN U19315 ( .A(n19254), .B(n19255), .Z(n18871) );
  NAND U19316 ( .A(n18872), .B(n18871), .Z(n18875) );
  AND U19317 ( .A(b[8]), .B(a[63]), .Z(n18876) );
  OR U19318 ( .A(n18875), .B(n18876), .Z(n18878) );
  XNOR U19319 ( .A(n18874), .B(n18873), .Z(n18886) );
  XOR U19320 ( .A(n18876), .B(n18875), .Z(n18885) );
  NANDN U19321 ( .A(n18886), .B(n18885), .Z(n18877) );
  NAND U19322 ( .A(n18878), .B(n18877), .Z(n18883) );
  OR U19323 ( .A(n18884), .B(n18883), .Z(n18882) );
  XOR U19324 ( .A(n18880), .B(n18879), .Z(n18881) );
  NAND U19325 ( .A(n18882), .B(n18881), .Z(n21937) );
  XNOR U19326 ( .A(n18882), .B(n18881), .Z(n24116) );
  XOR U19327 ( .A(n18884), .B(n18883), .Z(n21932) );
  XNOR U19328 ( .A(n18886), .B(n18885), .Z(n19638) );
  NAND U19329 ( .A(a[60]), .B(b[7]), .Z(n19240) );
  ANDN U19330 ( .B(b[7]), .A(n201), .Z(n19197) );
  ANDN U19331 ( .B(b[7]), .A(n199), .Z(n19185) );
  ANDN U19332 ( .B(b[7]), .A(n197), .Z(n19173) );
  ANDN U19333 ( .B(b[7]), .A(n195), .Z(n19161) );
  ANDN U19334 ( .B(b[7]), .A(n193), .Z(n19149) );
  ANDN U19335 ( .B(b[7]), .A(n191), .Z(n19137) );
  ANDN U19336 ( .B(b[7]), .A(n189), .Z(n19125) );
  ANDN U19337 ( .B(b[7]), .A(n187), .Z(n19113) );
  ANDN U19338 ( .B(b[7]), .A(n21772), .Z(n19101) );
  ANDN U19339 ( .B(b[7]), .A(n184), .Z(n19089) );
  ANDN U19340 ( .B(b[7]), .A(n21751), .Z(n19077) );
  ANDN U19341 ( .B(b[7]), .A(n21740), .Z(n19065) );
  ANDN U19342 ( .B(b[7]), .A(n21727), .Z(n19053) );
  ANDN U19343 ( .B(b[7]), .A(n21716), .Z(n19041) );
  ANDN U19344 ( .B(b[7]), .A(n21703), .Z(n19029) );
  ANDN U19345 ( .B(b[7]), .A(n21692), .Z(n19017) );
  ANDN U19346 ( .B(b[7]), .A(n21681), .Z(n19005) );
  XNOR U19347 ( .A(n18888), .B(n18887), .Z(n19001) );
  ANDN U19348 ( .B(b[7]), .A(n21670), .Z(n18995) );
  NAND U19349 ( .A(a[17]), .B(b[7]), .Z(n18983) );
  ANDN U19350 ( .B(b[7]), .A(n172), .Z(n18971) );
  ANDN U19351 ( .B(b[7]), .A(n170), .Z(n18959) );
  ANDN U19352 ( .B(b[7]), .A(n21164), .Z(n18947) );
  ANDN U19353 ( .B(b[7]), .A(n21615), .Z(n18935) );
  ANDN U19354 ( .B(b[7]), .A(n166), .Z(n18923) );
  NAND U19355 ( .A(a[6]), .B(b[7]), .Z(n18918) );
  XOR U19356 ( .A(n18890), .B(n18889), .Z(n18919) );
  NANDN U19357 ( .A(n18918), .B(n18919), .Z(n18921) );
  ANDN U19358 ( .B(b[7]), .A(n164), .Z(n18913) );
  ANDN U19359 ( .B(b[7]), .A(n21580), .Z(n18900) );
  NAND U19360 ( .A(b[8]), .B(a[1]), .Z(n18895) );
  NANDN U19361 ( .A(n18895), .B(a[0]), .Z(n18891) );
  XNOR U19362 ( .A(a[2]), .B(n18891), .Z(n18892) );
  NAND U19363 ( .A(b[7]), .B(n18892), .Z(n19277) );
  AND U19364 ( .A(a[1]), .B(b[8]), .Z(n18893) );
  XOR U19365 ( .A(n18894), .B(n18893), .Z(n19278) );
  OR U19366 ( .A(n19277), .B(n19278), .Z(n18899) );
  AND U19367 ( .A(b[7]), .B(a[0]), .Z(n19654) );
  NANDN U19368 ( .A(n18895), .B(n19654), .Z(n18897) );
  NAND U19369 ( .A(a[2]), .B(b[7]), .Z(n18896) );
  AND U19370 ( .A(n18897), .B(n18896), .Z(n18898) );
  ANDN U19371 ( .B(n18899), .A(n18898), .Z(n18901) );
  OR U19372 ( .A(n18900), .B(n18901), .Z(n18905) );
  XNOR U19373 ( .A(n18901), .B(n18900), .Z(n19282) );
  XNOR U19374 ( .A(n18903), .B(n18902), .Z(n19281) );
  OR U19375 ( .A(n19282), .B(n19281), .Z(n18904) );
  NAND U19376 ( .A(n18905), .B(n18904), .Z(n18909) );
  XOR U19377 ( .A(n18907), .B(n18906), .Z(n18908) );
  OR U19378 ( .A(n18909), .B(n18908), .Z(n18911) );
  NAND U19379 ( .A(a[4]), .B(b[7]), .Z(n19290) );
  XOR U19380 ( .A(n18909), .B(n18908), .Z(n19289) );
  NANDN U19381 ( .A(n19290), .B(n19289), .Z(n18910) );
  NAND U19382 ( .A(n18911), .B(n18910), .Z(n18912) );
  OR U19383 ( .A(n18913), .B(n18912), .Z(n18917) );
  XNOR U19384 ( .A(n18913), .B(n18912), .Z(n19264) );
  XOR U19385 ( .A(n18915), .B(n18914), .Z(n19265) );
  NANDN U19386 ( .A(n19264), .B(n19265), .Z(n18916) );
  NAND U19387 ( .A(n18917), .B(n18916), .Z(n19299) );
  XNOR U19388 ( .A(n18919), .B(n18918), .Z(n19300) );
  NANDN U19389 ( .A(n19299), .B(n19300), .Z(n18920) );
  NAND U19390 ( .A(n18921), .B(n18920), .Z(n18922) );
  OR U19391 ( .A(n18923), .B(n18922), .Z(n18927) );
  XNOR U19392 ( .A(n18923), .B(n18922), .Z(n19262) );
  XOR U19393 ( .A(n18925), .B(n18924), .Z(n19263) );
  NANDN U19394 ( .A(n19262), .B(n19263), .Z(n18926) );
  NAND U19395 ( .A(n18927), .B(n18926), .Z(n18930) );
  XOR U19396 ( .A(n18929), .B(n18928), .Z(n18931) );
  NANDN U19397 ( .A(n18930), .B(n18931), .Z(n18933) );
  NAND U19398 ( .A(a[8]), .B(b[7]), .Z(n19309) );
  XNOR U19399 ( .A(n18931), .B(n18930), .Z(n19310) );
  NANDN U19400 ( .A(n19309), .B(n19310), .Z(n18932) );
  NAND U19401 ( .A(n18933), .B(n18932), .Z(n18934) );
  OR U19402 ( .A(n18935), .B(n18934), .Z(n18939) );
  XNOR U19403 ( .A(n18935), .B(n18934), .Z(n19260) );
  XOR U19404 ( .A(n18937), .B(n18936), .Z(n19261) );
  NANDN U19405 ( .A(n19260), .B(n19261), .Z(n18938) );
  NAND U19406 ( .A(n18939), .B(n18938), .Z(n18942) );
  XOR U19407 ( .A(n18941), .B(n18940), .Z(n18943) );
  NANDN U19408 ( .A(n18942), .B(n18943), .Z(n18945) );
  NAND U19409 ( .A(a[10]), .B(b[7]), .Z(n19319) );
  XNOR U19410 ( .A(n18943), .B(n18942), .Z(n19320) );
  NANDN U19411 ( .A(n19319), .B(n19320), .Z(n18944) );
  NAND U19412 ( .A(n18945), .B(n18944), .Z(n18946) );
  OR U19413 ( .A(n18947), .B(n18946), .Z(n18951) );
  XNOR U19414 ( .A(n18947), .B(n18946), .Z(n19323) );
  XOR U19415 ( .A(n18949), .B(n18948), .Z(n19324) );
  NANDN U19416 ( .A(n19323), .B(n19324), .Z(n18950) );
  NAND U19417 ( .A(n18951), .B(n18950), .Z(n18954) );
  XOR U19418 ( .A(n18953), .B(n18952), .Z(n18955) );
  NANDN U19419 ( .A(n18954), .B(n18955), .Z(n18957) );
  NAND U19420 ( .A(a[12]), .B(b[7]), .Z(n19331) );
  XNOR U19421 ( .A(n18955), .B(n18954), .Z(n19332) );
  NANDN U19422 ( .A(n19331), .B(n19332), .Z(n18956) );
  NAND U19423 ( .A(n18957), .B(n18956), .Z(n18958) );
  OR U19424 ( .A(n18959), .B(n18958), .Z(n18963) );
  XNOR U19425 ( .A(n18959), .B(n18958), .Z(n19335) );
  XOR U19426 ( .A(n18961), .B(n18960), .Z(n19336) );
  NANDN U19427 ( .A(n19335), .B(n19336), .Z(n18962) );
  NAND U19428 ( .A(n18963), .B(n18962), .Z(n18965) );
  NAND U19429 ( .A(a[14]), .B(b[7]), .Z(n18964) );
  OR U19430 ( .A(n18965), .B(n18964), .Z(n18969) );
  XOR U19431 ( .A(n18965), .B(n18964), .Z(n19341) );
  NAND U19432 ( .A(n19341), .B(n19342), .Z(n18968) );
  NAND U19433 ( .A(n18969), .B(n18968), .Z(n18970) );
  OR U19434 ( .A(n18971), .B(n18970), .Z(n18975) );
  XNOR U19435 ( .A(n18971), .B(n18970), .Z(n19347) );
  XOR U19436 ( .A(n18973), .B(n18972), .Z(n19348) );
  NANDN U19437 ( .A(n19347), .B(n19348), .Z(n18974) );
  NAND U19438 ( .A(n18975), .B(n18974), .Z(n18978) );
  XOR U19439 ( .A(n18977), .B(n18976), .Z(n18979) );
  NANDN U19440 ( .A(n18978), .B(n18979), .Z(n18981) );
  NAND U19441 ( .A(a[16]), .B(b[7]), .Z(n19355) );
  XNOR U19442 ( .A(n18979), .B(n18978), .Z(n19356) );
  NANDN U19443 ( .A(n19355), .B(n19356), .Z(n18980) );
  NAND U19444 ( .A(n18981), .B(n18980), .Z(n18982) );
  NANDN U19445 ( .A(n18983), .B(n18982), .Z(n18987) );
  NAND U19446 ( .A(n19361), .B(n19362), .Z(n18986) );
  NAND U19447 ( .A(n18987), .B(n18986), .Z(n18991) );
  XOR U19448 ( .A(n18989), .B(n18988), .Z(n18990) );
  NANDN U19449 ( .A(n18991), .B(n18990), .Z(n18993) );
  ANDN U19450 ( .B(b[7]), .A(n175), .Z(n19366) );
  XOR U19451 ( .A(n18991), .B(n18990), .Z(n19365) );
  OR U19452 ( .A(n19366), .B(n19365), .Z(n18992) );
  AND U19453 ( .A(n18993), .B(n18992), .Z(n18994) );
  OR U19454 ( .A(n18995), .B(n18994), .Z(n18999) );
  XNOR U19455 ( .A(n18995), .B(n18994), .Z(n19371) );
  XOR U19456 ( .A(n18997), .B(n18996), .Z(n19372) );
  NANDN U19457 ( .A(n19371), .B(n19372), .Z(n18998) );
  NAND U19458 ( .A(n18999), .B(n18998), .Z(n19000) );
  NANDN U19459 ( .A(n19001), .B(n19000), .Z(n19003) );
  ANDN U19460 ( .B(b[7]), .A(n176), .Z(n19378) );
  NANDN U19461 ( .A(n19378), .B(n19377), .Z(n19002) );
  NAND U19462 ( .A(n19003), .B(n19002), .Z(n19004) );
  NANDN U19463 ( .A(n19005), .B(n19004), .Z(n19009) );
  XOR U19464 ( .A(n19007), .B(n19006), .Z(n19383) );
  NANDN U19465 ( .A(n19384), .B(n19383), .Z(n19008) );
  NAND U19466 ( .A(n19009), .B(n19008), .Z(n19012) );
  XOR U19467 ( .A(n19011), .B(n19010), .Z(n19013) );
  NANDN U19468 ( .A(n19012), .B(n19013), .Z(n19015) );
  NAND U19469 ( .A(a[22]), .B(b[7]), .Z(n19391) );
  XNOR U19470 ( .A(n19013), .B(n19012), .Z(n19392) );
  NANDN U19471 ( .A(n19391), .B(n19392), .Z(n19014) );
  NAND U19472 ( .A(n19015), .B(n19014), .Z(n19016) );
  OR U19473 ( .A(n19017), .B(n19016), .Z(n19021) );
  XNOR U19474 ( .A(n19017), .B(n19016), .Z(n19395) );
  XOR U19475 ( .A(n19019), .B(n19018), .Z(n19396) );
  NANDN U19476 ( .A(n19395), .B(n19396), .Z(n19020) );
  NAND U19477 ( .A(n19021), .B(n19020), .Z(n19024) );
  XOR U19478 ( .A(n19023), .B(n19022), .Z(n19025) );
  NANDN U19479 ( .A(n19024), .B(n19025), .Z(n19027) );
  NAND U19480 ( .A(a[24]), .B(b[7]), .Z(n19403) );
  XNOR U19481 ( .A(n19025), .B(n19024), .Z(n19404) );
  NANDN U19482 ( .A(n19403), .B(n19404), .Z(n19026) );
  NAND U19483 ( .A(n19027), .B(n19026), .Z(n19028) );
  OR U19484 ( .A(n19029), .B(n19028), .Z(n19033) );
  XNOR U19485 ( .A(n19029), .B(n19028), .Z(n19407) );
  XOR U19486 ( .A(n19031), .B(n19030), .Z(n19408) );
  NANDN U19487 ( .A(n19407), .B(n19408), .Z(n19032) );
  NAND U19488 ( .A(n19033), .B(n19032), .Z(n19036) );
  XOR U19489 ( .A(n19035), .B(n19034), .Z(n19037) );
  NANDN U19490 ( .A(n19036), .B(n19037), .Z(n19039) );
  NAND U19491 ( .A(a[26]), .B(b[7]), .Z(n19415) );
  XNOR U19492 ( .A(n19037), .B(n19036), .Z(n19416) );
  NANDN U19493 ( .A(n19415), .B(n19416), .Z(n19038) );
  NAND U19494 ( .A(n19039), .B(n19038), .Z(n19040) );
  OR U19495 ( .A(n19041), .B(n19040), .Z(n19045) );
  XNOR U19496 ( .A(n19041), .B(n19040), .Z(n19419) );
  XOR U19497 ( .A(n19043), .B(n19042), .Z(n19420) );
  NANDN U19498 ( .A(n19419), .B(n19420), .Z(n19044) );
  NAND U19499 ( .A(n19045), .B(n19044), .Z(n19048) );
  XOR U19500 ( .A(n19047), .B(n19046), .Z(n19049) );
  NANDN U19501 ( .A(n19048), .B(n19049), .Z(n19051) );
  NAND U19502 ( .A(a[28]), .B(b[7]), .Z(n19427) );
  XNOR U19503 ( .A(n19049), .B(n19048), .Z(n19428) );
  NANDN U19504 ( .A(n19427), .B(n19428), .Z(n19050) );
  NAND U19505 ( .A(n19051), .B(n19050), .Z(n19052) );
  OR U19506 ( .A(n19053), .B(n19052), .Z(n19057) );
  XNOR U19507 ( .A(n19053), .B(n19052), .Z(n19431) );
  XOR U19508 ( .A(n19055), .B(n19054), .Z(n19432) );
  NANDN U19509 ( .A(n19431), .B(n19432), .Z(n19056) );
  NAND U19510 ( .A(n19057), .B(n19056), .Z(n19060) );
  XOR U19511 ( .A(n19059), .B(n19058), .Z(n19061) );
  NANDN U19512 ( .A(n19060), .B(n19061), .Z(n19063) );
  NAND U19513 ( .A(a[30]), .B(b[7]), .Z(n19439) );
  XNOR U19514 ( .A(n19061), .B(n19060), .Z(n19440) );
  NANDN U19515 ( .A(n19439), .B(n19440), .Z(n19062) );
  NAND U19516 ( .A(n19063), .B(n19062), .Z(n19064) );
  OR U19517 ( .A(n19065), .B(n19064), .Z(n19069) );
  XNOR U19518 ( .A(n19065), .B(n19064), .Z(n19443) );
  XOR U19519 ( .A(n19067), .B(n19066), .Z(n19444) );
  NANDN U19520 ( .A(n19443), .B(n19444), .Z(n19068) );
  NAND U19521 ( .A(n19069), .B(n19068), .Z(n19072) );
  XOR U19522 ( .A(n19071), .B(n19070), .Z(n19073) );
  NANDN U19523 ( .A(n19072), .B(n19073), .Z(n19075) );
  NAND U19524 ( .A(a[32]), .B(b[7]), .Z(n19451) );
  XNOR U19525 ( .A(n19073), .B(n19072), .Z(n19452) );
  NANDN U19526 ( .A(n19451), .B(n19452), .Z(n19074) );
  NAND U19527 ( .A(n19075), .B(n19074), .Z(n19076) );
  OR U19528 ( .A(n19077), .B(n19076), .Z(n19081) );
  XNOR U19529 ( .A(n19077), .B(n19076), .Z(n19455) );
  XOR U19530 ( .A(n19079), .B(n19078), .Z(n19456) );
  NANDN U19531 ( .A(n19455), .B(n19456), .Z(n19080) );
  NAND U19532 ( .A(n19081), .B(n19080), .Z(n19084) );
  XOR U19533 ( .A(n19083), .B(n19082), .Z(n19085) );
  NANDN U19534 ( .A(n19084), .B(n19085), .Z(n19087) );
  NAND U19535 ( .A(a[34]), .B(b[7]), .Z(n19463) );
  XNOR U19536 ( .A(n19085), .B(n19084), .Z(n19464) );
  NANDN U19537 ( .A(n19463), .B(n19464), .Z(n19086) );
  NAND U19538 ( .A(n19087), .B(n19086), .Z(n19088) );
  OR U19539 ( .A(n19089), .B(n19088), .Z(n19093) );
  XNOR U19540 ( .A(n19089), .B(n19088), .Z(n19467) );
  XOR U19541 ( .A(n19091), .B(n19090), .Z(n19468) );
  NANDN U19542 ( .A(n19467), .B(n19468), .Z(n19092) );
  NAND U19543 ( .A(n19093), .B(n19092), .Z(n19096) );
  XOR U19544 ( .A(n19095), .B(n19094), .Z(n19097) );
  NANDN U19545 ( .A(n19096), .B(n19097), .Z(n19099) );
  NAND U19546 ( .A(a[36]), .B(b[7]), .Z(n19475) );
  XNOR U19547 ( .A(n19097), .B(n19096), .Z(n19476) );
  NANDN U19548 ( .A(n19475), .B(n19476), .Z(n19098) );
  NAND U19549 ( .A(n19099), .B(n19098), .Z(n19100) );
  OR U19550 ( .A(n19101), .B(n19100), .Z(n19105) );
  XNOR U19551 ( .A(n19101), .B(n19100), .Z(n19479) );
  XOR U19552 ( .A(n19103), .B(n19102), .Z(n19480) );
  NANDN U19553 ( .A(n19479), .B(n19480), .Z(n19104) );
  NAND U19554 ( .A(n19105), .B(n19104), .Z(n19108) );
  XOR U19555 ( .A(n19107), .B(n19106), .Z(n19109) );
  NANDN U19556 ( .A(n19108), .B(n19109), .Z(n19111) );
  NAND U19557 ( .A(a[38]), .B(b[7]), .Z(n19487) );
  XNOR U19558 ( .A(n19109), .B(n19108), .Z(n19488) );
  NANDN U19559 ( .A(n19487), .B(n19488), .Z(n19110) );
  NAND U19560 ( .A(n19111), .B(n19110), .Z(n19112) );
  OR U19561 ( .A(n19113), .B(n19112), .Z(n19117) );
  XNOR U19562 ( .A(n19113), .B(n19112), .Z(n19491) );
  XOR U19563 ( .A(n19115), .B(n19114), .Z(n19492) );
  NANDN U19564 ( .A(n19491), .B(n19492), .Z(n19116) );
  NAND U19565 ( .A(n19117), .B(n19116), .Z(n19120) );
  XOR U19566 ( .A(n19119), .B(n19118), .Z(n19121) );
  NANDN U19567 ( .A(n19120), .B(n19121), .Z(n19123) );
  NAND U19568 ( .A(a[40]), .B(b[7]), .Z(n19499) );
  XNOR U19569 ( .A(n19121), .B(n19120), .Z(n19500) );
  NANDN U19570 ( .A(n19499), .B(n19500), .Z(n19122) );
  NAND U19571 ( .A(n19123), .B(n19122), .Z(n19124) );
  OR U19572 ( .A(n19125), .B(n19124), .Z(n19129) );
  XNOR U19573 ( .A(n19125), .B(n19124), .Z(n19503) );
  XOR U19574 ( .A(n19127), .B(n19126), .Z(n19504) );
  NANDN U19575 ( .A(n19503), .B(n19504), .Z(n19128) );
  NAND U19576 ( .A(n19129), .B(n19128), .Z(n19132) );
  XOR U19577 ( .A(n19131), .B(n19130), .Z(n19133) );
  NANDN U19578 ( .A(n19132), .B(n19133), .Z(n19135) );
  NAND U19579 ( .A(a[42]), .B(b[7]), .Z(n19511) );
  XNOR U19580 ( .A(n19133), .B(n19132), .Z(n19512) );
  NANDN U19581 ( .A(n19511), .B(n19512), .Z(n19134) );
  NAND U19582 ( .A(n19135), .B(n19134), .Z(n19136) );
  OR U19583 ( .A(n19137), .B(n19136), .Z(n19141) );
  XNOR U19584 ( .A(n19137), .B(n19136), .Z(n19515) );
  XOR U19585 ( .A(n19139), .B(n19138), .Z(n19516) );
  NANDN U19586 ( .A(n19515), .B(n19516), .Z(n19140) );
  NAND U19587 ( .A(n19141), .B(n19140), .Z(n19144) );
  XOR U19588 ( .A(n19143), .B(n19142), .Z(n19145) );
  NANDN U19589 ( .A(n19144), .B(n19145), .Z(n19147) );
  NAND U19590 ( .A(a[44]), .B(b[7]), .Z(n19523) );
  XNOR U19591 ( .A(n19145), .B(n19144), .Z(n19524) );
  NANDN U19592 ( .A(n19523), .B(n19524), .Z(n19146) );
  NAND U19593 ( .A(n19147), .B(n19146), .Z(n19148) );
  OR U19594 ( .A(n19149), .B(n19148), .Z(n19153) );
  XNOR U19595 ( .A(n19149), .B(n19148), .Z(n19527) );
  XOR U19596 ( .A(n19151), .B(n19150), .Z(n19528) );
  NANDN U19597 ( .A(n19527), .B(n19528), .Z(n19152) );
  NAND U19598 ( .A(n19153), .B(n19152), .Z(n19156) );
  XOR U19599 ( .A(n19155), .B(n19154), .Z(n19157) );
  NANDN U19600 ( .A(n19156), .B(n19157), .Z(n19159) );
  NAND U19601 ( .A(a[46]), .B(b[7]), .Z(n19535) );
  XNOR U19602 ( .A(n19157), .B(n19156), .Z(n19536) );
  NANDN U19603 ( .A(n19535), .B(n19536), .Z(n19158) );
  NAND U19604 ( .A(n19159), .B(n19158), .Z(n19160) );
  OR U19605 ( .A(n19161), .B(n19160), .Z(n19165) );
  XNOR U19606 ( .A(n19161), .B(n19160), .Z(n19539) );
  XOR U19607 ( .A(n19163), .B(n19162), .Z(n19540) );
  NANDN U19608 ( .A(n19539), .B(n19540), .Z(n19164) );
  NAND U19609 ( .A(n19165), .B(n19164), .Z(n19168) );
  XOR U19610 ( .A(n19167), .B(n19166), .Z(n19169) );
  NANDN U19611 ( .A(n19168), .B(n19169), .Z(n19171) );
  NAND U19612 ( .A(a[48]), .B(b[7]), .Z(n19547) );
  XNOR U19613 ( .A(n19169), .B(n19168), .Z(n19548) );
  NANDN U19614 ( .A(n19547), .B(n19548), .Z(n19170) );
  NAND U19615 ( .A(n19171), .B(n19170), .Z(n19172) );
  OR U19616 ( .A(n19173), .B(n19172), .Z(n19177) );
  XNOR U19617 ( .A(n19173), .B(n19172), .Z(n19551) );
  XOR U19618 ( .A(n19175), .B(n19174), .Z(n19552) );
  NANDN U19619 ( .A(n19551), .B(n19552), .Z(n19176) );
  NAND U19620 ( .A(n19177), .B(n19176), .Z(n19180) );
  XOR U19621 ( .A(n19179), .B(n19178), .Z(n19181) );
  NANDN U19622 ( .A(n19180), .B(n19181), .Z(n19183) );
  NAND U19623 ( .A(a[50]), .B(b[7]), .Z(n19559) );
  XNOR U19624 ( .A(n19181), .B(n19180), .Z(n19560) );
  NANDN U19625 ( .A(n19559), .B(n19560), .Z(n19182) );
  NAND U19626 ( .A(n19183), .B(n19182), .Z(n19184) );
  OR U19627 ( .A(n19185), .B(n19184), .Z(n19189) );
  XNOR U19628 ( .A(n19185), .B(n19184), .Z(n19563) );
  XOR U19629 ( .A(n19187), .B(n19186), .Z(n19564) );
  NANDN U19630 ( .A(n19563), .B(n19564), .Z(n19188) );
  NAND U19631 ( .A(n19189), .B(n19188), .Z(n19192) );
  XOR U19632 ( .A(n19191), .B(n19190), .Z(n19193) );
  NANDN U19633 ( .A(n19192), .B(n19193), .Z(n19195) );
  NAND U19634 ( .A(a[52]), .B(b[7]), .Z(n19571) );
  XNOR U19635 ( .A(n19193), .B(n19192), .Z(n19572) );
  NANDN U19636 ( .A(n19571), .B(n19572), .Z(n19194) );
  NAND U19637 ( .A(n19195), .B(n19194), .Z(n19196) );
  OR U19638 ( .A(n19197), .B(n19196), .Z(n19201) );
  XNOR U19639 ( .A(n19197), .B(n19196), .Z(n19575) );
  XOR U19640 ( .A(n19199), .B(n19198), .Z(n19576) );
  NANDN U19641 ( .A(n19575), .B(n19576), .Z(n19200) );
  NAND U19642 ( .A(n19201), .B(n19200), .Z(n19204) );
  XOR U19643 ( .A(n19203), .B(n19202), .Z(n19205) );
  NANDN U19644 ( .A(n19204), .B(n19205), .Z(n19207) );
  NAND U19645 ( .A(a[54]), .B(b[7]), .Z(n19583) );
  XNOR U19646 ( .A(n19205), .B(n19204), .Z(n19584) );
  NANDN U19647 ( .A(n19583), .B(n19584), .Z(n19206) );
  NAND U19648 ( .A(n19207), .B(n19206), .Z(n19210) );
  ANDN U19649 ( .B(b[7]), .A(n203), .Z(n19211) );
  OR U19650 ( .A(n19210), .B(n19211), .Z(n19213) );
  XOR U19651 ( .A(n19209), .B(n19208), .Z(n19588) );
  XOR U19652 ( .A(n19211), .B(n19210), .Z(n19587) );
  NANDN U19653 ( .A(n19588), .B(n19587), .Z(n19212) );
  NAND U19654 ( .A(n19213), .B(n19212), .Z(n19216) );
  XNOR U19655 ( .A(n19215), .B(n19214), .Z(n19217) );
  OR U19656 ( .A(n19216), .B(n19217), .Z(n19219) );
  XNOR U19657 ( .A(n19217), .B(n19216), .Z(n19594) );
  NAND U19658 ( .A(a[56]), .B(b[7]), .Z(n19593) );
  OR U19659 ( .A(n19594), .B(n19593), .Z(n19218) );
  NAND U19660 ( .A(n19219), .B(n19218), .Z(n19222) );
  ANDN U19661 ( .B(b[7]), .A(n205), .Z(n19223) );
  OR U19662 ( .A(n19222), .B(n19223), .Z(n19225) );
  XOR U19663 ( .A(n19223), .B(n19222), .Z(n19601) );
  NANDN U19664 ( .A(n19602), .B(n19601), .Z(n19224) );
  NAND U19665 ( .A(n19225), .B(n19224), .Z(n19229) );
  NAND U19666 ( .A(a[58]), .B(b[7]), .Z(n19228) );
  OR U19667 ( .A(n19229), .B(n19228), .Z(n19231) );
  XOR U19668 ( .A(n19227), .B(n19226), .Z(n19605) );
  XOR U19669 ( .A(n19229), .B(n19228), .Z(n19606) );
  NAND U19670 ( .A(n19605), .B(n19606), .Z(n19230) );
  NAND U19671 ( .A(n19231), .B(n19230), .Z(n19235) );
  XOR U19672 ( .A(n19233), .B(n19232), .Z(n19234) );
  NAND U19673 ( .A(n19235), .B(n19234), .Z(n19237) );
  XNOR U19674 ( .A(n19235), .B(n19234), .Z(n19612) );
  NAND U19675 ( .A(a[59]), .B(b[7]), .Z(n19611) );
  OR U19676 ( .A(n19612), .B(n19611), .Z(n19236) );
  NAND U19677 ( .A(n19237), .B(n19236), .Z(n19241) );
  NANDN U19678 ( .A(n19240), .B(n19241), .Z(n19243) );
  XNOR U19679 ( .A(n19239), .B(n19238), .Z(n19618) );
  XNOR U19680 ( .A(n19241), .B(n19240), .Z(n19617) );
  NANDN U19681 ( .A(n19618), .B(n19617), .Z(n19242) );
  NAND U19682 ( .A(n19243), .B(n19242), .Z(n19246) );
  XOR U19683 ( .A(n19245), .B(n19244), .Z(n19247) );
  AND U19684 ( .A(b[7]), .B(a[61]), .Z(n19624) );
  XOR U19685 ( .A(n19247), .B(n19246), .Z(n19623) );
  NAND U19686 ( .A(a[62]), .B(b[7]), .Z(n19250) );
  OR U19687 ( .A(n19251), .B(n19250), .Z(n19253) );
  XNOR U19688 ( .A(n19249), .B(n19248), .Z(n19630) );
  XOR U19689 ( .A(n19251), .B(n19250), .Z(n19629) );
  NANDN U19690 ( .A(n19630), .B(n19629), .Z(n19252) );
  NAND U19691 ( .A(n19253), .B(n19252), .Z(n19257) );
  XNOR U19692 ( .A(n19255), .B(n19254), .Z(n19256) );
  NAND U19693 ( .A(n19257), .B(n19256), .Z(n19259) );
  XNOR U19694 ( .A(n19257), .B(n19256), .Z(n19636) );
  NAND U19695 ( .A(a[63]), .B(b[7]), .Z(n19635) );
  OR U19696 ( .A(n19636), .B(n19635), .Z(n19258) );
  AND U19697 ( .A(n19259), .B(n19258), .Z(n19637) );
  OR U19698 ( .A(n19638), .B(n19637), .Z(n21933) );
  NANDN U19699 ( .A(n21932), .B(n21933), .Z(n21935) );
  NAND U19700 ( .A(a[60]), .B(b[6]), .Z(n19613) );
  ANDN U19701 ( .B(b[6]), .A(n203), .Z(n19582) );
  ANDN U19702 ( .B(b[6]), .A(n201), .Z(n19570) );
  ANDN U19703 ( .B(b[6]), .A(n199), .Z(n19558) );
  ANDN U19704 ( .B(b[6]), .A(n197), .Z(n19546) );
  ANDN U19705 ( .B(b[6]), .A(n195), .Z(n19534) );
  ANDN U19706 ( .B(b[6]), .A(n193), .Z(n19522) );
  ANDN U19707 ( .B(b[6]), .A(n191), .Z(n19510) );
  ANDN U19708 ( .B(b[6]), .A(n189), .Z(n19498) );
  ANDN U19709 ( .B(b[6]), .A(n187), .Z(n19486) );
  ANDN U19710 ( .B(b[6]), .A(n21772), .Z(n19474) );
  ANDN U19711 ( .B(b[6]), .A(n184), .Z(n19462) );
  ANDN U19712 ( .B(b[6]), .A(n21751), .Z(n19450) );
  ANDN U19713 ( .B(b[6]), .A(n21740), .Z(n19438) );
  ANDN U19714 ( .B(b[6]), .A(n21727), .Z(n19426) );
  ANDN U19715 ( .B(b[6]), .A(n21716), .Z(n19414) );
  ANDN U19716 ( .B(b[6]), .A(n21703), .Z(n19402) );
  ANDN U19717 ( .B(b[6]), .A(n21692), .Z(n19390) );
  ANDN U19718 ( .B(b[6]), .A(n21681), .Z(n19380) );
  ANDN U19719 ( .B(b[6]), .A(n21670), .Z(n19368) );
  NAND U19720 ( .A(a[18]), .B(b[6]), .Z(n19360) );
  NAND U19721 ( .A(a[17]), .B(b[6]), .Z(n19354) );
  ANDN U19722 ( .B(b[6]), .A(n172), .Z(n19344) );
  ANDN U19723 ( .B(b[6]), .A(n170), .Z(n19330) );
  ANDN U19724 ( .B(b[6]), .A(n21164), .Z(n19318) );
  NAND U19725 ( .A(a[10]), .B(b[6]), .Z(n19313) );
  XOR U19726 ( .A(n19261), .B(n19260), .Z(n19314) );
  NANDN U19727 ( .A(n19313), .B(n19314), .Z(n19316) );
  ANDN U19728 ( .B(b[6]), .A(n21615), .Z(n19308) );
  NAND U19729 ( .A(a[8]), .B(b[6]), .Z(n19303) );
  XOR U19730 ( .A(n19263), .B(n19262), .Z(n19304) );
  NANDN U19731 ( .A(n19303), .B(n19304), .Z(n19306) );
  ANDN U19732 ( .B(b[6]), .A(n166), .Z(n19298) );
  NAND U19733 ( .A(a[6]), .B(b[6]), .Z(n19293) );
  XOR U19734 ( .A(n19265), .B(n19264), .Z(n19294) );
  NANDN U19735 ( .A(n19293), .B(n19294), .Z(n19296) );
  ANDN U19736 ( .B(b[6]), .A(n21580), .Z(n19275) );
  NAND U19737 ( .A(b[7]), .B(a[1]), .Z(n19270) );
  NANDN U19738 ( .A(n19270), .B(a[0]), .Z(n19266) );
  XNOR U19739 ( .A(a[2]), .B(n19266), .Z(n19267) );
  NAND U19740 ( .A(b[6]), .B(n19267), .Z(n19662) );
  AND U19741 ( .A(a[1]), .B(b[7]), .Z(n19268) );
  XOR U19742 ( .A(n19269), .B(n19268), .Z(n19663) );
  OR U19743 ( .A(n19662), .B(n19663), .Z(n19274) );
  AND U19744 ( .A(b[6]), .B(a[0]), .Z(n20035) );
  NANDN U19745 ( .A(n19270), .B(n20035), .Z(n19272) );
  NAND U19746 ( .A(a[2]), .B(b[6]), .Z(n19271) );
  AND U19747 ( .A(n19272), .B(n19271), .Z(n19273) );
  ANDN U19748 ( .B(n19274), .A(n19273), .Z(n19276) );
  OR U19749 ( .A(n19275), .B(n19276), .Z(n19280) );
  XNOR U19750 ( .A(n19276), .B(n19275), .Z(n19667) );
  XNOR U19751 ( .A(n19278), .B(n19277), .Z(n19666) );
  OR U19752 ( .A(n19667), .B(n19666), .Z(n19279) );
  NAND U19753 ( .A(n19280), .B(n19279), .Z(n19284) );
  XOR U19754 ( .A(n19282), .B(n19281), .Z(n19283) );
  OR U19755 ( .A(n19284), .B(n19283), .Z(n19286) );
  NAND U19756 ( .A(a[4]), .B(b[6]), .Z(n19675) );
  XOR U19757 ( .A(n19284), .B(n19283), .Z(n19674) );
  NANDN U19758 ( .A(n19675), .B(n19674), .Z(n19285) );
  NAND U19759 ( .A(n19286), .B(n19285), .Z(n19287) );
  ANDN U19760 ( .B(b[6]), .A(n164), .Z(n19288) );
  OR U19761 ( .A(n19287), .B(n19288), .Z(n19292) );
  XNOR U19762 ( .A(n19288), .B(n19287), .Z(n19678) );
  OR U19763 ( .A(n19678), .B(n19679), .Z(n19291) );
  NAND U19764 ( .A(n19292), .B(n19291), .Z(n19686) );
  XNOR U19765 ( .A(n19294), .B(n19293), .Z(n19687) );
  NANDN U19766 ( .A(n19686), .B(n19687), .Z(n19295) );
  NAND U19767 ( .A(n19296), .B(n19295), .Z(n19297) );
  OR U19768 ( .A(n19298), .B(n19297), .Z(n19302) );
  XNOR U19769 ( .A(n19298), .B(n19297), .Z(n19649) );
  XOR U19770 ( .A(n19300), .B(n19299), .Z(n19650) );
  NANDN U19771 ( .A(n19649), .B(n19650), .Z(n19301) );
  NAND U19772 ( .A(n19302), .B(n19301), .Z(n19696) );
  XNOR U19773 ( .A(n19304), .B(n19303), .Z(n19697) );
  NANDN U19774 ( .A(n19696), .B(n19697), .Z(n19305) );
  NAND U19775 ( .A(n19306), .B(n19305), .Z(n19307) );
  OR U19776 ( .A(n19308), .B(n19307), .Z(n19312) );
  XNOR U19777 ( .A(n19308), .B(n19307), .Z(n19647) );
  XOR U19778 ( .A(n19310), .B(n19309), .Z(n19648) );
  NANDN U19779 ( .A(n19647), .B(n19648), .Z(n19311) );
  NAND U19780 ( .A(n19312), .B(n19311), .Z(n19706) );
  XNOR U19781 ( .A(n19314), .B(n19313), .Z(n19707) );
  NANDN U19782 ( .A(n19706), .B(n19707), .Z(n19315) );
  NAND U19783 ( .A(n19316), .B(n19315), .Z(n19317) );
  OR U19784 ( .A(n19318), .B(n19317), .Z(n19322) );
  XNOR U19785 ( .A(n19318), .B(n19317), .Z(n19710) );
  XOR U19786 ( .A(n19320), .B(n19319), .Z(n19711) );
  NANDN U19787 ( .A(n19710), .B(n19711), .Z(n19321) );
  NAND U19788 ( .A(n19322), .B(n19321), .Z(n19326) );
  NAND U19789 ( .A(a[12]), .B(b[6]), .Z(n19325) );
  OR U19790 ( .A(n19326), .B(n19325), .Z(n19328) );
  XOR U19791 ( .A(n19324), .B(n19323), .Z(n19717) );
  XOR U19792 ( .A(n19326), .B(n19325), .Z(n19716) );
  NAND U19793 ( .A(n19717), .B(n19716), .Z(n19327) );
  NAND U19794 ( .A(n19328), .B(n19327), .Z(n19329) );
  OR U19795 ( .A(n19330), .B(n19329), .Z(n19334) );
  XNOR U19796 ( .A(n19330), .B(n19329), .Z(n19722) );
  XOR U19797 ( .A(n19332), .B(n19331), .Z(n19723) );
  NANDN U19798 ( .A(n19722), .B(n19723), .Z(n19333) );
  NAND U19799 ( .A(n19334), .B(n19333), .Z(n19337) );
  XOR U19800 ( .A(n19336), .B(n19335), .Z(n19338) );
  NANDN U19801 ( .A(n19337), .B(n19338), .Z(n19340) );
  NAND U19802 ( .A(a[14]), .B(b[6]), .Z(n19730) );
  XNOR U19803 ( .A(n19338), .B(n19337), .Z(n19731) );
  NANDN U19804 ( .A(n19730), .B(n19731), .Z(n19339) );
  NAND U19805 ( .A(n19340), .B(n19339), .Z(n19343) );
  OR U19806 ( .A(n19344), .B(n19343), .Z(n19346) );
  XOR U19807 ( .A(n19344), .B(n19343), .Z(n19734) );
  NANDN U19808 ( .A(n19735), .B(n19734), .Z(n19345) );
  NAND U19809 ( .A(n19346), .B(n19345), .Z(n19349) );
  XOR U19810 ( .A(n19348), .B(n19347), .Z(n19350) );
  NANDN U19811 ( .A(n19349), .B(n19350), .Z(n19352) );
  NAND U19812 ( .A(a[16]), .B(b[6]), .Z(n19742) );
  XNOR U19813 ( .A(n19350), .B(n19349), .Z(n19743) );
  NANDN U19814 ( .A(n19742), .B(n19743), .Z(n19351) );
  NAND U19815 ( .A(n19352), .B(n19351), .Z(n19353) );
  NANDN U19816 ( .A(n19354), .B(n19353), .Z(n19358) );
  XNOR U19817 ( .A(n19356), .B(n19355), .Z(n19749) );
  NAND U19818 ( .A(n19748), .B(n19749), .Z(n19357) );
  NAND U19819 ( .A(n19358), .B(n19357), .Z(n19359) );
  NANDN U19820 ( .A(n19360), .B(n19359), .Z(n19364) );
  NAND U19821 ( .A(n19752), .B(n19753), .Z(n19363) );
  NAND U19822 ( .A(n19364), .B(n19363), .Z(n19367) );
  OR U19823 ( .A(n19368), .B(n19367), .Z(n19370) );
  XNOR U19824 ( .A(n19366), .B(n19365), .Z(n19646) );
  XOR U19825 ( .A(n19368), .B(n19367), .Z(n19645) );
  NANDN U19826 ( .A(n19646), .B(n19645), .Z(n19369) );
  NAND U19827 ( .A(n19370), .B(n19369), .Z(n19373) );
  XOR U19828 ( .A(n19372), .B(n19371), .Z(n19374) );
  NANDN U19829 ( .A(n19373), .B(n19374), .Z(n19376) );
  NAND U19830 ( .A(a[20]), .B(b[6]), .Z(n19764) );
  XNOR U19831 ( .A(n19374), .B(n19373), .Z(n19765) );
  NANDN U19832 ( .A(n19764), .B(n19765), .Z(n19375) );
  NAND U19833 ( .A(n19376), .B(n19375), .Z(n19379) );
  OR U19834 ( .A(n19380), .B(n19379), .Z(n19382) );
  XOR U19835 ( .A(n19378), .B(n19377), .Z(n19768) );
  XOR U19836 ( .A(n19380), .B(n19379), .Z(n19769) );
  NANDN U19837 ( .A(n19768), .B(n19769), .Z(n19381) );
  NAND U19838 ( .A(n19382), .B(n19381), .Z(n19385) );
  NANDN U19839 ( .A(n19385), .B(n19386), .Z(n19388) );
  NAND U19840 ( .A(a[22]), .B(b[6]), .Z(n19774) );
  XNOR U19841 ( .A(n19386), .B(n19385), .Z(n19775) );
  NANDN U19842 ( .A(n19774), .B(n19775), .Z(n19387) );
  NAND U19843 ( .A(n19388), .B(n19387), .Z(n19389) );
  OR U19844 ( .A(n19390), .B(n19389), .Z(n19394) );
  XNOR U19845 ( .A(n19390), .B(n19389), .Z(n19780) );
  XOR U19846 ( .A(n19392), .B(n19391), .Z(n19781) );
  NANDN U19847 ( .A(n19780), .B(n19781), .Z(n19393) );
  NAND U19848 ( .A(n19394), .B(n19393), .Z(n19397) );
  XOR U19849 ( .A(n19396), .B(n19395), .Z(n19398) );
  NANDN U19850 ( .A(n19397), .B(n19398), .Z(n19400) );
  NAND U19851 ( .A(a[24]), .B(b[6]), .Z(n19788) );
  XNOR U19852 ( .A(n19398), .B(n19397), .Z(n19789) );
  NANDN U19853 ( .A(n19788), .B(n19789), .Z(n19399) );
  NAND U19854 ( .A(n19400), .B(n19399), .Z(n19401) );
  OR U19855 ( .A(n19402), .B(n19401), .Z(n19406) );
  XNOR U19856 ( .A(n19402), .B(n19401), .Z(n19792) );
  XOR U19857 ( .A(n19404), .B(n19403), .Z(n19793) );
  NANDN U19858 ( .A(n19792), .B(n19793), .Z(n19405) );
  NAND U19859 ( .A(n19406), .B(n19405), .Z(n19409) );
  XOR U19860 ( .A(n19408), .B(n19407), .Z(n19410) );
  NANDN U19861 ( .A(n19409), .B(n19410), .Z(n19412) );
  NAND U19862 ( .A(a[26]), .B(b[6]), .Z(n19800) );
  XNOR U19863 ( .A(n19410), .B(n19409), .Z(n19801) );
  NANDN U19864 ( .A(n19800), .B(n19801), .Z(n19411) );
  NAND U19865 ( .A(n19412), .B(n19411), .Z(n19413) );
  OR U19866 ( .A(n19414), .B(n19413), .Z(n19418) );
  XNOR U19867 ( .A(n19414), .B(n19413), .Z(n19804) );
  XOR U19868 ( .A(n19416), .B(n19415), .Z(n19805) );
  NANDN U19869 ( .A(n19804), .B(n19805), .Z(n19417) );
  NAND U19870 ( .A(n19418), .B(n19417), .Z(n19421) );
  XOR U19871 ( .A(n19420), .B(n19419), .Z(n19422) );
  NANDN U19872 ( .A(n19421), .B(n19422), .Z(n19424) );
  NAND U19873 ( .A(a[28]), .B(b[6]), .Z(n19812) );
  XNOR U19874 ( .A(n19422), .B(n19421), .Z(n19813) );
  NANDN U19875 ( .A(n19812), .B(n19813), .Z(n19423) );
  NAND U19876 ( .A(n19424), .B(n19423), .Z(n19425) );
  OR U19877 ( .A(n19426), .B(n19425), .Z(n19430) );
  XNOR U19878 ( .A(n19426), .B(n19425), .Z(n19816) );
  XOR U19879 ( .A(n19428), .B(n19427), .Z(n19817) );
  NANDN U19880 ( .A(n19816), .B(n19817), .Z(n19429) );
  NAND U19881 ( .A(n19430), .B(n19429), .Z(n19433) );
  XOR U19882 ( .A(n19432), .B(n19431), .Z(n19434) );
  NANDN U19883 ( .A(n19433), .B(n19434), .Z(n19436) );
  NAND U19884 ( .A(a[30]), .B(b[6]), .Z(n19824) );
  XNOR U19885 ( .A(n19434), .B(n19433), .Z(n19825) );
  NANDN U19886 ( .A(n19824), .B(n19825), .Z(n19435) );
  NAND U19887 ( .A(n19436), .B(n19435), .Z(n19437) );
  OR U19888 ( .A(n19438), .B(n19437), .Z(n19442) );
  XNOR U19889 ( .A(n19438), .B(n19437), .Z(n19828) );
  XOR U19890 ( .A(n19440), .B(n19439), .Z(n19829) );
  NANDN U19891 ( .A(n19828), .B(n19829), .Z(n19441) );
  NAND U19892 ( .A(n19442), .B(n19441), .Z(n19445) );
  XOR U19893 ( .A(n19444), .B(n19443), .Z(n19446) );
  NANDN U19894 ( .A(n19445), .B(n19446), .Z(n19448) );
  NAND U19895 ( .A(a[32]), .B(b[6]), .Z(n19836) );
  XNOR U19896 ( .A(n19446), .B(n19445), .Z(n19837) );
  NANDN U19897 ( .A(n19836), .B(n19837), .Z(n19447) );
  NAND U19898 ( .A(n19448), .B(n19447), .Z(n19449) );
  OR U19899 ( .A(n19450), .B(n19449), .Z(n19454) );
  XNOR U19900 ( .A(n19450), .B(n19449), .Z(n19840) );
  XOR U19901 ( .A(n19452), .B(n19451), .Z(n19841) );
  NANDN U19902 ( .A(n19840), .B(n19841), .Z(n19453) );
  NAND U19903 ( .A(n19454), .B(n19453), .Z(n19457) );
  XOR U19904 ( .A(n19456), .B(n19455), .Z(n19458) );
  NANDN U19905 ( .A(n19457), .B(n19458), .Z(n19460) );
  NAND U19906 ( .A(a[34]), .B(b[6]), .Z(n19848) );
  XNOR U19907 ( .A(n19458), .B(n19457), .Z(n19849) );
  NANDN U19908 ( .A(n19848), .B(n19849), .Z(n19459) );
  NAND U19909 ( .A(n19460), .B(n19459), .Z(n19461) );
  OR U19910 ( .A(n19462), .B(n19461), .Z(n19466) );
  XNOR U19911 ( .A(n19462), .B(n19461), .Z(n19852) );
  XOR U19912 ( .A(n19464), .B(n19463), .Z(n19853) );
  NANDN U19913 ( .A(n19852), .B(n19853), .Z(n19465) );
  NAND U19914 ( .A(n19466), .B(n19465), .Z(n19469) );
  XOR U19915 ( .A(n19468), .B(n19467), .Z(n19470) );
  NANDN U19916 ( .A(n19469), .B(n19470), .Z(n19472) );
  NAND U19917 ( .A(a[36]), .B(b[6]), .Z(n19860) );
  XNOR U19918 ( .A(n19470), .B(n19469), .Z(n19861) );
  NANDN U19919 ( .A(n19860), .B(n19861), .Z(n19471) );
  NAND U19920 ( .A(n19472), .B(n19471), .Z(n19473) );
  OR U19921 ( .A(n19474), .B(n19473), .Z(n19478) );
  XNOR U19922 ( .A(n19474), .B(n19473), .Z(n19864) );
  XOR U19923 ( .A(n19476), .B(n19475), .Z(n19865) );
  NANDN U19924 ( .A(n19864), .B(n19865), .Z(n19477) );
  NAND U19925 ( .A(n19478), .B(n19477), .Z(n19481) );
  XOR U19926 ( .A(n19480), .B(n19479), .Z(n19482) );
  NANDN U19927 ( .A(n19481), .B(n19482), .Z(n19484) );
  NAND U19928 ( .A(a[38]), .B(b[6]), .Z(n19872) );
  XNOR U19929 ( .A(n19482), .B(n19481), .Z(n19873) );
  NANDN U19930 ( .A(n19872), .B(n19873), .Z(n19483) );
  NAND U19931 ( .A(n19484), .B(n19483), .Z(n19485) );
  OR U19932 ( .A(n19486), .B(n19485), .Z(n19490) );
  XNOR U19933 ( .A(n19486), .B(n19485), .Z(n19876) );
  XOR U19934 ( .A(n19488), .B(n19487), .Z(n19877) );
  NANDN U19935 ( .A(n19876), .B(n19877), .Z(n19489) );
  NAND U19936 ( .A(n19490), .B(n19489), .Z(n19493) );
  XOR U19937 ( .A(n19492), .B(n19491), .Z(n19494) );
  NANDN U19938 ( .A(n19493), .B(n19494), .Z(n19496) );
  NAND U19939 ( .A(a[40]), .B(b[6]), .Z(n19884) );
  XNOR U19940 ( .A(n19494), .B(n19493), .Z(n19885) );
  NANDN U19941 ( .A(n19884), .B(n19885), .Z(n19495) );
  NAND U19942 ( .A(n19496), .B(n19495), .Z(n19497) );
  OR U19943 ( .A(n19498), .B(n19497), .Z(n19502) );
  XNOR U19944 ( .A(n19498), .B(n19497), .Z(n19888) );
  XOR U19945 ( .A(n19500), .B(n19499), .Z(n19889) );
  NANDN U19946 ( .A(n19888), .B(n19889), .Z(n19501) );
  NAND U19947 ( .A(n19502), .B(n19501), .Z(n19505) );
  XOR U19948 ( .A(n19504), .B(n19503), .Z(n19506) );
  NANDN U19949 ( .A(n19505), .B(n19506), .Z(n19508) );
  NAND U19950 ( .A(a[42]), .B(b[6]), .Z(n19896) );
  XNOR U19951 ( .A(n19506), .B(n19505), .Z(n19897) );
  NANDN U19952 ( .A(n19896), .B(n19897), .Z(n19507) );
  NAND U19953 ( .A(n19508), .B(n19507), .Z(n19509) );
  OR U19954 ( .A(n19510), .B(n19509), .Z(n19514) );
  XNOR U19955 ( .A(n19510), .B(n19509), .Z(n19900) );
  XOR U19956 ( .A(n19512), .B(n19511), .Z(n19901) );
  NANDN U19957 ( .A(n19900), .B(n19901), .Z(n19513) );
  NAND U19958 ( .A(n19514), .B(n19513), .Z(n19517) );
  XOR U19959 ( .A(n19516), .B(n19515), .Z(n19518) );
  NANDN U19960 ( .A(n19517), .B(n19518), .Z(n19520) );
  NAND U19961 ( .A(a[44]), .B(b[6]), .Z(n19908) );
  XNOR U19962 ( .A(n19518), .B(n19517), .Z(n19909) );
  NANDN U19963 ( .A(n19908), .B(n19909), .Z(n19519) );
  NAND U19964 ( .A(n19520), .B(n19519), .Z(n19521) );
  OR U19965 ( .A(n19522), .B(n19521), .Z(n19526) );
  XNOR U19966 ( .A(n19522), .B(n19521), .Z(n19912) );
  XOR U19967 ( .A(n19524), .B(n19523), .Z(n19913) );
  NANDN U19968 ( .A(n19912), .B(n19913), .Z(n19525) );
  NAND U19969 ( .A(n19526), .B(n19525), .Z(n19529) );
  XOR U19970 ( .A(n19528), .B(n19527), .Z(n19530) );
  NANDN U19971 ( .A(n19529), .B(n19530), .Z(n19532) );
  NAND U19972 ( .A(a[46]), .B(b[6]), .Z(n19920) );
  XNOR U19973 ( .A(n19530), .B(n19529), .Z(n19921) );
  NANDN U19974 ( .A(n19920), .B(n19921), .Z(n19531) );
  NAND U19975 ( .A(n19532), .B(n19531), .Z(n19533) );
  OR U19976 ( .A(n19534), .B(n19533), .Z(n19538) );
  XNOR U19977 ( .A(n19534), .B(n19533), .Z(n19924) );
  XOR U19978 ( .A(n19536), .B(n19535), .Z(n19925) );
  NANDN U19979 ( .A(n19924), .B(n19925), .Z(n19537) );
  NAND U19980 ( .A(n19538), .B(n19537), .Z(n19541) );
  XOR U19981 ( .A(n19540), .B(n19539), .Z(n19542) );
  NANDN U19982 ( .A(n19541), .B(n19542), .Z(n19544) );
  NAND U19983 ( .A(a[48]), .B(b[6]), .Z(n19932) );
  XNOR U19984 ( .A(n19542), .B(n19541), .Z(n19933) );
  NANDN U19985 ( .A(n19932), .B(n19933), .Z(n19543) );
  NAND U19986 ( .A(n19544), .B(n19543), .Z(n19545) );
  OR U19987 ( .A(n19546), .B(n19545), .Z(n19550) );
  XNOR U19988 ( .A(n19546), .B(n19545), .Z(n19936) );
  XOR U19989 ( .A(n19548), .B(n19547), .Z(n19937) );
  NANDN U19990 ( .A(n19936), .B(n19937), .Z(n19549) );
  NAND U19991 ( .A(n19550), .B(n19549), .Z(n19553) );
  XOR U19992 ( .A(n19552), .B(n19551), .Z(n19554) );
  NANDN U19993 ( .A(n19553), .B(n19554), .Z(n19556) );
  NAND U19994 ( .A(a[50]), .B(b[6]), .Z(n19944) );
  XNOR U19995 ( .A(n19554), .B(n19553), .Z(n19945) );
  NANDN U19996 ( .A(n19944), .B(n19945), .Z(n19555) );
  NAND U19997 ( .A(n19556), .B(n19555), .Z(n19557) );
  OR U19998 ( .A(n19558), .B(n19557), .Z(n19562) );
  XNOR U19999 ( .A(n19558), .B(n19557), .Z(n19948) );
  XOR U20000 ( .A(n19560), .B(n19559), .Z(n19949) );
  NANDN U20001 ( .A(n19948), .B(n19949), .Z(n19561) );
  NAND U20002 ( .A(n19562), .B(n19561), .Z(n19565) );
  XOR U20003 ( .A(n19564), .B(n19563), .Z(n19566) );
  NANDN U20004 ( .A(n19565), .B(n19566), .Z(n19568) );
  NAND U20005 ( .A(a[52]), .B(b[6]), .Z(n19956) );
  XNOR U20006 ( .A(n19566), .B(n19565), .Z(n19957) );
  NANDN U20007 ( .A(n19956), .B(n19957), .Z(n19567) );
  NAND U20008 ( .A(n19568), .B(n19567), .Z(n19569) );
  OR U20009 ( .A(n19570), .B(n19569), .Z(n19574) );
  XNOR U20010 ( .A(n19570), .B(n19569), .Z(n19960) );
  XOR U20011 ( .A(n19572), .B(n19571), .Z(n19961) );
  NANDN U20012 ( .A(n19960), .B(n19961), .Z(n19573) );
  NAND U20013 ( .A(n19574), .B(n19573), .Z(n19577) );
  XOR U20014 ( .A(n19576), .B(n19575), .Z(n19578) );
  NANDN U20015 ( .A(n19577), .B(n19578), .Z(n19580) );
  NAND U20016 ( .A(a[54]), .B(b[6]), .Z(n19968) );
  XNOR U20017 ( .A(n19578), .B(n19577), .Z(n19969) );
  NANDN U20018 ( .A(n19968), .B(n19969), .Z(n19579) );
  NAND U20019 ( .A(n19580), .B(n19579), .Z(n19581) );
  OR U20020 ( .A(n19582), .B(n19581), .Z(n19586) );
  XNOR U20021 ( .A(n19582), .B(n19581), .Z(n19972) );
  XOR U20022 ( .A(n19584), .B(n19583), .Z(n19973) );
  NANDN U20023 ( .A(n19972), .B(n19973), .Z(n19585) );
  NAND U20024 ( .A(n19586), .B(n19585), .Z(n19589) );
  XNOR U20025 ( .A(n19588), .B(n19587), .Z(n19590) );
  OR U20026 ( .A(n19589), .B(n19590), .Z(n19592) );
  XNOR U20027 ( .A(n19590), .B(n19589), .Z(n19979) );
  NAND U20028 ( .A(a[56]), .B(b[6]), .Z(n19978) );
  OR U20029 ( .A(n19979), .B(n19978), .Z(n19591) );
  NAND U20030 ( .A(n19592), .B(n19591), .Z(n19595) );
  ANDN U20031 ( .B(b[6]), .A(n205), .Z(n19596) );
  OR U20032 ( .A(n19595), .B(n19596), .Z(n19598) );
  XOR U20033 ( .A(n19594), .B(n19593), .Z(n19985) );
  XOR U20034 ( .A(n19596), .B(n19595), .Z(n19984) );
  NANDN U20035 ( .A(n19985), .B(n19984), .Z(n19597) );
  NAND U20036 ( .A(n19598), .B(n19597), .Z(n19600) );
  AND U20037 ( .A(b[6]), .B(a[58]), .Z(n19599) );
  NANDN U20038 ( .A(n19600), .B(n19599), .Z(n19604) );
  XNOR U20039 ( .A(n19600), .B(n19599), .Z(n19990) );
  NAND U20040 ( .A(n19990), .B(n19991), .Z(n19603) );
  NAND U20041 ( .A(n19604), .B(n19603), .Z(n19608) );
  XOR U20042 ( .A(n19606), .B(n19605), .Z(n19607) );
  NAND U20043 ( .A(n19608), .B(n19607), .Z(n19610) );
  XNOR U20044 ( .A(n19608), .B(n19607), .Z(n19997) );
  NAND U20045 ( .A(a[59]), .B(b[6]), .Z(n19996) );
  OR U20046 ( .A(n19997), .B(n19996), .Z(n19609) );
  NAND U20047 ( .A(n19610), .B(n19609), .Z(n19614) );
  NANDN U20048 ( .A(n19613), .B(n19614), .Z(n19616) );
  XOR U20049 ( .A(n19612), .B(n19611), .Z(n20002) );
  XNOR U20050 ( .A(n19614), .B(n19613), .Z(n20003) );
  NAND U20051 ( .A(n20002), .B(n20003), .Z(n19615) );
  NAND U20052 ( .A(n19616), .B(n19615), .Z(n19619) );
  AND U20053 ( .A(b[6]), .B(a[61]), .Z(n19620) );
  OR U20054 ( .A(n19619), .B(n19620), .Z(n19622) );
  XNOR U20055 ( .A(n19618), .B(n19617), .Z(n20009) );
  XOR U20056 ( .A(n19620), .B(n19619), .Z(n20008) );
  NANDN U20057 ( .A(n20009), .B(n20008), .Z(n19621) );
  NAND U20058 ( .A(n19622), .B(n19621), .Z(n19626) );
  NAND U20059 ( .A(a[62]), .B(b[6]), .Z(n19625) );
  OR U20060 ( .A(n19626), .B(n19625), .Z(n19628) );
  XOR U20061 ( .A(n19624), .B(n19623), .Z(n20015) );
  XOR U20062 ( .A(n19626), .B(n19625), .Z(n20014) );
  NAND U20063 ( .A(n20015), .B(n20014), .Z(n19627) );
  NAND U20064 ( .A(n19628), .B(n19627), .Z(n19631) );
  AND U20065 ( .A(b[6]), .B(a[63]), .Z(n19632) );
  OR U20066 ( .A(n19631), .B(n19632), .Z(n19634) );
  XNOR U20067 ( .A(n19630), .B(n19629), .Z(n19644) );
  XOR U20068 ( .A(n19632), .B(n19631), .Z(n19643) );
  NANDN U20069 ( .A(n19644), .B(n19643), .Z(n19633) );
  NAND U20070 ( .A(n19634), .B(n19633), .Z(n19641) );
  XOR U20071 ( .A(n19636), .B(n19635), .Z(n19642) );
  NANDN U20072 ( .A(n19641), .B(n19642), .Z(n19639) );
  XOR U20073 ( .A(n19638), .B(n19637), .Z(n19640) );
  NANDN U20074 ( .A(n19639), .B(n19640), .Z(n21931) );
  XOR U20075 ( .A(n19640), .B(n19639), .Z(n24112) );
  XNOR U20076 ( .A(n19642), .B(n19641), .Z(n21926) );
  XNOR U20077 ( .A(n19644), .B(n19643), .Z(n20021) );
  NAND U20078 ( .A(a[62]), .B(b[5]), .Z(n20010) );
  ANDN U20079 ( .B(b[5]), .A(n203), .Z(n19967) );
  ANDN U20080 ( .B(b[5]), .A(n201), .Z(n19955) );
  ANDN U20081 ( .B(b[5]), .A(n199), .Z(n19943) );
  ANDN U20082 ( .B(b[5]), .A(n197), .Z(n19931) );
  ANDN U20083 ( .B(b[5]), .A(n195), .Z(n19919) );
  ANDN U20084 ( .B(b[5]), .A(n193), .Z(n19907) );
  ANDN U20085 ( .B(b[5]), .A(n191), .Z(n19895) );
  ANDN U20086 ( .B(b[5]), .A(n189), .Z(n19883) );
  ANDN U20087 ( .B(b[5]), .A(n187), .Z(n19871) );
  ANDN U20088 ( .B(b[5]), .A(n21772), .Z(n19859) );
  ANDN U20089 ( .B(b[5]), .A(n184), .Z(n19847) );
  ANDN U20090 ( .B(b[5]), .A(n21751), .Z(n19835) );
  ANDN U20091 ( .B(b[5]), .A(n21740), .Z(n19823) );
  ANDN U20092 ( .B(b[5]), .A(n21727), .Z(n19811) );
  ANDN U20093 ( .B(b[5]), .A(n21716), .Z(n19799) );
  ANDN U20094 ( .B(b[5]), .A(n21703), .Z(n19787) );
  ANDN U20095 ( .B(b[5]), .A(n21692), .Z(n19777) );
  ANDN U20096 ( .B(b[5]), .A(n21681), .Z(n19763) );
  XOR U20097 ( .A(n19646), .B(n19645), .Z(n19758) );
  ANDN U20098 ( .B(b[5]), .A(n21670), .Z(n19755) );
  NAND U20099 ( .A(a[18]), .B(b[5]), .Z(n19747) );
  NAND U20100 ( .A(a[17]), .B(b[5]), .Z(n19741) );
  ANDN U20101 ( .B(b[5]), .A(n172), .Z(n19729) );
  ANDN U20102 ( .B(b[5]), .A(n170), .Z(n19719) );
  ANDN U20103 ( .B(b[5]), .A(n21164), .Z(n19705) );
  NAND U20104 ( .A(a[10]), .B(b[5]), .Z(n19700) );
  XOR U20105 ( .A(n19648), .B(n19647), .Z(n19701) );
  NANDN U20106 ( .A(n19700), .B(n19701), .Z(n19703) );
  ANDN U20107 ( .B(b[5]), .A(n21615), .Z(n19695) );
  NAND U20108 ( .A(a[8]), .B(b[5]), .Z(n19690) );
  XOR U20109 ( .A(n19650), .B(n19649), .Z(n19691) );
  NANDN U20110 ( .A(n19690), .B(n19691), .Z(n19693) );
  ANDN U20111 ( .B(b[5]), .A(n166), .Z(n19685) );
  ANDN U20112 ( .B(b[5]), .A(n21580), .Z(n19660) );
  NAND U20113 ( .A(b[6]), .B(a[1]), .Z(n19655) );
  NANDN U20114 ( .A(n19655), .B(a[0]), .Z(n19651) );
  XNOR U20115 ( .A(a[2]), .B(n19651), .Z(n19652) );
  NAND U20116 ( .A(b[5]), .B(n19652), .Z(n20043) );
  AND U20117 ( .A(a[1]), .B(b[6]), .Z(n19653) );
  XOR U20118 ( .A(n19654), .B(n19653), .Z(n20044) );
  OR U20119 ( .A(n20043), .B(n20044), .Z(n19659) );
  AND U20120 ( .A(b[5]), .B(a[0]), .Z(n20415) );
  NANDN U20121 ( .A(n19655), .B(n20415), .Z(n19657) );
  NAND U20122 ( .A(a[2]), .B(b[5]), .Z(n19656) );
  AND U20123 ( .A(n19657), .B(n19656), .Z(n19658) );
  ANDN U20124 ( .B(n19659), .A(n19658), .Z(n19661) );
  OR U20125 ( .A(n19660), .B(n19661), .Z(n19665) );
  XNOR U20126 ( .A(n19661), .B(n19660), .Z(n20048) );
  XNOR U20127 ( .A(n19663), .B(n19662), .Z(n20047) );
  OR U20128 ( .A(n20048), .B(n20047), .Z(n19664) );
  NAND U20129 ( .A(n19665), .B(n19664), .Z(n19669) );
  XOR U20130 ( .A(n19667), .B(n19666), .Z(n19668) );
  OR U20131 ( .A(n19669), .B(n19668), .Z(n19671) );
  NAND U20132 ( .A(a[4]), .B(b[5]), .Z(n20056) );
  XOR U20133 ( .A(n19669), .B(n19668), .Z(n20055) );
  NANDN U20134 ( .A(n20056), .B(n20055), .Z(n19670) );
  NAND U20135 ( .A(n19671), .B(n19670), .Z(n19672) );
  ANDN U20136 ( .B(b[5]), .A(n164), .Z(n19673) );
  OR U20137 ( .A(n19672), .B(n19673), .Z(n19677) );
  XNOR U20138 ( .A(n19673), .B(n19672), .Z(n20059) );
  OR U20139 ( .A(n20059), .B(n20060), .Z(n19676) );
  AND U20140 ( .A(n19677), .B(n19676), .Z(n19681) );
  XOR U20141 ( .A(n19679), .B(n19678), .Z(n19680) );
  NANDN U20142 ( .A(n19681), .B(n19680), .Z(n19683) );
  XOR U20143 ( .A(n19681), .B(n19680), .Z(n20068) );
  ANDN U20144 ( .B(b[5]), .A(n165), .Z(n20067) );
  OR U20145 ( .A(n20068), .B(n20067), .Z(n19682) );
  NAND U20146 ( .A(n19683), .B(n19682), .Z(n19684) );
  NANDN U20147 ( .A(n19685), .B(n19684), .Z(n19689) );
  XOR U20148 ( .A(n19687), .B(n19686), .Z(n20071) );
  NANDN U20149 ( .A(n20072), .B(n20071), .Z(n19688) );
  NAND U20150 ( .A(n19689), .B(n19688), .Z(n20079) );
  XNOR U20151 ( .A(n19691), .B(n19690), .Z(n20080) );
  NANDN U20152 ( .A(n20079), .B(n20080), .Z(n19692) );
  NAND U20153 ( .A(n19693), .B(n19692), .Z(n19694) );
  OR U20154 ( .A(n19695), .B(n19694), .Z(n19699) );
  XNOR U20155 ( .A(n19695), .B(n19694), .Z(n20030) );
  XOR U20156 ( .A(n19697), .B(n19696), .Z(n20031) );
  NANDN U20157 ( .A(n20030), .B(n20031), .Z(n19698) );
  NAND U20158 ( .A(n19699), .B(n19698), .Z(n20089) );
  XNOR U20159 ( .A(n19701), .B(n19700), .Z(n20090) );
  NANDN U20160 ( .A(n20089), .B(n20090), .Z(n19702) );
  NAND U20161 ( .A(n19703), .B(n19702), .Z(n19704) );
  OR U20162 ( .A(n19705), .B(n19704), .Z(n19709) );
  XNOR U20163 ( .A(n19705), .B(n19704), .Z(n20026) );
  XOR U20164 ( .A(n19707), .B(n19706), .Z(n20027) );
  NANDN U20165 ( .A(n20026), .B(n20027), .Z(n19708) );
  NAND U20166 ( .A(n19709), .B(n19708), .Z(n19712) );
  XOR U20167 ( .A(n19711), .B(n19710), .Z(n19713) );
  NANDN U20168 ( .A(n19712), .B(n19713), .Z(n19715) );
  NAND U20169 ( .A(a[12]), .B(b[5]), .Z(n20097) );
  XNOR U20170 ( .A(n19713), .B(n19712), .Z(n20098) );
  NANDN U20171 ( .A(n20097), .B(n20098), .Z(n19714) );
  NAND U20172 ( .A(n19715), .B(n19714), .Z(n19718) );
  OR U20173 ( .A(n19719), .B(n19718), .Z(n19721) );
  XOR U20174 ( .A(n19717), .B(n19716), .Z(n20102) );
  XOR U20175 ( .A(n19719), .B(n19718), .Z(n20101) );
  NANDN U20176 ( .A(n20102), .B(n20101), .Z(n19720) );
  NAND U20177 ( .A(n19721), .B(n19720), .Z(n19724) );
  XOR U20178 ( .A(n19723), .B(n19722), .Z(n19725) );
  NANDN U20179 ( .A(n19724), .B(n19725), .Z(n19727) );
  NAND U20180 ( .A(a[14]), .B(b[5]), .Z(n20107) );
  XNOR U20181 ( .A(n19725), .B(n19724), .Z(n20108) );
  NANDN U20182 ( .A(n20107), .B(n20108), .Z(n19726) );
  NAND U20183 ( .A(n19727), .B(n19726), .Z(n19728) );
  OR U20184 ( .A(n19729), .B(n19728), .Z(n19733) );
  XNOR U20185 ( .A(n19729), .B(n19728), .Z(n20113) );
  XOR U20186 ( .A(n19731), .B(n19730), .Z(n20114) );
  NANDN U20187 ( .A(n20113), .B(n20114), .Z(n19732) );
  NAND U20188 ( .A(n19733), .B(n19732), .Z(n19736) );
  NANDN U20189 ( .A(n19736), .B(n19737), .Z(n19739) );
  NAND U20190 ( .A(a[16]), .B(b[5]), .Z(n20121) );
  XNOR U20191 ( .A(n19737), .B(n19736), .Z(n20122) );
  NANDN U20192 ( .A(n20121), .B(n20122), .Z(n19738) );
  NAND U20193 ( .A(n19739), .B(n19738), .Z(n19740) );
  NANDN U20194 ( .A(n19741), .B(n19740), .Z(n19745) );
  XNOR U20195 ( .A(n19743), .B(n19742), .Z(n20128) );
  NAND U20196 ( .A(n20127), .B(n20128), .Z(n19744) );
  NAND U20197 ( .A(n19745), .B(n19744), .Z(n19746) );
  NANDN U20198 ( .A(n19747), .B(n19746), .Z(n19751) );
  NAND U20199 ( .A(n20131), .B(n20132), .Z(n19750) );
  NAND U20200 ( .A(n19751), .B(n19750), .Z(n19754) );
  OR U20201 ( .A(n19755), .B(n19754), .Z(n19757) );
  XOR U20202 ( .A(n19755), .B(n19754), .Z(n20137) );
  NANDN U20203 ( .A(n20138), .B(n20137), .Z(n19756) );
  NAND U20204 ( .A(n19757), .B(n19756), .Z(n19759) );
  NANDN U20205 ( .A(n19758), .B(n19759), .Z(n19761) );
  ANDN U20206 ( .B(b[5]), .A(n176), .Z(n20144) );
  XOR U20207 ( .A(n19759), .B(n19758), .Z(n20143) );
  OR U20208 ( .A(n20144), .B(n20143), .Z(n19760) );
  AND U20209 ( .A(n19761), .B(n19760), .Z(n19762) );
  OR U20210 ( .A(n19763), .B(n19762), .Z(n19767) );
  XNOR U20211 ( .A(n19763), .B(n19762), .Z(n20149) );
  XOR U20212 ( .A(n19765), .B(n19764), .Z(n20150) );
  NANDN U20213 ( .A(n20149), .B(n20150), .Z(n19766) );
  NAND U20214 ( .A(n19767), .B(n19766), .Z(n19771) );
  XOR U20215 ( .A(n19769), .B(n19768), .Z(n19770) );
  NANDN U20216 ( .A(n19771), .B(n19770), .Z(n19773) );
  NAND U20217 ( .A(a[22]), .B(b[5]), .Z(n20155) );
  NANDN U20218 ( .A(n20155), .B(n20156), .Z(n19772) );
  NAND U20219 ( .A(n19773), .B(n19772), .Z(n19776) );
  OR U20220 ( .A(n19777), .B(n19776), .Z(n19779) );
  XOR U20221 ( .A(n19775), .B(n19774), .Z(n20025) );
  XOR U20222 ( .A(n19777), .B(n19776), .Z(n20024) );
  NAND U20223 ( .A(n20025), .B(n20024), .Z(n19778) );
  NAND U20224 ( .A(n19779), .B(n19778), .Z(n19782) );
  XOR U20225 ( .A(n19781), .B(n19780), .Z(n19783) );
  NANDN U20226 ( .A(n19782), .B(n19783), .Z(n19785) );
  NAND U20227 ( .A(a[24]), .B(b[5]), .Z(n20167) );
  XNOR U20228 ( .A(n19783), .B(n19782), .Z(n20168) );
  NANDN U20229 ( .A(n20167), .B(n20168), .Z(n19784) );
  NAND U20230 ( .A(n19785), .B(n19784), .Z(n19786) );
  OR U20231 ( .A(n19787), .B(n19786), .Z(n19791) );
  XNOR U20232 ( .A(n19787), .B(n19786), .Z(n20171) );
  XOR U20233 ( .A(n19789), .B(n19788), .Z(n20172) );
  NANDN U20234 ( .A(n20171), .B(n20172), .Z(n19790) );
  NAND U20235 ( .A(n19791), .B(n19790), .Z(n19794) );
  XOR U20236 ( .A(n19793), .B(n19792), .Z(n19795) );
  NANDN U20237 ( .A(n19794), .B(n19795), .Z(n19797) );
  NAND U20238 ( .A(a[26]), .B(b[5]), .Z(n20179) );
  XNOR U20239 ( .A(n19795), .B(n19794), .Z(n20180) );
  NANDN U20240 ( .A(n20179), .B(n20180), .Z(n19796) );
  NAND U20241 ( .A(n19797), .B(n19796), .Z(n19798) );
  OR U20242 ( .A(n19799), .B(n19798), .Z(n19803) );
  XNOR U20243 ( .A(n19799), .B(n19798), .Z(n20183) );
  XOR U20244 ( .A(n19801), .B(n19800), .Z(n20184) );
  NANDN U20245 ( .A(n20183), .B(n20184), .Z(n19802) );
  NAND U20246 ( .A(n19803), .B(n19802), .Z(n19806) );
  XOR U20247 ( .A(n19805), .B(n19804), .Z(n19807) );
  NANDN U20248 ( .A(n19806), .B(n19807), .Z(n19809) );
  NAND U20249 ( .A(a[28]), .B(b[5]), .Z(n20191) );
  XNOR U20250 ( .A(n19807), .B(n19806), .Z(n20192) );
  NANDN U20251 ( .A(n20191), .B(n20192), .Z(n19808) );
  NAND U20252 ( .A(n19809), .B(n19808), .Z(n19810) );
  OR U20253 ( .A(n19811), .B(n19810), .Z(n19815) );
  XNOR U20254 ( .A(n19811), .B(n19810), .Z(n20195) );
  XOR U20255 ( .A(n19813), .B(n19812), .Z(n20196) );
  NANDN U20256 ( .A(n20195), .B(n20196), .Z(n19814) );
  NAND U20257 ( .A(n19815), .B(n19814), .Z(n19818) );
  XOR U20258 ( .A(n19817), .B(n19816), .Z(n19819) );
  NANDN U20259 ( .A(n19818), .B(n19819), .Z(n19821) );
  NAND U20260 ( .A(a[30]), .B(b[5]), .Z(n20203) );
  XNOR U20261 ( .A(n19819), .B(n19818), .Z(n20204) );
  NANDN U20262 ( .A(n20203), .B(n20204), .Z(n19820) );
  NAND U20263 ( .A(n19821), .B(n19820), .Z(n19822) );
  OR U20264 ( .A(n19823), .B(n19822), .Z(n19827) );
  XNOR U20265 ( .A(n19823), .B(n19822), .Z(n20207) );
  XOR U20266 ( .A(n19825), .B(n19824), .Z(n20208) );
  NANDN U20267 ( .A(n20207), .B(n20208), .Z(n19826) );
  NAND U20268 ( .A(n19827), .B(n19826), .Z(n19830) );
  XOR U20269 ( .A(n19829), .B(n19828), .Z(n19831) );
  NANDN U20270 ( .A(n19830), .B(n19831), .Z(n19833) );
  NAND U20271 ( .A(a[32]), .B(b[5]), .Z(n20215) );
  XNOR U20272 ( .A(n19831), .B(n19830), .Z(n20216) );
  NANDN U20273 ( .A(n20215), .B(n20216), .Z(n19832) );
  NAND U20274 ( .A(n19833), .B(n19832), .Z(n19834) );
  OR U20275 ( .A(n19835), .B(n19834), .Z(n19839) );
  XNOR U20276 ( .A(n19835), .B(n19834), .Z(n20219) );
  XOR U20277 ( .A(n19837), .B(n19836), .Z(n20220) );
  NANDN U20278 ( .A(n20219), .B(n20220), .Z(n19838) );
  NAND U20279 ( .A(n19839), .B(n19838), .Z(n19842) );
  XOR U20280 ( .A(n19841), .B(n19840), .Z(n19843) );
  NANDN U20281 ( .A(n19842), .B(n19843), .Z(n19845) );
  NAND U20282 ( .A(a[34]), .B(b[5]), .Z(n20227) );
  XNOR U20283 ( .A(n19843), .B(n19842), .Z(n20228) );
  NANDN U20284 ( .A(n20227), .B(n20228), .Z(n19844) );
  NAND U20285 ( .A(n19845), .B(n19844), .Z(n19846) );
  OR U20286 ( .A(n19847), .B(n19846), .Z(n19851) );
  XNOR U20287 ( .A(n19847), .B(n19846), .Z(n20231) );
  XOR U20288 ( .A(n19849), .B(n19848), .Z(n20232) );
  NANDN U20289 ( .A(n20231), .B(n20232), .Z(n19850) );
  NAND U20290 ( .A(n19851), .B(n19850), .Z(n19854) );
  XOR U20291 ( .A(n19853), .B(n19852), .Z(n19855) );
  NANDN U20292 ( .A(n19854), .B(n19855), .Z(n19857) );
  NAND U20293 ( .A(a[36]), .B(b[5]), .Z(n20239) );
  XNOR U20294 ( .A(n19855), .B(n19854), .Z(n20240) );
  NANDN U20295 ( .A(n20239), .B(n20240), .Z(n19856) );
  NAND U20296 ( .A(n19857), .B(n19856), .Z(n19858) );
  OR U20297 ( .A(n19859), .B(n19858), .Z(n19863) );
  XNOR U20298 ( .A(n19859), .B(n19858), .Z(n20243) );
  XOR U20299 ( .A(n19861), .B(n19860), .Z(n20244) );
  NANDN U20300 ( .A(n20243), .B(n20244), .Z(n19862) );
  NAND U20301 ( .A(n19863), .B(n19862), .Z(n19866) );
  XOR U20302 ( .A(n19865), .B(n19864), .Z(n19867) );
  NANDN U20303 ( .A(n19866), .B(n19867), .Z(n19869) );
  NAND U20304 ( .A(a[38]), .B(b[5]), .Z(n20251) );
  XNOR U20305 ( .A(n19867), .B(n19866), .Z(n20252) );
  NANDN U20306 ( .A(n20251), .B(n20252), .Z(n19868) );
  NAND U20307 ( .A(n19869), .B(n19868), .Z(n19870) );
  OR U20308 ( .A(n19871), .B(n19870), .Z(n19875) );
  XNOR U20309 ( .A(n19871), .B(n19870), .Z(n20255) );
  XOR U20310 ( .A(n19873), .B(n19872), .Z(n20256) );
  NANDN U20311 ( .A(n20255), .B(n20256), .Z(n19874) );
  NAND U20312 ( .A(n19875), .B(n19874), .Z(n19878) );
  XOR U20313 ( .A(n19877), .B(n19876), .Z(n19879) );
  NANDN U20314 ( .A(n19878), .B(n19879), .Z(n19881) );
  NAND U20315 ( .A(a[40]), .B(b[5]), .Z(n20263) );
  XNOR U20316 ( .A(n19879), .B(n19878), .Z(n20264) );
  NANDN U20317 ( .A(n20263), .B(n20264), .Z(n19880) );
  NAND U20318 ( .A(n19881), .B(n19880), .Z(n19882) );
  OR U20319 ( .A(n19883), .B(n19882), .Z(n19887) );
  XNOR U20320 ( .A(n19883), .B(n19882), .Z(n20267) );
  XOR U20321 ( .A(n19885), .B(n19884), .Z(n20268) );
  NANDN U20322 ( .A(n20267), .B(n20268), .Z(n19886) );
  NAND U20323 ( .A(n19887), .B(n19886), .Z(n19890) );
  XOR U20324 ( .A(n19889), .B(n19888), .Z(n19891) );
  NANDN U20325 ( .A(n19890), .B(n19891), .Z(n19893) );
  NAND U20326 ( .A(a[42]), .B(b[5]), .Z(n20275) );
  XNOR U20327 ( .A(n19891), .B(n19890), .Z(n20276) );
  NANDN U20328 ( .A(n20275), .B(n20276), .Z(n19892) );
  NAND U20329 ( .A(n19893), .B(n19892), .Z(n19894) );
  OR U20330 ( .A(n19895), .B(n19894), .Z(n19899) );
  XNOR U20331 ( .A(n19895), .B(n19894), .Z(n20279) );
  XOR U20332 ( .A(n19897), .B(n19896), .Z(n20280) );
  NANDN U20333 ( .A(n20279), .B(n20280), .Z(n19898) );
  NAND U20334 ( .A(n19899), .B(n19898), .Z(n19902) );
  XOR U20335 ( .A(n19901), .B(n19900), .Z(n19903) );
  NANDN U20336 ( .A(n19902), .B(n19903), .Z(n19905) );
  NAND U20337 ( .A(a[44]), .B(b[5]), .Z(n20287) );
  XNOR U20338 ( .A(n19903), .B(n19902), .Z(n20288) );
  NANDN U20339 ( .A(n20287), .B(n20288), .Z(n19904) );
  NAND U20340 ( .A(n19905), .B(n19904), .Z(n19906) );
  OR U20341 ( .A(n19907), .B(n19906), .Z(n19911) );
  XNOR U20342 ( .A(n19907), .B(n19906), .Z(n20291) );
  XOR U20343 ( .A(n19909), .B(n19908), .Z(n20292) );
  NANDN U20344 ( .A(n20291), .B(n20292), .Z(n19910) );
  NAND U20345 ( .A(n19911), .B(n19910), .Z(n19914) );
  XOR U20346 ( .A(n19913), .B(n19912), .Z(n19915) );
  NANDN U20347 ( .A(n19914), .B(n19915), .Z(n19917) );
  NAND U20348 ( .A(a[46]), .B(b[5]), .Z(n20299) );
  XNOR U20349 ( .A(n19915), .B(n19914), .Z(n20300) );
  NANDN U20350 ( .A(n20299), .B(n20300), .Z(n19916) );
  NAND U20351 ( .A(n19917), .B(n19916), .Z(n19918) );
  OR U20352 ( .A(n19919), .B(n19918), .Z(n19923) );
  XNOR U20353 ( .A(n19919), .B(n19918), .Z(n20303) );
  XOR U20354 ( .A(n19921), .B(n19920), .Z(n20304) );
  NANDN U20355 ( .A(n20303), .B(n20304), .Z(n19922) );
  NAND U20356 ( .A(n19923), .B(n19922), .Z(n19926) );
  XOR U20357 ( .A(n19925), .B(n19924), .Z(n19927) );
  NANDN U20358 ( .A(n19926), .B(n19927), .Z(n19929) );
  NAND U20359 ( .A(a[48]), .B(b[5]), .Z(n20311) );
  XNOR U20360 ( .A(n19927), .B(n19926), .Z(n20312) );
  NANDN U20361 ( .A(n20311), .B(n20312), .Z(n19928) );
  NAND U20362 ( .A(n19929), .B(n19928), .Z(n19930) );
  OR U20363 ( .A(n19931), .B(n19930), .Z(n19935) );
  XNOR U20364 ( .A(n19931), .B(n19930), .Z(n20315) );
  XOR U20365 ( .A(n19933), .B(n19932), .Z(n20316) );
  NANDN U20366 ( .A(n20315), .B(n20316), .Z(n19934) );
  NAND U20367 ( .A(n19935), .B(n19934), .Z(n19938) );
  XOR U20368 ( .A(n19937), .B(n19936), .Z(n19939) );
  NANDN U20369 ( .A(n19938), .B(n19939), .Z(n19941) );
  NAND U20370 ( .A(a[50]), .B(b[5]), .Z(n20323) );
  XNOR U20371 ( .A(n19939), .B(n19938), .Z(n20324) );
  NANDN U20372 ( .A(n20323), .B(n20324), .Z(n19940) );
  NAND U20373 ( .A(n19941), .B(n19940), .Z(n19942) );
  OR U20374 ( .A(n19943), .B(n19942), .Z(n19947) );
  XNOR U20375 ( .A(n19943), .B(n19942), .Z(n20327) );
  XOR U20376 ( .A(n19945), .B(n19944), .Z(n20328) );
  NANDN U20377 ( .A(n20327), .B(n20328), .Z(n19946) );
  NAND U20378 ( .A(n19947), .B(n19946), .Z(n19950) );
  XOR U20379 ( .A(n19949), .B(n19948), .Z(n19951) );
  NANDN U20380 ( .A(n19950), .B(n19951), .Z(n19953) );
  NAND U20381 ( .A(a[52]), .B(b[5]), .Z(n20335) );
  XNOR U20382 ( .A(n19951), .B(n19950), .Z(n20336) );
  NANDN U20383 ( .A(n20335), .B(n20336), .Z(n19952) );
  NAND U20384 ( .A(n19953), .B(n19952), .Z(n19954) );
  OR U20385 ( .A(n19955), .B(n19954), .Z(n19959) );
  XNOR U20386 ( .A(n19955), .B(n19954), .Z(n20339) );
  XOR U20387 ( .A(n19957), .B(n19956), .Z(n20340) );
  NANDN U20388 ( .A(n20339), .B(n20340), .Z(n19958) );
  NAND U20389 ( .A(n19959), .B(n19958), .Z(n19962) );
  XOR U20390 ( .A(n19961), .B(n19960), .Z(n19963) );
  NANDN U20391 ( .A(n19962), .B(n19963), .Z(n19965) );
  NAND U20392 ( .A(a[54]), .B(b[5]), .Z(n20347) );
  XNOR U20393 ( .A(n19963), .B(n19962), .Z(n20348) );
  NANDN U20394 ( .A(n20347), .B(n20348), .Z(n19964) );
  NAND U20395 ( .A(n19965), .B(n19964), .Z(n19966) );
  OR U20396 ( .A(n19967), .B(n19966), .Z(n19971) );
  XNOR U20397 ( .A(n19967), .B(n19966), .Z(n20351) );
  XOR U20398 ( .A(n19969), .B(n19968), .Z(n20352) );
  NANDN U20399 ( .A(n20351), .B(n20352), .Z(n19970) );
  NAND U20400 ( .A(n19971), .B(n19970), .Z(n19974) );
  XOR U20401 ( .A(n19973), .B(n19972), .Z(n19975) );
  NANDN U20402 ( .A(n19974), .B(n19975), .Z(n19977) );
  NAND U20403 ( .A(a[56]), .B(b[5]), .Z(n20359) );
  XNOR U20404 ( .A(n19975), .B(n19974), .Z(n20360) );
  NANDN U20405 ( .A(n20359), .B(n20360), .Z(n19976) );
  NAND U20406 ( .A(n19977), .B(n19976), .Z(n19980) );
  ANDN U20407 ( .B(b[5]), .A(n205), .Z(n19981) );
  OR U20408 ( .A(n19980), .B(n19981), .Z(n19983) );
  XOR U20409 ( .A(n19979), .B(n19978), .Z(n20364) );
  XOR U20410 ( .A(n19981), .B(n19980), .Z(n20363) );
  NANDN U20411 ( .A(n20364), .B(n20363), .Z(n19982) );
  NAND U20412 ( .A(n19983), .B(n19982), .Z(n19986) );
  XNOR U20413 ( .A(n19985), .B(n19984), .Z(n19987) );
  OR U20414 ( .A(n19986), .B(n19987), .Z(n19989) );
  XNOR U20415 ( .A(n19987), .B(n19986), .Z(n20370) );
  NAND U20416 ( .A(a[58]), .B(b[5]), .Z(n20369) );
  OR U20417 ( .A(n20370), .B(n20369), .Z(n19988) );
  NAND U20418 ( .A(n19989), .B(n19988), .Z(n19992) );
  ANDN U20419 ( .B(b[5]), .A(n207), .Z(n19993) );
  OR U20420 ( .A(n19992), .B(n19993), .Z(n19995) );
  XOR U20421 ( .A(n19993), .B(n19992), .Z(n20377) );
  NANDN U20422 ( .A(n20378), .B(n20377), .Z(n19994) );
  NAND U20423 ( .A(n19995), .B(n19994), .Z(n19999) );
  NAND U20424 ( .A(a[60]), .B(b[5]), .Z(n19998) );
  OR U20425 ( .A(n19999), .B(n19998), .Z(n20001) );
  XOR U20426 ( .A(n19997), .B(n19996), .Z(n20381) );
  XOR U20427 ( .A(n19999), .B(n19998), .Z(n20382) );
  NAND U20428 ( .A(n20381), .B(n20382), .Z(n20000) );
  NAND U20429 ( .A(n20001), .B(n20000), .Z(n20005) );
  XOR U20430 ( .A(n20003), .B(n20002), .Z(n20004) );
  NAND U20431 ( .A(n20005), .B(n20004), .Z(n20007) );
  XNOR U20432 ( .A(n20005), .B(n20004), .Z(n20386) );
  NAND U20433 ( .A(a[61]), .B(b[5]), .Z(n20385) );
  OR U20434 ( .A(n20386), .B(n20385), .Z(n20006) );
  NAND U20435 ( .A(n20007), .B(n20006), .Z(n20011) );
  NANDN U20436 ( .A(n20010), .B(n20011), .Z(n20013) );
  XNOR U20437 ( .A(n20009), .B(n20008), .Z(n20388) );
  XNOR U20438 ( .A(n20011), .B(n20010), .Z(n20387) );
  NANDN U20439 ( .A(n20388), .B(n20387), .Z(n20012) );
  NAND U20440 ( .A(n20013), .B(n20012), .Z(n20017) );
  XOR U20441 ( .A(n20015), .B(n20014), .Z(n20016) );
  NAND U20442 ( .A(n20017), .B(n20016), .Z(n20019) );
  XNOR U20443 ( .A(n20017), .B(n20016), .Z(n20023) );
  NAND U20444 ( .A(a[63]), .B(b[5]), .Z(n20022) );
  OR U20445 ( .A(n20023), .B(n20022), .Z(n20018) );
  AND U20446 ( .A(n20019), .B(n20018), .Z(n20020) );
  OR U20447 ( .A(n20021), .B(n20020), .Z(n21927) );
  NANDN U20448 ( .A(n21926), .B(n21927), .Z(n21929) );
  XNOR U20449 ( .A(n20021), .B(n20020), .Z(n24106) );
  XOR U20450 ( .A(n20023), .B(n20022), .Z(n20394) );
  NAND U20451 ( .A(a[62]), .B(b[4]), .Z(n20383) );
  ANDN U20452 ( .B(b[4]), .A(n205), .Z(n20358) );
  ANDN U20453 ( .B(b[4]), .A(n203), .Z(n20346) );
  ANDN U20454 ( .B(b[4]), .A(n201), .Z(n20334) );
  ANDN U20455 ( .B(b[4]), .A(n199), .Z(n20322) );
  ANDN U20456 ( .B(b[4]), .A(n197), .Z(n20310) );
  ANDN U20457 ( .B(b[4]), .A(n195), .Z(n20298) );
  ANDN U20458 ( .B(b[4]), .A(n193), .Z(n20286) );
  ANDN U20459 ( .B(b[4]), .A(n191), .Z(n20274) );
  ANDN U20460 ( .B(b[4]), .A(n189), .Z(n20262) );
  ANDN U20461 ( .B(b[4]), .A(n187), .Z(n20250) );
  ANDN U20462 ( .B(b[4]), .A(n21772), .Z(n20238) );
  ANDN U20463 ( .B(b[4]), .A(n184), .Z(n20226) );
  ANDN U20464 ( .B(b[4]), .A(n21751), .Z(n20214) );
  ANDN U20465 ( .B(b[4]), .A(n21740), .Z(n20202) );
  ANDN U20466 ( .B(b[4]), .A(n21727), .Z(n20190) );
  ANDN U20467 ( .B(b[4]), .A(n21716), .Z(n20178) );
  NAND U20468 ( .A(a[25]), .B(b[4]), .Z(n20166) );
  XNOR U20469 ( .A(n20025), .B(n20024), .Z(n20162) );
  ANDN U20470 ( .B(b[4]), .A(n21692), .Z(n20158) );
  ANDN U20471 ( .B(b[4]), .A(n21681), .Z(n20146) );
  ANDN U20472 ( .B(b[4]), .A(n21670), .Z(n20134) );
  ANDN U20473 ( .B(b[4]), .A(n174), .Z(n20120) );
  ANDN U20474 ( .B(b[4]), .A(n172), .Z(n20110) );
  ANDN U20475 ( .B(b[4]), .A(n170), .Z(n20096) );
  NAND U20476 ( .A(a[12]), .B(b[4]), .Z(n20028) );
  XOR U20477 ( .A(n20027), .B(n20026), .Z(n20029) );
  NANDN U20478 ( .A(n20028), .B(n20029), .Z(n20094) );
  XOR U20479 ( .A(n20029), .B(n20028), .Z(n20477) );
  ANDN U20480 ( .B(b[4]), .A(n21164), .Z(n20088) );
  NAND U20481 ( .A(a[10]), .B(b[4]), .Z(n20083) );
  XOR U20482 ( .A(n20031), .B(n20030), .Z(n20084) );
  NANDN U20483 ( .A(n20083), .B(n20084), .Z(n20086) );
  ANDN U20484 ( .B(b[4]), .A(n21615), .Z(n20078) );
  ANDN U20485 ( .B(b[4]), .A(n166), .Z(n20065) );
  NAND U20486 ( .A(b[5]), .B(a[1]), .Z(n20036) );
  NANDN U20487 ( .A(n20036), .B(a[0]), .Z(n20032) );
  XNOR U20488 ( .A(a[2]), .B(n20032), .Z(n20033) );
  NAND U20489 ( .A(b[4]), .B(n20033), .Z(n20420) );
  AND U20490 ( .A(a[1]), .B(b[5]), .Z(n20034) );
  XOR U20491 ( .A(n20035), .B(n20034), .Z(n20421) );
  OR U20492 ( .A(n20420), .B(n20421), .Z(n20040) );
  AND U20493 ( .A(b[4]), .B(a[0]), .Z(n20785) );
  NANDN U20494 ( .A(n20036), .B(n20785), .Z(n20038) );
  NAND U20495 ( .A(a[2]), .B(b[4]), .Z(n20037) );
  AND U20496 ( .A(n20038), .B(n20037), .Z(n20039) );
  ANDN U20497 ( .B(n20040), .A(n20039), .Z(n20042) );
  NANDN U20498 ( .A(n21580), .B(b[4]), .Z(n20041) );
  NANDN U20499 ( .A(n20042), .B(n20041), .Z(n20046) );
  XOR U20500 ( .A(n20042), .B(n20041), .Z(n20425) );
  XNOR U20501 ( .A(n20044), .B(n20043), .Z(n20424) );
  OR U20502 ( .A(n20425), .B(n20424), .Z(n20045) );
  NAND U20503 ( .A(n20046), .B(n20045), .Z(n20050) );
  XOR U20504 ( .A(n20048), .B(n20047), .Z(n20049) );
  OR U20505 ( .A(n20050), .B(n20049), .Z(n20052) );
  NAND U20506 ( .A(a[4]), .B(b[4]), .Z(n20431) );
  XOR U20507 ( .A(n20050), .B(n20049), .Z(n20430) );
  NANDN U20508 ( .A(n20431), .B(n20430), .Z(n20051) );
  NAND U20509 ( .A(n20052), .B(n20051), .Z(n20053) );
  ANDN U20510 ( .B(b[4]), .A(n164), .Z(n20054) );
  OR U20511 ( .A(n20053), .B(n20054), .Z(n20058) );
  XNOR U20512 ( .A(n20054), .B(n20053), .Z(n20434) );
  OR U20513 ( .A(n20434), .B(n20435), .Z(n20057) );
  AND U20514 ( .A(n20058), .B(n20057), .Z(n20062) );
  XOR U20515 ( .A(n20060), .B(n20059), .Z(n20061) );
  NANDN U20516 ( .A(n20062), .B(n20061), .Z(n20064) );
  XOR U20517 ( .A(n20062), .B(n20061), .Z(n20443) );
  ANDN U20518 ( .B(b[4]), .A(n165), .Z(n20442) );
  OR U20519 ( .A(n20443), .B(n20442), .Z(n20063) );
  AND U20520 ( .A(n20064), .B(n20063), .Z(n20066) );
  OR U20521 ( .A(n20065), .B(n20066), .Z(n20070) );
  XNOR U20522 ( .A(n20066), .B(n20065), .Z(n20447) );
  XNOR U20523 ( .A(n20068), .B(n20067), .Z(n20446) );
  OR U20524 ( .A(n20447), .B(n20446), .Z(n20069) );
  NAND U20525 ( .A(n20070), .B(n20069), .Z(n20073) );
  NANDN U20526 ( .A(n20073), .B(n20074), .Z(n20076) );
  NAND U20527 ( .A(a[8]), .B(b[4]), .Z(n20454) );
  XNOR U20528 ( .A(n20074), .B(n20073), .Z(n20455) );
  NANDN U20529 ( .A(n20454), .B(n20455), .Z(n20075) );
  NAND U20530 ( .A(n20076), .B(n20075), .Z(n20077) );
  OR U20531 ( .A(n20078), .B(n20077), .Z(n20082) );
  XNOR U20532 ( .A(n20078), .B(n20077), .Z(n20407) );
  XOR U20533 ( .A(n20080), .B(n20079), .Z(n20408) );
  NANDN U20534 ( .A(n20407), .B(n20408), .Z(n20081) );
  NAND U20535 ( .A(n20082), .B(n20081), .Z(n20464) );
  XNOR U20536 ( .A(n20084), .B(n20083), .Z(n20465) );
  NANDN U20537 ( .A(n20464), .B(n20465), .Z(n20085) );
  NAND U20538 ( .A(n20086), .B(n20085), .Z(n20087) );
  OR U20539 ( .A(n20088), .B(n20087), .Z(n20092) );
  XNOR U20540 ( .A(n20088), .B(n20087), .Z(n20468) );
  XOR U20541 ( .A(n20090), .B(n20089), .Z(n20469) );
  NANDN U20542 ( .A(n20468), .B(n20469), .Z(n20091) );
  NAND U20543 ( .A(n20092), .B(n20091), .Z(n20476) );
  OR U20544 ( .A(n20477), .B(n20476), .Z(n20093) );
  NAND U20545 ( .A(n20094), .B(n20093), .Z(n20095) );
  OR U20546 ( .A(n20096), .B(n20095), .Z(n20100) );
  XNOR U20547 ( .A(n20096), .B(n20095), .Z(n20403) );
  XOR U20548 ( .A(n20098), .B(n20097), .Z(n20404) );
  NANDN U20549 ( .A(n20403), .B(n20404), .Z(n20099) );
  NAND U20550 ( .A(n20100), .B(n20099), .Z(n20103) );
  XNOR U20551 ( .A(n20102), .B(n20101), .Z(n20104) );
  OR U20552 ( .A(n20103), .B(n20104), .Z(n20106) );
  NAND U20553 ( .A(a[14]), .B(b[4]), .Z(n20484) );
  XOR U20554 ( .A(n20104), .B(n20103), .Z(n20485) );
  NANDN U20555 ( .A(n20484), .B(n20485), .Z(n20105) );
  NAND U20556 ( .A(n20106), .B(n20105), .Z(n20109) );
  OR U20557 ( .A(n20110), .B(n20109), .Z(n20112) );
  XOR U20558 ( .A(n20108), .B(n20107), .Z(n20402) );
  XOR U20559 ( .A(n20110), .B(n20109), .Z(n20401) );
  NAND U20560 ( .A(n20402), .B(n20401), .Z(n20111) );
  NAND U20561 ( .A(n20112), .B(n20111), .Z(n20115) );
  XOR U20562 ( .A(n20114), .B(n20113), .Z(n20116) );
  NANDN U20563 ( .A(n20115), .B(n20116), .Z(n20118) );
  NAND U20564 ( .A(a[16]), .B(b[4]), .Z(n20494) );
  XNOR U20565 ( .A(n20116), .B(n20115), .Z(n20495) );
  NANDN U20566 ( .A(n20494), .B(n20495), .Z(n20117) );
  NAND U20567 ( .A(n20118), .B(n20117), .Z(n20119) );
  OR U20568 ( .A(n20120), .B(n20119), .Z(n20124) );
  XNOR U20569 ( .A(n20120), .B(n20119), .Z(n20498) );
  XOR U20570 ( .A(n20122), .B(n20121), .Z(n20499) );
  NANDN U20571 ( .A(n20498), .B(n20499), .Z(n20123) );
  NAND U20572 ( .A(n20124), .B(n20123), .Z(n20126) );
  NAND U20573 ( .A(a[18]), .B(b[4]), .Z(n20125) );
  OR U20574 ( .A(n20126), .B(n20125), .Z(n20130) );
  XOR U20575 ( .A(n20126), .B(n20125), .Z(n20504) );
  NAND U20576 ( .A(n20504), .B(n20505), .Z(n20129) );
  NAND U20577 ( .A(n20130), .B(n20129), .Z(n20133) );
  OR U20578 ( .A(n20134), .B(n20133), .Z(n20136) );
  XOR U20579 ( .A(n20134), .B(n20133), .Z(n20510) );
  NANDN U20580 ( .A(n20511), .B(n20510), .Z(n20135) );
  NAND U20581 ( .A(n20136), .B(n20135), .Z(n20139) );
  NANDN U20582 ( .A(n20139), .B(n20140), .Z(n20142) );
  NAND U20583 ( .A(a[20]), .B(b[4]), .Z(n20518) );
  XNOR U20584 ( .A(n20140), .B(n20139), .Z(n20519) );
  NANDN U20585 ( .A(n20518), .B(n20519), .Z(n20141) );
  NAND U20586 ( .A(n20142), .B(n20141), .Z(n20145) );
  OR U20587 ( .A(n20146), .B(n20145), .Z(n20148) );
  XOR U20588 ( .A(n20144), .B(n20143), .Z(n20399) );
  XOR U20589 ( .A(n20146), .B(n20145), .Z(n20400) );
  NAND U20590 ( .A(n20399), .B(n20400), .Z(n20147) );
  NAND U20591 ( .A(n20148), .B(n20147), .Z(n20151) );
  XOR U20592 ( .A(n20150), .B(n20149), .Z(n20152) );
  NANDN U20593 ( .A(n20151), .B(n20152), .Z(n20154) );
  NAND U20594 ( .A(a[22]), .B(b[4]), .Z(n20526) );
  XNOR U20595 ( .A(n20152), .B(n20151), .Z(n20527) );
  NANDN U20596 ( .A(n20526), .B(n20527), .Z(n20153) );
  NAND U20597 ( .A(n20154), .B(n20153), .Z(n20157) );
  OR U20598 ( .A(n20158), .B(n20157), .Z(n20160) );
  XOR U20599 ( .A(n20156), .B(n20155), .Z(n20398) );
  XOR U20600 ( .A(n20158), .B(n20157), .Z(n20397) );
  NAND U20601 ( .A(n20398), .B(n20397), .Z(n20159) );
  NAND U20602 ( .A(n20160), .B(n20159), .Z(n20161) );
  NANDN U20603 ( .A(n20162), .B(n20161), .Z(n20164) );
  ANDN U20604 ( .B(b[4]), .A(n178), .Z(n20539) );
  NANDN U20605 ( .A(n20539), .B(n20538), .Z(n20163) );
  AND U20606 ( .A(n20164), .B(n20163), .Z(n20165) );
  NANDN U20607 ( .A(n20166), .B(n20165), .Z(n20170) );
  XNOR U20608 ( .A(n20168), .B(n20167), .Z(n20396) );
  NAND U20609 ( .A(n20395), .B(n20396), .Z(n20169) );
  AND U20610 ( .A(n20170), .B(n20169), .Z(n20173) );
  XOR U20611 ( .A(n20172), .B(n20171), .Z(n20174) );
  NANDN U20612 ( .A(n20173), .B(n20174), .Z(n20176) );
  NAND U20613 ( .A(a[26]), .B(b[4]), .Z(n20548) );
  XNOR U20614 ( .A(n20174), .B(n20173), .Z(n20549) );
  NANDN U20615 ( .A(n20548), .B(n20549), .Z(n20175) );
  NAND U20616 ( .A(n20176), .B(n20175), .Z(n20177) );
  OR U20617 ( .A(n20178), .B(n20177), .Z(n20182) );
  XNOR U20618 ( .A(n20178), .B(n20177), .Z(n20552) );
  XOR U20619 ( .A(n20180), .B(n20179), .Z(n20553) );
  NANDN U20620 ( .A(n20552), .B(n20553), .Z(n20181) );
  NAND U20621 ( .A(n20182), .B(n20181), .Z(n20185) );
  XOR U20622 ( .A(n20184), .B(n20183), .Z(n20186) );
  NANDN U20623 ( .A(n20185), .B(n20186), .Z(n20188) );
  NAND U20624 ( .A(a[28]), .B(b[4]), .Z(n20560) );
  XNOR U20625 ( .A(n20186), .B(n20185), .Z(n20561) );
  NANDN U20626 ( .A(n20560), .B(n20561), .Z(n20187) );
  NAND U20627 ( .A(n20188), .B(n20187), .Z(n20189) );
  OR U20628 ( .A(n20190), .B(n20189), .Z(n20194) );
  XNOR U20629 ( .A(n20190), .B(n20189), .Z(n20564) );
  XOR U20630 ( .A(n20192), .B(n20191), .Z(n20565) );
  NANDN U20631 ( .A(n20564), .B(n20565), .Z(n20193) );
  NAND U20632 ( .A(n20194), .B(n20193), .Z(n20197) );
  XOR U20633 ( .A(n20196), .B(n20195), .Z(n20198) );
  NANDN U20634 ( .A(n20197), .B(n20198), .Z(n20200) );
  NAND U20635 ( .A(a[30]), .B(b[4]), .Z(n20572) );
  XNOR U20636 ( .A(n20198), .B(n20197), .Z(n20573) );
  NANDN U20637 ( .A(n20572), .B(n20573), .Z(n20199) );
  NAND U20638 ( .A(n20200), .B(n20199), .Z(n20201) );
  OR U20639 ( .A(n20202), .B(n20201), .Z(n20206) );
  XNOR U20640 ( .A(n20202), .B(n20201), .Z(n20576) );
  XOR U20641 ( .A(n20204), .B(n20203), .Z(n20577) );
  NANDN U20642 ( .A(n20576), .B(n20577), .Z(n20205) );
  NAND U20643 ( .A(n20206), .B(n20205), .Z(n20209) );
  XOR U20644 ( .A(n20208), .B(n20207), .Z(n20210) );
  NANDN U20645 ( .A(n20209), .B(n20210), .Z(n20212) );
  NAND U20646 ( .A(a[32]), .B(b[4]), .Z(n20584) );
  XNOR U20647 ( .A(n20210), .B(n20209), .Z(n20585) );
  NANDN U20648 ( .A(n20584), .B(n20585), .Z(n20211) );
  NAND U20649 ( .A(n20212), .B(n20211), .Z(n20213) );
  OR U20650 ( .A(n20214), .B(n20213), .Z(n20218) );
  XNOR U20651 ( .A(n20214), .B(n20213), .Z(n20588) );
  XOR U20652 ( .A(n20216), .B(n20215), .Z(n20589) );
  NANDN U20653 ( .A(n20588), .B(n20589), .Z(n20217) );
  NAND U20654 ( .A(n20218), .B(n20217), .Z(n20221) );
  XOR U20655 ( .A(n20220), .B(n20219), .Z(n20222) );
  NANDN U20656 ( .A(n20221), .B(n20222), .Z(n20224) );
  NAND U20657 ( .A(a[34]), .B(b[4]), .Z(n20596) );
  XNOR U20658 ( .A(n20222), .B(n20221), .Z(n20597) );
  NANDN U20659 ( .A(n20596), .B(n20597), .Z(n20223) );
  NAND U20660 ( .A(n20224), .B(n20223), .Z(n20225) );
  OR U20661 ( .A(n20226), .B(n20225), .Z(n20230) );
  XNOR U20662 ( .A(n20226), .B(n20225), .Z(n20600) );
  XOR U20663 ( .A(n20228), .B(n20227), .Z(n20601) );
  NANDN U20664 ( .A(n20600), .B(n20601), .Z(n20229) );
  NAND U20665 ( .A(n20230), .B(n20229), .Z(n20233) );
  XOR U20666 ( .A(n20232), .B(n20231), .Z(n20234) );
  NANDN U20667 ( .A(n20233), .B(n20234), .Z(n20236) );
  NAND U20668 ( .A(a[36]), .B(b[4]), .Z(n20608) );
  XNOR U20669 ( .A(n20234), .B(n20233), .Z(n20609) );
  NANDN U20670 ( .A(n20608), .B(n20609), .Z(n20235) );
  NAND U20671 ( .A(n20236), .B(n20235), .Z(n20237) );
  OR U20672 ( .A(n20238), .B(n20237), .Z(n20242) );
  XNOR U20673 ( .A(n20238), .B(n20237), .Z(n20612) );
  XOR U20674 ( .A(n20240), .B(n20239), .Z(n20613) );
  NANDN U20675 ( .A(n20612), .B(n20613), .Z(n20241) );
  NAND U20676 ( .A(n20242), .B(n20241), .Z(n20245) );
  XOR U20677 ( .A(n20244), .B(n20243), .Z(n20246) );
  NANDN U20678 ( .A(n20245), .B(n20246), .Z(n20248) );
  NAND U20679 ( .A(a[38]), .B(b[4]), .Z(n20620) );
  XNOR U20680 ( .A(n20246), .B(n20245), .Z(n20621) );
  NANDN U20681 ( .A(n20620), .B(n20621), .Z(n20247) );
  NAND U20682 ( .A(n20248), .B(n20247), .Z(n20249) );
  OR U20683 ( .A(n20250), .B(n20249), .Z(n20254) );
  XNOR U20684 ( .A(n20250), .B(n20249), .Z(n20624) );
  XOR U20685 ( .A(n20252), .B(n20251), .Z(n20625) );
  NANDN U20686 ( .A(n20624), .B(n20625), .Z(n20253) );
  NAND U20687 ( .A(n20254), .B(n20253), .Z(n20257) );
  XOR U20688 ( .A(n20256), .B(n20255), .Z(n20258) );
  NANDN U20689 ( .A(n20257), .B(n20258), .Z(n20260) );
  NAND U20690 ( .A(a[40]), .B(b[4]), .Z(n20632) );
  XNOR U20691 ( .A(n20258), .B(n20257), .Z(n20633) );
  NANDN U20692 ( .A(n20632), .B(n20633), .Z(n20259) );
  NAND U20693 ( .A(n20260), .B(n20259), .Z(n20261) );
  OR U20694 ( .A(n20262), .B(n20261), .Z(n20266) );
  XNOR U20695 ( .A(n20262), .B(n20261), .Z(n20636) );
  XOR U20696 ( .A(n20264), .B(n20263), .Z(n20637) );
  NANDN U20697 ( .A(n20636), .B(n20637), .Z(n20265) );
  NAND U20698 ( .A(n20266), .B(n20265), .Z(n20269) );
  XOR U20699 ( .A(n20268), .B(n20267), .Z(n20270) );
  NANDN U20700 ( .A(n20269), .B(n20270), .Z(n20272) );
  NAND U20701 ( .A(a[42]), .B(b[4]), .Z(n20644) );
  XNOR U20702 ( .A(n20270), .B(n20269), .Z(n20645) );
  NANDN U20703 ( .A(n20644), .B(n20645), .Z(n20271) );
  NAND U20704 ( .A(n20272), .B(n20271), .Z(n20273) );
  OR U20705 ( .A(n20274), .B(n20273), .Z(n20278) );
  XNOR U20706 ( .A(n20274), .B(n20273), .Z(n20648) );
  XOR U20707 ( .A(n20276), .B(n20275), .Z(n20649) );
  NANDN U20708 ( .A(n20648), .B(n20649), .Z(n20277) );
  NAND U20709 ( .A(n20278), .B(n20277), .Z(n20281) );
  XOR U20710 ( .A(n20280), .B(n20279), .Z(n20282) );
  NANDN U20711 ( .A(n20281), .B(n20282), .Z(n20284) );
  NAND U20712 ( .A(a[44]), .B(b[4]), .Z(n20656) );
  XNOR U20713 ( .A(n20282), .B(n20281), .Z(n20657) );
  NANDN U20714 ( .A(n20656), .B(n20657), .Z(n20283) );
  NAND U20715 ( .A(n20284), .B(n20283), .Z(n20285) );
  OR U20716 ( .A(n20286), .B(n20285), .Z(n20290) );
  XNOR U20717 ( .A(n20286), .B(n20285), .Z(n20660) );
  XOR U20718 ( .A(n20288), .B(n20287), .Z(n20661) );
  NANDN U20719 ( .A(n20660), .B(n20661), .Z(n20289) );
  NAND U20720 ( .A(n20290), .B(n20289), .Z(n20293) );
  XOR U20721 ( .A(n20292), .B(n20291), .Z(n20294) );
  NANDN U20722 ( .A(n20293), .B(n20294), .Z(n20296) );
  NAND U20723 ( .A(a[46]), .B(b[4]), .Z(n20668) );
  XNOR U20724 ( .A(n20294), .B(n20293), .Z(n20669) );
  NANDN U20725 ( .A(n20668), .B(n20669), .Z(n20295) );
  NAND U20726 ( .A(n20296), .B(n20295), .Z(n20297) );
  OR U20727 ( .A(n20298), .B(n20297), .Z(n20302) );
  XNOR U20728 ( .A(n20298), .B(n20297), .Z(n20672) );
  XOR U20729 ( .A(n20300), .B(n20299), .Z(n20673) );
  NANDN U20730 ( .A(n20672), .B(n20673), .Z(n20301) );
  NAND U20731 ( .A(n20302), .B(n20301), .Z(n20305) );
  XOR U20732 ( .A(n20304), .B(n20303), .Z(n20306) );
  NANDN U20733 ( .A(n20305), .B(n20306), .Z(n20308) );
  NAND U20734 ( .A(a[48]), .B(b[4]), .Z(n20680) );
  XNOR U20735 ( .A(n20306), .B(n20305), .Z(n20681) );
  NANDN U20736 ( .A(n20680), .B(n20681), .Z(n20307) );
  NAND U20737 ( .A(n20308), .B(n20307), .Z(n20309) );
  OR U20738 ( .A(n20310), .B(n20309), .Z(n20314) );
  XNOR U20739 ( .A(n20310), .B(n20309), .Z(n20684) );
  XOR U20740 ( .A(n20312), .B(n20311), .Z(n20685) );
  NANDN U20741 ( .A(n20684), .B(n20685), .Z(n20313) );
  NAND U20742 ( .A(n20314), .B(n20313), .Z(n20317) );
  XOR U20743 ( .A(n20316), .B(n20315), .Z(n20318) );
  NANDN U20744 ( .A(n20317), .B(n20318), .Z(n20320) );
  NAND U20745 ( .A(a[50]), .B(b[4]), .Z(n20692) );
  XNOR U20746 ( .A(n20318), .B(n20317), .Z(n20693) );
  NANDN U20747 ( .A(n20692), .B(n20693), .Z(n20319) );
  NAND U20748 ( .A(n20320), .B(n20319), .Z(n20321) );
  OR U20749 ( .A(n20322), .B(n20321), .Z(n20326) );
  XNOR U20750 ( .A(n20322), .B(n20321), .Z(n20696) );
  XOR U20751 ( .A(n20324), .B(n20323), .Z(n20697) );
  NANDN U20752 ( .A(n20696), .B(n20697), .Z(n20325) );
  NAND U20753 ( .A(n20326), .B(n20325), .Z(n20329) );
  XOR U20754 ( .A(n20328), .B(n20327), .Z(n20330) );
  NANDN U20755 ( .A(n20329), .B(n20330), .Z(n20332) );
  NAND U20756 ( .A(a[52]), .B(b[4]), .Z(n20704) );
  XNOR U20757 ( .A(n20330), .B(n20329), .Z(n20705) );
  NANDN U20758 ( .A(n20704), .B(n20705), .Z(n20331) );
  NAND U20759 ( .A(n20332), .B(n20331), .Z(n20333) );
  OR U20760 ( .A(n20334), .B(n20333), .Z(n20338) );
  XNOR U20761 ( .A(n20334), .B(n20333), .Z(n20708) );
  XOR U20762 ( .A(n20336), .B(n20335), .Z(n20709) );
  NANDN U20763 ( .A(n20708), .B(n20709), .Z(n20337) );
  NAND U20764 ( .A(n20338), .B(n20337), .Z(n20341) );
  XOR U20765 ( .A(n20340), .B(n20339), .Z(n20342) );
  NANDN U20766 ( .A(n20341), .B(n20342), .Z(n20344) );
  NAND U20767 ( .A(a[54]), .B(b[4]), .Z(n20716) );
  XNOR U20768 ( .A(n20342), .B(n20341), .Z(n20717) );
  NANDN U20769 ( .A(n20716), .B(n20717), .Z(n20343) );
  NAND U20770 ( .A(n20344), .B(n20343), .Z(n20345) );
  OR U20771 ( .A(n20346), .B(n20345), .Z(n20350) );
  XNOR U20772 ( .A(n20346), .B(n20345), .Z(n20720) );
  XOR U20773 ( .A(n20348), .B(n20347), .Z(n20721) );
  NANDN U20774 ( .A(n20720), .B(n20721), .Z(n20349) );
  NAND U20775 ( .A(n20350), .B(n20349), .Z(n20353) );
  XOR U20776 ( .A(n20352), .B(n20351), .Z(n20354) );
  NANDN U20777 ( .A(n20353), .B(n20354), .Z(n20356) );
  NAND U20778 ( .A(a[56]), .B(b[4]), .Z(n20728) );
  XNOR U20779 ( .A(n20354), .B(n20353), .Z(n20729) );
  NANDN U20780 ( .A(n20728), .B(n20729), .Z(n20355) );
  NAND U20781 ( .A(n20356), .B(n20355), .Z(n20357) );
  OR U20782 ( .A(n20358), .B(n20357), .Z(n20362) );
  XNOR U20783 ( .A(n20358), .B(n20357), .Z(n20732) );
  XOR U20784 ( .A(n20360), .B(n20359), .Z(n20733) );
  NANDN U20785 ( .A(n20732), .B(n20733), .Z(n20361) );
  NAND U20786 ( .A(n20362), .B(n20361), .Z(n20365) );
  XNOR U20787 ( .A(n20364), .B(n20363), .Z(n20366) );
  OR U20788 ( .A(n20365), .B(n20366), .Z(n20368) );
  XNOR U20789 ( .A(n20366), .B(n20365), .Z(n20739) );
  NAND U20790 ( .A(a[58]), .B(b[4]), .Z(n20738) );
  OR U20791 ( .A(n20739), .B(n20738), .Z(n20367) );
  NAND U20792 ( .A(n20368), .B(n20367), .Z(n20371) );
  ANDN U20793 ( .B(b[4]), .A(n207), .Z(n20372) );
  OR U20794 ( .A(n20371), .B(n20372), .Z(n20374) );
  XOR U20795 ( .A(n20370), .B(n20369), .Z(n20745) );
  XOR U20796 ( .A(n20372), .B(n20371), .Z(n20744) );
  NANDN U20797 ( .A(n20745), .B(n20744), .Z(n20373) );
  NAND U20798 ( .A(n20374), .B(n20373), .Z(n20376) );
  AND U20799 ( .A(b[4]), .B(a[60]), .Z(n20375) );
  NANDN U20800 ( .A(n20376), .B(n20375), .Z(n20380) );
  XNOR U20801 ( .A(n20376), .B(n20375), .Z(n20750) );
  NAND U20802 ( .A(n20750), .B(n20751), .Z(n20379) );
  AND U20803 ( .A(n20380), .B(n20379), .Z(n20757) );
  XOR U20804 ( .A(n20382), .B(n20381), .Z(n20756) );
  NAND U20805 ( .A(a[61]), .B(b[4]), .Z(n20759) );
  XOR U20806 ( .A(n20384), .B(n20383), .Z(n20761) );
  XOR U20807 ( .A(n20386), .B(n20385), .Z(n20760) );
  AND U20808 ( .A(b[4]), .B(a[63]), .Z(n20390) );
  OR U20809 ( .A(n20389), .B(n20390), .Z(n20392) );
  XOR U20810 ( .A(n20388), .B(n20387), .Z(n20767) );
  XOR U20811 ( .A(n20390), .B(n20389), .Z(n20766) );
  NAND U20812 ( .A(n20767), .B(n20766), .Z(n20391) );
  NAND U20813 ( .A(n20392), .B(n20391), .Z(n20393) );
  NANDN U20814 ( .A(n24106), .B(n24105), .Z(n20768) );
  XOR U20815 ( .A(n20394), .B(n20393), .Z(n24095) );
  ANDN U20816 ( .B(b[3]), .A(n205), .Z(n20727) );
  ANDN U20817 ( .B(b[3]), .A(n203), .Z(n20715) );
  ANDN U20818 ( .B(b[3]), .A(n201), .Z(n20703) );
  ANDN U20819 ( .B(b[3]), .A(n199), .Z(n20691) );
  ANDN U20820 ( .B(b[3]), .A(n197), .Z(n20679) );
  ANDN U20821 ( .B(b[3]), .A(n195), .Z(n20667) );
  ANDN U20822 ( .B(b[3]), .A(n193), .Z(n20655) );
  ANDN U20823 ( .B(b[3]), .A(n191), .Z(n20643) );
  ANDN U20824 ( .B(b[3]), .A(n189), .Z(n20631) );
  ANDN U20825 ( .B(b[3]), .A(n187), .Z(n20619) );
  ANDN U20826 ( .B(b[3]), .A(n21772), .Z(n20607) );
  ANDN U20827 ( .B(b[3]), .A(n184), .Z(n20595) );
  ANDN U20828 ( .B(b[3]), .A(n21751), .Z(n20583) );
  ANDN U20829 ( .B(b[3]), .A(n21740), .Z(n20571) );
  ANDN U20830 ( .B(b[3]), .A(n21727), .Z(n20559) );
  NAND U20831 ( .A(a[27]), .B(b[3]), .Z(n20547) );
  ANDN U20832 ( .B(b[3]), .A(n21703), .Z(n20536) );
  XNOR U20833 ( .A(n20398), .B(n20397), .Z(n20533) );
  ANDN U20834 ( .B(b[3]), .A(n21692), .Z(n20529) );
  ANDN U20835 ( .B(b[3]), .A(n21681), .Z(n20517) );
  ANDN U20836 ( .B(b[3]), .A(n21670), .Z(n20507) );
  ANDN U20837 ( .B(b[3]), .A(n174), .Z(n20493) );
  XNOR U20838 ( .A(n20402), .B(n20401), .Z(n20489) );
  ANDN U20839 ( .B(b[3]), .A(n172), .Z(n20483) );
  NAND U20840 ( .A(a[14]), .B(b[3]), .Z(n20405) );
  XOR U20841 ( .A(n20404), .B(n20403), .Z(n20406) );
  NANDN U20842 ( .A(n20405), .B(n20406), .Z(n20481) );
  XOR U20843 ( .A(n20406), .B(n20405), .Z(n20857) );
  NAND U20844 ( .A(a[13]), .B(b[3]), .Z(n20475) );
  NAND U20845 ( .A(a[12]), .B(b[3]), .Z(n20471) );
  ANDN U20846 ( .B(b[3]), .A(n21164), .Z(n20463) );
  NAND U20847 ( .A(a[10]), .B(b[3]), .Z(n20458) );
  XOR U20848 ( .A(n20408), .B(n20407), .Z(n20459) );
  NANDN U20849 ( .A(n20458), .B(n20459), .Z(n20461) );
  ANDN U20850 ( .B(b[3]), .A(n21615), .Z(n20453) );
  ANDN U20851 ( .B(b[3]), .A(n166), .Z(n20440) );
  NAND U20852 ( .A(b[4]), .B(a[1]), .Z(n20411) );
  AND U20853 ( .A(b[3]), .B(a[0]), .Z(n21171) );
  NANDN U20854 ( .A(n20411), .B(n21171), .Z(n20410) );
  NAND U20855 ( .A(b[3]), .B(a[2]), .Z(n20409) );
  AND U20856 ( .A(n20410), .B(n20409), .Z(n20417) );
  NANDN U20857 ( .A(n20411), .B(a[0]), .Z(n20412) );
  XNOR U20858 ( .A(a[2]), .B(n20412), .Z(n20413) );
  NAND U20859 ( .A(b[3]), .B(n20413), .Z(n20790) );
  AND U20860 ( .A(a[1]), .B(b[4]), .Z(n20414) );
  XNOR U20861 ( .A(n20415), .B(n20414), .Z(n20791) );
  NANDN U20862 ( .A(n20790), .B(n20791), .Z(n20416) );
  NANDN U20863 ( .A(n20417), .B(n20416), .Z(n20419) );
  NANDN U20864 ( .A(n152), .B(a[3]), .Z(n20418) );
  NAND U20865 ( .A(n20419), .B(n20418), .Z(n20423) );
  XNOR U20866 ( .A(n20419), .B(n20418), .Z(n20795) );
  XNOR U20867 ( .A(n20421), .B(n20420), .Z(n20794) );
  OR U20868 ( .A(n20795), .B(n20794), .Z(n20422) );
  NAND U20869 ( .A(n20423), .B(n20422), .Z(n20427) );
  XOR U20870 ( .A(n20425), .B(n20424), .Z(n20426) );
  NAND U20871 ( .A(a[4]), .B(b[3]), .Z(n20802) );
  XOR U20872 ( .A(n20427), .B(n20426), .Z(n20803) );
  ANDN U20873 ( .B(b[3]), .A(n164), .Z(n20429) );
  OR U20874 ( .A(n20428), .B(n20429), .Z(n20433) );
  XNOR U20875 ( .A(n20429), .B(n20428), .Z(n20804) );
  OR U20876 ( .A(n20804), .B(n20805), .Z(n20432) );
  AND U20877 ( .A(n20433), .B(n20432), .Z(n20437) );
  XOR U20878 ( .A(n20435), .B(n20434), .Z(n20436) );
  NANDN U20879 ( .A(n20437), .B(n20436), .Z(n20439) );
  XOR U20880 ( .A(n20437), .B(n20436), .Z(n20813) );
  ANDN U20881 ( .B(b[3]), .A(n165), .Z(n20812) );
  OR U20882 ( .A(n20813), .B(n20812), .Z(n20438) );
  AND U20883 ( .A(n20439), .B(n20438), .Z(n20441) );
  OR U20884 ( .A(n20440), .B(n20441), .Z(n20445) );
  XNOR U20885 ( .A(n20441), .B(n20440), .Z(n20817) );
  XNOR U20886 ( .A(n20443), .B(n20442), .Z(n20816) );
  OR U20887 ( .A(n20817), .B(n20816), .Z(n20444) );
  NAND U20888 ( .A(n20445), .B(n20444), .Z(n20449) );
  XOR U20889 ( .A(n20447), .B(n20446), .Z(n20448) );
  OR U20890 ( .A(n20449), .B(n20448), .Z(n20451) );
  NAND U20891 ( .A(a[8]), .B(b[3]), .Z(n20825) );
  XOR U20892 ( .A(n20449), .B(n20448), .Z(n20824) );
  NANDN U20893 ( .A(n20825), .B(n20824), .Z(n20450) );
  NAND U20894 ( .A(n20451), .B(n20450), .Z(n20452) );
  OR U20895 ( .A(n20453), .B(n20452), .Z(n20457) );
  XNOR U20896 ( .A(n20453), .B(n20452), .Z(n20828) );
  XOR U20897 ( .A(n20455), .B(n20454), .Z(n20829) );
  NANDN U20898 ( .A(n20828), .B(n20829), .Z(n20456) );
  NAND U20899 ( .A(n20457), .B(n20456), .Z(n20836) );
  XNOR U20900 ( .A(n20459), .B(n20458), .Z(n20837) );
  NANDN U20901 ( .A(n20836), .B(n20837), .Z(n20460) );
  NAND U20902 ( .A(n20461), .B(n20460), .Z(n20462) );
  OR U20903 ( .A(n20463), .B(n20462), .Z(n20467) );
  XNOR U20904 ( .A(n20463), .B(n20462), .Z(n20777) );
  XOR U20905 ( .A(n20465), .B(n20464), .Z(n20778) );
  NANDN U20906 ( .A(n20777), .B(n20778), .Z(n20466) );
  AND U20907 ( .A(n20467), .B(n20466), .Z(n20470) );
  NANDN U20908 ( .A(n20471), .B(n20470), .Z(n20473) );
  XOR U20909 ( .A(n20469), .B(n20468), .Z(n20845) );
  NAND U20910 ( .A(n20845), .B(n20844), .Z(n20472) );
  NAND U20911 ( .A(n20473), .B(n20472), .Z(n20474) );
  NANDN U20912 ( .A(n20475), .B(n20474), .Z(n20479) );
  XOR U20913 ( .A(n20477), .B(n20476), .Z(n20853) );
  NAND U20914 ( .A(n20852), .B(n20853), .Z(n20478) );
  NAND U20915 ( .A(n20479), .B(n20478), .Z(n20856) );
  NANDN U20916 ( .A(n20857), .B(n20856), .Z(n20480) );
  NAND U20917 ( .A(n20481), .B(n20480), .Z(n20482) );
  OR U20918 ( .A(n20483), .B(n20482), .Z(n20487) );
  XNOR U20919 ( .A(n20483), .B(n20482), .Z(n20773) );
  XOR U20920 ( .A(n20485), .B(n20484), .Z(n20774) );
  NANDN U20921 ( .A(n20773), .B(n20774), .Z(n20486) );
  NAND U20922 ( .A(n20487), .B(n20486), .Z(n20488) );
  NANDN U20923 ( .A(n20489), .B(n20488), .Z(n20491) );
  ANDN U20924 ( .B(b[3]), .A(n173), .Z(n20865) );
  NANDN U20925 ( .A(n20865), .B(n20864), .Z(n20490) );
  AND U20926 ( .A(n20491), .B(n20490), .Z(n20492) );
  OR U20927 ( .A(n20493), .B(n20492), .Z(n20497) );
  XNOR U20928 ( .A(n20493), .B(n20492), .Z(n20870) );
  XOR U20929 ( .A(n20495), .B(n20494), .Z(n20871) );
  NANDN U20930 ( .A(n20870), .B(n20871), .Z(n20496) );
  NAND U20931 ( .A(n20497), .B(n20496), .Z(n20500) );
  XOR U20932 ( .A(n20499), .B(n20498), .Z(n20501) );
  NANDN U20933 ( .A(n20500), .B(n20501), .Z(n20503) );
  NAND U20934 ( .A(a[18]), .B(b[3]), .Z(n20878) );
  XNOR U20935 ( .A(n20501), .B(n20500), .Z(n20879) );
  NANDN U20936 ( .A(n20878), .B(n20879), .Z(n20502) );
  NAND U20937 ( .A(n20503), .B(n20502), .Z(n20506) );
  OR U20938 ( .A(n20507), .B(n20506), .Z(n20509) );
  XOR U20939 ( .A(n20507), .B(n20506), .Z(n20882) );
  NANDN U20940 ( .A(n20883), .B(n20882), .Z(n20508) );
  NAND U20941 ( .A(n20509), .B(n20508), .Z(n20512) );
  NANDN U20942 ( .A(n20512), .B(n20513), .Z(n20515) );
  NAND U20943 ( .A(a[20]), .B(b[3]), .Z(n20890) );
  XNOR U20944 ( .A(n20513), .B(n20512), .Z(n20891) );
  NANDN U20945 ( .A(n20890), .B(n20891), .Z(n20514) );
  NAND U20946 ( .A(n20515), .B(n20514), .Z(n20516) );
  OR U20947 ( .A(n20517), .B(n20516), .Z(n20521) );
  XNOR U20948 ( .A(n20517), .B(n20516), .Z(n20894) );
  XOR U20949 ( .A(n20519), .B(n20518), .Z(n20895) );
  NANDN U20950 ( .A(n20894), .B(n20895), .Z(n20520) );
  NAND U20951 ( .A(n20521), .B(n20520), .Z(n20522) );
  OR U20952 ( .A(n20523), .B(n20522), .Z(n20525) );
  NAND U20953 ( .A(b[3]), .B(a[22]), .Z(n20902) );
  XOR U20954 ( .A(n20523), .B(n20522), .Z(n20903) );
  NANDN U20955 ( .A(n20902), .B(n20903), .Z(n20524) );
  NAND U20956 ( .A(n20525), .B(n20524), .Z(n20528) );
  OR U20957 ( .A(n20529), .B(n20528), .Z(n20531) );
  XOR U20958 ( .A(n20527), .B(n20526), .Z(n20772) );
  XOR U20959 ( .A(n20529), .B(n20528), .Z(n20771) );
  NAND U20960 ( .A(n20772), .B(n20771), .Z(n20530) );
  NAND U20961 ( .A(n20531), .B(n20530), .Z(n20532) );
  NANDN U20962 ( .A(n20533), .B(n20532), .Z(n20535) );
  ANDN U20963 ( .B(b[3]), .A(n178), .Z(n20911) );
  NANDN U20964 ( .A(n20911), .B(n20910), .Z(n20534) );
  NAND U20965 ( .A(n20535), .B(n20534), .Z(n20537) );
  NANDN U20966 ( .A(n20536), .B(n20537), .Z(n20541) );
  XOR U20967 ( .A(n20537), .B(n20536), .Z(n20917) );
  XOR U20968 ( .A(n20539), .B(n20538), .Z(n20916) );
  OR U20969 ( .A(n20917), .B(n20916), .Z(n20540) );
  AND U20970 ( .A(n20541), .B(n20540), .Z(n20542) );
  OR U20971 ( .A(n20543), .B(n20542), .Z(n20545) );
  ANDN U20972 ( .B(b[3]), .A(n179), .Z(n20923) );
  XOR U20973 ( .A(n20543), .B(n20542), .Z(n20922) );
  NANDN U20974 ( .A(n20923), .B(n20922), .Z(n20544) );
  AND U20975 ( .A(n20545), .B(n20544), .Z(n20546) );
  NANDN U20976 ( .A(n20547), .B(n20546), .Z(n20551) );
  XNOR U20977 ( .A(n20549), .B(n20548), .Z(n20770) );
  NAND U20978 ( .A(n20769), .B(n20770), .Z(n20550) );
  AND U20979 ( .A(n20551), .B(n20550), .Z(n20554) );
  XOR U20980 ( .A(n20553), .B(n20552), .Z(n20555) );
  NANDN U20981 ( .A(n20554), .B(n20555), .Z(n20557) );
  NAND U20982 ( .A(b[3]), .B(a[28]), .Z(n20934) );
  XNOR U20983 ( .A(n20555), .B(n20554), .Z(n20935) );
  NANDN U20984 ( .A(n20934), .B(n20935), .Z(n20556) );
  NAND U20985 ( .A(n20557), .B(n20556), .Z(n20558) );
  OR U20986 ( .A(n20559), .B(n20558), .Z(n20563) );
  XNOR U20987 ( .A(n20559), .B(n20558), .Z(n20938) );
  XOR U20988 ( .A(n20561), .B(n20560), .Z(n20939) );
  NANDN U20989 ( .A(n20938), .B(n20939), .Z(n20562) );
  NAND U20990 ( .A(n20563), .B(n20562), .Z(n20566) );
  XOR U20991 ( .A(n20565), .B(n20564), .Z(n20567) );
  NANDN U20992 ( .A(n20566), .B(n20567), .Z(n20569) );
  NAND U20993 ( .A(a[30]), .B(b[3]), .Z(n20946) );
  XNOR U20994 ( .A(n20567), .B(n20566), .Z(n20947) );
  NANDN U20995 ( .A(n20946), .B(n20947), .Z(n20568) );
  NAND U20996 ( .A(n20569), .B(n20568), .Z(n20570) );
  OR U20997 ( .A(n20571), .B(n20570), .Z(n20575) );
  XNOR U20998 ( .A(n20571), .B(n20570), .Z(n20950) );
  XOR U20999 ( .A(n20573), .B(n20572), .Z(n20951) );
  NANDN U21000 ( .A(n20950), .B(n20951), .Z(n20574) );
  NAND U21001 ( .A(n20575), .B(n20574), .Z(n20578) );
  XOR U21002 ( .A(n20577), .B(n20576), .Z(n20579) );
  NANDN U21003 ( .A(n20578), .B(n20579), .Z(n20581) );
  NAND U21004 ( .A(a[32]), .B(b[3]), .Z(n20958) );
  XNOR U21005 ( .A(n20579), .B(n20578), .Z(n20959) );
  NANDN U21006 ( .A(n20958), .B(n20959), .Z(n20580) );
  NAND U21007 ( .A(n20581), .B(n20580), .Z(n20582) );
  OR U21008 ( .A(n20583), .B(n20582), .Z(n20587) );
  XNOR U21009 ( .A(n20583), .B(n20582), .Z(n20962) );
  XOR U21010 ( .A(n20585), .B(n20584), .Z(n20963) );
  NANDN U21011 ( .A(n20962), .B(n20963), .Z(n20586) );
  NAND U21012 ( .A(n20587), .B(n20586), .Z(n20590) );
  XOR U21013 ( .A(n20589), .B(n20588), .Z(n20591) );
  NANDN U21014 ( .A(n20590), .B(n20591), .Z(n20593) );
  NAND U21015 ( .A(a[34]), .B(b[3]), .Z(n20970) );
  XNOR U21016 ( .A(n20591), .B(n20590), .Z(n20971) );
  NANDN U21017 ( .A(n20970), .B(n20971), .Z(n20592) );
  NAND U21018 ( .A(n20593), .B(n20592), .Z(n20594) );
  OR U21019 ( .A(n20595), .B(n20594), .Z(n20599) );
  XNOR U21020 ( .A(n20595), .B(n20594), .Z(n20974) );
  XOR U21021 ( .A(n20597), .B(n20596), .Z(n20975) );
  NANDN U21022 ( .A(n20974), .B(n20975), .Z(n20598) );
  NAND U21023 ( .A(n20599), .B(n20598), .Z(n20602) );
  XOR U21024 ( .A(n20601), .B(n20600), .Z(n20603) );
  NANDN U21025 ( .A(n20602), .B(n20603), .Z(n20605) );
  NAND U21026 ( .A(a[36]), .B(b[3]), .Z(n20982) );
  XNOR U21027 ( .A(n20603), .B(n20602), .Z(n20983) );
  NANDN U21028 ( .A(n20982), .B(n20983), .Z(n20604) );
  NAND U21029 ( .A(n20605), .B(n20604), .Z(n20606) );
  OR U21030 ( .A(n20607), .B(n20606), .Z(n20611) );
  XNOR U21031 ( .A(n20607), .B(n20606), .Z(n20986) );
  XOR U21032 ( .A(n20609), .B(n20608), .Z(n20987) );
  NANDN U21033 ( .A(n20986), .B(n20987), .Z(n20610) );
  NAND U21034 ( .A(n20611), .B(n20610), .Z(n20614) );
  XOR U21035 ( .A(n20613), .B(n20612), .Z(n20615) );
  NANDN U21036 ( .A(n20614), .B(n20615), .Z(n20617) );
  NAND U21037 ( .A(a[38]), .B(b[3]), .Z(n20994) );
  XNOR U21038 ( .A(n20615), .B(n20614), .Z(n20995) );
  NANDN U21039 ( .A(n20994), .B(n20995), .Z(n20616) );
  NAND U21040 ( .A(n20617), .B(n20616), .Z(n20618) );
  OR U21041 ( .A(n20619), .B(n20618), .Z(n20623) );
  XNOR U21042 ( .A(n20619), .B(n20618), .Z(n20998) );
  XOR U21043 ( .A(n20621), .B(n20620), .Z(n20999) );
  NANDN U21044 ( .A(n20998), .B(n20999), .Z(n20622) );
  NAND U21045 ( .A(n20623), .B(n20622), .Z(n20626) );
  XOR U21046 ( .A(n20625), .B(n20624), .Z(n20627) );
  NANDN U21047 ( .A(n20626), .B(n20627), .Z(n20629) );
  NAND U21048 ( .A(a[40]), .B(b[3]), .Z(n21006) );
  XNOR U21049 ( .A(n20627), .B(n20626), .Z(n21007) );
  NANDN U21050 ( .A(n21006), .B(n21007), .Z(n20628) );
  NAND U21051 ( .A(n20629), .B(n20628), .Z(n20630) );
  OR U21052 ( .A(n20631), .B(n20630), .Z(n20635) );
  XNOR U21053 ( .A(n20631), .B(n20630), .Z(n21010) );
  XOR U21054 ( .A(n20633), .B(n20632), .Z(n21011) );
  NANDN U21055 ( .A(n21010), .B(n21011), .Z(n20634) );
  NAND U21056 ( .A(n20635), .B(n20634), .Z(n20638) );
  XOR U21057 ( .A(n20637), .B(n20636), .Z(n20639) );
  NANDN U21058 ( .A(n20638), .B(n20639), .Z(n20641) );
  NAND U21059 ( .A(a[42]), .B(b[3]), .Z(n21018) );
  XNOR U21060 ( .A(n20639), .B(n20638), .Z(n21019) );
  NANDN U21061 ( .A(n21018), .B(n21019), .Z(n20640) );
  NAND U21062 ( .A(n20641), .B(n20640), .Z(n20642) );
  OR U21063 ( .A(n20643), .B(n20642), .Z(n20647) );
  XNOR U21064 ( .A(n20643), .B(n20642), .Z(n21022) );
  XOR U21065 ( .A(n20645), .B(n20644), .Z(n21023) );
  NANDN U21066 ( .A(n21022), .B(n21023), .Z(n20646) );
  NAND U21067 ( .A(n20647), .B(n20646), .Z(n20650) );
  XOR U21068 ( .A(n20649), .B(n20648), .Z(n20651) );
  NANDN U21069 ( .A(n20650), .B(n20651), .Z(n20653) );
  NAND U21070 ( .A(a[44]), .B(b[3]), .Z(n21030) );
  XNOR U21071 ( .A(n20651), .B(n20650), .Z(n21031) );
  NANDN U21072 ( .A(n21030), .B(n21031), .Z(n20652) );
  NAND U21073 ( .A(n20653), .B(n20652), .Z(n20654) );
  OR U21074 ( .A(n20655), .B(n20654), .Z(n20659) );
  XNOR U21075 ( .A(n20655), .B(n20654), .Z(n21034) );
  XOR U21076 ( .A(n20657), .B(n20656), .Z(n21035) );
  NANDN U21077 ( .A(n21034), .B(n21035), .Z(n20658) );
  NAND U21078 ( .A(n20659), .B(n20658), .Z(n20662) );
  XOR U21079 ( .A(n20661), .B(n20660), .Z(n20663) );
  NANDN U21080 ( .A(n20662), .B(n20663), .Z(n20665) );
  NAND U21081 ( .A(a[46]), .B(b[3]), .Z(n21042) );
  XNOR U21082 ( .A(n20663), .B(n20662), .Z(n21043) );
  NANDN U21083 ( .A(n21042), .B(n21043), .Z(n20664) );
  NAND U21084 ( .A(n20665), .B(n20664), .Z(n20666) );
  OR U21085 ( .A(n20667), .B(n20666), .Z(n20671) );
  XNOR U21086 ( .A(n20667), .B(n20666), .Z(n21046) );
  XOR U21087 ( .A(n20669), .B(n20668), .Z(n21047) );
  NANDN U21088 ( .A(n21046), .B(n21047), .Z(n20670) );
  NAND U21089 ( .A(n20671), .B(n20670), .Z(n20674) );
  XOR U21090 ( .A(n20673), .B(n20672), .Z(n20675) );
  NANDN U21091 ( .A(n20674), .B(n20675), .Z(n20677) );
  NAND U21092 ( .A(a[48]), .B(b[3]), .Z(n21054) );
  XNOR U21093 ( .A(n20675), .B(n20674), .Z(n21055) );
  NANDN U21094 ( .A(n21054), .B(n21055), .Z(n20676) );
  NAND U21095 ( .A(n20677), .B(n20676), .Z(n20678) );
  OR U21096 ( .A(n20679), .B(n20678), .Z(n20683) );
  XNOR U21097 ( .A(n20679), .B(n20678), .Z(n21058) );
  XOR U21098 ( .A(n20681), .B(n20680), .Z(n21059) );
  NANDN U21099 ( .A(n21058), .B(n21059), .Z(n20682) );
  NAND U21100 ( .A(n20683), .B(n20682), .Z(n20686) );
  XOR U21101 ( .A(n20685), .B(n20684), .Z(n20687) );
  NANDN U21102 ( .A(n20686), .B(n20687), .Z(n20689) );
  NAND U21103 ( .A(a[50]), .B(b[3]), .Z(n21066) );
  XNOR U21104 ( .A(n20687), .B(n20686), .Z(n21067) );
  NANDN U21105 ( .A(n21066), .B(n21067), .Z(n20688) );
  NAND U21106 ( .A(n20689), .B(n20688), .Z(n20690) );
  OR U21107 ( .A(n20691), .B(n20690), .Z(n20695) );
  XNOR U21108 ( .A(n20691), .B(n20690), .Z(n21070) );
  XOR U21109 ( .A(n20693), .B(n20692), .Z(n21071) );
  NANDN U21110 ( .A(n21070), .B(n21071), .Z(n20694) );
  NAND U21111 ( .A(n20695), .B(n20694), .Z(n20698) );
  XOR U21112 ( .A(n20697), .B(n20696), .Z(n20699) );
  NANDN U21113 ( .A(n20698), .B(n20699), .Z(n20701) );
  NAND U21114 ( .A(a[52]), .B(b[3]), .Z(n21078) );
  XNOR U21115 ( .A(n20699), .B(n20698), .Z(n21079) );
  NANDN U21116 ( .A(n21078), .B(n21079), .Z(n20700) );
  NAND U21117 ( .A(n20701), .B(n20700), .Z(n20702) );
  OR U21118 ( .A(n20703), .B(n20702), .Z(n20707) );
  XNOR U21119 ( .A(n20703), .B(n20702), .Z(n21082) );
  XOR U21120 ( .A(n20705), .B(n20704), .Z(n21083) );
  NANDN U21121 ( .A(n21082), .B(n21083), .Z(n20706) );
  NAND U21122 ( .A(n20707), .B(n20706), .Z(n20710) );
  XOR U21123 ( .A(n20709), .B(n20708), .Z(n20711) );
  NANDN U21124 ( .A(n20710), .B(n20711), .Z(n20713) );
  NAND U21125 ( .A(a[54]), .B(b[3]), .Z(n21090) );
  XNOR U21126 ( .A(n20711), .B(n20710), .Z(n21091) );
  NANDN U21127 ( .A(n21090), .B(n21091), .Z(n20712) );
  NAND U21128 ( .A(n20713), .B(n20712), .Z(n20714) );
  OR U21129 ( .A(n20715), .B(n20714), .Z(n20719) );
  XNOR U21130 ( .A(n20715), .B(n20714), .Z(n21094) );
  XOR U21131 ( .A(n20717), .B(n20716), .Z(n21095) );
  NANDN U21132 ( .A(n21094), .B(n21095), .Z(n20718) );
  NAND U21133 ( .A(n20719), .B(n20718), .Z(n20722) );
  XOR U21134 ( .A(n20721), .B(n20720), .Z(n20723) );
  NANDN U21135 ( .A(n20722), .B(n20723), .Z(n20725) );
  NAND U21136 ( .A(a[56]), .B(b[3]), .Z(n21102) );
  XNOR U21137 ( .A(n20723), .B(n20722), .Z(n21103) );
  NANDN U21138 ( .A(n21102), .B(n21103), .Z(n20724) );
  NAND U21139 ( .A(n20725), .B(n20724), .Z(n20726) );
  OR U21140 ( .A(n20727), .B(n20726), .Z(n20731) );
  XNOR U21141 ( .A(n20727), .B(n20726), .Z(n21106) );
  XOR U21142 ( .A(n20729), .B(n20728), .Z(n21107) );
  NANDN U21143 ( .A(n21106), .B(n21107), .Z(n20730) );
  NAND U21144 ( .A(n20731), .B(n20730), .Z(n20734) );
  XOR U21145 ( .A(n20733), .B(n20732), .Z(n20735) );
  NANDN U21146 ( .A(n20734), .B(n20735), .Z(n20737) );
  NAND U21147 ( .A(a[58]), .B(b[3]), .Z(n21114) );
  XNOR U21148 ( .A(n20735), .B(n20734), .Z(n21115) );
  NANDN U21149 ( .A(n21114), .B(n21115), .Z(n20736) );
  NAND U21150 ( .A(n20737), .B(n20736), .Z(n20740) );
  ANDN U21151 ( .B(b[3]), .A(n207), .Z(n20741) );
  OR U21152 ( .A(n20740), .B(n20741), .Z(n20743) );
  XOR U21153 ( .A(n20739), .B(n20738), .Z(n21119) );
  XOR U21154 ( .A(n20741), .B(n20740), .Z(n21118) );
  NANDN U21155 ( .A(n21119), .B(n21118), .Z(n20742) );
  NAND U21156 ( .A(n20743), .B(n20742), .Z(n20746) );
  XNOR U21157 ( .A(n20745), .B(n20744), .Z(n20747) );
  OR U21158 ( .A(n20746), .B(n20747), .Z(n20749) );
  XNOR U21159 ( .A(n20747), .B(n20746), .Z(n21125) );
  NAND U21160 ( .A(a[60]), .B(b[3]), .Z(n21124) );
  OR U21161 ( .A(n21125), .B(n21124), .Z(n20748) );
  NAND U21162 ( .A(n20749), .B(n20748), .Z(n20752) );
  ANDN U21163 ( .B(b[3]), .A(n209), .Z(n20753) );
  OR U21164 ( .A(n20752), .B(n20753), .Z(n20755) );
  XOR U21165 ( .A(n20753), .B(n20752), .Z(n21132) );
  NANDN U21166 ( .A(n21133), .B(n21132), .Z(n20754) );
  AND U21167 ( .A(n20755), .B(n20754), .Z(n21136) );
  ANDN U21168 ( .B(a[62]), .A(n152), .Z(n21137) );
  XNOR U21169 ( .A(n20757), .B(n20756), .Z(n20758) );
  XNOR U21170 ( .A(n20759), .B(n20758), .Z(n21139) );
  XNOR U21171 ( .A(n20761), .B(n20760), .Z(n20762) );
  NANDN U21172 ( .A(n20763), .B(n20762), .Z(n20765) );
  XOR U21173 ( .A(n20763), .B(n20762), .Z(n21141) );
  NAND U21174 ( .A(b[3]), .B(a[63]), .Z(n21140) );
  OR U21175 ( .A(n21141), .B(n21140), .Z(n20764) );
  AND U21176 ( .A(n20765), .B(n20764), .Z(n21142) );
  XNOR U21177 ( .A(n20767), .B(n20766), .Z(n21143) );
  NANDN U21178 ( .A(n21142), .B(n21143), .Z(n24096) );
  NOR U21179 ( .A(n24095), .B(n24096), .Z(n24103) );
  ANDN U21180 ( .B(n20768), .A(n24103), .Z(n21923) );
  AND U21181 ( .A(n24095), .B(n24096), .Z(n21921) );
  ANDN U21182 ( .B(b[2]), .A(n207), .Z(n21113) );
  ANDN U21183 ( .B(b[2]), .A(n205), .Z(n21101) );
  ANDN U21184 ( .B(b[2]), .A(n203), .Z(n21089) );
  ANDN U21185 ( .B(b[2]), .A(n201), .Z(n21077) );
  ANDN U21186 ( .B(b[2]), .A(n199), .Z(n21065) );
  ANDN U21187 ( .B(b[2]), .A(n197), .Z(n21053) );
  ANDN U21188 ( .B(b[2]), .A(n195), .Z(n21041) );
  ANDN U21189 ( .B(b[2]), .A(n193), .Z(n21029) );
  ANDN U21190 ( .B(b[2]), .A(n191), .Z(n21017) );
  ANDN U21191 ( .B(b[2]), .A(n189), .Z(n21005) );
  ANDN U21192 ( .B(b[2]), .A(n187), .Z(n20993) );
  ANDN U21193 ( .B(b[2]), .A(n21772), .Z(n20981) );
  ANDN U21194 ( .B(b[2]), .A(n184), .Z(n20969) );
  ANDN U21195 ( .B(b[2]), .A(n21751), .Z(n20957) );
  ANDN U21196 ( .B(b[2]), .A(n21740), .Z(n20945) );
  NAND U21197 ( .A(a[29]), .B(b[2]), .Z(n20933) );
  ANDN U21198 ( .B(b[2]), .A(n21716), .Z(n20925) );
  ANDN U21199 ( .B(b[2]), .A(n178), .Z(n20907) );
  XNOR U21200 ( .A(n20772), .B(n20771), .Z(n20906) );
  OR U21201 ( .A(n20907), .B(n20906), .Z(n20909) );
  NAND U21202 ( .A(a[23]), .B(b[2]), .Z(n20901) );
  ANDN U21203 ( .B(b[2]), .A(n21681), .Z(n20889) );
  ANDN U21204 ( .B(b[2]), .A(n21670), .Z(n20877) );
  ANDN U21205 ( .B(b[2]), .A(n174), .Z(n20867) );
  NAND U21206 ( .A(a[16]), .B(b[2]), .Z(n20775) );
  XOR U21207 ( .A(n20774), .B(n20773), .Z(n20776) );
  NANDN U21208 ( .A(n20775), .B(n20776), .Z(n20863) );
  XOR U21209 ( .A(n20776), .B(n20775), .Z(n21251) );
  ANDN U21210 ( .B(b[2]), .A(n172), .Z(n20859) );
  ANDN U21211 ( .B(b[2]), .A(n170), .Z(n20847) );
  NAND U21212 ( .A(a[12]), .B(b[2]), .Z(n20840) );
  XOR U21213 ( .A(n20778), .B(n20777), .Z(n20841) );
  NANDN U21214 ( .A(n20840), .B(n20841), .Z(n20843) );
  ANDN U21215 ( .B(b[2]), .A(n21164), .Z(n20835) );
  ANDN U21216 ( .B(b[2]), .A(n166), .Z(n20810) );
  NAND U21217 ( .A(b[3]), .B(a[1]), .Z(n20781) );
  AND U21218 ( .A(b[2]), .B(a[0]), .Z(n21574) );
  NANDN U21219 ( .A(n20781), .B(n21574), .Z(n20780) );
  NAND U21220 ( .A(b[2]), .B(a[2]), .Z(n20779) );
  AND U21221 ( .A(n20780), .B(n20779), .Z(n20787) );
  NANDN U21222 ( .A(n20781), .B(a[0]), .Z(n20782) );
  XNOR U21223 ( .A(a[2]), .B(n20782), .Z(n20783) );
  NAND U21224 ( .A(b[2]), .B(n20783), .Z(n21176) );
  AND U21225 ( .A(a[1]), .B(b[3]), .Z(n20784) );
  XNOR U21226 ( .A(n20785), .B(n20784), .Z(n21177) );
  NANDN U21227 ( .A(n21176), .B(n21177), .Z(n20786) );
  NANDN U21228 ( .A(n20787), .B(n20786), .Z(n20789) );
  NANDN U21229 ( .A(n151), .B(a[3]), .Z(n20788) );
  NAND U21230 ( .A(n20789), .B(n20788), .Z(n20793) );
  XNOR U21231 ( .A(n20789), .B(n20788), .Z(n21181) );
  XNOR U21232 ( .A(n20791), .B(n20790), .Z(n21180) );
  NANDN U21233 ( .A(n21181), .B(n21180), .Z(n20792) );
  NAND U21234 ( .A(n20793), .B(n20792), .Z(n20796) );
  XNOR U21235 ( .A(n20795), .B(n20794), .Z(n20797) );
  NANDN U21236 ( .A(n20796), .B(n20797), .Z(n20799) );
  NAND U21237 ( .A(a[4]), .B(b[2]), .Z(n21186) );
  XNOR U21238 ( .A(n20797), .B(n20796), .Z(n21187) );
  NANDN U21239 ( .A(n21186), .B(n21187), .Z(n20798) );
  NAND U21240 ( .A(n20799), .B(n20798), .Z(n20800) );
  NANDN U21241 ( .A(n151), .B(a[5]), .Z(n20801) );
  XOR U21242 ( .A(n20801), .B(n20800), .Z(n21192) );
  XNOR U21243 ( .A(n20803), .B(n20802), .Z(n21193) );
  XOR U21244 ( .A(n20805), .B(n20804), .Z(n20806) );
  NANDN U21245 ( .A(n20807), .B(n20806), .Z(n20809) );
  XOR U21246 ( .A(n20807), .B(n20806), .Z(n21200) );
  AND U21247 ( .A(a[6]), .B(b[2]), .Z(n21201) );
  OR U21248 ( .A(n21200), .B(n21201), .Z(n20808) );
  AND U21249 ( .A(n20809), .B(n20808), .Z(n20811) );
  OR U21250 ( .A(n20810), .B(n20811), .Z(n20815) );
  XNOR U21251 ( .A(n20811), .B(n20810), .Z(n21205) );
  XNOR U21252 ( .A(n20813), .B(n20812), .Z(n21204) );
  OR U21253 ( .A(n21205), .B(n21204), .Z(n20814) );
  NAND U21254 ( .A(n20815), .B(n20814), .Z(n20819) );
  XOR U21255 ( .A(n20817), .B(n20816), .Z(n20818) );
  OR U21256 ( .A(n20819), .B(n20818), .Z(n20821) );
  NAND U21257 ( .A(a[8]), .B(b[2]), .Z(n21211) );
  XOR U21258 ( .A(n20819), .B(n20818), .Z(n21210) );
  NANDN U21259 ( .A(n21211), .B(n21210), .Z(n20820) );
  NAND U21260 ( .A(n20821), .B(n20820), .Z(n20822) );
  ANDN U21261 ( .B(b[2]), .A(n21615), .Z(n20823) );
  OR U21262 ( .A(n20822), .B(n20823), .Z(n20827) );
  XNOR U21263 ( .A(n20823), .B(n20822), .Z(n21216) );
  OR U21264 ( .A(n21216), .B(n21217), .Z(n20826) );
  NAND U21265 ( .A(n20827), .B(n20826), .Z(n20830) );
  XOR U21266 ( .A(n20829), .B(n20828), .Z(n20831) );
  NANDN U21267 ( .A(n20830), .B(n20831), .Z(n20833) );
  NAND U21268 ( .A(a[10]), .B(b[2]), .Z(n21224) );
  XNOR U21269 ( .A(n20831), .B(n20830), .Z(n21225) );
  NANDN U21270 ( .A(n21224), .B(n21225), .Z(n20832) );
  NAND U21271 ( .A(n20833), .B(n20832), .Z(n20834) );
  OR U21272 ( .A(n20835), .B(n20834), .Z(n20839) );
  XNOR U21273 ( .A(n20835), .B(n20834), .Z(n21160) );
  XOR U21274 ( .A(n20837), .B(n20836), .Z(n21161) );
  NANDN U21275 ( .A(n21160), .B(n21161), .Z(n20838) );
  NAND U21276 ( .A(n20839), .B(n20838), .Z(n21230) );
  XNOR U21277 ( .A(n20841), .B(n20840), .Z(n21231) );
  NANDN U21278 ( .A(n21230), .B(n21231), .Z(n20842) );
  NAND U21279 ( .A(n20843), .B(n20842), .Z(n20846) );
  OR U21280 ( .A(n20847), .B(n20846), .Z(n20849) );
  XOR U21281 ( .A(n20845), .B(n20844), .Z(n21159) );
  XOR U21282 ( .A(n20847), .B(n20846), .Z(n21158) );
  NANDN U21283 ( .A(n21159), .B(n21158), .Z(n20848) );
  NAND U21284 ( .A(n20849), .B(n20848), .Z(n20851) );
  NAND U21285 ( .A(b[2]), .B(a[14]), .Z(n20850) );
  OR U21286 ( .A(n20851), .B(n20850), .Z(n20855) );
  XOR U21287 ( .A(n20851), .B(n20850), .Z(n21240) );
  NAND U21288 ( .A(n21240), .B(n21241), .Z(n20854) );
  NAND U21289 ( .A(n20855), .B(n20854), .Z(n20858) );
  OR U21290 ( .A(n20859), .B(n20858), .Z(n20861) );
  XOR U21291 ( .A(n20859), .B(n20858), .Z(n21156) );
  NAND U21292 ( .A(n21157), .B(n21156), .Z(n20860) );
  AND U21293 ( .A(n20861), .B(n20860), .Z(n21250) );
  NANDN U21294 ( .A(n21251), .B(n21250), .Z(n20862) );
  NAND U21295 ( .A(n20863), .B(n20862), .Z(n20866) );
  OR U21296 ( .A(n20867), .B(n20866), .Z(n20869) );
  XOR U21297 ( .A(n20865), .B(n20864), .Z(n21154) );
  XOR U21298 ( .A(n20867), .B(n20866), .Z(n21155) );
  NANDN U21299 ( .A(n21154), .B(n21155), .Z(n20868) );
  NAND U21300 ( .A(n20869), .B(n20868), .Z(n20872) );
  XOR U21301 ( .A(n20871), .B(n20870), .Z(n20873) );
  NANDN U21302 ( .A(n20872), .B(n20873), .Z(n20875) );
  NAND U21303 ( .A(b[2]), .B(a[18]), .Z(n21260) );
  XNOR U21304 ( .A(n20873), .B(n20872), .Z(n21261) );
  NANDN U21305 ( .A(n21260), .B(n21261), .Z(n20874) );
  NAND U21306 ( .A(n20875), .B(n20874), .Z(n20876) );
  OR U21307 ( .A(n20877), .B(n20876), .Z(n20881) );
  XNOR U21308 ( .A(n20877), .B(n20876), .Z(n21150) );
  XOR U21309 ( .A(n20879), .B(n20878), .Z(n21151) );
  NANDN U21310 ( .A(n21150), .B(n21151), .Z(n20880) );
  NAND U21311 ( .A(n20881), .B(n20880), .Z(n20884) );
  NANDN U21312 ( .A(n20884), .B(n20885), .Z(n20887) );
  NAND U21313 ( .A(a[20]), .B(b[2]), .Z(n21268) );
  XNOR U21314 ( .A(n20885), .B(n20884), .Z(n21269) );
  NANDN U21315 ( .A(n21268), .B(n21269), .Z(n20886) );
  NAND U21316 ( .A(n20887), .B(n20886), .Z(n20888) );
  OR U21317 ( .A(n20889), .B(n20888), .Z(n20893) );
  XNOR U21318 ( .A(n20889), .B(n20888), .Z(n21274) );
  XOR U21319 ( .A(n20891), .B(n20890), .Z(n21275) );
  NANDN U21320 ( .A(n21274), .B(n21275), .Z(n20892) );
  NAND U21321 ( .A(n20893), .B(n20892), .Z(n20896) );
  XOR U21322 ( .A(n20895), .B(n20894), .Z(n20897) );
  NANDN U21323 ( .A(n20896), .B(n20897), .Z(n20899) );
  NAND U21324 ( .A(b[2]), .B(a[22]), .Z(n21280) );
  XNOR U21325 ( .A(n20897), .B(n20896), .Z(n21281) );
  NANDN U21326 ( .A(n21280), .B(n21281), .Z(n20898) );
  NAND U21327 ( .A(n20899), .B(n20898), .Z(n20900) );
  NANDN U21328 ( .A(n20901), .B(n20900), .Z(n20905) );
  XNOR U21329 ( .A(n20903), .B(n20902), .Z(n21287) );
  NAND U21330 ( .A(n21286), .B(n21287), .Z(n20904) );
  AND U21331 ( .A(n20905), .B(n20904), .Z(n21292) );
  XOR U21332 ( .A(n20907), .B(n20906), .Z(n21293) );
  NAND U21333 ( .A(n21292), .B(n21293), .Z(n20908) );
  NAND U21334 ( .A(n20909), .B(n20908), .Z(n20913) );
  NAND U21335 ( .A(b[2]), .B(a[25]), .Z(n20912) );
  OR U21336 ( .A(n20913), .B(n20912), .Z(n20915) );
  XOR U21337 ( .A(n20913), .B(n20912), .Z(n21148) );
  NAND U21338 ( .A(n21149), .B(n21148), .Z(n20914) );
  AND U21339 ( .A(n20915), .B(n20914), .Z(n20919) );
  XNOR U21340 ( .A(n20917), .B(n20916), .Z(n20918) );
  NANDN U21341 ( .A(n20919), .B(n20918), .Z(n20921) );
  NAND U21342 ( .A(b[2]), .B(a[26]), .Z(n21302) );
  NANDN U21343 ( .A(n21302), .B(n21303), .Z(n20920) );
  NAND U21344 ( .A(n20921), .B(n20920), .Z(n20924) );
  OR U21345 ( .A(n20925), .B(n20924), .Z(n20927) );
  XOR U21346 ( .A(n20923), .B(n20922), .Z(n21308) );
  XOR U21347 ( .A(n20925), .B(n20924), .Z(n21309) );
  NANDN U21348 ( .A(n21308), .B(n21309), .Z(n20926) );
  AND U21349 ( .A(n20927), .B(n20926), .Z(n20928) );
  OR U21350 ( .A(n20929), .B(n20928), .Z(n20931) );
  ANDN U21351 ( .B(b[2]), .A(n180), .Z(n21317) );
  XNOR U21352 ( .A(n20929), .B(n20928), .Z(n21316) );
  OR U21353 ( .A(n21317), .B(n21316), .Z(n20930) );
  AND U21354 ( .A(n20931), .B(n20930), .Z(n20932) );
  NANDN U21355 ( .A(n20933), .B(n20932), .Z(n20937) );
  XNOR U21356 ( .A(n20935), .B(n20934), .Z(n21147) );
  NAND U21357 ( .A(n21146), .B(n21147), .Z(n20936) );
  AND U21358 ( .A(n20937), .B(n20936), .Z(n20940) );
  XOR U21359 ( .A(n20939), .B(n20938), .Z(n20941) );
  NANDN U21360 ( .A(n20940), .B(n20941), .Z(n20943) );
  NAND U21361 ( .A(b[2]), .B(a[30]), .Z(n21324) );
  XNOR U21362 ( .A(n20941), .B(n20940), .Z(n21325) );
  NANDN U21363 ( .A(n21324), .B(n21325), .Z(n20942) );
  NAND U21364 ( .A(n20943), .B(n20942), .Z(n20944) );
  OR U21365 ( .A(n20945), .B(n20944), .Z(n20949) );
  XNOR U21366 ( .A(n20945), .B(n20944), .Z(n21330) );
  XOR U21367 ( .A(n20947), .B(n20946), .Z(n21331) );
  NANDN U21368 ( .A(n21330), .B(n21331), .Z(n20948) );
  NAND U21369 ( .A(n20949), .B(n20948), .Z(n20952) );
  XOR U21370 ( .A(n20951), .B(n20950), .Z(n20953) );
  NANDN U21371 ( .A(n20952), .B(n20953), .Z(n20955) );
  NAND U21372 ( .A(a[32]), .B(b[2]), .Z(n21336) );
  XNOR U21373 ( .A(n20953), .B(n20952), .Z(n21337) );
  NANDN U21374 ( .A(n21336), .B(n21337), .Z(n20954) );
  NAND U21375 ( .A(n20955), .B(n20954), .Z(n20956) );
  OR U21376 ( .A(n20957), .B(n20956), .Z(n20961) );
  XNOR U21377 ( .A(n20957), .B(n20956), .Z(n21342) );
  XOR U21378 ( .A(n20959), .B(n20958), .Z(n21343) );
  NANDN U21379 ( .A(n21342), .B(n21343), .Z(n20960) );
  NAND U21380 ( .A(n20961), .B(n20960), .Z(n20964) );
  XOR U21381 ( .A(n20963), .B(n20962), .Z(n20965) );
  NANDN U21382 ( .A(n20964), .B(n20965), .Z(n20967) );
  NAND U21383 ( .A(a[34]), .B(b[2]), .Z(n21348) );
  XNOR U21384 ( .A(n20965), .B(n20964), .Z(n21349) );
  NANDN U21385 ( .A(n21348), .B(n21349), .Z(n20966) );
  NAND U21386 ( .A(n20967), .B(n20966), .Z(n20968) );
  OR U21387 ( .A(n20969), .B(n20968), .Z(n20973) );
  XNOR U21388 ( .A(n20969), .B(n20968), .Z(n21354) );
  XOR U21389 ( .A(n20971), .B(n20970), .Z(n21355) );
  NANDN U21390 ( .A(n21354), .B(n21355), .Z(n20972) );
  NAND U21391 ( .A(n20973), .B(n20972), .Z(n20976) );
  XOR U21392 ( .A(n20975), .B(n20974), .Z(n20977) );
  NANDN U21393 ( .A(n20976), .B(n20977), .Z(n20979) );
  NAND U21394 ( .A(a[36]), .B(b[2]), .Z(n21360) );
  XNOR U21395 ( .A(n20977), .B(n20976), .Z(n21361) );
  NANDN U21396 ( .A(n21360), .B(n21361), .Z(n20978) );
  NAND U21397 ( .A(n20979), .B(n20978), .Z(n20980) );
  OR U21398 ( .A(n20981), .B(n20980), .Z(n20985) );
  XNOR U21399 ( .A(n20981), .B(n20980), .Z(n21366) );
  XOR U21400 ( .A(n20983), .B(n20982), .Z(n21367) );
  NANDN U21401 ( .A(n21366), .B(n21367), .Z(n20984) );
  NAND U21402 ( .A(n20985), .B(n20984), .Z(n20988) );
  XOR U21403 ( .A(n20987), .B(n20986), .Z(n20989) );
  NANDN U21404 ( .A(n20988), .B(n20989), .Z(n20991) );
  NAND U21405 ( .A(a[38]), .B(b[2]), .Z(n21372) );
  XNOR U21406 ( .A(n20989), .B(n20988), .Z(n21373) );
  NANDN U21407 ( .A(n21372), .B(n21373), .Z(n20990) );
  NAND U21408 ( .A(n20991), .B(n20990), .Z(n20992) );
  OR U21409 ( .A(n20993), .B(n20992), .Z(n20997) );
  XNOR U21410 ( .A(n20993), .B(n20992), .Z(n21378) );
  XOR U21411 ( .A(n20995), .B(n20994), .Z(n21379) );
  NANDN U21412 ( .A(n21378), .B(n21379), .Z(n20996) );
  NAND U21413 ( .A(n20997), .B(n20996), .Z(n21000) );
  XOR U21414 ( .A(n20999), .B(n20998), .Z(n21001) );
  NANDN U21415 ( .A(n21000), .B(n21001), .Z(n21003) );
  NAND U21416 ( .A(a[40]), .B(b[2]), .Z(n21384) );
  XNOR U21417 ( .A(n21001), .B(n21000), .Z(n21385) );
  NANDN U21418 ( .A(n21384), .B(n21385), .Z(n21002) );
  NAND U21419 ( .A(n21003), .B(n21002), .Z(n21004) );
  OR U21420 ( .A(n21005), .B(n21004), .Z(n21009) );
  XNOR U21421 ( .A(n21005), .B(n21004), .Z(n21390) );
  XOR U21422 ( .A(n21007), .B(n21006), .Z(n21391) );
  NANDN U21423 ( .A(n21390), .B(n21391), .Z(n21008) );
  NAND U21424 ( .A(n21009), .B(n21008), .Z(n21012) );
  XOR U21425 ( .A(n21011), .B(n21010), .Z(n21013) );
  NANDN U21426 ( .A(n21012), .B(n21013), .Z(n21015) );
  NAND U21427 ( .A(a[42]), .B(b[2]), .Z(n21396) );
  XNOR U21428 ( .A(n21013), .B(n21012), .Z(n21397) );
  NANDN U21429 ( .A(n21396), .B(n21397), .Z(n21014) );
  NAND U21430 ( .A(n21015), .B(n21014), .Z(n21016) );
  OR U21431 ( .A(n21017), .B(n21016), .Z(n21021) );
  XNOR U21432 ( .A(n21017), .B(n21016), .Z(n21402) );
  XOR U21433 ( .A(n21019), .B(n21018), .Z(n21403) );
  NANDN U21434 ( .A(n21402), .B(n21403), .Z(n21020) );
  NAND U21435 ( .A(n21021), .B(n21020), .Z(n21024) );
  XOR U21436 ( .A(n21023), .B(n21022), .Z(n21025) );
  NANDN U21437 ( .A(n21024), .B(n21025), .Z(n21027) );
  NAND U21438 ( .A(a[44]), .B(b[2]), .Z(n21408) );
  XNOR U21439 ( .A(n21025), .B(n21024), .Z(n21409) );
  NANDN U21440 ( .A(n21408), .B(n21409), .Z(n21026) );
  NAND U21441 ( .A(n21027), .B(n21026), .Z(n21028) );
  OR U21442 ( .A(n21029), .B(n21028), .Z(n21033) );
  XNOR U21443 ( .A(n21029), .B(n21028), .Z(n21414) );
  XOR U21444 ( .A(n21031), .B(n21030), .Z(n21415) );
  NANDN U21445 ( .A(n21414), .B(n21415), .Z(n21032) );
  NAND U21446 ( .A(n21033), .B(n21032), .Z(n21036) );
  XOR U21447 ( .A(n21035), .B(n21034), .Z(n21037) );
  NANDN U21448 ( .A(n21036), .B(n21037), .Z(n21039) );
  NAND U21449 ( .A(a[46]), .B(b[2]), .Z(n21420) );
  XNOR U21450 ( .A(n21037), .B(n21036), .Z(n21421) );
  NANDN U21451 ( .A(n21420), .B(n21421), .Z(n21038) );
  NAND U21452 ( .A(n21039), .B(n21038), .Z(n21040) );
  OR U21453 ( .A(n21041), .B(n21040), .Z(n21045) );
  XNOR U21454 ( .A(n21041), .B(n21040), .Z(n21426) );
  XOR U21455 ( .A(n21043), .B(n21042), .Z(n21427) );
  NANDN U21456 ( .A(n21426), .B(n21427), .Z(n21044) );
  NAND U21457 ( .A(n21045), .B(n21044), .Z(n21048) );
  XOR U21458 ( .A(n21047), .B(n21046), .Z(n21049) );
  NANDN U21459 ( .A(n21048), .B(n21049), .Z(n21051) );
  NAND U21460 ( .A(a[48]), .B(b[2]), .Z(n21432) );
  XNOR U21461 ( .A(n21049), .B(n21048), .Z(n21433) );
  NANDN U21462 ( .A(n21432), .B(n21433), .Z(n21050) );
  NAND U21463 ( .A(n21051), .B(n21050), .Z(n21052) );
  OR U21464 ( .A(n21053), .B(n21052), .Z(n21057) );
  XNOR U21465 ( .A(n21053), .B(n21052), .Z(n21438) );
  XOR U21466 ( .A(n21055), .B(n21054), .Z(n21439) );
  NANDN U21467 ( .A(n21438), .B(n21439), .Z(n21056) );
  NAND U21468 ( .A(n21057), .B(n21056), .Z(n21060) );
  XOR U21469 ( .A(n21059), .B(n21058), .Z(n21061) );
  NANDN U21470 ( .A(n21060), .B(n21061), .Z(n21063) );
  NAND U21471 ( .A(a[50]), .B(b[2]), .Z(n21444) );
  XNOR U21472 ( .A(n21061), .B(n21060), .Z(n21445) );
  NANDN U21473 ( .A(n21444), .B(n21445), .Z(n21062) );
  NAND U21474 ( .A(n21063), .B(n21062), .Z(n21064) );
  OR U21475 ( .A(n21065), .B(n21064), .Z(n21069) );
  XNOR U21476 ( .A(n21065), .B(n21064), .Z(n21450) );
  XOR U21477 ( .A(n21067), .B(n21066), .Z(n21451) );
  NANDN U21478 ( .A(n21450), .B(n21451), .Z(n21068) );
  NAND U21479 ( .A(n21069), .B(n21068), .Z(n21072) );
  XOR U21480 ( .A(n21071), .B(n21070), .Z(n21073) );
  NANDN U21481 ( .A(n21072), .B(n21073), .Z(n21075) );
  NAND U21482 ( .A(a[52]), .B(b[2]), .Z(n21456) );
  XNOR U21483 ( .A(n21073), .B(n21072), .Z(n21457) );
  NANDN U21484 ( .A(n21456), .B(n21457), .Z(n21074) );
  NAND U21485 ( .A(n21075), .B(n21074), .Z(n21076) );
  OR U21486 ( .A(n21077), .B(n21076), .Z(n21081) );
  XNOR U21487 ( .A(n21077), .B(n21076), .Z(n21462) );
  XOR U21488 ( .A(n21079), .B(n21078), .Z(n21463) );
  NANDN U21489 ( .A(n21462), .B(n21463), .Z(n21080) );
  NAND U21490 ( .A(n21081), .B(n21080), .Z(n21084) );
  XOR U21491 ( .A(n21083), .B(n21082), .Z(n21085) );
  NANDN U21492 ( .A(n21084), .B(n21085), .Z(n21087) );
  NAND U21493 ( .A(a[54]), .B(b[2]), .Z(n21468) );
  XNOR U21494 ( .A(n21085), .B(n21084), .Z(n21469) );
  NANDN U21495 ( .A(n21468), .B(n21469), .Z(n21086) );
  NAND U21496 ( .A(n21087), .B(n21086), .Z(n21088) );
  OR U21497 ( .A(n21089), .B(n21088), .Z(n21093) );
  XNOR U21498 ( .A(n21089), .B(n21088), .Z(n21474) );
  XOR U21499 ( .A(n21091), .B(n21090), .Z(n21475) );
  NANDN U21500 ( .A(n21474), .B(n21475), .Z(n21092) );
  NAND U21501 ( .A(n21093), .B(n21092), .Z(n21096) );
  XOR U21502 ( .A(n21095), .B(n21094), .Z(n21097) );
  NANDN U21503 ( .A(n21096), .B(n21097), .Z(n21099) );
  NAND U21504 ( .A(a[56]), .B(b[2]), .Z(n21480) );
  XNOR U21505 ( .A(n21097), .B(n21096), .Z(n21481) );
  NANDN U21506 ( .A(n21480), .B(n21481), .Z(n21098) );
  NAND U21507 ( .A(n21099), .B(n21098), .Z(n21100) );
  OR U21508 ( .A(n21101), .B(n21100), .Z(n21105) );
  XNOR U21509 ( .A(n21101), .B(n21100), .Z(n21486) );
  XOR U21510 ( .A(n21103), .B(n21102), .Z(n21487) );
  NANDN U21511 ( .A(n21486), .B(n21487), .Z(n21104) );
  NAND U21512 ( .A(n21105), .B(n21104), .Z(n21108) );
  XOR U21513 ( .A(n21107), .B(n21106), .Z(n21109) );
  NANDN U21514 ( .A(n21108), .B(n21109), .Z(n21111) );
  NAND U21515 ( .A(a[58]), .B(b[2]), .Z(n21492) );
  XNOR U21516 ( .A(n21109), .B(n21108), .Z(n21493) );
  NANDN U21517 ( .A(n21492), .B(n21493), .Z(n21110) );
  NAND U21518 ( .A(n21111), .B(n21110), .Z(n21112) );
  OR U21519 ( .A(n21113), .B(n21112), .Z(n21117) );
  XNOR U21520 ( .A(n21113), .B(n21112), .Z(n21498) );
  XOR U21521 ( .A(n21115), .B(n21114), .Z(n21499) );
  NANDN U21522 ( .A(n21498), .B(n21499), .Z(n21116) );
  NAND U21523 ( .A(n21117), .B(n21116), .Z(n21120) );
  XNOR U21524 ( .A(n21119), .B(n21118), .Z(n21121) );
  OR U21525 ( .A(n21120), .B(n21121), .Z(n21123) );
  XNOR U21526 ( .A(n21121), .B(n21120), .Z(n21507) );
  NAND U21527 ( .A(a[60]), .B(b[2]), .Z(n21506) );
  OR U21528 ( .A(n21507), .B(n21506), .Z(n21122) );
  NAND U21529 ( .A(n21123), .B(n21122), .Z(n21126) );
  ANDN U21530 ( .B(b[2]), .A(n209), .Z(n21127) );
  OR U21531 ( .A(n21126), .B(n21127), .Z(n21129) );
  XOR U21532 ( .A(n21125), .B(n21124), .Z(n21511) );
  XOR U21533 ( .A(n21127), .B(n21126), .Z(n21510) );
  NANDN U21534 ( .A(n21511), .B(n21510), .Z(n21128) );
  NAND U21535 ( .A(n21129), .B(n21128), .Z(n21131) );
  AND U21536 ( .A(a[62]), .B(b[2]), .Z(n21130) );
  NANDN U21537 ( .A(n21131), .B(n21130), .Z(n21135) );
  XNOR U21538 ( .A(n21131), .B(n21130), .Z(n21516) );
  NAND U21539 ( .A(n21516), .B(n21517), .Z(n21134) );
  AND U21540 ( .A(n21135), .B(n21134), .Z(n21523) );
  XNOR U21541 ( .A(n21137), .B(n21136), .Z(n21138) );
  XNOR U21542 ( .A(n21139), .B(n21138), .Z(n21522) );
  NAND U21543 ( .A(b[2]), .B(a[63]), .Z(n21525) );
  XOR U21544 ( .A(n21141), .B(n21140), .Z(n21144) );
  AND U21545 ( .A(n21145), .B(n21144), .Z(n24092) );
  XNOR U21546 ( .A(n21143), .B(n21142), .Z(n21917) );
  AND U21547 ( .A(n24092), .B(n21917), .Z(n24100) );
  XNOR U21548 ( .A(n21145), .B(n21144), .Z(n24091) );
  ANDN U21549 ( .B(b[1]), .A(n207), .Z(n21495) );
  ANDN U21550 ( .B(b[1]), .A(n205), .Z(n21483) );
  ANDN U21551 ( .B(b[1]), .A(n203), .Z(n21471) );
  ANDN U21552 ( .B(b[1]), .A(n201), .Z(n21459) );
  ANDN U21553 ( .B(b[1]), .A(n199), .Z(n21447) );
  ANDN U21554 ( .B(b[1]), .A(n197), .Z(n21435) );
  ANDN U21555 ( .B(b[1]), .A(n195), .Z(n21423) );
  ANDN U21556 ( .B(b[1]), .A(n193), .Z(n21411) );
  ANDN U21557 ( .B(b[1]), .A(n191), .Z(n21399) );
  ANDN U21558 ( .B(b[1]), .A(n189), .Z(n21387) );
  ANDN U21559 ( .B(b[1]), .A(n187), .Z(n21375) );
  ANDN U21560 ( .B(b[1]), .A(n21772), .Z(n21363) );
  ANDN U21561 ( .B(b[1]), .A(n184), .Z(n21351) );
  ANDN U21562 ( .B(b[1]), .A(n21751), .Z(n21339) );
  NAND U21563 ( .A(a[31]), .B(b[1]), .Z(n21327) );
  ANDN U21564 ( .B(b[1]), .A(n21727), .Z(n21315) );
  NAND U21565 ( .A(a[27]), .B(b[1]), .Z(n21305) );
  XOR U21566 ( .A(n21149), .B(n21148), .Z(n21299) );
  ANDN U21567 ( .B(b[1]), .A(n21703), .Z(n21295) );
  NAND U21568 ( .A(a[24]), .B(b[1]), .Z(n21289) );
  NAND U21569 ( .A(a[23]), .B(b[1]), .Z(n21283) );
  ANDN U21570 ( .B(b[1]), .A(n21681), .Z(n21271) );
  NAND U21571 ( .A(a[20]), .B(b[1]), .Z(n21152) );
  XOR U21572 ( .A(n21151), .B(n21150), .Z(n21153) );
  NANDN U21573 ( .A(n21152), .B(n21153), .Z(n21267) );
  XOR U21574 ( .A(n21153), .B(n21152), .Z(n21684) );
  NAND U21575 ( .A(a[19]), .B(b[1]), .Z(n21263) );
  NAND U21576 ( .A(a[18]), .B(b[1]), .Z(n21257) );
  XOR U21577 ( .A(n21155), .B(n21154), .Z(n21256) );
  NANDN U21578 ( .A(n21257), .B(n21256), .Z(n21259) );
  NAND U21579 ( .A(a[17]), .B(b[1]), .Z(n21253) );
  NAND U21580 ( .A(a[16]), .B(b[1]), .Z(n21246) );
  XOR U21581 ( .A(n21157), .B(n21156), .Z(n21247) );
  OR U21582 ( .A(n21246), .B(n21247), .Z(n21249) );
  ANDN U21583 ( .B(b[1]), .A(n172), .Z(n21243) );
  NAND U21584 ( .A(a[14]), .B(b[1]), .Z(n21236) );
  XNOR U21585 ( .A(n21159), .B(n21158), .Z(n21237) );
  OR U21586 ( .A(n21236), .B(n21237), .Z(n21239) );
  ANDN U21587 ( .B(b[1]), .A(n170), .Z(n21233) );
  NAND U21588 ( .A(a[12]), .B(b[1]), .Z(n21162) );
  XOR U21589 ( .A(n21161), .B(n21160), .Z(n21163) );
  NANDN U21590 ( .A(n21162), .B(n21163), .Z(n21229) );
  XOR U21591 ( .A(n21163), .B(n21162), .Z(n21643) );
  ANDN U21592 ( .B(b[1]), .A(n21164), .Z(n21222) );
  NAND U21593 ( .A(b[2]), .B(a[1]), .Z(n21167) );
  AND U21594 ( .A(b[1]), .B(a[0]), .Z(n24341) );
  NANDN U21595 ( .A(n21167), .B(n24341), .Z(n21166) );
  NAND U21596 ( .A(b[1]), .B(a[2]), .Z(n21165) );
  AND U21597 ( .A(n21166), .B(n21165), .Z(n21173) );
  NANDN U21598 ( .A(n21167), .B(a[0]), .Z(n21168) );
  XNOR U21599 ( .A(a[2]), .B(n21168), .Z(n21169) );
  NAND U21600 ( .A(b[1]), .B(n21169), .Z(n21583) );
  AND U21601 ( .A(a[1]), .B(b[2]), .Z(n21170) );
  XNOR U21602 ( .A(n21171), .B(n21170), .Z(n21584) );
  NANDN U21603 ( .A(n21583), .B(n21584), .Z(n21172) );
  NANDN U21604 ( .A(n21173), .B(n21172), .Z(n21175) );
  NANDN U21605 ( .A(n150), .B(a[3]), .Z(n21174) );
  NAND U21606 ( .A(n21175), .B(n21174), .Z(n21179) );
  XNOR U21607 ( .A(n21175), .B(n21174), .Z(n21588) );
  XNOR U21608 ( .A(n21177), .B(n21176), .Z(n21587) );
  NANDN U21609 ( .A(n21588), .B(n21587), .Z(n21178) );
  NAND U21610 ( .A(n21179), .B(n21178), .Z(n21182) );
  XOR U21611 ( .A(n21181), .B(n21180), .Z(n21183) );
  NANDN U21612 ( .A(n21182), .B(n21183), .Z(n21185) );
  NAND U21613 ( .A(a[4]), .B(b[1]), .Z(n21595) );
  XNOR U21614 ( .A(n21183), .B(n21182), .Z(n21596) );
  NANDN U21615 ( .A(n21595), .B(n21596), .Z(n21184) );
  NAND U21616 ( .A(n21185), .B(n21184), .Z(n21188) );
  AND U21617 ( .A(a[5]), .B(b[1]), .Z(n21189) );
  OR U21618 ( .A(n21188), .B(n21189), .Z(n21191) );
  XOR U21619 ( .A(n21187), .B(n21186), .Z(n21571) );
  XOR U21620 ( .A(n21189), .B(n21188), .Z(n21570) );
  NAND U21621 ( .A(n21571), .B(n21570), .Z(n21190) );
  NAND U21622 ( .A(n21191), .B(n21190), .Z(n21195) );
  XOR U21623 ( .A(n21193), .B(n21192), .Z(n21194) );
  NAND U21624 ( .A(n21195), .B(n21194), .Z(n21197) );
  XNOR U21625 ( .A(n21195), .B(n21194), .Z(n21605) );
  AND U21626 ( .A(a[6]), .B(b[1]), .Z(n21606) );
  OR U21627 ( .A(n21605), .B(n21606), .Z(n21196) );
  NAND U21628 ( .A(n21197), .B(n21196), .Z(n21199) );
  NANDN U21629 ( .A(n150), .B(a[7]), .Z(n21198) );
  NAND U21630 ( .A(n21199), .B(n21198), .Z(n21203) );
  XNOR U21631 ( .A(n21199), .B(n21198), .Z(n21610) );
  XOR U21632 ( .A(n21201), .B(n21200), .Z(n21609) );
  NANDN U21633 ( .A(n21610), .B(n21609), .Z(n21202) );
  NAND U21634 ( .A(n21203), .B(n21202), .Z(n21206) );
  XNOR U21635 ( .A(n21205), .B(n21204), .Z(n21207) );
  NANDN U21636 ( .A(n21206), .B(n21207), .Z(n21209) );
  XOR U21637 ( .A(n21207), .B(n21206), .Z(n21619) );
  NAND U21638 ( .A(a[8]), .B(b[1]), .Z(n21618) );
  OR U21639 ( .A(n21619), .B(n21618), .Z(n21208) );
  NAND U21640 ( .A(n21209), .B(n21208), .Z(n21212) );
  AND U21641 ( .A(a[9]), .B(b[1]), .Z(n21213) );
  OR U21642 ( .A(n21212), .B(n21213), .Z(n21215) );
  XNOR U21643 ( .A(n21211), .B(n21210), .Z(n21623) );
  XOR U21644 ( .A(n21213), .B(n21212), .Z(n21622) );
  NANDN U21645 ( .A(n21623), .B(n21622), .Z(n21214) );
  AND U21646 ( .A(n21215), .B(n21214), .Z(n21219) );
  XOR U21647 ( .A(n21217), .B(n21216), .Z(n21218) );
  NANDN U21648 ( .A(n21219), .B(n21218), .Z(n21221) );
  XOR U21649 ( .A(n21219), .B(n21218), .Z(n21629) );
  ANDN U21650 ( .B(b[1]), .A(n168), .Z(n21628) );
  OR U21651 ( .A(n21629), .B(n21628), .Z(n21220) );
  NAND U21652 ( .A(n21221), .B(n21220), .Z(n21223) );
  NANDN U21653 ( .A(n21222), .B(n21223), .Z(n21227) );
  XOR U21654 ( .A(n21223), .B(n21222), .Z(n21635) );
  XOR U21655 ( .A(n21225), .B(n21224), .Z(n21634) );
  NANDN U21656 ( .A(n21635), .B(n21634), .Z(n21226) );
  NAND U21657 ( .A(n21227), .B(n21226), .Z(n21642) );
  OR U21658 ( .A(n21643), .B(n21642), .Z(n21228) );
  NAND U21659 ( .A(n21229), .B(n21228), .Z(n21232) );
  OR U21660 ( .A(n21233), .B(n21232), .Z(n21235) );
  XOR U21661 ( .A(n21231), .B(n21230), .Z(n21569) );
  XOR U21662 ( .A(n21233), .B(n21232), .Z(n21568) );
  NAND U21663 ( .A(n21569), .B(n21568), .Z(n21234) );
  NAND U21664 ( .A(n21235), .B(n21234), .Z(n21652) );
  XOR U21665 ( .A(n21237), .B(n21236), .Z(n21653) );
  NANDN U21666 ( .A(n21652), .B(n21653), .Z(n21238) );
  NAND U21667 ( .A(n21239), .B(n21238), .Z(n21242) );
  OR U21668 ( .A(n21243), .B(n21242), .Z(n21245) );
  XOR U21669 ( .A(n21243), .B(n21242), .Z(n21566) );
  NANDN U21670 ( .A(n21567), .B(n21566), .Z(n21244) );
  NAND U21671 ( .A(n21245), .B(n21244), .Z(n21662) );
  XOR U21672 ( .A(n21247), .B(n21246), .Z(n21663) );
  NANDN U21673 ( .A(n21662), .B(n21663), .Z(n21248) );
  NAND U21674 ( .A(n21249), .B(n21248), .Z(n21252) );
  NANDN U21675 ( .A(n21253), .B(n21252), .Z(n21255) );
  XOR U21676 ( .A(n21251), .B(n21250), .Z(n21564) );
  NANDN U21677 ( .A(n21564), .B(n21565), .Z(n21254) );
  NAND U21678 ( .A(n21255), .B(n21254), .Z(n21674) );
  NAND U21679 ( .A(n21674), .B(n21673), .Z(n21258) );
  NAND U21680 ( .A(n21259), .B(n21258), .Z(n21262) );
  NANDN U21681 ( .A(n21263), .B(n21262), .Z(n21265) );
  XOR U21682 ( .A(n21261), .B(n21260), .Z(n21562) );
  NANDN U21683 ( .A(n21562), .B(n21563), .Z(n21264) );
  NAND U21684 ( .A(n21265), .B(n21264), .Z(n21685) );
  NANDN U21685 ( .A(n21684), .B(n21685), .Z(n21266) );
  NAND U21686 ( .A(n21267), .B(n21266), .Z(n21270) );
  OR U21687 ( .A(n21271), .B(n21270), .Z(n21273) );
  XOR U21688 ( .A(n21269), .B(n21268), .Z(n21561) );
  XOR U21689 ( .A(n21271), .B(n21270), .Z(n21560) );
  NAND U21690 ( .A(n21561), .B(n21560), .Z(n21272) );
  NAND U21691 ( .A(n21273), .B(n21272), .Z(n21276) );
  XOR U21692 ( .A(n21275), .B(n21274), .Z(n21277) );
  NANDN U21693 ( .A(n21276), .B(n21277), .Z(n21279) );
  XOR U21694 ( .A(n21277), .B(n21276), .Z(n21696) );
  NAND U21695 ( .A(a[22]), .B(b[1]), .Z(n21695) );
  OR U21696 ( .A(n21696), .B(n21695), .Z(n21278) );
  NAND U21697 ( .A(n21279), .B(n21278), .Z(n21282) );
  NANDN U21698 ( .A(n21283), .B(n21282), .Z(n21285) );
  XOR U21699 ( .A(n21281), .B(n21280), .Z(n21558) );
  NANDN U21700 ( .A(n21558), .B(n21559), .Z(n21284) );
  NAND U21701 ( .A(n21285), .B(n21284), .Z(n21288) );
  NANDN U21702 ( .A(n21289), .B(n21288), .Z(n21291) );
  NAND U21703 ( .A(n21706), .B(n21707), .Z(n21290) );
  NAND U21704 ( .A(n21291), .B(n21290), .Z(n21294) );
  OR U21705 ( .A(n21295), .B(n21294), .Z(n21297) );
  XNOR U21706 ( .A(n21293), .B(n21292), .Z(n21711) );
  XOR U21707 ( .A(n21295), .B(n21294), .Z(n21710) );
  NANDN U21708 ( .A(n21711), .B(n21710), .Z(n21296) );
  AND U21709 ( .A(n21297), .B(n21296), .Z(n21298) );
  OR U21710 ( .A(n21299), .B(n21298), .Z(n21301) );
  ANDN U21711 ( .B(b[1]), .A(n179), .Z(n21720) );
  XOR U21712 ( .A(n21299), .B(n21298), .Z(n21719) );
  NANDN U21713 ( .A(n21720), .B(n21719), .Z(n21300) );
  AND U21714 ( .A(n21301), .B(n21300), .Z(n21304) );
  NANDN U21715 ( .A(n21305), .B(n21304), .Z(n21307) );
  XOR U21716 ( .A(n21303), .B(n21302), .Z(n21556) );
  NANDN U21717 ( .A(n21556), .B(n21557), .Z(n21306) );
  AND U21718 ( .A(n21307), .B(n21306), .Z(n21311) );
  XOR U21719 ( .A(n21309), .B(n21308), .Z(n21310) );
  NANDN U21720 ( .A(n21311), .B(n21310), .Z(n21313) );
  NAND U21721 ( .A(a[28]), .B(b[1]), .Z(n21730) );
  NANDN U21722 ( .A(n21730), .B(n21731), .Z(n21312) );
  NAND U21723 ( .A(n21313), .B(n21312), .Z(n21314) );
  OR U21724 ( .A(n21315), .B(n21314), .Z(n21319) );
  XOR U21725 ( .A(n21315), .B(n21314), .Z(n21734) );
  XOR U21726 ( .A(n21317), .B(n21316), .Z(n21735) );
  NAND U21727 ( .A(n21734), .B(n21735), .Z(n21318) );
  AND U21728 ( .A(n21319), .B(n21318), .Z(n21320) );
  OR U21729 ( .A(n21321), .B(n21320), .Z(n21323) );
  ANDN U21730 ( .B(b[1]), .A(n181), .Z(n21742) );
  XOR U21731 ( .A(n21321), .B(n21320), .Z(n21741) );
  NANDN U21732 ( .A(n21742), .B(n21741), .Z(n21322) );
  AND U21733 ( .A(n21323), .B(n21322), .Z(n21326) );
  NANDN U21734 ( .A(n21327), .B(n21326), .Z(n21329) );
  XOR U21735 ( .A(n21325), .B(n21324), .Z(n21554) );
  NANDN U21736 ( .A(n21554), .B(n21555), .Z(n21328) );
  AND U21737 ( .A(n21329), .B(n21328), .Z(n21332) );
  XOR U21738 ( .A(n21331), .B(n21330), .Z(n21333) );
  NANDN U21739 ( .A(n21332), .B(n21333), .Z(n21335) );
  XOR U21740 ( .A(n21333), .B(n21332), .Z(n21755) );
  NAND U21741 ( .A(a[32]), .B(b[1]), .Z(n21754) );
  OR U21742 ( .A(n21755), .B(n21754), .Z(n21334) );
  NAND U21743 ( .A(n21335), .B(n21334), .Z(n21338) );
  OR U21744 ( .A(n21339), .B(n21338), .Z(n21341) );
  XOR U21745 ( .A(n21337), .B(n21336), .Z(n21553) );
  XOR U21746 ( .A(n21339), .B(n21338), .Z(n21552) );
  NAND U21747 ( .A(n21553), .B(n21552), .Z(n21340) );
  NAND U21748 ( .A(n21341), .B(n21340), .Z(n21344) );
  XOR U21749 ( .A(n21343), .B(n21342), .Z(n21345) );
  NANDN U21750 ( .A(n21344), .B(n21345), .Z(n21347) );
  XOR U21751 ( .A(n21345), .B(n21344), .Z(n21765) );
  NAND U21752 ( .A(a[34]), .B(b[1]), .Z(n21764) );
  OR U21753 ( .A(n21765), .B(n21764), .Z(n21346) );
  NAND U21754 ( .A(n21347), .B(n21346), .Z(n21350) );
  OR U21755 ( .A(n21351), .B(n21350), .Z(n21353) );
  XOR U21756 ( .A(n21349), .B(n21348), .Z(n21551) );
  XOR U21757 ( .A(n21351), .B(n21350), .Z(n21550) );
  NAND U21758 ( .A(n21551), .B(n21550), .Z(n21352) );
  NAND U21759 ( .A(n21353), .B(n21352), .Z(n21356) );
  XOR U21760 ( .A(n21355), .B(n21354), .Z(n21357) );
  NANDN U21761 ( .A(n21356), .B(n21357), .Z(n21359) );
  XOR U21762 ( .A(n21357), .B(n21356), .Z(n21776) );
  NAND U21763 ( .A(a[36]), .B(b[1]), .Z(n21775) );
  OR U21764 ( .A(n21776), .B(n21775), .Z(n21358) );
  NAND U21765 ( .A(n21359), .B(n21358), .Z(n21362) );
  OR U21766 ( .A(n21363), .B(n21362), .Z(n21365) );
  XOR U21767 ( .A(n21361), .B(n21360), .Z(n21549) );
  XOR U21768 ( .A(n21363), .B(n21362), .Z(n21548) );
  NAND U21769 ( .A(n21549), .B(n21548), .Z(n21364) );
  NAND U21770 ( .A(n21365), .B(n21364), .Z(n21368) );
  XOR U21771 ( .A(n21367), .B(n21366), .Z(n21369) );
  NANDN U21772 ( .A(n21368), .B(n21369), .Z(n21371) );
  XOR U21773 ( .A(n21369), .B(n21368), .Z(n21786) );
  NAND U21774 ( .A(a[38]), .B(b[1]), .Z(n21785) );
  OR U21775 ( .A(n21786), .B(n21785), .Z(n21370) );
  NAND U21776 ( .A(n21371), .B(n21370), .Z(n21374) );
  OR U21777 ( .A(n21375), .B(n21374), .Z(n21377) );
  XOR U21778 ( .A(n21373), .B(n21372), .Z(n21547) );
  XOR U21779 ( .A(n21375), .B(n21374), .Z(n21546) );
  NAND U21780 ( .A(n21547), .B(n21546), .Z(n21376) );
  NAND U21781 ( .A(n21377), .B(n21376), .Z(n21380) );
  XOR U21782 ( .A(n21379), .B(n21378), .Z(n21381) );
  NANDN U21783 ( .A(n21380), .B(n21381), .Z(n21383) );
  XOR U21784 ( .A(n21381), .B(n21380), .Z(n21796) );
  NAND U21785 ( .A(a[40]), .B(b[1]), .Z(n21795) );
  OR U21786 ( .A(n21796), .B(n21795), .Z(n21382) );
  NAND U21787 ( .A(n21383), .B(n21382), .Z(n21386) );
  OR U21788 ( .A(n21387), .B(n21386), .Z(n21389) );
  XOR U21789 ( .A(n21385), .B(n21384), .Z(n21545) );
  XOR U21790 ( .A(n21387), .B(n21386), .Z(n21544) );
  NAND U21791 ( .A(n21545), .B(n21544), .Z(n21388) );
  NAND U21792 ( .A(n21389), .B(n21388), .Z(n21392) );
  XOR U21793 ( .A(n21391), .B(n21390), .Z(n21393) );
  NANDN U21794 ( .A(n21392), .B(n21393), .Z(n21395) );
  XOR U21795 ( .A(n21393), .B(n21392), .Z(n21806) );
  NAND U21796 ( .A(a[42]), .B(b[1]), .Z(n21805) );
  OR U21797 ( .A(n21806), .B(n21805), .Z(n21394) );
  NAND U21798 ( .A(n21395), .B(n21394), .Z(n21398) );
  OR U21799 ( .A(n21399), .B(n21398), .Z(n21401) );
  XOR U21800 ( .A(n21397), .B(n21396), .Z(n21543) );
  XOR U21801 ( .A(n21399), .B(n21398), .Z(n21542) );
  NAND U21802 ( .A(n21543), .B(n21542), .Z(n21400) );
  NAND U21803 ( .A(n21401), .B(n21400), .Z(n21404) );
  XOR U21804 ( .A(n21403), .B(n21402), .Z(n21405) );
  NANDN U21805 ( .A(n21404), .B(n21405), .Z(n21407) );
  XOR U21806 ( .A(n21405), .B(n21404), .Z(n21816) );
  NAND U21807 ( .A(a[44]), .B(b[1]), .Z(n21815) );
  OR U21808 ( .A(n21816), .B(n21815), .Z(n21406) );
  NAND U21809 ( .A(n21407), .B(n21406), .Z(n21410) );
  OR U21810 ( .A(n21411), .B(n21410), .Z(n21413) );
  XOR U21811 ( .A(n21409), .B(n21408), .Z(n21541) );
  XOR U21812 ( .A(n21411), .B(n21410), .Z(n21540) );
  NAND U21813 ( .A(n21541), .B(n21540), .Z(n21412) );
  NAND U21814 ( .A(n21413), .B(n21412), .Z(n21416) );
  XOR U21815 ( .A(n21415), .B(n21414), .Z(n21417) );
  NANDN U21816 ( .A(n21416), .B(n21417), .Z(n21419) );
  XOR U21817 ( .A(n21417), .B(n21416), .Z(n21826) );
  NAND U21818 ( .A(a[46]), .B(b[1]), .Z(n21825) );
  OR U21819 ( .A(n21826), .B(n21825), .Z(n21418) );
  NAND U21820 ( .A(n21419), .B(n21418), .Z(n21422) );
  OR U21821 ( .A(n21423), .B(n21422), .Z(n21425) );
  XOR U21822 ( .A(n21421), .B(n21420), .Z(n21539) );
  XOR U21823 ( .A(n21423), .B(n21422), .Z(n21538) );
  NAND U21824 ( .A(n21539), .B(n21538), .Z(n21424) );
  NAND U21825 ( .A(n21425), .B(n21424), .Z(n21428) );
  XOR U21826 ( .A(n21427), .B(n21426), .Z(n21429) );
  NANDN U21827 ( .A(n21428), .B(n21429), .Z(n21431) );
  XOR U21828 ( .A(n21429), .B(n21428), .Z(n21836) );
  NAND U21829 ( .A(a[48]), .B(b[1]), .Z(n21835) );
  OR U21830 ( .A(n21836), .B(n21835), .Z(n21430) );
  NAND U21831 ( .A(n21431), .B(n21430), .Z(n21434) );
  OR U21832 ( .A(n21435), .B(n21434), .Z(n21437) );
  XOR U21833 ( .A(n21433), .B(n21432), .Z(n21537) );
  XOR U21834 ( .A(n21435), .B(n21434), .Z(n21536) );
  NAND U21835 ( .A(n21537), .B(n21536), .Z(n21436) );
  NAND U21836 ( .A(n21437), .B(n21436), .Z(n21440) );
  XOR U21837 ( .A(n21439), .B(n21438), .Z(n21441) );
  NANDN U21838 ( .A(n21440), .B(n21441), .Z(n21443) );
  XOR U21839 ( .A(n21441), .B(n21440), .Z(n21846) );
  NAND U21840 ( .A(a[50]), .B(b[1]), .Z(n21845) );
  OR U21841 ( .A(n21846), .B(n21845), .Z(n21442) );
  NAND U21842 ( .A(n21443), .B(n21442), .Z(n21446) );
  OR U21843 ( .A(n21447), .B(n21446), .Z(n21449) );
  XOR U21844 ( .A(n21445), .B(n21444), .Z(n21535) );
  XOR U21845 ( .A(n21447), .B(n21446), .Z(n21534) );
  NAND U21846 ( .A(n21535), .B(n21534), .Z(n21448) );
  NAND U21847 ( .A(n21449), .B(n21448), .Z(n21452) );
  XOR U21848 ( .A(n21451), .B(n21450), .Z(n21453) );
  NANDN U21849 ( .A(n21452), .B(n21453), .Z(n21455) );
  XOR U21850 ( .A(n21453), .B(n21452), .Z(n21856) );
  NAND U21851 ( .A(a[52]), .B(b[1]), .Z(n21855) );
  OR U21852 ( .A(n21856), .B(n21855), .Z(n21454) );
  NAND U21853 ( .A(n21455), .B(n21454), .Z(n21458) );
  OR U21854 ( .A(n21459), .B(n21458), .Z(n21461) );
  XOR U21855 ( .A(n21457), .B(n21456), .Z(n21533) );
  XOR U21856 ( .A(n21459), .B(n21458), .Z(n21532) );
  NAND U21857 ( .A(n21533), .B(n21532), .Z(n21460) );
  NAND U21858 ( .A(n21461), .B(n21460), .Z(n21464) );
  XOR U21859 ( .A(n21463), .B(n21462), .Z(n21465) );
  NANDN U21860 ( .A(n21464), .B(n21465), .Z(n21467) );
  XOR U21861 ( .A(n21465), .B(n21464), .Z(n21866) );
  NAND U21862 ( .A(a[54]), .B(b[1]), .Z(n21865) );
  OR U21863 ( .A(n21866), .B(n21865), .Z(n21466) );
  NAND U21864 ( .A(n21467), .B(n21466), .Z(n21470) );
  OR U21865 ( .A(n21471), .B(n21470), .Z(n21473) );
  XOR U21866 ( .A(n21469), .B(n21468), .Z(n21531) );
  XOR U21867 ( .A(n21471), .B(n21470), .Z(n21530) );
  NAND U21868 ( .A(n21531), .B(n21530), .Z(n21472) );
  NAND U21869 ( .A(n21473), .B(n21472), .Z(n21476) );
  XOR U21870 ( .A(n21475), .B(n21474), .Z(n21477) );
  NANDN U21871 ( .A(n21476), .B(n21477), .Z(n21479) );
  XOR U21872 ( .A(n21477), .B(n21476), .Z(n21876) );
  NAND U21873 ( .A(a[56]), .B(b[1]), .Z(n21875) );
  OR U21874 ( .A(n21876), .B(n21875), .Z(n21478) );
  NAND U21875 ( .A(n21479), .B(n21478), .Z(n21482) );
  OR U21876 ( .A(n21483), .B(n21482), .Z(n21485) );
  XOR U21877 ( .A(n21481), .B(n21480), .Z(n21529) );
  XOR U21878 ( .A(n21483), .B(n21482), .Z(n21528) );
  NAND U21879 ( .A(n21529), .B(n21528), .Z(n21484) );
  NAND U21880 ( .A(n21485), .B(n21484), .Z(n21488) );
  XOR U21881 ( .A(n21487), .B(n21486), .Z(n21489) );
  NANDN U21882 ( .A(n21488), .B(n21489), .Z(n21491) );
  XOR U21883 ( .A(n21489), .B(n21488), .Z(n21886) );
  NAND U21884 ( .A(a[58]), .B(b[1]), .Z(n21885) );
  OR U21885 ( .A(n21886), .B(n21885), .Z(n21490) );
  NAND U21886 ( .A(n21491), .B(n21490), .Z(n21494) );
  OR U21887 ( .A(n21495), .B(n21494), .Z(n21497) );
  XOR U21888 ( .A(n21493), .B(n21492), .Z(n21527) );
  XOR U21889 ( .A(n21495), .B(n21494), .Z(n21526) );
  NAND U21890 ( .A(n21527), .B(n21526), .Z(n21496) );
  NAND U21891 ( .A(n21497), .B(n21496), .Z(n21500) );
  XOR U21892 ( .A(n21499), .B(n21498), .Z(n21501) );
  NANDN U21893 ( .A(n21500), .B(n21501), .Z(n21503) );
  XOR U21894 ( .A(n21501), .B(n21500), .Z(n21896) );
  NAND U21895 ( .A(a[60]), .B(b[1]), .Z(n21895) );
  OR U21896 ( .A(n21896), .B(n21895), .Z(n21502) );
  NAND U21897 ( .A(n21503), .B(n21502), .Z(n21504) );
  ANDN U21898 ( .B(b[1]), .A(n209), .Z(n21505) );
  OR U21899 ( .A(n21504), .B(n21505), .Z(n21509) );
  XNOR U21900 ( .A(n21505), .B(n21504), .Z(n21899) );
  XOR U21901 ( .A(n21507), .B(n21506), .Z(n21900) );
  OR U21902 ( .A(n21899), .B(n21900), .Z(n21508) );
  NAND U21903 ( .A(n21509), .B(n21508), .Z(n21512) );
  XNOR U21904 ( .A(n21511), .B(n21510), .Z(n21513) );
  OR U21905 ( .A(n21512), .B(n21513), .Z(n21515) );
  XNOR U21906 ( .A(n21513), .B(n21512), .Z(n21908) );
  NAND U21907 ( .A(a[62]), .B(b[1]), .Z(n21907) );
  OR U21908 ( .A(n21908), .B(n21907), .Z(n21514) );
  NAND U21909 ( .A(n21515), .B(n21514), .Z(n21518) );
  ANDN U21910 ( .B(b[1]), .A(n210), .Z(n21519) );
  OR U21911 ( .A(n21518), .B(n21519), .Z(n21521) );
  XOR U21912 ( .A(n21519), .B(n21518), .Z(n21911) );
  NANDN U21913 ( .A(n21912), .B(n21911), .Z(n21520) );
  AND U21914 ( .A(n21521), .B(n21520), .Z(n21913) );
  XNOR U21915 ( .A(n21523), .B(n21522), .Z(n21524) );
  XNOR U21916 ( .A(n21525), .B(n21524), .Z(n21914) );
  NAND U21917 ( .A(n21913), .B(n21914), .Z(n21916) );
  XNOR U21918 ( .A(n21527), .B(n21526), .Z(n21889) );
  XNOR U21919 ( .A(n21529), .B(n21528), .Z(n21879) );
  XNOR U21920 ( .A(n21531), .B(n21530), .Z(n21869) );
  XNOR U21921 ( .A(n21533), .B(n21532), .Z(n21859) );
  XNOR U21922 ( .A(n21535), .B(n21534), .Z(n21849) );
  XNOR U21923 ( .A(n21537), .B(n21536), .Z(n21839) );
  XNOR U21924 ( .A(n21539), .B(n21538), .Z(n21829) );
  XNOR U21925 ( .A(n21541), .B(n21540), .Z(n21819) );
  XNOR U21926 ( .A(n21543), .B(n21542), .Z(n21809) );
  XNOR U21927 ( .A(n21545), .B(n21544), .Z(n21799) );
  XNOR U21928 ( .A(n21547), .B(n21546), .Z(n21789) );
  XNOR U21929 ( .A(n21549), .B(n21548), .Z(n21779) );
  XNOR U21930 ( .A(n21551), .B(n21550), .Z(n21768) );
  XNOR U21931 ( .A(n21553), .B(n21552), .Z(n21758) );
  XNOR U21932 ( .A(n21555), .B(n21554), .Z(n21747) );
  XNOR U21933 ( .A(n21557), .B(n21556), .Z(n21723) );
  XNOR U21934 ( .A(n21559), .B(n21558), .Z(n21699) );
  XNOR U21935 ( .A(n21561), .B(n21560), .Z(n21688) );
  XNOR U21936 ( .A(n21563), .B(n21562), .Z(n21677) );
  XNOR U21937 ( .A(n21565), .B(n21564), .Z(n21666) );
  XOR U21938 ( .A(n21567), .B(n21566), .Z(n21656) );
  XNOR U21939 ( .A(n21569), .B(n21568), .Z(n21646) );
  AND U21940 ( .A(b[0]), .B(a[11]), .Z(n21630) );
  XNOR U21941 ( .A(n21571), .B(n21570), .Z(n21599) );
  NAND U21942 ( .A(a[2]), .B(b[0]), .Z(n21572) );
  ANDN U21943 ( .B(b[0]), .A(n161), .Z(c[0]) );
  AND U21944 ( .A(a[1]), .B(b[1]), .Z(n21573) );
  AND U21945 ( .A(c[0]), .B(n21573), .Z(n21575) );
  ANDN U21946 ( .B(n21572), .A(n21575), .Z(n21579) );
  XOR U21947 ( .A(n21574), .B(n21573), .Z(n24215) );
  XOR U21948 ( .A(a[2]), .B(n21575), .Z(n21577) );
  NANDN U21949 ( .A(b[0]), .B(a[2]), .Z(n21576) );
  AND U21950 ( .A(n21577), .B(n21576), .Z(n24214) );
  NANDN U21951 ( .A(n24215), .B(n24214), .Z(n21578) );
  NANDN U21952 ( .A(n21579), .B(n21578), .Z(n21582) );
  NANDN U21953 ( .A(n21580), .B(b[0]), .Z(n21581) );
  NAND U21954 ( .A(n21582), .B(n21581), .Z(n21586) );
  XNOR U21955 ( .A(n21582), .B(n21581), .Z(n24237) );
  XNOR U21956 ( .A(n21584), .B(n21583), .Z(n24236) );
  NANDN U21957 ( .A(n24237), .B(n24236), .Z(n21585) );
  NAND U21958 ( .A(n21586), .B(n21585), .Z(n21590) );
  XNOR U21959 ( .A(n21588), .B(n21587), .Z(n21589) );
  NAND U21960 ( .A(n21590), .B(n21589), .Z(n21592) );
  AND U21961 ( .A(b[0]), .B(a[4]), .Z(n24258) );
  XNOR U21962 ( .A(n21590), .B(n21589), .Z(n24259) );
  OR U21963 ( .A(n24258), .B(n24259), .Z(n21591) );
  NAND U21964 ( .A(n21592), .B(n21591), .Z(n21594) );
  NANDN U21965 ( .A(n164), .B(b[0]), .Z(n21593) );
  NAND U21966 ( .A(n21594), .B(n21593), .Z(n21598) );
  XNOR U21967 ( .A(n21594), .B(n21593), .Z(n24281) );
  XNOR U21968 ( .A(n21596), .B(n21595), .Z(n24280) );
  OR U21969 ( .A(n24281), .B(n24280), .Z(n21597) );
  NAND U21970 ( .A(n21598), .B(n21597), .Z(n21600) );
  NANDN U21971 ( .A(n21599), .B(n21600), .Z(n21602) );
  AND U21972 ( .A(b[0]), .B(a[6]), .Z(n24302) );
  XNOR U21973 ( .A(n21600), .B(n21599), .Z(n24303) );
  NANDN U21974 ( .A(n24302), .B(n24303), .Z(n21601) );
  NAND U21975 ( .A(n21602), .B(n21601), .Z(n21604) );
  NANDN U21976 ( .A(n166), .B(b[0]), .Z(n21603) );
  NAND U21977 ( .A(n21604), .B(n21603), .Z(n21608) );
  XNOR U21978 ( .A(n21604), .B(n21603), .Z(n24324) );
  XOR U21979 ( .A(n21606), .B(n21605), .Z(n24325) );
  NANDN U21980 ( .A(n24324), .B(n24325), .Z(n21607) );
  NAND U21981 ( .A(n21608), .B(n21607), .Z(n21612) );
  XNOR U21982 ( .A(n21610), .B(n21609), .Z(n21611) );
  NAND U21983 ( .A(n21612), .B(n21611), .Z(n21614) );
  AND U21984 ( .A(b[0]), .B(a[8]), .Z(n24332) );
  XNOR U21985 ( .A(n21612), .B(n21611), .Z(n24333) );
  OR U21986 ( .A(n24332), .B(n24333), .Z(n21613) );
  NAND U21987 ( .A(n21614), .B(n21613), .Z(n21617) );
  NANDN U21988 ( .A(n21615), .B(b[0]), .Z(n21616) );
  NAND U21989 ( .A(n21617), .B(n21616), .Z(n21621) );
  XNOR U21990 ( .A(n21617), .B(n21616), .Z(n24335) );
  XOR U21991 ( .A(n21619), .B(n21618), .Z(n24334) );
  OR U21992 ( .A(n24335), .B(n24334), .Z(n21620) );
  NAND U21993 ( .A(n21621), .B(n21620), .Z(n21625) );
  XNOR U21994 ( .A(n21623), .B(n21622), .Z(n21624) );
  NAND U21995 ( .A(n21625), .B(n21624), .Z(n21627) );
  AND U21996 ( .A(b[0]), .B(a[10]), .Z(n24336) );
  XNOR U21997 ( .A(n21625), .B(n21624), .Z(n24337) );
  OR U21998 ( .A(n24336), .B(n24337), .Z(n21626) );
  AND U21999 ( .A(n21627), .B(n21626), .Z(n21631) );
  OR U22000 ( .A(n21630), .B(n21631), .Z(n21633) );
  XNOR U22001 ( .A(n21629), .B(n21628), .Z(n24339) );
  XNOR U22002 ( .A(n21631), .B(n21630), .Z(n24338) );
  OR U22003 ( .A(n24339), .B(n24338), .Z(n21632) );
  NAND U22004 ( .A(n21633), .B(n21632), .Z(n21637) );
  NAND U22005 ( .A(n21637), .B(n21636), .Z(n21639) );
  AND U22006 ( .A(b[0]), .B(a[12]), .Z(n24216) );
  XNOR U22007 ( .A(n21637), .B(n21636), .Z(n24217) );
  OR U22008 ( .A(n24216), .B(n24217), .Z(n21638) );
  NAND U22009 ( .A(n21639), .B(n21638), .Z(n21641) );
  NANDN U22010 ( .A(n170), .B(b[0]), .Z(n21640) );
  NAND U22011 ( .A(n21641), .B(n21640), .Z(n21645) );
  XNOR U22012 ( .A(n21641), .B(n21640), .Z(n24219) );
  XOR U22013 ( .A(n21643), .B(n21642), .Z(n24218) );
  OR U22014 ( .A(n24219), .B(n24218), .Z(n21644) );
  NAND U22015 ( .A(n21645), .B(n21644), .Z(n21647) );
  NANDN U22016 ( .A(n21646), .B(n21647), .Z(n21649) );
  AND U22017 ( .A(b[0]), .B(a[14]), .Z(n24220) );
  XNOR U22018 ( .A(n21647), .B(n21646), .Z(n24221) );
  NANDN U22019 ( .A(n24220), .B(n24221), .Z(n21648) );
  NAND U22020 ( .A(n21649), .B(n21648), .Z(n21651) );
  NANDN U22021 ( .A(n172), .B(b[0]), .Z(n21650) );
  NAND U22022 ( .A(n21651), .B(n21650), .Z(n21655) );
  XNOR U22023 ( .A(n21651), .B(n21650), .Z(n24223) );
  XNOR U22024 ( .A(n21653), .B(n21652), .Z(n24222) );
  OR U22025 ( .A(n24223), .B(n24222), .Z(n21654) );
  NAND U22026 ( .A(n21655), .B(n21654), .Z(n21657) );
  NANDN U22027 ( .A(n21656), .B(n21657), .Z(n21659) );
  AND U22028 ( .A(b[0]), .B(a[16]), .Z(n24224) );
  XNOR U22029 ( .A(n21657), .B(n21656), .Z(n24225) );
  NANDN U22030 ( .A(n24224), .B(n24225), .Z(n21658) );
  NAND U22031 ( .A(n21659), .B(n21658), .Z(n21661) );
  NANDN U22032 ( .A(n174), .B(b[0]), .Z(n21660) );
  NAND U22033 ( .A(n21661), .B(n21660), .Z(n21665) );
  XNOR U22034 ( .A(n21661), .B(n21660), .Z(n24227) );
  XNOR U22035 ( .A(n21663), .B(n21662), .Z(n24226) );
  OR U22036 ( .A(n24227), .B(n24226), .Z(n21664) );
  NAND U22037 ( .A(n21665), .B(n21664), .Z(n21667) );
  NANDN U22038 ( .A(n21666), .B(n21667), .Z(n21669) );
  AND U22039 ( .A(b[0]), .B(a[18]), .Z(n24228) );
  XNOR U22040 ( .A(n21667), .B(n21666), .Z(n24229) );
  NANDN U22041 ( .A(n24228), .B(n24229), .Z(n21668) );
  NAND U22042 ( .A(n21669), .B(n21668), .Z(n21672) );
  NANDN U22043 ( .A(n21670), .B(b[0]), .Z(n21671) );
  NAND U22044 ( .A(n21672), .B(n21671), .Z(n21676) );
  XNOR U22045 ( .A(n21672), .B(n21671), .Z(n24231) );
  XOR U22046 ( .A(n21674), .B(n21673), .Z(n24230) );
  OR U22047 ( .A(n24231), .B(n24230), .Z(n21675) );
  NAND U22048 ( .A(n21676), .B(n21675), .Z(n21678) );
  NANDN U22049 ( .A(n21677), .B(n21678), .Z(n21680) );
  AND U22050 ( .A(b[0]), .B(a[20]), .Z(n24232) );
  XNOR U22051 ( .A(n21678), .B(n21677), .Z(n24233) );
  NANDN U22052 ( .A(n24232), .B(n24233), .Z(n21679) );
  NAND U22053 ( .A(n21680), .B(n21679), .Z(n21683) );
  NANDN U22054 ( .A(n21681), .B(b[0]), .Z(n21682) );
  NAND U22055 ( .A(n21683), .B(n21682), .Z(n21687) );
  XNOR U22056 ( .A(n21683), .B(n21682), .Z(n24235) );
  XNOR U22057 ( .A(n21685), .B(n21684), .Z(n24234) );
  OR U22058 ( .A(n24235), .B(n24234), .Z(n21686) );
  NAND U22059 ( .A(n21687), .B(n21686), .Z(n21689) );
  NANDN U22060 ( .A(n21688), .B(n21689), .Z(n21691) );
  AND U22061 ( .A(b[0]), .B(a[22]), .Z(n24238) );
  XNOR U22062 ( .A(n21689), .B(n21688), .Z(n24239) );
  NANDN U22063 ( .A(n24238), .B(n24239), .Z(n21690) );
  NAND U22064 ( .A(n21691), .B(n21690), .Z(n21694) );
  NANDN U22065 ( .A(n21692), .B(b[0]), .Z(n21693) );
  NAND U22066 ( .A(n21694), .B(n21693), .Z(n21698) );
  XNOR U22067 ( .A(n21694), .B(n21693), .Z(n24241) );
  XOR U22068 ( .A(n21696), .B(n21695), .Z(n24240) );
  OR U22069 ( .A(n24241), .B(n24240), .Z(n21697) );
  NAND U22070 ( .A(n21698), .B(n21697), .Z(n21700) );
  NANDN U22071 ( .A(n21699), .B(n21700), .Z(n21702) );
  AND U22072 ( .A(b[0]), .B(a[24]), .Z(n24242) );
  XNOR U22073 ( .A(n21700), .B(n21699), .Z(n24243) );
  NANDN U22074 ( .A(n24242), .B(n24243), .Z(n21701) );
  NAND U22075 ( .A(n21702), .B(n21701), .Z(n21705) );
  NANDN U22076 ( .A(n21703), .B(b[0]), .Z(n21704) );
  NAND U22077 ( .A(n21705), .B(n21704), .Z(n21709) );
  XNOR U22078 ( .A(n21705), .B(n21704), .Z(n24245) );
  XOR U22079 ( .A(n21707), .B(n21706), .Z(n24244) );
  OR U22080 ( .A(n24245), .B(n24244), .Z(n21708) );
  NAND U22081 ( .A(n21709), .B(n21708), .Z(n21713) );
  XNOR U22082 ( .A(n21711), .B(n21710), .Z(n21712) );
  NAND U22083 ( .A(n21713), .B(n21712), .Z(n21715) );
  AND U22084 ( .A(b[0]), .B(a[26]), .Z(n24246) );
  XNOR U22085 ( .A(n21713), .B(n21712), .Z(n24247) );
  OR U22086 ( .A(n24246), .B(n24247), .Z(n21714) );
  NAND U22087 ( .A(n21715), .B(n21714), .Z(n21718) );
  NANDN U22088 ( .A(n21716), .B(b[0]), .Z(n21717) );
  NAND U22089 ( .A(n21718), .B(n21717), .Z(n21722) );
  XNOR U22090 ( .A(n21718), .B(n21717), .Z(n24249) );
  XOR U22091 ( .A(n21720), .B(n21719), .Z(n24248) );
  OR U22092 ( .A(n24249), .B(n24248), .Z(n21721) );
  NAND U22093 ( .A(n21722), .B(n21721), .Z(n21724) );
  NANDN U22094 ( .A(n21723), .B(n21724), .Z(n21726) );
  AND U22095 ( .A(b[0]), .B(a[28]), .Z(n24250) );
  XNOR U22096 ( .A(n21724), .B(n21723), .Z(n24251) );
  NANDN U22097 ( .A(n24250), .B(n24251), .Z(n21725) );
  NAND U22098 ( .A(n21726), .B(n21725), .Z(n21729) );
  NANDN U22099 ( .A(n21727), .B(b[0]), .Z(n21728) );
  NAND U22100 ( .A(n21729), .B(n21728), .Z(n21733) );
  XNOR U22101 ( .A(n21729), .B(n21728), .Z(n24253) );
  XNOR U22102 ( .A(n21731), .B(n21730), .Z(n24252) );
  OR U22103 ( .A(n24253), .B(n24252), .Z(n21732) );
  NAND U22104 ( .A(n21733), .B(n21732), .Z(n21737) );
  NAND U22105 ( .A(n21737), .B(n21736), .Z(n21739) );
  AND U22106 ( .A(b[0]), .B(a[30]), .Z(n24254) );
  XNOR U22107 ( .A(n21737), .B(n21736), .Z(n24255) );
  OR U22108 ( .A(n24254), .B(n24255), .Z(n21738) );
  NAND U22109 ( .A(n21739), .B(n21738), .Z(n21744) );
  NANDN U22110 ( .A(n21740), .B(b[0]), .Z(n21743) );
  NAND U22111 ( .A(n21744), .B(n21743), .Z(n21746) );
  XOR U22112 ( .A(n21742), .B(n21741), .Z(n24257) );
  XNOR U22113 ( .A(n21744), .B(n21743), .Z(n24256) );
  OR U22114 ( .A(n24257), .B(n24256), .Z(n21745) );
  NAND U22115 ( .A(n21746), .B(n21745), .Z(n21748) );
  NANDN U22116 ( .A(n21747), .B(n21748), .Z(n21750) );
  AND U22117 ( .A(b[0]), .B(a[32]), .Z(n24260) );
  XNOR U22118 ( .A(n21748), .B(n21747), .Z(n24261) );
  NANDN U22119 ( .A(n24260), .B(n24261), .Z(n21749) );
  NAND U22120 ( .A(n21750), .B(n21749), .Z(n21753) );
  NANDN U22121 ( .A(n21751), .B(b[0]), .Z(n21752) );
  NAND U22122 ( .A(n21753), .B(n21752), .Z(n21757) );
  XNOR U22123 ( .A(n21753), .B(n21752), .Z(n24263) );
  XOR U22124 ( .A(n21755), .B(n21754), .Z(n24262) );
  OR U22125 ( .A(n24263), .B(n24262), .Z(n21756) );
  NAND U22126 ( .A(n21757), .B(n21756), .Z(n21759) );
  NANDN U22127 ( .A(n21758), .B(n21759), .Z(n21761) );
  AND U22128 ( .A(b[0]), .B(a[34]), .Z(n24264) );
  XNOR U22129 ( .A(n21759), .B(n21758), .Z(n24265) );
  NANDN U22130 ( .A(n24264), .B(n24265), .Z(n21760) );
  NAND U22131 ( .A(n21761), .B(n21760), .Z(n21763) );
  NANDN U22132 ( .A(n184), .B(b[0]), .Z(n21762) );
  NAND U22133 ( .A(n21763), .B(n21762), .Z(n21767) );
  XNOR U22134 ( .A(n21763), .B(n21762), .Z(n24267) );
  XOR U22135 ( .A(n21765), .B(n21764), .Z(n24266) );
  OR U22136 ( .A(n24267), .B(n24266), .Z(n21766) );
  NAND U22137 ( .A(n21767), .B(n21766), .Z(n21769) );
  NANDN U22138 ( .A(n21768), .B(n21769), .Z(n21771) );
  AND U22139 ( .A(b[0]), .B(a[36]), .Z(n24268) );
  XNOR U22140 ( .A(n21769), .B(n21768), .Z(n24269) );
  NANDN U22141 ( .A(n24268), .B(n24269), .Z(n21770) );
  NAND U22142 ( .A(n21771), .B(n21770), .Z(n21774) );
  NANDN U22143 ( .A(n21772), .B(b[0]), .Z(n21773) );
  NAND U22144 ( .A(n21774), .B(n21773), .Z(n21778) );
  XNOR U22145 ( .A(n21774), .B(n21773), .Z(n24271) );
  XOR U22146 ( .A(n21776), .B(n21775), .Z(n24270) );
  OR U22147 ( .A(n24271), .B(n24270), .Z(n21777) );
  NAND U22148 ( .A(n21778), .B(n21777), .Z(n21780) );
  NANDN U22149 ( .A(n21779), .B(n21780), .Z(n21782) );
  AND U22150 ( .A(b[0]), .B(a[38]), .Z(n24272) );
  XNOR U22151 ( .A(n21780), .B(n21779), .Z(n24273) );
  NANDN U22152 ( .A(n24272), .B(n24273), .Z(n21781) );
  NAND U22153 ( .A(n21782), .B(n21781), .Z(n21784) );
  NANDN U22154 ( .A(n187), .B(b[0]), .Z(n21783) );
  NAND U22155 ( .A(n21784), .B(n21783), .Z(n21788) );
  XNOR U22156 ( .A(n21784), .B(n21783), .Z(n24275) );
  XOR U22157 ( .A(n21786), .B(n21785), .Z(n24274) );
  OR U22158 ( .A(n24275), .B(n24274), .Z(n21787) );
  NAND U22159 ( .A(n21788), .B(n21787), .Z(n21790) );
  NANDN U22160 ( .A(n21789), .B(n21790), .Z(n21792) );
  AND U22161 ( .A(b[0]), .B(a[40]), .Z(n24276) );
  XNOR U22162 ( .A(n21790), .B(n21789), .Z(n24277) );
  NANDN U22163 ( .A(n24276), .B(n24277), .Z(n21791) );
  NAND U22164 ( .A(n21792), .B(n21791), .Z(n21794) );
  NANDN U22165 ( .A(n189), .B(b[0]), .Z(n21793) );
  NAND U22166 ( .A(n21794), .B(n21793), .Z(n21798) );
  XNOR U22167 ( .A(n21794), .B(n21793), .Z(n24279) );
  XOR U22168 ( .A(n21796), .B(n21795), .Z(n24278) );
  OR U22169 ( .A(n24279), .B(n24278), .Z(n21797) );
  NAND U22170 ( .A(n21798), .B(n21797), .Z(n21800) );
  NANDN U22171 ( .A(n21799), .B(n21800), .Z(n21802) );
  AND U22172 ( .A(b[0]), .B(a[42]), .Z(n24282) );
  XNOR U22173 ( .A(n21800), .B(n21799), .Z(n24283) );
  NANDN U22174 ( .A(n24282), .B(n24283), .Z(n21801) );
  NAND U22175 ( .A(n21802), .B(n21801), .Z(n21804) );
  NANDN U22176 ( .A(n191), .B(b[0]), .Z(n21803) );
  NAND U22177 ( .A(n21804), .B(n21803), .Z(n21808) );
  XNOR U22178 ( .A(n21804), .B(n21803), .Z(n24285) );
  XOR U22179 ( .A(n21806), .B(n21805), .Z(n24284) );
  OR U22180 ( .A(n24285), .B(n24284), .Z(n21807) );
  NAND U22181 ( .A(n21808), .B(n21807), .Z(n21810) );
  NANDN U22182 ( .A(n21809), .B(n21810), .Z(n21812) );
  AND U22183 ( .A(b[0]), .B(a[44]), .Z(n24286) );
  XNOR U22184 ( .A(n21810), .B(n21809), .Z(n24287) );
  NANDN U22185 ( .A(n24286), .B(n24287), .Z(n21811) );
  NAND U22186 ( .A(n21812), .B(n21811), .Z(n21814) );
  NANDN U22187 ( .A(n193), .B(b[0]), .Z(n21813) );
  NAND U22188 ( .A(n21814), .B(n21813), .Z(n21818) );
  XNOR U22189 ( .A(n21814), .B(n21813), .Z(n24289) );
  XOR U22190 ( .A(n21816), .B(n21815), .Z(n24288) );
  OR U22191 ( .A(n24289), .B(n24288), .Z(n21817) );
  NAND U22192 ( .A(n21818), .B(n21817), .Z(n21820) );
  NANDN U22193 ( .A(n21819), .B(n21820), .Z(n21822) );
  AND U22194 ( .A(b[0]), .B(a[46]), .Z(n24290) );
  XNOR U22195 ( .A(n21820), .B(n21819), .Z(n24291) );
  NANDN U22196 ( .A(n24290), .B(n24291), .Z(n21821) );
  NAND U22197 ( .A(n21822), .B(n21821), .Z(n21824) );
  NANDN U22198 ( .A(n195), .B(b[0]), .Z(n21823) );
  NAND U22199 ( .A(n21824), .B(n21823), .Z(n21828) );
  XNOR U22200 ( .A(n21824), .B(n21823), .Z(n24293) );
  XOR U22201 ( .A(n21826), .B(n21825), .Z(n24292) );
  OR U22202 ( .A(n24293), .B(n24292), .Z(n21827) );
  NAND U22203 ( .A(n21828), .B(n21827), .Z(n21830) );
  NANDN U22204 ( .A(n21829), .B(n21830), .Z(n21832) );
  AND U22205 ( .A(b[0]), .B(a[48]), .Z(n24294) );
  XNOR U22206 ( .A(n21830), .B(n21829), .Z(n24295) );
  NANDN U22207 ( .A(n24294), .B(n24295), .Z(n21831) );
  NAND U22208 ( .A(n21832), .B(n21831), .Z(n21834) );
  NANDN U22209 ( .A(n197), .B(b[0]), .Z(n21833) );
  NAND U22210 ( .A(n21834), .B(n21833), .Z(n21838) );
  XNOR U22211 ( .A(n21834), .B(n21833), .Z(n24297) );
  XOR U22212 ( .A(n21836), .B(n21835), .Z(n24296) );
  OR U22213 ( .A(n24297), .B(n24296), .Z(n21837) );
  NAND U22214 ( .A(n21838), .B(n21837), .Z(n21840) );
  NANDN U22215 ( .A(n21839), .B(n21840), .Z(n21842) );
  AND U22216 ( .A(b[0]), .B(a[50]), .Z(n24298) );
  XNOR U22217 ( .A(n21840), .B(n21839), .Z(n24299) );
  NANDN U22218 ( .A(n24298), .B(n24299), .Z(n21841) );
  NAND U22219 ( .A(n21842), .B(n21841), .Z(n21844) );
  NANDN U22220 ( .A(n199), .B(b[0]), .Z(n21843) );
  NAND U22221 ( .A(n21844), .B(n21843), .Z(n21848) );
  XNOR U22222 ( .A(n21844), .B(n21843), .Z(n24301) );
  XOR U22223 ( .A(n21846), .B(n21845), .Z(n24300) );
  OR U22224 ( .A(n24301), .B(n24300), .Z(n21847) );
  NAND U22225 ( .A(n21848), .B(n21847), .Z(n21850) );
  NANDN U22226 ( .A(n21849), .B(n21850), .Z(n21852) );
  AND U22227 ( .A(b[0]), .B(a[52]), .Z(n24304) );
  XNOR U22228 ( .A(n21850), .B(n21849), .Z(n24305) );
  NANDN U22229 ( .A(n24304), .B(n24305), .Z(n21851) );
  NAND U22230 ( .A(n21852), .B(n21851), .Z(n21854) );
  NANDN U22231 ( .A(n201), .B(b[0]), .Z(n21853) );
  NAND U22232 ( .A(n21854), .B(n21853), .Z(n21858) );
  XNOR U22233 ( .A(n21854), .B(n21853), .Z(n24307) );
  XOR U22234 ( .A(n21856), .B(n21855), .Z(n24306) );
  OR U22235 ( .A(n24307), .B(n24306), .Z(n21857) );
  NAND U22236 ( .A(n21858), .B(n21857), .Z(n21860) );
  NANDN U22237 ( .A(n21859), .B(n21860), .Z(n21862) );
  AND U22238 ( .A(b[0]), .B(a[54]), .Z(n24308) );
  XNOR U22239 ( .A(n21860), .B(n21859), .Z(n24309) );
  NANDN U22240 ( .A(n24308), .B(n24309), .Z(n21861) );
  NAND U22241 ( .A(n21862), .B(n21861), .Z(n21864) );
  NANDN U22242 ( .A(n203), .B(b[0]), .Z(n21863) );
  NAND U22243 ( .A(n21864), .B(n21863), .Z(n21868) );
  XNOR U22244 ( .A(n21864), .B(n21863), .Z(n24311) );
  XOR U22245 ( .A(n21866), .B(n21865), .Z(n24310) );
  OR U22246 ( .A(n24311), .B(n24310), .Z(n21867) );
  NAND U22247 ( .A(n21868), .B(n21867), .Z(n21870) );
  NANDN U22248 ( .A(n21869), .B(n21870), .Z(n21872) );
  AND U22249 ( .A(b[0]), .B(a[56]), .Z(n24312) );
  XNOR U22250 ( .A(n21870), .B(n21869), .Z(n24313) );
  NANDN U22251 ( .A(n24312), .B(n24313), .Z(n21871) );
  NAND U22252 ( .A(n21872), .B(n21871), .Z(n21874) );
  NANDN U22253 ( .A(n205), .B(b[0]), .Z(n21873) );
  NAND U22254 ( .A(n21874), .B(n21873), .Z(n21878) );
  XNOR U22255 ( .A(n21874), .B(n21873), .Z(n24315) );
  XOR U22256 ( .A(n21876), .B(n21875), .Z(n24314) );
  OR U22257 ( .A(n24315), .B(n24314), .Z(n21877) );
  NAND U22258 ( .A(n21878), .B(n21877), .Z(n21880) );
  NANDN U22259 ( .A(n21879), .B(n21880), .Z(n21882) );
  AND U22260 ( .A(b[0]), .B(a[58]), .Z(n24316) );
  XNOR U22261 ( .A(n21880), .B(n21879), .Z(n24317) );
  NANDN U22262 ( .A(n24316), .B(n24317), .Z(n21881) );
  NAND U22263 ( .A(n21882), .B(n21881), .Z(n21884) );
  NANDN U22264 ( .A(n207), .B(b[0]), .Z(n21883) );
  NAND U22265 ( .A(n21884), .B(n21883), .Z(n21888) );
  XNOR U22266 ( .A(n21884), .B(n21883), .Z(n24319) );
  XOR U22267 ( .A(n21886), .B(n21885), .Z(n24318) );
  OR U22268 ( .A(n24319), .B(n24318), .Z(n21887) );
  NAND U22269 ( .A(n21888), .B(n21887), .Z(n21890) );
  NANDN U22270 ( .A(n21889), .B(n21890), .Z(n21892) );
  AND U22271 ( .A(b[0]), .B(a[60]), .Z(n24320) );
  XNOR U22272 ( .A(n21890), .B(n21889), .Z(n24321) );
  NANDN U22273 ( .A(n24320), .B(n24321), .Z(n21891) );
  NAND U22274 ( .A(n21892), .B(n21891), .Z(n21894) );
  NANDN U22275 ( .A(n209), .B(b[0]), .Z(n21893) );
  NAND U22276 ( .A(n21894), .B(n21893), .Z(n21898) );
  XNOR U22277 ( .A(n21894), .B(n21893), .Z(n24323) );
  XOR U22278 ( .A(n21896), .B(n21895), .Z(n24322) );
  OR U22279 ( .A(n24323), .B(n24322), .Z(n21897) );
  NAND U22280 ( .A(n21898), .B(n21897), .Z(n21902) );
  XOR U22281 ( .A(n21900), .B(n21899), .Z(n21901) );
  NAND U22282 ( .A(n21902), .B(n21901), .Z(n21904) );
  AND U22283 ( .A(b[0]), .B(a[62]), .Z(n24326) );
  XNOR U22284 ( .A(n21902), .B(n21901), .Z(n24327) );
  OR U22285 ( .A(n24326), .B(n24327), .Z(n21903) );
  NAND U22286 ( .A(n21904), .B(n21903), .Z(n21906) );
  NANDN U22287 ( .A(n210), .B(b[0]), .Z(n21905) );
  NAND U22288 ( .A(n21906), .B(n21905), .Z(n21910) );
  XNOR U22289 ( .A(n21906), .B(n21905), .Z(n24329) );
  XOR U22290 ( .A(n21908), .B(n21907), .Z(n24328) );
  OR U22291 ( .A(n24329), .B(n24328), .Z(n21909) );
  NAND U22292 ( .A(n21910), .B(n21909), .Z(n24331) );
  XNOR U22293 ( .A(n21912), .B(n21911), .Z(n24330) );
  OR U22294 ( .A(n24331), .B(n24330), .Z(n24089) );
  XNOR U22295 ( .A(n21914), .B(n21913), .Z(n24088) );
  OR U22296 ( .A(n24089), .B(n24088), .Z(n21915) );
  AND U22297 ( .A(n21916), .B(n21915), .Z(n24090) );
  NOR U22298 ( .A(n24091), .B(n24090), .Z(n24097) );
  IV U22299 ( .A(n24097), .Z(n24094) );
  NANDN U22300 ( .A(n24100), .B(n24094), .Z(n21919) );
  IV U22301 ( .A(n21917), .Z(n24093) );
  ANDN U22302 ( .B(n24093), .A(n24092), .Z(n21918) );
  ANDN U22303 ( .B(n21919), .A(n21918), .Z(n21920) );
  NANDN U22304 ( .A(n21921), .B(n21920), .Z(n21922) );
  NAND U22305 ( .A(n21923), .B(n21922), .Z(n21925) );
  ANDN U22306 ( .B(n24106), .A(n24105), .Z(n21924) );
  ANDN U22307 ( .B(n21925), .A(n21924), .Z(n24109) );
  XNOR U22308 ( .A(n21927), .B(n21926), .Z(n24110) );
  NANDN U22309 ( .A(n24109), .B(n24110), .Z(n21928) );
  NAND U22310 ( .A(n21929), .B(n21928), .Z(n24111) );
  OR U22311 ( .A(n24112), .B(n24111), .Z(n21930) );
  NAND U22312 ( .A(n21931), .B(n21930), .Z(n24114) );
  XNOR U22313 ( .A(n21933), .B(n21932), .Z(n24113) );
  NANDN U22314 ( .A(n24114), .B(n24113), .Z(n21934) );
  AND U22315 ( .A(n21935), .B(n21934), .Z(n24115) );
  OR U22316 ( .A(n24116), .B(n24115), .Z(n21936) );
  AND U22317 ( .A(n21937), .B(n21936), .Z(n24120) );
  NANDN U22318 ( .A(n21938), .B(n24120), .Z(n21949) );
  ANDN U22319 ( .B(n24138), .A(n24139), .Z(n21940) );
  NOR U22320 ( .A(n21939), .B(n24132), .Z(n24137) );
  NOR U22321 ( .A(n21940), .B(n24137), .Z(n21947) );
  AND U22322 ( .A(n21942), .B(n21941), .Z(n21945) );
  NOR U22323 ( .A(n24117), .B(n24119), .Z(n24121) );
  NANDN U22324 ( .A(n24121), .B(n24123), .Z(n21943) );
  ANDN U22325 ( .B(n21943), .A(n24132), .Z(n21944) );
  NANDN U22326 ( .A(n21945), .B(n21944), .Z(n21946) );
  AND U22327 ( .A(n21947), .B(n21946), .Z(n21948) );
  NAND U22328 ( .A(n21949), .B(n21948), .Z(n21950) );
  NANDN U22329 ( .A(n21951), .B(n21950), .Z(n21955) );
  OR U22330 ( .A(n21953), .B(n21952), .Z(n21954) );
  AND U22331 ( .A(n21955), .B(n21954), .Z(n24142) );
  XNOR U22332 ( .A(n21957), .B(n21956), .Z(n24143) );
  NANDN U22333 ( .A(n24142), .B(n24143), .Z(n24145) );
  OR U22334 ( .A(n24144), .B(n24145), .Z(n21958) );
  AND U22335 ( .A(n21959), .B(n21958), .Z(n24146) );
  XNOR U22336 ( .A(n21961), .B(n21960), .Z(n24147) );
  XOR U22337 ( .A(n21963), .B(n21962), .Z(n24148) );
  NANDN U22338 ( .A(n24149), .B(n24148), .Z(n21964) );
  AND U22339 ( .A(n21965), .B(n21964), .Z(n24153) );
  NAND U22340 ( .A(n24166), .B(n24167), .Z(n21966) );
  AND U22341 ( .A(n21967), .B(n21966), .Z(n24168) );
  XOR U22342 ( .A(n21969), .B(n21968), .Z(n24169) );
  XOR U22343 ( .A(n21971), .B(n21970), .Z(n24171) );
  OR U22344 ( .A(n24173), .B(n24172), .Z(n21972) );
  AND U22345 ( .A(n21973), .B(n21972), .Z(n24176) );
  IV U22346 ( .A(n21974), .Z(n24180) );
  NOR U22347 ( .A(n21976), .B(n24175), .Z(n24179) );
  XNOR U22348 ( .A(n21979), .B(n21978), .Z(n24193) );
  AND U22349 ( .A(n21981), .B(n21980), .Z(n24192) );
  XNOR U22350 ( .A(n21983), .B(n21982), .Z(n24197) );
  NANDN U22351 ( .A(n24196), .B(n24197), .Z(n21984) );
  NAND U22352 ( .A(n21985), .B(n21984), .Z(n24199) );
  OR U22353 ( .A(n24198), .B(n24199), .Z(n21986) );
  NAND U22354 ( .A(n21987), .B(n21986), .Z(n24200) );
  XNOR U22355 ( .A(n21989), .B(n21988), .Z(n24201) );
  NANDN U22356 ( .A(n24200), .B(n24201), .Z(n21990) );
  AND U22357 ( .A(n21991), .B(n21990), .Z(n24202) );
  XOR U22358 ( .A(n21993), .B(n21992), .Z(n24203) );
  XOR U22359 ( .A(n21995), .B(n21994), .Z(n24205) );
  NANDN U22360 ( .A(n24204), .B(n24205), .Z(n21996) );
  NAND U22361 ( .A(n21997), .B(n21996), .Z(n24207) );
  XOR U22362 ( .A(n21999), .B(n21998), .Z(n24206) );
  OR U22363 ( .A(n24209), .B(n24208), .Z(n22000) );
  NAND U22364 ( .A(n22001), .B(n22000), .Z(n24213) );
  NANDN U22365 ( .A(n22002), .B(n24213), .Z(n22003) );
  NAND U22366 ( .A(n22004), .B(n22003), .Z(n22297) );
  OR U22367 ( .A(n22006), .B(n22005), .Z(n22295) );
  AND U22368 ( .A(a[61]), .B(b[41]), .Z(n22282) );
  OR U22369 ( .A(n22008), .B(n22007), .Z(n22012) );
  NANDN U22370 ( .A(n22010), .B(n22009), .Z(n22011) );
  NAND U22371 ( .A(n22012), .B(n22011), .Z(n22268) );
  OR U22372 ( .A(n22014), .B(n22013), .Z(n22018) );
  NANDN U22373 ( .A(n22016), .B(n22015), .Z(n22017) );
  NAND U22374 ( .A(n22018), .B(n22017), .Z(n22256) );
  AND U22375 ( .A(a[55]), .B(b[47]), .Z(n22248) );
  OR U22376 ( .A(n22020), .B(n22019), .Z(n22024) );
  NANDN U22377 ( .A(n22022), .B(n22021), .Z(n22023) );
  NAND U22378 ( .A(n22024), .B(n22023), .Z(n22234) );
  OR U22379 ( .A(n22026), .B(n22025), .Z(n22030) );
  NANDN U22380 ( .A(n22028), .B(n22027), .Z(n22029) );
  NAND U22381 ( .A(n22030), .B(n22029), .Z(n22222) );
  AND U22382 ( .A(a[49]), .B(b[53]), .Z(n22214) );
  OR U22383 ( .A(n22032), .B(n22031), .Z(n22036) );
  NANDN U22384 ( .A(n22034), .B(n22033), .Z(n22035) );
  NAND U22385 ( .A(n22036), .B(n22035), .Z(n22200) );
  AND U22386 ( .A(a[45]), .B(b[57]), .Z(n22192) );
  OR U22387 ( .A(n22038), .B(n22037), .Z(n22042) );
  NANDN U22388 ( .A(n22040), .B(n22039), .Z(n22041) );
  NAND U22389 ( .A(n22042), .B(n22041), .Z(n22178) );
  AND U22390 ( .A(a[41]), .B(b[61]), .Z(n22168) );
  OR U22391 ( .A(n22044), .B(n22043), .Z(n22048) );
  OR U22392 ( .A(n22046), .B(n22045), .Z(n22047) );
  NAND U22393 ( .A(n22048), .B(n22047), .Z(n22160) );
  NAND U22394 ( .A(a[40]), .B(b[62]), .Z(n22159) );
  XOR U22395 ( .A(n22160), .B(n22159), .Z(n22161) );
  NAND U22396 ( .A(a[39]), .B(b[63]), .Z(n22162) );
  XOR U22397 ( .A(n22161), .B(n22162), .Z(n22165) );
  OR U22398 ( .A(n22050), .B(n22049), .Z(n22054) );
  OR U22399 ( .A(n22052), .B(n22051), .Z(n22053) );
  AND U22400 ( .A(n22054), .B(n22053), .Z(n22166) );
  XNOR U22401 ( .A(n22165), .B(n22166), .Z(n22167) );
  XOR U22402 ( .A(n22168), .B(n22167), .Z(n22174) );
  OR U22403 ( .A(n22056), .B(n22055), .Z(n22060) );
  OR U22404 ( .A(n22058), .B(n22057), .Z(n22059) );
  NAND U22405 ( .A(n22060), .B(n22059), .Z(n22172) );
  NAND U22406 ( .A(b[60]), .B(a[42]), .Z(n22171) );
  XOR U22407 ( .A(n22172), .B(n22171), .Z(n22173) );
  XOR U22408 ( .A(n22174), .B(n22173), .Z(n22177) );
  XNOR U22409 ( .A(n22178), .B(n22177), .Z(n22180) );
  NAND U22410 ( .A(b[59]), .B(a[43]), .Z(n22179) );
  XOR U22411 ( .A(n22180), .B(n22179), .Z(n22185) );
  OR U22412 ( .A(n22062), .B(n22061), .Z(n22066) );
  NANDN U22413 ( .A(n22064), .B(n22063), .Z(n22065) );
  NAND U22414 ( .A(n22066), .B(n22065), .Z(n22184) );
  NAND U22415 ( .A(b[58]), .B(a[44]), .Z(n22183) );
  XOR U22416 ( .A(n22184), .B(n22183), .Z(n22186) );
  XOR U22417 ( .A(n22185), .B(n22186), .Z(n22189) );
  OR U22418 ( .A(n22068), .B(n22067), .Z(n22072) );
  NANDN U22419 ( .A(n22070), .B(n22069), .Z(n22071) );
  NAND U22420 ( .A(n22072), .B(n22071), .Z(n22190) );
  XOR U22421 ( .A(n22189), .B(n22190), .Z(n22191) );
  XOR U22422 ( .A(n22192), .B(n22191), .Z(n22196) );
  OR U22423 ( .A(n22074), .B(n22073), .Z(n22078) );
  NANDN U22424 ( .A(n22076), .B(n22075), .Z(n22077) );
  NAND U22425 ( .A(n22078), .B(n22077), .Z(n22193) );
  NAND U22426 ( .A(a[46]), .B(b[56]), .Z(n22194) );
  XNOR U22427 ( .A(n22193), .B(n22194), .Z(n22195) );
  XOR U22428 ( .A(n22196), .B(n22195), .Z(n22199) );
  XOR U22429 ( .A(n22200), .B(n22199), .Z(n22202) );
  NAND U22430 ( .A(b[55]), .B(a[47]), .Z(n22201) );
  XOR U22431 ( .A(n22202), .B(n22201), .Z(n22207) );
  OR U22432 ( .A(n22080), .B(n22079), .Z(n22084) );
  OR U22433 ( .A(n22082), .B(n22081), .Z(n22083) );
  NAND U22434 ( .A(n22084), .B(n22083), .Z(n22206) );
  NAND U22435 ( .A(b[54]), .B(a[48]), .Z(n22205) );
  XOR U22436 ( .A(n22206), .B(n22205), .Z(n22208) );
  XOR U22437 ( .A(n22207), .B(n22208), .Z(n22211) );
  OR U22438 ( .A(n22086), .B(n22085), .Z(n22090) );
  NANDN U22439 ( .A(n22088), .B(n22087), .Z(n22089) );
  NAND U22440 ( .A(n22090), .B(n22089), .Z(n22212) );
  XOR U22441 ( .A(n22211), .B(n22212), .Z(n22213) );
  XOR U22442 ( .A(n22214), .B(n22213), .Z(n22218) );
  OR U22443 ( .A(n22092), .B(n22091), .Z(n22096) );
  NANDN U22444 ( .A(n22094), .B(n22093), .Z(n22095) );
  NAND U22445 ( .A(n22096), .B(n22095), .Z(n22215) );
  NAND U22446 ( .A(a[50]), .B(b[52]), .Z(n22216) );
  XNOR U22447 ( .A(n22215), .B(n22216), .Z(n22217) );
  XOR U22448 ( .A(n22218), .B(n22217), .Z(n22221) );
  XOR U22449 ( .A(n22222), .B(n22221), .Z(n22224) );
  NAND U22450 ( .A(b[51]), .B(a[51]), .Z(n22223) );
  XOR U22451 ( .A(n22224), .B(n22223), .Z(n22229) );
  OR U22452 ( .A(n22098), .B(n22097), .Z(n22102) );
  OR U22453 ( .A(n22100), .B(n22099), .Z(n22101) );
  NAND U22454 ( .A(n22102), .B(n22101), .Z(n22228) );
  NAND U22455 ( .A(b[50]), .B(a[52]), .Z(n22227) );
  XOR U22456 ( .A(n22228), .B(n22227), .Z(n22230) );
  XOR U22457 ( .A(n22229), .B(n22230), .Z(n22233) );
  XNOR U22458 ( .A(n22234), .B(n22233), .Z(n22236) );
  NAND U22459 ( .A(b[49]), .B(a[53]), .Z(n22235) );
  XOR U22460 ( .A(n22236), .B(n22235), .Z(n22241) );
  OR U22461 ( .A(n22104), .B(n22103), .Z(n22108) );
  OR U22462 ( .A(n22106), .B(n22105), .Z(n22107) );
  NAND U22463 ( .A(n22108), .B(n22107), .Z(n22240) );
  NAND U22464 ( .A(b[48]), .B(a[54]), .Z(n22239) );
  XOR U22465 ( .A(n22240), .B(n22239), .Z(n22242) );
  XOR U22466 ( .A(n22241), .B(n22242), .Z(n22245) );
  NANDN U22467 ( .A(n22110), .B(n22109), .Z(n22114) );
  NANDN U22468 ( .A(n22112), .B(n22111), .Z(n22113) );
  AND U22469 ( .A(n22114), .B(n22113), .Z(n22246) );
  XOR U22470 ( .A(n22245), .B(n22246), .Z(n22247) );
  XOR U22471 ( .A(n22248), .B(n22247), .Z(n22252) );
  OR U22472 ( .A(n22116), .B(n22115), .Z(n22120) );
  OR U22473 ( .A(n22118), .B(n22117), .Z(n22119) );
  NAND U22474 ( .A(n22120), .B(n22119), .Z(n22250) );
  NAND U22475 ( .A(b[46]), .B(a[56]), .Z(n22249) );
  XOR U22476 ( .A(n22250), .B(n22249), .Z(n22251) );
  XOR U22477 ( .A(n22252), .B(n22251), .Z(n22255) );
  XNOR U22478 ( .A(n22256), .B(n22255), .Z(n22258) );
  NAND U22479 ( .A(b[45]), .B(a[57]), .Z(n22257) );
  XOR U22480 ( .A(n22258), .B(n22257), .Z(n22263) );
  OR U22481 ( .A(n22122), .B(n22121), .Z(n22126) );
  OR U22482 ( .A(n22124), .B(n22123), .Z(n22125) );
  NAND U22483 ( .A(n22126), .B(n22125), .Z(n22261) );
  NAND U22484 ( .A(a[58]), .B(b[44]), .Z(n22262) );
  XNOR U22485 ( .A(n22261), .B(n22262), .Z(n22264) );
  XOR U22486 ( .A(n22263), .B(n22264), .Z(n22267) );
  XOR U22487 ( .A(n22268), .B(n22267), .Z(n22270) );
  NAND U22488 ( .A(b[43]), .B(a[59]), .Z(n22269) );
  XOR U22489 ( .A(n22270), .B(n22269), .Z(n22275) );
  OR U22490 ( .A(n22128), .B(n22127), .Z(n22132) );
  OR U22491 ( .A(n22130), .B(n22129), .Z(n22131) );
  NAND U22492 ( .A(n22132), .B(n22131), .Z(n22274) );
  NAND U22493 ( .A(b[42]), .B(a[60]), .Z(n22273) );
  XOR U22494 ( .A(n22274), .B(n22273), .Z(n22276) );
  XOR U22495 ( .A(n22275), .B(n22276), .Z(n22279) );
  OR U22496 ( .A(n22134), .B(n22133), .Z(n22138) );
  NANDN U22497 ( .A(n22136), .B(n22135), .Z(n22137) );
  NAND U22498 ( .A(n22138), .B(n22137), .Z(n22280) );
  XOR U22499 ( .A(n22279), .B(n22280), .Z(n22281) );
  XOR U22500 ( .A(n22282), .B(n22281), .Z(n22286) );
  OR U22501 ( .A(n22140), .B(n22139), .Z(n22144) );
  NANDN U22502 ( .A(n22142), .B(n22141), .Z(n22143) );
  NAND U22503 ( .A(n22144), .B(n22143), .Z(n22283) );
  NAND U22504 ( .A(a[62]), .B(b[40]), .Z(n22284) );
  XNOR U22505 ( .A(n22283), .B(n22284), .Z(n22285) );
  XOR U22506 ( .A(n22286), .B(n22285), .Z(n22289) );
  OR U22507 ( .A(n22146), .B(n22145), .Z(n22150) );
  NANDN U22508 ( .A(n22148), .B(n22147), .Z(n22149) );
  AND U22509 ( .A(n22150), .B(n22149), .Z(n22290) );
  XNOR U22510 ( .A(n22289), .B(n22290), .Z(n22292) );
  NAND U22511 ( .A(b[39]), .B(a[63]), .Z(n22291) );
  XNOR U22512 ( .A(n22292), .B(n22291), .Z(n22158) );
  OR U22513 ( .A(n22152), .B(n22151), .Z(n22156) );
  OR U22514 ( .A(n22154), .B(n22153), .Z(n22155) );
  NAND U22515 ( .A(n22156), .B(n22155), .Z(n22157) );
  XOR U22516 ( .A(n22158), .B(n22157), .Z(n22296) );
  XNOR U22517 ( .A(n22295), .B(n22296), .Z(n22298) );
  XNOR U22518 ( .A(n22297), .B(n22298), .Z(c[102]) );
  NOR U22519 ( .A(n22158), .B(n22157), .Z(n22441) );
  AND U22520 ( .A(b[63]), .B(a[40]), .Z(n22402) );
  AND U22521 ( .A(b[62]), .B(a[41]), .Z(n22399) );
  OR U22522 ( .A(n22160), .B(n22159), .Z(n22164) );
  NANDN U22523 ( .A(n22162), .B(n22161), .Z(n22163) );
  NAND U22524 ( .A(n22164), .B(n22163), .Z(n22400) );
  XOR U22525 ( .A(n22399), .B(n22400), .Z(n22401) );
  XOR U22526 ( .A(n22402), .B(n22401), .Z(n22396) );
  NANDN U22527 ( .A(n22166), .B(n22165), .Z(n22170) );
  NANDN U22528 ( .A(n22168), .B(n22167), .Z(n22169) );
  NAND U22529 ( .A(n22170), .B(n22169), .Z(n22394) );
  NAND U22530 ( .A(b[61]), .B(a[42]), .Z(n22393) );
  XOR U22531 ( .A(n22394), .B(n22393), .Z(n22395) );
  XOR U22532 ( .A(n22396), .B(n22395), .Z(n22408) );
  AND U22533 ( .A(a[43]), .B(b[60]), .Z(n22405) );
  OR U22534 ( .A(n22172), .B(n22171), .Z(n22176) );
  NAND U22535 ( .A(n22174), .B(n22173), .Z(n22175) );
  NAND U22536 ( .A(n22176), .B(n22175), .Z(n22406) );
  XOR U22537 ( .A(n22405), .B(n22406), .Z(n22407) );
  XNOR U22538 ( .A(n22408), .B(n22407), .Z(n22390) );
  NAND U22539 ( .A(n22178), .B(n22177), .Z(n22182) );
  OR U22540 ( .A(n22180), .B(n22179), .Z(n22181) );
  NAND U22541 ( .A(n22182), .B(n22181), .Z(n22387) );
  NAND U22542 ( .A(a[44]), .B(b[59]), .Z(n22388) );
  XNOR U22543 ( .A(n22387), .B(n22388), .Z(n22389) );
  XNOR U22544 ( .A(n22390), .B(n22389), .Z(n22384) );
  AND U22545 ( .A(a[45]), .B(b[58]), .Z(n22381) );
  OR U22546 ( .A(n22184), .B(n22183), .Z(n22188) );
  NAND U22547 ( .A(n22186), .B(n22185), .Z(n22187) );
  NAND U22548 ( .A(n22188), .B(n22187), .Z(n22382) );
  XOR U22549 ( .A(n22381), .B(n22382), .Z(n22383) );
  XNOR U22550 ( .A(n22384), .B(n22383), .Z(n22414) );
  NAND U22551 ( .A(b[57]), .B(a[46]), .Z(n22411) );
  XOR U22552 ( .A(n22412), .B(n22411), .Z(n22413) );
  XNOR U22553 ( .A(n22414), .B(n22413), .Z(n22420) );
  AND U22554 ( .A(a[47]), .B(b[56]), .Z(n22417) );
  NANDN U22555 ( .A(n22194), .B(n22193), .Z(n22198) );
  NAND U22556 ( .A(n22196), .B(n22195), .Z(n22197) );
  NAND U22557 ( .A(n22198), .B(n22197), .Z(n22418) );
  XOR U22558 ( .A(n22417), .B(n22418), .Z(n22419) );
  XNOR U22559 ( .A(n22420), .B(n22419), .Z(n22378) );
  NANDN U22560 ( .A(n22200), .B(n22199), .Z(n22204) );
  OR U22561 ( .A(n22202), .B(n22201), .Z(n22203) );
  NAND U22562 ( .A(n22204), .B(n22203), .Z(n22375) );
  NAND U22563 ( .A(a[48]), .B(b[55]), .Z(n22376) );
  XNOR U22564 ( .A(n22375), .B(n22376), .Z(n22377) );
  XNOR U22565 ( .A(n22378), .B(n22377), .Z(n22372) );
  AND U22566 ( .A(a[49]), .B(b[54]), .Z(n22369) );
  OR U22567 ( .A(n22206), .B(n22205), .Z(n22210) );
  NAND U22568 ( .A(n22208), .B(n22207), .Z(n22209) );
  NAND U22569 ( .A(n22210), .B(n22209), .Z(n22370) );
  XOR U22570 ( .A(n22369), .B(n22370), .Z(n22371) );
  XNOR U22571 ( .A(n22372), .B(n22371), .Z(n22366) );
  NAND U22572 ( .A(b[53]), .B(a[50]), .Z(n22363) );
  XOR U22573 ( .A(n22364), .B(n22363), .Z(n22365) );
  XNOR U22574 ( .A(n22366), .B(n22365), .Z(n22360) );
  AND U22575 ( .A(a[51]), .B(b[52]), .Z(n22357) );
  NANDN U22576 ( .A(n22216), .B(n22215), .Z(n22220) );
  NAND U22577 ( .A(n22218), .B(n22217), .Z(n22219) );
  NAND U22578 ( .A(n22220), .B(n22219), .Z(n22358) );
  XOR U22579 ( .A(n22357), .B(n22358), .Z(n22359) );
  XNOR U22580 ( .A(n22360), .B(n22359), .Z(n22354) );
  NANDN U22581 ( .A(n22222), .B(n22221), .Z(n22226) );
  OR U22582 ( .A(n22224), .B(n22223), .Z(n22225) );
  NAND U22583 ( .A(n22226), .B(n22225), .Z(n22351) );
  NAND U22584 ( .A(a[52]), .B(b[51]), .Z(n22352) );
  XNOR U22585 ( .A(n22351), .B(n22352), .Z(n22353) );
  XNOR U22586 ( .A(n22354), .B(n22353), .Z(n22348) );
  AND U22587 ( .A(a[53]), .B(b[50]), .Z(n22345) );
  OR U22588 ( .A(n22228), .B(n22227), .Z(n22232) );
  NAND U22589 ( .A(n22230), .B(n22229), .Z(n22231) );
  NAND U22590 ( .A(n22232), .B(n22231), .Z(n22346) );
  XOR U22591 ( .A(n22345), .B(n22346), .Z(n22347) );
  XNOR U22592 ( .A(n22348), .B(n22347), .Z(n22342) );
  NAND U22593 ( .A(n22234), .B(n22233), .Z(n22238) );
  OR U22594 ( .A(n22236), .B(n22235), .Z(n22237) );
  NAND U22595 ( .A(n22238), .B(n22237), .Z(n22339) );
  NAND U22596 ( .A(a[54]), .B(b[49]), .Z(n22340) );
  XNOR U22597 ( .A(n22339), .B(n22340), .Z(n22341) );
  XNOR U22598 ( .A(n22342), .B(n22341), .Z(n22336) );
  AND U22599 ( .A(a[55]), .B(b[48]), .Z(n22333) );
  OR U22600 ( .A(n22240), .B(n22239), .Z(n22244) );
  NAND U22601 ( .A(n22242), .B(n22241), .Z(n22243) );
  NAND U22602 ( .A(n22244), .B(n22243), .Z(n22334) );
  XOR U22603 ( .A(n22333), .B(n22334), .Z(n22335) );
  XNOR U22604 ( .A(n22336), .B(n22335), .Z(n22330) );
  NAND U22605 ( .A(b[47]), .B(a[56]), .Z(n22327) );
  XOR U22606 ( .A(n22328), .B(n22327), .Z(n22329) );
  XNOR U22607 ( .A(n22330), .B(n22329), .Z(n22426) );
  AND U22608 ( .A(a[57]), .B(b[46]), .Z(n22423) );
  OR U22609 ( .A(n22250), .B(n22249), .Z(n22254) );
  NAND U22610 ( .A(n22252), .B(n22251), .Z(n22253) );
  NAND U22611 ( .A(n22254), .B(n22253), .Z(n22424) );
  XOR U22612 ( .A(n22423), .B(n22424), .Z(n22425) );
  XNOR U22613 ( .A(n22426), .B(n22425), .Z(n22324) );
  NAND U22614 ( .A(n22256), .B(n22255), .Z(n22260) );
  OR U22615 ( .A(n22258), .B(n22257), .Z(n22259) );
  NAND U22616 ( .A(n22260), .B(n22259), .Z(n22321) );
  NAND U22617 ( .A(a[58]), .B(b[45]), .Z(n22322) );
  XNOR U22618 ( .A(n22321), .B(n22322), .Z(n22323) );
  XNOR U22619 ( .A(n22324), .B(n22323), .Z(n22318) );
  AND U22620 ( .A(a[59]), .B(b[44]), .Z(n22315) );
  NANDN U22621 ( .A(n22262), .B(n22261), .Z(n22266) );
  NAND U22622 ( .A(n22264), .B(n22263), .Z(n22265) );
  NAND U22623 ( .A(n22266), .B(n22265), .Z(n22316) );
  XOR U22624 ( .A(n22315), .B(n22316), .Z(n22317) );
  XNOR U22625 ( .A(n22318), .B(n22317), .Z(n22312) );
  NANDN U22626 ( .A(n22268), .B(n22267), .Z(n22272) );
  OR U22627 ( .A(n22270), .B(n22269), .Z(n22271) );
  NAND U22628 ( .A(n22272), .B(n22271), .Z(n22309) );
  NAND U22629 ( .A(a[60]), .B(b[43]), .Z(n22310) );
  XNOR U22630 ( .A(n22309), .B(n22310), .Z(n22311) );
  XNOR U22631 ( .A(n22312), .B(n22311), .Z(n22306) );
  AND U22632 ( .A(a[61]), .B(b[42]), .Z(n22303) );
  OR U22633 ( .A(n22274), .B(n22273), .Z(n22278) );
  NAND U22634 ( .A(n22276), .B(n22275), .Z(n22277) );
  NAND U22635 ( .A(n22278), .B(n22277), .Z(n22304) );
  XOR U22636 ( .A(n22303), .B(n22304), .Z(n22305) );
  XNOR U22637 ( .A(n22306), .B(n22305), .Z(n22432) );
  NAND U22638 ( .A(b[41]), .B(a[62]), .Z(n22429) );
  XOR U22639 ( .A(n22430), .B(n22429), .Z(n22431) );
  XNOR U22640 ( .A(n22432), .B(n22431), .Z(n22438) );
  AND U22641 ( .A(a[63]), .B(b[40]), .Z(n22435) );
  NANDN U22642 ( .A(n22284), .B(n22283), .Z(n22288) );
  NAND U22643 ( .A(n22286), .B(n22285), .Z(n22287) );
  NAND U22644 ( .A(n22288), .B(n22287), .Z(n22436) );
  XOR U22645 ( .A(n22435), .B(n22436), .Z(n22437) );
  XNOR U22646 ( .A(n22438), .B(n22437), .Z(n22301) );
  NAND U22647 ( .A(n22290), .B(n22289), .Z(n22294) );
  OR U22648 ( .A(n22292), .B(n22291), .Z(n22293) );
  NAND U22649 ( .A(n22294), .B(n22293), .Z(n22302) );
  XNOR U22650 ( .A(n22301), .B(n22302), .Z(n22442) );
  XOR U22651 ( .A(n22441), .B(n22442), .Z(n22443) );
  NANDN U22652 ( .A(n22296), .B(n22295), .Z(n22300) );
  NAND U22653 ( .A(n22298), .B(n22297), .Z(n22299) );
  AND U22654 ( .A(n22300), .B(n22299), .Z(n22444) );
  XOR U22655 ( .A(n22443), .B(n22444), .Z(c[103]) );
  ANDN U22656 ( .B(n22302), .A(n22301), .Z(n22577) );
  NAND U22657 ( .A(a[63]), .B(b[41]), .Z(n22574) );
  OR U22658 ( .A(n22304), .B(n22303), .Z(n22308) );
  NANDN U22659 ( .A(n22306), .B(n22305), .Z(n22307) );
  NAND U22660 ( .A(n22308), .B(n22307), .Z(n22566) );
  NAND U22661 ( .A(b[42]), .B(a[62]), .Z(n22565) );
  XOR U22662 ( .A(n22566), .B(n22565), .Z(n22567) );
  NANDN U22663 ( .A(n22310), .B(n22309), .Z(n22314) );
  NANDN U22664 ( .A(n22312), .B(n22311), .Z(n22313) );
  NAND U22665 ( .A(n22314), .B(n22313), .Z(n22560) );
  OR U22666 ( .A(n22316), .B(n22315), .Z(n22320) );
  NANDN U22667 ( .A(n22318), .B(n22317), .Z(n22319) );
  NAND U22668 ( .A(n22320), .B(n22319), .Z(n22554) );
  NAND U22669 ( .A(b[44]), .B(a[60]), .Z(n22553) );
  XOR U22670 ( .A(n22554), .B(n22553), .Z(n22555) );
  NANDN U22671 ( .A(n22322), .B(n22321), .Z(n22326) );
  NANDN U22672 ( .A(n22324), .B(n22323), .Z(n22325) );
  NAND U22673 ( .A(n22326), .B(n22325), .Z(n22548) );
  OR U22674 ( .A(n22328), .B(n22327), .Z(n22332) );
  NANDN U22675 ( .A(n22330), .B(n22329), .Z(n22331) );
  NAND U22676 ( .A(n22332), .B(n22331), .Z(n22536) );
  OR U22677 ( .A(n22334), .B(n22333), .Z(n22338) );
  NANDN U22678 ( .A(n22336), .B(n22335), .Z(n22337) );
  NAND U22679 ( .A(n22338), .B(n22337), .Z(n22530) );
  NAND U22680 ( .A(b[48]), .B(a[56]), .Z(n22529) );
  XOR U22681 ( .A(n22530), .B(n22529), .Z(n22531) );
  NANDN U22682 ( .A(n22340), .B(n22339), .Z(n22344) );
  NANDN U22683 ( .A(n22342), .B(n22341), .Z(n22343) );
  NAND U22684 ( .A(n22344), .B(n22343), .Z(n22524) );
  OR U22685 ( .A(n22346), .B(n22345), .Z(n22350) );
  NANDN U22686 ( .A(n22348), .B(n22347), .Z(n22349) );
  NAND U22687 ( .A(n22350), .B(n22349), .Z(n22518) );
  NAND U22688 ( .A(b[50]), .B(a[54]), .Z(n22517) );
  XOR U22689 ( .A(n22518), .B(n22517), .Z(n22519) );
  NANDN U22690 ( .A(n22352), .B(n22351), .Z(n22356) );
  NANDN U22691 ( .A(n22354), .B(n22353), .Z(n22355) );
  NAND U22692 ( .A(n22356), .B(n22355), .Z(n22512) );
  OR U22693 ( .A(n22358), .B(n22357), .Z(n22362) );
  NANDN U22694 ( .A(n22360), .B(n22359), .Z(n22361) );
  NAND U22695 ( .A(n22362), .B(n22361), .Z(n22506) );
  NAND U22696 ( .A(b[52]), .B(a[52]), .Z(n22505) );
  XOR U22697 ( .A(n22506), .B(n22505), .Z(n22507) );
  OR U22698 ( .A(n22364), .B(n22363), .Z(n22368) );
  NANDN U22699 ( .A(n22366), .B(n22365), .Z(n22367) );
  NAND U22700 ( .A(n22368), .B(n22367), .Z(n22500) );
  OR U22701 ( .A(n22370), .B(n22369), .Z(n22374) );
  NANDN U22702 ( .A(n22372), .B(n22371), .Z(n22373) );
  NAND U22703 ( .A(n22374), .B(n22373), .Z(n22494) );
  NAND U22704 ( .A(b[54]), .B(a[50]), .Z(n22493) );
  XOR U22705 ( .A(n22494), .B(n22493), .Z(n22495) );
  NANDN U22706 ( .A(n22376), .B(n22375), .Z(n22380) );
  NANDN U22707 ( .A(n22378), .B(n22377), .Z(n22379) );
  NAND U22708 ( .A(n22380), .B(n22379), .Z(n22488) );
  OR U22709 ( .A(n22382), .B(n22381), .Z(n22386) );
  NANDN U22710 ( .A(n22384), .B(n22383), .Z(n22385) );
  NAND U22711 ( .A(n22386), .B(n22385), .Z(n22472) );
  NAND U22712 ( .A(b[58]), .B(a[46]), .Z(n22471) );
  XOR U22713 ( .A(n22472), .B(n22471), .Z(n22473) );
  NANDN U22714 ( .A(n22388), .B(n22387), .Z(n22392) );
  NANDN U22715 ( .A(n22390), .B(n22389), .Z(n22391) );
  NAND U22716 ( .A(n22392), .B(n22391), .Z(n22466) );
  OR U22717 ( .A(n22394), .B(n22393), .Z(n22398) );
  NAND U22718 ( .A(n22396), .B(n22395), .Z(n22397) );
  NAND U22719 ( .A(n22398), .B(n22397), .Z(n22453) );
  NAND U22720 ( .A(a[43]), .B(b[61]), .Z(n22454) );
  XNOR U22721 ( .A(n22453), .B(n22454), .Z(n22455) );
  OR U22722 ( .A(n22400), .B(n22399), .Z(n22404) );
  NANDN U22723 ( .A(n22402), .B(n22401), .Z(n22403) );
  NAND U22724 ( .A(n22404), .B(n22403), .Z(n22448) );
  NAND U22725 ( .A(a[42]), .B(b[62]), .Z(n22447) );
  XOR U22726 ( .A(n22448), .B(n22447), .Z(n22449) );
  NAND U22727 ( .A(b[63]), .B(a[41]), .Z(n22450) );
  XOR U22728 ( .A(n22449), .B(n22450), .Z(n22456) );
  XNOR U22729 ( .A(n22455), .B(n22456), .Z(n22461) );
  OR U22730 ( .A(n22406), .B(n22405), .Z(n22410) );
  NANDN U22731 ( .A(n22408), .B(n22407), .Z(n22409) );
  NAND U22732 ( .A(n22410), .B(n22409), .Z(n22460) );
  NAND U22733 ( .A(b[60]), .B(a[44]), .Z(n22459) );
  XOR U22734 ( .A(n22460), .B(n22459), .Z(n22462) );
  XOR U22735 ( .A(n22461), .B(n22462), .Z(n22465) );
  XNOR U22736 ( .A(n22466), .B(n22465), .Z(n22468) );
  NAND U22737 ( .A(b[59]), .B(a[45]), .Z(n22467) );
  XOR U22738 ( .A(n22468), .B(n22467), .Z(n22474) );
  XOR U22739 ( .A(n22473), .B(n22474), .Z(n22479) );
  AND U22740 ( .A(a[47]), .B(b[57]), .Z(n22477) );
  OR U22741 ( .A(n22412), .B(n22411), .Z(n22416) );
  NANDN U22742 ( .A(n22414), .B(n22413), .Z(n22415) );
  NAND U22743 ( .A(n22416), .B(n22415), .Z(n22478) );
  XOR U22744 ( .A(n22477), .B(n22478), .Z(n22480) );
  XOR U22745 ( .A(n22479), .B(n22480), .Z(n22484) );
  OR U22746 ( .A(n22418), .B(n22417), .Z(n22422) );
  NANDN U22747 ( .A(n22420), .B(n22419), .Z(n22421) );
  NAND U22748 ( .A(n22422), .B(n22421), .Z(n22482) );
  NAND U22749 ( .A(b[56]), .B(a[48]), .Z(n22481) );
  XOR U22750 ( .A(n22482), .B(n22481), .Z(n22483) );
  XOR U22751 ( .A(n22484), .B(n22483), .Z(n22487) );
  XNOR U22752 ( .A(n22488), .B(n22487), .Z(n22490) );
  NAND U22753 ( .A(b[55]), .B(a[49]), .Z(n22489) );
  XOR U22754 ( .A(n22490), .B(n22489), .Z(n22496) );
  XOR U22755 ( .A(n22495), .B(n22496), .Z(n22499) );
  XNOR U22756 ( .A(n22500), .B(n22499), .Z(n22502) );
  NAND U22757 ( .A(b[53]), .B(a[51]), .Z(n22501) );
  XOR U22758 ( .A(n22502), .B(n22501), .Z(n22508) );
  XOR U22759 ( .A(n22507), .B(n22508), .Z(n22511) );
  XNOR U22760 ( .A(n22512), .B(n22511), .Z(n22514) );
  NAND U22761 ( .A(b[51]), .B(a[53]), .Z(n22513) );
  XOR U22762 ( .A(n22514), .B(n22513), .Z(n22520) );
  XOR U22763 ( .A(n22519), .B(n22520), .Z(n22523) );
  XNOR U22764 ( .A(n22524), .B(n22523), .Z(n22526) );
  NAND U22765 ( .A(b[49]), .B(a[55]), .Z(n22525) );
  XOR U22766 ( .A(n22526), .B(n22525), .Z(n22532) );
  XOR U22767 ( .A(n22531), .B(n22532), .Z(n22535) );
  XNOR U22768 ( .A(n22536), .B(n22535), .Z(n22538) );
  NAND U22769 ( .A(b[47]), .B(a[57]), .Z(n22537) );
  XOR U22770 ( .A(n22538), .B(n22537), .Z(n22543) );
  OR U22771 ( .A(n22424), .B(n22423), .Z(n22428) );
  NANDN U22772 ( .A(n22426), .B(n22425), .Z(n22427) );
  NAND U22773 ( .A(n22428), .B(n22427), .Z(n22542) );
  NAND U22774 ( .A(b[46]), .B(a[58]), .Z(n22541) );
  XOR U22775 ( .A(n22542), .B(n22541), .Z(n22544) );
  XOR U22776 ( .A(n22543), .B(n22544), .Z(n22547) );
  XNOR U22777 ( .A(n22548), .B(n22547), .Z(n22550) );
  NAND U22778 ( .A(b[45]), .B(a[59]), .Z(n22549) );
  XOR U22779 ( .A(n22550), .B(n22549), .Z(n22556) );
  XOR U22780 ( .A(n22555), .B(n22556), .Z(n22559) );
  XNOR U22781 ( .A(n22560), .B(n22559), .Z(n22562) );
  NAND U22782 ( .A(b[43]), .B(a[61]), .Z(n22561) );
  XOR U22783 ( .A(n22562), .B(n22561), .Z(n22568) );
  XOR U22784 ( .A(n22567), .B(n22568), .Z(n22571) );
  OR U22785 ( .A(n22430), .B(n22429), .Z(n22434) );
  NANDN U22786 ( .A(n22432), .B(n22431), .Z(n22433) );
  NAND U22787 ( .A(n22434), .B(n22433), .Z(n22572) );
  XOR U22788 ( .A(n22571), .B(n22572), .Z(n22573) );
  XOR U22789 ( .A(n22574), .B(n22573), .Z(n22446) );
  OR U22790 ( .A(n22436), .B(n22435), .Z(n22440) );
  NANDN U22791 ( .A(n22438), .B(n22437), .Z(n22439) );
  NAND U22792 ( .A(n22440), .B(n22439), .Z(n22445) );
  XOR U22793 ( .A(n22446), .B(n22445), .Z(n22578) );
  XOR U22794 ( .A(n22577), .B(n22578), .Z(n22579) );
  XOR U22795 ( .A(n22579), .B(n22580), .Z(c[104]) );
  NOR U22796 ( .A(n22446), .B(n22445), .Z(n22581) );
  AND U22797 ( .A(b[63]), .B(a[42]), .Z(n22668) );
  AND U22798 ( .A(b[62]), .B(a[43]), .Z(n22665) );
  OR U22799 ( .A(n22448), .B(n22447), .Z(n22452) );
  NANDN U22800 ( .A(n22450), .B(n22449), .Z(n22451) );
  NAND U22801 ( .A(n22452), .B(n22451), .Z(n22666) );
  XOR U22802 ( .A(n22665), .B(n22666), .Z(n22667) );
  XOR U22803 ( .A(n22668), .B(n22667), .Z(n22662) );
  NANDN U22804 ( .A(n22454), .B(n22453), .Z(n22458) );
  NANDN U22805 ( .A(n22456), .B(n22455), .Z(n22457) );
  NAND U22806 ( .A(n22458), .B(n22457), .Z(n22659) );
  NAND U22807 ( .A(a[44]), .B(b[61]), .Z(n22660) );
  XNOR U22808 ( .A(n22659), .B(n22660), .Z(n22661) );
  XOR U22809 ( .A(n22662), .B(n22661), .Z(n22656) );
  AND U22810 ( .A(a[45]), .B(b[60]), .Z(n22653) );
  OR U22811 ( .A(n22460), .B(n22459), .Z(n22464) );
  NAND U22812 ( .A(n22462), .B(n22461), .Z(n22463) );
  NAND U22813 ( .A(n22464), .B(n22463), .Z(n22654) );
  XOR U22814 ( .A(n22653), .B(n22654), .Z(n22655) );
  XNOR U22815 ( .A(n22656), .B(n22655), .Z(n22650) );
  NAND U22816 ( .A(n22466), .B(n22465), .Z(n22470) );
  OR U22817 ( .A(n22468), .B(n22467), .Z(n22469) );
  NAND U22818 ( .A(n22470), .B(n22469), .Z(n22647) );
  NAND U22819 ( .A(a[46]), .B(b[59]), .Z(n22648) );
  XNOR U22820 ( .A(n22647), .B(n22648), .Z(n22649) );
  XNOR U22821 ( .A(n22650), .B(n22649), .Z(n22644) );
  AND U22822 ( .A(a[47]), .B(b[58]), .Z(n22641) );
  OR U22823 ( .A(n22472), .B(n22471), .Z(n22476) );
  NAND U22824 ( .A(n22474), .B(n22473), .Z(n22475) );
  NAND U22825 ( .A(n22476), .B(n22475), .Z(n22642) );
  XOR U22826 ( .A(n22641), .B(n22642), .Z(n22643) );
  XNOR U22827 ( .A(n22644), .B(n22643), .Z(n22638) );
  NAND U22828 ( .A(b[57]), .B(a[48]), .Z(n22635) );
  XOR U22829 ( .A(n22636), .B(n22635), .Z(n22637) );
  XNOR U22830 ( .A(n22638), .B(n22637), .Z(n22632) );
  AND U22831 ( .A(a[49]), .B(b[56]), .Z(n22629) );
  OR U22832 ( .A(n22482), .B(n22481), .Z(n22486) );
  NAND U22833 ( .A(n22484), .B(n22483), .Z(n22485) );
  NAND U22834 ( .A(n22486), .B(n22485), .Z(n22630) );
  XOR U22835 ( .A(n22629), .B(n22630), .Z(n22631) );
  XNOR U22836 ( .A(n22632), .B(n22631), .Z(n22626) );
  NAND U22837 ( .A(n22488), .B(n22487), .Z(n22492) );
  OR U22838 ( .A(n22490), .B(n22489), .Z(n22491) );
  NAND U22839 ( .A(n22492), .B(n22491), .Z(n22623) );
  NAND U22840 ( .A(a[50]), .B(b[55]), .Z(n22624) );
  XNOR U22841 ( .A(n22623), .B(n22624), .Z(n22625) );
  XNOR U22842 ( .A(n22626), .B(n22625), .Z(n22620) );
  AND U22843 ( .A(a[51]), .B(b[54]), .Z(n22617) );
  OR U22844 ( .A(n22494), .B(n22493), .Z(n22498) );
  NAND U22845 ( .A(n22496), .B(n22495), .Z(n22497) );
  NAND U22846 ( .A(n22498), .B(n22497), .Z(n22618) );
  XOR U22847 ( .A(n22617), .B(n22618), .Z(n22619) );
  XNOR U22848 ( .A(n22620), .B(n22619), .Z(n22674) );
  NAND U22849 ( .A(n22500), .B(n22499), .Z(n22504) );
  OR U22850 ( .A(n22502), .B(n22501), .Z(n22503) );
  NAND U22851 ( .A(n22504), .B(n22503), .Z(n22671) );
  NAND U22852 ( .A(a[52]), .B(b[53]), .Z(n22672) );
  XNOR U22853 ( .A(n22671), .B(n22672), .Z(n22673) );
  XNOR U22854 ( .A(n22674), .B(n22673), .Z(n22680) );
  AND U22855 ( .A(a[53]), .B(b[52]), .Z(n22677) );
  OR U22856 ( .A(n22506), .B(n22505), .Z(n22510) );
  NAND U22857 ( .A(n22508), .B(n22507), .Z(n22509) );
  NAND U22858 ( .A(n22510), .B(n22509), .Z(n22678) );
  XOR U22859 ( .A(n22677), .B(n22678), .Z(n22679) );
  XNOR U22860 ( .A(n22680), .B(n22679), .Z(n22686) );
  NAND U22861 ( .A(n22512), .B(n22511), .Z(n22516) );
  OR U22862 ( .A(n22514), .B(n22513), .Z(n22515) );
  NAND U22863 ( .A(n22516), .B(n22515), .Z(n22683) );
  NAND U22864 ( .A(a[54]), .B(b[51]), .Z(n22684) );
  XNOR U22865 ( .A(n22683), .B(n22684), .Z(n22685) );
  XNOR U22866 ( .A(n22686), .B(n22685), .Z(n22692) );
  AND U22867 ( .A(a[55]), .B(b[50]), .Z(n22689) );
  OR U22868 ( .A(n22518), .B(n22517), .Z(n22522) );
  NAND U22869 ( .A(n22520), .B(n22519), .Z(n22521) );
  NAND U22870 ( .A(n22522), .B(n22521), .Z(n22690) );
  XOR U22871 ( .A(n22689), .B(n22690), .Z(n22691) );
  XNOR U22872 ( .A(n22692), .B(n22691), .Z(n22614) );
  NAND U22873 ( .A(n22524), .B(n22523), .Z(n22528) );
  OR U22874 ( .A(n22526), .B(n22525), .Z(n22527) );
  NAND U22875 ( .A(n22528), .B(n22527), .Z(n22611) );
  NAND U22876 ( .A(a[56]), .B(b[49]), .Z(n22612) );
  XNOR U22877 ( .A(n22611), .B(n22612), .Z(n22613) );
  XNOR U22878 ( .A(n22614), .B(n22613), .Z(n22698) );
  AND U22879 ( .A(a[57]), .B(b[48]), .Z(n22695) );
  OR U22880 ( .A(n22530), .B(n22529), .Z(n22534) );
  NAND U22881 ( .A(n22532), .B(n22531), .Z(n22533) );
  NAND U22882 ( .A(n22534), .B(n22533), .Z(n22696) );
  XOR U22883 ( .A(n22695), .B(n22696), .Z(n22697) );
  XNOR U22884 ( .A(n22698), .B(n22697), .Z(n22608) );
  NAND U22885 ( .A(n22536), .B(n22535), .Z(n22540) );
  OR U22886 ( .A(n22538), .B(n22537), .Z(n22539) );
  NAND U22887 ( .A(n22540), .B(n22539), .Z(n22605) );
  NAND U22888 ( .A(a[58]), .B(b[47]), .Z(n22606) );
  XNOR U22889 ( .A(n22605), .B(n22606), .Z(n22607) );
  XNOR U22890 ( .A(n22608), .B(n22607), .Z(n22602) );
  AND U22891 ( .A(a[59]), .B(b[46]), .Z(n22599) );
  OR U22892 ( .A(n22542), .B(n22541), .Z(n22546) );
  NAND U22893 ( .A(n22544), .B(n22543), .Z(n22545) );
  NAND U22894 ( .A(n22546), .B(n22545), .Z(n22600) );
  XOR U22895 ( .A(n22599), .B(n22600), .Z(n22601) );
  XNOR U22896 ( .A(n22602), .B(n22601), .Z(n22596) );
  NAND U22897 ( .A(n22548), .B(n22547), .Z(n22552) );
  OR U22898 ( .A(n22550), .B(n22549), .Z(n22551) );
  NAND U22899 ( .A(n22552), .B(n22551), .Z(n22593) );
  NAND U22900 ( .A(a[60]), .B(b[45]), .Z(n22594) );
  XNOR U22901 ( .A(n22593), .B(n22594), .Z(n22595) );
  XNOR U22902 ( .A(n22596), .B(n22595), .Z(n22590) );
  AND U22903 ( .A(a[61]), .B(b[44]), .Z(n22587) );
  OR U22904 ( .A(n22554), .B(n22553), .Z(n22558) );
  NAND U22905 ( .A(n22556), .B(n22555), .Z(n22557) );
  NAND U22906 ( .A(n22558), .B(n22557), .Z(n22588) );
  XOR U22907 ( .A(n22587), .B(n22588), .Z(n22589) );
  XNOR U22908 ( .A(n22590), .B(n22589), .Z(n22704) );
  NAND U22909 ( .A(n22560), .B(n22559), .Z(n22564) );
  OR U22910 ( .A(n22562), .B(n22561), .Z(n22563) );
  NAND U22911 ( .A(n22564), .B(n22563), .Z(n22701) );
  NAND U22912 ( .A(a[62]), .B(b[43]), .Z(n22702) );
  XNOR U22913 ( .A(n22701), .B(n22702), .Z(n22703) );
  XOR U22914 ( .A(n22704), .B(n22703), .Z(n22709) );
  NAND U22915 ( .A(b[42]), .B(a[63]), .Z(n22708) );
  OR U22916 ( .A(n22566), .B(n22565), .Z(n22570) );
  NAND U22917 ( .A(n22568), .B(n22567), .Z(n22569) );
  AND U22918 ( .A(n22570), .B(n22569), .Z(n22707) );
  XNOR U22919 ( .A(n22708), .B(n22707), .Z(n22710) );
  XNOR U22920 ( .A(n22709), .B(n22710), .Z(n22585) );
  NAND U22921 ( .A(n22572), .B(n22571), .Z(n22576) );
  NANDN U22922 ( .A(n22574), .B(n22573), .Z(n22575) );
  NAND U22923 ( .A(n22576), .B(n22575), .Z(n22586) );
  XNOR U22924 ( .A(n22585), .B(n22586), .Z(n22582) );
  XOR U22925 ( .A(n22581), .B(n22582), .Z(n22583) );
  XOR U22926 ( .A(n22583), .B(n22584), .Z(c[105]) );
  ANDN U22927 ( .B(n22586), .A(n22585), .Z(n22955) );
  NANDN U22928 ( .A(n156), .B(a[63]), .Z(n22833) );
  OR U22929 ( .A(n22588), .B(n22587), .Z(n22592) );
  NANDN U22930 ( .A(n22590), .B(n22589), .Z(n22591) );
  NAND U22931 ( .A(n22592), .B(n22591), .Z(n22825) );
  NAND U22932 ( .A(b[44]), .B(a[62]), .Z(n22824) );
  XOR U22933 ( .A(n22825), .B(n22824), .Z(n22826) );
  NANDN U22934 ( .A(n22594), .B(n22593), .Z(n22598) );
  NANDN U22935 ( .A(n22596), .B(n22595), .Z(n22597) );
  NAND U22936 ( .A(n22598), .B(n22597), .Z(n22819) );
  OR U22937 ( .A(n22600), .B(n22599), .Z(n22604) );
  NANDN U22938 ( .A(n22602), .B(n22601), .Z(n22603) );
  NAND U22939 ( .A(n22604), .B(n22603), .Z(n22813) );
  NAND U22940 ( .A(b[46]), .B(a[60]), .Z(n22812) );
  XOR U22941 ( .A(n22813), .B(n22812), .Z(n22814) );
  NANDN U22942 ( .A(n22606), .B(n22605), .Z(n22610) );
  NANDN U22943 ( .A(n22608), .B(n22607), .Z(n22609) );
  NAND U22944 ( .A(n22610), .B(n22609), .Z(n22807) );
  NANDN U22945 ( .A(n22612), .B(n22611), .Z(n22616) );
  NANDN U22946 ( .A(n22614), .B(n22613), .Z(n22615) );
  NAND U22947 ( .A(n22616), .B(n22615), .Z(n22795) );
  AND U22948 ( .A(a[55]), .B(b[51]), .Z(n22785) );
  AND U22949 ( .A(a[53]), .B(b[53]), .Z(n22775) );
  OR U22950 ( .A(n22618), .B(n22617), .Z(n22622) );
  NANDN U22951 ( .A(n22620), .B(n22619), .Z(n22621) );
  NAND U22952 ( .A(n22622), .B(n22621), .Z(n22767) );
  NAND U22953 ( .A(b[54]), .B(a[52]), .Z(n22766) );
  XOR U22954 ( .A(n22767), .B(n22766), .Z(n22768) );
  NANDN U22955 ( .A(n22624), .B(n22623), .Z(n22628) );
  NANDN U22956 ( .A(n22626), .B(n22625), .Z(n22627) );
  NAND U22957 ( .A(n22628), .B(n22627), .Z(n22761) );
  OR U22958 ( .A(n22630), .B(n22629), .Z(n22634) );
  NANDN U22959 ( .A(n22632), .B(n22631), .Z(n22633) );
  NAND U22960 ( .A(n22634), .B(n22633), .Z(n22755) );
  NAND U22961 ( .A(b[56]), .B(a[50]), .Z(n22754) );
  XOR U22962 ( .A(n22755), .B(n22754), .Z(n22756) );
  OR U22963 ( .A(n22636), .B(n22635), .Z(n22640) );
  NANDN U22964 ( .A(n22638), .B(n22637), .Z(n22639) );
  NAND U22965 ( .A(n22640), .B(n22639), .Z(n22748) );
  NAND U22966 ( .A(a[49]), .B(b[57]), .Z(n22749) );
  XNOR U22967 ( .A(n22748), .B(n22749), .Z(n22750) );
  OR U22968 ( .A(n22642), .B(n22641), .Z(n22646) );
  NANDN U22969 ( .A(n22644), .B(n22643), .Z(n22645) );
  NAND U22970 ( .A(n22646), .B(n22645), .Z(n22743) );
  NAND U22971 ( .A(b[58]), .B(a[48]), .Z(n22742) );
  XOR U22972 ( .A(n22743), .B(n22742), .Z(n22744) );
  NANDN U22973 ( .A(n22648), .B(n22647), .Z(n22652) );
  NANDN U22974 ( .A(n22650), .B(n22649), .Z(n22651) );
  NAND U22975 ( .A(n22652), .B(n22651), .Z(n22737) );
  OR U22976 ( .A(n22654), .B(n22653), .Z(n22658) );
  NANDN U22977 ( .A(n22656), .B(n22655), .Z(n22657) );
  NAND U22978 ( .A(n22658), .B(n22657), .Z(n22731) );
  NAND U22979 ( .A(b[60]), .B(a[46]), .Z(n22730) );
  XOR U22980 ( .A(n22731), .B(n22730), .Z(n22732) );
  NANDN U22981 ( .A(n22660), .B(n22659), .Z(n22664) );
  NAND U22982 ( .A(n22662), .B(n22661), .Z(n22663) );
  NAND U22983 ( .A(n22664), .B(n22663), .Z(n22727) );
  NAND U22984 ( .A(a[45]), .B(b[61]), .Z(n22724) );
  OR U22985 ( .A(n22666), .B(n22665), .Z(n22670) );
  NANDN U22986 ( .A(n22668), .B(n22667), .Z(n22669) );
  NAND U22987 ( .A(n22670), .B(n22669), .Z(n22719) );
  NAND U22988 ( .A(a[44]), .B(b[62]), .Z(n22718) );
  XOR U22989 ( .A(n22719), .B(n22718), .Z(n22720) );
  NAND U22990 ( .A(b[63]), .B(a[43]), .Z(n22721) );
  XOR U22991 ( .A(n22720), .B(n22721), .Z(n22725) );
  XOR U22992 ( .A(n22724), .B(n22725), .Z(n22726) );
  XOR U22993 ( .A(n22727), .B(n22726), .Z(n22733) );
  XOR U22994 ( .A(n22732), .B(n22733), .Z(n22736) );
  XNOR U22995 ( .A(n22737), .B(n22736), .Z(n22739) );
  NAND U22996 ( .A(b[59]), .B(a[47]), .Z(n22738) );
  XOR U22997 ( .A(n22739), .B(n22738), .Z(n22745) );
  XOR U22998 ( .A(n22744), .B(n22745), .Z(n22751) );
  XOR U22999 ( .A(n22750), .B(n22751), .Z(n22757) );
  XOR U23000 ( .A(n22756), .B(n22757), .Z(n22760) );
  XNOR U23001 ( .A(n22761), .B(n22760), .Z(n22763) );
  NAND U23002 ( .A(b[55]), .B(a[51]), .Z(n22762) );
  XOR U23003 ( .A(n22763), .B(n22762), .Z(n22769) );
  XOR U23004 ( .A(n22768), .B(n22769), .Z(n22772) );
  NANDN U23005 ( .A(n22672), .B(n22671), .Z(n22676) );
  NANDN U23006 ( .A(n22674), .B(n22673), .Z(n22675) );
  NAND U23007 ( .A(n22676), .B(n22675), .Z(n22773) );
  XOR U23008 ( .A(n22772), .B(n22773), .Z(n22774) );
  XOR U23009 ( .A(n22775), .B(n22774), .Z(n22779) );
  OR U23010 ( .A(n22678), .B(n22677), .Z(n22682) );
  NANDN U23011 ( .A(n22680), .B(n22679), .Z(n22681) );
  NAND U23012 ( .A(n22682), .B(n22681), .Z(n22777) );
  NAND U23013 ( .A(b[52]), .B(a[54]), .Z(n22776) );
  XOR U23014 ( .A(n22777), .B(n22776), .Z(n22778) );
  XOR U23015 ( .A(n22779), .B(n22778), .Z(n22782) );
  NANDN U23016 ( .A(n22684), .B(n22683), .Z(n22688) );
  NANDN U23017 ( .A(n22686), .B(n22685), .Z(n22687) );
  NAND U23018 ( .A(n22688), .B(n22687), .Z(n22783) );
  XOR U23019 ( .A(n22782), .B(n22783), .Z(n22784) );
  XOR U23020 ( .A(n22785), .B(n22784), .Z(n22791) );
  OR U23021 ( .A(n22690), .B(n22689), .Z(n22694) );
  NANDN U23022 ( .A(n22692), .B(n22691), .Z(n22693) );
  NAND U23023 ( .A(n22694), .B(n22693), .Z(n22789) );
  NAND U23024 ( .A(b[50]), .B(a[56]), .Z(n22788) );
  XOR U23025 ( .A(n22789), .B(n22788), .Z(n22790) );
  XOR U23026 ( .A(n22791), .B(n22790), .Z(n22794) );
  XNOR U23027 ( .A(n22795), .B(n22794), .Z(n22797) );
  NAND U23028 ( .A(b[49]), .B(a[57]), .Z(n22796) );
  XOR U23029 ( .A(n22797), .B(n22796), .Z(n22802) );
  OR U23030 ( .A(n22696), .B(n22695), .Z(n22700) );
  NANDN U23031 ( .A(n22698), .B(n22697), .Z(n22699) );
  NAND U23032 ( .A(n22700), .B(n22699), .Z(n22801) );
  NAND U23033 ( .A(b[48]), .B(a[58]), .Z(n22800) );
  XOR U23034 ( .A(n22801), .B(n22800), .Z(n22803) );
  XOR U23035 ( .A(n22802), .B(n22803), .Z(n22806) );
  XNOR U23036 ( .A(n22807), .B(n22806), .Z(n22809) );
  NAND U23037 ( .A(b[47]), .B(a[59]), .Z(n22808) );
  XOR U23038 ( .A(n22809), .B(n22808), .Z(n22815) );
  XOR U23039 ( .A(n22814), .B(n22815), .Z(n22818) );
  XNOR U23040 ( .A(n22819), .B(n22818), .Z(n22821) );
  NAND U23041 ( .A(b[45]), .B(a[61]), .Z(n22820) );
  XOR U23042 ( .A(n22821), .B(n22820), .Z(n22827) );
  XOR U23043 ( .A(n22826), .B(n22827), .Z(n22830) );
  NANDN U23044 ( .A(n22702), .B(n22701), .Z(n22706) );
  NANDN U23045 ( .A(n22704), .B(n22703), .Z(n22705) );
  NAND U23046 ( .A(n22706), .B(n22705), .Z(n22831) );
  XOR U23047 ( .A(n22830), .B(n22831), .Z(n22832) );
  XOR U23048 ( .A(n22833), .B(n22832), .Z(n22717) );
  NAND U23049 ( .A(n22708), .B(n22707), .Z(n22712) );
  NANDN U23050 ( .A(n22710), .B(n22709), .Z(n22711) );
  NAND U23051 ( .A(n22712), .B(n22711), .Z(n22716) );
  XNOR U23052 ( .A(n22717), .B(n22716), .Z(n22714) );
  XNOR U23053 ( .A(n22955), .B(n22714), .Z(n22713) );
  XNOR U23054 ( .A(n22952), .B(n22713), .Z(c[106]) );
  NAND U23055 ( .A(n22713), .B(n22952), .Z(n22715) );
  IV U23056 ( .A(n22714), .Z(n22954) );
  NOR U23057 ( .A(n22954), .B(n22955), .Z(n22953) );
  ANDN U23058 ( .B(n22715), .A(n22953), .Z(n22835) );
  OR U23059 ( .A(n22717), .B(n22716), .Z(n22961) );
  AND U23060 ( .A(b[63]), .B(a[44]), .Z(n22893) );
  AND U23061 ( .A(b[62]), .B(a[45]), .Z(n22891) );
  OR U23062 ( .A(n22719), .B(n22718), .Z(n22723) );
  NANDN U23063 ( .A(n22721), .B(n22720), .Z(n22722) );
  AND U23064 ( .A(n22723), .B(n22722), .Z(n22890) );
  XNOR U23065 ( .A(n22891), .B(n22890), .Z(n22892) );
  XOR U23066 ( .A(n22893), .B(n22892), .Z(n22899) );
  OR U23067 ( .A(n22725), .B(n22724), .Z(n22729) );
  NAND U23068 ( .A(n22727), .B(n22726), .Z(n22728) );
  NAND U23069 ( .A(n22729), .B(n22728), .Z(n22896) );
  NAND U23070 ( .A(a[46]), .B(b[61]), .Z(n22897) );
  XNOR U23071 ( .A(n22896), .B(n22897), .Z(n22898) );
  XOR U23072 ( .A(n22899), .B(n22898), .Z(n22905) );
  AND U23073 ( .A(a[47]), .B(b[60]), .Z(n22902) );
  OR U23074 ( .A(n22731), .B(n22730), .Z(n22735) );
  NAND U23075 ( .A(n22733), .B(n22732), .Z(n22734) );
  NAND U23076 ( .A(n22735), .B(n22734), .Z(n22903) );
  XOR U23077 ( .A(n22902), .B(n22903), .Z(n22904) );
  XNOR U23078 ( .A(n22905), .B(n22904), .Z(n22887) );
  NAND U23079 ( .A(n22737), .B(n22736), .Z(n22741) );
  OR U23080 ( .A(n22739), .B(n22738), .Z(n22740) );
  NAND U23081 ( .A(n22741), .B(n22740), .Z(n22884) );
  NAND U23082 ( .A(a[48]), .B(b[59]), .Z(n22885) );
  XNOR U23083 ( .A(n22884), .B(n22885), .Z(n22886) );
  XNOR U23084 ( .A(n22887), .B(n22886), .Z(n22881) );
  AND U23085 ( .A(a[49]), .B(b[58]), .Z(n22878) );
  OR U23086 ( .A(n22743), .B(n22742), .Z(n22747) );
  NAND U23087 ( .A(n22745), .B(n22744), .Z(n22746) );
  NAND U23088 ( .A(n22747), .B(n22746), .Z(n22879) );
  XOR U23089 ( .A(n22878), .B(n22879), .Z(n22880) );
  XNOR U23090 ( .A(n22881), .B(n22880), .Z(n22911) );
  NANDN U23091 ( .A(n22749), .B(n22748), .Z(n22753) );
  NAND U23092 ( .A(n22751), .B(n22750), .Z(n22752) );
  NAND U23093 ( .A(n22753), .B(n22752), .Z(n22908) );
  NAND U23094 ( .A(a[50]), .B(b[57]), .Z(n22909) );
  XNOR U23095 ( .A(n22908), .B(n22909), .Z(n22910) );
  XNOR U23096 ( .A(n22911), .B(n22910), .Z(n22917) );
  AND U23097 ( .A(a[51]), .B(b[56]), .Z(n22914) );
  OR U23098 ( .A(n22755), .B(n22754), .Z(n22759) );
  NAND U23099 ( .A(n22757), .B(n22756), .Z(n22758) );
  NAND U23100 ( .A(n22759), .B(n22758), .Z(n22915) );
  XOR U23101 ( .A(n22914), .B(n22915), .Z(n22916) );
  XNOR U23102 ( .A(n22917), .B(n22916), .Z(n22923) );
  NAND U23103 ( .A(n22761), .B(n22760), .Z(n22765) );
  OR U23104 ( .A(n22763), .B(n22762), .Z(n22764) );
  NAND U23105 ( .A(n22765), .B(n22764), .Z(n22920) );
  NAND U23106 ( .A(a[52]), .B(b[55]), .Z(n22921) );
  XNOR U23107 ( .A(n22920), .B(n22921), .Z(n22922) );
  XNOR U23108 ( .A(n22923), .B(n22922), .Z(n22929) );
  AND U23109 ( .A(a[53]), .B(b[54]), .Z(n22926) );
  OR U23110 ( .A(n22767), .B(n22766), .Z(n22771) );
  NAND U23111 ( .A(n22769), .B(n22768), .Z(n22770) );
  NAND U23112 ( .A(n22771), .B(n22770), .Z(n22927) );
  XOR U23113 ( .A(n22926), .B(n22927), .Z(n22928) );
  XNOR U23114 ( .A(n22929), .B(n22928), .Z(n22875) );
  NAND U23115 ( .A(b[53]), .B(a[54]), .Z(n22872) );
  XOR U23116 ( .A(n22873), .B(n22872), .Z(n22874) );
  XNOR U23117 ( .A(n22875), .B(n22874), .Z(n22869) );
  AND U23118 ( .A(a[55]), .B(b[52]), .Z(n22866) );
  OR U23119 ( .A(n22777), .B(n22776), .Z(n22781) );
  NAND U23120 ( .A(n22779), .B(n22778), .Z(n22780) );
  NAND U23121 ( .A(n22781), .B(n22780), .Z(n22867) );
  XOR U23122 ( .A(n22866), .B(n22867), .Z(n22868) );
  XNOR U23123 ( .A(n22869), .B(n22868), .Z(n22863) );
  OR U23124 ( .A(n22783), .B(n22782), .Z(n22787) );
  NANDN U23125 ( .A(n22785), .B(n22784), .Z(n22786) );
  NAND U23126 ( .A(n22787), .B(n22786), .Z(n22861) );
  NAND U23127 ( .A(b[51]), .B(a[56]), .Z(n22860) );
  XOR U23128 ( .A(n22861), .B(n22860), .Z(n22862) );
  XNOR U23129 ( .A(n22863), .B(n22862), .Z(n22857) );
  AND U23130 ( .A(a[57]), .B(b[50]), .Z(n22854) );
  OR U23131 ( .A(n22789), .B(n22788), .Z(n22793) );
  NAND U23132 ( .A(n22791), .B(n22790), .Z(n22792) );
  NAND U23133 ( .A(n22793), .B(n22792), .Z(n22855) );
  XOR U23134 ( .A(n22854), .B(n22855), .Z(n22856) );
  XNOR U23135 ( .A(n22857), .B(n22856), .Z(n22851) );
  NAND U23136 ( .A(n22795), .B(n22794), .Z(n22799) );
  OR U23137 ( .A(n22797), .B(n22796), .Z(n22798) );
  NAND U23138 ( .A(n22799), .B(n22798), .Z(n22848) );
  NAND U23139 ( .A(a[58]), .B(b[49]), .Z(n22849) );
  XNOR U23140 ( .A(n22848), .B(n22849), .Z(n22850) );
  XNOR U23141 ( .A(n22851), .B(n22850), .Z(n22845) );
  AND U23142 ( .A(a[59]), .B(b[48]), .Z(n22842) );
  OR U23143 ( .A(n22801), .B(n22800), .Z(n22805) );
  NAND U23144 ( .A(n22803), .B(n22802), .Z(n22804) );
  NAND U23145 ( .A(n22805), .B(n22804), .Z(n22843) );
  XOR U23146 ( .A(n22842), .B(n22843), .Z(n22844) );
  XNOR U23147 ( .A(n22845), .B(n22844), .Z(n22935) );
  NAND U23148 ( .A(n22807), .B(n22806), .Z(n22811) );
  OR U23149 ( .A(n22809), .B(n22808), .Z(n22810) );
  NAND U23150 ( .A(n22811), .B(n22810), .Z(n22932) );
  NAND U23151 ( .A(a[60]), .B(b[47]), .Z(n22933) );
  XNOR U23152 ( .A(n22932), .B(n22933), .Z(n22934) );
  XNOR U23153 ( .A(n22935), .B(n22934), .Z(n22941) );
  AND U23154 ( .A(a[61]), .B(b[46]), .Z(n22938) );
  OR U23155 ( .A(n22813), .B(n22812), .Z(n22817) );
  NAND U23156 ( .A(n22815), .B(n22814), .Z(n22816) );
  NAND U23157 ( .A(n22817), .B(n22816), .Z(n22939) );
  XOR U23158 ( .A(n22938), .B(n22939), .Z(n22940) );
  XNOR U23159 ( .A(n22941), .B(n22940), .Z(n22839) );
  NAND U23160 ( .A(n22819), .B(n22818), .Z(n22823) );
  OR U23161 ( .A(n22821), .B(n22820), .Z(n22822) );
  NAND U23162 ( .A(n22823), .B(n22822), .Z(n22836) );
  NAND U23163 ( .A(a[62]), .B(b[45]), .Z(n22837) );
  XNOR U23164 ( .A(n22836), .B(n22837), .Z(n22838) );
  XNOR U23165 ( .A(n22839), .B(n22838), .Z(n22947) );
  AND U23166 ( .A(a[63]), .B(b[44]), .Z(n22944) );
  OR U23167 ( .A(n22825), .B(n22824), .Z(n22829) );
  NAND U23168 ( .A(n22827), .B(n22826), .Z(n22828) );
  NAND U23169 ( .A(n22829), .B(n22828), .Z(n22945) );
  XOR U23170 ( .A(n22944), .B(n22945), .Z(n22946) );
  XNOR U23171 ( .A(n22947), .B(n22946), .Z(n22950) );
  XOR U23172 ( .A(n22950), .B(n22951), .Z(n22959) );
  XOR U23173 ( .A(n22961), .B(n22959), .Z(n22834) );
  XNOR U23174 ( .A(n22835), .B(n22834), .Z(c[107]) );
  NANDN U23175 ( .A(n22837), .B(n22836), .Z(n22841) );
  NANDN U23176 ( .A(n22839), .B(n22838), .Z(n22840) );
  NAND U23177 ( .A(n22841), .B(n22840), .Z(n23071) );
  AND U23178 ( .A(a[61]), .B(b[47]), .Z(n23063) );
  OR U23179 ( .A(n22843), .B(n22842), .Z(n22847) );
  NANDN U23180 ( .A(n22845), .B(n22844), .Z(n22846) );
  NAND U23181 ( .A(n22847), .B(n22846), .Z(n23055) );
  NAND U23182 ( .A(b[48]), .B(a[60]), .Z(n23054) );
  XOR U23183 ( .A(n23055), .B(n23054), .Z(n23056) );
  NANDN U23184 ( .A(n22849), .B(n22848), .Z(n22853) );
  NANDN U23185 ( .A(n22851), .B(n22850), .Z(n22852) );
  NAND U23186 ( .A(n22853), .B(n22852), .Z(n23049) );
  OR U23187 ( .A(n22855), .B(n22854), .Z(n22859) );
  NANDN U23188 ( .A(n22857), .B(n22856), .Z(n22858) );
  NAND U23189 ( .A(n22859), .B(n22858), .Z(n23043) );
  NAND U23190 ( .A(b[50]), .B(a[58]), .Z(n23042) );
  XOR U23191 ( .A(n23043), .B(n23042), .Z(n23044) );
  OR U23192 ( .A(n22861), .B(n22860), .Z(n22865) );
  NANDN U23193 ( .A(n22863), .B(n22862), .Z(n22864) );
  NAND U23194 ( .A(n22865), .B(n22864), .Z(n23037) );
  OR U23195 ( .A(n22867), .B(n22866), .Z(n22871) );
  NANDN U23196 ( .A(n22869), .B(n22868), .Z(n22870) );
  NAND U23197 ( .A(n22871), .B(n22870), .Z(n23031) );
  NAND U23198 ( .A(b[52]), .B(a[56]), .Z(n23030) );
  XOR U23199 ( .A(n23031), .B(n23030), .Z(n23032) );
  OR U23200 ( .A(n22873), .B(n22872), .Z(n22877) );
  NANDN U23201 ( .A(n22875), .B(n22874), .Z(n22876) );
  NAND U23202 ( .A(n22877), .B(n22876), .Z(n23025) );
  AND U23203 ( .A(a[53]), .B(b[55]), .Z(n23015) );
  AND U23204 ( .A(a[51]), .B(b[57]), .Z(n23005) );
  OR U23205 ( .A(n22879), .B(n22878), .Z(n22883) );
  NANDN U23206 ( .A(n22881), .B(n22880), .Z(n22882) );
  NAND U23207 ( .A(n22883), .B(n22882), .Z(n22997) );
  NAND U23208 ( .A(b[58]), .B(a[50]), .Z(n22996) );
  XOR U23209 ( .A(n22997), .B(n22996), .Z(n22998) );
  NANDN U23210 ( .A(n22885), .B(n22884), .Z(n22889) );
  NANDN U23211 ( .A(n22887), .B(n22886), .Z(n22888) );
  NAND U23212 ( .A(n22889), .B(n22888), .Z(n22991) );
  AND U23213 ( .A(a[47]), .B(b[61]), .Z(n22981) );
  NANDN U23214 ( .A(n22891), .B(n22890), .Z(n22895) );
  NANDN U23215 ( .A(n22893), .B(n22892), .Z(n22894) );
  NAND U23216 ( .A(n22895), .B(n22894), .Z(n22973) );
  NAND U23217 ( .A(a[46]), .B(b[62]), .Z(n22972) );
  XOR U23218 ( .A(n22973), .B(n22972), .Z(n22974) );
  NAND U23219 ( .A(a[45]), .B(b[63]), .Z(n22975) );
  XOR U23220 ( .A(n22974), .B(n22975), .Z(n22978) );
  NANDN U23221 ( .A(n22897), .B(n22896), .Z(n22901) );
  NAND U23222 ( .A(n22899), .B(n22898), .Z(n22900) );
  NAND U23223 ( .A(n22901), .B(n22900), .Z(n22979) );
  XNOR U23224 ( .A(n22978), .B(n22979), .Z(n22980) );
  XOR U23225 ( .A(n22981), .B(n22980), .Z(n22987) );
  OR U23226 ( .A(n22903), .B(n22902), .Z(n22907) );
  NANDN U23227 ( .A(n22905), .B(n22904), .Z(n22906) );
  NAND U23228 ( .A(n22907), .B(n22906), .Z(n22985) );
  NAND U23229 ( .A(b[60]), .B(a[48]), .Z(n22984) );
  XOR U23230 ( .A(n22985), .B(n22984), .Z(n22986) );
  XOR U23231 ( .A(n22987), .B(n22986), .Z(n22990) );
  XNOR U23232 ( .A(n22991), .B(n22990), .Z(n22993) );
  NAND U23233 ( .A(b[59]), .B(a[49]), .Z(n22992) );
  XOR U23234 ( .A(n22993), .B(n22992), .Z(n22999) );
  XOR U23235 ( .A(n22998), .B(n22999), .Z(n23002) );
  NANDN U23236 ( .A(n22909), .B(n22908), .Z(n22913) );
  NANDN U23237 ( .A(n22911), .B(n22910), .Z(n22912) );
  NAND U23238 ( .A(n22913), .B(n22912), .Z(n23003) );
  XOR U23239 ( .A(n23002), .B(n23003), .Z(n23004) );
  XOR U23240 ( .A(n23005), .B(n23004), .Z(n23009) );
  OR U23241 ( .A(n22915), .B(n22914), .Z(n22919) );
  NANDN U23242 ( .A(n22917), .B(n22916), .Z(n22918) );
  NAND U23243 ( .A(n22919), .B(n22918), .Z(n23007) );
  NAND U23244 ( .A(b[56]), .B(a[52]), .Z(n23006) );
  XOR U23245 ( .A(n23007), .B(n23006), .Z(n23008) );
  XOR U23246 ( .A(n23009), .B(n23008), .Z(n23012) );
  NANDN U23247 ( .A(n22921), .B(n22920), .Z(n22925) );
  NANDN U23248 ( .A(n22923), .B(n22922), .Z(n22924) );
  NAND U23249 ( .A(n22925), .B(n22924), .Z(n23013) );
  XOR U23250 ( .A(n23012), .B(n23013), .Z(n23014) );
  XOR U23251 ( .A(n23015), .B(n23014), .Z(n23021) );
  OR U23252 ( .A(n22927), .B(n22926), .Z(n22931) );
  NANDN U23253 ( .A(n22929), .B(n22928), .Z(n22930) );
  NAND U23254 ( .A(n22931), .B(n22930), .Z(n23019) );
  NAND U23255 ( .A(b[54]), .B(a[54]), .Z(n23018) );
  XOR U23256 ( .A(n23019), .B(n23018), .Z(n23020) );
  XOR U23257 ( .A(n23021), .B(n23020), .Z(n23024) );
  XNOR U23258 ( .A(n23025), .B(n23024), .Z(n23027) );
  NAND U23259 ( .A(b[53]), .B(a[55]), .Z(n23026) );
  XOR U23260 ( .A(n23027), .B(n23026), .Z(n23033) );
  XOR U23261 ( .A(n23032), .B(n23033), .Z(n23036) );
  XNOR U23262 ( .A(n23037), .B(n23036), .Z(n23039) );
  NAND U23263 ( .A(b[51]), .B(a[57]), .Z(n23038) );
  XOR U23264 ( .A(n23039), .B(n23038), .Z(n23045) );
  XOR U23265 ( .A(n23044), .B(n23045), .Z(n23048) );
  XNOR U23266 ( .A(n23049), .B(n23048), .Z(n23051) );
  NAND U23267 ( .A(b[49]), .B(a[59]), .Z(n23050) );
  XOR U23268 ( .A(n23051), .B(n23050), .Z(n23057) );
  XOR U23269 ( .A(n23056), .B(n23057), .Z(n23060) );
  NANDN U23270 ( .A(n22933), .B(n22932), .Z(n22937) );
  NANDN U23271 ( .A(n22935), .B(n22934), .Z(n22936) );
  NAND U23272 ( .A(n22937), .B(n22936), .Z(n23061) );
  XOR U23273 ( .A(n23060), .B(n23061), .Z(n23062) );
  XOR U23274 ( .A(n23063), .B(n23062), .Z(n23067) );
  OR U23275 ( .A(n22939), .B(n22938), .Z(n22943) );
  NANDN U23276 ( .A(n22941), .B(n22940), .Z(n22942) );
  NAND U23277 ( .A(n22943), .B(n22942), .Z(n23065) );
  NAND U23278 ( .A(b[46]), .B(a[62]), .Z(n23064) );
  XOR U23279 ( .A(n23065), .B(n23064), .Z(n23066) );
  XOR U23280 ( .A(n23067), .B(n23066), .Z(n23070) );
  XNOR U23281 ( .A(n23071), .B(n23070), .Z(n23073) );
  NAND U23282 ( .A(b[45]), .B(a[63]), .Z(n23072) );
  XOR U23283 ( .A(n23073), .B(n23072), .Z(n22970) );
  OR U23284 ( .A(n22945), .B(n22944), .Z(n22949) );
  NANDN U23285 ( .A(n22947), .B(n22946), .Z(n22948) );
  AND U23286 ( .A(n22949), .B(n22948), .Z(n22971) );
  XNOR U23287 ( .A(n22970), .B(n22971), .Z(n22965) );
  NOR U23288 ( .A(n22951), .B(n22950), .Z(n22964) );
  XOR U23289 ( .A(n22965), .B(n22964), .Z(n22967) );
  NOR U23290 ( .A(n22953), .B(n22952), .Z(n22958) );
  AND U23291 ( .A(n22955), .B(n22954), .Z(n22956) );
  OR U23292 ( .A(n22958), .B(n22956), .Z(n22957) );
  NAND U23293 ( .A(n22957), .B(n22959), .Z(n22963) );
  OR U23294 ( .A(n22959), .B(n22958), .Z(n22960) );
  NANDN U23295 ( .A(n22961), .B(n22960), .Z(n22962) );
  AND U23296 ( .A(n22963), .B(n22962), .Z(n22966) );
  XOR U23297 ( .A(n22967), .B(n22966), .Z(c[108]) );
  NANDN U23298 ( .A(n22965), .B(n22964), .Z(n22969) );
  OR U23299 ( .A(n22967), .B(n22966), .Z(n22968) );
  NAND U23300 ( .A(n22969), .B(n22968), .Z(n23183) );
  AND U23301 ( .A(n22971), .B(n22970), .Z(n23180) );
  AND U23302 ( .A(b[63]), .B(a[46]), .Z(n23105) );
  AND U23303 ( .A(b[62]), .B(a[47]), .Z(n23103) );
  OR U23304 ( .A(n22973), .B(n22972), .Z(n22977) );
  NANDN U23305 ( .A(n22975), .B(n22974), .Z(n22976) );
  AND U23306 ( .A(n22977), .B(n22976), .Z(n23102) );
  XNOR U23307 ( .A(n23103), .B(n23102), .Z(n23104) );
  XOR U23308 ( .A(n23105), .B(n23104), .Z(n23111) );
  NANDN U23309 ( .A(n22979), .B(n22978), .Z(n22983) );
  NANDN U23310 ( .A(n22981), .B(n22980), .Z(n22982) );
  NAND U23311 ( .A(n22983), .B(n22982), .Z(n23109) );
  NAND U23312 ( .A(b[61]), .B(a[48]), .Z(n23108) );
  XOR U23313 ( .A(n23109), .B(n23108), .Z(n23110) );
  XOR U23314 ( .A(n23111), .B(n23110), .Z(n23117) );
  AND U23315 ( .A(a[49]), .B(b[60]), .Z(n23114) );
  OR U23316 ( .A(n22985), .B(n22984), .Z(n22989) );
  NAND U23317 ( .A(n22987), .B(n22986), .Z(n22988) );
  NAND U23318 ( .A(n22989), .B(n22988), .Z(n23115) );
  XOR U23319 ( .A(n23114), .B(n23115), .Z(n23116) );
  XNOR U23320 ( .A(n23117), .B(n23116), .Z(n23099) );
  NAND U23321 ( .A(n22991), .B(n22990), .Z(n22995) );
  OR U23322 ( .A(n22993), .B(n22992), .Z(n22994) );
  NAND U23323 ( .A(n22995), .B(n22994), .Z(n23096) );
  NAND U23324 ( .A(a[50]), .B(b[59]), .Z(n23097) );
  XNOR U23325 ( .A(n23096), .B(n23097), .Z(n23098) );
  XNOR U23326 ( .A(n23099), .B(n23098), .Z(n23093) );
  AND U23327 ( .A(a[51]), .B(b[58]), .Z(n23090) );
  OR U23328 ( .A(n22997), .B(n22996), .Z(n23001) );
  NAND U23329 ( .A(n22999), .B(n22998), .Z(n23000) );
  NAND U23330 ( .A(n23001), .B(n23000), .Z(n23091) );
  XOR U23331 ( .A(n23090), .B(n23091), .Z(n23092) );
  XNOR U23332 ( .A(n23093), .B(n23092), .Z(n23123) );
  NAND U23333 ( .A(b[57]), .B(a[52]), .Z(n23120) );
  XOR U23334 ( .A(n23121), .B(n23120), .Z(n23122) );
  XNOR U23335 ( .A(n23123), .B(n23122), .Z(n23129) );
  AND U23336 ( .A(a[53]), .B(b[56]), .Z(n23126) );
  OR U23337 ( .A(n23007), .B(n23006), .Z(n23011) );
  NAND U23338 ( .A(n23009), .B(n23008), .Z(n23010) );
  NAND U23339 ( .A(n23011), .B(n23010), .Z(n23127) );
  XOR U23340 ( .A(n23126), .B(n23127), .Z(n23128) );
  XNOR U23341 ( .A(n23129), .B(n23128), .Z(n23087) );
  OR U23342 ( .A(n23013), .B(n23012), .Z(n23017) );
  NANDN U23343 ( .A(n23015), .B(n23014), .Z(n23016) );
  NAND U23344 ( .A(n23017), .B(n23016), .Z(n23085) );
  NAND U23345 ( .A(b[55]), .B(a[54]), .Z(n23084) );
  XOR U23346 ( .A(n23085), .B(n23084), .Z(n23086) );
  XNOR U23347 ( .A(n23087), .B(n23086), .Z(n23081) );
  AND U23348 ( .A(a[55]), .B(b[54]), .Z(n23078) );
  OR U23349 ( .A(n23019), .B(n23018), .Z(n23023) );
  NAND U23350 ( .A(n23021), .B(n23020), .Z(n23022) );
  NAND U23351 ( .A(n23023), .B(n23022), .Z(n23079) );
  XOR U23352 ( .A(n23078), .B(n23079), .Z(n23080) );
  XNOR U23353 ( .A(n23081), .B(n23080), .Z(n23135) );
  NAND U23354 ( .A(n23025), .B(n23024), .Z(n23029) );
  OR U23355 ( .A(n23027), .B(n23026), .Z(n23028) );
  NAND U23356 ( .A(n23029), .B(n23028), .Z(n23132) );
  NAND U23357 ( .A(a[56]), .B(b[53]), .Z(n23133) );
  XNOR U23358 ( .A(n23132), .B(n23133), .Z(n23134) );
  XNOR U23359 ( .A(n23135), .B(n23134), .Z(n23141) );
  AND U23360 ( .A(a[57]), .B(b[52]), .Z(n23138) );
  OR U23361 ( .A(n23031), .B(n23030), .Z(n23035) );
  NAND U23362 ( .A(n23033), .B(n23032), .Z(n23034) );
  NAND U23363 ( .A(n23035), .B(n23034), .Z(n23139) );
  XOR U23364 ( .A(n23138), .B(n23139), .Z(n23140) );
  XNOR U23365 ( .A(n23141), .B(n23140), .Z(n23147) );
  NAND U23366 ( .A(n23037), .B(n23036), .Z(n23041) );
  OR U23367 ( .A(n23039), .B(n23038), .Z(n23040) );
  NAND U23368 ( .A(n23041), .B(n23040), .Z(n23144) );
  NAND U23369 ( .A(a[58]), .B(b[51]), .Z(n23145) );
  XNOR U23370 ( .A(n23144), .B(n23145), .Z(n23146) );
  XNOR U23371 ( .A(n23147), .B(n23146), .Z(n23153) );
  AND U23372 ( .A(a[59]), .B(b[50]), .Z(n23150) );
  OR U23373 ( .A(n23043), .B(n23042), .Z(n23047) );
  NAND U23374 ( .A(n23045), .B(n23044), .Z(n23046) );
  NAND U23375 ( .A(n23047), .B(n23046), .Z(n23151) );
  XOR U23376 ( .A(n23150), .B(n23151), .Z(n23152) );
  XNOR U23377 ( .A(n23153), .B(n23152), .Z(n23159) );
  NAND U23378 ( .A(n23049), .B(n23048), .Z(n23053) );
  OR U23379 ( .A(n23051), .B(n23050), .Z(n23052) );
  NAND U23380 ( .A(n23053), .B(n23052), .Z(n23156) );
  NAND U23381 ( .A(a[60]), .B(b[49]), .Z(n23157) );
  XNOR U23382 ( .A(n23156), .B(n23157), .Z(n23158) );
  XNOR U23383 ( .A(n23159), .B(n23158), .Z(n23165) );
  AND U23384 ( .A(a[61]), .B(b[48]), .Z(n23162) );
  OR U23385 ( .A(n23055), .B(n23054), .Z(n23059) );
  NAND U23386 ( .A(n23057), .B(n23056), .Z(n23058) );
  NAND U23387 ( .A(n23059), .B(n23058), .Z(n23163) );
  XOR U23388 ( .A(n23162), .B(n23163), .Z(n23164) );
  XNOR U23389 ( .A(n23165), .B(n23164), .Z(n23171) );
  NAND U23390 ( .A(b[47]), .B(a[62]), .Z(n23168) );
  XOR U23391 ( .A(n23169), .B(n23168), .Z(n23170) );
  XNOR U23392 ( .A(n23171), .B(n23170), .Z(n23177) );
  AND U23393 ( .A(a[63]), .B(b[46]), .Z(n23174) );
  OR U23394 ( .A(n23065), .B(n23064), .Z(n23069) );
  NAND U23395 ( .A(n23067), .B(n23066), .Z(n23068) );
  NAND U23396 ( .A(n23069), .B(n23068), .Z(n23175) );
  XOR U23397 ( .A(n23174), .B(n23175), .Z(n23176) );
  XNOR U23398 ( .A(n23177), .B(n23176), .Z(n23076) );
  NAND U23399 ( .A(n23071), .B(n23070), .Z(n23075) );
  OR U23400 ( .A(n23073), .B(n23072), .Z(n23074) );
  NAND U23401 ( .A(n23075), .B(n23074), .Z(n23077) );
  XNOR U23402 ( .A(n23076), .B(n23077), .Z(n23181) );
  XOR U23403 ( .A(n23180), .B(n23181), .Z(n23182) );
  XOR U23404 ( .A(n23183), .B(n23182), .Z(c[109]) );
  ANDN U23405 ( .B(n23077), .A(n23076), .Z(n23278) );
  AND U23406 ( .A(a[63]), .B(b[47]), .Z(n23275) );
  AND U23407 ( .A(a[61]), .B(b[49]), .Z(n23263) );
  AND U23408 ( .A(a[59]), .B(b[51]), .Z(n23251) );
  AND U23409 ( .A(a[57]), .B(b[53]), .Z(n23241) );
  OR U23410 ( .A(n23079), .B(n23078), .Z(n23083) );
  NANDN U23411 ( .A(n23081), .B(n23080), .Z(n23082) );
  NAND U23412 ( .A(n23083), .B(n23082), .Z(n23233) );
  NAND U23413 ( .A(b[54]), .B(a[56]), .Z(n23232) );
  XOR U23414 ( .A(n23233), .B(n23232), .Z(n23234) );
  OR U23415 ( .A(n23085), .B(n23084), .Z(n23089) );
  NANDN U23416 ( .A(n23087), .B(n23086), .Z(n23088) );
  NAND U23417 ( .A(n23089), .B(n23088), .Z(n23227) );
  AND U23418 ( .A(a[53]), .B(b[57]), .Z(n23219) );
  OR U23419 ( .A(n23091), .B(n23090), .Z(n23095) );
  NANDN U23420 ( .A(n23093), .B(n23092), .Z(n23094) );
  NAND U23421 ( .A(n23095), .B(n23094), .Z(n23211) );
  NAND U23422 ( .A(b[58]), .B(a[52]), .Z(n23210) );
  XOR U23423 ( .A(n23211), .B(n23210), .Z(n23212) );
  NANDN U23424 ( .A(n23097), .B(n23096), .Z(n23101) );
  NANDN U23425 ( .A(n23099), .B(n23098), .Z(n23100) );
  NAND U23426 ( .A(n23101), .B(n23100), .Z(n23205) );
  AND U23427 ( .A(a[49]), .B(b[61]), .Z(n23195) );
  NANDN U23428 ( .A(n23103), .B(n23102), .Z(n23107) );
  NANDN U23429 ( .A(n23105), .B(n23104), .Z(n23106) );
  NAND U23430 ( .A(n23107), .B(n23106), .Z(n23187) );
  NAND U23431 ( .A(a[48]), .B(b[62]), .Z(n23186) );
  XOR U23432 ( .A(n23187), .B(n23186), .Z(n23188) );
  NAND U23433 ( .A(a[47]), .B(b[63]), .Z(n23189) );
  XOR U23434 ( .A(n23188), .B(n23189), .Z(n23192) );
  OR U23435 ( .A(n23109), .B(n23108), .Z(n23113) );
  NAND U23436 ( .A(n23111), .B(n23110), .Z(n23112) );
  NAND U23437 ( .A(n23113), .B(n23112), .Z(n23193) );
  XNOR U23438 ( .A(n23192), .B(n23193), .Z(n23194) );
  XOR U23439 ( .A(n23195), .B(n23194), .Z(n23201) );
  OR U23440 ( .A(n23115), .B(n23114), .Z(n23119) );
  NANDN U23441 ( .A(n23117), .B(n23116), .Z(n23118) );
  NAND U23442 ( .A(n23119), .B(n23118), .Z(n23199) );
  NAND U23443 ( .A(b[60]), .B(a[50]), .Z(n23198) );
  XOR U23444 ( .A(n23199), .B(n23198), .Z(n23200) );
  XOR U23445 ( .A(n23201), .B(n23200), .Z(n23204) );
  XNOR U23446 ( .A(n23205), .B(n23204), .Z(n23207) );
  NAND U23447 ( .A(b[59]), .B(a[51]), .Z(n23206) );
  XOR U23448 ( .A(n23207), .B(n23206), .Z(n23213) );
  XOR U23449 ( .A(n23212), .B(n23213), .Z(n23216) );
  OR U23450 ( .A(n23121), .B(n23120), .Z(n23125) );
  NANDN U23451 ( .A(n23123), .B(n23122), .Z(n23124) );
  NAND U23452 ( .A(n23125), .B(n23124), .Z(n23217) );
  XOR U23453 ( .A(n23216), .B(n23217), .Z(n23218) );
  XOR U23454 ( .A(n23219), .B(n23218), .Z(n23223) );
  OR U23455 ( .A(n23127), .B(n23126), .Z(n23131) );
  NANDN U23456 ( .A(n23129), .B(n23128), .Z(n23130) );
  NAND U23457 ( .A(n23131), .B(n23130), .Z(n23221) );
  NAND U23458 ( .A(b[56]), .B(a[54]), .Z(n23220) );
  XOR U23459 ( .A(n23221), .B(n23220), .Z(n23222) );
  XOR U23460 ( .A(n23223), .B(n23222), .Z(n23226) );
  XNOR U23461 ( .A(n23227), .B(n23226), .Z(n23229) );
  NAND U23462 ( .A(b[55]), .B(a[55]), .Z(n23228) );
  XOR U23463 ( .A(n23229), .B(n23228), .Z(n23235) );
  XOR U23464 ( .A(n23234), .B(n23235), .Z(n23238) );
  NANDN U23465 ( .A(n23133), .B(n23132), .Z(n23137) );
  NANDN U23466 ( .A(n23135), .B(n23134), .Z(n23136) );
  NAND U23467 ( .A(n23137), .B(n23136), .Z(n23239) );
  XOR U23468 ( .A(n23238), .B(n23239), .Z(n23240) );
  XOR U23469 ( .A(n23241), .B(n23240), .Z(n23245) );
  OR U23470 ( .A(n23139), .B(n23138), .Z(n23143) );
  NANDN U23471 ( .A(n23141), .B(n23140), .Z(n23142) );
  NAND U23472 ( .A(n23143), .B(n23142), .Z(n23243) );
  NAND U23473 ( .A(b[52]), .B(a[58]), .Z(n23242) );
  XOR U23474 ( .A(n23243), .B(n23242), .Z(n23244) );
  XOR U23475 ( .A(n23245), .B(n23244), .Z(n23248) );
  NANDN U23476 ( .A(n23145), .B(n23144), .Z(n23149) );
  NANDN U23477 ( .A(n23147), .B(n23146), .Z(n23148) );
  NAND U23478 ( .A(n23149), .B(n23148), .Z(n23249) );
  XOR U23479 ( .A(n23248), .B(n23249), .Z(n23250) );
  XOR U23480 ( .A(n23251), .B(n23250), .Z(n23257) );
  OR U23481 ( .A(n23151), .B(n23150), .Z(n23155) );
  NANDN U23482 ( .A(n23153), .B(n23152), .Z(n23154) );
  NAND U23483 ( .A(n23155), .B(n23154), .Z(n23255) );
  NAND U23484 ( .A(b[50]), .B(a[60]), .Z(n23254) );
  XOR U23485 ( .A(n23255), .B(n23254), .Z(n23256) );
  XOR U23486 ( .A(n23257), .B(n23256), .Z(n23260) );
  NANDN U23487 ( .A(n23157), .B(n23156), .Z(n23161) );
  NANDN U23488 ( .A(n23159), .B(n23158), .Z(n23160) );
  NAND U23489 ( .A(n23161), .B(n23160), .Z(n23261) );
  XOR U23490 ( .A(n23260), .B(n23261), .Z(n23262) );
  XOR U23491 ( .A(n23263), .B(n23262), .Z(n23269) );
  OR U23492 ( .A(n23163), .B(n23162), .Z(n23167) );
  NANDN U23493 ( .A(n23165), .B(n23164), .Z(n23166) );
  NAND U23494 ( .A(n23167), .B(n23166), .Z(n23267) );
  NAND U23495 ( .A(b[48]), .B(a[62]), .Z(n23266) );
  XOR U23496 ( .A(n23267), .B(n23266), .Z(n23268) );
  XOR U23497 ( .A(n23269), .B(n23268), .Z(n23272) );
  OR U23498 ( .A(n23169), .B(n23168), .Z(n23173) );
  NANDN U23499 ( .A(n23171), .B(n23170), .Z(n23172) );
  NAND U23500 ( .A(n23173), .B(n23172), .Z(n23273) );
  XOR U23501 ( .A(n23272), .B(n23273), .Z(n23274) );
  XOR U23502 ( .A(n23275), .B(n23274), .Z(n23184) );
  OR U23503 ( .A(n23175), .B(n23174), .Z(n23179) );
  NANDN U23504 ( .A(n23177), .B(n23176), .Z(n23178) );
  AND U23505 ( .A(n23179), .B(n23178), .Z(n23185) );
  XOR U23506 ( .A(n23184), .B(n23185), .Z(n23279) );
  XOR U23507 ( .A(n23278), .B(n23279), .Z(n23280) );
  XOR U23508 ( .A(n23280), .B(n23281), .Z(c[110]) );
  AND U23509 ( .A(n23185), .B(n23184), .Z(n23374) );
  AND U23510 ( .A(b[63]), .B(a[48]), .Z(n23323) );
  AND U23511 ( .A(b[62]), .B(a[49]), .Z(n23321) );
  OR U23512 ( .A(n23187), .B(n23186), .Z(n23191) );
  NANDN U23513 ( .A(n23189), .B(n23188), .Z(n23190) );
  AND U23514 ( .A(n23191), .B(n23190), .Z(n23320) );
  XNOR U23515 ( .A(n23321), .B(n23320), .Z(n23322) );
  XOR U23516 ( .A(n23323), .B(n23322), .Z(n23329) );
  NANDN U23517 ( .A(n23193), .B(n23192), .Z(n23197) );
  NANDN U23518 ( .A(n23195), .B(n23194), .Z(n23196) );
  NAND U23519 ( .A(n23197), .B(n23196), .Z(n23327) );
  NAND U23520 ( .A(b[61]), .B(a[50]), .Z(n23326) );
  XOR U23521 ( .A(n23327), .B(n23326), .Z(n23328) );
  XOR U23522 ( .A(n23329), .B(n23328), .Z(n23335) );
  AND U23523 ( .A(a[51]), .B(b[60]), .Z(n23332) );
  OR U23524 ( .A(n23199), .B(n23198), .Z(n23203) );
  NAND U23525 ( .A(n23201), .B(n23200), .Z(n23202) );
  NAND U23526 ( .A(n23203), .B(n23202), .Z(n23333) );
  XOR U23527 ( .A(n23332), .B(n23333), .Z(n23334) );
  XNOR U23528 ( .A(n23335), .B(n23334), .Z(n23317) );
  NAND U23529 ( .A(n23205), .B(n23204), .Z(n23209) );
  OR U23530 ( .A(n23207), .B(n23206), .Z(n23208) );
  NAND U23531 ( .A(n23209), .B(n23208), .Z(n23314) );
  NAND U23532 ( .A(a[52]), .B(b[59]), .Z(n23315) );
  XNOR U23533 ( .A(n23314), .B(n23315), .Z(n23316) );
  XNOR U23534 ( .A(n23317), .B(n23316), .Z(n23311) );
  AND U23535 ( .A(a[53]), .B(b[58]), .Z(n23308) );
  OR U23536 ( .A(n23211), .B(n23210), .Z(n23215) );
  NAND U23537 ( .A(n23213), .B(n23212), .Z(n23214) );
  NAND U23538 ( .A(n23215), .B(n23214), .Z(n23309) );
  XOR U23539 ( .A(n23308), .B(n23309), .Z(n23310) );
  XNOR U23540 ( .A(n23311), .B(n23310), .Z(n23341) );
  NAND U23541 ( .A(b[57]), .B(a[54]), .Z(n23338) );
  XOR U23542 ( .A(n23339), .B(n23338), .Z(n23340) );
  XNOR U23543 ( .A(n23341), .B(n23340), .Z(n23347) );
  AND U23544 ( .A(a[55]), .B(b[56]), .Z(n23344) );
  OR U23545 ( .A(n23221), .B(n23220), .Z(n23225) );
  NAND U23546 ( .A(n23223), .B(n23222), .Z(n23224) );
  NAND U23547 ( .A(n23225), .B(n23224), .Z(n23345) );
  XOR U23548 ( .A(n23344), .B(n23345), .Z(n23346) );
  XNOR U23549 ( .A(n23347), .B(n23346), .Z(n23353) );
  NAND U23550 ( .A(n23227), .B(n23226), .Z(n23231) );
  OR U23551 ( .A(n23229), .B(n23228), .Z(n23230) );
  NAND U23552 ( .A(n23231), .B(n23230), .Z(n23350) );
  NAND U23553 ( .A(a[56]), .B(b[55]), .Z(n23351) );
  XNOR U23554 ( .A(n23350), .B(n23351), .Z(n23352) );
  XNOR U23555 ( .A(n23353), .B(n23352), .Z(n23359) );
  AND U23556 ( .A(a[57]), .B(b[54]), .Z(n23356) );
  OR U23557 ( .A(n23233), .B(n23232), .Z(n23237) );
  NAND U23558 ( .A(n23235), .B(n23234), .Z(n23236) );
  NAND U23559 ( .A(n23237), .B(n23236), .Z(n23357) );
  XOR U23560 ( .A(n23356), .B(n23357), .Z(n23358) );
  XNOR U23561 ( .A(n23359), .B(n23358), .Z(n23305) );
  NAND U23562 ( .A(b[53]), .B(a[58]), .Z(n23302) );
  XOR U23563 ( .A(n23303), .B(n23302), .Z(n23304) );
  XNOR U23564 ( .A(n23305), .B(n23304), .Z(n23299) );
  AND U23565 ( .A(a[59]), .B(b[52]), .Z(n23296) );
  OR U23566 ( .A(n23243), .B(n23242), .Z(n23247) );
  NAND U23567 ( .A(n23245), .B(n23244), .Z(n23246) );
  NAND U23568 ( .A(n23247), .B(n23246), .Z(n23297) );
  XOR U23569 ( .A(n23296), .B(n23297), .Z(n23298) );
  XNOR U23570 ( .A(n23299), .B(n23298), .Z(n23293) );
  OR U23571 ( .A(n23249), .B(n23248), .Z(n23253) );
  NANDN U23572 ( .A(n23251), .B(n23250), .Z(n23252) );
  NAND U23573 ( .A(n23253), .B(n23252), .Z(n23291) );
  NAND U23574 ( .A(b[51]), .B(a[60]), .Z(n23290) );
  XOR U23575 ( .A(n23291), .B(n23290), .Z(n23292) );
  XNOR U23576 ( .A(n23293), .B(n23292), .Z(n23287) );
  AND U23577 ( .A(a[61]), .B(b[50]), .Z(n23284) );
  OR U23578 ( .A(n23255), .B(n23254), .Z(n23259) );
  NAND U23579 ( .A(n23257), .B(n23256), .Z(n23258) );
  NAND U23580 ( .A(n23259), .B(n23258), .Z(n23285) );
  XOR U23581 ( .A(n23284), .B(n23285), .Z(n23286) );
  XNOR U23582 ( .A(n23287), .B(n23286), .Z(n23365) );
  OR U23583 ( .A(n23261), .B(n23260), .Z(n23265) );
  NANDN U23584 ( .A(n23263), .B(n23262), .Z(n23264) );
  NAND U23585 ( .A(n23265), .B(n23264), .Z(n23363) );
  NAND U23586 ( .A(b[49]), .B(a[62]), .Z(n23362) );
  XOR U23587 ( .A(n23363), .B(n23362), .Z(n23364) );
  XNOR U23588 ( .A(n23365), .B(n23364), .Z(n23371) );
  AND U23589 ( .A(a[63]), .B(b[48]), .Z(n23368) );
  OR U23590 ( .A(n23267), .B(n23266), .Z(n23271) );
  NAND U23591 ( .A(n23269), .B(n23268), .Z(n23270) );
  NAND U23592 ( .A(n23271), .B(n23270), .Z(n23369) );
  XOR U23593 ( .A(n23368), .B(n23369), .Z(n23370) );
  XNOR U23594 ( .A(n23371), .B(n23370), .Z(n23282) );
  OR U23595 ( .A(n23273), .B(n23272), .Z(n23277) );
  NANDN U23596 ( .A(n23275), .B(n23274), .Z(n23276) );
  AND U23597 ( .A(n23277), .B(n23276), .Z(n23283) );
  XNOR U23598 ( .A(n23282), .B(n23283), .Z(n23375) );
  XOR U23599 ( .A(n23374), .B(n23375), .Z(n23376) );
  XOR U23600 ( .A(n23376), .B(n23377), .Z(c[111]) );
  ANDN U23601 ( .B(n23283), .A(n23282), .Z(n23460) );
  AND U23602 ( .A(a[63]), .B(b[49]), .Z(n23459) );
  OR U23603 ( .A(n23285), .B(n23284), .Z(n23289) );
  NANDN U23604 ( .A(n23287), .B(n23286), .Z(n23288) );
  NAND U23605 ( .A(n23289), .B(n23288), .Z(n23451) );
  NAND U23606 ( .A(b[50]), .B(a[62]), .Z(n23450) );
  XOR U23607 ( .A(n23451), .B(n23450), .Z(n23452) );
  OR U23608 ( .A(n23291), .B(n23290), .Z(n23295) );
  NANDN U23609 ( .A(n23293), .B(n23292), .Z(n23294) );
  NAND U23610 ( .A(n23295), .B(n23294), .Z(n23445) );
  OR U23611 ( .A(n23297), .B(n23296), .Z(n23301) );
  NANDN U23612 ( .A(n23299), .B(n23298), .Z(n23300) );
  NAND U23613 ( .A(n23301), .B(n23300), .Z(n23439) );
  NAND U23614 ( .A(b[52]), .B(a[60]), .Z(n23438) );
  XOR U23615 ( .A(n23439), .B(n23438), .Z(n23440) );
  OR U23616 ( .A(n23303), .B(n23302), .Z(n23307) );
  NANDN U23617 ( .A(n23305), .B(n23304), .Z(n23306) );
  NAND U23618 ( .A(n23307), .B(n23306), .Z(n23433) );
  AND U23619 ( .A(a[57]), .B(b[55]), .Z(n23423) );
  AND U23620 ( .A(a[55]), .B(b[57]), .Z(n23413) );
  OR U23621 ( .A(n23309), .B(n23308), .Z(n23313) );
  NANDN U23622 ( .A(n23311), .B(n23310), .Z(n23312) );
  NAND U23623 ( .A(n23313), .B(n23312), .Z(n23405) );
  NAND U23624 ( .A(b[58]), .B(a[54]), .Z(n23404) );
  XOR U23625 ( .A(n23405), .B(n23404), .Z(n23406) );
  NANDN U23626 ( .A(n23315), .B(n23314), .Z(n23319) );
  NANDN U23627 ( .A(n23317), .B(n23316), .Z(n23318) );
  NAND U23628 ( .A(n23319), .B(n23318), .Z(n23399) );
  AND U23629 ( .A(a[51]), .B(b[61]), .Z(n23389) );
  NANDN U23630 ( .A(n23321), .B(n23320), .Z(n23325) );
  NANDN U23631 ( .A(n23323), .B(n23322), .Z(n23324) );
  NAND U23632 ( .A(n23325), .B(n23324), .Z(n23381) );
  NAND U23633 ( .A(a[50]), .B(b[62]), .Z(n23380) );
  XOR U23634 ( .A(n23381), .B(n23380), .Z(n23382) );
  NAND U23635 ( .A(a[49]), .B(b[63]), .Z(n23383) );
  XOR U23636 ( .A(n23382), .B(n23383), .Z(n23386) );
  OR U23637 ( .A(n23327), .B(n23326), .Z(n23331) );
  NAND U23638 ( .A(n23329), .B(n23328), .Z(n23330) );
  NAND U23639 ( .A(n23331), .B(n23330), .Z(n23387) );
  XNOR U23640 ( .A(n23386), .B(n23387), .Z(n23388) );
  XOR U23641 ( .A(n23389), .B(n23388), .Z(n23395) );
  OR U23642 ( .A(n23333), .B(n23332), .Z(n23337) );
  NANDN U23643 ( .A(n23335), .B(n23334), .Z(n23336) );
  NAND U23644 ( .A(n23337), .B(n23336), .Z(n23393) );
  NAND U23645 ( .A(b[60]), .B(a[52]), .Z(n23392) );
  XOR U23646 ( .A(n23393), .B(n23392), .Z(n23394) );
  XOR U23647 ( .A(n23395), .B(n23394), .Z(n23398) );
  XNOR U23648 ( .A(n23399), .B(n23398), .Z(n23401) );
  NAND U23649 ( .A(b[59]), .B(a[53]), .Z(n23400) );
  XOR U23650 ( .A(n23401), .B(n23400), .Z(n23407) );
  XOR U23651 ( .A(n23406), .B(n23407), .Z(n23410) );
  OR U23652 ( .A(n23339), .B(n23338), .Z(n23343) );
  NANDN U23653 ( .A(n23341), .B(n23340), .Z(n23342) );
  NAND U23654 ( .A(n23343), .B(n23342), .Z(n23411) );
  XOR U23655 ( .A(n23410), .B(n23411), .Z(n23412) );
  XOR U23656 ( .A(n23413), .B(n23412), .Z(n23417) );
  OR U23657 ( .A(n23345), .B(n23344), .Z(n23349) );
  NANDN U23658 ( .A(n23347), .B(n23346), .Z(n23348) );
  NAND U23659 ( .A(n23349), .B(n23348), .Z(n23415) );
  NAND U23660 ( .A(b[56]), .B(a[56]), .Z(n23414) );
  XOR U23661 ( .A(n23415), .B(n23414), .Z(n23416) );
  XOR U23662 ( .A(n23417), .B(n23416), .Z(n23420) );
  NANDN U23663 ( .A(n23351), .B(n23350), .Z(n23355) );
  NANDN U23664 ( .A(n23353), .B(n23352), .Z(n23354) );
  NAND U23665 ( .A(n23355), .B(n23354), .Z(n23421) );
  XOR U23666 ( .A(n23420), .B(n23421), .Z(n23422) );
  XOR U23667 ( .A(n23423), .B(n23422), .Z(n23429) );
  OR U23668 ( .A(n23357), .B(n23356), .Z(n23361) );
  NANDN U23669 ( .A(n23359), .B(n23358), .Z(n23360) );
  NAND U23670 ( .A(n23361), .B(n23360), .Z(n23427) );
  NAND U23671 ( .A(b[54]), .B(a[58]), .Z(n23426) );
  XOR U23672 ( .A(n23427), .B(n23426), .Z(n23428) );
  XOR U23673 ( .A(n23429), .B(n23428), .Z(n23432) );
  XNOR U23674 ( .A(n23433), .B(n23432), .Z(n23435) );
  NAND U23675 ( .A(b[53]), .B(a[59]), .Z(n23434) );
  XOR U23676 ( .A(n23435), .B(n23434), .Z(n23441) );
  XOR U23677 ( .A(n23440), .B(n23441), .Z(n23444) );
  XNOR U23678 ( .A(n23445), .B(n23444), .Z(n23447) );
  NAND U23679 ( .A(b[51]), .B(a[61]), .Z(n23446) );
  XOR U23680 ( .A(n23447), .B(n23446), .Z(n23453) );
  XOR U23681 ( .A(n23452), .B(n23453), .Z(n23456) );
  OR U23682 ( .A(n23363), .B(n23362), .Z(n23367) );
  NANDN U23683 ( .A(n23365), .B(n23364), .Z(n23366) );
  NAND U23684 ( .A(n23367), .B(n23366), .Z(n23457) );
  XOR U23685 ( .A(n23456), .B(n23457), .Z(n23458) );
  XOR U23686 ( .A(n23459), .B(n23458), .Z(n23378) );
  OR U23687 ( .A(n23369), .B(n23368), .Z(n23373) );
  NANDN U23688 ( .A(n23371), .B(n23370), .Z(n23372) );
  AND U23689 ( .A(n23373), .B(n23372), .Z(n23379) );
  XOR U23690 ( .A(n23378), .B(n23379), .Z(n23461) );
  XOR U23691 ( .A(n23460), .B(n23461), .Z(n23462) );
  XOR U23692 ( .A(n23462), .B(n23463), .Z(c[112]) );
  AND U23693 ( .A(n23379), .B(n23378), .Z(n23544) );
  AND U23694 ( .A(b[63]), .B(a[50]), .Z(n23493) );
  AND U23695 ( .A(b[62]), .B(a[51]), .Z(n23491) );
  OR U23696 ( .A(n23381), .B(n23380), .Z(n23385) );
  NANDN U23697 ( .A(n23383), .B(n23382), .Z(n23384) );
  AND U23698 ( .A(n23385), .B(n23384), .Z(n23490) );
  XNOR U23699 ( .A(n23491), .B(n23490), .Z(n23492) );
  XOR U23700 ( .A(n23493), .B(n23492), .Z(n23499) );
  NANDN U23701 ( .A(n23387), .B(n23386), .Z(n23391) );
  NANDN U23702 ( .A(n23389), .B(n23388), .Z(n23390) );
  NAND U23703 ( .A(n23391), .B(n23390), .Z(n23497) );
  NAND U23704 ( .A(b[61]), .B(a[52]), .Z(n23496) );
  XOR U23705 ( .A(n23497), .B(n23496), .Z(n23498) );
  XOR U23706 ( .A(n23499), .B(n23498), .Z(n23505) );
  AND U23707 ( .A(a[53]), .B(b[60]), .Z(n23502) );
  OR U23708 ( .A(n23393), .B(n23392), .Z(n23397) );
  NAND U23709 ( .A(n23395), .B(n23394), .Z(n23396) );
  NAND U23710 ( .A(n23397), .B(n23396), .Z(n23503) );
  XOR U23711 ( .A(n23502), .B(n23503), .Z(n23504) );
  XNOR U23712 ( .A(n23505), .B(n23504), .Z(n23487) );
  NAND U23713 ( .A(n23399), .B(n23398), .Z(n23403) );
  OR U23714 ( .A(n23401), .B(n23400), .Z(n23402) );
  NAND U23715 ( .A(n23403), .B(n23402), .Z(n23484) );
  NAND U23716 ( .A(a[54]), .B(b[59]), .Z(n23485) );
  XNOR U23717 ( .A(n23484), .B(n23485), .Z(n23486) );
  XNOR U23718 ( .A(n23487), .B(n23486), .Z(n23481) );
  AND U23719 ( .A(a[55]), .B(b[58]), .Z(n23478) );
  OR U23720 ( .A(n23405), .B(n23404), .Z(n23409) );
  NAND U23721 ( .A(n23407), .B(n23406), .Z(n23408) );
  NAND U23722 ( .A(n23409), .B(n23408), .Z(n23479) );
  XOR U23723 ( .A(n23478), .B(n23479), .Z(n23480) );
  XNOR U23724 ( .A(n23481), .B(n23480), .Z(n23511) );
  NAND U23725 ( .A(b[57]), .B(a[56]), .Z(n23508) );
  XOR U23726 ( .A(n23509), .B(n23508), .Z(n23510) );
  XNOR U23727 ( .A(n23511), .B(n23510), .Z(n23517) );
  AND U23728 ( .A(a[57]), .B(b[56]), .Z(n23514) );
  OR U23729 ( .A(n23415), .B(n23414), .Z(n23419) );
  NAND U23730 ( .A(n23417), .B(n23416), .Z(n23418) );
  NAND U23731 ( .A(n23419), .B(n23418), .Z(n23515) );
  XOR U23732 ( .A(n23514), .B(n23515), .Z(n23516) );
  XNOR U23733 ( .A(n23517), .B(n23516), .Z(n23475) );
  OR U23734 ( .A(n23421), .B(n23420), .Z(n23425) );
  NANDN U23735 ( .A(n23423), .B(n23422), .Z(n23424) );
  NAND U23736 ( .A(n23425), .B(n23424), .Z(n23473) );
  NAND U23737 ( .A(b[55]), .B(a[58]), .Z(n23472) );
  XOR U23738 ( .A(n23473), .B(n23472), .Z(n23474) );
  XNOR U23739 ( .A(n23475), .B(n23474), .Z(n23469) );
  AND U23740 ( .A(a[59]), .B(b[54]), .Z(n23466) );
  OR U23741 ( .A(n23427), .B(n23426), .Z(n23431) );
  NAND U23742 ( .A(n23429), .B(n23428), .Z(n23430) );
  NAND U23743 ( .A(n23431), .B(n23430), .Z(n23467) );
  XOR U23744 ( .A(n23466), .B(n23467), .Z(n23468) );
  XNOR U23745 ( .A(n23469), .B(n23468), .Z(n23523) );
  NAND U23746 ( .A(n23433), .B(n23432), .Z(n23437) );
  OR U23747 ( .A(n23435), .B(n23434), .Z(n23436) );
  NAND U23748 ( .A(n23437), .B(n23436), .Z(n23520) );
  NAND U23749 ( .A(a[60]), .B(b[53]), .Z(n23521) );
  XNOR U23750 ( .A(n23520), .B(n23521), .Z(n23522) );
  XNOR U23751 ( .A(n23523), .B(n23522), .Z(n23529) );
  AND U23752 ( .A(a[61]), .B(b[52]), .Z(n23526) );
  OR U23753 ( .A(n23439), .B(n23438), .Z(n23443) );
  NAND U23754 ( .A(n23441), .B(n23440), .Z(n23442) );
  NAND U23755 ( .A(n23443), .B(n23442), .Z(n23527) );
  XOR U23756 ( .A(n23526), .B(n23527), .Z(n23528) );
  XNOR U23757 ( .A(n23529), .B(n23528), .Z(n23535) );
  NAND U23758 ( .A(n23445), .B(n23444), .Z(n23449) );
  OR U23759 ( .A(n23447), .B(n23446), .Z(n23448) );
  NAND U23760 ( .A(n23449), .B(n23448), .Z(n23532) );
  NAND U23761 ( .A(a[62]), .B(b[51]), .Z(n23533) );
  XNOR U23762 ( .A(n23532), .B(n23533), .Z(n23534) );
  XNOR U23763 ( .A(n23535), .B(n23534), .Z(n23541) );
  AND U23764 ( .A(a[63]), .B(b[50]), .Z(n23538) );
  OR U23765 ( .A(n23451), .B(n23450), .Z(n23455) );
  NAND U23766 ( .A(n23453), .B(n23452), .Z(n23454) );
  NAND U23767 ( .A(n23455), .B(n23454), .Z(n23539) );
  XOR U23768 ( .A(n23538), .B(n23539), .Z(n23540) );
  XNOR U23769 ( .A(n23541), .B(n23540), .Z(n23464) );
  XNOR U23770 ( .A(n23464), .B(n23465), .Z(n23545) );
  XOR U23771 ( .A(n23544), .B(n23545), .Z(n23546) );
  XOR U23772 ( .A(n23546), .B(n23547), .Z(c[113]) );
  ANDN U23773 ( .B(n23465), .A(n23464), .Z(n23618) );
  AND U23774 ( .A(a[63]), .B(b[51]), .Z(n23615) );
  AND U23775 ( .A(a[61]), .B(b[53]), .Z(n23605) );
  OR U23776 ( .A(n23467), .B(n23466), .Z(n23471) );
  NANDN U23777 ( .A(n23469), .B(n23468), .Z(n23470) );
  NAND U23778 ( .A(n23471), .B(n23470), .Z(n23597) );
  NAND U23779 ( .A(b[54]), .B(a[60]), .Z(n23596) );
  XOR U23780 ( .A(n23597), .B(n23596), .Z(n23598) );
  OR U23781 ( .A(n23473), .B(n23472), .Z(n23477) );
  NANDN U23782 ( .A(n23475), .B(n23474), .Z(n23476) );
  NAND U23783 ( .A(n23477), .B(n23476), .Z(n23591) );
  AND U23784 ( .A(a[57]), .B(b[57]), .Z(n23583) );
  OR U23785 ( .A(n23479), .B(n23478), .Z(n23483) );
  NANDN U23786 ( .A(n23481), .B(n23480), .Z(n23482) );
  NAND U23787 ( .A(n23483), .B(n23482), .Z(n23575) );
  NAND U23788 ( .A(b[58]), .B(a[56]), .Z(n23574) );
  XOR U23789 ( .A(n23575), .B(n23574), .Z(n23576) );
  NANDN U23790 ( .A(n23485), .B(n23484), .Z(n23489) );
  NANDN U23791 ( .A(n23487), .B(n23486), .Z(n23488) );
  NAND U23792 ( .A(n23489), .B(n23488), .Z(n23569) );
  AND U23793 ( .A(a[53]), .B(b[61]), .Z(n23559) );
  NANDN U23794 ( .A(n23491), .B(n23490), .Z(n23495) );
  NANDN U23795 ( .A(n23493), .B(n23492), .Z(n23494) );
  NAND U23796 ( .A(n23495), .B(n23494), .Z(n23551) );
  NAND U23797 ( .A(a[52]), .B(b[62]), .Z(n23550) );
  XOR U23798 ( .A(n23551), .B(n23550), .Z(n23552) );
  NAND U23799 ( .A(a[51]), .B(b[63]), .Z(n23553) );
  XOR U23800 ( .A(n23552), .B(n23553), .Z(n23556) );
  OR U23801 ( .A(n23497), .B(n23496), .Z(n23501) );
  NAND U23802 ( .A(n23499), .B(n23498), .Z(n23500) );
  NAND U23803 ( .A(n23501), .B(n23500), .Z(n23557) );
  XNOR U23804 ( .A(n23556), .B(n23557), .Z(n23558) );
  XOR U23805 ( .A(n23559), .B(n23558), .Z(n23565) );
  OR U23806 ( .A(n23503), .B(n23502), .Z(n23507) );
  NANDN U23807 ( .A(n23505), .B(n23504), .Z(n23506) );
  NAND U23808 ( .A(n23507), .B(n23506), .Z(n23563) );
  NAND U23809 ( .A(b[60]), .B(a[54]), .Z(n23562) );
  XOR U23810 ( .A(n23563), .B(n23562), .Z(n23564) );
  XOR U23811 ( .A(n23565), .B(n23564), .Z(n23568) );
  XNOR U23812 ( .A(n23569), .B(n23568), .Z(n23571) );
  NAND U23813 ( .A(b[59]), .B(a[55]), .Z(n23570) );
  XOR U23814 ( .A(n23571), .B(n23570), .Z(n23577) );
  XOR U23815 ( .A(n23576), .B(n23577), .Z(n23580) );
  OR U23816 ( .A(n23509), .B(n23508), .Z(n23513) );
  NANDN U23817 ( .A(n23511), .B(n23510), .Z(n23512) );
  NAND U23818 ( .A(n23513), .B(n23512), .Z(n23581) );
  XOR U23819 ( .A(n23580), .B(n23581), .Z(n23582) );
  XOR U23820 ( .A(n23583), .B(n23582), .Z(n23587) );
  OR U23821 ( .A(n23515), .B(n23514), .Z(n23519) );
  NANDN U23822 ( .A(n23517), .B(n23516), .Z(n23518) );
  NAND U23823 ( .A(n23519), .B(n23518), .Z(n23585) );
  NAND U23824 ( .A(b[56]), .B(a[58]), .Z(n23584) );
  XOR U23825 ( .A(n23585), .B(n23584), .Z(n23586) );
  XOR U23826 ( .A(n23587), .B(n23586), .Z(n23590) );
  XNOR U23827 ( .A(n23591), .B(n23590), .Z(n23593) );
  NAND U23828 ( .A(b[55]), .B(a[59]), .Z(n23592) );
  XOR U23829 ( .A(n23593), .B(n23592), .Z(n23599) );
  XOR U23830 ( .A(n23598), .B(n23599), .Z(n23602) );
  NANDN U23831 ( .A(n23521), .B(n23520), .Z(n23525) );
  NANDN U23832 ( .A(n23523), .B(n23522), .Z(n23524) );
  NAND U23833 ( .A(n23525), .B(n23524), .Z(n23603) );
  XOR U23834 ( .A(n23602), .B(n23603), .Z(n23604) );
  XOR U23835 ( .A(n23605), .B(n23604), .Z(n23609) );
  OR U23836 ( .A(n23527), .B(n23526), .Z(n23531) );
  NANDN U23837 ( .A(n23529), .B(n23528), .Z(n23530) );
  NAND U23838 ( .A(n23531), .B(n23530), .Z(n23607) );
  NAND U23839 ( .A(b[52]), .B(a[62]), .Z(n23606) );
  XOR U23840 ( .A(n23607), .B(n23606), .Z(n23608) );
  XOR U23841 ( .A(n23609), .B(n23608), .Z(n23612) );
  NANDN U23842 ( .A(n23533), .B(n23532), .Z(n23537) );
  NANDN U23843 ( .A(n23535), .B(n23534), .Z(n23536) );
  NAND U23844 ( .A(n23537), .B(n23536), .Z(n23613) );
  XOR U23845 ( .A(n23612), .B(n23613), .Z(n23614) );
  XOR U23846 ( .A(n23615), .B(n23614), .Z(n23548) );
  OR U23847 ( .A(n23539), .B(n23538), .Z(n23543) );
  NANDN U23848 ( .A(n23541), .B(n23540), .Z(n23542) );
  AND U23849 ( .A(n23543), .B(n23542), .Z(n23549) );
  XOR U23850 ( .A(n23548), .B(n23549), .Z(n23619) );
  XOR U23851 ( .A(n23618), .B(n23619), .Z(n23620) );
  XOR U23852 ( .A(n23620), .B(n23621), .Z(c[114]) );
  AND U23853 ( .A(n23549), .B(n23548), .Z(n23690) );
  AND U23854 ( .A(b[63]), .B(a[52]), .Z(n23639) );
  AND U23855 ( .A(b[62]), .B(a[53]), .Z(n23637) );
  OR U23856 ( .A(n23551), .B(n23550), .Z(n23555) );
  NANDN U23857 ( .A(n23553), .B(n23552), .Z(n23554) );
  AND U23858 ( .A(n23555), .B(n23554), .Z(n23636) );
  XNOR U23859 ( .A(n23637), .B(n23636), .Z(n23638) );
  XOR U23860 ( .A(n23639), .B(n23638), .Z(n23645) );
  NANDN U23861 ( .A(n23557), .B(n23556), .Z(n23561) );
  NANDN U23862 ( .A(n23559), .B(n23558), .Z(n23560) );
  NAND U23863 ( .A(n23561), .B(n23560), .Z(n23643) );
  NAND U23864 ( .A(b[61]), .B(a[54]), .Z(n23642) );
  XOR U23865 ( .A(n23643), .B(n23642), .Z(n23644) );
  XOR U23866 ( .A(n23645), .B(n23644), .Z(n23651) );
  AND U23867 ( .A(a[55]), .B(b[60]), .Z(n23648) );
  OR U23868 ( .A(n23563), .B(n23562), .Z(n23567) );
  NAND U23869 ( .A(n23565), .B(n23564), .Z(n23566) );
  NAND U23870 ( .A(n23567), .B(n23566), .Z(n23649) );
  XOR U23871 ( .A(n23648), .B(n23649), .Z(n23650) );
  XNOR U23872 ( .A(n23651), .B(n23650), .Z(n23633) );
  NAND U23873 ( .A(n23569), .B(n23568), .Z(n23573) );
  OR U23874 ( .A(n23571), .B(n23570), .Z(n23572) );
  NAND U23875 ( .A(n23573), .B(n23572), .Z(n23630) );
  NAND U23876 ( .A(a[56]), .B(b[59]), .Z(n23631) );
  XNOR U23877 ( .A(n23630), .B(n23631), .Z(n23632) );
  XNOR U23878 ( .A(n23633), .B(n23632), .Z(n23627) );
  AND U23879 ( .A(a[57]), .B(b[58]), .Z(n23624) );
  OR U23880 ( .A(n23575), .B(n23574), .Z(n23579) );
  NAND U23881 ( .A(n23577), .B(n23576), .Z(n23578) );
  NAND U23882 ( .A(n23579), .B(n23578), .Z(n23625) );
  XOR U23883 ( .A(n23624), .B(n23625), .Z(n23626) );
  XNOR U23884 ( .A(n23627), .B(n23626), .Z(n23657) );
  NAND U23885 ( .A(b[57]), .B(a[58]), .Z(n23654) );
  XOR U23886 ( .A(n23655), .B(n23654), .Z(n23656) );
  XNOR U23887 ( .A(n23657), .B(n23656), .Z(n23663) );
  AND U23888 ( .A(a[59]), .B(b[56]), .Z(n23660) );
  OR U23889 ( .A(n23585), .B(n23584), .Z(n23589) );
  NAND U23890 ( .A(n23587), .B(n23586), .Z(n23588) );
  NAND U23891 ( .A(n23589), .B(n23588), .Z(n23661) );
  XOR U23892 ( .A(n23660), .B(n23661), .Z(n23662) );
  XNOR U23893 ( .A(n23663), .B(n23662), .Z(n23669) );
  NAND U23894 ( .A(n23591), .B(n23590), .Z(n23595) );
  OR U23895 ( .A(n23593), .B(n23592), .Z(n23594) );
  NAND U23896 ( .A(n23595), .B(n23594), .Z(n23666) );
  NAND U23897 ( .A(a[60]), .B(b[55]), .Z(n23667) );
  XNOR U23898 ( .A(n23666), .B(n23667), .Z(n23668) );
  XNOR U23899 ( .A(n23669), .B(n23668), .Z(n23675) );
  AND U23900 ( .A(a[61]), .B(b[54]), .Z(n23672) );
  OR U23901 ( .A(n23597), .B(n23596), .Z(n23601) );
  NAND U23902 ( .A(n23599), .B(n23598), .Z(n23600) );
  NAND U23903 ( .A(n23601), .B(n23600), .Z(n23673) );
  XOR U23904 ( .A(n23672), .B(n23673), .Z(n23674) );
  XNOR U23905 ( .A(n23675), .B(n23674), .Z(n23681) );
  NAND U23906 ( .A(b[53]), .B(a[62]), .Z(n23678) );
  XOR U23907 ( .A(n23679), .B(n23678), .Z(n23680) );
  XNOR U23908 ( .A(n23681), .B(n23680), .Z(n23687) );
  AND U23909 ( .A(a[63]), .B(b[52]), .Z(n23684) );
  OR U23910 ( .A(n23607), .B(n23606), .Z(n23611) );
  NAND U23911 ( .A(n23609), .B(n23608), .Z(n23610) );
  NAND U23912 ( .A(n23611), .B(n23610), .Z(n23685) );
  XOR U23913 ( .A(n23684), .B(n23685), .Z(n23686) );
  XNOR U23914 ( .A(n23687), .B(n23686), .Z(n23622) );
  OR U23915 ( .A(n23613), .B(n23612), .Z(n23617) );
  NANDN U23916 ( .A(n23615), .B(n23614), .Z(n23616) );
  AND U23917 ( .A(n23617), .B(n23616), .Z(n23623) );
  XNOR U23918 ( .A(n23622), .B(n23623), .Z(n23691) );
  XOR U23919 ( .A(n23690), .B(n23691), .Z(n23692) );
  XOR U23920 ( .A(n23692), .B(n23693), .Z(c[115]) );
  ANDN U23921 ( .B(n23623), .A(n23622), .Z(n23754) );
  AND U23922 ( .A(a[63]), .B(b[53]), .Z(n23751) );
  AND U23923 ( .A(a[61]), .B(b[55]), .Z(n23739) );
  AND U23924 ( .A(a[59]), .B(b[57]), .Z(n23729) );
  OR U23925 ( .A(n23625), .B(n23624), .Z(n23629) );
  NANDN U23926 ( .A(n23627), .B(n23626), .Z(n23628) );
  NAND U23927 ( .A(n23629), .B(n23628), .Z(n23721) );
  NAND U23928 ( .A(b[58]), .B(a[58]), .Z(n23720) );
  XOR U23929 ( .A(n23721), .B(n23720), .Z(n23722) );
  NANDN U23930 ( .A(n23631), .B(n23630), .Z(n23635) );
  NANDN U23931 ( .A(n23633), .B(n23632), .Z(n23634) );
  NAND U23932 ( .A(n23635), .B(n23634), .Z(n23715) );
  AND U23933 ( .A(a[55]), .B(b[61]), .Z(n23705) );
  NANDN U23934 ( .A(n23637), .B(n23636), .Z(n23641) );
  NANDN U23935 ( .A(n23639), .B(n23638), .Z(n23640) );
  NAND U23936 ( .A(n23641), .B(n23640), .Z(n23697) );
  NAND U23937 ( .A(a[54]), .B(b[62]), .Z(n23696) );
  XOR U23938 ( .A(n23697), .B(n23696), .Z(n23698) );
  NAND U23939 ( .A(a[53]), .B(b[63]), .Z(n23699) );
  XOR U23940 ( .A(n23698), .B(n23699), .Z(n23702) );
  OR U23941 ( .A(n23643), .B(n23642), .Z(n23647) );
  NAND U23942 ( .A(n23645), .B(n23644), .Z(n23646) );
  NAND U23943 ( .A(n23647), .B(n23646), .Z(n23703) );
  XNOR U23944 ( .A(n23702), .B(n23703), .Z(n23704) );
  XOR U23945 ( .A(n23705), .B(n23704), .Z(n23711) );
  OR U23946 ( .A(n23649), .B(n23648), .Z(n23653) );
  NANDN U23947 ( .A(n23651), .B(n23650), .Z(n23652) );
  NAND U23948 ( .A(n23653), .B(n23652), .Z(n23709) );
  NAND U23949 ( .A(b[60]), .B(a[56]), .Z(n23708) );
  XOR U23950 ( .A(n23709), .B(n23708), .Z(n23710) );
  XOR U23951 ( .A(n23711), .B(n23710), .Z(n23714) );
  XNOR U23952 ( .A(n23715), .B(n23714), .Z(n23717) );
  NAND U23953 ( .A(b[59]), .B(a[57]), .Z(n23716) );
  XOR U23954 ( .A(n23717), .B(n23716), .Z(n23723) );
  XOR U23955 ( .A(n23722), .B(n23723), .Z(n23726) );
  OR U23956 ( .A(n23655), .B(n23654), .Z(n23659) );
  NANDN U23957 ( .A(n23657), .B(n23656), .Z(n23658) );
  NAND U23958 ( .A(n23659), .B(n23658), .Z(n23727) );
  XOR U23959 ( .A(n23726), .B(n23727), .Z(n23728) );
  XOR U23960 ( .A(n23729), .B(n23728), .Z(n23733) );
  OR U23961 ( .A(n23661), .B(n23660), .Z(n23665) );
  NANDN U23962 ( .A(n23663), .B(n23662), .Z(n23664) );
  NAND U23963 ( .A(n23665), .B(n23664), .Z(n23731) );
  NAND U23964 ( .A(b[56]), .B(a[60]), .Z(n23730) );
  XOR U23965 ( .A(n23731), .B(n23730), .Z(n23732) );
  XOR U23966 ( .A(n23733), .B(n23732), .Z(n23736) );
  NANDN U23967 ( .A(n23667), .B(n23666), .Z(n23671) );
  NANDN U23968 ( .A(n23669), .B(n23668), .Z(n23670) );
  NAND U23969 ( .A(n23671), .B(n23670), .Z(n23737) );
  XOR U23970 ( .A(n23736), .B(n23737), .Z(n23738) );
  XOR U23971 ( .A(n23739), .B(n23738), .Z(n23745) );
  OR U23972 ( .A(n23673), .B(n23672), .Z(n23677) );
  NANDN U23973 ( .A(n23675), .B(n23674), .Z(n23676) );
  NAND U23974 ( .A(n23677), .B(n23676), .Z(n23743) );
  NAND U23975 ( .A(b[54]), .B(a[62]), .Z(n23742) );
  XOR U23976 ( .A(n23743), .B(n23742), .Z(n23744) );
  XOR U23977 ( .A(n23745), .B(n23744), .Z(n23748) );
  OR U23978 ( .A(n23679), .B(n23678), .Z(n23683) );
  NANDN U23979 ( .A(n23681), .B(n23680), .Z(n23682) );
  NAND U23980 ( .A(n23683), .B(n23682), .Z(n23749) );
  XOR U23981 ( .A(n23748), .B(n23749), .Z(n23750) );
  XOR U23982 ( .A(n23751), .B(n23750), .Z(n23694) );
  OR U23983 ( .A(n23685), .B(n23684), .Z(n23689) );
  NANDN U23984 ( .A(n23687), .B(n23686), .Z(n23688) );
  AND U23985 ( .A(n23689), .B(n23688), .Z(n23695) );
  XOR U23986 ( .A(n23694), .B(n23695), .Z(n23755) );
  XOR U23987 ( .A(n23754), .B(n23755), .Z(n23756) );
  XOR U23988 ( .A(n23756), .B(n23757), .Z(c[116]) );
  AND U23989 ( .A(n23695), .B(n23694), .Z(n23814) );
  AND U23990 ( .A(b[63]), .B(a[54]), .Z(n23775) );
  AND U23991 ( .A(b[62]), .B(a[55]), .Z(n23773) );
  OR U23992 ( .A(n23697), .B(n23696), .Z(n23701) );
  NANDN U23993 ( .A(n23699), .B(n23698), .Z(n23700) );
  AND U23994 ( .A(n23701), .B(n23700), .Z(n23772) );
  XNOR U23995 ( .A(n23773), .B(n23772), .Z(n23774) );
  XOR U23996 ( .A(n23775), .B(n23774), .Z(n23781) );
  NANDN U23997 ( .A(n23703), .B(n23702), .Z(n23707) );
  NANDN U23998 ( .A(n23705), .B(n23704), .Z(n23706) );
  NAND U23999 ( .A(n23707), .B(n23706), .Z(n23779) );
  NAND U24000 ( .A(b[61]), .B(a[56]), .Z(n23778) );
  XOR U24001 ( .A(n23779), .B(n23778), .Z(n23780) );
  XOR U24002 ( .A(n23781), .B(n23780), .Z(n23787) );
  AND U24003 ( .A(a[57]), .B(b[60]), .Z(n23784) );
  OR U24004 ( .A(n23709), .B(n23708), .Z(n23713) );
  NAND U24005 ( .A(n23711), .B(n23710), .Z(n23712) );
  NAND U24006 ( .A(n23713), .B(n23712), .Z(n23785) );
  XOR U24007 ( .A(n23784), .B(n23785), .Z(n23786) );
  XNOR U24008 ( .A(n23787), .B(n23786), .Z(n23769) );
  NAND U24009 ( .A(n23715), .B(n23714), .Z(n23719) );
  OR U24010 ( .A(n23717), .B(n23716), .Z(n23718) );
  NAND U24011 ( .A(n23719), .B(n23718), .Z(n23766) );
  NAND U24012 ( .A(a[58]), .B(b[59]), .Z(n23767) );
  XNOR U24013 ( .A(n23766), .B(n23767), .Z(n23768) );
  XNOR U24014 ( .A(n23769), .B(n23768), .Z(n23763) );
  AND U24015 ( .A(a[59]), .B(b[58]), .Z(n23760) );
  OR U24016 ( .A(n23721), .B(n23720), .Z(n23725) );
  NAND U24017 ( .A(n23723), .B(n23722), .Z(n23724) );
  NAND U24018 ( .A(n23725), .B(n23724), .Z(n23761) );
  XOR U24019 ( .A(n23760), .B(n23761), .Z(n23762) );
  XNOR U24020 ( .A(n23763), .B(n23762), .Z(n23793) );
  NAND U24021 ( .A(b[57]), .B(a[60]), .Z(n23790) );
  XOR U24022 ( .A(n23791), .B(n23790), .Z(n23792) );
  XNOR U24023 ( .A(n23793), .B(n23792), .Z(n23799) );
  AND U24024 ( .A(a[61]), .B(b[56]), .Z(n23796) );
  OR U24025 ( .A(n23731), .B(n23730), .Z(n23735) );
  NAND U24026 ( .A(n23733), .B(n23732), .Z(n23734) );
  NAND U24027 ( .A(n23735), .B(n23734), .Z(n23797) );
  XOR U24028 ( .A(n23796), .B(n23797), .Z(n23798) );
  XNOR U24029 ( .A(n23799), .B(n23798), .Z(n23805) );
  OR U24030 ( .A(n23737), .B(n23736), .Z(n23741) );
  NANDN U24031 ( .A(n23739), .B(n23738), .Z(n23740) );
  NAND U24032 ( .A(n23741), .B(n23740), .Z(n23803) );
  NAND U24033 ( .A(b[55]), .B(a[62]), .Z(n23802) );
  XOR U24034 ( .A(n23803), .B(n23802), .Z(n23804) );
  XNOR U24035 ( .A(n23805), .B(n23804), .Z(n23811) );
  AND U24036 ( .A(a[63]), .B(b[54]), .Z(n23808) );
  OR U24037 ( .A(n23743), .B(n23742), .Z(n23747) );
  NAND U24038 ( .A(n23745), .B(n23744), .Z(n23746) );
  NAND U24039 ( .A(n23747), .B(n23746), .Z(n23809) );
  XOR U24040 ( .A(n23808), .B(n23809), .Z(n23810) );
  XNOR U24041 ( .A(n23811), .B(n23810), .Z(n23758) );
  OR U24042 ( .A(n23749), .B(n23748), .Z(n23753) );
  NANDN U24043 ( .A(n23751), .B(n23750), .Z(n23752) );
  AND U24044 ( .A(n23753), .B(n23752), .Z(n23759) );
  XNOR U24045 ( .A(n23758), .B(n23759), .Z(n23815) );
  XOR U24046 ( .A(n23814), .B(n23815), .Z(n23816) );
  XOR U24047 ( .A(n23816), .B(n23817), .Z(c[117]) );
  ANDN U24048 ( .B(n23759), .A(n23758), .Z(n23866) );
  AND U24049 ( .A(a[63]), .B(b[55]), .Z(n23863) );
  AND U24050 ( .A(a[61]), .B(b[57]), .Z(n23853) );
  OR U24051 ( .A(n23761), .B(n23760), .Z(n23765) );
  NANDN U24052 ( .A(n23763), .B(n23762), .Z(n23764) );
  NAND U24053 ( .A(n23765), .B(n23764), .Z(n23845) );
  NAND U24054 ( .A(b[58]), .B(a[60]), .Z(n23844) );
  XOR U24055 ( .A(n23845), .B(n23844), .Z(n23846) );
  NANDN U24056 ( .A(n23767), .B(n23766), .Z(n23771) );
  NANDN U24057 ( .A(n23769), .B(n23768), .Z(n23770) );
  NAND U24058 ( .A(n23771), .B(n23770), .Z(n23839) );
  AND U24059 ( .A(a[57]), .B(b[61]), .Z(n23829) );
  NANDN U24060 ( .A(n23773), .B(n23772), .Z(n23777) );
  NANDN U24061 ( .A(n23775), .B(n23774), .Z(n23776) );
  NAND U24062 ( .A(n23777), .B(n23776), .Z(n23821) );
  NAND U24063 ( .A(a[56]), .B(b[62]), .Z(n23820) );
  XOR U24064 ( .A(n23821), .B(n23820), .Z(n23822) );
  NAND U24065 ( .A(a[55]), .B(b[63]), .Z(n23823) );
  XOR U24066 ( .A(n23822), .B(n23823), .Z(n23826) );
  OR U24067 ( .A(n23779), .B(n23778), .Z(n23783) );
  NAND U24068 ( .A(n23781), .B(n23780), .Z(n23782) );
  NAND U24069 ( .A(n23783), .B(n23782), .Z(n23827) );
  XNOR U24070 ( .A(n23826), .B(n23827), .Z(n23828) );
  XOR U24071 ( .A(n23829), .B(n23828), .Z(n23835) );
  OR U24072 ( .A(n23785), .B(n23784), .Z(n23789) );
  NANDN U24073 ( .A(n23787), .B(n23786), .Z(n23788) );
  NAND U24074 ( .A(n23789), .B(n23788), .Z(n23833) );
  NAND U24075 ( .A(b[60]), .B(a[58]), .Z(n23832) );
  XOR U24076 ( .A(n23833), .B(n23832), .Z(n23834) );
  XOR U24077 ( .A(n23835), .B(n23834), .Z(n23838) );
  XNOR U24078 ( .A(n23839), .B(n23838), .Z(n23841) );
  NAND U24079 ( .A(b[59]), .B(a[59]), .Z(n23840) );
  XOR U24080 ( .A(n23841), .B(n23840), .Z(n23847) );
  XOR U24081 ( .A(n23846), .B(n23847), .Z(n23850) );
  OR U24082 ( .A(n23791), .B(n23790), .Z(n23795) );
  NANDN U24083 ( .A(n23793), .B(n23792), .Z(n23794) );
  NAND U24084 ( .A(n23795), .B(n23794), .Z(n23851) );
  XOR U24085 ( .A(n23850), .B(n23851), .Z(n23852) );
  XOR U24086 ( .A(n23853), .B(n23852), .Z(n23857) );
  OR U24087 ( .A(n23797), .B(n23796), .Z(n23801) );
  NANDN U24088 ( .A(n23799), .B(n23798), .Z(n23800) );
  NAND U24089 ( .A(n23801), .B(n23800), .Z(n23855) );
  NAND U24090 ( .A(b[56]), .B(a[62]), .Z(n23854) );
  XOR U24091 ( .A(n23855), .B(n23854), .Z(n23856) );
  XOR U24092 ( .A(n23857), .B(n23856), .Z(n23860) );
  OR U24093 ( .A(n23803), .B(n23802), .Z(n23807) );
  NANDN U24094 ( .A(n23805), .B(n23804), .Z(n23806) );
  NAND U24095 ( .A(n23807), .B(n23806), .Z(n23861) );
  XOR U24096 ( .A(n23860), .B(n23861), .Z(n23862) );
  XOR U24097 ( .A(n23863), .B(n23862), .Z(n23818) );
  OR U24098 ( .A(n23809), .B(n23808), .Z(n23813) );
  NANDN U24099 ( .A(n23811), .B(n23810), .Z(n23812) );
  AND U24100 ( .A(n23813), .B(n23812), .Z(n23819) );
  XOR U24101 ( .A(n23818), .B(n23819), .Z(n23867) );
  XOR U24102 ( .A(n23866), .B(n23867), .Z(n23868) );
  XOR U24103 ( .A(n23868), .B(n23869), .Z(c[118]) );
  AND U24104 ( .A(n23819), .B(n23818), .Z(n23914) );
  AND U24105 ( .A(b[63]), .B(a[56]), .Z(n23887) );
  AND U24106 ( .A(b[62]), .B(a[57]), .Z(n23885) );
  OR U24107 ( .A(n23821), .B(n23820), .Z(n23825) );
  NANDN U24108 ( .A(n23823), .B(n23822), .Z(n23824) );
  AND U24109 ( .A(n23825), .B(n23824), .Z(n23884) );
  XNOR U24110 ( .A(n23885), .B(n23884), .Z(n23886) );
  XOR U24111 ( .A(n23887), .B(n23886), .Z(n23893) );
  NANDN U24112 ( .A(n23827), .B(n23826), .Z(n23831) );
  NANDN U24113 ( .A(n23829), .B(n23828), .Z(n23830) );
  NAND U24114 ( .A(n23831), .B(n23830), .Z(n23891) );
  NAND U24115 ( .A(b[61]), .B(a[58]), .Z(n23890) );
  XOR U24116 ( .A(n23891), .B(n23890), .Z(n23892) );
  XOR U24117 ( .A(n23893), .B(n23892), .Z(n23899) );
  AND U24118 ( .A(a[59]), .B(b[60]), .Z(n23896) );
  OR U24119 ( .A(n23833), .B(n23832), .Z(n23837) );
  NAND U24120 ( .A(n23835), .B(n23834), .Z(n23836) );
  NAND U24121 ( .A(n23837), .B(n23836), .Z(n23897) );
  XOR U24122 ( .A(n23896), .B(n23897), .Z(n23898) );
  XNOR U24123 ( .A(n23899), .B(n23898), .Z(n23881) );
  NAND U24124 ( .A(n23839), .B(n23838), .Z(n23843) );
  OR U24125 ( .A(n23841), .B(n23840), .Z(n23842) );
  NAND U24126 ( .A(n23843), .B(n23842), .Z(n23878) );
  NAND U24127 ( .A(a[60]), .B(b[59]), .Z(n23879) );
  XNOR U24128 ( .A(n23878), .B(n23879), .Z(n23880) );
  XNOR U24129 ( .A(n23881), .B(n23880), .Z(n23875) );
  AND U24130 ( .A(a[61]), .B(b[58]), .Z(n23872) );
  OR U24131 ( .A(n23845), .B(n23844), .Z(n23849) );
  NAND U24132 ( .A(n23847), .B(n23846), .Z(n23848) );
  NAND U24133 ( .A(n23849), .B(n23848), .Z(n23873) );
  XOR U24134 ( .A(n23872), .B(n23873), .Z(n23874) );
  XNOR U24135 ( .A(n23875), .B(n23874), .Z(n23905) );
  NAND U24136 ( .A(b[57]), .B(a[62]), .Z(n23902) );
  XOR U24137 ( .A(n23903), .B(n23902), .Z(n23904) );
  XNOR U24138 ( .A(n23905), .B(n23904), .Z(n23911) );
  AND U24139 ( .A(a[63]), .B(b[56]), .Z(n23908) );
  OR U24140 ( .A(n23855), .B(n23854), .Z(n23859) );
  NAND U24141 ( .A(n23857), .B(n23856), .Z(n23858) );
  NAND U24142 ( .A(n23859), .B(n23858), .Z(n23909) );
  XOR U24143 ( .A(n23908), .B(n23909), .Z(n23910) );
  XNOR U24144 ( .A(n23911), .B(n23910), .Z(n23870) );
  OR U24145 ( .A(n23861), .B(n23860), .Z(n23865) );
  NANDN U24146 ( .A(n23863), .B(n23862), .Z(n23864) );
  AND U24147 ( .A(n23865), .B(n23864), .Z(n23871) );
  XNOR U24148 ( .A(n23870), .B(n23871), .Z(n23915) );
  XOR U24149 ( .A(n23914), .B(n23915), .Z(n23916) );
  XOR U24150 ( .A(n23916), .B(n23917), .Z(c[119]) );
  ANDN U24151 ( .B(n23871), .A(n23870), .Z(n23954) );
  AND U24152 ( .A(a[63]), .B(b[57]), .Z(n23953) );
  OR U24153 ( .A(n23873), .B(n23872), .Z(n23877) );
  NANDN U24154 ( .A(n23875), .B(n23874), .Z(n23876) );
  NAND U24155 ( .A(n23877), .B(n23876), .Z(n23945) );
  NAND U24156 ( .A(b[58]), .B(a[62]), .Z(n23944) );
  XOR U24157 ( .A(n23945), .B(n23944), .Z(n23946) );
  NANDN U24158 ( .A(n23879), .B(n23878), .Z(n23883) );
  NANDN U24159 ( .A(n23881), .B(n23880), .Z(n23882) );
  NAND U24160 ( .A(n23883), .B(n23882), .Z(n23939) );
  AND U24161 ( .A(a[59]), .B(b[61]), .Z(n23929) );
  NANDN U24162 ( .A(n23885), .B(n23884), .Z(n23889) );
  NANDN U24163 ( .A(n23887), .B(n23886), .Z(n23888) );
  NAND U24164 ( .A(n23889), .B(n23888), .Z(n23921) );
  NAND U24165 ( .A(a[58]), .B(b[62]), .Z(n23920) );
  XOR U24166 ( .A(n23921), .B(n23920), .Z(n23922) );
  NAND U24167 ( .A(a[57]), .B(b[63]), .Z(n23923) );
  XOR U24168 ( .A(n23922), .B(n23923), .Z(n23926) );
  OR U24169 ( .A(n23891), .B(n23890), .Z(n23895) );
  NAND U24170 ( .A(n23893), .B(n23892), .Z(n23894) );
  NAND U24171 ( .A(n23895), .B(n23894), .Z(n23927) );
  XNOR U24172 ( .A(n23926), .B(n23927), .Z(n23928) );
  XOR U24173 ( .A(n23929), .B(n23928), .Z(n23935) );
  OR U24174 ( .A(n23897), .B(n23896), .Z(n23901) );
  NANDN U24175 ( .A(n23899), .B(n23898), .Z(n23900) );
  NAND U24176 ( .A(n23901), .B(n23900), .Z(n23933) );
  NAND U24177 ( .A(b[60]), .B(a[60]), .Z(n23932) );
  XOR U24178 ( .A(n23933), .B(n23932), .Z(n23934) );
  XOR U24179 ( .A(n23935), .B(n23934), .Z(n23938) );
  XNOR U24180 ( .A(n23939), .B(n23938), .Z(n23941) );
  NAND U24181 ( .A(b[59]), .B(a[61]), .Z(n23940) );
  XOR U24182 ( .A(n23941), .B(n23940), .Z(n23947) );
  XOR U24183 ( .A(n23946), .B(n23947), .Z(n23950) );
  OR U24184 ( .A(n23903), .B(n23902), .Z(n23907) );
  NANDN U24185 ( .A(n23905), .B(n23904), .Z(n23906) );
  NAND U24186 ( .A(n23907), .B(n23906), .Z(n23951) );
  XOR U24187 ( .A(n23950), .B(n23951), .Z(n23952) );
  XOR U24188 ( .A(n23953), .B(n23952), .Z(n23918) );
  OR U24189 ( .A(n23909), .B(n23908), .Z(n23913) );
  NANDN U24190 ( .A(n23911), .B(n23910), .Z(n23912) );
  AND U24191 ( .A(n23913), .B(n23912), .Z(n23919) );
  XOR U24192 ( .A(n23918), .B(n23919), .Z(n23955) );
  XOR U24193 ( .A(n23954), .B(n23955), .Z(n23956) );
  XOR U24194 ( .A(n23956), .B(n23957), .Z(c[120]) );
  AND U24195 ( .A(n23919), .B(n23918), .Z(n23990) );
  AND U24196 ( .A(b[63]), .B(a[58]), .Z(n23963) );
  AND U24197 ( .A(b[62]), .B(a[59]), .Z(n23961) );
  OR U24198 ( .A(n23921), .B(n23920), .Z(n23925) );
  NANDN U24199 ( .A(n23923), .B(n23922), .Z(n23924) );
  AND U24200 ( .A(n23925), .B(n23924), .Z(n23960) );
  XNOR U24201 ( .A(n23961), .B(n23960), .Z(n23962) );
  XOR U24202 ( .A(n23963), .B(n23962), .Z(n23969) );
  NANDN U24203 ( .A(n23927), .B(n23926), .Z(n23931) );
  NANDN U24204 ( .A(n23929), .B(n23928), .Z(n23930) );
  NAND U24205 ( .A(n23931), .B(n23930), .Z(n23967) );
  NAND U24206 ( .A(b[61]), .B(a[60]), .Z(n23966) );
  XOR U24207 ( .A(n23967), .B(n23966), .Z(n23968) );
  XOR U24208 ( .A(n23969), .B(n23968), .Z(n23975) );
  AND U24209 ( .A(a[61]), .B(b[60]), .Z(n23972) );
  OR U24210 ( .A(n23933), .B(n23932), .Z(n23937) );
  NAND U24211 ( .A(n23935), .B(n23934), .Z(n23936) );
  NAND U24212 ( .A(n23937), .B(n23936), .Z(n23973) );
  XOR U24213 ( .A(n23972), .B(n23973), .Z(n23974) );
  XNOR U24214 ( .A(n23975), .B(n23974), .Z(n23981) );
  NAND U24215 ( .A(n23939), .B(n23938), .Z(n23943) );
  OR U24216 ( .A(n23941), .B(n23940), .Z(n23942) );
  NAND U24217 ( .A(n23943), .B(n23942), .Z(n23978) );
  NAND U24218 ( .A(a[62]), .B(b[59]), .Z(n23979) );
  XNOR U24219 ( .A(n23978), .B(n23979), .Z(n23980) );
  XNOR U24220 ( .A(n23981), .B(n23980), .Z(n23987) );
  AND U24221 ( .A(a[63]), .B(b[58]), .Z(n23984) );
  OR U24222 ( .A(n23945), .B(n23944), .Z(n23949) );
  NAND U24223 ( .A(n23947), .B(n23946), .Z(n23948) );
  NAND U24224 ( .A(n23949), .B(n23948), .Z(n23985) );
  XOR U24225 ( .A(n23984), .B(n23985), .Z(n23986) );
  XNOR U24226 ( .A(n23987), .B(n23986), .Z(n23958) );
  XNOR U24227 ( .A(n23958), .B(n23959), .Z(n23991) );
  XOR U24228 ( .A(n23990), .B(n23991), .Z(n23992) );
  XOR U24229 ( .A(n23992), .B(n23993), .Z(c[121]) );
  ANDN U24230 ( .B(n23959), .A(n23958), .Z(n24020) );
  AND U24231 ( .A(a[63]), .B(b[59]), .Z(n24017) );
  AND U24232 ( .A(a[61]), .B(b[61]), .Z(n24005) );
  NANDN U24233 ( .A(n23961), .B(n23960), .Z(n23965) );
  NANDN U24234 ( .A(n23963), .B(n23962), .Z(n23964) );
  NAND U24235 ( .A(n23965), .B(n23964), .Z(n23997) );
  NAND U24236 ( .A(a[60]), .B(b[62]), .Z(n23996) );
  XOR U24237 ( .A(n23997), .B(n23996), .Z(n23998) );
  NAND U24238 ( .A(a[59]), .B(b[63]), .Z(n23999) );
  XOR U24239 ( .A(n23998), .B(n23999), .Z(n24002) );
  OR U24240 ( .A(n23967), .B(n23966), .Z(n23971) );
  NAND U24241 ( .A(n23969), .B(n23968), .Z(n23970) );
  NAND U24242 ( .A(n23971), .B(n23970), .Z(n24003) );
  XNOR U24243 ( .A(n24002), .B(n24003), .Z(n24004) );
  XOR U24244 ( .A(n24005), .B(n24004), .Z(n24011) );
  OR U24245 ( .A(n23973), .B(n23972), .Z(n23977) );
  NANDN U24246 ( .A(n23975), .B(n23974), .Z(n23976) );
  NAND U24247 ( .A(n23977), .B(n23976), .Z(n24009) );
  NAND U24248 ( .A(b[60]), .B(a[62]), .Z(n24008) );
  XOR U24249 ( .A(n24009), .B(n24008), .Z(n24010) );
  XOR U24250 ( .A(n24011), .B(n24010), .Z(n24014) );
  NANDN U24251 ( .A(n23979), .B(n23978), .Z(n23983) );
  NANDN U24252 ( .A(n23981), .B(n23980), .Z(n23982) );
  NAND U24253 ( .A(n23983), .B(n23982), .Z(n24015) );
  XOR U24254 ( .A(n24014), .B(n24015), .Z(n24016) );
  XOR U24255 ( .A(n24017), .B(n24016), .Z(n23994) );
  OR U24256 ( .A(n23985), .B(n23984), .Z(n23989) );
  NANDN U24257 ( .A(n23987), .B(n23986), .Z(n23988) );
  AND U24258 ( .A(n23989), .B(n23988), .Z(n23995) );
  XOR U24259 ( .A(n23994), .B(n23995), .Z(n24021) );
  XOR U24260 ( .A(n24020), .B(n24021), .Z(n24022) );
  XOR U24261 ( .A(n24022), .B(n24023), .Z(c[122]) );
  AND U24262 ( .A(n23995), .B(n23994), .Z(n24044) );
  AND U24263 ( .A(b[63]), .B(a[60]), .Z(n24029) );
  AND U24264 ( .A(b[62]), .B(a[61]), .Z(n24027) );
  OR U24265 ( .A(n23997), .B(n23996), .Z(n24001) );
  NANDN U24266 ( .A(n23999), .B(n23998), .Z(n24000) );
  AND U24267 ( .A(n24001), .B(n24000), .Z(n24026) );
  XNOR U24268 ( .A(n24027), .B(n24026), .Z(n24028) );
  XOR U24269 ( .A(n24029), .B(n24028), .Z(n24035) );
  NANDN U24270 ( .A(n24003), .B(n24002), .Z(n24007) );
  NANDN U24271 ( .A(n24005), .B(n24004), .Z(n24006) );
  NAND U24272 ( .A(n24007), .B(n24006), .Z(n24033) );
  NAND U24273 ( .A(b[61]), .B(a[62]), .Z(n24032) );
  XOR U24274 ( .A(n24033), .B(n24032), .Z(n24034) );
  XOR U24275 ( .A(n24035), .B(n24034), .Z(n24041) );
  AND U24276 ( .A(a[63]), .B(b[60]), .Z(n24038) );
  OR U24277 ( .A(n24009), .B(n24008), .Z(n24013) );
  NAND U24278 ( .A(n24011), .B(n24010), .Z(n24012) );
  NAND U24279 ( .A(n24013), .B(n24012), .Z(n24039) );
  XOR U24280 ( .A(n24038), .B(n24039), .Z(n24040) );
  XNOR U24281 ( .A(n24041), .B(n24040), .Z(n24024) );
  OR U24282 ( .A(n24015), .B(n24014), .Z(n24019) );
  NANDN U24283 ( .A(n24017), .B(n24016), .Z(n24018) );
  AND U24284 ( .A(n24019), .B(n24018), .Z(n24025) );
  XNOR U24285 ( .A(n24024), .B(n24025), .Z(n24045) );
  XOR U24286 ( .A(n24044), .B(n24045), .Z(n24046) );
  XOR U24287 ( .A(n24046), .B(n24047), .Z(c[123]) );
  ANDN U24288 ( .B(n24025), .A(n24024), .Z(n24062) );
  AND U24289 ( .A(a[63]), .B(b[61]), .Z(n24059) );
  NANDN U24290 ( .A(n24027), .B(n24026), .Z(n24031) );
  NANDN U24291 ( .A(n24029), .B(n24028), .Z(n24030) );
  NAND U24292 ( .A(n24031), .B(n24030), .Z(n24051) );
  NAND U24293 ( .A(a[62]), .B(b[62]), .Z(n24050) );
  XOR U24294 ( .A(n24051), .B(n24050), .Z(n24052) );
  NAND U24295 ( .A(a[61]), .B(b[63]), .Z(n24053) );
  XOR U24296 ( .A(n24052), .B(n24053), .Z(n24056) );
  OR U24297 ( .A(n24033), .B(n24032), .Z(n24037) );
  NAND U24298 ( .A(n24035), .B(n24034), .Z(n24036) );
  NAND U24299 ( .A(n24037), .B(n24036), .Z(n24057) );
  XNOR U24300 ( .A(n24056), .B(n24057), .Z(n24058) );
  XOR U24301 ( .A(n24059), .B(n24058), .Z(n24048) );
  OR U24302 ( .A(n24039), .B(n24038), .Z(n24043) );
  NANDN U24303 ( .A(n24041), .B(n24040), .Z(n24042) );
  AND U24304 ( .A(n24043), .B(n24042), .Z(n24049) );
  XOR U24305 ( .A(n24048), .B(n24049), .Z(n24063) );
  XOR U24306 ( .A(n24062), .B(n24063), .Z(n24064) );
  XOR U24307 ( .A(n24064), .B(n24065), .Z(c[124]) );
  AND U24308 ( .A(n24049), .B(n24048), .Z(n24075) );
  AND U24309 ( .A(b[63]), .B(a[62]), .Z(n24071) );
  AND U24310 ( .A(a[63]), .B(b[62]), .Z(n24069) );
  OR U24311 ( .A(n24051), .B(n24050), .Z(n24055) );
  NANDN U24312 ( .A(n24053), .B(n24052), .Z(n24054) );
  AND U24313 ( .A(n24055), .B(n24054), .Z(n24068) );
  XNOR U24314 ( .A(n24069), .B(n24068), .Z(n24070) );
  XOR U24315 ( .A(n24071), .B(n24070), .Z(n24066) );
  NANDN U24316 ( .A(n24057), .B(n24056), .Z(n24061) );
  NANDN U24317 ( .A(n24059), .B(n24058), .Z(n24060) );
  AND U24318 ( .A(n24061), .B(n24060), .Z(n24067) );
  XOR U24319 ( .A(n24066), .B(n24067), .Z(n24076) );
  XOR U24320 ( .A(n24075), .B(n24076), .Z(n24077) );
  XOR U24321 ( .A(n24077), .B(n24078), .Z(c[125]) );
  AND U24322 ( .A(n24067), .B(n24066), .Z(n24082) );
  NANDN U24323 ( .A(n24069), .B(n24068), .Z(n24073) );
  NANDN U24324 ( .A(n24071), .B(n24070), .Z(n24072) );
  AND U24325 ( .A(n24073), .B(n24072), .Z(n24079) );
  NAND U24326 ( .A(a[63]), .B(b[63]), .Z(n24074) );
  XNOR U24327 ( .A(n24079), .B(n24074), .Z(n24083) );
  XNOR U24328 ( .A(n24082), .B(n24083), .Z(n24081) );
  XNOR U24329 ( .A(n24081), .B(n24080), .Z(c[126]) );
  AND U24330 ( .A(n24079), .B(a[63]), .Z(n24087) );
  OR U24331 ( .A(n24081), .B(n24080), .Z(n24085) );
  OR U24332 ( .A(n24083), .B(n24082), .Z(n24084) );
  NAND U24333 ( .A(n24085), .B(n24084), .Z(n24086) );
  XNOR U24334 ( .A(n24087), .B(n24086), .Z(c[127]) );
  XOR U24335 ( .A(n24089), .B(n24088), .Z(c[65]) );
  XOR U24336 ( .A(n24091), .B(n24090), .Z(c[66]) );
  XOR U24337 ( .A(n24093), .B(n24092), .Z(n24098) );
  XOR U24338 ( .A(n24098), .B(n24094), .Z(c[67]) );
  XOR U24339 ( .A(n24096), .B(n24095), .Z(n24101) );
  NANDN U24340 ( .A(n24098), .B(n24097), .Z(n24099) );
  NANDN U24341 ( .A(n24100), .B(n24099), .Z(n24102) );
  XOR U24342 ( .A(n24101), .B(n24102), .Z(c[68]) );
  NAND U24343 ( .A(n24102), .B(n24101), .Z(n24104) );
  ANDN U24344 ( .B(n24104), .A(n24103), .Z(n24108) );
  XOR U24345 ( .A(n24106), .B(n24105), .Z(n24107) );
  XOR U24346 ( .A(n24108), .B(n24107), .Z(c[69]) );
  XOR U24347 ( .A(n24110), .B(n24109), .Z(c[70]) );
  XOR U24348 ( .A(n24112), .B(n24111), .Z(c[71]) );
  XOR U24349 ( .A(n24114), .B(n24113), .Z(c[72]) );
  XNOR U24350 ( .A(n24116), .B(n24115), .Z(c[73]) );
  XNOR U24351 ( .A(n24117), .B(n24120), .Z(n24118) );
  XNOR U24352 ( .A(n24119), .B(n24118), .Z(c[74]) );
  OR U24353 ( .A(n24121), .B(n24120), .Z(n24128) );
  AND U24354 ( .A(n24128), .B(n24122), .Z(n24125) );
  XOR U24355 ( .A(n24123), .B(n24126), .Z(n24124) );
  XNOR U24356 ( .A(n24125), .B(n24124), .Z(c[75]) );
  NAND U24357 ( .A(n24127), .B(n24126), .Z(n24131) );
  NANDN U24358 ( .A(n24129), .B(n24128), .Z(n24130) );
  NAND U24359 ( .A(n24131), .B(n24130), .Z(n24134) );
  XOR U24360 ( .A(n24133), .B(n24132), .Z(n24135) );
  XNOR U24361 ( .A(n24134), .B(n24135), .Z(c[76]) );
  NANDN U24362 ( .A(n24135), .B(n24134), .Z(n24136) );
  NANDN U24363 ( .A(n24137), .B(n24136), .Z(n24141) );
  XOR U24364 ( .A(n24139), .B(n24138), .Z(n24140) );
  XNOR U24365 ( .A(n24141), .B(n24140), .Z(c[77]) );
  XNOR U24366 ( .A(n24143), .B(n24142), .Z(c[78]) );
  XOR U24367 ( .A(n24145), .B(n24144), .Z(c[79]) );
  XNOR U24368 ( .A(n24147), .B(n24146), .Z(c[80]) );
  XOR U24369 ( .A(n24149), .B(n24148), .Z(c[81]) );
  XOR U24370 ( .A(n24151), .B(n24150), .Z(n24152) );
  XOR U24371 ( .A(n24153), .B(n24152), .Z(c[82]) );
  XOR U24372 ( .A(n24155), .B(n24154), .Z(n24156) );
  XOR U24373 ( .A(n24157), .B(n24156), .Z(c[83]) );
  XNOR U24374 ( .A(n24159), .B(n24158), .Z(n24160) );
  XNOR U24375 ( .A(n24161), .B(n24160), .Z(c[84]) );
  XNOR U24376 ( .A(n24163), .B(n24162), .Z(n24164) );
  XOR U24377 ( .A(n24165), .B(n24164), .Z(c[85]) );
  XNOR U24378 ( .A(n24167), .B(n24166), .Z(c[86]) );
  XOR U24379 ( .A(n24169), .B(n24168), .Z(c[87]) );
  XOR U24380 ( .A(n24171), .B(n24170), .Z(c[88]) );
  XNOR U24381 ( .A(n24173), .B(n24172), .Z(c[89]) );
  XOR U24382 ( .A(n24175), .B(n24174), .Z(n24177) );
  XNOR U24383 ( .A(n24177), .B(n24176), .Z(c[90]) );
  NANDN U24384 ( .A(n24177), .B(n24176), .Z(n24178) );
  NANDN U24385 ( .A(n24179), .B(n24178), .Z(n24185) );
  XNOR U24386 ( .A(n24181), .B(n24180), .Z(n24184) );
  XOR U24387 ( .A(n24185), .B(n24184), .Z(c[91]) );
  XOR U24388 ( .A(n24183), .B(n24182), .Z(n24188) );
  NANDN U24389 ( .A(n24185), .B(n24184), .Z(n24186) );
  NANDN U24390 ( .A(n24187), .B(n24186), .Z(n24189) );
  XNOR U24391 ( .A(n24188), .B(n24189), .Z(c[92]) );
  NAND U24392 ( .A(n24189), .B(n24188), .Z(n24191) );
  AND U24393 ( .A(n24191), .B(n24190), .Z(n24195) );
  XOR U24394 ( .A(n24193), .B(n24192), .Z(n24194) );
  XNOR U24395 ( .A(n24195), .B(n24194), .Z(c[93]) );
  XOR U24396 ( .A(n24197), .B(n24196), .Z(c[94]) );
  XOR U24397 ( .A(n24199), .B(n24198), .Z(c[95]) );
  XOR U24398 ( .A(n24201), .B(n24200), .Z(c[96]) );
  XOR U24399 ( .A(n24203), .B(n24202), .Z(c[97]) );
  XNOR U24400 ( .A(n24205), .B(n24204), .Z(c[98]) );
  XOR U24401 ( .A(n24207), .B(n24206), .Z(c[99]) );
  XNOR U24402 ( .A(n24209), .B(n24208), .Z(c[100]) );
  XNOR U24403 ( .A(n24211), .B(n24210), .Z(n24212) );
  XOR U24404 ( .A(n24213), .B(n24212), .Z(c[101]) );
  XOR U24405 ( .A(n24215), .B(n24214), .Z(c[2]) );
  XNOR U24406 ( .A(n24217), .B(n24216), .Z(c[12]) );
  XNOR U24407 ( .A(n24219), .B(n24218), .Z(c[13]) );
  XOR U24408 ( .A(n24221), .B(n24220), .Z(c[14]) );
  XNOR U24409 ( .A(n24223), .B(n24222), .Z(c[15]) );
  XOR U24410 ( .A(n24225), .B(n24224), .Z(c[16]) );
  XNOR U24411 ( .A(n24227), .B(n24226), .Z(c[17]) );
  XOR U24412 ( .A(n24229), .B(n24228), .Z(c[18]) );
  XNOR U24413 ( .A(n24231), .B(n24230), .Z(c[19]) );
  XOR U24414 ( .A(n24233), .B(n24232), .Z(c[20]) );
  XNOR U24415 ( .A(n24235), .B(n24234), .Z(c[21]) );
  XOR U24416 ( .A(n24237), .B(n24236), .Z(c[3]) );
  XOR U24417 ( .A(n24239), .B(n24238), .Z(c[22]) );
  XNOR U24418 ( .A(n24241), .B(n24240), .Z(c[23]) );
  XOR U24419 ( .A(n24243), .B(n24242), .Z(c[24]) );
  XNOR U24420 ( .A(n24245), .B(n24244), .Z(c[25]) );
  XNOR U24421 ( .A(n24247), .B(n24246), .Z(c[26]) );
  XNOR U24422 ( .A(n24249), .B(n24248), .Z(c[27]) );
  XOR U24423 ( .A(n24251), .B(n24250), .Z(c[28]) );
  XNOR U24424 ( .A(n24253), .B(n24252), .Z(c[29]) );
  XNOR U24425 ( .A(n24255), .B(n24254), .Z(c[30]) );
  XNOR U24426 ( .A(n24257), .B(n24256), .Z(c[31]) );
  XNOR U24427 ( .A(n24259), .B(n24258), .Z(c[4]) );
  XOR U24428 ( .A(n24261), .B(n24260), .Z(c[32]) );
  XNOR U24429 ( .A(n24263), .B(n24262), .Z(c[33]) );
  XOR U24430 ( .A(n24265), .B(n24264), .Z(c[34]) );
  XNOR U24431 ( .A(n24267), .B(n24266), .Z(c[35]) );
  XOR U24432 ( .A(n24269), .B(n24268), .Z(c[36]) );
  XNOR U24433 ( .A(n24271), .B(n24270), .Z(c[37]) );
  XOR U24434 ( .A(n24273), .B(n24272), .Z(c[38]) );
  XNOR U24435 ( .A(n24275), .B(n24274), .Z(c[39]) );
  XOR U24436 ( .A(n24277), .B(n24276), .Z(c[40]) );
  XNOR U24437 ( .A(n24279), .B(n24278), .Z(c[41]) );
  XNOR U24438 ( .A(n24281), .B(n24280), .Z(c[5]) );
  XOR U24439 ( .A(n24283), .B(n24282), .Z(c[42]) );
  XNOR U24440 ( .A(n24285), .B(n24284), .Z(c[43]) );
  XOR U24441 ( .A(n24287), .B(n24286), .Z(c[44]) );
  XNOR U24442 ( .A(n24289), .B(n24288), .Z(c[45]) );
  XOR U24443 ( .A(n24291), .B(n24290), .Z(c[46]) );
  XNOR U24444 ( .A(n24293), .B(n24292), .Z(c[47]) );
  XOR U24445 ( .A(n24295), .B(n24294), .Z(c[48]) );
  XNOR U24446 ( .A(n24297), .B(n24296), .Z(c[49]) );
  XOR U24447 ( .A(n24299), .B(n24298), .Z(c[50]) );
  XNOR U24448 ( .A(n24301), .B(n24300), .Z(c[51]) );
  XOR U24449 ( .A(n24303), .B(n24302), .Z(c[6]) );
  XOR U24450 ( .A(n24305), .B(n24304), .Z(c[52]) );
  XNOR U24451 ( .A(n24307), .B(n24306), .Z(c[53]) );
  XOR U24452 ( .A(n24309), .B(n24308), .Z(c[54]) );
  XNOR U24453 ( .A(n24311), .B(n24310), .Z(c[55]) );
  XOR U24454 ( .A(n24313), .B(n24312), .Z(c[56]) );
  XNOR U24455 ( .A(n24315), .B(n24314), .Z(c[57]) );
  XOR U24456 ( .A(n24317), .B(n24316), .Z(c[58]) );
  XNOR U24457 ( .A(n24319), .B(n24318), .Z(c[59]) );
  XOR U24458 ( .A(n24321), .B(n24320), .Z(c[60]) );
  XNOR U24459 ( .A(n24323), .B(n24322), .Z(c[61]) );
  XOR U24460 ( .A(n24325), .B(n24324), .Z(c[7]) );
  XNOR U24461 ( .A(n24327), .B(n24326), .Z(c[62]) );
  XNOR U24462 ( .A(n24329), .B(n24328), .Z(c[63]) );
  XOR U24463 ( .A(n24331), .B(n24330), .Z(c[64]) );
  XNOR U24464 ( .A(n24333), .B(n24332), .Z(c[8]) );
  XNOR U24465 ( .A(n24335), .B(n24334), .Z(c[9]) );
  XNOR U24466 ( .A(n24337), .B(n24336), .Z(c[10]) );
  XNOR U24467 ( .A(n24339), .B(n24338), .Z(c[11]) );
  NAND U24468 ( .A(a[1]), .B(b[0]), .Z(n24340) );
  XNOR U24469 ( .A(n24341), .B(n24340), .Z(c[1]) );
endmodule

