
module stackMachine_N32 ( clk, rst, x, opcode, o );
  input [31:0] x;
  input [2:0] opcode;
  output [31:0] o;
  input clk, rst;
  wire   \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_1 , \C3/DATA5_3 , \C3/DATA5_4 , \C3/DATA5_5 ,
         \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 , \C3/DATA5_10 ,
         \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 , \C3/DATA5_14 ,
         \C3/DATA5_15 , \C3/DATA5_16 , \C3/DATA5_17 , \C3/DATA5_18 ,
         \C3/DATA5_19 , \C3/DATA5_20 , \C3/DATA5_21 , \C3/DATA5_22 ,
         \C3/DATA5_23 , \C3/DATA5_24 , \C3/DATA5_25 , \C3/DATA5_26 ,
         \C3/DATA5_27 , \C3/DATA5_28 , \C3/DATA5_29 , \C3/DATA5_30 ,
         \C3/DATA5_31 , n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, \C1/Z_0 ,
         \U1/RSOP_16/C3/Z_31 , \U1/RSOP_16/C3/Z_30 , \U1/RSOP_16/C3/Z_29 ,
         \U1/RSOP_16/C3/Z_28 , \U1/RSOP_16/C3/Z_27 , \U1/RSOP_16/C3/Z_26 ,
         \U1/RSOP_16/C3/Z_25 , \U1/RSOP_16/C3/Z_24 , \U1/RSOP_16/C3/Z_23 ,
         \U1/RSOP_16/C3/Z_22 , \U1/RSOP_16/C3/Z_21 , \U1/RSOP_16/C3/Z_20 ,
         \U1/RSOP_16/C3/Z_19 , \U1/RSOP_16/C3/Z_18 , \U1/RSOP_16/C3/Z_17 ,
         \U1/RSOP_16/C3/Z_16 , \U1/RSOP_16/C3/Z_15 , \U1/RSOP_16/C3/Z_14 ,
         \U1/RSOP_16/C3/Z_13 , \U1/RSOP_16/C3/Z_12 , \U1/RSOP_16/C3/Z_11 ,
         \U1/RSOP_16/C3/Z_10 , \U1/RSOP_16/C3/Z_9 , \U1/RSOP_16/C3/Z_8 ,
         \U1/RSOP_16/C3/Z_7 , \U1/RSOP_16/C3/Z_6 , \U1/RSOP_16/C3/Z_5 ,
         \U1/RSOP_16/C3/Z_4 , \U1/RSOP_16/C3/Z_3 , \U1/RSOP_16/C3/Z_2 ,
         \U1/RSOP_16/C3/Z_1 , \U1/RSOP_16/C3/Z_0 , \U1/RSOP_16/C2/Z_31 ,
         \U1/RSOP_16/C2/Z_30 , \U1/RSOP_16/C2/Z_29 , \U1/RSOP_16/C2/Z_28 ,
         \U1/RSOP_16/C2/Z_27 , \U1/RSOP_16/C2/Z_26 , \U1/RSOP_16/C2/Z_25 ,
         \U1/RSOP_16/C2/Z_24 , \U1/RSOP_16/C2/Z_23 , \U1/RSOP_16/C2/Z_22 ,
         \U1/RSOP_16/C2/Z_21 , \U1/RSOP_16/C2/Z_20 , \U1/RSOP_16/C2/Z_19 ,
         \U1/RSOP_16/C2/Z_18 , \U1/RSOP_16/C2/Z_17 , \U1/RSOP_16/C2/Z_16 ,
         \U1/RSOP_16/C2/Z_15 , \U1/RSOP_16/C2/Z_14 , \U1/RSOP_16/C2/Z_13 ,
         \U1/RSOP_16/C2/Z_12 , \U1/RSOP_16/C2/Z_11 , \U1/RSOP_16/C2/Z_10 ,
         \U1/RSOP_16/C2/Z_9 , \U1/RSOP_16/C2/Z_8 , \U1/RSOP_16/C2/Z_7 ,
         \U1/RSOP_16/C2/Z_6 , \U1/RSOP_16/C2/Z_5 , \U1/RSOP_16/C2/Z_4 ,
         \U1/RSOP_16/C2/Z_3 , \U1/RSOP_16/C2/Z_2 , \U1/RSOP_16/C2/Z_1 ,
         \U1/RSOP_16/C2/Z_0 , \DP_OP_25_64_5665/n336 , \DP_OP_25_64_5665/n335 ,
         \DP_OP_25_64_5665/n334 , \DP_OP_25_64_5665/n333 ,
         \DP_OP_25_64_5665/n332 , \DP_OP_25_64_5665/n331 ,
         \DP_OP_25_64_5665/n330 , \DP_OP_25_64_5665/n329 ,
         \DP_OP_25_64_5665/n328 , \DP_OP_25_64_5665/n327 ,
         \DP_OP_25_64_5665/n326 , \DP_OP_25_64_5665/n325 ,
         \DP_OP_25_64_5665/n324 , \DP_OP_25_64_5665/n323 ,
         \DP_OP_25_64_5665/n322 , \DP_OP_25_64_5665/n321 ,
         \DP_OP_25_64_5665/n320 , \DP_OP_25_64_5665/n319 ,
         \DP_OP_25_64_5665/n318 , \DP_OP_25_64_5665/n317 ,
         \DP_OP_25_64_5665/n316 , \DP_OP_25_64_5665/n315 ,
         \DP_OP_25_64_5665/n314 , \DP_OP_25_64_5665/n313 ,
         \DP_OP_25_64_5665/n312 , \DP_OP_25_64_5665/n311 ,
         \DP_OP_25_64_5665/n310 , \DP_OP_25_64_5665/n309 ,
         \DP_OP_25_64_5665/n308 , \DP_OP_25_64_5665/n307 ,
         \DP_OP_25_64_5665/n306 , \DP_OP_25_64_5665/n305 ,
         \DP_OP_25_64_5665/n300 , \DP_OP_25_64_5665/n299 ,
         \DP_OP_25_64_5665/n298 , \DP_OP_25_64_5665/n297 ,
         \DP_OP_25_64_5665/n296 , \DP_OP_25_64_5665/n295 ,
         \DP_OP_25_64_5665/n294 , \DP_OP_25_64_5665/n293 ,
         \DP_OP_25_64_5665/n292 , \DP_OP_25_64_5665/n291 ,
         \DP_OP_25_64_5665/n290 , \DP_OP_25_64_5665/n289 ,
         \DP_OP_25_64_5665/n288 , \DP_OP_25_64_5665/n287 ,
         \DP_OP_25_64_5665/n286 , \DP_OP_25_64_5665/n285 ,
         \DP_OP_25_64_5665/n284 , \DP_OP_25_64_5665/n283 ,
         \DP_OP_25_64_5665/n282 , \DP_OP_25_64_5665/n281 ,
         \DP_OP_25_64_5665/n280 , \DP_OP_25_64_5665/n279 ,
         \DP_OP_25_64_5665/n278 , \DP_OP_25_64_5665/n277 ,
         \DP_OP_25_64_5665/n276 , \DP_OP_25_64_5665/n275 ,
         \DP_OP_25_64_5665/n274 , \DP_OP_25_64_5665/n273 ,
         \DP_OP_25_64_5665/n272 , \DP_OP_25_64_5665/n271 ,
         \DP_OP_25_64_5665/n270 , \DP_OP_25_64_5665/n269 ,
         \DP_OP_25_64_5665/n268 , \DP_OP_25_64_5665/n267 ,
         \DP_OP_25_64_5665/n266 , \DP_OP_25_64_5665/n265 ,
         \DP_OP_25_64_5665/n264 , \DP_OP_25_64_5665/n263 ,
         \DP_OP_25_64_5665/n262 , \DP_OP_25_64_5665/n261 ,
         \DP_OP_25_64_5665/n260 , \DP_OP_25_64_5665/n259 ,
         \DP_OP_25_64_5665/n258 , \DP_OP_25_64_5665/n257 ,
         \DP_OP_25_64_5665/n256 , \DP_OP_25_64_5665/n255 ,
         \DP_OP_25_64_5665/n254 , \DP_OP_25_64_5665/n253 ,
         \DP_OP_25_64_5665/n252 , \DP_OP_25_64_5665/n251 ,
         \DP_OP_25_64_5665/n250 , \DP_OP_25_64_5665/n249 ,
         \DP_OP_25_64_5665/n248 , \DP_OP_25_64_5665/n247 ,
         \DP_OP_25_64_5665/n246 , \DP_OP_25_64_5665/n245 ,
         \DP_OP_25_64_5665/n244 , \DP_OP_25_64_5665/n243 ,
         \DP_OP_25_64_5665/n242 , \DP_OP_25_64_5665/n241 ,
         \DP_OP_25_64_5665/n240 , \DP_OP_25_64_5665/n239 ,
         \DP_OP_25_64_5665/n238 , \DP_OP_25_64_5665/n236 ,
         \DP_OP_25_64_5665/n235 , \DP_OP_25_64_5665/n229 ,
         \DP_OP_25_64_5665/n228 , \DP_OP_25_64_5665/n222 ,
         \DP_OP_25_64_5665/n221 , \DP_OP_25_64_5665/n215 ,
         \DP_OP_25_64_5665/n214 , \DP_OP_25_64_5665/n208 ,
         \DP_OP_25_64_5665/n207 , \DP_OP_25_64_5665/n201 ,
         \DP_OP_25_64_5665/n200 , \DP_OP_25_64_5665/n194 ,
         \DP_OP_25_64_5665/n193 , \DP_OP_25_64_5665/n187 ,
         \DP_OP_25_64_5665/n186 , \DP_OP_25_64_5665/n180 ,
         \DP_OP_25_64_5665/n179 , \DP_OP_25_64_5665/n173 ,
         \DP_OP_25_64_5665/n172 , \DP_OP_25_64_5665/n166 ,
         \DP_OP_25_64_5665/n165 , \DP_OP_25_64_5665/n159 ,
         \DP_OP_25_64_5665/n158 , \DP_OP_25_64_5665/n152 ,
         \DP_OP_25_64_5665/n151 , \DP_OP_25_64_5665/n145 ,
         \DP_OP_25_64_5665/n144 , \DP_OP_25_64_5665/n138 ,
         \DP_OP_25_64_5665/n137 , \DP_OP_25_64_5665/n131 ,
         \DP_OP_25_64_5665/n130 , \DP_OP_25_64_5665/n124 ,
         \DP_OP_25_64_5665/n123 , \DP_OP_25_64_5665/n117 ,
         \DP_OP_25_64_5665/n116 , \DP_OP_25_64_5665/n110 ,
         \DP_OP_25_64_5665/n109 , \DP_OP_25_64_5665/n103 ,
         \DP_OP_25_64_5665/n102 , \DP_OP_25_64_5665/n96 ,
         \DP_OP_25_64_5665/n95 , \DP_OP_25_64_5665/n89 ,
         \DP_OP_25_64_5665/n88 , \DP_OP_25_64_5665/n82 ,
         \DP_OP_25_64_5665/n81 , \DP_OP_25_64_5665/n57 ,
         \DP_OP_25_64_5665/n56 , \DP_OP_25_64_5665/n50 ,
         \DP_OP_25_64_5665/n49 , \DP_OP_25_64_5665/n43 ,
         \DP_OP_25_64_5665/n42 , \DP_OP_25_64_5665/n36 ,
         \DP_OP_25_64_5665/n35 , \DP_OP_25_64_5665/n29 ,
         \DP_OP_25_64_5665/n28 , \DP_OP_25_64_5665/n22 ,
         \DP_OP_25_64_5665/n21 , \DP_OP_25_64_5665/n15 ,
         \DP_OP_25_64_5665/n14 , \DP_OP_25_64_5665/n8 , \DP_OP_25_64_5665/n5 ,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606;

  DFF \stack_reg[0][0]  ( .D(n1318), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n1317), .CLK(clk), .RST(rst), .Q(\stack[1][0] )
         );
  DFF \stack_reg[0][1]  ( .D(n1316), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n1315), .CLK(clk), .RST(rst), .Q(\stack[1][1] )
         );
  DFF \stack_reg[2][1]  ( .D(n1314), .CLK(clk), .RST(rst), .Q(\stack[2][1] )
         );
  DFF \stack_reg[3][1]  ( .D(n1313), .CLK(clk), .RST(rst), .Q(\stack[3][1] )
         );
  DFF \stack_reg[4][1]  ( .D(n1312), .CLK(clk), .RST(rst), .Q(\stack[4][1] )
         );
  DFF \stack_reg[5][1]  ( .D(n1311), .CLK(clk), .RST(rst), .Q(\stack[5][1] )
         );
  DFF \stack_reg[6][1]  ( .D(n1310), .CLK(clk), .RST(rst), .Q(\stack[6][1] )
         );
  DFF \stack_reg[7][1]  ( .D(n1309), .CLK(clk), .RST(rst), .Q(\stack[7][1] )
         );
  DFF \stack_reg[0][2]  ( .D(n1308), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n1307), .CLK(clk), .RST(rst), .Q(\stack[1][2] )
         );
  DFF \stack_reg[2][2]  ( .D(n1306), .CLK(clk), .RST(rst), .Q(\stack[2][2] )
         );
  DFF \stack_reg[3][2]  ( .D(n1305), .CLK(clk), .RST(rst), .Q(\stack[3][2] )
         );
  DFF \stack_reg[4][2]  ( .D(n1304), .CLK(clk), .RST(rst), .Q(\stack[4][2] )
         );
  DFF \stack_reg[5][2]  ( .D(n1303), .CLK(clk), .RST(rst), .Q(\stack[5][2] )
         );
  DFF \stack_reg[6][2]  ( .D(n1302), .CLK(clk), .RST(rst), .Q(\stack[6][2] )
         );
  DFF \stack_reg[7][2]  ( .D(n1301), .CLK(clk), .RST(rst), .Q(\stack[7][2] )
         );
  DFF \stack_reg[0][3]  ( .D(n1300), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n1299), .CLK(clk), .RST(rst), .Q(\stack[1][3] )
         );
  DFF \stack_reg[2][3]  ( .D(n1298), .CLK(clk), .RST(rst), .Q(\stack[2][3] )
         );
  DFF \stack_reg[3][3]  ( .D(n1297), .CLK(clk), .RST(rst), .Q(\stack[3][3] )
         );
  DFF \stack_reg[4][3]  ( .D(n1296), .CLK(clk), .RST(rst), .Q(\stack[4][3] )
         );
  DFF \stack_reg[5][3]  ( .D(n1295), .CLK(clk), .RST(rst), .Q(\stack[5][3] )
         );
  DFF \stack_reg[6][3]  ( .D(n1294), .CLK(clk), .RST(rst), .Q(\stack[6][3] )
         );
  DFF \stack_reg[7][3]  ( .D(n1293), .CLK(clk), .RST(rst), .Q(\stack[7][3] )
         );
  DFF \stack_reg[0][4]  ( .D(n1292), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n1291), .CLK(clk), .RST(rst), .Q(\stack[1][4] )
         );
  DFF \stack_reg[2][4]  ( .D(n1290), .CLK(clk), .RST(rst), .Q(\stack[2][4] )
         );
  DFF \stack_reg[3][4]  ( .D(n1289), .CLK(clk), .RST(rst), .Q(\stack[3][4] )
         );
  DFF \stack_reg[4][4]  ( .D(n1288), .CLK(clk), .RST(rst), .Q(\stack[4][4] )
         );
  DFF \stack_reg[5][4]  ( .D(n1287), .CLK(clk), .RST(rst), .Q(\stack[5][4] )
         );
  DFF \stack_reg[6][4]  ( .D(n1286), .CLK(clk), .RST(rst), .Q(\stack[6][4] )
         );
  DFF \stack_reg[7][4]  ( .D(n1285), .CLK(clk), .RST(rst), .Q(\stack[7][4] )
         );
  DFF \stack_reg[0][5]  ( .D(n1284), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n1283), .CLK(clk), .RST(rst), .Q(\stack[1][5] )
         );
  DFF \stack_reg[2][5]  ( .D(n1282), .CLK(clk), .RST(rst), .Q(\stack[2][5] )
         );
  DFF \stack_reg[3][5]  ( .D(n1281), .CLK(clk), .RST(rst), .Q(\stack[3][5] )
         );
  DFF \stack_reg[4][5]  ( .D(n1280), .CLK(clk), .RST(rst), .Q(\stack[4][5] )
         );
  DFF \stack_reg[5][5]  ( .D(n1279), .CLK(clk), .RST(rst), .Q(\stack[5][5] )
         );
  DFF \stack_reg[6][5]  ( .D(n1278), .CLK(clk), .RST(rst), .Q(\stack[6][5] )
         );
  DFF \stack_reg[7][5]  ( .D(n1277), .CLK(clk), .RST(rst), .Q(\stack[7][5] )
         );
  DFF \stack_reg[0][6]  ( .D(n1276), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n1275), .CLK(clk), .RST(rst), .Q(\stack[1][6] )
         );
  DFF \stack_reg[2][6]  ( .D(n1274), .CLK(clk), .RST(rst), .Q(\stack[2][6] )
         );
  DFF \stack_reg[3][6]  ( .D(n1273), .CLK(clk), .RST(rst), .Q(\stack[3][6] )
         );
  DFF \stack_reg[4][6]  ( .D(n1272), .CLK(clk), .RST(rst), .Q(\stack[4][6] )
         );
  DFF \stack_reg[5][6]  ( .D(n1271), .CLK(clk), .RST(rst), .Q(\stack[5][6] )
         );
  DFF \stack_reg[6][6]  ( .D(n1270), .CLK(clk), .RST(rst), .Q(\stack[6][6] )
         );
  DFF \stack_reg[7][6]  ( .D(n1269), .CLK(clk), .RST(rst), .Q(\stack[7][6] )
         );
  DFF \stack_reg[0][7]  ( .D(n1268), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n1267), .CLK(clk), .RST(rst), .Q(\stack[1][7] )
         );
  DFF \stack_reg[2][7]  ( .D(n1266), .CLK(clk), .RST(rst), .Q(\stack[2][7] )
         );
  DFF \stack_reg[3][7]  ( .D(n1265), .CLK(clk), .RST(rst), .Q(\stack[3][7] )
         );
  DFF \stack_reg[4][7]  ( .D(n1264), .CLK(clk), .RST(rst), .Q(\stack[4][7] )
         );
  DFF \stack_reg[5][7]  ( .D(n1263), .CLK(clk), .RST(rst), .Q(\stack[5][7] )
         );
  DFF \stack_reg[6][7]  ( .D(n1262), .CLK(clk), .RST(rst), .Q(\stack[6][7] )
         );
  DFF \stack_reg[7][7]  ( .D(n1261), .CLK(clk), .RST(rst), .Q(\stack[7][7] )
         );
  DFF \stack_reg[0][8]  ( .D(n1260), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n1259), .CLK(clk), .RST(rst), .Q(\stack[1][8] )
         );
  DFF \stack_reg[2][8]  ( .D(n1258), .CLK(clk), .RST(rst), .Q(\stack[2][8] )
         );
  DFF \stack_reg[3][8]  ( .D(n1257), .CLK(clk), .RST(rst), .Q(\stack[3][8] )
         );
  DFF \stack_reg[4][8]  ( .D(n1256), .CLK(clk), .RST(rst), .Q(\stack[4][8] )
         );
  DFF \stack_reg[5][8]  ( .D(n1255), .CLK(clk), .RST(rst), .Q(\stack[5][8] )
         );
  DFF \stack_reg[6][8]  ( .D(n1254), .CLK(clk), .RST(rst), .Q(\stack[6][8] )
         );
  DFF \stack_reg[7][8]  ( .D(n1253), .CLK(clk), .RST(rst), .Q(\stack[7][8] )
         );
  DFF \stack_reg[0][9]  ( .D(n1252), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n1251), .CLK(clk), .RST(rst), .Q(\stack[1][9] )
         );
  DFF \stack_reg[2][9]  ( .D(n1250), .CLK(clk), .RST(rst), .Q(\stack[2][9] )
         );
  DFF \stack_reg[3][9]  ( .D(n1249), .CLK(clk), .RST(rst), .Q(\stack[3][9] )
         );
  DFF \stack_reg[4][9]  ( .D(n1248), .CLK(clk), .RST(rst), .Q(\stack[4][9] )
         );
  DFF \stack_reg[5][9]  ( .D(n1247), .CLK(clk), .RST(rst), .Q(\stack[5][9] )
         );
  DFF \stack_reg[6][9]  ( .D(n1246), .CLK(clk), .RST(rst), .Q(\stack[6][9] )
         );
  DFF \stack_reg[7][9]  ( .D(n1245), .CLK(clk), .RST(rst), .Q(\stack[7][9] )
         );
  DFF \stack_reg[0][10]  ( .D(n1244), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n1243), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n1242), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n1241), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n1240), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n1239), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n1238), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n1237), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n1236), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n1235), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n1234), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n1233), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n1232), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n1231), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n1230), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n1229), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n1228), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n1227), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n1226), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n1225), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n1224), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n1223), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n1222), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n1221), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n1220), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n1219), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n1218), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n1217), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n1216), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n1215), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n1214), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n1213), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n1212), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n1211), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n1210), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n1209), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n1208), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n1207), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n1206), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n1205), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n1204), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n1203), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n1202), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n1201), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n1200), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n1199), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n1198), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n1197), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[0][16]  ( .D(n1196), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \stack_reg[1][16]  ( .D(n1195), .CLK(clk), .RST(rst), .Q(\stack[1][16] )
         );
  DFF \stack_reg[2][16]  ( .D(n1194), .CLK(clk), .RST(rst), .Q(\stack[2][16] )
         );
  DFF \stack_reg[3][16]  ( .D(n1193), .CLK(clk), .RST(rst), .Q(\stack[3][16] )
         );
  DFF \stack_reg[4][16]  ( .D(n1192), .CLK(clk), .RST(rst), .Q(\stack[4][16] )
         );
  DFF \stack_reg[5][16]  ( .D(n1191), .CLK(clk), .RST(rst), .Q(\stack[5][16] )
         );
  DFF \stack_reg[6][16]  ( .D(n1190), .CLK(clk), .RST(rst), .Q(\stack[6][16] )
         );
  DFF \stack_reg[7][16]  ( .D(n1189), .CLK(clk), .RST(rst), .Q(\stack[7][16] )
         );
  DFF \stack_reg[0][17]  ( .D(n1188), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \stack_reg[1][17]  ( .D(n1187), .CLK(clk), .RST(rst), .Q(\stack[1][17] )
         );
  DFF \stack_reg[2][17]  ( .D(n1186), .CLK(clk), .RST(rst), .Q(\stack[2][17] )
         );
  DFF \stack_reg[3][17]  ( .D(n1185), .CLK(clk), .RST(rst), .Q(\stack[3][17] )
         );
  DFF \stack_reg[4][17]  ( .D(n1184), .CLK(clk), .RST(rst), .Q(\stack[4][17] )
         );
  DFF \stack_reg[5][17]  ( .D(n1183), .CLK(clk), .RST(rst), .Q(\stack[5][17] )
         );
  DFF \stack_reg[6][17]  ( .D(n1182), .CLK(clk), .RST(rst), .Q(\stack[6][17] )
         );
  DFF \stack_reg[7][17]  ( .D(n1181), .CLK(clk), .RST(rst), .Q(\stack[7][17] )
         );
  DFF \stack_reg[0][18]  ( .D(n1180), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \stack_reg[1][18]  ( .D(n1179), .CLK(clk), .RST(rst), .Q(\stack[1][18] )
         );
  DFF \stack_reg[2][18]  ( .D(n1178), .CLK(clk), .RST(rst), .Q(\stack[2][18] )
         );
  DFF \stack_reg[3][18]  ( .D(n1177), .CLK(clk), .RST(rst), .Q(\stack[3][18] )
         );
  DFF \stack_reg[4][18]  ( .D(n1176), .CLK(clk), .RST(rst), .Q(\stack[4][18] )
         );
  DFF \stack_reg[5][18]  ( .D(n1175), .CLK(clk), .RST(rst), .Q(\stack[5][18] )
         );
  DFF \stack_reg[6][18]  ( .D(n1174), .CLK(clk), .RST(rst), .Q(\stack[6][18] )
         );
  DFF \stack_reg[7][18]  ( .D(n1173), .CLK(clk), .RST(rst), .Q(\stack[7][18] )
         );
  DFF \stack_reg[0][19]  ( .D(n1172), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \stack_reg[1][19]  ( .D(n1171), .CLK(clk), .RST(rst), .Q(\stack[1][19] )
         );
  DFF \stack_reg[2][19]  ( .D(n1170), .CLK(clk), .RST(rst), .Q(\stack[2][19] )
         );
  DFF \stack_reg[3][19]  ( .D(n1169), .CLK(clk), .RST(rst), .Q(\stack[3][19] )
         );
  DFF \stack_reg[4][19]  ( .D(n1168), .CLK(clk), .RST(rst), .Q(\stack[4][19] )
         );
  DFF \stack_reg[5][19]  ( .D(n1167), .CLK(clk), .RST(rst), .Q(\stack[5][19] )
         );
  DFF \stack_reg[6][19]  ( .D(n1166), .CLK(clk), .RST(rst), .Q(\stack[6][19] )
         );
  DFF \stack_reg[7][19]  ( .D(n1165), .CLK(clk), .RST(rst), .Q(\stack[7][19] )
         );
  DFF \stack_reg[0][20]  ( .D(n1164), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \stack_reg[1][20]  ( .D(n1163), .CLK(clk), .RST(rst), .Q(\stack[1][20] )
         );
  DFF \stack_reg[2][20]  ( .D(n1162), .CLK(clk), .RST(rst), .Q(\stack[2][20] )
         );
  DFF \stack_reg[3][20]  ( .D(n1161), .CLK(clk), .RST(rst), .Q(\stack[3][20] )
         );
  DFF \stack_reg[4][20]  ( .D(n1160), .CLK(clk), .RST(rst), .Q(\stack[4][20] )
         );
  DFF \stack_reg[5][20]  ( .D(n1159), .CLK(clk), .RST(rst), .Q(\stack[5][20] )
         );
  DFF \stack_reg[6][20]  ( .D(n1158), .CLK(clk), .RST(rst), .Q(\stack[6][20] )
         );
  DFF \stack_reg[7][20]  ( .D(n1157), .CLK(clk), .RST(rst), .Q(\stack[7][20] )
         );
  DFF \stack_reg[0][21]  ( .D(n1156), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \stack_reg[1][21]  ( .D(n1155), .CLK(clk), .RST(rst), .Q(\stack[1][21] )
         );
  DFF \stack_reg[2][21]  ( .D(n1154), .CLK(clk), .RST(rst), .Q(\stack[2][21] )
         );
  DFF \stack_reg[3][21]  ( .D(n1153), .CLK(clk), .RST(rst), .Q(\stack[3][21] )
         );
  DFF \stack_reg[4][21]  ( .D(n1152), .CLK(clk), .RST(rst), .Q(\stack[4][21] )
         );
  DFF \stack_reg[5][21]  ( .D(n1151), .CLK(clk), .RST(rst), .Q(\stack[5][21] )
         );
  DFF \stack_reg[6][21]  ( .D(n1150), .CLK(clk), .RST(rst), .Q(\stack[6][21] )
         );
  DFF \stack_reg[7][21]  ( .D(n1149), .CLK(clk), .RST(rst), .Q(\stack[7][21] )
         );
  DFF \stack_reg[0][22]  ( .D(n1148), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \stack_reg[1][22]  ( .D(n1147), .CLK(clk), .RST(rst), .Q(\stack[1][22] )
         );
  DFF \stack_reg[2][22]  ( .D(n1146), .CLK(clk), .RST(rst), .Q(\stack[2][22] )
         );
  DFF \stack_reg[3][22]  ( .D(n1145), .CLK(clk), .RST(rst), .Q(\stack[3][22] )
         );
  DFF \stack_reg[4][22]  ( .D(n1144), .CLK(clk), .RST(rst), .Q(\stack[4][22] )
         );
  DFF \stack_reg[5][22]  ( .D(n1143), .CLK(clk), .RST(rst), .Q(\stack[5][22] )
         );
  DFF \stack_reg[6][22]  ( .D(n1142), .CLK(clk), .RST(rst), .Q(\stack[6][22] )
         );
  DFF \stack_reg[7][22]  ( .D(n1141), .CLK(clk), .RST(rst), .Q(\stack[7][22] )
         );
  DFF \stack_reg[0][23]  ( .D(n1140), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \stack_reg[1][23]  ( .D(n1139), .CLK(clk), .RST(rst), .Q(\stack[1][23] )
         );
  DFF \stack_reg[2][23]  ( .D(n1138), .CLK(clk), .RST(rst), .Q(\stack[2][23] )
         );
  DFF \stack_reg[3][23]  ( .D(n1137), .CLK(clk), .RST(rst), .Q(\stack[3][23] )
         );
  DFF \stack_reg[4][23]  ( .D(n1136), .CLK(clk), .RST(rst), .Q(\stack[4][23] )
         );
  DFF \stack_reg[5][23]  ( .D(n1135), .CLK(clk), .RST(rst), .Q(\stack[5][23] )
         );
  DFF \stack_reg[6][23]  ( .D(n1134), .CLK(clk), .RST(rst), .Q(\stack[6][23] )
         );
  DFF \stack_reg[7][23]  ( .D(n1133), .CLK(clk), .RST(rst), .Q(\stack[7][23] )
         );
  DFF \stack_reg[0][24]  ( .D(n1132), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \stack_reg[1][24]  ( .D(n1131), .CLK(clk), .RST(rst), .Q(\stack[1][24] )
         );
  DFF \stack_reg[2][24]  ( .D(n1130), .CLK(clk), .RST(rst), .Q(\stack[2][24] )
         );
  DFF \stack_reg[3][24]  ( .D(n1129), .CLK(clk), .RST(rst), .Q(\stack[3][24] )
         );
  DFF \stack_reg[4][24]  ( .D(n1128), .CLK(clk), .RST(rst), .Q(\stack[4][24] )
         );
  DFF \stack_reg[5][24]  ( .D(n1127), .CLK(clk), .RST(rst), .Q(\stack[5][24] )
         );
  DFF \stack_reg[6][24]  ( .D(n1126), .CLK(clk), .RST(rst), .Q(\stack[6][24] )
         );
  DFF \stack_reg[7][24]  ( .D(n1125), .CLK(clk), .RST(rst), .Q(\stack[7][24] )
         );
  DFF \stack_reg[0][25]  ( .D(n1124), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \stack_reg[1][25]  ( .D(n1123), .CLK(clk), .RST(rst), .Q(\stack[1][25] )
         );
  DFF \stack_reg[2][25]  ( .D(n1122), .CLK(clk), .RST(rst), .Q(\stack[2][25] )
         );
  DFF \stack_reg[3][25]  ( .D(n1121), .CLK(clk), .RST(rst), .Q(\stack[3][25] )
         );
  DFF \stack_reg[4][25]  ( .D(n1120), .CLK(clk), .RST(rst), .Q(\stack[4][25] )
         );
  DFF \stack_reg[5][25]  ( .D(n1119), .CLK(clk), .RST(rst), .Q(\stack[5][25] )
         );
  DFF \stack_reg[6][25]  ( .D(n1118), .CLK(clk), .RST(rst), .Q(\stack[6][25] )
         );
  DFF \stack_reg[7][25]  ( .D(n1117), .CLK(clk), .RST(rst), .Q(\stack[7][25] )
         );
  DFF \stack_reg[0][26]  ( .D(n1116), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \stack_reg[1][26]  ( .D(n1115), .CLK(clk), .RST(rst), .Q(\stack[1][26] )
         );
  DFF \stack_reg[2][26]  ( .D(n1114), .CLK(clk), .RST(rst), .Q(\stack[2][26] )
         );
  DFF \stack_reg[3][26]  ( .D(n1113), .CLK(clk), .RST(rst), .Q(\stack[3][26] )
         );
  DFF \stack_reg[4][26]  ( .D(n1112), .CLK(clk), .RST(rst), .Q(\stack[4][26] )
         );
  DFF \stack_reg[5][26]  ( .D(n1111), .CLK(clk), .RST(rst), .Q(\stack[5][26] )
         );
  DFF \stack_reg[6][26]  ( .D(n1110), .CLK(clk), .RST(rst), .Q(\stack[6][26] )
         );
  DFF \stack_reg[7][26]  ( .D(n1109), .CLK(clk), .RST(rst), .Q(\stack[7][26] )
         );
  DFF \stack_reg[0][27]  ( .D(n1108), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \stack_reg[1][27]  ( .D(n1107), .CLK(clk), .RST(rst), .Q(\stack[1][27] )
         );
  DFF \stack_reg[2][27]  ( .D(n1106), .CLK(clk), .RST(rst), .Q(\stack[2][27] )
         );
  DFF \stack_reg[3][27]  ( .D(n1105), .CLK(clk), .RST(rst), .Q(\stack[3][27] )
         );
  DFF \stack_reg[4][27]  ( .D(n1104), .CLK(clk), .RST(rst), .Q(\stack[4][27] )
         );
  DFF \stack_reg[5][27]  ( .D(n1103), .CLK(clk), .RST(rst), .Q(\stack[5][27] )
         );
  DFF \stack_reg[6][27]  ( .D(n1102), .CLK(clk), .RST(rst), .Q(\stack[6][27] )
         );
  DFF \stack_reg[7][27]  ( .D(n1101), .CLK(clk), .RST(rst), .Q(\stack[7][27] )
         );
  DFF \stack_reg[0][28]  ( .D(n1100), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \stack_reg[1][28]  ( .D(n1099), .CLK(clk), .RST(rst), .Q(\stack[1][28] )
         );
  DFF \stack_reg[2][28]  ( .D(n1098), .CLK(clk), .RST(rst), .Q(\stack[2][28] )
         );
  DFF \stack_reg[3][28]  ( .D(n1097), .CLK(clk), .RST(rst), .Q(\stack[3][28] )
         );
  DFF \stack_reg[4][28]  ( .D(n1096), .CLK(clk), .RST(rst), .Q(\stack[4][28] )
         );
  DFF \stack_reg[5][28]  ( .D(n1095), .CLK(clk), .RST(rst), .Q(\stack[5][28] )
         );
  DFF \stack_reg[6][28]  ( .D(n1094), .CLK(clk), .RST(rst), .Q(\stack[6][28] )
         );
  DFF \stack_reg[7][28]  ( .D(n1093), .CLK(clk), .RST(rst), .Q(\stack[7][28] )
         );
  DFF \stack_reg[0][29]  ( .D(n1092), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \stack_reg[1][29]  ( .D(n1091), .CLK(clk), .RST(rst), .Q(\stack[1][29] )
         );
  DFF \stack_reg[2][29]  ( .D(n1090), .CLK(clk), .RST(rst), .Q(\stack[2][29] )
         );
  DFF \stack_reg[3][29]  ( .D(n1089), .CLK(clk), .RST(rst), .Q(\stack[3][29] )
         );
  DFF \stack_reg[4][29]  ( .D(n1088), .CLK(clk), .RST(rst), .Q(\stack[4][29] )
         );
  DFF \stack_reg[5][29]  ( .D(n1087), .CLK(clk), .RST(rst), .Q(\stack[5][29] )
         );
  DFF \stack_reg[6][29]  ( .D(n1086), .CLK(clk), .RST(rst), .Q(\stack[6][29] )
         );
  DFF \stack_reg[7][29]  ( .D(n1085), .CLK(clk), .RST(rst), .Q(\stack[7][29] )
         );
  DFF \stack_reg[0][30]  ( .D(n1084), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \stack_reg[1][30]  ( .D(n1083), .CLK(clk), .RST(rst), .Q(\stack[1][30] )
         );
  DFF \stack_reg[2][30]  ( .D(n1082), .CLK(clk), .RST(rst), .Q(\stack[2][30] )
         );
  DFF \stack_reg[3][30]  ( .D(n1081), .CLK(clk), .RST(rst), .Q(\stack[3][30] )
         );
  DFF \stack_reg[4][30]  ( .D(n1080), .CLK(clk), .RST(rst), .Q(\stack[4][30] )
         );
  DFF \stack_reg[5][30]  ( .D(n1079), .CLK(clk), .RST(rst), .Q(\stack[5][30] )
         );
  DFF \stack_reg[6][30]  ( .D(n1078), .CLK(clk), .RST(rst), .Q(\stack[6][30] )
         );
  DFF \stack_reg[7][30]  ( .D(n1077), .CLK(clk), .RST(rst), .Q(\stack[7][30] )
         );
  DFF \stack_reg[0][31]  ( .D(n1076), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \stack_reg[1][31]  ( .D(n1075), .CLK(clk), .RST(rst), .Q(\stack[1][31] )
         );
  DFF \stack_reg[2][31]  ( .D(n1074), .CLK(clk), .RST(rst), .Q(\stack[2][31] )
         );
  DFF \stack_reg[3][31]  ( .D(n1073), .CLK(clk), .RST(rst), .Q(\stack[3][31] )
         );
  DFF \stack_reg[4][31]  ( .D(n1072), .CLK(clk), .RST(rst), .Q(\stack[4][31] )
         );
  DFF \stack_reg[5][31]  ( .D(n1071), .CLK(clk), .RST(rst), .Q(\stack[5][31] )
         );
  DFF \stack_reg[6][31]  ( .D(n1070), .CLK(clk), .RST(rst), .Q(\stack[6][31] )
         );
  DFF \stack_reg[7][31]  ( .D(n1069), .CLK(clk), .RST(rst), .Q(\stack[7][31] )
         );
  DFF \stack_reg[2][0]  ( .D(n1068), .CLK(clk), .RST(rst), .Q(\stack[2][0] )
         );
  DFF \stack_reg[3][0]  ( .D(n1067), .CLK(clk), .RST(rst), .Q(\stack[3][0] )
         );
  DFF \stack_reg[4][0]  ( .D(n1066), .CLK(clk), .RST(rst), .Q(\stack[4][0] )
         );
  DFF \stack_reg[5][0]  ( .D(n1065), .CLK(clk), .RST(rst), .Q(\stack[5][0] )
         );
  DFF \stack_reg[6][0]  ( .D(n1064), .CLK(clk), .RST(rst), .Q(\stack[6][0] )
         );
  DFF \stack_reg[7][0]  ( .D(n1063), .CLK(clk), .RST(rst), .Q(\stack[7][0] )
         );
  XOR \DP_OP_25_64_5665/U149  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_5665/n336 ) );
  XOR \DP_OP_25_64_5665/U148  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_5665/n335 ) );
  XOR \DP_OP_25_64_5665/U147  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_5665/n334 ) );
  XOR \DP_OP_25_64_5665/U146  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_5665/n333 ) );
  XOR \DP_OP_25_64_5665/U145  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_5665/n332 ) );
  XOR \DP_OP_25_64_5665/U144  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_5665/n331 ) );
  XOR \DP_OP_25_64_5665/U143  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_5665/n330 ) );
  XOR \DP_OP_25_64_5665/U142  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_5665/n329 ) );
  XOR \DP_OP_25_64_5665/U141  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_5665/n328 ) );
  XOR \DP_OP_25_64_5665/U140  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_5665/n327 ) );
  XOR \DP_OP_25_64_5665/U139  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_5665/n326 ) );
  XOR \DP_OP_25_64_5665/U138  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_5665/n325 ) );
  XOR \DP_OP_25_64_5665/U137  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_5665/n324 ) );
  XOR \DP_OP_25_64_5665/U136  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_5665/n323 ) );
  XOR \DP_OP_25_64_5665/U135  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_5665/n322 ) );
  XOR \DP_OP_25_64_5665/U134  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_5665/n321 ) );
  XOR \DP_OP_25_64_5665/U133  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_16 ), .Z(
        \DP_OP_25_64_5665/n320 ) );
  XOR \DP_OP_25_64_5665/U132  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_17 ), .Z(
        \DP_OP_25_64_5665/n319 ) );
  XOR \DP_OP_25_64_5665/U131  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_18 ), .Z(
        \DP_OP_25_64_5665/n318 ) );
  XOR \DP_OP_25_64_5665/U109  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_19 ), .Z(
        \DP_OP_25_64_5665/n317 ) );
  XOR \DP_OP_25_64_5665/U108  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_20 ), .Z(
        \DP_OP_25_64_5665/n316 ) );
  XOR \DP_OP_25_64_5665/U107  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_21 ), .Z(
        \DP_OP_25_64_5665/n315 ) );
  XOR \DP_OP_25_64_5665/U106  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_22 ), .Z(
        \DP_OP_25_64_5665/n314 ) );
  XOR \DP_OP_25_64_5665/U105  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_23 ), .Z(
        \DP_OP_25_64_5665/n313 ) );
  XOR \DP_OP_25_64_5665/U104  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_24 ), .Z(
        \DP_OP_25_64_5665/n312 ) );
  XOR \DP_OP_25_64_5665/U103  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_25 ), .Z(
        \DP_OP_25_64_5665/n311 ) );
  XOR \DP_OP_25_64_5665/U102  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_26 ), .Z(
        \DP_OP_25_64_5665/n310 ) );
  XOR \DP_OP_25_64_5665/U101  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_27 ), .Z(
        \DP_OP_25_64_5665/n309 ) );
  XOR \DP_OP_25_64_5665/U100  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_28 ), .Z(
        \DP_OP_25_64_5665/n308 ) );
  XOR \DP_OP_25_64_5665/U99  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_29 ), .Z(
        \DP_OP_25_64_5665/n307 ) );
  XOR \DP_OP_25_64_5665/U98  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_30 ), .Z(
        \DP_OP_25_64_5665/n306 ) );
  XOR \DP_OP_25_64_5665/U97  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_31 ), .Z(
        \DP_OP_25_64_5665/n305 ) );
  XOR \DP_OP_25_64_5665/U94  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_5665/n269 ) );
  XOR \DP_OP_25_64_5665/U93  ( .A(\DP_OP_25_64_5665/n269 ), .B(
        \DP_OP_25_64_5665/n336 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_5665/U92  ( .A(\DP_OP_25_64_5665/n335 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_5665/n268 ) );
  XOR \DP_OP_25_64_5665/U91  ( .A(\DP_OP_25_64_5665/n300 ), .B(
        \DP_OP_25_64_5665/n268 ), .Z(\C3/DATA5_1 ) );
  XOR \DP_OP_25_64_5665/U90  ( .A(\DP_OP_25_64_5665/n334 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_5665/n267 ) );
  XOR \DP_OP_25_64_5665/U88  ( .A(\DP_OP_25_64_5665/n333 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_5665/n266 ) );
  XOR \DP_OP_25_64_5665/U87  ( .A(\DP_OP_25_64_5665/n298 ), .B(
        \DP_OP_25_64_5665/n266 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_5665/U86  ( .A(\DP_OP_25_64_5665/n332 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_5665/n265 ) );
  XOR \DP_OP_25_64_5665/U85  ( .A(\DP_OP_25_64_5665/n297 ), .B(
        \DP_OP_25_64_5665/n265 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_5665/U84  ( .A(\DP_OP_25_64_5665/n331 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_5665/n264 ) );
  XOR \DP_OP_25_64_5665/U83  ( .A(\DP_OP_25_64_5665/n296 ), .B(
        \DP_OP_25_64_5665/n264 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_5665/U82  ( .A(\DP_OP_25_64_5665/n330 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_5665/n263 ) );
  XOR \DP_OP_25_64_5665/U81  ( .A(\DP_OP_25_64_5665/n295 ), .B(
        \DP_OP_25_64_5665/n263 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_5665/U80  ( .A(\DP_OP_25_64_5665/n329 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_5665/n262 ) );
  XOR \DP_OP_25_64_5665/U79  ( .A(\DP_OP_25_64_5665/n294 ), .B(
        \DP_OP_25_64_5665/n262 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_5665/U78  ( .A(\DP_OP_25_64_5665/n328 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_5665/n261 ) );
  XOR \DP_OP_25_64_5665/U77  ( .A(\DP_OP_25_64_5665/n293 ), .B(
        \DP_OP_25_64_5665/n261 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_5665/U76  ( .A(\DP_OP_25_64_5665/n327 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_5665/n260 ) );
  XOR \DP_OP_25_64_5665/U75  ( .A(\DP_OP_25_64_5665/n292 ), .B(
        \DP_OP_25_64_5665/n260 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_5665/U74  ( .A(\DP_OP_25_64_5665/n326 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_5665/n259 ) );
  XOR \DP_OP_25_64_5665/U73  ( .A(\DP_OP_25_64_5665/n291 ), .B(
        \DP_OP_25_64_5665/n259 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_5665/U72  ( .A(\DP_OP_25_64_5665/n325 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_5665/n258 ) );
  XOR \DP_OP_25_64_5665/U71  ( .A(\DP_OP_25_64_5665/n290 ), .B(
        \DP_OP_25_64_5665/n258 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_5665/U70  ( .A(\DP_OP_25_64_5665/n324 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_5665/n257 ) );
  XOR \DP_OP_25_64_5665/U69  ( .A(\DP_OP_25_64_5665/n289 ), .B(
        \DP_OP_25_64_5665/n257 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_5665/U68  ( .A(\DP_OP_25_64_5665/n323 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_5665/n256 ) );
  XOR \DP_OP_25_64_5665/U67  ( .A(\DP_OP_25_64_5665/n288 ), .B(
        \DP_OP_25_64_5665/n256 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_5665/U66  ( .A(\DP_OP_25_64_5665/n322 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_5665/n255 ) );
  XOR \DP_OP_25_64_5665/U65  ( .A(\DP_OP_25_64_5665/n287 ), .B(
        \DP_OP_25_64_5665/n255 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_5665/U64  ( .A(\DP_OP_25_64_5665/n321 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_5665/n254 ) );
  XOR \DP_OP_25_64_5665/U63  ( .A(\DP_OP_25_64_5665/n286 ), .B(
        \DP_OP_25_64_5665/n254 ), .Z(\C3/DATA5_15 ) );
  XOR \DP_OP_25_64_5665/U62  ( .A(\DP_OP_25_64_5665/n320 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_5665/n253 ) );
  XOR \DP_OP_25_64_5665/U61  ( .A(\DP_OP_25_64_5665/n285 ), .B(
        \DP_OP_25_64_5665/n253 ), .Z(\C3/DATA5_16 ) );
  XOR \DP_OP_25_64_5665/U60  ( .A(\DP_OP_25_64_5665/n319 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_5665/n252 ) );
  XOR \DP_OP_25_64_5665/U59  ( .A(\DP_OP_25_64_5665/n284 ), .B(
        \DP_OP_25_64_5665/n252 ), .Z(\C3/DATA5_17 ) );
  XOR \DP_OP_25_64_5665/U58  ( .A(\DP_OP_25_64_5665/n318 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_5665/n251 ) );
  XOR \DP_OP_25_64_5665/U57  ( .A(\DP_OP_25_64_5665/n283 ), .B(
        \DP_OP_25_64_5665/n251 ), .Z(\C3/DATA5_18 ) );
  XOR \DP_OP_25_64_5665/U56  ( .A(\DP_OP_25_64_5665/n317 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_5665/n250 ) );
  XOR \DP_OP_25_64_5665/U55  ( .A(\DP_OP_25_64_5665/n282 ), .B(
        \DP_OP_25_64_5665/n250 ), .Z(\C3/DATA5_19 ) );
  XOR \DP_OP_25_64_5665/U54  ( .A(\DP_OP_25_64_5665/n316 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_5665/n249 ) );
  XOR \DP_OP_25_64_5665/U53  ( .A(\DP_OP_25_64_5665/n281 ), .B(
        \DP_OP_25_64_5665/n249 ), .Z(\C3/DATA5_20 ) );
  XOR \DP_OP_25_64_5665/U52  ( .A(\DP_OP_25_64_5665/n315 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_5665/n248 ) );
  XOR \DP_OP_25_64_5665/U51  ( .A(\DP_OP_25_64_5665/n280 ), .B(
        \DP_OP_25_64_5665/n248 ), .Z(\C3/DATA5_21 ) );
  XOR \DP_OP_25_64_5665/U50  ( .A(\DP_OP_25_64_5665/n314 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_5665/n247 ) );
  XOR \DP_OP_25_64_5665/U49  ( .A(\DP_OP_25_64_5665/n279 ), .B(
        \DP_OP_25_64_5665/n247 ), .Z(\C3/DATA5_22 ) );
  XOR \DP_OP_25_64_5665/U48  ( .A(\DP_OP_25_64_5665/n313 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_5665/n246 ) );
  XOR \DP_OP_25_64_5665/U47  ( .A(\DP_OP_25_64_5665/n278 ), .B(
        \DP_OP_25_64_5665/n246 ), .Z(\C3/DATA5_23 ) );
  XOR \DP_OP_25_64_5665/U46  ( .A(\DP_OP_25_64_5665/n312 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_5665/n245 ) );
  XOR \DP_OP_25_64_5665/U45  ( .A(\DP_OP_25_64_5665/n277 ), .B(
        \DP_OP_25_64_5665/n245 ), .Z(\C3/DATA5_24 ) );
  XOR \DP_OP_25_64_5665/U44  ( .A(\DP_OP_25_64_5665/n311 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_5665/n244 ) );
  XOR \DP_OP_25_64_5665/U43  ( .A(\DP_OP_25_64_5665/n276 ), .B(
        \DP_OP_25_64_5665/n244 ), .Z(\C3/DATA5_25 ) );
  XOR \DP_OP_25_64_5665/U42  ( .A(\DP_OP_25_64_5665/n310 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_5665/n243 ) );
  XOR \DP_OP_25_64_5665/U41  ( .A(\DP_OP_25_64_5665/n275 ), .B(
        \DP_OP_25_64_5665/n243 ), .Z(\C3/DATA5_26 ) );
  XOR \DP_OP_25_64_5665/U40  ( .A(\DP_OP_25_64_5665/n309 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_5665/n242 ) );
  XOR \DP_OP_25_64_5665/U30  ( .A(\DP_OP_25_64_5665/n274 ), .B(
        \DP_OP_25_64_5665/n242 ), .Z(\C3/DATA5_27 ) );
  XOR \DP_OP_25_64_5665/U20  ( .A(\DP_OP_25_64_5665/n308 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_5665/n241 ) );
  XOR \DP_OP_25_64_5665/U10  ( .A(\DP_OP_25_64_5665/n273 ), .B(
        \DP_OP_25_64_5665/n241 ), .Z(\C3/DATA5_28 ) );
  XOR \DP_OP_25_64_5665/U9  ( .A(\DP_OP_25_64_5665/n307 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_5665/n240 ) );
  XOR \DP_OP_25_64_5665/U8  ( .A(\DP_OP_25_64_5665/n272 ), .B(
        \DP_OP_25_64_5665/n240 ), .Z(\C3/DATA5_29 ) );
  XOR \DP_OP_25_64_5665/U7  ( .A(\DP_OP_25_64_5665/n306 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_5665/n239 ) );
  XOR \DP_OP_25_64_5665/U6  ( .A(\DP_OP_25_64_5665/n271 ), .B(
        \DP_OP_25_64_5665/n239 ), .Z(\C3/DATA5_30 ) );
  XOR \DP_OP_25_64_5665/U5  ( .A(\DP_OP_25_64_5665/n305 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_5665/n238 ) );
  XOR \DP_OP_25_64_5665/U4  ( .A(\DP_OP_25_64_5665/n270 ), .B(
        \DP_OP_25_64_5665/n238 ), .Z(\C3/DATA5_31 ) );
  NAND \DP_OP_25_64_5665/U130  ( .A(\DP_OP_25_64_5665/n306 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_5665/n5 ) );
  NAND \DP_OP_25_64_5665/U230  ( .A(\DP_OP_25_64_5665/n271 ), .B(
        \DP_OP_25_64_5665/n239 ), .Z(\DP_OP_25_64_5665/n8 ) );
  NAND \DP_OP_25_64_5665/U330  ( .A(\DP_OP_25_64_5665/n5 ), .B(
        \DP_OP_25_64_5665/n8 ), .Z(\DP_OP_25_64_5665/n270 ) );
  NAND \DP_OP_25_64_5665/U129  ( .A(\DP_OP_25_64_5665/n307 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_5665/n14 ) );
  NAND \DP_OP_25_64_5665/U229  ( .A(\DP_OP_25_64_5665/n272 ), .B(
        \DP_OP_25_64_5665/n240 ), .Z(\DP_OP_25_64_5665/n15 ) );
  NAND \DP_OP_25_64_5665/U329  ( .A(\DP_OP_25_64_5665/n14 ), .B(
        \DP_OP_25_64_5665/n15 ), .Z(\DP_OP_25_64_5665/n271 ) );
  NAND \DP_OP_25_64_5665/U128  ( .A(\DP_OP_25_64_5665/n308 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_5665/n21 ) );
  NAND \DP_OP_25_64_5665/U228  ( .A(\DP_OP_25_64_5665/n273 ), .B(
        \DP_OP_25_64_5665/n241 ), .Z(\DP_OP_25_64_5665/n22 ) );
  NAND \DP_OP_25_64_5665/U328  ( .A(\DP_OP_25_64_5665/n21 ), .B(
        \DP_OP_25_64_5665/n22 ), .Z(\DP_OP_25_64_5665/n272 ) );
  NAND \DP_OP_25_64_5665/U127  ( .A(\DP_OP_25_64_5665/n309 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_5665/n28 ) );
  NAND \DP_OP_25_64_5665/U227  ( .A(\DP_OP_25_64_5665/n274 ), .B(
        \DP_OP_25_64_5665/n242 ), .Z(\DP_OP_25_64_5665/n29 ) );
  NAND \DP_OP_25_64_5665/U327  ( .A(\DP_OP_25_64_5665/n28 ), .B(
        \DP_OP_25_64_5665/n29 ), .Z(\DP_OP_25_64_5665/n273 ) );
  NAND \DP_OP_25_64_5665/U126  ( .A(\DP_OP_25_64_5665/n310 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_5665/n35 ) );
  NAND \DP_OP_25_64_5665/U226  ( .A(\DP_OP_25_64_5665/n275 ), .B(
        \DP_OP_25_64_5665/n243 ), .Z(\DP_OP_25_64_5665/n36 ) );
  NAND \DP_OP_25_64_5665/U326  ( .A(\DP_OP_25_64_5665/n35 ), .B(
        \DP_OP_25_64_5665/n36 ), .Z(\DP_OP_25_64_5665/n274 ) );
  NAND \DP_OP_25_64_5665/U125  ( .A(\DP_OP_25_64_5665/n311 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_5665/n42 ) );
  NAND \DP_OP_25_64_5665/U225  ( .A(\DP_OP_25_64_5665/n276 ), .B(
        \DP_OP_25_64_5665/n244 ), .Z(\DP_OP_25_64_5665/n43 ) );
  NAND \DP_OP_25_64_5665/U325  ( .A(\DP_OP_25_64_5665/n42 ), .B(
        \DP_OP_25_64_5665/n43 ), .Z(\DP_OP_25_64_5665/n275 ) );
  NAND \DP_OP_25_64_5665/U124  ( .A(\DP_OP_25_64_5665/n312 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_5665/n49 ) );
  NAND \DP_OP_25_64_5665/U224  ( .A(\DP_OP_25_64_5665/n277 ), .B(
        \DP_OP_25_64_5665/n245 ), .Z(\DP_OP_25_64_5665/n50 ) );
  NAND \DP_OP_25_64_5665/U324  ( .A(\DP_OP_25_64_5665/n49 ), .B(
        \DP_OP_25_64_5665/n50 ), .Z(\DP_OP_25_64_5665/n276 ) );
  NAND \DP_OP_25_64_5665/U123  ( .A(\DP_OP_25_64_5665/n313 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_5665/n56 ) );
  NAND \DP_OP_25_64_5665/U223  ( .A(\DP_OP_25_64_5665/n278 ), .B(
        \DP_OP_25_64_5665/n246 ), .Z(\DP_OP_25_64_5665/n57 ) );
  NAND \DP_OP_25_64_5665/U323  ( .A(\DP_OP_25_64_5665/n56 ), .B(
        \DP_OP_25_64_5665/n57 ), .Z(\DP_OP_25_64_5665/n277 ) );
  NAND \DP_OP_25_64_5665/U122  ( .A(\DP_OP_25_64_5665/n314 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_5665/n81 ) );
  NAND \DP_OP_25_64_5665/U222  ( .A(\DP_OP_25_64_5665/n279 ), .B(
        \DP_OP_25_64_5665/n247 ), .Z(\DP_OP_25_64_5665/n82 ) );
  NAND \DP_OP_25_64_5665/U322  ( .A(\DP_OP_25_64_5665/n81 ), .B(
        \DP_OP_25_64_5665/n82 ), .Z(\DP_OP_25_64_5665/n278 ) );
  NAND \DP_OP_25_64_5665/U121  ( .A(\DP_OP_25_64_5665/n315 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_5665/n88 ) );
  NAND \DP_OP_25_64_5665/U221  ( .A(\DP_OP_25_64_5665/n280 ), .B(
        \DP_OP_25_64_5665/n248 ), .Z(\DP_OP_25_64_5665/n89 ) );
  NAND \DP_OP_25_64_5665/U321  ( .A(\DP_OP_25_64_5665/n88 ), .B(
        \DP_OP_25_64_5665/n89 ), .Z(\DP_OP_25_64_5665/n279 ) );
  NAND \DP_OP_25_64_5665/U120  ( .A(\DP_OP_25_64_5665/n316 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_5665/n95 ) );
  NAND \DP_OP_25_64_5665/U220  ( .A(\DP_OP_25_64_5665/n281 ), .B(
        \DP_OP_25_64_5665/n249 ), .Z(\DP_OP_25_64_5665/n96 ) );
  NAND \DP_OP_25_64_5665/U320  ( .A(\DP_OP_25_64_5665/n95 ), .B(
        \DP_OP_25_64_5665/n96 ), .Z(\DP_OP_25_64_5665/n280 ) );
  NAND \DP_OP_25_64_5665/U119  ( .A(\DP_OP_25_64_5665/n317 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_5665/n102 ) );
  NAND \DP_OP_25_64_5665/U219  ( .A(\DP_OP_25_64_5665/n282 ), .B(
        \DP_OP_25_64_5665/n250 ), .Z(\DP_OP_25_64_5665/n103 ) );
  NAND \DP_OP_25_64_5665/U319  ( .A(\DP_OP_25_64_5665/n102 ), .B(
        \DP_OP_25_64_5665/n103 ), .Z(\DP_OP_25_64_5665/n281 ) );
  NAND \DP_OP_25_64_5665/U118  ( .A(\DP_OP_25_64_5665/n318 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_5665/n109 ) );
  NAND \DP_OP_25_64_5665/U218  ( .A(\DP_OP_25_64_5665/n283 ), .B(
        \DP_OP_25_64_5665/n251 ), .Z(\DP_OP_25_64_5665/n110 ) );
  NAND \DP_OP_25_64_5665/U318  ( .A(\DP_OP_25_64_5665/n109 ), .B(
        \DP_OP_25_64_5665/n110 ), .Z(\DP_OP_25_64_5665/n282 ) );
  NAND \DP_OP_25_64_5665/U117  ( .A(\DP_OP_25_64_5665/n319 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_5665/n116 ) );
  NAND \DP_OP_25_64_5665/U217  ( .A(\DP_OP_25_64_5665/n284 ), .B(
        \DP_OP_25_64_5665/n252 ), .Z(\DP_OP_25_64_5665/n117 ) );
  NAND \DP_OP_25_64_5665/U317  ( .A(\DP_OP_25_64_5665/n116 ), .B(
        \DP_OP_25_64_5665/n117 ), .Z(\DP_OP_25_64_5665/n283 ) );
  NAND \DP_OP_25_64_5665/U116  ( .A(\DP_OP_25_64_5665/n320 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_5665/n123 ) );
  NAND \DP_OP_25_64_5665/U216  ( .A(\DP_OP_25_64_5665/n285 ), .B(
        \DP_OP_25_64_5665/n253 ), .Z(\DP_OP_25_64_5665/n124 ) );
  NAND \DP_OP_25_64_5665/U316  ( .A(\DP_OP_25_64_5665/n123 ), .B(
        \DP_OP_25_64_5665/n124 ), .Z(\DP_OP_25_64_5665/n284 ) );
  NAND \DP_OP_25_64_5665/U115  ( .A(\DP_OP_25_64_5665/n321 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_5665/n130 ) );
  NAND \DP_OP_25_64_5665/U215  ( .A(\DP_OP_25_64_5665/n286 ), .B(
        \DP_OP_25_64_5665/n254 ), .Z(\DP_OP_25_64_5665/n131 ) );
  NAND \DP_OP_25_64_5665/U315  ( .A(\DP_OP_25_64_5665/n130 ), .B(
        \DP_OP_25_64_5665/n131 ), .Z(\DP_OP_25_64_5665/n285 ) );
  NAND \DP_OP_25_64_5665/U114  ( .A(\DP_OP_25_64_5665/n322 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_5665/n137 ) );
  NAND \DP_OP_25_64_5665/U214  ( .A(\DP_OP_25_64_5665/n287 ), .B(
        \DP_OP_25_64_5665/n255 ), .Z(\DP_OP_25_64_5665/n138 ) );
  NAND \DP_OP_25_64_5665/U314  ( .A(\DP_OP_25_64_5665/n137 ), .B(
        \DP_OP_25_64_5665/n138 ), .Z(\DP_OP_25_64_5665/n286 ) );
  NAND \DP_OP_25_64_5665/U113  ( .A(\DP_OP_25_64_5665/n323 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_5665/n144 ) );
  NAND \DP_OP_25_64_5665/U213  ( .A(\DP_OP_25_64_5665/n288 ), .B(
        \DP_OP_25_64_5665/n256 ), .Z(\DP_OP_25_64_5665/n145 ) );
  NAND \DP_OP_25_64_5665/U313  ( .A(\DP_OP_25_64_5665/n144 ), .B(
        \DP_OP_25_64_5665/n145 ), .Z(\DP_OP_25_64_5665/n287 ) );
  NAND \DP_OP_25_64_5665/U112  ( .A(\DP_OP_25_64_5665/n324 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_5665/n151 ) );
  NAND \DP_OP_25_64_5665/U212  ( .A(\DP_OP_25_64_5665/n289 ), .B(
        \DP_OP_25_64_5665/n257 ), .Z(\DP_OP_25_64_5665/n152 ) );
  NAND \DP_OP_25_64_5665/U312  ( .A(\DP_OP_25_64_5665/n151 ), .B(
        \DP_OP_25_64_5665/n152 ), .Z(\DP_OP_25_64_5665/n288 ) );
  NAND \DP_OP_25_64_5665/U111  ( .A(\DP_OP_25_64_5665/n325 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_5665/n158 ) );
  NAND \DP_OP_25_64_5665/U211  ( .A(\DP_OP_25_64_5665/n290 ), .B(
        \DP_OP_25_64_5665/n258 ), .Z(\DP_OP_25_64_5665/n159 ) );
  NAND \DP_OP_25_64_5665/U311  ( .A(\DP_OP_25_64_5665/n158 ), .B(
        \DP_OP_25_64_5665/n159 ), .Z(\DP_OP_25_64_5665/n289 ) );
  NAND \DP_OP_25_64_5665/U110  ( .A(\DP_OP_25_64_5665/n326 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_5665/n165 ) );
  NAND \DP_OP_25_64_5665/U210  ( .A(\DP_OP_25_64_5665/n291 ), .B(
        \DP_OP_25_64_5665/n259 ), .Z(\DP_OP_25_64_5665/n166 ) );
  NAND \DP_OP_25_64_5665/U310  ( .A(\DP_OP_25_64_5665/n165 ), .B(
        \DP_OP_25_64_5665/n166 ), .Z(\DP_OP_25_64_5665/n290 ) );
  NAND \DP_OP_25_64_5665/U19  ( .A(\DP_OP_25_64_5665/n327 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_5665/n172 ) );
  NAND \DP_OP_25_64_5665/U29  ( .A(\DP_OP_25_64_5665/n292 ), .B(
        \DP_OP_25_64_5665/n260 ), .Z(\DP_OP_25_64_5665/n173 ) );
  NAND \DP_OP_25_64_5665/U39  ( .A(\DP_OP_25_64_5665/n172 ), .B(
        \DP_OP_25_64_5665/n173 ), .Z(\DP_OP_25_64_5665/n291 ) );
  NAND \DP_OP_25_64_5665/U18  ( .A(\DP_OP_25_64_5665/n328 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_5665/n179 ) );
  NAND \DP_OP_25_64_5665/U28  ( .A(\DP_OP_25_64_5665/n293 ), .B(
        \DP_OP_25_64_5665/n261 ), .Z(\DP_OP_25_64_5665/n180 ) );
  NAND \DP_OP_25_64_5665/U38  ( .A(\DP_OP_25_64_5665/n179 ), .B(
        \DP_OP_25_64_5665/n180 ), .Z(\DP_OP_25_64_5665/n292 ) );
  NAND \DP_OP_25_64_5665/U17  ( .A(\DP_OP_25_64_5665/n329 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_5665/n186 ) );
  NAND \DP_OP_25_64_5665/U27  ( .A(\DP_OP_25_64_5665/n294 ), .B(
        \DP_OP_25_64_5665/n262 ), .Z(\DP_OP_25_64_5665/n187 ) );
  NAND \DP_OP_25_64_5665/U37  ( .A(\DP_OP_25_64_5665/n186 ), .B(
        \DP_OP_25_64_5665/n187 ), .Z(\DP_OP_25_64_5665/n293 ) );
  NAND \DP_OP_25_64_5665/U16  ( .A(\DP_OP_25_64_5665/n330 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_5665/n193 ) );
  NAND \DP_OP_25_64_5665/U26  ( .A(\DP_OP_25_64_5665/n295 ), .B(
        \DP_OP_25_64_5665/n263 ), .Z(\DP_OP_25_64_5665/n194 ) );
  NAND \DP_OP_25_64_5665/U36  ( .A(\DP_OP_25_64_5665/n193 ), .B(
        \DP_OP_25_64_5665/n194 ), .Z(\DP_OP_25_64_5665/n294 ) );
  NAND \DP_OP_25_64_5665/U15  ( .A(\DP_OP_25_64_5665/n331 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_5665/n200 ) );
  NAND \DP_OP_25_64_5665/U25  ( .A(\DP_OP_25_64_5665/n296 ), .B(
        \DP_OP_25_64_5665/n264 ), .Z(\DP_OP_25_64_5665/n201 ) );
  NAND \DP_OP_25_64_5665/U35  ( .A(\DP_OP_25_64_5665/n200 ), .B(
        \DP_OP_25_64_5665/n201 ), .Z(\DP_OP_25_64_5665/n295 ) );
  NAND \DP_OP_25_64_5665/U14  ( .A(\DP_OP_25_64_5665/n332 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_5665/n207 ) );
  NAND \DP_OP_25_64_5665/U24  ( .A(\DP_OP_25_64_5665/n297 ), .B(
        \DP_OP_25_64_5665/n265 ), .Z(\DP_OP_25_64_5665/n208 ) );
  NAND \DP_OP_25_64_5665/U34  ( .A(\DP_OP_25_64_5665/n207 ), .B(
        \DP_OP_25_64_5665/n208 ), .Z(\DP_OP_25_64_5665/n296 ) );
  NAND \DP_OP_25_64_5665/U13  ( .A(\DP_OP_25_64_5665/n333 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_5665/n214 ) );
  NAND \DP_OP_25_64_5665/U23  ( .A(\DP_OP_25_64_5665/n298 ), .B(
        \DP_OP_25_64_5665/n266 ), .Z(\DP_OP_25_64_5665/n215 ) );
  NAND \DP_OP_25_64_5665/U33  ( .A(\DP_OP_25_64_5665/n214 ), .B(
        \DP_OP_25_64_5665/n215 ), .Z(\DP_OP_25_64_5665/n297 ) );
  NAND \DP_OP_25_64_5665/U12  ( .A(\DP_OP_25_64_5665/n334 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_5665/n221 ) );
  NAND \DP_OP_25_64_5665/U22  ( .A(\DP_OP_25_64_5665/n299 ), .B(
        \DP_OP_25_64_5665/n267 ), .Z(\DP_OP_25_64_5665/n222 ) );
  NAND \DP_OP_25_64_5665/U32  ( .A(\DP_OP_25_64_5665/n221 ), .B(
        \DP_OP_25_64_5665/n222 ), .Z(\DP_OP_25_64_5665/n298 ) );
  NAND \DP_OP_25_64_5665/U11  ( .A(\DP_OP_25_64_5665/n335 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_5665/n228 ) );
  NAND \DP_OP_25_64_5665/U21  ( .A(\DP_OP_25_64_5665/n300 ), .B(
        \DP_OP_25_64_5665/n268 ), .Z(\DP_OP_25_64_5665/n229 ) );
  NAND \DP_OP_25_64_5665/U31  ( .A(\DP_OP_25_64_5665/n228 ), .B(
        \DP_OP_25_64_5665/n229 ), .Z(\DP_OP_25_64_5665/n299 ) );
  NAND \DP_OP_25_64_5665/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_5665/n235 ) );
  NAND \DP_OP_25_64_5665/U2  ( .A(\DP_OP_25_64_5665/n269 ), .B(
        \DP_OP_25_64_5665/n336 ), .Z(\DP_OP_25_64_5665/n236 ) );
  NAND \DP_OP_25_64_5665/U3  ( .A(\DP_OP_25_64_5665/n235 ), .B(
        \DP_OP_25_64_5665/n236 ), .Z(\DP_OP_25_64_5665/n300 ) );
  XOR U1492 ( .A(n2180), .B(n2181), .Z(n2183) );
  XOR U1493 ( .A(n2550), .B(n2551), .Z(n2887) );
  XOR U1494 ( .A(n2537), .B(n2538), .Z(n2540) );
  XOR U1495 ( .A(n2899), .B(n2900), .Z(n3025) );
  XOR U1496 ( .A(n3710), .B(n3711), .Z(n3756) );
  XOR U1497 ( .A(n3662), .B(n3663), .Z(n3759) );
  XOR U1498 ( .A(n2945), .B(n2946), .Z(n2956) );
  XOR U1499 ( .A(n3888), .B(n3889), .Z(n4062) );
  XOR U1500 ( .A(n3878), .B(n3879), .Z(n4049) );
  XOR U1501 ( .A(n4045), .B(n4046), .Z(n4209) );
  XOR U1502 ( .A(n4019), .B(n4020), .Z(n4186) );
  XOR U1503 ( .A(n3949), .B(n3950), .Z(n3952) );
  XOR U1504 ( .A(n4069), .B(n4070), .Z(n4233) );
  XOR U1505 ( .A(n2098), .B(n2099), .Z(n2154) );
  XOR U1506 ( .A(n2172), .B(n2173), .Z(n2432) );
  XOR U1507 ( .A(n2459), .B(n2460), .Z(n2559) );
  XOR U1508 ( .A(n2447), .B(n2448), .Z(n2551) );
  XOR U1509 ( .A(n2428), .B(n2429), .Z(n2511) );
  XOR U1510 ( .A(n2549), .B(n5315), .Z(n2888) );
  XOR U1511 ( .A(n2539), .B(n2540), .Z(n2876) );
  XOR U1512 ( .A(n2529), .B(n2530), .Z(n2863) );
  XOR U1513 ( .A(n2857), .B(n2858), .Z(n2964) );
  XOR U1514 ( .A(n3034), .B(n3035), .Z(n3301) );
  XOR U1515 ( .A(n2895), .B(n2896), .Z(n3017) );
  XOR U1516 ( .A(n3012), .B(n3013), .Z(n3221) );
  XOR U1517 ( .A(n2981), .B(n2982), .Z(n3243) );
  XOR U1518 ( .A(n3046), .B(n3047), .Z(n3313) );
  XOR U1519 ( .A(n3256), .B(n3257), .Z(n3653) );
  XOR U1520 ( .A(n3239), .B(n3240), .Z(n3612) );
  XOR U1521 ( .A(n3326), .B(n3327), .Z(n3724) );
  XOR U1522 ( .A(n3720), .B(n3721), .Z(n3871) );
  XOR U1523 ( .A(n3274), .B(n3275), .Z(n3667) );
  XOR U1524 ( .A(n3660), .B(n3661), .Z(n3760) );
  XOR U1525 ( .A(n3650), .B(n3651), .Z(n3805) );
  XOR U1526 ( .A(n3630), .B(n3631), .Z(n3780) );
  XOR U1527 ( .A(n3794), .B(n3795), .Z(n3964) );
  XOR U1528 ( .A(n3774), .B(n3775), .Z(n3925) );
  XOR U1529 ( .A(n4055), .B(n4056), .Z(n4222) );
  XOR U1530 ( .A(n4043), .B(n4044), .Z(n4210) );
  XOR U1531 ( .A(n4033), .B(n4034), .Z(n4197) );
  XOR U1532 ( .A(n4021), .B(n4022), .Z(n4185) );
  XOR U1533 ( .A(n4007), .B(n4008), .Z(n4174) );
  XOR U1534 ( .A(n3997), .B(n3998), .Z(n4161) );
  XOR U1535 ( .A(n3985), .B(n3986), .Z(n4081) );
  XOR U1536 ( .A(n3961), .B(n3962), .Z(n4130) );
  XOR U1537 ( .A(n3951), .B(n3952), .Z(n4118) );
  XOR U1538 ( .A(n3941), .B(n3942), .Z(n4105) );
  XOR U1539 ( .A(n3196), .B(n3195), .Z(n3202) );
  XOR U1540 ( .A(n4093), .B(n4094), .Z(n4096) );
  XOR U1541 ( .A(n4067), .B(n4068), .Z(n4234) );
  XOR U1542 ( .A(n4141), .B(n4142), .Z(n4324) );
  XOR U1543 ( .A(n2090), .B(n2091), .Z(n2093) );
  XOR U1544 ( .A(n1908), .B(n1909), .Z(n2099) );
  XOR U1545 ( .A(n2182), .B(n2183), .Z(n2446) );
  XOR U1546 ( .A(n2420), .B(n2421), .Z(n2423) );
  XOR U1547 ( .A(n2439), .B(n2440), .Z(n2442) );
  XOR U1548 ( .A(n2192), .B(n2193), .Z(n2458) );
  XOR U1549 ( .A(n2560), .B(n2561), .Z(n2841) );
  XOR U1550 ( .A(n2570), .B(n2571), .Z(n2910) );
  XOR U1551 ( .A(n1934), .B(n1935), .Z(n2127) );
  XOR U1552 ( .A(n2875), .B(n2876), .Z(n2878) );
  XOR U1553 ( .A(n2889), .B(n2890), .Z(n3011) );
  XOR U1554 ( .A(n2869), .B(n2870), .Z(n2872) );
  XOR U1555 ( .A(n3024), .B(n3025), .Z(n3288) );
  XOR U1556 ( .A(n2989), .B(n2990), .Z(n2992) );
  XOR U1557 ( .A(n3314), .B(n3315), .Z(n3709) );
  XOR U1558 ( .A(n3302), .B(n3303), .Z(n3697) );
  XOR U1559 ( .A(n3018), .B(n3019), .Z(n3283) );
  XOR U1560 ( .A(n3268), .B(n3269), .Z(n3661) );
  XOR U1561 ( .A(n3249), .B(n3250), .Z(n3252) );
  XOR U1562 ( .A(n3237), .B(n3238), .Z(n3613) );
  XNOR U1563 ( .A(n3320), .B(n3321), .Z(n3715) );
  XOR U1564 ( .A(n3698), .B(n3699), .Z(n3848) );
  XOR U1565 ( .A(n3684), .B(n3685), .Z(n3837) );
  XOR U1566 ( .A(n3284), .B(n3285), .Z(n3678) );
  XOR U1567 ( .A(n3674), .B(n3675), .Z(n3757) );
  XOR U1568 ( .A(n3640), .B(n3641), .Z(n3793) );
  XOR U1569 ( .A(n3622), .B(n3623), .Z(n3625) );
  XOR U1570 ( .A(n2697), .B(n2696), .Z(n2699) );
  XOR U1571 ( .A(n3733), .B(n3734), .Z(n3883) );
  XNOR U1572 ( .A(n2754), .B(n2753), .Z(n2798) );
  XOR U1573 ( .A(n3668), .B(n3669), .Z(n3821) );
  XOR U1574 ( .A(n3890), .B(n3891), .Z(n4061) );
  XOR U1575 ( .A(n3876), .B(n3877), .Z(n4050) );
  XOR U1576 ( .A(n3866), .B(n3867), .Z(n4037) );
  XOR U1577 ( .A(n3856), .B(n3857), .Z(n4025) );
  XOR U1578 ( .A(n3832), .B(n3833), .Z(n4002) );
  XOR U1579 ( .A(n3822), .B(n3823), .Z(n3989) );
  XOR U1580 ( .A(n3812), .B(n3813), .Z(n3978) );
  XOR U1581 ( .A(n3971), .B(n3972), .Z(n4084) );
  XOR U1582 ( .A(n3788), .B(n3789), .Z(n3955) );
  XOR U1583 ( .A(n3096), .B(n3095), .Z(n3208) );
  XOR U1584 ( .A(n3945), .B(n3946), .Z(n4112) );
  XOR U1585 ( .A(n3350), .B(n3351), .Z(n3609) );
  XOR U1586 ( .A(n4235), .B(n4236), .Z(n4246) );
  XOR U1587 ( .A(n4223), .B(n4224), .Z(n4248) );
  XOR U1588 ( .A(n4211), .B(n4212), .Z(n4250) );
  XOR U1589 ( .A(n4199), .B(n4200), .Z(n4252) );
  XOR U1590 ( .A(n4187), .B(n4188), .Z(n4254) );
  XOR U1591 ( .A(n4175), .B(n4176), .Z(n4256) );
  XOR U1592 ( .A(n4163), .B(n4164), .Z(n4258) );
  XOR U1593 ( .A(n4151), .B(n4152), .Z(n4260) );
  XOR U1594 ( .A(n4131), .B(n4132), .Z(n4262) );
  XOR U1595 ( .A(n4119), .B(n4120), .Z(n4301) );
  XOR U1596 ( .A(n4107), .B(n4108), .Z(n4264) );
  XOR U1597 ( .A(n4095), .B(n4096), .Z(n4266) );
  XOR U1598 ( .A(n4422), .B(n4421), .Z(n4420) );
  XOR U1599 ( .A(n4323), .B(n4324), .Z(n4326) );
  XOR U1600 ( .A(n1914), .B(n1915), .Z(n2102) );
  XOR U1601 ( .A(n2096), .B(n2097), .Z(n2155) );
  XOR U1602 ( .A(n1856), .B(n1857), .Z(n1912) );
  XOR U1603 ( .A(n2164), .B(n2165), .Z(n2167) );
  XOR U1604 ( .A(n2445), .B(n2446), .Z(n2448) );
  XNOR U1605 ( .A(n1726), .B(n1727), .Z(n1728) );
  XOR U1606 ( .A(n2422), .B(n2423), .Z(n2527) );
  XOR U1607 ( .A(n2558), .B(n2559), .Z(n2842) );
  XOR U1608 ( .A(n2441), .B(n2442), .Z(n2543) );
  XOR U1609 ( .A(n2521), .B(n2522), .Z(n2524) );
  XOR U1610 ( .A(n2469), .B(n2470), .Z(n2573) );
  XOR U1611 ( .A(n2564), .B(n2565), .Z(n2567) );
  XOR U1612 ( .A(n2533), .B(n2534), .Z(n2870) );
  XOR U1613 ( .A(n2851), .B(n2852), .Z(n2854) );
  XOR U1614 ( .A(n2554), .B(n2555), .Z(n2894) );
  XOR U1615 ( .A(n2877), .B(n2878), .Z(n3003) );
  XNOR U1616 ( .A(n2150), .B(n2151), .Z(n2208) );
  XOR U1617 ( .A(n1838), .B(n1839), .Z(n1885) );
  XOR U1618 ( .A(n1955), .B(n1954), .Z(n1957) );
  XOR U1619 ( .A(n3036), .B(n3037), .Z(n3300) );
  XOR U1620 ( .A(n2905), .B(n2906), .Z(n3028) );
  XOR U1621 ( .A(n3022), .B(n3023), .Z(n3289) );
  XOR U1622 ( .A(n2973), .B(n2974), .Z(n2976) );
  XOR U1623 ( .A(n2019), .B(n2018), .Z(n2063) );
  XOR U1624 ( .A(n3040), .B(n3041), .Z(n3043) );
  XOR U1625 ( .A(n2985), .B(n2986), .Z(n3250) );
  XOR U1626 ( .A(n3231), .B(n3232), .Z(n3234) );
  XOR U1627 ( .A(n2074), .B(n2075), .Z(n2145) );
  XOR U1628 ( .A(n2241), .B(n2240), .Z(n2243) );
  XOR U1629 ( .A(n2299), .B(n2298), .Z(n2301) );
  XOR U1630 ( .A(n3278), .B(n3279), .Z(n3675) );
  XOR U1631 ( .A(n3006), .B(n3007), .Z(n3273) );
  XOR U1632 ( .A(n2997), .B(n2998), .Z(n3260) );
  XOR U1633 ( .A(n3245), .B(n3246), .Z(n3638) );
  XOR U1634 ( .A(n3318), .B(n3319), .Z(n3714) );
  XOR U1635 ( .A(n3296), .B(n3297), .Z(n3690) );
  XOR U1636 ( .A(n3282), .B(n3283), .Z(n3679) );
  XOR U1637 ( .A(n3672), .B(n3673), .Z(n3758) );
  XOR U1638 ( .A(n3262), .B(n3263), .Z(n3610) );
  XOR U1639 ( .A(n3652), .B(n3653), .Z(n3804) );
  XOR U1640 ( .A(n2327), .B(n2326), .Z(n2395) );
  XOR U1641 ( .A(n2685), .B(n2684), .Z(n2687) );
  XOR U1642 ( .A(n3634), .B(n3635), .Z(n3787) );
  XOR U1643 ( .A(n3624), .B(n3625), .Z(n3777) );
  XOR U1644 ( .A(n3768), .B(n3769), .Z(n3771) );
  XOR U1645 ( .A(n2798), .B(n2797), .Z(n2800) );
  XOR U1646 ( .A(n3729), .B(n3730), .Z(n3877) );
  XOR U1647 ( .A(n3704), .B(n3705), .Z(n3854) );
  XOR U1648 ( .A(n3850), .B(n3851), .Z(n4020) );
  XOR U1649 ( .A(n3838), .B(n3839), .Z(n4010) );
  XOR U1650 ( .A(n3646), .B(n3647), .Z(n3798) );
  XOR U1651 ( .A(n3782), .B(n3783), .Z(n3950) );
  XNOR U1652 ( .A(n2736), .B(n2735), .Z(n2816) );
  XOR U1653 ( .A(n4031), .B(n4032), .Z(n4198) );
  XOR U1654 ( .A(n3995), .B(n3996), .Z(n4162) );
  XOR U1655 ( .A(n3820), .B(n3821), .Z(n3990) );
  XOR U1656 ( .A(n3983), .B(n3984), .Z(n4082) );
  XOR U1657 ( .A(n3973), .B(n3974), .Z(n4083) );
  XOR U1658 ( .A(n3800), .B(n3801), .Z(n3922) );
  XOR U1659 ( .A(n3963), .B(n3964), .Z(n4129) );
  XOR U1660 ( .A(n3747), .B(n3748), .Z(n3894) );
  XOR U1661 ( .A(n3090), .B(n3089), .Z(n3214) );
  XOR U1662 ( .A(n4001), .B(n4002), .Z(n4004) );
  XOR U1663 ( .A(n3977), .B(n3978), .Z(n3980) );
  XOR U1664 ( .A(n3933), .B(n3934), .Z(n3936) );
  XNOR U1665 ( .A(n3553), .B(n3552), .Z(n3579) );
  XOR U1666 ( .A(n3957), .B(n3958), .Z(n4124) );
  XOR U1667 ( .A(n4111), .B(n4112), .Z(n4114) );
  XOR U1668 ( .A(n4239), .B(n4240), .Z(n4412) );
  XOR U1669 ( .A(n4215), .B(n4216), .Z(n4392) );
  XOR U1670 ( .A(n4191), .B(n4192), .Z(n4372) );
  XOR U1671 ( .A(n4179), .B(n4180), .Z(n4362) );
  XOR U1672 ( .A(n4125), .B(n4126), .Z(n4309) );
  XOR U1673 ( .A(n4416), .B(n4415), .Z(n4480) );
  XOR U1674 ( .A(n4405), .B(n4406), .Z(n4556) );
  XOR U1675 ( .A(n4395), .B(n4396), .Z(n4632) );
  XOR U1676 ( .A(n4385), .B(n4386), .Z(n4708) );
  XOR U1677 ( .A(n4375), .B(n4376), .Z(n4784) );
  XOR U1678 ( .A(n4365), .B(n4366), .Z(n4860) );
  XOR U1679 ( .A(n4355), .B(n4356), .Z(n4936) );
  XOR U1680 ( .A(n4345), .B(n4346), .Z(n5012) );
  XOR U1681 ( .A(n4335), .B(n4336), .Z(n5090) );
  XOR U1682 ( .A(n4325), .B(n4326), .Z(n5166) );
  XOR U1683 ( .A(n4313), .B(n4314), .Z(n5242) );
  XOR U1684 ( .A(n4303), .B(n4304), .Z(n5319) );
  XOR U1685 ( .A(n4291), .B(n4292), .Z(n5397) );
  XOR U1686 ( .A(n4281), .B(n4282), .Z(n5473) );
  XOR U1687 ( .A(n1906), .B(n1907), .Z(n1909) );
  XOR U1688 ( .A(n2092), .B(n2093), .Z(n2170) );
  XOR U1689 ( .A(n2104), .B(n2105), .Z(n2181) );
  XOR U1690 ( .A(n2176), .B(n2177), .Z(n2440) );
  XOR U1691 ( .A(n2166), .B(n2167), .Z(n2429) );
  XOR U1692 ( .A(n1728), .B(n1729), .Z(n1843) );
  XOR U1693 ( .A(n2188), .B(n2189), .Z(n2451) );
  XOR U1694 ( .A(n2426), .B(n2427), .Z(n2512) );
  XOR U1695 ( .A(n1692), .B(n1693), .Z(n1719) );
  XOR U1696 ( .A(n2453), .B(n2454), .Z(n2509) );
  XOR U1697 ( .A(n2198), .B(n2199), .Z(n2464) );
  XOR U1698 ( .A(n2523), .B(n2524), .Z(n2860) );
  XOR U1699 ( .A(n1878), .B(n1879), .Z(n1889) );
  XOR U1700 ( .A(n2911), .B(n2912), .Z(n3035) );
  XOR U1701 ( .A(n2566), .B(n2567), .Z(n2903) );
  XOR U1702 ( .A(n2545), .B(n2546), .Z(n2881) );
  XOR U1703 ( .A(n2853), .B(n2854), .Z(n2979) );
  XOR U1704 ( .A(n2408), .B(n2409), .Z(n2480) );
  XNOR U1705 ( .A(n1951), .B(n1950), .Z(n1944) );
  XOR U1706 ( .A(n3010), .B(n3011), .Z(n3222) );
  XOR U1707 ( .A(n2883), .B(n2884), .Z(n2961) );
  XOR U1708 ( .A(n3001), .B(n3002), .Z(n3267) );
  XOR U1709 ( .A(n2871), .B(n2872), .Z(n2995) );
  XOR U1710 ( .A(n2991), .B(n2992), .Z(n3255) );
  XOR U1711 ( .A(n2031), .B(n2030), .Z(n2047) );
  XOR U1712 ( .A(n3016), .B(n3017), .Z(n3019) );
  XOR U1713 ( .A(n2975), .B(n2976), .Z(n3240) );
  XNOR U1714 ( .A(n2307), .B(n2306), .Z(n2247) );
  XOR U1715 ( .A(n3052), .B(n3053), .Z(n3321) );
  XOR U1716 ( .A(n3042), .B(n3043), .Z(n3306) );
  XOR U1717 ( .A(n3290), .B(n3291), .Z(n3687) );
  XOR U1718 ( .A(n3233), .B(n3234), .Z(n3628) );
  XOR U1719 ( .A(n2255), .B(n2254), .Z(n2295) );
  XOR U1720 ( .A(n2389), .B(n2388), .Z(n2391) );
  XOR U1721 ( .A(n2351), .B(n2350), .Z(n2367) );
  XOR U1722 ( .A(n3308), .B(n3309), .Z(n3702) );
  XOR U1723 ( .A(n3696), .B(n3697), .Z(n3849) );
  XOR U1724 ( .A(n3294), .B(n3295), .Z(n3691) );
  XOR U1725 ( .A(n3251), .B(n3252), .Z(n3644) );
  XOR U1726 ( .A(n2237), .B(n2236), .Z(n2228) );
  XOR U1727 ( .A(n2705), .B(n2704), .Z(n2620) );
  XOR U1728 ( .A(n2693), .B(n2692), .Z(n2633) );
  XOR U1729 ( .A(n2766), .B(n2765), .Z(n2782) );
  XNOR U1730 ( .A(n3755), .B(n3756), .Z(n3861) );
  XOR U1731 ( .A(n3666), .B(n3667), .Z(n3669) );
  XOR U1732 ( .A(n3792), .B(n3793), .Z(n3795) );
  XOR U1733 ( .A(n3126), .B(n3125), .Z(n3166) );
  XOR U1734 ( .A(n3219), .B(n3220), .Z(n3337) );
  XOR U1735 ( .A(n3884), .B(n3885), .Z(n4058) );
  XOR U1736 ( .A(n3872), .B(n3873), .Z(n4046) );
  XOR U1737 ( .A(n3680), .B(n3681), .Z(n3831) );
  XOR U1738 ( .A(n3826), .B(n3827), .Z(n3998) );
  XOR U1739 ( .A(n3816), .B(n3817), .Z(n3984) );
  XOR U1740 ( .A(n3656), .B(n3657), .Z(n3811) );
  XOR U1741 ( .A(n3806), .B(n3807), .Z(n3972) );
  XOR U1742 ( .A(n3786), .B(n3787), .Z(n3789) );
  XOR U1743 ( .A(n3776), .B(n3777), .Z(n3924) );
  XOR U1744 ( .A(n3770), .B(n3771), .Z(n3939) );
  XOR U1745 ( .A(n2816), .B(n2815), .Z(n2818) );
  XOR U1746 ( .A(n2748), .B(n2747), .Z(n2804) );
  XOR U1747 ( .A(n3190), .B(n3189), .Z(n3105) );
  XOR U1748 ( .A(n3397), .B(n3396), .Z(n3490) );
  XOR U1749 ( .A(n3178), .B(n3177), .Z(n3117) );
  XOR U1750 ( .A(n3844), .B(n3845), .Z(n4013) );
  XOR U1751 ( .A(n3896), .B(n3897), .Z(n4068) );
  XOR U1752 ( .A(n3519), .B(n3520), .Z(n3518) );
  XOR U1753 ( .A(n4117), .B(n4118), .Z(n4120) );
  XOR U1754 ( .A(n3579), .B(n3578), .Z(n3577) );
  XOR U1755 ( .A(n4051), .B(n4052), .Z(n4216) );
  XOR U1756 ( .A(n4039), .B(n4040), .Z(n4203) );
  XOR U1757 ( .A(n4027), .B(n4028), .Z(n4192) );
  XOR U1758 ( .A(n4003), .B(n4004), .Z(n4167) );
  XOR U1759 ( .A(n3991), .B(n3992), .Z(n4156) );
  XOR U1760 ( .A(n3979), .B(n3980), .Z(n4145) );
  XOR U1761 ( .A(n3967), .B(n3968), .Z(n4136) );
  XOR U1762 ( .A(n3935), .B(n3936), .Z(n4099) );
  XOR U1763 ( .A(n4075), .B(n4076), .Z(n4240) );
  XOR U1764 ( .A(n3911), .B(n3910), .Z(n3907) );
  XOR U1765 ( .A(n4241), .B(n4242), .Z(n4411) );
  XOR U1766 ( .A(n4229), .B(n4230), .Z(n4401) );
  XOR U1767 ( .A(n4217), .B(n4218), .Z(n4391) );
  XOR U1768 ( .A(n4205), .B(n4206), .Z(n4381) );
  XOR U1769 ( .A(n4193), .B(n4194), .Z(n4371) );
  XOR U1770 ( .A(n4181), .B(n4182), .Z(n4361) );
  XOR U1771 ( .A(n4169), .B(n4170), .Z(n4351) );
  XOR U1772 ( .A(n4157), .B(n4158), .Z(n4341) );
  XOR U1773 ( .A(n4147), .B(n4148), .Z(n4331) );
  XOR U1774 ( .A(n4137), .B(n4138), .Z(n4319) );
  XOR U1775 ( .A(n4123), .B(n4124), .Z(n4310) );
  XOR U1776 ( .A(n4113), .B(n4114), .Z(n4297) );
  XOR U1777 ( .A(n4101), .B(n4102), .Z(n4287) );
  XOR U1778 ( .A(n4409), .B(n4410), .Z(n4517) );
  XOR U1779 ( .A(n4399), .B(n4400), .Z(n4593) );
  XOR U1780 ( .A(n4389), .B(n4390), .Z(n4669) );
  XOR U1781 ( .A(n4379), .B(n4380), .Z(n4745) );
  XOR U1782 ( .A(n4369), .B(n4370), .Z(n4821) );
  XOR U1783 ( .A(n4359), .B(n4360), .Z(n4897) );
  XOR U1784 ( .A(n4349), .B(n4350), .Z(n4973) );
  XOR U1785 ( .A(n4339), .B(n4340), .Z(n5050) );
  XOR U1786 ( .A(n4329), .B(n4330), .Z(n5128) );
  XOR U1787 ( .A(n4317), .B(n4318), .Z(n5204) );
  XOR U1788 ( .A(n4307), .B(n4308), .Z(n5280) );
  XOR U1789 ( .A(n4295), .B(n4296), .Z(n5358) );
  XOR U1790 ( .A(n4285), .B(n4286), .Z(n5435) );
  XOR U1791 ( .A(n4275), .B(n4276), .Z(n5511) );
  NAND U1792 ( .A(n5594), .B(o[2]), .Z(n1491) );
  NANDN U1793 ( .A(n5598), .B(n1491), .Z(n1492) );
  NAND U1794 ( .A(\stack[1][2] ), .B(n1492), .Z(n1493) );
  NAND U1795 ( .A(x[2]), .B(n5603), .Z(n1494) );
  AND U1796 ( .A(n1493), .B(n1494), .Z(n1495) );
  XOR U1797 ( .A(\DP_OP_25_64_5665/n299 ), .B(\DP_OP_25_64_5665/n267 ), .Z(
        n1496) );
  AND U1798 ( .A(n1601), .B(n1496), .Z(n1497) );
  ANDN U1799 ( .B(n1495), .A(n1497), .Z(n1498) );
  NANDN U1800 ( .A(n5597), .B(o[2]), .Z(n1499) );
  NAND U1801 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U1802 ( .A(n5547), .B(n5546), .Z(n1501) );
  NAND U1803 ( .A(n5578), .B(n1501), .Z(n1502) );
  NANDN U1804 ( .A(n1500), .B(n1502), .Z(n1308) );
  ANDN U1805 ( .B(opcode[0]), .A(opcode[1]), .Z(n1570) );
  ANDN U1806 ( .B(n1570), .A(opcode[2]), .Z(n1604) );
  ANDN U1807 ( .B(opcode[1]), .A(opcode[0]), .Z(n1603) );
  NANDN U1808 ( .A(opcode[2]), .B(n1603), .Z(n1569) );
  NANDN U1809 ( .A(n1604), .B(n1569), .Z(n1565) );
  AND U1810 ( .A(o[31]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_31 ) );
  AND U1811 ( .A(o[30]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_30 ) );
  AND U1812 ( .A(o[29]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_29 ) );
  AND U1813 ( .A(o[28]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_28 ) );
  AND U1814 ( .A(o[27]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_27 ) );
  AND U1815 ( .A(o[26]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_26 ) );
  AND U1816 ( .A(o[25]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_25 ) );
  AND U1817 ( .A(o[24]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_24 ) );
  AND U1818 ( .A(o[23]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_23 ) );
  AND U1819 ( .A(o[22]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_22 ) );
  AND U1820 ( .A(o[21]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_21 ) );
  AND U1821 ( .A(o[20]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_20 ) );
  AND U1822 ( .A(o[19]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_19 ) );
  AND U1823 ( .A(o[18]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_18 ) );
  AND U1824 ( .A(o[17]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_17 ) );
  AND U1825 ( .A(o[16]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_16 ) );
  AND U1826 ( .A(o[15]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U1827 ( .A(o[14]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U1828 ( .A(o[13]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U1829 ( .A(o[12]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U1830 ( .A(o[11]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U1831 ( .A(o[10]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U1832 ( .A(o[9]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U1833 ( .A(o[8]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U1834 ( .A(o[7]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U1835 ( .A(o[6]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U1836 ( .A(o[5]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U1837 ( .A(o[4]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U1838 ( .A(o[3]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U1839 ( .A(o[2]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U1840 ( .A(o[1]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U1841 ( .A(o[0]), .B(n1565), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U1842 ( .A(n1570), .B(opcode[2]), .Z(n1568) );
  NAND U1843 ( .A(n1568), .B(o[31]), .Z(n1504) );
  NAND U1844 ( .A(\stack[1][31] ), .B(n1565), .Z(n1503) );
  NAND U1845 ( .A(n1504), .B(n1503), .Z(\U1/RSOP_16/C3/Z_31 ) );
  NAND U1846 ( .A(n1568), .B(o[30]), .Z(n1506) );
  NAND U1847 ( .A(\stack[1][30] ), .B(n1565), .Z(n1505) );
  NAND U1848 ( .A(n1506), .B(n1505), .Z(\U1/RSOP_16/C3/Z_30 ) );
  NAND U1849 ( .A(n1568), .B(o[29]), .Z(n1508) );
  NAND U1850 ( .A(\stack[1][29] ), .B(n1565), .Z(n1507) );
  NAND U1851 ( .A(n1508), .B(n1507), .Z(\U1/RSOP_16/C3/Z_29 ) );
  NAND U1852 ( .A(n1568), .B(o[28]), .Z(n1510) );
  NAND U1853 ( .A(\stack[1][28] ), .B(n1565), .Z(n1509) );
  NAND U1854 ( .A(n1510), .B(n1509), .Z(\U1/RSOP_16/C3/Z_28 ) );
  NAND U1855 ( .A(n1568), .B(o[27]), .Z(n1512) );
  NAND U1856 ( .A(\stack[1][27] ), .B(n1565), .Z(n1511) );
  NAND U1857 ( .A(n1512), .B(n1511), .Z(\U1/RSOP_16/C3/Z_27 ) );
  NAND U1858 ( .A(n1568), .B(o[26]), .Z(n1514) );
  NAND U1859 ( .A(\stack[1][26] ), .B(n1565), .Z(n1513) );
  NAND U1860 ( .A(n1514), .B(n1513), .Z(\U1/RSOP_16/C3/Z_26 ) );
  NAND U1861 ( .A(n1568), .B(o[25]), .Z(n1516) );
  NAND U1862 ( .A(\stack[1][25] ), .B(n1565), .Z(n1515) );
  NAND U1863 ( .A(n1516), .B(n1515), .Z(\U1/RSOP_16/C3/Z_25 ) );
  NAND U1864 ( .A(n1568), .B(o[24]), .Z(n1518) );
  NAND U1865 ( .A(\stack[1][24] ), .B(n1565), .Z(n1517) );
  NAND U1866 ( .A(n1518), .B(n1517), .Z(\U1/RSOP_16/C3/Z_24 ) );
  NAND U1867 ( .A(n1568), .B(o[23]), .Z(n1520) );
  NAND U1868 ( .A(\stack[1][23] ), .B(n1565), .Z(n1519) );
  NAND U1869 ( .A(n1520), .B(n1519), .Z(\U1/RSOP_16/C3/Z_23 ) );
  NAND U1870 ( .A(n1568), .B(o[22]), .Z(n1522) );
  NAND U1871 ( .A(\stack[1][22] ), .B(n1565), .Z(n1521) );
  NAND U1872 ( .A(n1522), .B(n1521), .Z(\U1/RSOP_16/C3/Z_22 ) );
  NAND U1873 ( .A(n1568), .B(o[21]), .Z(n1524) );
  NAND U1874 ( .A(\stack[1][21] ), .B(n1565), .Z(n1523) );
  NAND U1875 ( .A(n1524), .B(n1523), .Z(\U1/RSOP_16/C3/Z_21 ) );
  NAND U1876 ( .A(n1568), .B(o[20]), .Z(n1526) );
  NAND U1877 ( .A(\stack[1][20] ), .B(n1565), .Z(n1525) );
  NAND U1878 ( .A(n1526), .B(n1525), .Z(\U1/RSOP_16/C3/Z_20 ) );
  NAND U1879 ( .A(n1568), .B(o[19]), .Z(n1528) );
  NAND U1880 ( .A(\stack[1][19] ), .B(n1565), .Z(n1527) );
  NAND U1881 ( .A(n1528), .B(n1527), .Z(\U1/RSOP_16/C3/Z_19 ) );
  NAND U1882 ( .A(n1568), .B(o[18]), .Z(n1530) );
  NAND U1883 ( .A(\stack[1][18] ), .B(n1565), .Z(n1529) );
  NAND U1884 ( .A(n1530), .B(n1529), .Z(\U1/RSOP_16/C3/Z_18 ) );
  NAND U1885 ( .A(n1568), .B(o[17]), .Z(n1532) );
  NAND U1886 ( .A(\stack[1][17] ), .B(n1565), .Z(n1531) );
  NAND U1887 ( .A(n1532), .B(n1531), .Z(\U1/RSOP_16/C3/Z_17 ) );
  NAND U1888 ( .A(n1568), .B(o[16]), .Z(n1534) );
  NAND U1889 ( .A(\stack[1][16] ), .B(n1565), .Z(n1533) );
  NAND U1890 ( .A(n1534), .B(n1533), .Z(\U1/RSOP_16/C3/Z_16 ) );
  NAND U1891 ( .A(n1568), .B(o[15]), .Z(n1536) );
  NAND U1892 ( .A(\stack[1][15] ), .B(n1565), .Z(n1535) );
  NAND U1893 ( .A(n1536), .B(n1535), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U1894 ( .A(n1568), .B(o[14]), .Z(n1538) );
  NAND U1895 ( .A(\stack[1][14] ), .B(n1565), .Z(n1537) );
  NAND U1896 ( .A(n1538), .B(n1537), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U1897 ( .A(n1568), .B(o[13]), .Z(n1540) );
  NAND U1898 ( .A(\stack[1][13] ), .B(n1565), .Z(n1539) );
  NAND U1899 ( .A(n1540), .B(n1539), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U1900 ( .A(n1568), .B(o[12]), .Z(n1542) );
  NAND U1901 ( .A(\stack[1][12] ), .B(n1565), .Z(n1541) );
  NAND U1902 ( .A(n1542), .B(n1541), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U1903 ( .A(n1568), .B(o[11]), .Z(n1544) );
  NAND U1904 ( .A(\stack[1][11] ), .B(n1565), .Z(n1543) );
  NAND U1905 ( .A(n1544), .B(n1543), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U1906 ( .A(n1568), .B(o[10]), .Z(n1546) );
  NAND U1907 ( .A(\stack[1][10] ), .B(n1565), .Z(n1545) );
  NAND U1908 ( .A(n1546), .B(n1545), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U1909 ( .A(n1568), .B(o[9]), .Z(n1548) );
  NAND U1910 ( .A(\stack[1][9] ), .B(n1565), .Z(n1547) );
  NAND U1911 ( .A(n1548), .B(n1547), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U1912 ( .A(n1568), .B(o[8]), .Z(n1550) );
  NAND U1913 ( .A(\stack[1][8] ), .B(n1565), .Z(n1549) );
  NAND U1914 ( .A(n1550), .B(n1549), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U1915 ( .A(n1568), .B(o[7]), .Z(n1552) );
  NAND U1916 ( .A(\stack[1][7] ), .B(n1565), .Z(n1551) );
  NAND U1917 ( .A(n1552), .B(n1551), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U1918 ( .A(n1568), .B(o[6]), .Z(n1554) );
  NAND U1919 ( .A(\stack[1][6] ), .B(n1565), .Z(n1553) );
  NAND U1920 ( .A(n1554), .B(n1553), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U1921 ( .A(n1568), .B(o[5]), .Z(n1556) );
  NAND U1922 ( .A(\stack[1][5] ), .B(n1565), .Z(n1555) );
  NAND U1923 ( .A(n1556), .B(n1555), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U1924 ( .A(n1568), .B(o[4]), .Z(n1558) );
  NAND U1925 ( .A(\stack[1][4] ), .B(n1565), .Z(n1557) );
  NAND U1926 ( .A(n1558), .B(n1557), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U1927 ( .A(n1568), .B(o[3]), .Z(n1560) );
  NAND U1928 ( .A(\stack[1][3] ), .B(n1565), .Z(n1559) );
  NAND U1929 ( .A(n1560), .B(n1559), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U1930 ( .A(n1568), .B(o[2]), .Z(n1562) );
  NAND U1931 ( .A(\stack[1][2] ), .B(n1565), .Z(n1561) );
  NAND U1932 ( .A(n1562), .B(n1561), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U1933 ( .A(n1568), .B(o[1]), .Z(n1564) );
  NAND U1934 ( .A(\stack[1][1] ), .B(n1565), .Z(n1563) );
  NAND U1935 ( .A(n1564), .B(n1563), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U1936 ( .A(n1568), .B(o[0]), .Z(n1567) );
  NAND U1937 ( .A(\stack[1][0] ), .B(n1565), .Z(n1566) );
  NAND U1938 ( .A(n1567), .B(n1566), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U1939 ( .A(n1568), .B(n1569), .Z(\C1/Z_0 ) );
  NANDN U1940 ( .A(n1570), .B(n1569), .Z(n1601) );
  NAND U1941 ( .A(\C3/DATA5_31 ), .B(n1601), .Z(n1571) );
  ANDN U1942 ( .B(n1571), .A(n4448), .Z(n4449) );
  NAND U1943 ( .A(\C3/DATA5_30 ), .B(n1601), .Z(n1572) );
  AND U1944 ( .A(n4479), .B(n1572), .Z(n4484) );
  NAND U1945 ( .A(\C3/DATA5_29 ), .B(n1601), .Z(n1573) );
  ANDN U1946 ( .B(n1573), .A(n4524), .Z(n4525) );
  NAND U1947 ( .A(\C3/DATA5_28 ), .B(n1601), .Z(n1574) );
  AND U1948 ( .A(n4555), .B(n1574), .Z(n4560) );
  NAND U1949 ( .A(\C3/DATA5_27 ), .B(n1601), .Z(n1575) );
  ANDN U1950 ( .B(n1575), .A(n4600), .Z(n4601) );
  NAND U1951 ( .A(\C3/DATA5_26 ), .B(n1601), .Z(n1576) );
  AND U1952 ( .A(n4631), .B(n1576), .Z(n4636) );
  NAND U1953 ( .A(\C3/DATA5_25 ), .B(n1601), .Z(n1577) );
  ANDN U1954 ( .B(n1577), .A(n4676), .Z(n4677) );
  NAND U1955 ( .A(\C3/DATA5_24 ), .B(n1601), .Z(n1578) );
  AND U1956 ( .A(n4707), .B(n1578), .Z(n4712) );
  NAND U1957 ( .A(\C3/DATA5_23 ), .B(n1601), .Z(n1579) );
  ANDN U1958 ( .B(n1579), .A(n4752), .Z(n4753) );
  NAND U1959 ( .A(\C3/DATA5_22 ), .B(n1601), .Z(n1580) );
  AND U1960 ( .A(n4783), .B(n1580), .Z(n4788) );
  NAND U1961 ( .A(\C3/DATA5_21 ), .B(n1601), .Z(n1581) );
  ANDN U1962 ( .B(n1581), .A(n4828), .Z(n4829) );
  NAND U1963 ( .A(\C3/DATA5_20 ), .B(n1601), .Z(n1582) );
  AND U1964 ( .A(n4859), .B(n1582), .Z(n4864) );
  NAND U1965 ( .A(\C3/DATA5_19 ), .B(n1601), .Z(n1583) );
  ANDN U1966 ( .B(n1583), .A(n4904), .Z(n4905) );
  NAND U1967 ( .A(\C3/DATA5_18 ), .B(n1601), .Z(n1584) );
  AND U1968 ( .A(n4935), .B(n1584), .Z(n4940) );
  NAND U1969 ( .A(\C3/DATA5_17 ), .B(n1601), .Z(n1585) );
  ANDN U1970 ( .B(n1585), .A(n4980), .Z(n4981) );
  NAND U1971 ( .A(\C3/DATA5_16 ), .B(n1601), .Z(n1586) );
  AND U1972 ( .A(n5011), .B(n1586), .Z(n5016) );
  NAND U1973 ( .A(\C3/DATA5_15 ), .B(n1601), .Z(n1587) );
  ANDN U1974 ( .B(n1587), .A(n5057), .Z(n5058) );
  NAND U1975 ( .A(\C3/DATA5_14 ), .B(n1601), .Z(n1588) );
  AND U1976 ( .A(n5089), .B(n1588), .Z(n5094) );
  NAND U1977 ( .A(\C3/DATA5_13 ), .B(n1601), .Z(n1589) );
  AND U1978 ( .A(n5127), .B(n1589), .Z(n5132) );
  NAND U1979 ( .A(\C3/DATA5_12 ), .B(n1601), .Z(n1590) );
  AND U1980 ( .A(n5165), .B(n1590), .Z(n5170) );
  NAND U1981 ( .A(\C3/DATA5_11 ), .B(n1601), .Z(n1591) );
  AND U1982 ( .A(n5203), .B(n1591), .Z(n5208) );
  NAND U1983 ( .A(\C3/DATA5_10 ), .B(n1601), .Z(n1592) );
  AND U1984 ( .A(n5241), .B(n1592), .Z(n5246) );
  NAND U1985 ( .A(\C3/DATA5_9 ), .B(n1601), .Z(n1593) );
  AND U1986 ( .A(n5279), .B(n1593), .Z(n5284) );
  NAND U1987 ( .A(\C3/DATA5_8 ), .B(n1601), .Z(n1594) );
  AND U1988 ( .A(n5318), .B(n1594), .Z(n5323) );
  NAND U1989 ( .A(\C3/DATA5_7 ), .B(n1601), .Z(n1595) );
  AND U1990 ( .A(n5357), .B(n1595), .Z(n5362) );
  NAND U1991 ( .A(\C3/DATA5_6 ), .B(n1601), .Z(n1596) );
  AND U1992 ( .A(n5396), .B(n1596), .Z(n5401) );
  NAND U1993 ( .A(\C3/DATA5_5 ), .B(n1601), .Z(n1597) );
  AND U1994 ( .A(n5434), .B(n1597), .Z(n5439) );
  NAND U1995 ( .A(\C3/DATA5_4 ), .B(n1601), .Z(n1598) );
  AND U1996 ( .A(n5472), .B(n1598), .Z(n5477) );
  NAND U1997 ( .A(\C3/DATA5_3 ), .B(n1601), .Z(n1599) );
  AND U1998 ( .A(n5510), .B(n1599), .Z(n5515) );
  NAND U1999 ( .A(\C3/DATA5_1 ), .B(n1601), .Z(n1600) );
  NAND U2000 ( .A(n5574), .B(n1600), .Z(n5587) );
  NAND U2001 ( .A(\C3/DATA5_0 ), .B(n1601), .Z(n1602) );
  AND U2002 ( .A(n5604), .B(n1602), .Z(n5605) );
  ANDN U2003 ( .B(opcode[2]), .A(opcode[0]), .Z(n1609) );
  ANDN U2004 ( .B(n1609), .A(opcode[1]), .Z(n5603) );
  NAND U2005 ( .A(\stack[6][0] ), .B(n5603), .Z(n1606) );
  NANDN U2006 ( .A(n5603), .B(\stack[7][0] ), .Z(n1605) );
  NAND U2007 ( .A(n1606), .B(n1605), .Z(n1063) );
  NAND U2008 ( .A(\stack[5][0] ), .B(n5603), .Z(n1608) );
  NOR U2009 ( .A(opcode[1]), .B(n1604), .Z(n5588) );
  NANDN U2010 ( .A(n5588), .B(\stack[7][0] ), .Z(n1607) );
  AND U2011 ( .A(n1608), .B(n1607), .Z(n1611) );
  ANDN U2012 ( .B(n5588), .A(n1609), .Z(n5591) );
  NAND U2013 ( .A(n5591), .B(\stack[6][0] ), .Z(n1610) );
  NAND U2014 ( .A(n1611), .B(n1610), .Z(n1064) );
  NAND U2015 ( .A(\stack[4][0] ), .B(n5603), .Z(n1613) );
  NANDN U2016 ( .A(n5588), .B(\stack[6][0] ), .Z(n1612) );
  AND U2017 ( .A(n1613), .B(n1612), .Z(n1615) );
  NAND U2018 ( .A(n5591), .B(\stack[5][0] ), .Z(n1614) );
  NAND U2019 ( .A(n1615), .B(n1614), .Z(n1065) );
  NAND U2020 ( .A(\stack[3][0] ), .B(n5603), .Z(n1617) );
  NANDN U2021 ( .A(n5588), .B(\stack[5][0] ), .Z(n1616) );
  AND U2022 ( .A(n1617), .B(n1616), .Z(n1619) );
  NAND U2023 ( .A(n5591), .B(\stack[4][0] ), .Z(n1618) );
  NAND U2024 ( .A(n1619), .B(n1618), .Z(n1066) );
  NAND U2025 ( .A(\stack[2][0] ), .B(n5603), .Z(n1621) );
  NANDN U2026 ( .A(n5588), .B(\stack[4][0] ), .Z(n1620) );
  AND U2027 ( .A(n1621), .B(n1620), .Z(n1623) );
  NAND U2028 ( .A(n5591), .B(\stack[3][0] ), .Z(n1622) );
  NAND U2029 ( .A(n1623), .B(n1622), .Z(n1067) );
  NAND U2030 ( .A(n5603), .B(\stack[1][0] ), .Z(n1625) );
  NANDN U2031 ( .A(n5588), .B(\stack[3][0] ), .Z(n1624) );
  AND U2032 ( .A(n1625), .B(n1624), .Z(n1627) );
  NAND U2033 ( .A(n5591), .B(\stack[2][0] ), .Z(n1626) );
  NAND U2034 ( .A(n1627), .B(n1626), .Z(n1068) );
  NAND U2035 ( .A(\stack[6][31] ), .B(n5603), .Z(n1629) );
  NANDN U2036 ( .A(n5603), .B(\stack[7][31] ), .Z(n1628) );
  NAND U2037 ( .A(n1629), .B(n1628), .Z(n1069) );
  NAND U2038 ( .A(\stack[5][31] ), .B(n5603), .Z(n1631) );
  NANDN U2039 ( .A(n5588), .B(\stack[7][31] ), .Z(n1630) );
  AND U2040 ( .A(n1631), .B(n1630), .Z(n1633) );
  NAND U2041 ( .A(n5591), .B(\stack[6][31] ), .Z(n1632) );
  NAND U2042 ( .A(n1633), .B(n1632), .Z(n1070) );
  NAND U2043 ( .A(\stack[4][31] ), .B(n5603), .Z(n1635) );
  NANDN U2044 ( .A(n5588), .B(\stack[6][31] ), .Z(n1634) );
  AND U2045 ( .A(n1635), .B(n1634), .Z(n1637) );
  NAND U2046 ( .A(n5591), .B(\stack[5][31] ), .Z(n1636) );
  NAND U2047 ( .A(n1637), .B(n1636), .Z(n1071) );
  NAND U2048 ( .A(\stack[3][31] ), .B(n5603), .Z(n1639) );
  NANDN U2049 ( .A(n5588), .B(\stack[5][31] ), .Z(n1638) );
  AND U2050 ( .A(n1639), .B(n1638), .Z(n1641) );
  NAND U2051 ( .A(n5591), .B(\stack[4][31] ), .Z(n1640) );
  NAND U2052 ( .A(n1641), .B(n1640), .Z(n1072) );
  NAND U2053 ( .A(\stack[2][31] ), .B(n5603), .Z(n1643) );
  NANDN U2054 ( .A(n5588), .B(\stack[4][31] ), .Z(n1642) );
  AND U2055 ( .A(n1643), .B(n1642), .Z(n1645) );
  NAND U2056 ( .A(n5591), .B(\stack[3][31] ), .Z(n1644) );
  NAND U2057 ( .A(n1645), .B(n1644), .Z(n1073) );
  NAND U2058 ( .A(n5603), .B(\stack[1][31] ), .Z(n1647) );
  NANDN U2059 ( .A(n5588), .B(\stack[3][31] ), .Z(n1646) );
  AND U2060 ( .A(n1647), .B(n1646), .Z(n1649) );
  NAND U2061 ( .A(n5591), .B(\stack[2][31] ), .Z(n1648) );
  NAND U2062 ( .A(n1649), .B(n1648), .Z(n1074) );
  NAND U2063 ( .A(n5603), .B(o[31]), .Z(n1651) );
  NANDN U2064 ( .A(n5588), .B(\stack[2][31] ), .Z(n1650) );
  AND U2065 ( .A(n1651), .B(n1650), .Z(n1653) );
  NAND U2066 ( .A(\stack[1][31] ), .B(n5591), .Z(n1652) );
  NAND U2067 ( .A(n1653), .B(n1652), .Z(n1075) );
  AND U2068 ( .A(opcode[1]), .B(opcode[0]), .Z(n5595) );
  ANDN U2069 ( .B(n5595), .A(opcode[2]), .Z(n5578) );
  AND U2070 ( .A(\stack[1][8] ), .B(o[21]), .Z(n3089) );
  AND U2071 ( .A(\stack[1][8] ), .B(o[20]), .Z(n2612) );
  AND U2072 ( .A(\stack[1][10] ), .B(o[17]), .Z(n2617) );
  AND U2073 ( .A(\stack[1][12] ), .B(o[12]), .Z(n2006) );
  AND U2074 ( .A(o[8]), .B(\stack[1][14] ), .Z(n1760) );
  AND U2075 ( .A(o[6]), .B(\stack[1][15] ), .Z(n1793) );
  AND U2076 ( .A(o[1]), .B(\stack[1][19] ), .Z(n1671) );
  NAND U2077 ( .A(\stack[1][20] ), .B(o[0]), .Z(n1654) );
  XNOR U2078 ( .A(n1671), .B(n1654), .Z(n1675) );
  NAND U2079 ( .A(n1671), .B(o[0]), .Z(n1655) );
  XNOR U2080 ( .A(o[2]), .B(n1655), .Z(n1656) );
  AND U2081 ( .A(\stack[1][18] ), .B(n1656), .Z(n1674) );
  XOR U2082 ( .A(n1675), .B(n1674), .Z(n1664) );
  AND U2083 ( .A(o[0]), .B(\stack[1][17] ), .Z(n1657) );
  AND U2084 ( .A(o[1]), .B(\stack[1][18] ), .Z(n1661) );
  AND U2085 ( .A(n1657), .B(n1661), .Z(n1658) );
  NAND U2086 ( .A(o[2]), .B(n1658), .Z(n1663) );
  NAND U2087 ( .A(n1661), .B(o[0]), .Z(n1659) );
  XNOR U2088 ( .A(o[2]), .B(n1659), .Z(n1660) );
  AND U2089 ( .A(\stack[1][17] ), .B(n1660), .Z(n1679) );
  AND U2090 ( .A(o[0]), .B(\stack[1][19] ), .Z(n1769) );
  XOR U2091 ( .A(n1661), .B(n1769), .Z(n1678) );
  NAND U2092 ( .A(n1679), .B(n1678), .Z(n1662) );
  NAND U2093 ( .A(n1663), .B(n1662), .Z(n1665) );
  NAND U2094 ( .A(n1664), .B(n1665), .Z(n1667) );
  XOR U2095 ( .A(n1665), .B(n1664), .Z(n1692) );
  AND U2096 ( .A(o[3]), .B(\stack[1][17] ), .Z(n1693) );
  NAND U2097 ( .A(n1692), .B(n1693), .Z(n1666) );
  NAND U2098 ( .A(n1667), .B(n1666), .Z(n1762) );
  AND U2099 ( .A(o[4]), .B(\stack[1][17] ), .Z(n1763) );
  XOR U2100 ( .A(n1762), .B(n1763), .Z(n1765) );
  AND U2101 ( .A(o[1]), .B(\stack[1][20] ), .Z(n1768) );
  NAND U2102 ( .A(\stack[1][21] ), .B(o[0]), .Z(n1668) );
  XNOR U2103 ( .A(n1768), .B(n1668), .Z(n1772) );
  NAND U2104 ( .A(n1768), .B(o[0]), .Z(n1669) );
  XNOR U2105 ( .A(o[2]), .B(n1669), .Z(n1670) );
  AND U2106 ( .A(\stack[1][19] ), .B(n1670), .Z(n1771) );
  XOR U2107 ( .A(n1772), .B(n1771), .Z(n1779) );
  AND U2108 ( .A(o[0]), .B(\stack[1][18] ), .Z(n1672) );
  AND U2109 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U2110 ( .A(o[2]), .B(n1673), .Z(n1677) );
  NAND U2111 ( .A(n1675), .B(n1674), .Z(n1676) );
  NAND U2112 ( .A(n1677), .B(n1676), .Z(n1778) );
  XOR U2113 ( .A(n1779), .B(n1778), .Z(n1781) );
  AND U2114 ( .A(o[3]), .B(\stack[1][18] ), .Z(n1780) );
  XOR U2115 ( .A(n1781), .B(n1780), .Z(n1764) );
  XOR U2116 ( .A(n1765), .B(n1764), .Z(n1785) );
  AND U2117 ( .A(o[5]), .B(\stack[1][16] ), .Z(n1784) );
  XOR U2118 ( .A(n1785), .B(n1784), .Z(n1787) );
  AND U2119 ( .A(o[4]), .B(\stack[1][16] ), .Z(n1695) );
  XOR U2120 ( .A(n1679), .B(n1678), .Z(n1689) );
  AND U2121 ( .A(o[0]), .B(\stack[1][16] ), .Z(n1680) );
  AND U2122 ( .A(o[1]), .B(\stack[1][17] ), .Z(n1683) );
  AND U2123 ( .A(n1680), .B(n1683), .Z(n1681) );
  NAND U2124 ( .A(o[2]), .B(n1681), .Z(n1687) );
  NAND U2125 ( .A(\stack[1][18] ), .B(o[0]), .Z(n1682) );
  XNOR U2126 ( .A(n1683), .B(n1682), .Z(n1699) );
  NAND U2127 ( .A(n1683), .B(o[0]), .Z(n1684) );
  XNOR U2128 ( .A(o[2]), .B(n1684), .Z(n1685) );
  AND U2129 ( .A(\stack[1][16] ), .B(n1685), .Z(n1698) );
  NAND U2130 ( .A(n1699), .B(n1698), .Z(n1686) );
  NAND U2131 ( .A(n1687), .B(n1686), .Z(n1688) );
  NAND U2132 ( .A(n1689), .B(n1688), .Z(n1691) );
  XOR U2133 ( .A(n1689), .B(n1688), .Z(n1713) );
  AND U2134 ( .A(o[3]), .B(\stack[1][16] ), .Z(n1712) );
  NAND U2135 ( .A(n1713), .B(n1712), .Z(n1690) );
  NAND U2136 ( .A(n1691), .B(n1690), .Z(n1694) );
  NAND U2137 ( .A(n1695), .B(n1694), .Z(n1697) );
  XOR U2138 ( .A(n1695), .B(n1694), .Z(n1718) );
  NAND U2139 ( .A(n1719), .B(n1718), .Z(n1696) );
  NAND U2140 ( .A(n1697), .B(n1696), .Z(n1786) );
  XOR U2141 ( .A(n1787), .B(n1786), .Z(n1791) );
  XOR U2142 ( .A(n1699), .B(n1698), .Z(n1708) );
  AND U2143 ( .A(o[0]), .B(\stack[1][15] ), .Z(n1700) );
  AND U2144 ( .A(o[1]), .B(\stack[1][16] ), .Z(n1703) );
  AND U2145 ( .A(n1700), .B(n1703), .Z(n1701) );
  NAND U2146 ( .A(o[2]), .B(n1701), .Z(n1707) );
  NAND U2147 ( .A(\stack[1][17] ), .B(o[0]), .Z(n1702) );
  XNOR U2148 ( .A(n1703), .B(n1702), .Z(n1731) );
  NAND U2149 ( .A(n1703), .B(o[0]), .Z(n1704) );
  XNOR U2150 ( .A(o[2]), .B(n1704), .Z(n1705) );
  AND U2151 ( .A(\stack[1][15] ), .B(n1705), .Z(n1730) );
  NAND U2152 ( .A(n1731), .B(n1730), .Z(n1706) );
  NAND U2153 ( .A(n1707), .B(n1706), .Z(n1709) );
  NAND U2154 ( .A(n1708), .B(n1709), .Z(n1711) );
  XOR U2155 ( .A(n1709), .B(n1708), .Z(n1745) );
  AND U2156 ( .A(o[3]), .B(\stack[1][15] ), .Z(n1744) );
  NAND U2157 ( .A(n1745), .B(n1744), .Z(n1710) );
  AND U2158 ( .A(n1711), .B(n1710), .Z(n1715) );
  NAND U2159 ( .A(o[4]), .B(\stack[1][15] ), .Z(n1714) );
  NAND U2160 ( .A(n1715), .B(n1714), .Z(n1717) );
  XNOR U2161 ( .A(n1713), .B(n1712), .Z(n1726) );
  XOR U2162 ( .A(n1715), .B(n1714), .Z(n1727) );
  NAND U2163 ( .A(n1726), .B(n1727), .Z(n1716) );
  AND U2164 ( .A(n1717), .B(n1716), .Z(n1721) );
  XOR U2165 ( .A(n1719), .B(n1718), .Z(n1720) );
  NAND U2166 ( .A(n1721), .B(n1720), .Z(n1723) );
  XOR U2167 ( .A(n1721), .B(n1720), .Z(n1725) );
  AND U2168 ( .A(o[5]), .B(\stack[1][15] ), .Z(n1724) );
  NAND U2169 ( .A(n1725), .B(n1724), .Z(n1722) );
  NAND U2170 ( .A(n1723), .B(n1722), .Z(n1790) );
  XOR U2171 ( .A(n1791), .B(n1790), .Z(n1792) );
  XOR U2172 ( .A(n1793), .B(n1792), .Z(n1756) );
  XOR U2173 ( .A(n1725), .B(n1724), .Z(n1753) );
  AND U2174 ( .A(o[5]), .B(\stack[1][14] ), .Z(n1729) );
  NAND U2175 ( .A(n1728), .B(n1729), .Z(n1751) );
  AND U2176 ( .A(o[4]), .B(\stack[1][14] ), .Z(n1747) );
  XOR U2177 ( .A(n1731), .B(n1730), .Z(n1741) );
  AND U2178 ( .A(o[0]), .B(\stack[1][14] ), .Z(n1732) );
  AND U2179 ( .A(o[1]), .B(\stack[1][15] ), .Z(n1735) );
  AND U2180 ( .A(n1732), .B(n1735), .Z(n1733) );
  NAND U2181 ( .A(o[2]), .B(n1733), .Z(n1739) );
  NAND U2182 ( .A(\stack[1][16] ), .B(o[0]), .Z(n1734) );
  XNOR U2183 ( .A(n1735), .B(n1734), .Z(n1855) );
  NAND U2184 ( .A(n1735), .B(o[0]), .Z(n1736) );
  XNOR U2185 ( .A(o[2]), .B(n1736), .Z(n1737) );
  AND U2186 ( .A(\stack[1][14] ), .B(n1737), .Z(n1854) );
  NAND U2187 ( .A(n1855), .B(n1854), .Z(n1738) );
  NAND U2188 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U2189 ( .A(n1741), .B(n1740), .Z(n1743) );
  XOR U2190 ( .A(n1741), .B(n1740), .Z(n1863) );
  AND U2191 ( .A(o[3]), .B(\stack[1][14] ), .Z(n1862) );
  NAND U2192 ( .A(n1863), .B(n1862), .Z(n1742) );
  NAND U2193 ( .A(n1743), .B(n1742), .Z(n1746) );
  NAND U2194 ( .A(n1747), .B(n1746), .Z(n1749) );
  XOR U2195 ( .A(n1745), .B(n1744), .Z(n1845) );
  XOR U2196 ( .A(n1747), .B(n1746), .Z(n1844) );
  NAND U2197 ( .A(n1845), .B(n1844), .Z(n1748) );
  NAND U2198 ( .A(n1749), .B(n1748), .Z(n1842) );
  NAND U2199 ( .A(n1843), .B(n1842), .Z(n1750) );
  NAND U2200 ( .A(n1751), .B(n1750), .Z(n1752) );
  NAND U2201 ( .A(n1753), .B(n1752), .Z(n1755) );
  XOR U2202 ( .A(n1753), .B(n1752), .Z(n1841) );
  AND U2203 ( .A(o[6]), .B(\stack[1][14] ), .Z(n1840) );
  NAND U2204 ( .A(n1841), .B(n1840), .Z(n1754) );
  NAND U2205 ( .A(n1755), .B(n1754), .Z(n1757) );
  NAND U2206 ( .A(n1756), .B(n1757), .Z(n1759) );
  XOR U2207 ( .A(n1757), .B(n1756), .Z(n1878) );
  AND U2208 ( .A(o[7]), .B(\stack[1][14] ), .Z(n1879) );
  NAND U2209 ( .A(n1878), .B(n1879), .Z(n1758) );
  NAND U2210 ( .A(n1759), .B(n1758), .Z(n1761) );
  NAND U2211 ( .A(n1760), .B(n1761), .Z(n1797) );
  XOR U2212 ( .A(n1761), .B(n1760), .Z(n1838) );
  NAND U2213 ( .A(n1763), .B(n1762), .Z(n1767) );
  NAND U2214 ( .A(n1765), .B(n1764), .Z(n1766) );
  NAND U2215 ( .A(n1767), .B(n1766), .Z(n1826) );
  AND U2216 ( .A(n1769), .B(n1768), .Z(n1770) );
  NAND U2217 ( .A(o[2]), .B(n1770), .Z(n1774) );
  NAND U2218 ( .A(n1772), .B(n1771), .Z(n1773) );
  NAND U2219 ( .A(n1774), .B(n1773), .Z(n1804) );
  AND U2220 ( .A(o[1]), .B(\stack[1][21] ), .Z(n1813) );
  NAND U2221 ( .A(\stack[1][22] ), .B(o[0]), .Z(n1775) );
  XNOR U2222 ( .A(n1813), .B(n1775), .Z(n1817) );
  NAND U2223 ( .A(n1813), .B(o[0]), .Z(n1776) );
  XNOR U2224 ( .A(o[2]), .B(n1776), .Z(n1777) );
  AND U2225 ( .A(\stack[1][20] ), .B(n1777), .Z(n1816) );
  XOR U2226 ( .A(n1817), .B(n1816), .Z(n1805) );
  XOR U2227 ( .A(n1804), .B(n1805), .Z(n1807) );
  AND U2228 ( .A(o[3]), .B(\stack[1][19] ), .Z(n1806) );
  XOR U2229 ( .A(n1807), .B(n1806), .Z(n1823) );
  AND U2230 ( .A(o[4]), .B(\stack[1][18] ), .Z(n1821) );
  NAND U2231 ( .A(n1779), .B(n1778), .Z(n1783) );
  NAND U2232 ( .A(n1781), .B(n1780), .Z(n1782) );
  NAND U2233 ( .A(n1783), .B(n1782), .Z(n1820) );
  XOR U2234 ( .A(n1821), .B(n1820), .Z(n1822) );
  XOR U2235 ( .A(n1823), .B(n1822), .Z(n1827) );
  XOR U2236 ( .A(n1826), .B(n1827), .Z(n1829) );
  AND U2237 ( .A(o[5]), .B(\stack[1][17] ), .Z(n1828) );
  XOR U2238 ( .A(n1829), .B(n1828), .Z(n1799) );
  NAND U2239 ( .A(n1785), .B(n1784), .Z(n1789) );
  NAND U2240 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U2241 ( .A(n1789), .B(n1788), .Z(n1798) );
  XOR U2242 ( .A(n1799), .B(n1798), .Z(n1801) );
  AND U2243 ( .A(o[6]), .B(\stack[1][16] ), .Z(n1800) );
  XOR U2244 ( .A(n1801), .B(n1800), .Z(n1833) );
  NAND U2245 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U2246 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U2247 ( .A(n1795), .B(n1794), .Z(n1832) );
  XOR U2248 ( .A(n1833), .B(n1832), .Z(n1835) );
  AND U2249 ( .A(o[7]), .B(\stack[1][15] ), .Z(n1834) );
  XOR U2250 ( .A(n1835), .B(n1834), .Z(n1839) );
  NAND U2251 ( .A(n1838), .B(n1839), .Z(n1796) );
  AND U2252 ( .A(n1797), .B(n1796), .Z(n1954) );
  NAND U2253 ( .A(n1799), .B(n1798), .Z(n1803) );
  NAND U2254 ( .A(n1801), .B(n1800), .Z(n1802) );
  NAND U2255 ( .A(n1803), .B(n1802), .Z(n1994) );
  AND U2256 ( .A(o[6]), .B(\stack[1][17] ), .Z(n1991) );
  NAND U2257 ( .A(n1805), .B(n1804), .Z(n1809) );
  NAND U2258 ( .A(n1807), .B(n1806), .Z(n1808) );
  NAND U2259 ( .A(n1809), .B(n1808), .Z(n1960) );
  AND U2260 ( .A(o[4]), .B(\stack[1][19] ), .Z(n1961) );
  XOR U2261 ( .A(n1960), .B(n1961), .Z(n1963) );
  AND U2262 ( .A(o[1]), .B(\stack[1][22] ), .Z(n1966) );
  NAND U2263 ( .A(\stack[1][23] ), .B(o[0]), .Z(n1810) );
  XNOR U2264 ( .A(n1966), .B(n1810), .Z(n1970) );
  NAND U2265 ( .A(n1966), .B(o[0]), .Z(n1811) );
  XNOR U2266 ( .A(o[2]), .B(n1811), .Z(n1812) );
  AND U2267 ( .A(\stack[1][21] ), .B(n1812), .Z(n1969) );
  XOR U2268 ( .A(n1970), .B(n1969), .Z(n1977) );
  AND U2269 ( .A(o[0]), .B(\stack[1][20] ), .Z(n1814) );
  AND U2270 ( .A(n1814), .B(n1813), .Z(n1815) );
  NAND U2271 ( .A(o[2]), .B(n1815), .Z(n1819) );
  NAND U2272 ( .A(n1817), .B(n1816), .Z(n1818) );
  NAND U2273 ( .A(n1819), .B(n1818), .Z(n1976) );
  XOR U2274 ( .A(n1977), .B(n1976), .Z(n1979) );
  AND U2275 ( .A(o[3]), .B(\stack[1][20] ), .Z(n1978) );
  XOR U2276 ( .A(n1979), .B(n1978), .Z(n1962) );
  XOR U2277 ( .A(n1963), .B(n1962), .Z(n1983) );
  AND U2278 ( .A(o[5]), .B(\stack[1][18] ), .Z(n1982) );
  XOR U2279 ( .A(n1983), .B(n1982), .Z(n1985) );
  NAND U2280 ( .A(n1821), .B(n1820), .Z(n1825) );
  NAND U2281 ( .A(n1823), .B(n1822), .Z(n1824) );
  NAND U2282 ( .A(n1825), .B(n1824), .Z(n1984) );
  XOR U2283 ( .A(n1985), .B(n1984), .Z(n1989) );
  NAND U2284 ( .A(n1827), .B(n1826), .Z(n1831) );
  NAND U2285 ( .A(n1829), .B(n1828), .Z(n1830) );
  NAND U2286 ( .A(n1831), .B(n1830), .Z(n1988) );
  XOR U2287 ( .A(n1989), .B(n1988), .Z(n1990) );
  XOR U2288 ( .A(n1991), .B(n1990), .Z(n1995) );
  XOR U2289 ( .A(n1994), .B(n1995), .Z(n1997) );
  AND U2290 ( .A(o[7]), .B(\stack[1][16] ), .Z(n1996) );
  XOR U2291 ( .A(n1997), .B(n1996), .Z(n2003) );
  AND U2292 ( .A(o[8]), .B(\stack[1][15] ), .Z(n2001) );
  NAND U2293 ( .A(n1833), .B(n1832), .Z(n1837) );
  NAND U2294 ( .A(n1835), .B(n1834), .Z(n1836) );
  NAND U2295 ( .A(n1837), .B(n1836), .Z(n2000) );
  XOR U2296 ( .A(n2001), .B(n2000), .Z(n2002) );
  XNOR U2297 ( .A(n2003), .B(n2002), .Z(n1955) );
  NAND U2298 ( .A(o[9]), .B(\stack[1][14] ), .Z(n1956) );
  XNOR U2299 ( .A(n1957), .B(n1956), .Z(n1951) );
  AND U2300 ( .A(o[10]), .B(\stack[1][13] ), .Z(n1949) );
  AND U2301 ( .A(o[8]), .B(\stack[1][13] ), .Z(n1881) );
  XOR U2302 ( .A(n1841), .B(n1840), .Z(n1875) );
  XOR U2303 ( .A(n1843), .B(n1842), .Z(n1871) );
  XOR U2304 ( .A(n1845), .B(n1844), .Z(n1866) );
  AND U2305 ( .A(o[4]), .B(\stack[1][13] ), .Z(n1860) );
  AND U2306 ( .A(o[0]), .B(\stack[1][13] ), .Z(n1846) );
  AND U2307 ( .A(o[1]), .B(\stack[1][14] ), .Z(n1851) );
  AND U2308 ( .A(n1846), .B(n1851), .Z(n1847) );
  NAND U2309 ( .A(o[2]), .B(n1847), .Z(n1853) );
  NAND U2310 ( .A(n1851), .B(o[0]), .Z(n1848) );
  XNOR U2311 ( .A(o[2]), .B(n1848), .Z(n1849) );
  AND U2312 ( .A(\stack[1][13] ), .B(n1849), .Z(n1906) );
  NAND U2313 ( .A(\stack[1][15] ), .B(o[0]), .Z(n1850) );
  XNOR U2314 ( .A(n1851), .B(n1850), .Z(n1907) );
  NAND U2315 ( .A(n1906), .B(n1907), .Z(n1852) );
  NAND U2316 ( .A(n1853), .B(n1852), .Z(n1856) );
  XOR U2317 ( .A(n1855), .B(n1854), .Z(n1857) );
  NAND U2318 ( .A(n1856), .B(n1857), .Z(n1859) );
  AND U2319 ( .A(o[3]), .B(\stack[1][13] ), .Z(n1913) );
  NAND U2320 ( .A(n1913), .B(n1912), .Z(n1858) );
  NAND U2321 ( .A(n1859), .B(n1858), .Z(n1861) );
  NAND U2322 ( .A(n1860), .B(n1861), .Z(n1865) );
  XOR U2323 ( .A(n1861), .B(n1860), .Z(n1895) );
  XOR U2324 ( .A(n1863), .B(n1862), .Z(n1894) );
  NAND U2325 ( .A(n1895), .B(n1894), .Z(n1864) );
  NAND U2326 ( .A(n1865), .B(n1864), .Z(n1867) );
  NAND U2327 ( .A(n1866), .B(n1867), .Z(n1869) );
  XOR U2328 ( .A(n1867), .B(n1866), .Z(n1893) );
  AND U2329 ( .A(o[5]), .B(\stack[1][13] ), .Z(n1892) );
  NAND U2330 ( .A(n1893), .B(n1892), .Z(n1868) );
  NAND U2331 ( .A(n1869), .B(n1868), .Z(n1870) );
  NAND U2332 ( .A(n1871), .B(n1870), .Z(n1873) );
  AND U2333 ( .A(o[6]), .B(\stack[1][13] ), .Z(n1891) );
  XOR U2334 ( .A(n1871), .B(n1870), .Z(n1890) );
  NAND U2335 ( .A(n1891), .B(n1890), .Z(n1872) );
  NAND U2336 ( .A(n1873), .B(n1872), .Z(n1874) );
  NAND U2337 ( .A(n1875), .B(n1874), .Z(n1877) );
  XOR U2338 ( .A(n1875), .B(n1874), .Z(n1931) );
  AND U2339 ( .A(o[7]), .B(\stack[1][13] ), .Z(n1930) );
  NAND U2340 ( .A(n1931), .B(n1930), .Z(n1876) );
  NAND U2341 ( .A(n1877), .B(n1876), .Z(n1880) );
  NAND U2342 ( .A(n1881), .B(n1880), .Z(n1883) );
  XOR U2343 ( .A(n1881), .B(n1880), .Z(n1888) );
  NAND U2344 ( .A(n1889), .B(n1888), .Z(n1882) );
  NAND U2345 ( .A(n1883), .B(n1882), .Z(n1884) );
  NAND U2346 ( .A(n1885), .B(n1884), .Z(n1887) );
  XOR U2347 ( .A(n1885), .B(n1884), .Z(n1941) );
  AND U2348 ( .A(o[9]), .B(\stack[1][13] ), .Z(n1940) );
  NAND U2349 ( .A(n1941), .B(n1940), .Z(n1886) );
  NAND U2350 ( .A(n1887), .B(n1886), .Z(n1948) );
  XOR U2351 ( .A(n1949), .B(n1948), .Z(n1950) );
  XNOR U2352 ( .A(n1889), .B(n1888), .Z(n1934) );
  AND U2353 ( .A(o[8]), .B(\stack[1][12] ), .Z(n1928) );
  XOR U2354 ( .A(n1891), .B(n1890), .Z(n1924) );
  XOR U2355 ( .A(n1893), .B(n1892), .Z(n1921) );
  XOR U2356 ( .A(n1895), .B(n1894), .Z(n1897) );
  AND U2357 ( .A(o[5]), .B(\stack[1][12] ), .Z(n1896) );
  NAND U2358 ( .A(n1897), .B(n1896), .Z(n1919) );
  XOR U2359 ( .A(n1897), .B(n1896), .Z(n2081) );
  AND U2360 ( .A(o[0]), .B(\stack[1][12] ), .Z(n1898) );
  AND U2361 ( .A(o[1]), .B(\stack[1][13] ), .Z(n1903) );
  AND U2362 ( .A(n1898), .B(n1903), .Z(n1899) );
  NAND U2363 ( .A(o[2]), .B(n1899), .Z(n1905) );
  NAND U2364 ( .A(n1903), .B(o[0]), .Z(n1900) );
  XNOR U2365 ( .A(o[2]), .B(n1900), .Z(n1901) );
  AND U2366 ( .A(\stack[1][12] ), .B(n1901), .Z(n2090) );
  NAND U2367 ( .A(\stack[1][14] ), .B(o[0]), .Z(n1902) );
  XNOR U2368 ( .A(n1903), .B(n1902), .Z(n2091) );
  NAND U2369 ( .A(n2090), .B(n2091), .Z(n1904) );
  NAND U2370 ( .A(n1905), .B(n1904), .Z(n1908) );
  NAND U2371 ( .A(n1908), .B(n1909), .Z(n1911) );
  AND U2372 ( .A(o[3]), .B(\stack[1][12] ), .Z(n2098) );
  NAND U2373 ( .A(n2098), .B(n2099), .Z(n1910) );
  NAND U2374 ( .A(n1911), .B(n1910), .Z(n1914) );
  AND U2375 ( .A(o[4]), .B(\stack[1][12] ), .Z(n1915) );
  NAND U2376 ( .A(n1914), .B(n1915), .Z(n1917) );
  XOR U2377 ( .A(n1913), .B(n1912), .Z(n2103) );
  NAND U2378 ( .A(n2103), .B(n2102), .Z(n1916) );
  NAND U2379 ( .A(n1917), .B(n1916), .Z(n2080) );
  NAND U2380 ( .A(n2081), .B(n2080), .Z(n1918) );
  NAND U2381 ( .A(n1919), .B(n1918), .Z(n1920) );
  NAND U2382 ( .A(n1921), .B(n1920), .Z(n1923) );
  AND U2383 ( .A(o[6]), .B(\stack[1][12] ), .Z(n2079) );
  XOR U2384 ( .A(n1921), .B(n1920), .Z(n2078) );
  NAND U2385 ( .A(n2079), .B(n2078), .Z(n1922) );
  NAND U2386 ( .A(n1923), .B(n1922), .Z(n1925) );
  NAND U2387 ( .A(n1924), .B(n1925), .Z(n1927) );
  XOR U2388 ( .A(n1925), .B(n1924), .Z(n2117) );
  AND U2389 ( .A(o[7]), .B(\stack[1][12] ), .Z(n2116) );
  NAND U2390 ( .A(n2117), .B(n2116), .Z(n1926) );
  NAND U2391 ( .A(n1927), .B(n1926), .Z(n1929) );
  NAND U2392 ( .A(n1928), .B(n1929), .Z(n1933) );
  XOR U2393 ( .A(n1929), .B(n1928), .Z(n2077) );
  XOR U2394 ( .A(n1931), .B(n1930), .Z(n2076) );
  NAND U2395 ( .A(n2077), .B(n2076), .Z(n1932) );
  AND U2396 ( .A(n1933), .B(n1932), .Z(n1935) );
  NAND U2397 ( .A(n1934), .B(n1935), .Z(n1937) );
  NAND U2398 ( .A(o[9]), .B(\stack[1][12] ), .Z(n2126) );
  NAND U2399 ( .A(n2127), .B(n2126), .Z(n1936) );
  NAND U2400 ( .A(n1937), .B(n1936), .Z(n1939) );
  NAND U2401 ( .A(o[10]), .B(\stack[1][12] ), .Z(n1938) );
  NAND U2402 ( .A(n1939), .B(n1938), .Z(n1943) );
  XOR U2403 ( .A(n1939), .B(n1938), .Z(n2133) );
  XNOR U2404 ( .A(n1941), .B(n1940), .Z(n2132) );
  NAND U2405 ( .A(n2133), .B(n2132), .Z(n1942) );
  AND U2406 ( .A(n1943), .B(n1942), .Z(n1945) );
  NANDN U2407 ( .A(n1944), .B(n1945), .Z(n1947) );
  XNOR U2408 ( .A(n1945), .B(n1944), .Z(n2139) );
  AND U2409 ( .A(\stack[1][12] ), .B(o[11]), .Z(n2138) );
  NAND U2410 ( .A(n2139), .B(n2138), .Z(n1946) );
  NAND U2411 ( .A(n1947), .B(n1946), .Z(n2007) );
  NAND U2412 ( .A(n2006), .B(n2007), .Z(n2009) );
  NAND U2413 ( .A(n1949), .B(n1948), .Z(n1953) );
  NAND U2414 ( .A(n1951), .B(n1950), .Z(n1952) );
  AND U2415 ( .A(n1953), .B(n1952), .Z(n2069) );
  NAND U2416 ( .A(n1955), .B(n1954), .Z(n1959) );
  NAND U2417 ( .A(n1957), .B(n1956), .Z(n1958) );
  NAND U2418 ( .A(n1959), .B(n1958), .Z(n2011) );
  NAND U2419 ( .A(o[10]), .B(\stack[1][14] ), .Z(n2010) );
  XOR U2420 ( .A(n2011), .B(n2010), .Z(n2013) );
  AND U2421 ( .A(o[6]), .B(\stack[1][18] ), .Z(n2025) );
  NAND U2422 ( .A(n1961), .B(n1960), .Z(n1965) );
  NAND U2423 ( .A(n1963), .B(n1962), .Z(n1964) );
  NAND U2424 ( .A(n1965), .B(n1964), .Z(n2050) );
  AND U2425 ( .A(o[3]), .B(\stack[1][21] ), .Z(n2030) );
  AND U2426 ( .A(o[0]), .B(\stack[1][21] ), .Z(n1967) );
  AND U2427 ( .A(n1967), .B(n1966), .Z(n1968) );
  NAND U2428 ( .A(o[2]), .B(n1968), .Z(n1972) );
  NAND U2429 ( .A(n1970), .B(n1969), .Z(n1971) );
  NAND U2430 ( .A(n1972), .B(n1971), .Z(n2028) );
  AND U2431 ( .A(o[1]), .B(\stack[1][23] ), .Z(n2037) );
  NAND U2432 ( .A(\stack[1][24] ), .B(o[0]), .Z(n1973) );
  XNOR U2433 ( .A(n2037), .B(n1973), .Z(n2041) );
  NAND U2434 ( .A(n2037), .B(o[0]), .Z(n1974) );
  XNOR U2435 ( .A(o[2]), .B(n1974), .Z(n1975) );
  AND U2436 ( .A(\stack[1][22] ), .B(n1975), .Z(n2040) );
  XOR U2437 ( .A(n2041), .B(n2040), .Z(n2029) );
  XOR U2438 ( .A(n2028), .B(n2029), .Z(n2031) );
  AND U2439 ( .A(o[4]), .B(\stack[1][20] ), .Z(n2045) );
  NAND U2440 ( .A(n1977), .B(n1976), .Z(n1981) );
  NAND U2441 ( .A(n1979), .B(n1978), .Z(n1980) );
  NAND U2442 ( .A(n1981), .B(n1980), .Z(n2044) );
  XOR U2443 ( .A(n2045), .B(n2044), .Z(n2046) );
  XOR U2444 ( .A(n2047), .B(n2046), .Z(n2051) );
  XOR U2445 ( .A(n2050), .B(n2051), .Z(n2053) );
  AND U2446 ( .A(o[5]), .B(\stack[1][19] ), .Z(n2052) );
  XOR U2447 ( .A(n2053), .B(n2052), .Z(n2023) );
  NAND U2448 ( .A(n1983), .B(n1982), .Z(n1987) );
  NAND U2449 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U2450 ( .A(n1987), .B(n1986), .Z(n2022) );
  XOR U2451 ( .A(n2023), .B(n2022), .Z(n2024) );
  XOR U2452 ( .A(n2025), .B(n2024), .Z(n2057) );
  NAND U2453 ( .A(n1989), .B(n1988), .Z(n1993) );
  NAND U2454 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U2455 ( .A(n1993), .B(n1992), .Z(n2056) );
  XOR U2456 ( .A(n2057), .B(n2056), .Z(n2059) );
  AND U2457 ( .A(o[7]), .B(\stack[1][17] ), .Z(n2058) );
  XOR U2458 ( .A(n2059), .B(n2058), .Z(n2018) );
  NAND U2459 ( .A(n1995), .B(n1994), .Z(n1999) );
  NAND U2460 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U2461 ( .A(n1999), .B(n1998), .Z(n2016) );
  AND U2462 ( .A(o[8]), .B(\stack[1][16] ), .Z(n2017) );
  XOR U2463 ( .A(n2016), .B(n2017), .Z(n2019) );
  NAND U2464 ( .A(n2001), .B(n2000), .Z(n2005) );
  NAND U2465 ( .A(n2003), .B(n2002), .Z(n2004) );
  NAND U2466 ( .A(n2005), .B(n2004), .Z(n2062) );
  XOR U2467 ( .A(n2063), .B(n2062), .Z(n2065) );
  AND U2468 ( .A(o[9]), .B(\stack[1][15] ), .Z(n2064) );
  XNOR U2469 ( .A(n2065), .B(n2064), .Z(n2012) );
  XOR U2470 ( .A(n2013), .B(n2012), .Z(n2068) );
  XOR U2471 ( .A(n2069), .B(n2068), .Z(n2071) );
  NAND U2472 ( .A(\stack[1][13] ), .B(o[11]), .Z(n2070) );
  XNOR U2473 ( .A(n2071), .B(n2070), .Z(n2074) );
  XOR U2474 ( .A(n2007), .B(n2006), .Z(n2075) );
  NAND U2475 ( .A(n2074), .B(n2075), .Z(n2008) );
  AND U2476 ( .A(n2009), .B(n2008), .Z(n2240) );
  NAND U2477 ( .A(n2011), .B(n2010), .Z(n2015) );
  NAND U2478 ( .A(n2013), .B(n2012), .Z(n2014) );
  AND U2479 ( .A(n2015), .B(n2014), .Z(n2246) );
  NAND U2480 ( .A(n2017), .B(n2016), .Z(n2021) );
  NAND U2481 ( .A(n2019), .B(n2018), .Z(n2020) );
  AND U2482 ( .A(n2021), .B(n2020), .Z(n2298) );
  AND U2483 ( .A(o[7]), .B(\stack[1][18] ), .Z(n2254) );
  NAND U2484 ( .A(n2023), .B(n2022), .Z(n2027) );
  NAND U2485 ( .A(n2025), .B(n2024), .Z(n2026) );
  NAND U2486 ( .A(n2027), .B(n2026), .Z(n2252) );
  AND U2487 ( .A(o[6]), .B(\stack[1][19] ), .Z(n2289) );
  NAND U2488 ( .A(n2029), .B(n2028), .Z(n2033) );
  NAND U2489 ( .A(n2031), .B(n2030), .Z(n2032) );
  NAND U2490 ( .A(n2033), .B(n2032), .Z(n2258) );
  AND U2491 ( .A(o[4]), .B(\stack[1][21] ), .Z(n2259) );
  XOR U2492 ( .A(n2258), .B(n2259), .Z(n2261) );
  AND U2493 ( .A(o[1]), .B(\stack[1][24] ), .Z(n2264) );
  NAND U2494 ( .A(\stack[1][25] ), .B(o[0]), .Z(n2034) );
  XNOR U2495 ( .A(n2264), .B(n2034), .Z(n2268) );
  NAND U2496 ( .A(n2264), .B(o[0]), .Z(n2035) );
  XNOR U2497 ( .A(o[2]), .B(n2035), .Z(n2036) );
  AND U2498 ( .A(\stack[1][23] ), .B(n2036), .Z(n2267) );
  XOR U2499 ( .A(n2268), .B(n2267), .Z(n2275) );
  AND U2500 ( .A(o[0]), .B(\stack[1][22] ), .Z(n2038) );
  AND U2501 ( .A(n2038), .B(n2037), .Z(n2039) );
  NAND U2502 ( .A(o[2]), .B(n2039), .Z(n2043) );
  NAND U2503 ( .A(n2041), .B(n2040), .Z(n2042) );
  NAND U2504 ( .A(n2043), .B(n2042), .Z(n2274) );
  XOR U2505 ( .A(n2275), .B(n2274), .Z(n2277) );
  AND U2506 ( .A(o[3]), .B(\stack[1][22] ), .Z(n2276) );
  XOR U2507 ( .A(n2277), .B(n2276), .Z(n2260) );
  XOR U2508 ( .A(n2261), .B(n2260), .Z(n2281) );
  AND U2509 ( .A(o[5]), .B(\stack[1][20] ), .Z(n2280) );
  XOR U2510 ( .A(n2281), .B(n2280), .Z(n2283) );
  NAND U2511 ( .A(n2045), .B(n2044), .Z(n2049) );
  NAND U2512 ( .A(n2047), .B(n2046), .Z(n2048) );
  NAND U2513 ( .A(n2049), .B(n2048), .Z(n2282) );
  XOR U2514 ( .A(n2283), .B(n2282), .Z(n2287) );
  NAND U2515 ( .A(n2051), .B(n2050), .Z(n2055) );
  NAND U2516 ( .A(n2053), .B(n2052), .Z(n2054) );
  NAND U2517 ( .A(n2055), .B(n2054), .Z(n2286) );
  XOR U2518 ( .A(n2287), .B(n2286), .Z(n2288) );
  XOR U2519 ( .A(n2289), .B(n2288), .Z(n2253) );
  XOR U2520 ( .A(n2252), .B(n2253), .Z(n2255) );
  AND U2521 ( .A(o[8]), .B(\stack[1][17] ), .Z(n2293) );
  NAND U2522 ( .A(n2057), .B(n2056), .Z(n2061) );
  NAND U2523 ( .A(n2059), .B(n2058), .Z(n2060) );
  NAND U2524 ( .A(n2061), .B(n2060), .Z(n2292) );
  XOR U2525 ( .A(n2293), .B(n2292), .Z(n2294) );
  XNOR U2526 ( .A(n2295), .B(n2294), .Z(n2299) );
  NAND U2527 ( .A(o[9]), .B(\stack[1][16] ), .Z(n2300) );
  XNOR U2528 ( .A(n2301), .B(n2300), .Z(n2307) );
  AND U2529 ( .A(o[10]), .B(\stack[1][15] ), .Z(n2305) );
  NAND U2530 ( .A(n2063), .B(n2062), .Z(n2067) );
  NAND U2531 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U2532 ( .A(n2067), .B(n2066), .Z(n2304) );
  XOR U2533 ( .A(n2305), .B(n2304), .Z(n2306) );
  XNOR U2534 ( .A(n2246), .B(n2247), .Z(n2249) );
  AND U2535 ( .A(o[11]), .B(\stack[1][14] ), .Z(n2248) );
  XOR U2536 ( .A(n2249), .B(n2248), .Z(n2313) );
  AND U2537 ( .A(\stack[1][13] ), .B(o[12]), .Z(n2311) );
  NAND U2538 ( .A(n2069), .B(n2068), .Z(n2073) );
  NAND U2539 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2540 ( .A(n2073), .B(n2072), .Z(n2310) );
  XOR U2541 ( .A(n2311), .B(n2310), .Z(n2312) );
  XNOR U2542 ( .A(n2313), .B(n2312), .Z(n2241) );
  NAND U2543 ( .A(\stack[1][12] ), .B(o[13]), .Z(n2242) );
  XNOR U2544 ( .A(n2243), .B(n2242), .Z(n2237) );
  AND U2545 ( .A(\stack[1][11] ), .B(o[14]), .Z(n2235) );
  AND U2546 ( .A(\stack[1][11] ), .B(o[12]), .Z(n2141) );
  AND U2547 ( .A(o[10]), .B(\stack[1][11] ), .Z(n2129) );
  XOR U2548 ( .A(n2077), .B(n2076), .Z(n2123) );
  AND U2549 ( .A(o[8]), .B(\stack[1][11] ), .Z(n2119) );
  XOR U2550 ( .A(n2079), .B(n2078), .Z(n2113) );
  XOR U2551 ( .A(n2081), .B(n2080), .Z(n2109) );
  AND U2552 ( .A(o[0]), .B(\stack[1][11] ), .Z(n2082) );
  AND U2553 ( .A(o[1]), .B(\stack[1][12] ), .Z(n2087) );
  AND U2554 ( .A(n2082), .B(n2087), .Z(n2083) );
  NAND U2555 ( .A(o[2]), .B(n2083), .Z(n2089) );
  NAND U2556 ( .A(n2087), .B(o[0]), .Z(n2084) );
  XNOR U2557 ( .A(o[2]), .B(n2084), .Z(n2085) );
  AND U2558 ( .A(\stack[1][11] ), .B(n2085), .Z(n2164) );
  NAND U2559 ( .A(\stack[1][13] ), .B(o[0]), .Z(n2086) );
  XNOR U2560 ( .A(n2087), .B(n2086), .Z(n2165) );
  NAND U2561 ( .A(n2164), .B(n2165), .Z(n2088) );
  NAND U2562 ( .A(n2089), .B(n2088), .Z(n2092) );
  NAND U2563 ( .A(n2092), .B(n2093), .Z(n2095) );
  AND U2564 ( .A(o[3]), .B(\stack[1][11] ), .Z(n2171) );
  NAND U2565 ( .A(n2171), .B(n2170), .Z(n2094) );
  NAND U2566 ( .A(n2095), .B(n2094), .Z(n2096) );
  AND U2567 ( .A(o[4]), .B(\stack[1][11] ), .Z(n2097) );
  NAND U2568 ( .A(n2096), .B(n2097), .Z(n2101) );
  NAND U2569 ( .A(n2155), .B(n2154), .Z(n2100) );
  NAND U2570 ( .A(n2101), .B(n2100), .Z(n2104) );
  XOR U2571 ( .A(n2103), .B(n2102), .Z(n2105) );
  NAND U2572 ( .A(n2104), .B(n2105), .Z(n2107) );
  AND U2573 ( .A(o[5]), .B(\stack[1][11] ), .Z(n2180) );
  NAND U2574 ( .A(n2180), .B(n2181), .Z(n2106) );
  NAND U2575 ( .A(n2107), .B(n2106), .Z(n2108) );
  NAND U2576 ( .A(n2109), .B(n2108), .Z(n2111) );
  AND U2577 ( .A(o[6]), .B(\stack[1][11] ), .Z(n2187) );
  XOR U2578 ( .A(n2109), .B(n2108), .Z(n2186) );
  NAND U2579 ( .A(n2187), .B(n2186), .Z(n2110) );
  NAND U2580 ( .A(n2111), .B(n2110), .Z(n2112) );
  NAND U2581 ( .A(n2113), .B(n2112), .Z(n2115) );
  XOR U2582 ( .A(n2113), .B(n2112), .Z(n2195) );
  AND U2583 ( .A(o[7]), .B(\stack[1][11] ), .Z(n2194) );
  NAND U2584 ( .A(n2195), .B(n2194), .Z(n2114) );
  NAND U2585 ( .A(n2115), .B(n2114), .Z(n2118) );
  NAND U2586 ( .A(n2119), .B(n2118), .Z(n2121) );
  XOR U2587 ( .A(n2117), .B(n2116), .Z(n2153) );
  XOR U2588 ( .A(n2119), .B(n2118), .Z(n2152) );
  NAND U2589 ( .A(n2153), .B(n2152), .Z(n2120) );
  NAND U2590 ( .A(n2121), .B(n2120), .Z(n2122) );
  NAND U2591 ( .A(n2123), .B(n2122), .Z(n2125) );
  XOR U2592 ( .A(n2123), .B(n2122), .Z(n2205) );
  AND U2593 ( .A(\stack[1][11] ), .B(o[9]), .Z(n2204) );
  NAND U2594 ( .A(n2205), .B(n2204), .Z(n2124) );
  NAND U2595 ( .A(n2125), .B(n2124), .Z(n2128) );
  NAND U2596 ( .A(n2129), .B(n2128), .Z(n2131) );
  XNOR U2597 ( .A(n2127), .B(n2126), .Z(n2150) );
  XOR U2598 ( .A(n2129), .B(n2128), .Z(n2151) );
  NAND U2599 ( .A(n2150), .B(n2151), .Z(n2130) );
  AND U2600 ( .A(n2131), .B(n2130), .Z(n2135) );
  XOR U2601 ( .A(n2133), .B(n2132), .Z(n2134) );
  NAND U2602 ( .A(n2135), .B(n2134), .Z(n2137) );
  XOR U2603 ( .A(n2135), .B(n2134), .Z(n2212) );
  NAND U2604 ( .A(\stack[1][11] ), .B(o[11]), .Z(n2213) );
  NAND U2605 ( .A(n2212), .B(n2213), .Z(n2136) );
  AND U2606 ( .A(n2137), .B(n2136), .Z(n2140) );
  NAND U2607 ( .A(n2141), .B(n2140), .Z(n2143) );
  XOR U2608 ( .A(n2139), .B(n2138), .Z(n2149) );
  XOR U2609 ( .A(n2141), .B(n2140), .Z(n2148) );
  NAND U2610 ( .A(n2149), .B(n2148), .Z(n2142) );
  NAND U2611 ( .A(n2143), .B(n2142), .Z(n2144) );
  NAND U2612 ( .A(n2145), .B(n2144), .Z(n2147) );
  XOR U2613 ( .A(n2145), .B(n2144), .Z(n2225) );
  AND U2614 ( .A(\stack[1][11] ), .B(o[13]), .Z(n2224) );
  NAND U2615 ( .A(n2225), .B(n2224), .Z(n2146) );
  NAND U2616 ( .A(n2147), .B(n2146), .Z(n2234) );
  XOR U2617 ( .A(n2235), .B(n2234), .Z(n2236) );
  AND U2618 ( .A(\stack[1][10] ), .B(o[14]), .Z(n2222) );
  XOR U2619 ( .A(n2149), .B(n2148), .Z(n2218) );
  AND U2620 ( .A(\stack[1][10] ), .B(o[12]), .Z(n2214) );
  AND U2621 ( .A(o[10]), .B(\stack[1][10] ), .Z(n2203) );
  XNOR U2622 ( .A(n2153), .B(n2152), .Z(n2198) );
  AND U2623 ( .A(o[5]), .B(\stack[1][10] ), .Z(n2176) );
  XOR U2624 ( .A(n2155), .B(n2154), .Z(n2177) );
  NAND U2625 ( .A(n2176), .B(n2177), .Z(n2179) );
  AND U2626 ( .A(o[0]), .B(\stack[1][10] ), .Z(n2156) );
  AND U2627 ( .A(o[1]), .B(\stack[1][11] ), .Z(n2161) );
  AND U2628 ( .A(n2156), .B(n2161), .Z(n2157) );
  NAND U2629 ( .A(o[2]), .B(n2157), .Z(n2163) );
  NAND U2630 ( .A(n2161), .B(o[0]), .Z(n2158) );
  XNOR U2631 ( .A(o[2]), .B(n2158), .Z(n2159) );
  AND U2632 ( .A(\stack[1][10] ), .B(n2159), .Z(n2420) );
  NAND U2633 ( .A(\stack[1][12] ), .B(o[0]), .Z(n2160) );
  XNOR U2634 ( .A(n2161), .B(n2160), .Z(n2421) );
  NAND U2635 ( .A(n2420), .B(n2421), .Z(n2162) );
  NAND U2636 ( .A(n2163), .B(n2162), .Z(n2166) );
  NAND U2637 ( .A(n2166), .B(n2167), .Z(n2169) );
  AND U2638 ( .A(o[3]), .B(\stack[1][10] ), .Z(n2428) );
  NAND U2639 ( .A(n2428), .B(n2429), .Z(n2168) );
  NAND U2640 ( .A(n2169), .B(n2168), .Z(n2172) );
  AND U2641 ( .A(o[4]), .B(\stack[1][10] ), .Z(n2173) );
  NAND U2642 ( .A(n2172), .B(n2173), .Z(n2175) );
  XOR U2643 ( .A(n2171), .B(n2170), .Z(n2433) );
  NAND U2644 ( .A(n2433), .B(n2432), .Z(n2174) );
  NAND U2645 ( .A(n2175), .B(n2174), .Z(n2439) );
  NAND U2646 ( .A(n2439), .B(n2440), .Z(n2178) );
  NAND U2647 ( .A(n2179), .B(n2178), .Z(n2182) );
  NAND U2648 ( .A(n2182), .B(n2183), .Z(n2185) );
  AND U2649 ( .A(o[6]), .B(\stack[1][10] ), .Z(n2445) );
  NAND U2650 ( .A(n2445), .B(n2446), .Z(n2184) );
  NAND U2651 ( .A(n2185), .B(n2184), .Z(n2188) );
  XOR U2652 ( .A(n2187), .B(n2186), .Z(n2189) );
  NAND U2653 ( .A(n2188), .B(n2189), .Z(n2191) );
  AND U2654 ( .A(o[7]), .B(\stack[1][10] ), .Z(n2452) );
  NAND U2655 ( .A(n2452), .B(n2451), .Z(n2190) );
  NAND U2656 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U2657 ( .A(o[8]), .B(\stack[1][10] ), .Z(n2193) );
  NAND U2658 ( .A(n2192), .B(n2193), .Z(n2197) );
  XOR U2659 ( .A(n2195), .B(n2194), .Z(n2457) );
  NAND U2660 ( .A(n2458), .B(n2457), .Z(n2196) );
  AND U2661 ( .A(n2197), .B(n2196), .Z(n2199) );
  NAND U2662 ( .A(n2198), .B(n2199), .Z(n2201) );
  NAND U2663 ( .A(\stack[1][10] ), .B(o[9]), .Z(n2463) );
  NAND U2664 ( .A(n2464), .B(n2463), .Z(n2200) );
  AND U2665 ( .A(n2201), .B(n2200), .Z(n2202) );
  NAND U2666 ( .A(n2203), .B(n2202), .Z(n2207) );
  XOR U2667 ( .A(n2203), .B(n2202), .Z(n2411) );
  XOR U2668 ( .A(n2205), .B(n2204), .Z(n2410) );
  NAND U2669 ( .A(n2411), .B(n2410), .Z(n2206) );
  NAND U2670 ( .A(n2207), .B(n2206), .Z(n2209) );
  NANDN U2671 ( .A(n2208), .B(n2209), .Z(n2211) );
  XOR U2672 ( .A(n2209), .B(n2208), .Z(n2473) );
  AND U2673 ( .A(\stack[1][10] ), .B(o[11]), .Z(n2474) );
  NANDN U2674 ( .A(n2473), .B(n2474), .Z(n2210) );
  NAND U2675 ( .A(n2211), .B(n2210), .Z(n2215) );
  NAND U2676 ( .A(n2214), .B(n2215), .Z(n2217) );
  XNOR U2677 ( .A(n2213), .B(n2212), .Z(n2408) );
  XOR U2678 ( .A(n2215), .B(n2214), .Z(n2409) );
  NAND U2679 ( .A(n2408), .B(n2409), .Z(n2216) );
  NAND U2680 ( .A(n2217), .B(n2216), .Z(n2219) );
  NAND U2681 ( .A(n2218), .B(n2219), .Z(n2221) );
  XOR U2682 ( .A(n2219), .B(n2218), .Z(n2484) );
  AND U2683 ( .A(\stack[1][10] ), .B(o[13]), .Z(n2483) );
  NAND U2684 ( .A(n2484), .B(n2483), .Z(n2220) );
  NAND U2685 ( .A(n2221), .B(n2220), .Z(n2223) );
  NAND U2686 ( .A(n2222), .B(n2223), .Z(n2227) );
  XOR U2687 ( .A(n2223), .B(n2222), .Z(n2407) );
  XOR U2688 ( .A(n2225), .B(n2224), .Z(n2406) );
  NAND U2689 ( .A(n2407), .B(n2406), .Z(n2226) );
  NAND U2690 ( .A(n2227), .B(n2226), .Z(n2229) );
  NAND U2691 ( .A(n2228), .B(n2229), .Z(n2231) );
  XOR U2692 ( .A(n2229), .B(n2228), .Z(n2494) );
  AND U2693 ( .A(\stack[1][10] ), .B(o[15]), .Z(n2493) );
  NAND U2694 ( .A(n2494), .B(n2493), .Z(n2230) );
  AND U2695 ( .A(n2231), .B(n2230), .Z(n2233) );
  NAND U2696 ( .A(\stack[1][10] ), .B(o[16]), .Z(n2232) );
  NAND U2697 ( .A(n2233), .B(n2232), .Z(n2317) );
  XOR U2698 ( .A(n2233), .B(n2232), .Z(n2500) );
  NAND U2699 ( .A(n2235), .B(n2234), .Z(n2239) );
  NAND U2700 ( .A(n2237), .B(n2236), .Z(n2238) );
  NAND U2701 ( .A(n2239), .B(n2238), .Z(n2401) );
  NAND U2702 ( .A(n2241), .B(n2240), .Z(n2245) );
  NAND U2703 ( .A(n2243), .B(n2242), .Z(n2244) );
  NAND U2704 ( .A(n2245), .B(n2244), .Z(n2319) );
  NAND U2705 ( .A(\stack[1][12] ), .B(o[14]), .Z(n2318) );
  XOR U2706 ( .A(n2319), .B(n2318), .Z(n2321) );
  NANDN U2707 ( .A(n2247), .B(n2246), .Z(n2251) );
  NAND U2708 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2709 ( .A(n2251), .B(n2250), .Z(n2324) );
  AND U2710 ( .A(o[12]), .B(\stack[1][14] ), .Z(n2325) );
  XOR U2711 ( .A(n2324), .B(n2325), .Z(n2326) );
  NAND U2712 ( .A(n2253), .B(n2252), .Z(n2257) );
  NAND U2713 ( .A(n2255), .B(n2254), .Z(n2256) );
  NAND U2714 ( .A(n2257), .B(n2256), .Z(n2336) );
  AND U2715 ( .A(o[8]), .B(\stack[1][18] ), .Z(n2337) );
  XOR U2716 ( .A(n2336), .B(n2337), .Z(n2339) );
  AND U2717 ( .A(o[6]), .B(\stack[1][20] ), .Z(n2345) );
  NAND U2718 ( .A(n2259), .B(n2258), .Z(n2263) );
  NAND U2719 ( .A(n2261), .B(n2260), .Z(n2262) );
  NAND U2720 ( .A(n2263), .B(n2262), .Z(n2370) );
  AND U2721 ( .A(o[3]), .B(\stack[1][23] ), .Z(n2350) );
  AND U2722 ( .A(o[0]), .B(\stack[1][23] ), .Z(n2265) );
  AND U2723 ( .A(n2265), .B(n2264), .Z(n2266) );
  NAND U2724 ( .A(o[2]), .B(n2266), .Z(n2270) );
  NAND U2725 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U2726 ( .A(n2270), .B(n2269), .Z(n2348) );
  AND U2727 ( .A(o[1]), .B(\stack[1][25] ), .Z(n2357) );
  NAND U2728 ( .A(\stack[1][26] ), .B(o[0]), .Z(n2271) );
  XNOR U2729 ( .A(n2357), .B(n2271), .Z(n2361) );
  NAND U2730 ( .A(n2357), .B(o[0]), .Z(n2272) );
  XNOR U2731 ( .A(o[2]), .B(n2272), .Z(n2273) );
  AND U2732 ( .A(\stack[1][24] ), .B(n2273), .Z(n2360) );
  XOR U2733 ( .A(n2361), .B(n2360), .Z(n2349) );
  XOR U2734 ( .A(n2348), .B(n2349), .Z(n2351) );
  AND U2735 ( .A(o[4]), .B(\stack[1][22] ), .Z(n2365) );
  NAND U2736 ( .A(n2275), .B(n2274), .Z(n2279) );
  NAND U2737 ( .A(n2277), .B(n2276), .Z(n2278) );
  NAND U2738 ( .A(n2279), .B(n2278), .Z(n2364) );
  XOR U2739 ( .A(n2365), .B(n2364), .Z(n2366) );
  XOR U2740 ( .A(n2367), .B(n2366), .Z(n2371) );
  XOR U2741 ( .A(n2370), .B(n2371), .Z(n2373) );
  AND U2742 ( .A(o[5]), .B(\stack[1][21] ), .Z(n2372) );
  XOR U2743 ( .A(n2373), .B(n2372), .Z(n2343) );
  NAND U2744 ( .A(n2281), .B(n2280), .Z(n2285) );
  NAND U2745 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U2746 ( .A(n2285), .B(n2284), .Z(n2342) );
  XOR U2747 ( .A(n2343), .B(n2342), .Z(n2344) );
  XOR U2748 ( .A(n2345), .B(n2344), .Z(n2377) );
  NAND U2749 ( .A(n2287), .B(n2286), .Z(n2291) );
  NAND U2750 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2751 ( .A(n2291), .B(n2290), .Z(n2376) );
  XOR U2752 ( .A(n2377), .B(n2376), .Z(n2379) );
  AND U2753 ( .A(o[7]), .B(\stack[1][19] ), .Z(n2378) );
  XOR U2754 ( .A(n2379), .B(n2378), .Z(n2338) );
  XOR U2755 ( .A(n2339), .B(n2338), .Z(n2383) );
  NAND U2756 ( .A(n2293), .B(n2292), .Z(n2297) );
  NAND U2757 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2758 ( .A(n2297), .B(n2296), .Z(n2382) );
  XOR U2759 ( .A(n2383), .B(n2382), .Z(n2385) );
  AND U2760 ( .A(o[9]), .B(\stack[1][17] ), .Z(n2384) );
  XOR U2761 ( .A(n2385), .B(n2384), .Z(n2333) );
  NAND U2762 ( .A(n2299), .B(n2298), .Z(n2303) );
  NAND U2763 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2764 ( .A(n2303), .B(n2302), .Z(n2331) );
  AND U2765 ( .A(o[10]), .B(\stack[1][16] ), .Z(n2330) );
  XOR U2766 ( .A(n2331), .B(n2330), .Z(n2332) );
  XNOR U2767 ( .A(n2333), .B(n2332), .Z(n2389) );
  NAND U2768 ( .A(n2305), .B(n2304), .Z(n2309) );
  NAND U2769 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U2770 ( .A(n2309), .B(n2308), .Z(n2388) );
  NAND U2771 ( .A(o[11]), .B(\stack[1][15] ), .Z(n2390) );
  XNOR U2772 ( .A(n2391), .B(n2390), .Z(n2327) );
  NAND U2773 ( .A(n2311), .B(n2310), .Z(n2315) );
  NAND U2774 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2775 ( .A(n2315), .B(n2314), .Z(n2394) );
  XOR U2776 ( .A(n2395), .B(n2394), .Z(n2397) );
  AND U2777 ( .A(\stack[1][13] ), .B(o[13]), .Z(n2396) );
  XNOR U2778 ( .A(n2397), .B(n2396), .Z(n2320) );
  XNOR U2779 ( .A(n2321), .B(n2320), .Z(n2400) );
  XOR U2780 ( .A(n2401), .B(n2400), .Z(n2403) );
  AND U2781 ( .A(\stack[1][11] ), .B(o[15]), .Z(n2402) );
  XNOR U2782 ( .A(n2403), .B(n2402), .Z(n2499) );
  NAND U2783 ( .A(n2500), .B(n2499), .Z(n2316) );
  AND U2784 ( .A(n2317), .B(n2316), .Z(n2615) );
  AND U2785 ( .A(\stack[1][12] ), .B(o[15]), .Z(n2623) );
  NAND U2786 ( .A(n2319), .B(n2318), .Z(n2323) );
  NAND U2787 ( .A(n2321), .B(n2320), .Z(n2322) );
  AND U2788 ( .A(n2323), .B(n2322), .Z(n2621) );
  NAND U2789 ( .A(n2325), .B(n2324), .Z(n2329) );
  NAND U2790 ( .A(n2327), .B(n2326), .Z(n2328) );
  AND U2791 ( .A(n2329), .B(n2328), .Z(n2696) );
  NAND U2792 ( .A(n2331), .B(n2330), .Z(n2335) );
  NAND U2793 ( .A(n2333), .B(n2332), .Z(n2334) );
  NAND U2794 ( .A(n2335), .B(n2334), .Z(n2632) );
  NAND U2795 ( .A(n2337), .B(n2336), .Z(n2341) );
  NAND U2796 ( .A(n2339), .B(n2338), .Z(n2340) );
  AND U2797 ( .A(n2341), .B(n2340), .Z(n2684) );
  NAND U2798 ( .A(n2343), .B(n2342), .Z(n2347) );
  NAND U2799 ( .A(n2345), .B(n2344), .Z(n2346) );
  NAND U2800 ( .A(n2347), .B(n2346), .Z(n2672) );
  AND U2801 ( .A(o[6]), .B(\stack[1][21] ), .Z(n2669) );
  NAND U2802 ( .A(n2349), .B(n2348), .Z(n2353) );
  NAND U2803 ( .A(n2351), .B(n2350), .Z(n2352) );
  NAND U2804 ( .A(n2353), .B(n2352), .Z(n2638) );
  AND U2805 ( .A(o[4]), .B(\stack[1][23] ), .Z(n2639) );
  XOR U2806 ( .A(n2638), .B(n2639), .Z(n2641) );
  AND U2807 ( .A(o[1]), .B(\stack[1][26] ), .Z(n2644) );
  NAND U2808 ( .A(\stack[1][27] ), .B(o[0]), .Z(n2354) );
  XNOR U2809 ( .A(n2644), .B(n2354), .Z(n2648) );
  NAND U2810 ( .A(n2644), .B(o[0]), .Z(n2355) );
  XNOR U2811 ( .A(o[2]), .B(n2355), .Z(n2356) );
  AND U2812 ( .A(\stack[1][25] ), .B(n2356), .Z(n2647) );
  XOR U2813 ( .A(n2648), .B(n2647), .Z(n2655) );
  AND U2814 ( .A(o[0]), .B(\stack[1][24] ), .Z(n2358) );
  AND U2815 ( .A(n2358), .B(n2357), .Z(n2359) );
  NAND U2816 ( .A(o[2]), .B(n2359), .Z(n2363) );
  NAND U2817 ( .A(n2361), .B(n2360), .Z(n2362) );
  NAND U2818 ( .A(n2363), .B(n2362), .Z(n2654) );
  XOR U2819 ( .A(n2655), .B(n2654), .Z(n2657) );
  AND U2820 ( .A(o[3]), .B(\stack[1][24] ), .Z(n2656) );
  XOR U2821 ( .A(n2657), .B(n2656), .Z(n2640) );
  XOR U2822 ( .A(n2641), .B(n2640), .Z(n2661) );
  AND U2823 ( .A(o[5]), .B(\stack[1][22] ), .Z(n2660) );
  XOR U2824 ( .A(n2661), .B(n2660), .Z(n2663) );
  NAND U2825 ( .A(n2365), .B(n2364), .Z(n2369) );
  NAND U2826 ( .A(n2367), .B(n2366), .Z(n2368) );
  NAND U2827 ( .A(n2369), .B(n2368), .Z(n2662) );
  XOR U2828 ( .A(n2663), .B(n2662), .Z(n2667) );
  NAND U2829 ( .A(n2371), .B(n2370), .Z(n2375) );
  NAND U2830 ( .A(n2373), .B(n2372), .Z(n2374) );
  NAND U2831 ( .A(n2375), .B(n2374), .Z(n2666) );
  XOR U2832 ( .A(n2667), .B(n2666), .Z(n2668) );
  XOR U2833 ( .A(n2669), .B(n2668), .Z(n2673) );
  XOR U2834 ( .A(n2672), .B(n2673), .Z(n2675) );
  AND U2835 ( .A(o[7]), .B(\stack[1][20] ), .Z(n2674) );
  XOR U2836 ( .A(n2675), .B(n2674), .Z(n2681) );
  AND U2837 ( .A(o[8]), .B(\stack[1][19] ), .Z(n2679) );
  NAND U2838 ( .A(n2377), .B(n2376), .Z(n2381) );
  NAND U2839 ( .A(n2379), .B(n2378), .Z(n2380) );
  NAND U2840 ( .A(n2381), .B(n2380), .Z(n2678) );
  XOR U2841 ( .A(n2679), .B(n2678), .Z(n2680) );
  XNOR U2842 ( .A(n2681), .B(n2680), .Z(n2685) );
  NAND U2843 ( .A(o[9]), .B(\stack[1][18] ), .Z(n2686) );
  XNOR U2844 ( .A(n2687), .B(n2686), .Z(n2693) );
  AND U2845 ( .A(o[10]), .B(\stack[1][17] ), .Z(n2691) );
  NAND U2846 ( .A(n2383), .B(n2382), .Z(n2387) );
  NAND U2847 ( .A(n2385), .B(n2384), .Z(n2386) );
  NAND U2848 ( .A(n2387), .B(n2386), .Z(n2690) );
  XOR U2849 ( .A(n2691), .B(n2690), .Z(n2692) );
  XOR U2850 ( .A(n2632), .B(n2633), .Z(n2635) );
  AND U2851 ( .A(o[11]), .B(\stack[1][16] ), .Z(n2634) );
  XOR U2852 ( .A(n2635), .B(n2634), .Z(n2629) );
  AND U2853 ( .A(o[12]), .B(\stack[1][15] ), .Z(n2627) );
  NAND U2854 ( .A(n2389), .B(n2388), .Z(n2393) );
  NAND U2855 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U2856 ( .A(n2393), .B(n2392), .Z(n2626) );
  XOR U2857 ( .A(n2627), .B(n2626), .Z(n2628) );
  XNOR U2858 ( .A(n2629), .B(n2628), .Z(n2697) );
  NAND U2859 ( .A(\stack[1][14] ), .B(o[13]), .Z(n2698) );
  XNOR U2860 ( .A(n2699), .B(n2698), .Z(n2705) );
  AND U2861 ( .A(\stack[1][13] ), .B(o[14]), .Z(n2703) );
  NAND U2862 ( .A(n2395), .B(n2394), .Z(n2399) );
  NAND U2863 ( .A(n2397), .B(n2396), .Z(n2398) );
  NAND U2864 ( .A(n2399), .B(n2398), .Z(n2702) );
  XOR U2865 ( .A(n2703), .B(n2702), .Z(n2704) );
  XOR U2866 ( .A(n2621), .B(n2620), .Z(n2622) );
  XOR U2867 ( .A(n2623), .B(n2622), .Z(n2711) );
  AND U2868 ( .A(\stack[1][11] ), .B(o[16]), .Z(n2709) );
  NAND U2869 ( .A(n2401), .B(n2400), .Z(n2405) );
  NAND U2870 ( .A(n2403), .B(n2402), .Z(n2404) );
  NAND U2871 ( .A(n2405), .B(n2404), .Z(n2708) );
  XOR U2872 ( .A(n2709), .B(n2708), .Z(n2710) );
  XOR U2873 ( .A(n2711), .B(n2710), .Z(n2614) );
  XOR U2874 ( .A(n2615), .B(n2614), .Z(n2616) );
  XOR U2875 ( .A(n2617), .B(n2616), .Z(n2717) );
  AND U2876 ( .A(\stack[1][9] ), .B(o[18]), .Z(n2715) );
  AND U2877 ( .A(\stack[1][9] ), .B(o[16]), .Z(n2496) );
  XOR U2878 ( .A(n2407), .B(n2406), .Z(n2490) );
  AND U2879 ( .A(\stack[1][9] ), .B(o[14]), .Z(n2486) );
  AND U2880 ( .A(\stack[1][9] ), .B(o[12]), .Z(n2476) );
  XNOR U2881 ( .A(n2411), .B(n2410), .Z(n2469) );
  AND U2882 ( .A(o[10]), .B(\stack[1][9] ), .Z(n2466) );
  AND U2883 ( .A(o[0]), .B(\stack[1][9] ), .Z(n2412) );
  AND U2884 ( .A(\stack[1][10] ), .B(o[1]), .Z(n2415) );
  AND U2885 ( .A(n2412), .B(n2415), .Z(n2413) );
  NAND U2886 ( .A(o[2]), .B(n2413), .Z(n2419) );
  NAND U2887 ( .A(\stack[1][11] ), .B(o[0]), .Z(n2414) );
  XNOR U2888 ( .A(n2415), .B(n2414), .Z(n2521) );
  NAND U2889 ( .A(n2415), .B(o[0]), .Z(n2416) );
  XNOR U2890 ( .A(o[2]), .B(n2416), .Z(n2417) );
  AND U2891 ( .A(\stack[1][9] ), .B(n2417), .Z(n2522) );
  NAND U2892 ( .A(n2521), .B(n2522), .Z(n2418) );
  NAND U2893 ( .A(n2419), .B(n2418), .Z(n2422) );
  NAND U2894 ( .A(n2422), .B(n2423), .Z(n2425) );
  AND U2895 ( .A(o[3]), .B(\stack[1][9] ), .Z(n2528) );
  NAND U2896 ( .A(n2528), .B(n2527), .Z(n2424) );
  NAND U2897 ( .A(n2425), .B(n2424), .Z(n2426) );
  AND U2898 ( .A(o[4]), .B(\stack[1][9] ), .Z(n2427) );
  NAND U2899 ( .A(n2426), .B(n2427), .Z(n2431) );
  NAND U2900 ( .A(n2512), .B(n2511), .Z(n2430) );
  NAND U2901 ( .A(n2431), .B(n2430), .Z(n2434) );
  XOR U2902 ( .A(n2433), .B(n2432), .Z(n2435) );
  NAND U2903 ( .A(n2434), .B(n2435), .Z(n2438) );
  AND U2904 ( .A(o[5]), .B(\stack[1][9] ), .Z(n2537) );
  IV U2905 ( .A(n2434), .Z(n2436) );
  XNOR U2906 ( .A(n2436), .B(n2435), .Z(n2538) );
  NAND U2907 ( .A(n2537), .B(n2538), .Z(n2437) );
  NAND U2908 ( .A(n2438), .B(n2437), .Z(n2441) );
  NAND U2909 ( .A(n2441), .B(n2442), .Z(n2444) );
  AND U2910 ( .A(o[6]), .B(\stack[1][9] ), .Z(n2544) );
  NAND U2911 ( .A(n2544), .B(n2543), .Z(n2443) );
  NAND U2912 ( .A(n2444), .B(n2443), .Z(n2447) );
  NAND U2913 ( .A(n2447), .B(n2448), .Z(n2450) );
  AND U2914 ( .A(\stack[1][9] ), .B(o[7]), .Z(n2550) );
  NAND U2915 ( .A(n2550), .B(n2551), .Z(n2449) );
  NAND U2916 ( .A(n2450), .B(n2449), .Z(n2453) );
  AND U2917 ( .A(\stack[1][9] ), .B(o[8]), .Z(n2454) );
  NAND U2918 ( .A(n2453), .B(n2454), .Z(n2456) );
  XOR U2919 ( .A(n2452), .B(n2451), .Z(n2510) );
  NAND U2920 ( .A(n2510), .B(n2509), .Z(n2455) );
  NAND U2921 ( .A(n2456), .B(n2455), .Z(n2459) );
  XOR U2922 ( .A(n2458), .B(n2457), .Z(n2460) );
  NAND U2923 ( .A(n2459), .B(n2460), .Z(n2462) );
  AND U2924 ( .A(\stack[1][9] ), .B(o[9]), .Z(n2558) );
  NAND U2925 ( .A(n2558), .B(n2559), .Z(n2461) );
  NAND U2926 ( .A(n2462), .B(n2461), .Z(n2465) );
  NAND U2927 ( .A(n2466), .B(n2465), .Z(n2468) );
  XNOR U2928 ( .A(n2464), .B(n2463), .Z(n2564) );
  XOR U2929 ( .A(n2466), .B(n2465), .Z(n2565) );
  NAND U2930 ( .A(n2564), .B(n2565), .Z(n2467) );
  AND U2931 ( .A(n2468), .B(n2467), .Z(n2470) );
  NAND U2932 ( .A(n2469), .B(n2470), .Z(n2472) );
  NAND U2933 ( .A(\stack[1][9] ), .B(o[11]), .Z(n2572) );
  NAND U2934 ( .A(n2573), .B(n2572), .Z(n2471) );
  AND U2935 ( .A(n2472), .B(n2471), .Z(n2475) );
  NAND U2936 ( .A(n2476), .B(n2475), .Z(n2478) );
  XNOR U2937 ( .A(n2474), .B(n2473), .Z(n2577) );
  XOR U2938 ( .A(n2476), .B(n2475), .Z(n2576) );
  NAND U2939 ( .A(n2577), .B(n2576), .Z(n2477) );
  NAND U2940 ( .A(n2478), .B(n2477), .Z(n2479) );
  NAND U2941 ( .A(n2480), .B(n2479), .Z(n2482) );
  XOR U2942 ( .A(n2480), .B(n2479), .Z(n2585) );
  AND U2943 ( .A(\stack[1][9] ), .B(o[13]), .Z(n2584) );
  NAND U2944 ( .A(n2585), .B(n2584), .Z(n2481) );
  NAND U2945 ( .A(n2482), .B(n2481), .Z(n2485) );
  NAND U2946 ( .A(n2486), .B(n2485), .Z(n2488) );
  XOR U2947 ( .A(n2484), .B(n2483), .Z(n2508) );
  XOR U2948 ( .A(n2486), .B(n2485), .Z(n2507) );
  NAND U2949 ( .A(n2508), .B(n2507), .Z(n2487) );
  NAND U2950 ( .A(n2488), .B(n2487), .Z(n2489) );
  NAND U2951 ( .A(n2490), .B(n2489), .Z(n2492) );
  XOR U2952 ( .A(n2490), .B(n2489), .Z(n2595) );
  AND U2953 ( .A(\stack[1][9] ), .B(o[15]), .Z(n2594) );
  NAND U2954 ( .A(n2595), .B(n2594), .Z(n2491) );
  NAND U2955 ( .A(n2492), .B(n2491), .Z(n2495) );
  NAND U2956 ( .A(n2496), .B(n2495), .Z(n2498) );
  XOR U2957 ( .A(n2494), .B(n2493), .Z(n2506) );
  XOR U2958 ( .A(n2496), .B(n2495), .Z(n2505) );
  NAND U2959 ( .A(n2506), .B(n2505), .Z(n2497) );
  NAND U2960 ( .A(n2498), .B(n2497), .Z(n2502) );
  XNOR U2961 ( .A(n2500), .B(n2499), .Z(n2501) );
  NAND U2962 ( .A(n2502), .B(n2501), .Z(n2504) );
  XOR U2963 ( .A(n2502), .B(n2501), .Z(n2605) );
  AND U2964 ( .A(\stack[1][9] ), .B(o[17]), .Z(n2604) );
  NAND U2965 ( .A(n2605), .B(n2604), .Z(n2503) );
  NAND U2966 ( .A(n2504), .B(n2503), .Z(n2714) );
  XOR U2967 ( .A(n2715), .B(n2714), .Z(n2716) );
  XOR U2968 ( .A(n2717), .B(n2716), .Z(n2608) );
  AND U2969 ( .A(\stack[1][8] ), .B(o[18]), .Z(n2602) );
  XOR U2970 ( .A(n2506), .B(n2505), .Z(n2598) );
  AND U2971 ( .A(\stack[1][8] ), .B(o[16]), .Z(n2592) );
  XOR U2972 ( .A(n2508), .B(n2507), .Z(n2588) );
  NAND U2973 ( .A(\stack[1][8] ), .B(o[12]), .Z(n2570) );
  AND U2974 ( .A(o[10]), .B(\stack[1][8] ), .Z(n2560) );
  XNOR U2975 ( .A(n2510), .B(n2509), .Z(n2554) );
  AND U2976 ( .A(\stack[1][8] ), .B(o[5]), .Z(n2533) );
  XOR U2977 ( .A(n2512), .B(n2511), .Z(n2534) );
  NAND U2978 ( .A(n2533), .B(n2534), .Z(n2536) );
  AND U2979 ( .A(o[0]), .B(\stack[1][8] ), .Z(n2513) );
  AND U2980 ( .A(o[1]), .B(\stack[1][9] ), .Z(n2518) );
  AND U2981 ( .A(n2513), .B(n2518), .Z(n2514) );
  NAND U2982 ( .A(o[2]), .B(n2514), .Z(n2520) );
  NAND U2983 ( .A(n2518), .B(o[0]), .Z(n2515) );
  XNOR U2984 ( .A(o[2]), .B(n2515), .Z(n2516) );
  AND U2985 ( .A(\stack[1][8] ), .B(n2516), .Z(n2851) );
  NAND U2986 ( .A(\stack[1][10] ), .B(o[0]), .Z(n2517) );
  XNOR U2987 ( .A(n2518), .B(n2517), .Z(n2852) );
  NAND U2988 ( .A(n2851), .B(n2852), .Z(n2519) );
  NAND U2989 ( .A(n2520), .B(n2519), .Z(n2523) );
  NAND U2990 ( .A(n2523), .B(n2524), .Z(n2526) );
  AND U2991 ( .A(o[3]), .B(\stack[1][8] ), .Z(n2859) );
  NAND U2992 ( .A(n2860), .B(n2859), .Z(n2525) );
  NAND U2993 ( .A(n2526), .B(n2525), .Z(n2529) );
  AND U2994 ( .A(o[4]), .B(\stack[1][8] ), .Z(n2530) );
  NAND U2995 ( .A(n2529), .B(n2530), .Z(n2532) );
  XOR U2996 ( .A(n2528), .B(n2527), .Z(n2864) );
  NAND U2997 ( .A(n2864), .B(n2863), .Z(n2531) );
  NAND U2998 ( .A(n2532), .B(n2531), .Z(n2869) );
  NAND U2999 ( .A(n2869), .B(n2870), .Z(n2535) );
  NAND U3000 ( .A(n2536), .B(n2535), .Z(n2539) );
  NAND U3001 ( .A(n2539), .B(n2540), .Z(n2542) );
  AND U3002 ( .A(\stack[1][8] ), .B(o[6]), .Z(n2875) );
  NAND U3003 ( .A(n2875), .B(n2876), .Z(n2541) );
  NAND U3004 ( .A(n2542), .B(n2541), .Z(n2545) );
  XOR U3005 ( .A(n2544), .B(n2543), .Z(n2546) );
  NAND U3006 ( .A(n2545), .B(n2546), .Z(n2548) );
  AND U3007 ( .A(\stack[1][8] ), .B(o[7]), .Z(n2882) );
  NAND U3008 ( .A(n2882), .B(n2881), .Z(n2547) );
  NAND U3009 ( .A(n2548), .B(n2547), .Z(n2549) );
  AND U3010 ( .A(\stack[1][8] ), .B(o[8]), .Z(n5315) );
  NAND U3011 ( .A(n2549), .B(n5315), .Z(n2553) );
  NAND U3012 ( .A(n2888), .B(n2887), .Z(n2552) );
  AND U3013 ( .A(n2553), .B(n2552), .Z(n2555) );
  NAND U3014 ( .A(n2554), .B(n2555), .Z(n2557) );
  NAND U3015 ( .A(\stack[1][8] ), .B(o[9]), .Z(n2893) );
  NAND U3016 ( .A(n2894), .B(n2893), .Z(n2556) );
  AND U3017 ( .A(n2557), .B(n2556), .Z(n2561) );
  NAND U3018 ( .A(n2560), .B(n2561), .Z(n2563) );
  NAND U3019 ( .A(n2842), .B(n2841), .Z(n2562) );
  NAND U3020 ( .A(n2563), .B(n2562), .Z(n2566) );
  NAND U3021 ( .A(n2566), .B(n2567), .Z(n2569) );
  AND U3022 ( .A(\stack[1][8] ), .B(o[11]), .Z(n2904) );
  NAND U3023 ( .A(n2904), .B(n2903), .Z(n2568) );
  AND U3024 ( .A(n2569), .B(n2568), .Z(n2571) );
  NAND U3025 ( .A(n2570), .B(n2571), .Z(n2575) );
  XOR U3026 ( .A(n2573), .B(n2572), .Z(n2909) );
  NAND U3027 ( .A(n2910), .B(n2909), .Z(n2574) );
  NAND U3028 ( .A(n2575), .B(n2574), .Z(n2579) );
  XNOR U3029 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U3030 ( .A(n2579), .B(n2578), .Z(n2581) );
  XOR U3031 ( .A(n2579), .B(n2578), .Z(n2916) );
  NAND U3032 ( .A(\stack[1][8] ), .B(o[13]), .Z(n2915) );
  NAND U3033 ( .A(n2916), .B(n2915), .Z(n2580) );
  AND U3034 ( .A(n2581), .B(n2580), .Z(n2583) );
  AND U3035 ( .A(\stack[1][8] ), .B(o[14]), .Z(n2582) );
  NAND U3036 ( .A(n2583), .B(n2582), .Z(n2587) );
  XOR U3037 ( .A(n2583), .B(n2582), .Z(n2840) );
  XOR U3038 ( .A(n2585), .B(n2584), .Z(n2839) );
  NAND U3039 ( .A(n2840), .B(n2839), .Z(n2586) );
  NAND U3040 ( .A(n2587), .B(n2586), .Z(n2589) );
  NAND U3041 ( .A(n2588), .B(n2589), .Z(n2591) );
  XOR U3042 ( .A(n2589), .B(n2588), .Z(n2926) );
  AND U3043 ( .A(\stack[1][8] ), .B(o[15]), .Z(n2925) );
  NAND U3044 ( .A(n2926), .B(n2925), .Z(n2590) );
  NAND U3045 ( .A(n2591), .B(n2590), .Z(n2593) );
  NAND U3046 ( .A(n2592), .B(n2593), .Z(n2597) );
  XOR U3047 ( .A(n2593), .B(n2592), .Z(n2838) );
  XOR U3048 ( .A(n2595), .B(n2594), .Z(n2837) );
  NAND U3049 ( .A(n2838), .B(n2837), .Z(n2596) );
  NAND U3050 ( .A(n2597), .B(n2596), .Z(n2599) );
  NAND U3051 ( .A(n2598), .B(n2599), .Z(n2601) );
  XOR U3052 ( .A(n2599), .B(n2598), .Z(n2936) );
  AND U3053 ( .A(\stack[1][8] ), .B(o[17]), .Z(n2935) );
  NAND U3054 ( .A(n2936), .B(n2935), .Z(n2600) );
  NAND U3055 ( .A(n2601), .B(n2600), .Z(n2603) );
  NAND U3056 ( .A(n2602), .B(n2603), .Z(n2607) );
  XOR U3057 ( .A(n2603), .B(n2602), .Z(n2836) );
  XOR U3058 ( .A(n2605), .B(n2604), .Z(n2835) );
  NAND U3059 ( .A(n2836), .B(n2835), .Z(n2606) );
  NAND U3060 ( .A(n2607), .B(n2606), .Z(n2609) );
  NAND U3061 ( .A(n2608), .B(n2609), .Z(n2611) );
  XOR U3062 ( .A(n2609), .B(n2608), .Z(n2945) );
  AND U3063 ( .A(\stack[1][8] ), .B(o[19]), .Z(n2946) );
  NAND U3064 ( .A(n2945), .B(n2946), .Z(n2610) );
  NAND U3065 ( .A(n2611), .B(n2610), .Z(n2613) );
  NAND U3066 ( .A(n2612), .B(n2613), .Z(n2721) );
  XOR U3067 ( .A(n2613), .B(n2612), .Z(n2834) );
  NAND U3068 ( .A(n2615), .B(n2614), .Z(n2619) );
  NAND U3069 ( .A(n2617), .B(n2616), .Z(n2618) );
  NAND U3070 ( .A(n2619), .B(n2618), .Z(n2722) );
  AND U3071 ( .A(\stack[1][10] ), .B(o[18]), .Z(n2723) );
  XOR U3072 ( .A(n2722), .B(n2723), .Z(n2725) );
  NAND U3073 ( .A(n2621), .B(n2620), .Z(n2625) );
  NAND U3074 ( .A(n2623), .B(n2622), .Z(n2624) );
  NAND U3075 ( .A(n2625), .B(n2624), .Z(n2728) );
  AND U3076 ( .A(\stack[1][12] ), .B(o[16]), .Z(n2729) );
  XOR U3077 ( .A(n2728), .B(n2729), .Z(n2731) );
  NAND U3078 ( .A(n2627), .B(n2626), .Z(n2631) );
  NAND U3079 ( .A(n2629), .B(n2628), .Z(n2630) );
  NAND U3080 ( .A(n2631), .B(n2630), .Z(n2810) );
  NAND U3081 ( .A(n2633), .B(n2632), .Z(n2637) );
  NAND U3082 ( .A(n2635), .B(n2634), .Z(n2636) );
  AND U3083 ( .A(n2637), .B(n2636), .Z(n2740) );
  NAND U3084 ( .A(o[12]), .B(\stack[1][16] ), .Z(n2739) );
  XOR U3085 ( .A(n2740), .B(n2739), .Z(n2742) );
  AND U3086 ( .A(o[6]), .B(\stack[1][22] ), .Z(n2760) );
  NAND U3087 ( .A(n2639), .B(n2638), .Z(n2643) );
  NAND U3088 ( .A(n2641), .B(n2640), .Z(n2642) );
  NAND U3089 ( .A(n2643), .B(n2642), .Z(n2785) );
  AND U3090 ( .A(o[3]), .B(\stack[1][25] ), .Z(n2765) );
  AND U3091 ( .A(o[0]), .B(\stack[1][25] ), .Z(n2645) );
  AND U3092 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U3093 ( .A(o[2]), .B(n2646), .Z(n2650) );
  NAND U3094 ( .A(n2648), .B(n2647), .Z(n2649) );
  NAND U3095 ( .A(n2650), .B(n2649), .Z(n2763) );
  AND U3096 ( .A(o[1]), .B(\stack[1][27] ), .Z(n2772) );
  NAND U3097 ( .A(\stack[1][28] ), .B(o[0]), .Z(n2651) );
  XNOR U3098 ( .A(n2772), .B(n2651), .Z(n2776) );
  NAND U3099 ( .A(n2772), .B(o[0]), .Z(n2652) );
  XNOR U3100 ( .A(o[2]), .B(n2652), .Z(n2653) );
  AND U3101 ( .A(\stack[1][26] ), .B(n2653), .Z(n2775) );
  XOR U3102 ( .A(n2776), .B(n2775), .Z(n2764) );
  XOR U3103 ( .A(n2763), .B(n2764), .Z(n2766) );
  AND U3104 ( .A(o[4]), .B(\stack[1][24] ), .Z(n2780) );
  NAND U3105 ( .A(n2655), .B(n2654), .Z(n2659) );
  NAND U3106 ( .A(n2657), .B(n2656), .Z(n2658) );
  NAND U3107 ( .A(n2659), .B(n2658), .Z(n2779) );
  XOR U3108 ( .A(n2780), .B(n2779), .Z(n2781) );
  XOR U3109 ( .A(n2782), .B(n2781), .Z(n2786) );
  XOR U3110 ( .A(n2785), .B(n2786), .Z(n2788) );
  AND U3111 ( .A(o[5]), .B(\stack[1][23] ), .Z(n2787) );
  XOR U3112 ( .A(n2788), .B(n2787), .Z(n2758) );
  NAND U3113 ( .A(n2661), .B(n2660), .Z(n2665) );
  NAND U3114 ( .A(n2663), .B(n2662), .Z(n2664) );
  NAND U3115 ( .A(n2665), .B(n2664), .Z(n2757) );
  XOR U3116 ( .A(n2758), .B(n2757), .Z(n2759) );
  XOR U3117 ( .A(n2760), .B(n2759), .Z(n2792) );
  NAND U3118 ( .A(n2667), .B(n2666), .Z(n2671) );
  NAND U3119 ( .A(n2669), .B(n2668), .Z(n2670) );
  NAND U3120 ( .A(n2671), .B(n2670), .Z(n2791) );
  XOR U3121 ( .A(n2792), .B(n2791), .Z(n2794) );
  AND U3122 ( .A(o[7]), .B(\stack[1][21] ), .Z(n2793) );
  XNOR U3123 ( .A(n2794), .B(n2793), .Z(n2754) );
  NAND U3124 ( .A(n2673), .B(n2672), .Z(n2677) );
  NAND U3125 ( .A(n2675), .B(n2674), .Z(n2676) );
  AND U3126 ( .A(n2677), .B(n2676), .Z(n2752) );
  NAND U3127 ( .A(o[8]), .B(\stack[1][20] ), .Z(n2751) );
  XOR U3128 ( .A(n2752), .B(n2751), .Z(n2753) );
  NAND U3129 ( .A(n2679), .B(n2678), .Z(n2683) );
  NAND U3130 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U3131 ( .A(n2683), .B(n2682), .Z(n2797) );
  AND U3132 ( .A(o[9]), .B(\stack[1][19] ), .Z(n2799) );
  XNOR U3133 ( .A(n2800), .B(n2799), .Z(n2748) );
  NAND U3134 ( .A(n2685), .B(n2684), .Z(n2689) );
  NAND U3135 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3136 ( .A(n2689), .B(n2688), .Z(n2746) );
  NAND U3137 ( .A(o[10]), .B(\stack[1][18] ), .Z(n2745) );
  XOR U3138 ( .A(n2746), .B(n2745), .Z(n2747) );
  NAND U3139 ( .A(n2691), .B(n2690), .Z(n2695) );
  NAND U3140 ( .A(n2693), .B(n2692), .Z(n2694) );
  AND U3141 ( .A(n2695), .B(n2694), .Z(n2803) );
  XOR U3142 ( .A(n2804), .B(n2803), .Z(n2806) );
  NAND U3143 ( .A(o[11]), .B(\stack[1][17] ), .Z(n2805) );
  XOR U3144 ( .A(n2806), .B(n2805), .Z(n2741) );
  XNOR U3145 ( .A(n2742), .B(n2741), .Z(n2809) );
  XOR U3146 ( .A(n2810), .B(n2809), .Z(n2812) );
  AND U3147 ( .A(\stack[1][15] ), .B(o[13]), .Z(n2811) );
  XNOR U3148 ( .A(n2812), .B(n2811), .Z(n2736) );
  NAND U3149 ( .A(\stack[1][14] ), .B(o[14]), .Z(n5088) );
  NAND U3150 ( .A(n2697), .B(n2696), .Z(n2701) );
  NAND U3151 ( .A(n2699), .B(n2698), .Z(n2700) );
  NAND U3152 ( .A(n2701), .B(n2700), .Z(n2734) );
  XOR U3153 ( .A(n5088), .B(n2734), .Z(n2735) );
  NAND U3154 ( .A(n2703), .B(n2702), .Z(n2707) );
  NAND U3155 ( .A(n2705), .B(n2704), .Z(n2706) );
  NAND U3156 ( .A(n2707), .B(n2706), .Z(n2815) );
  AND U3157 ( .A(\stack[1][13] ), .B(o[15]), .Z(n2817) );
  XOR U3158 ( .A(n2818), .B(n2817), .Z(n2730) );
  XOR U3159 ( .A(n2731), .B(n2730), .Z(n2822) );
  NAND U3160 ( .A(n2709), .B(n2708), .Z(n2713) );
  NAND U3161 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U3162 ( .A(n2713), .B(n2712), .Z(n2821) );
  XOR U3163 ( .A(n2822), .B(n2821), .Z(n2824) );
  AND U3164 ( .A(\stack[1][11] ), .B(o[17]), .Z(n2823) );
  XOR U3165 ( .A(n2824), .B(n2823), .Z(n2724) );
  XOR U3166 ( .A(n2725), .B(n2724), .Z(n2828) );
  NAND U3167 ( .A(n2715), .B(n2714), .Z(n2719) );
  NAND U3168 ( .A(n2717), .B(n2716), .Z(n2718) );
  NAND U3169 ( .A(n2719), .B(n2718), .Z(n2827) );
  XOR U3170 ( .A(n2828), .B(n2827), .Z(n2830) );
  AND U3171 ( .A(\stack[1][9] ), .B(o[19]), .Z(n2829) );
  XOR U3172 ( .A(n2830), .B(n2829), .Z(n2833) );
  NAND U3173 ( .A(n2834), .B(n2833), .Z(n2720) );
  NAND U3174 ( .A(n2721), .B(n2720), .Z(n3087) );
  AND U3175 ( .A(\stack[1][10] ), .B(o[19]), .Z(n3095) );
  NAND U3176 ( .A(n2723), .B(n2722), .Z(n2727) );
  NAND U3177 ( .A(n2725), .B(n2724), .Z(n2726) );
  NAND U3178 ( .A(n2727), .B(n2726), .Z(n3093) );
  AND U3179 ( .A(\stack[1][12] ), .B(o[17]), .Z(n3195) );
  NAND U3180 ( .A(n2729), .B(n2728), .Z(n2733) );
  NAND U3181 ( .A(n2731), .B(n2730), .Z(n2732) );
  NAND U3182 ( .A(n2733), .B(n2732), .Z(n3193) );
  AND U3183 ( .A(\stack[1][14] ), .B(o[15]), .Z(n3108) );
  NAND U3184 ( .A(n5088), .B(n2734), .Z(n2738) );
  NAND U3185 ( .A(n2736), .B(n2735), .Z(n2737) );
  AND U3186 ( .A(n2738), .B(n2737), .Z(n3106) );
  NAND U3187 ( .A(o[13]), .B(\stack[1][16] ), .Z(n3183) );
  NAND U3188 ( .A(n2740), .B(n2739), .Z(n2744) );
  NAND U3189 ( .A(n2742), .B(n2741), .Z(n2743) );
  NAND U3190 ( .A(n2744), .B(n2743), .Z(n3182) );
  AND U3191 ( .A(o[11]), .B(\stack[1][18] ), .Z(n3120) );
  NAND U3192 ( .A(n2746), .B(n2745), .Z(n2750) );
  NAND U3193 ( .A(n2748), .B(n2747), .Z(n2749) );
  AND U3194 ( .A(n2750), .B(n2749), .Z(n3118) );
  NAND U3195 ( .A(n2752), .B(n2751), .Z(n2756) );
  NAND U3196 ( .A(n2754), .B(n2753), .Z(n2755) );
  NAND U3197 ( .A(n2756), .B(n2755), .Z(n3170) );
  AND U3198 ( .A(o[7]), .B(\stack[1][22] ), .Z(n3125) );
  NAND U3199 ( .A(n2758), .B(n2757), .Z(n2762) );
  NAND U3200 ( .A(n2760), .B(n2759), .Z(n2761) );
  NAND U3201 ( .A(n2762), .B(n2761), .Z(n3123) );
  AND U3202 ( .A(o[6]), .B(\stack[1][23] ), .Z(n3160) );
  NAND U3203 ( .A(n2764), .B(n2763), .Z(n2768) );
  NAND U3204 ( .A(n2766), .B(n2765), .Z(n2767) );
  NAND U3205 ( .A(n2768), .B(n2767), .Z(n3129) );
  AND U3206 ( .A(o[4]), .B(\stack[1][25] ), .Z(n3130) );
  XOR U3207 ( .A(n3129), .B(n3130), .Z(n3132) );
  AND U3208 ( .A(o[1]), .B(\stack[1][28] ), .Z(n3135) );
  NAND U3209 ( .A(\stack[1][29] ), .B(o[0]), .Z(n2769) );
  XNOR U3210 ( .A(n3135), .B(n2769), .Z(n3139) );
  NAND U3211 ( .A(n3135), .B(o[0]), .Z(n2770) );
  XNOR U3212 ( .A(o[2]), .B(n2770), .Z(n2771) );
  AND U3213 ( .A(\stack[1][27] ), .B(n2771), .Z(n3138) );
  XOR U3214 ( .A(n3139), .B(n3138), .Z(n3148) );
  AND U3215 ( .A(o[0]), .B(\stack[1][26] ), .Z(n2773) );
  AND U3216 ( .A(n2773), .B(n2772), .Z(n2774) );
  NAND U3217 ( .A(o[2]), .B(n2774), .Z(n2778) );
  NAND U3218 ( .A(n2776), .B(n2775), .Z(n2777) );
  NAND U3219 ( .A(n2778), .B(n2777), .Z(n3145) );
  AND U3220 ( .A(o[3]), .B(\stack[1][26] ), .Z(n3146) );
  XOR U3221 ( .A(n3145), .B(n3146), .Z(n3147) );
  XOR U3222 ( .A(n3148), .B(n3147), .Z(n3131) );
  XOR U3223 ( .A(n3132), .B(n3131), .Z(n3152) );
  AND U3224 ( .A(o[5]), .B(\stack[1][24] ), .Z(n3151) );
  XOR U3225 ( .A(n3152), .B(n3151), .Z(n3154) );
  NAND U3226 ( .A(n2780), .B(n2779), .Z(n2784) );
  NAND U3227 ( .A(n2782), .B(n2781), .Z(n2783) );
  NAND U3228 ( .A(n2784), .B(n2783), .Z(n3153) );
  XOR U3229 ( .A(n3154), .B(n3153), .Z(n3158) );
  NAND U3230 ( .A(n2786), .B(n2785), .Z(n2790) );
  NAND U3231 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U3232 ( .A(n2790), .B(n2789), .Z(n3157) );
  XOR U3233 ( .A(n3158), .B(n3157), .Z(n3159) );
  XOR U3234 ( .A(n3160), .B(n3159), .Z(n3124) );
  XOR U3235 ( .A(n3123), .B(n3124), .Z(n3126) );
  AND U3236 ( .A(o[8]), .B(\stack[1][21] ), .Z(n3164) );
  NAND U3237 ( .A(n2792), .B(n2791), .Z(n2796) );
  NAND U3238 ( .A(n2794), .B(n2793), .Z(n2795) );
  NAND U3239 ( .A(n2796), .B(n2795), .Z(n3163) );
  XOR U3240 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U3241 ( .A(n3166), .B(n3165), .Z(n3169) );
  XOR U3242 ( .A(n3170), .B(n3169), .Z(n3172) );
  NAND U3243 ( .A(o[9]), .B(\stack[1][20] ), .Z(n3171) );
  XNOR U3244 ( .A(n3172), .B(n3171), .Z(n3178) );
  AND U3245 ( .A(o[10]), .B(\stack[1][19] ), .Z(n3176) );
  NAND U3246 ( .A(n2798), .B(n2797), .Z(n2802) );
  NAND U3247 ( .A(n2800), .B(n2799), .Z(n2801) );
  NAND U3248 ( .A(n2802), .B(n2801), .Z(n3175) );
  XOR U3249 ( .A(n3176), .B(n3175), .Z(n3177) );
  XOR U3250 ( .A(n3118), .B(n3117), .Z(n3119) );
  XOR U3251 ( .A(n3120), .B(n3119), .Z(n3114) );
  AND U3252 ( .A(o[12]), .B(\stack[1][17] ), .Z(n3112) );
  NAND U3253 ( .A(n2804), .B(n2803), .Z(n2808) );
  NAND U3254 ( .A(n2806), .B(n2805), .Z(n2807) );
  AND U3255 ( .A(n2808), .B(n2807), .Z(n3111) );
  XOR U3256 ( .A(n3112), .B(n3111), .Z(n3113) );
  XNOR U3257 ( .A(n3114), .B(n3113), .Z(n3181) );
  XOR U3258 ( .A(n3182), .B(n3181), .Z(n3184) );
  XNOR U3259 ( .A(n3183), .B(n3184), .Z(n3190) );
  AND U3260 ( .A(\stack[1][15] ), .B(o[14]), .Z(n3188) );
  NAND U3261 ( .A(n2810), .B(n2809), .Z(n2814) );
  NAND U3262 ( .A(n2812), .B(n2811), .Z(n2813) );
  NAND U3263 ( .A(n2814), .B(n2813), .Z(n3187) );
  XOR U3264 ( .A(n3188), .B(n3187), .Z(n3189) );
  XOR U3265 ( .A(n3106), .B(n3105), .Z(n3107) );
  XOR U3266 ( .A(n3108), .B(n3107), .Z(n3102) );
  AND U3267 ( .A(\stack[1][13] ), .B(o[16]), .Z(n3100) );
  NAND U3268 ( .A(n2816), .B(n2815), .Z(n2820) );
  NAND U3269 ( .A(n2818), .B(n2817), .Z(n2819) );
  NAND U3270 ( .A(n2820), .B(n2819), .Z(n3099) );
  XOR U3271 ( .A(n3100), .B(n3099), .Z(n3101) );
  XOR U3272 ( .A(n3102), .B(n3101), .Z(n3194) );
  XOR U3273 ( .A(n3193), .B(n3194), .Z(n3196) );
  AND U3274 ( .A(\stack[1][11] ), .B(o[18]), .Z(n3200) );
  NAND U3275 ( .A(n2822), .B(n2821), .Z(n2826) );
  NAND U3276 ( .A(n2824), .B(n2823), .Z(n2825) );
  NAND U3277 ( .A(n2826), .B(n2825), .Z(n3199) );
  XOR U3278 ( .A(n3200), .B(n3199), .Z(n3201) );
  XOR U3279 ( .A(n3202), .B(n3201), .Z(n3094) );
  XOR U3280 ( .A(n3093), .B(n3094), .Z(n3096) );
  AND U3281 ( .A(\stack[1][9] ), .B(o[20]), .Z(n3206) );
  NAND U3282 ( .A(n2828), .B(n2827), .Z(n2832) );
  NAND U3283 ( .A(n2830), .B(n2829), .Z(n2831) );
  NAND U3284 ( .A(n2832), .B(n2831), .Z(n3205) );
  XOR U3285 ( .A(n3206), .B(n3205), .Z(n3207) );
  XOR U3286 ( .A(n3208), .B(n3207), .Z(n3088) );
  XOR U3287 ( .A(n3087), .B(n3088), .Z(n3090) );
  AND U3288 ( .A(\stack[1][7] ), .B(o[22]), .Z(n3212) );
  XOR U3289 ( .A(n2834), .B(n2833), .Z(n2952) );
  AND U3290 ( .A(\stack[1][7] ), .B(o[20]), .Z(n2948) );
  XOR U3291 ( .A(n2836), .B(n2835), .Z(n2942) );
  AND U3292 ( .A(\stack[1][7] ), .B(o[18]), .Z(n2938) );
  XOR U3293 ( .A(n2838), .B(n2837), .Z(n2932) );
  AND U3294 ( .A(\stack[1][7] ), .B(o[16]), .Z(n2928) );
  XOR U3295 ( .A(n2840), .B(n2839), .Z(n2922) );
  AND U3296 ( .A(\stack[1][7] ), .B(o[14]), .Z(n2918) );
  XNOR U3297 ( .A(n2842), .B(n2841), .Z(n2899) );
  NAND U3298 ( .A(o[4]), .B(\stack[1][7] ), .Z(n2857) );
  AND U3299 ( .A(o[0]), .B(\stack[1][7] ), .Z(n2843) );
  AND U3300 ( .A(o[1]), .B(\stack[1][8] ), .Z(n2848) );
  AND U3301 ( .A(n2843), .B(n2848), .Z(n2844) );
  NAND U3302 ( .A(o[2]), .B(n2844), .Z(n2850) );
  NAND U3303 ( .A(n2848), .B(o[0]), .Z(n2845) );
  XNOR U3304 ( .A(o[2]), .B(n2845), .Z(n2846) );
  AND U3305 ( .A(\stack[1][7] ), .B(n2846), .Z(n2973) );
  NAND U3306 ( .A(\stack[1][9] ), .B(o[0]), .Z(n2847) );
  XNOR U3307 ( .A(n2848), .B(n2847), .Z(n2974) );
  NAND U3308 ( .A(n2973), .B(n2974), .Z(n2849) );
  NAND U3309 ( .A(n2850), .B(n2849), .Z(n2853) );
  NAND U3310 ( .A(n2853), .B(n2854), .Z(n2856) );
  AND U3311 ( .A(o[3]), .B(\stack[1][7] ), .Z(n2980) );
  NAND U3312 ( .A(n2980), .B(n2979), .Z(n2855) );
  AND U3313 ( .A(n2856), .B(n2855), .Z(n2858) );
  NAND U3314 ( .A(n2857), .B(n2858), .Z(n2862) );
  XNOR U3315 ( .A(n2860), .B(n2859), .Z(n2963) );
  NAND U3316 ( .A(n2964), .B(n2963), .Z(n2861) );
  AND U3317 ( .A(n2862), .B(n2861), .Z(n2866) );
  XOR U3318 ( .A(n2864), .B(n2863), .Z(n2865) );
  NAND U3319 ( .A(n2866), .B(n2865), .Z(n2868) );
  AND U3320 ( .A(\stack[1][7] ), .B(o[5]), .Z(n2989) );
  XOR U3321 ( .A(n2866), .B(n2865), .Z(n2990) );
  NAND U3322 ( .A(n2989), .B(n2990), .Z(n2867) );
  NAND U3323 ( .A(n2868), .B(n2867), .Z(n2871) );
  NAND U3324 ( .A(n2871), .B(n2872), .Z(n2874) );
  AND U3325 ( .A(\stack[1][7] ), .B(o[6]), .Z(n2996) );
  NAND U3326 ( .A(n2996), .B(n2995), .Z(n2873) );
  NAND U3327 ( .A(n2874), .B(n2873), .Z(n2877) );
  NAND U3328 ( .A(n2877), .B(n2878), .Z(n2880) );
  AND U3329 ( .A(\stack[1][7] ), .B(o[7]), .Z(n5354) );
  NAND U3330 ( .A(n5354), .B(n3003), .Z(n2879) );
  NAND U3331 ( .A(n2880), .B(n2879), .Z(n2883) );
  AND U3332 ( .A(\stack[1][7] ), .B(o[8]), .Z(n2884) );
  NAND U3333 ( .A(n2883), .B(n2884), .Z(n2886) );
  XOR U3334 ( .A(n2882), .B(n2881), .Z(n2962) );
  NAND U3335 ( .A(n2962), .B(n2961), .Z(n2885) );
  NAND U3336 ( .A(n2886), .B(n2885), .Z(n2889) );
  XOR U3337 ( .A(n2888), .B(n2887), .Z(n2890) );
  NAND U3338 ( .A(n2889), .B(n2890), .Z(n2892) );
  AND U3339 ( .A(\stack[1][7] ), .B(o[9]), .Z(n3010) );
  NAND U3340 ( .A(n3010), .B(n3011), .Z(n2891) );
  NAND U3341 ( .A(n2892), .B(n2891), .Z(n2895) );
  AND U3342 ( .A(o[10]), .B(\stack[1][7] ), .Z(n2896) );
  NAND U3343 ( .A(n2895), .B(n2896), .Z(n2898) );
  XNOR U3344 ( .A(n2894), .B(n2893), .Z(n3016) );
  NAND U3345 ( .A(n3016), .B(n3017), .Z(n2897) );
  AND U3346 ( .A(n2898), .B(n2897), .Z(n2900) );
  NAND U3347 ( .A(n2899), .B(n2900), .Z(n2902) );
  NAND U3348 ( .A(\stack[1][7] ), .B(o[11]), .Z(n3024) );
  NAND U3349 ( .A(n3024), .B(n3025), .Z(n2901) );
  AND U3350 ( .A(n2902), .B(n2901), .Z(n2905) );
  AND U3351 ( .A(\stack[1][7] ), .B(o[12]), .Z(n2906) );
  NAND U3352 ( .A(n2905), .B(n2906), .Z(n2908) );
  XOR U3353 ( .A(n2904), .B(n2903), .Z(n3029) );
  NAND U3354 ( .A(n3029), .B(n3028), .Z(n2907) );
  NAND U3355 ( .A(n2908), .B(n2907), .Z(n2911) );
  XNOR U3356 ( .A(n2910), .B(n2909), .Z(n2912) );
  NAND U3357 ( .A(n2911), .B(n2912), .Z(n2914) );
  AND U3358 ( .A(\stack[1][7] ), .B(o[13]), .Z(n3034) );
  NAND U3359 ( .A(n3034), .B(n3035), .Z(n2913) );
  NAND U3360 ( .A(n2914), .B(n2913), .Z(n2917) );
  NAND U3361 ( .A(n2918), .B(n2917), .Z(n2920) );
  XNOR U3362 ( .A(n2916), .B(n2915), .Z(n3040) );
  XOR U3363 ( .A(n2918), .B(n2917), .Z(n3041) );
  NAND U3364 ( .A(n3040), .B(n3041), .Z(n2919) );
  NAND U3365 ( .A(n2920), .B(n2919), .Z(n2921) );
  NAND U3366 ( .A(n2922), .B(n2921), .Z(n2924) );
  XOR U3367 ( .A(n2922), .B(n2921), .Z(n3049) );
  AND U3368 ( .A(\stack[1][7] ), .B(o[15]), .Z(n3048) );
  NAND U3369 ( .A(n3049), .B(n3048), .Z(n2923) );
  NAND U3370 ( .A(n2924), .B(n2923), .Z(n2927) );
  NAND U3371 ( .A(n2928), .B(n2927), .Z(n2930) );
  XOR U3372 ( .A(n2926), .B(n2925), .Z(n2960) );
  XOR U3373 ( .A(n2928), .B(n2927), .Z(n2959) );
  NAND U3374 ( .A(n2960), .B(n2959), .Z(n2929) );
  NAND U3375 ( .A(n2930), .B(n2929), .Z(n2931) );
  NAND U3376 ( .A(n2932), .B(n2931), .Z(n2934) );
  XOR U3377 ( .A(n2932), .B(n2931), .Z(n3060) );
  AND U3378 ( .A(\stack[1][7] ), .B(o[17]), .Z(n3059) );
  NAND U3379 ( .A(n3060), .B(n3059), .Z(n2933) );
  NAND U3380 ( .A(n2934), .B(n2933), .Z(n2937) );
  NAND U3381 ( .A(n2938), .B(n2937), .Z(n2940) );
  XOR U3382 ( .A(n2936), .B(n2935), .Z(n2958) );
  XOR U3383 ( .A(n2938), .B(n2937), .Z(n2957) );
  NAND U3384 ( .A(n2958), .B(n2957), .Z(n2939) );
  NAND U3385 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3386 ( .A(n2942), .B(n2941), .Z(n2944) );
  XOR U3387 ( .A(n2942), .B(n2941), .Z(n3070) );
  AND U3388 ( .A(\stack[1][7] ), .B(o[19]), .Z(n3069) );
  NAND U3389 ( .A(n3070), .B(n3069), .Z(n2943) );
  NAND U3390 ( .A(n2944), .B(n2943), .Z(n2947) );
  NAND U3391 ( .A(n2948), .B(n2947), .Z(n2950) );
  XOR U3392 ( .A(n2948), .B(n2947), .Z(n2955) );
  NAND U3393 ( .A(n2956), .B(n2955), .Z(n2949) );
  NAND U3394 ( .A(n2950), .B(n2949), .Z(n2951) );
  NAND U3395 ( .A(n2952), .B(n2951), .Z(n2954) );
  XOR U3396 ( .A(n2952), .B(n2951), .Z(n3080) );
  AND U3397 ( .A(\stack[1][7] ), .B(o[21]), .Z(n3079) );
  NAND U3398 ( .A(n3080), .B(n3079), .Z(n2953) );
  NAND U3399 ( .A(n2954), .B(n2953), .Z(n3211) );
  XOR U3400 ( .A(n3212), .B(n3211), .Z(n3213) );
  XOR U3401 ( .A(n3214), .B(n3213), .Z(n3083) );
  AND U3402 ( .A(\stack[1][6] ), .B(o[22]), .Z(n3077) );
  XOR U3403 ( .A(n2956), .B(n2955), .Z(n3073) );
  AND U3404 ( .A(\stack[1][6] ), .B(o[20]), .Z(n3067) );
  XOR U3405 ( .A(n2958), .B(n2957), .Z(n3063) );
  AND U3406 ( .A(\stack[1][6] ), .B(o[18]), .Z(n3056) );
  XNOR U3407 ( .A(n2960), .B(n2959), .Z(n3052) );
  NAND U3408 ( .A(\stack[1][6] ), .B(o[12]), .Z(n3022) );
  AND U3409 ( .A(o[10]), .B(\stack[1][6] ), .Z(n3012) );
  XNOR U3410 ( .A(n2962), .B(n2961), .Z(n3006) );
  XNOR U3411 ( .A(n2964), .B(n2963), .Z(n2985) );
  AND U3412 ( .A(\stack[1][6] ), .B(o[5]), .Z(n2986) );
  NAND U3413 ( .A(n2985), .B(n2986), .Z(n2988) );
  AND U3414 ( .A(o[0]), .B(\stack[1][6] ), .Z(n2965) );
  AND U3415 ( .A(o[1]), .B(\stack[1][7] ), .Z(n2970) );
  AND U3416 ( .A(n2965), .B(n2970), .Z(n2966) );
  NAND U3417 ( .A(o[2]), .B(n2966), .Z(n2972) );
  NAND U3418 ( .A(n2970), .B(o[0]), .Z(n2967) );
  XNOR U3419 ( .A(o[2]), .B(n2967), .Z(n2968) );
  AND U3420 ( .A(\stack[1][6] ), .B(n2968), .Z(n3231) );
  NAND U3421 ( .A(\stack[1][8] ), .B(o[0]), .Z(n2969) );
  XNOR U3422 ( .A(n2970), .B(n2969), .Z(n3232) );
  NAND U3423 ( .A(n3231), .B(n3232), .Z(n2971) );
  NAND U3424 ( .A(n2972), .B(n2971), .Z(n2975) );
  NAND U3425 ( .A(n2975), .B(n2976), .Z(n2978) );
  AND U3426 ( .A(\stack[1][6] ), .B(o[3]), .Z(n3239) );
  NAND U3427 ( .A(n3239), .B(n3240), .Z(n2977) );
  NAND U3428 ( .A(n2978), .B(n2977), .Z(n2981) );
  AND U3429 ( .A(\stack[1][6] ), .B(o[4]), .Z(n2982) );
  NAND U3430 ( .A(n2981), .B(n2982), .Z(n2984) );
  XOR U3431 ( .A(n2980), .B(n2979), .Z(n3244) );
  NAND U3432 ( .A(n3244), .B(n3243), .Z(n2983) );
  NAND U3433 ( .A(n2984), .B(n2983), .Z(n3249) );
  NAND U3434 ( .A(n3249), .B(n3250), .Z(n2987) );
  NAND U3435 ( .A(n2988), .B(n2987), .Z(n2991) );
  NAND U3436 ( .A(n2991), .B(n2992), .Z(n2994) );
  AND U3437 ( .A(\stack[1][6] ), .B(o[6]), .Z(n5395) );
  NAND U3438 ( .A(n5395), .B(n3255), .Z(n2993) );
  NAND U3439 ( .A(n2994), .B(n2993), .Z(n2997) );
  XOR U3440 ( .A(n2996), .B(n2995), .Z(n2998) );
  NAND U3441 ( .A(n2997), .B(n2998), .Z(n3000) );
  AND U3442 ( .A(\stack[1][6] ), .B(o[7]), .Z(n3261) );
  NAND U3443 ( .A(n3261), .B(n3260), .Z(n2999) );
  NAND U3444 ( .A(n3000), .B(n2999), .Z(n3001) );
  AND U3445 ( .A(\stack[1][6] ), .B(o[8]), .Z(n3002) );
  NAND U3446 ( .A(n3001), .B(n3002), .Z(n3005) );
  XOR U3447 ( .A(n5354), .B(n3003), .Z(n3266) );
  NAND U3448 ( .A(n3267), .B(n3266), .Z(n3004) );
  AND U3449 ( .A(n3005), .B(n3004), .Z(n3007) );
  NAND U3450 ( .A(n3006), .B(n3007), .Z(n3009) );
  NAND U3451 ( .A(\stack[1][6] ), .B(o[9]), .Z(n3272) );
  NAND U3452 ( .A(n3273), .B(n3272), .Z(n3008) );
  AND U3453 ( .A(n3009), .B(n3008), .Z(n3013) );
  NAND U3454 ( .A(n3012), .B(n3013), .Z(n3015) );
  NAND U3455 ( .A(n3222), .B(n3221), .Z(n3014) );
  NAND U3456 ( .A(n3015), .B(n3014), .Z(n3018) );
  NAND U3457 ( .A(n3018), .B(n3019), .Z(n3021) );
  AND U3458 ( .A(\stack[1][6] ), .B(o[11]), .Z(n3282) );
  NAND U3459 ( .A(n3282), .B(n3283), .Z(n3020) );
  AND U3460 ( .A(n3021), .B(n3020), .Z(n3023) );
  NAND U3461 ( .A(n3022), .B(n3023), .Z(n3027) );
  NAND U3462 ( .A(n3289), .B(n3288), .Z(n3026) );
  AND U3463 ( .A(n3027), .B(n3026), .Z(n3031) );
  XOR U3464 ( .A(n3029), .B(n3028), .Z(n3030) );
  NAND U3465 ( .A(n3031), .B(n3030), .Z(n3033) );
  AND U3466 ( .A(\stack[1][6] ), .B(o[13]), .Z(n3294) );
  XOR U3467 ( .A(n3031), .B(n3030), .Z(n3295) );
  NAND U3468 ( .A(n3294), .B(n3295), .Z(n3032) );
  NAND U3469 ( .A(n3033), .B(n3032), .Z(n3036) );
  AND U3470 ( .A(\stack[1][6] ), .B(o[14]), .Z(n3037) );
  NAND U3471 ( .A(n3036), .B(n3037), .Z(n3039) );
  NAND U3472 ( .A(n3301), .B(n3300), .Z(n3038) );
  NAND U3473 ( .A(n3039), .B(n3038), .Z(n3042) );
  NAND U3474 ( .A(n3042), .B(n3043), .Z(n3045) );
  AND U3475 ( .A(\stack[1][6] ), .B(o[15]), .Z(n3307) );
  NAND U3476 ( .A(n3307), .B(n3306), .Z(n3044) );
  NAND U3477 ( .A(n3045), .B(n3044), .Z(n3046) );
  AND U3478 ( .A(\stack[1][6] ), .B(o[16]), .Z(n3047) );
  NAND U3479 ( .A(n3046), .B(n3047), .Z(n3051) );
  XOR U3480 ( .A(n3049), .B(n3048), .Z(n3312) );
  NAND U3481 ( .A(n3313), .B(n3312), .Z(n3050) );
  AND U3482 ( .A(n3051), .B(n3050), .Z(n3053) );
  NAND U3483 ( .A(n3052), .B(n3053), .Z(n3055) );
  NAND U3484 ( .A(\stack[1][6] ), .B(o[17]), .Z(n3320) );
  NAND U3485 ( .A(n3320), .B(n3321), .Z(n3054) );
  AND U3486 ( .A(n3055), .B(n3054), .Z(n3058) );
  NAND U3487 ( .A(n3056), .B(n3058), .Z(n3062) );
  IV U3488 ( .A(n3056), .Z(n3057) );
  XNOR U3489 ( .A(n3058), .B(n3057), .Z(n3325) );
  XOR U3490 ( .A(n3060), .B(n3059), .Z(n3324) );
  NAND U3491 ( .A(n3325), .B(n3324), .Z(n3061) );
  NAND U3492 ( .A(n3062), .B(n3061), .Z(n3064) );
  NAND U3493 ( .A(n3063), .B(n3064), .Z(n3066) );
  XOR U3494 ( .A(n3064), .B(n3063), .Z(n3331) );
  AND U3495 ( .A(\stack[1][6] ), .B(o[19]), .Z(n3330) );
  NAND U3496 ( .A(n3331), .B(n3330), .Z(n3065) );
  NAND U3497 ( .A(n3066), .B(n3065), .Z(n3068) );
  NAND U3498 ( .A(n3067), .B(n3068), .Z(n3072) );
  XOR U3499 ( .A(n3068), .B(n3067), .Z(n3219) );
  XOR U3500 ( .A(n3070), .B(n3069), .Z(n3220) );
  NAND U3501 ( .A(n3219), .B(n3220), .Z(n3071) );
  NAND U3502 ( .A(n3072), .B(n3071), .Z(n3074) );
  NAND U3503 ( .A(n3073), .B(n3074), .Z(n3076) );
  XOR U3504 ( .A(n3074), .B(n3073), .Z(n3341) );
  AND U3505 ( .A(\stack[1][6] ), .B(o[21]), .Z(n3340) );
  NAND U3506 ( .A(n3341), .B(n3340), .Z(n3075) );
  NAND U3507 ( .A(n3076), .B(n3075), .Z(n3078) );
  NAND U3508 ( .A(n3077), .B(n3078), .Z(n3082) );
  XOR U3509 ( .A(n3078), .B(n3077), .Z(n3218) );
  XOR U3510 ( .A(n3080), .B(n3079), .Z(n3217) );
  NAND U3511 ( .A(n3218), .B(n3217), .Z(n3081) );
  NAND U3512 ( .A(n3082), .B(n3081), .Z(n3084) );
  NAND U3513 ( .A(n3083), .B(n3084), .Z(n3086) );
  XOR U3514 ( .A(n3084), .B(n3083), .Z(n3350) );
  AND U3515 ( .A(\stack[1][6] ), .B(o[23]), .Z(n3351) );
  NAND U3516 ( .A(n3350), .B(n3351), .Z(n3085) );
  NAND U3517 ( .A(n3086), .B(n3085), .Z(n3362) );
  AND U3518 ( .A(\stack[1][6] ), .B(o[24]), .Z(n3363) );
  XOR U3519 ( .A(n3362), .B(n3363), .Z(n3361) );
  NAND U3520 ( .A(n3088), .B(n3087), .Z(n3092) );
  NAND U3521 ( .A(n3090), .B(n3089), .Z(n3091) );
  NAND U3522 ( .A(n3092), .B(n3091), .Z(n3596) );
  AND U3523 ( .A(\stack[1][8] ), .B(o[22]), .Z(n3597) );
  XOR U3524 ( .A(n3596), .B(n3597), .Z(n3595) );
  NAND U3525 ( .A(n3094), .B(n3093), .Z(n3098) );
  NAND U3526 ( .A(n3096), .B(n3095), .Z(n3097) );
  NAND U3527 ( .A(n3098), .B(n3097), .Z(n3368) );
  AND U3528 ( .A(\stack[1][10] ), .B(o[20]), .Z(n3369) );
  XOR U3529 ( .A(n3368), .B(n3369), .Z(n3367) );
  NAND U3530 ( .A(n3100), .B(n3099), .Z(n3104) );
  NAND U3531 ( .A(n3102), .B(n3101), .Z(n3103) );
  NAND U3532 ( .A(n3104), .B(n3103), .Z(n3375) );
  NAND U3533 ( .A(n3106), .B(n3105), .Z(n3110) );
  NAND U3534 ( .A(n3108), .B(n3107), .Z(n3109) );
  AND U3535 ( .A(n3110), .B(n3109), .Z(n3561) );
  NAND U3536 ( .A(\stack[1][14] ), .B(o[16]), .Z(n3560) );
  XOR U3537 ( .A(n3561), .B(n3560), .Z(n3559) );
  AND U3538 ( .A(\stack[1][15] ), .B(o[15]), .Z(n5047) );
  NAND U3539 ( .A(n3112), .B(n3111), .Z(n3116) );
  NAND U3540 ( .A(n3114), .B(n3113), .Z(n3115) );
  NAND U3541 ( .A(n3116), .B(n3115), .Z(n3381) );
  NAND U3542 ( .A(n3118), .B(n3117), .Z(n3122) );
  NAND U3543 ( .A(n3120), .B(n3119), .Z(n3121) );
  AND U3544 ( .A(n3122), .B(n3121), .Z(n3387) );
  NAND U3545 ( .A(o[12]), .B(\stack[1][18] ), .Z(n3386) );
  XOR U3546 ( .A(n3387), .B(n3386), .Z(n3385) );
  NAND U3547 ( .A(n3124), .B(n3123), .Z(n3128) );
  NAND U3548 ( .A(n3126), .B(n3125), .Z(n3127) );
  NAND U3549 ( .A(n3128), .B(n3127), .Z(n3392) );
  AND U3550 ( .A(o[8]), .B(\stack[1][22] ), .Z(n3393) );
  XOR U3551 ( .A(n3392), .B(n3393), .Z(n3391) );
  AND U3552 ( .A(o[6]), .B(\stack[1][24] ), .Z(n3482) );
  NAND U3553 ( .A(n3130), .B(n3129), .Z(n3134) );
  NAND U3554 ( .A(n3132), .B(n3131), .Z(n3133) );
  NAND U3555 ( .A(n3134), .B(n3133), .Z(n3489) );
  AND U3556 ( .A(o[0]), .B(\stack[1][27] ), .Z(n3136) );
  AND U3557 ( .A(n3136), .B(n3135), .Z(n3137) );
  NAND U3558 ( .A(o[2]), .B(n3137), .Z(n3141) );
  NAND U3559 ( .A(n3139), .B(n3138), .Z(n3140) );
  NAND U3560 ( .A(n3141), .B(n3140), .Z(n3404) );
  AND U3561 ( .A(o[3]), .B(\stack[1][27] ), .Z(n3405) );
  XOR U3562 ( .A(n3404), .B(n3405), .Z(n3403) );
  AND U3563 ( .A(o[1]), .B(\stack[1][29] ), .Z(n3424) );
  NAND U3564 ( .A(\stack[1][30] ), .B(o[0]), .Z(n3142) );
  XNOR U3565 ( .A(n3424), .B(n3142), .Z(n3423) );
  NAND U3566 ( .A(n3424), .B(o[0]), .Z(n3143) );
  XNOR U3567 ( .A(o[2]), .B(n3143), .Z(n3144) );
  AND U3568 ( .A(\stack[1][28] ), .B(n3144), .Z(n3422) );
  XOR U3569 ( .A(n3423), .B(n3422), .Z(n3402) );
  XOR U3570 ( .A(n3403), .B(n3402), .Z(n3396) );
  NAND U3571 ( .A(n3146), .B(n3145), .Z(n3150) );
  NAND U3572 ( .A(n3148), .B(n3147), .Z(n3149) );
  NAND U3573 ( .A(n3150), .B(n3149), .Z(n3398) );
  AND U3574 ( .A(o[4]), .B(\stack[1][26] ), .Z(n3399) );
  XOR U3575 ( .A(n3398), .B(n3399), .Z(n3397) );
  XOR U3576 ( .A(n3489), .B(n3490), .Z(n3488) );
  AND U3577 ( .A(o[5]), .B(\stack[1][25] ), .Z(n3487) );
  XOR U3578 ( .A(n3488), .B(n3487), .Z(n3484) );
  NAND U3579 ( .A(n3152), .B(n3151), .Z(n3156) );
  NAND U3580 ( .A(n3154), .B(n3153), .Z(n3155) );
  NAND U3581 ( .A(n3156), .B(n3155), .Z(n3483) );
  XOR U3582 ( .A(n3484), .B(n3483), .Z(n3481) );
  XOR U3583 ( .A(n3482), .B(n3481), .Z(n3508) );
  NAND U3584 ( .A(n3158), .B(n3157), .Z(n3162) );
  NAND U3585 ( .A(n3160), .B(n3159), .Z(n3161) );
  NAND U3586 ( .A(n3162), .B(n3161), .Z(n3507) );
  XOR U3587 ( .A(n3508), .B(n3507), .Z(n3506) );
  AND U3588 ( .A(o[7]), .B(\stack[1][23] ), .Z(n3505) );
  XOR U3589 ( .A(n3506), .B(n3505), .Z(n3390) );
  XOR U3590 ( .A(n3391), .B(n3390), .Z(n3502) );
  NAND U3591 ( .A(n3164), .B(n3163), .Z(n3168) );
  NAND U3592 ( .A(n3166), .B(n3165), .Z(n3167) );
  NAND U3593 ( .A(n3168), .B(n3167), .Z(n3501) );
  XOR U3594 ( .A(n3502), .B(n3501), .Z(n3500) );
  AND U3595 ( .A(o[9]), .B(\stack[1][21] ), .Z(n3499) );
  XOR U3596 ( .A(n3500), .B(n3499), .Z(n3526) );
  AND U3597 ( .A(o[10]), .B(\stack[1][20] ), .Z(n3524) );
  NAND U3598 ( .A(n3170), .B(n3169), .Z(n3174) );
  NAND U3599 ( .A(n3172), .B(n3171), .Z(n3173) );
  AND U3600 ( .A(n3174), .B(n3173), .Z(n3523) );
  XOR U3601 ( .A(n3524), .B(n3523), .Z(n3525) );
  XNOR U3602 ( .A(n3526), .B(n3525), .Z(n3519) );
  NAND U3603 ( .A(n3176), .B(n3175), .Z(n3180) );
  NAND U3604 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3605 ( .A(n3180), .B(n3179), .Z(n3520) );
  NAND U3606 ( .A(o[11]), .B(\stack[1][19] ), .Z(n3517) );
  XOR U3607 ( .A(n3518), .B(n3517), .Z(n3384) );
  XNOR U3608 ( .A(n3385), .B(n3384), .Z(n3380) );
  XOR U3609 ( .A(n3381), .B(n3380), .Z(n3379) );
  AND U3610 ( .A(o[13]), .B(\stack[1][17] ), .Z(n3378) );
  XOR U3611 ( .A(n3379), .B(n3378), .Z(n3541) );
  NAND U3612 ( .A(n3182), .B(n3181), .Z(n3186) );
  NAND U3613 ( .A(n3184), .B(n3183), .Z(n3185) );
  AND U3614 ( .A(n3186), .B(n3185), .Z(n3543) );
  AND U3615 ( .A(o[14]), .B(\stack[1][16] ), .Z(n3542) );
  XOR U3616 ( .A(n3543), .B(n3542), .Z(n3540) );
  XOR U3617 ( .A(n3541), .B(n3540), .Z(n3537) );
  NAND U3618 ( .A(n3188), .B(n3187), .Z(n3192) );
  NAND U3619 ( .A(n3190), .B(n3189), .Z(n3191) );
  NAND U3620 ( .A(n3192), .B(n3191), .Z(n3536) );
  XOR U3621 ( .A(n3537), .B(n3536), .Z(n3535) );
  XNOR U3622 ( .A(n5047), .B(n3535), .Z(n3558) );
  XNOR U3623 ( .A(n3559), .B(n3558), .Z(n3374) );
  XOR U3624 ( .A(n3375), .B(n3374), .Z(n3373) );
  AND U3625 ( .A(\stack[1][13] ), .B(o[17]), .Z(n3372) );
  XNOR U3626 ( .A(n3373), .B(n3372), .Z(n3553) );
  NAND U3627 ( .A(n3194), .B(n3193), .Z(n3198) );
  NAND U3628 ( .A(n3196), .B(n3195), .Z(n3197) );
  AND U3629 ( .A(n3198), .B(n3197), .Z(n3555) );
  NAND U3630 ( .A(\stack[1][12] ), .B(o[18]), .Z(n3554) );
  XOR U3631 ( .A(n3555), .B(n3554), .Z(n3552) );
  NAND U3632 ( .A(n3200), .B(n3199), .Z(n3204) );
  NAND U3633 ( .A(n3202), .B(n3201), .Z(n3203) );
  NAND U3634 ( .A(n3204), .B(n3203), .Z(n3578) );
  AND U3635 ( .A(\stack[1][11] ), .B(o[19]), .Z(n3576) );
  XOR U3636 ( .A(n3577), .B(n3576), .Z(n3366) );
  XOR U3637 ( .A(n3367), .B(n3366), .Z(n3573) );
  NAND U3638 ( .A(n3206), .B(n3205), .Z(n3210) );
  NAND U3639 ( .A(n3208), .B(n3207), .Z(n3209) );
  NAND U3640 ( .A(n3210), .B(n3209), .Z(n3572) );
  XOR U3641 ( .A(n3573), .B(n3572), .Z(n3571) );
  AND U3642 ( .A(\stack[1][9] ), .B(o[21]), .Z(n3570) );
  XOR U3643 ( .A(n3571), .B(n3570), .Z(n3594) );
  XOR U3644 ( .A(n3595), .B(n3594), .Z(n3591) );
  NAND U3645 ( .A(n3212), .B(n3211), .Z(n3216) );
  NAND U3646 ( .A(n3214), .B(n3213), .Z(n3215) );
  NAND U3647 ( .A(n3216), .B(n3215), .Z(n3590) );
  XOR U3648 ( .A(n3591), .B(n3590), .Z(n3589) );
  AND U3649 ( .A(\stack[1][7] ), .B(o[23]), .Z(n3588) );
  XOR U3650 ( .A(n3589), .B(n3588), .Z(n3360) );
  XOR U3651 ( .A(n3361), .B(n3360), .Z(n3357) );
  AND U3652 ( .A(\stack[1][5] ), .B(o[24]), .Z(n3353) );
  XOR U3653 ( .A(n3218), .B(n3217), .Z(n3347) );
  AND U3654 ( .A(\stack[1][5] ), .B(o[22]), .Z(n3343) );
  AND U3655 ( .A(\stack[1][5] ), .B(o[20]), .Z(n3333) );
  XNOR U3656 ( .A(n3222), .B(n3221), .Z(n3278) );
  AND U3657 ( .A(o[0]), .B(\stack[1][5] ), .Z(n3223) );
  AND U3658 ( .A(o[1]), .B(\stack[1][6] ), .Z(n3228) );
  AND U3659 ( .A(n3223), .B(n3228), .Z(n3224) );
  NAND U3660 ( .A(n3224), .B(o[2]), .Z(n3230) );
  NAND U3661 ( .A(n3228), .B(o[0]), .Z(n3225) );
  XNOR U3662 ( .A(o[2]), .B(n3225), .Z(n3226) );
  AND U3663 ( .A(\stack[1][5] ), .B(n3226), .Z(n3622) );
  NAND U3664 ( .A(\stack[1][7] ), .B(o[0]), .Z(n3227) );
  XNOR U3665 ( .A(n3228), .B(n3227), .Z(n3623) );
  NAND U3666 ( .A(n3622), .B(n3623), .Z(n3229) );
  NAND U3667 ( .A(n3230), .B(n3229), .Z(n3233) );
  NAND U3668 ( .A(n3233), .B(n3234), .Z(n3236) );
  AND U3669 ( .A(\stack[1][5] ), .B(o[3]), .Z(n3629) );
  NAND U3670 ( .A(n3629), .B(n3628), .Z(n3235) );
  NAND U3671 ( .A(n3236), .B(n3235), .Z(n3237) );
  AND U3672 ( .A(\stack[1][5] ), .B(o[4]), .Z(n3238) );
  NAND U3673 ( .A(n3237), .B(n3238), .Z(n3242) );
  NAND U3674 ( .A(n3613), .B(n3612), .Z(n3241) );
  NAND U3675 ( .A(n3242), .B(n3241), .Z(n3245) );
  XOR U3676 ( .A(n3244), .B(n3243), .Z(n3246) );
  NAND U3677 ( .A(n3245), .B(n3246), .Z(n3248) );
  AND U3678 ( .A(\stack[1][5] ), .B(o[5]), .Z(n3639) );
  NAND U3679 ( .A(n3639), .B(n3638), .Z(n3247) );
  NAND U3680 ( .A(n3248), .B(n3247), .Z(n3251) );
  NAND U3681 ( .A(n3251), .B(n3252), .Z(n3254) );
  AND U3682 ( .A(\stack[1][5] ), .B(o[6]), .Z(n3645) );
  NAND U3683 ( .A(n3645), .B(n3644), .Z(n3253) );
  NAND U3684 ( .A(n3254), .B(n3253), .Z(n3256) );
  XOR U3685 ( .A(n5395), .B(n3255), .Z(n3257) );
  NAND U3686 ( .A(n3256), .B(n3257), .Z(n3259) );
  AND U3687 ( .A(\stack[1][5] ), .B(o[7]), .Z(n3652) );
  NAND U3688 ( .A(n3652), .B(n3653), .Z(n3258) );
  NAND U3689 ( .A(n3259), .B(n3258), .Z(n3262) );
  AND U3690 ( .A(\stack[1][5] ), .B(o[8]), .Z(n3263) );
  NAND U3691 ( .A(n3262), .B(n3263), .Z(n3265) );
  XOR U3692 ( .A(n3261), .B(n3260), .Z(n3611) );
  NAND U3693 ( .A(n3611), .B(n3610), .Z(n3264) );
  NAND U3694 ( .A(n3265), .B(n3264), .Z(n3268) );
  XOR U3695 ( .A(n3267), .B(n3266), .Z(n3269) );
  NAND U3696 ( .A(n3268), .B(n3269), .Z(n3271) );
  AND U3697 ( .A(\stack[1][5] ), .B(o[9]), .Z(n3660) );
  NAND U3698 ( .A(n3660), .B(n3661), .Z(n3270) );
  NAND U3699 ( .A(n3271), .B(n3270), .Z(n3274) );
  AND U3700 ( .A(o[10]), .B(\stack[1][5] ), .Z(n3275) );
  NAND U3701 ( .A(n3274), .B(n3275), .Z(n3277) );
  XNOR U3702 ( .A(n3273), .B(n3272), .Z(n3666) );
  NAND U3703 ( .A(n3666), .B(n3667), .Z(n3276) );
  AND U3704 ( .A(n3277), .B(n3276), .Z(n3279) );
  NAND U3705 ( .A(n3278), .B(n3279), .Z(n3281) );
  NAND U3706 ( .A(\stack[1][5] ), .B(o[11]), .Z(n3674) );
  NAND U3707 ( .A(n3674), .B(n3675), .Z(n3280) );
  AND U3708 ( .A(n3281), .B(n3280), .Z(n3284) );
  AND U3709 ( .A(\stack[1][5] ), .B(o[12]), .Z(n3285) );
  NAND U3710 ( .A(n3284), .B(n3285), .Z(n3287) );
  NAND U3711 ( .A(n3679), .B(n3678), .Z(n3286) );
  NAND U3712 ( .A(n3287), .B(n3286), .Z(n3290) );
  XNOR U3713 ( .A(n3289), .B(n3288), .Z(n3291) );
  NAND U3714 ( .A(n3290), .B(n3291), .Z(n3293) );
  AND U3715 ( .A(\stack[1][5] ), .B(o[13]), .Z(n3686) );
  NAND U3716 ( .A(n3687), .B(n3686), .Z(n3292) );
  NAND U3717 ( .A(n3293), .B(n3292), .Z(n3296) );
  AND U3718 ( .A(\stack[1][5] ), .B(o[14]), .Z(n3297) );
  NAND U3719 ( .A(n3296), .B(n3297), .Z(n3299) );
  NAND U3720 ( .A(n3691), .B(n3690), .Z(n3298) );
  NAND U3721 ( .A(n3299), .B(n3298), .Z(n3302) );
  XOR U3722 ( .A(n3301), .B(n3300), .Z(n3303) );
  NAND U3723 ( .A(n3302), .B(n3303), .Z(n3305) );
  AND U3724 ( .A(\stack[1][5] ), .B(o[15]), .Z(n3696) );
  NAND U3725 ( .A(n3696), .B(n3697), .Z(n3304) );
  NAND U3726 ( .A(n3305), .B(n3304), .Z(n3308) );
  AND U3727 ( .A(\stack[1][5] ), .B(o[16]), .Z(n3309) );
  NAND U3728 ( .A(n3308), .B(n3309), .Z(n3311) );
  XOR U3729 ( .A(n3307), .B(n3306), .Z(n3703) );
  NAND U3730 ( .A(n3703), .B(n3702), .Z(n3310) );
  NAND U3731 ( .A(n3311), .B(n3310), .Z(n3314) );
  XOR U3732 ( .A(n3313), .B(n3312), .Z(n3315) );
  NAND U3733 ( .A(n3314), .B(n3315), .Z(n3317) );
  AND U3734 ( .A(\stack[1][5] ), .B(o[17]), .Z(n3708) );
  NAND U3735 ( .A(n3709), .B(n3708), .Z(n3316) );
  NAND U3736 ( .A(n3317), .B(n3316), .Z(n3318) );
  AND U3737 ( .A(\stack[1][5] ), .B(o[18]), .Z(n3319) );
  NAND U3738 ( .A(n3318), .B(n3319), .Z(n3323) );
  NAND U3739 ( .A(n3714), .B(n3715), .Z(n3322) );
  NAND U3740 ( .A(n3323), .B(n3322), .Z(n3326) );
  XOR U3741 ( .A(n3325), .B(n3324), .Z(n3327) );
  NAND U3742 ( .A(n3326), .B(n3327), .Z(n3329) );
  AND U3743 ( .A(\stack[1][5] ), .B(o[19]), .Z(n3722) );
  NAND U3744 ( .A(n3722), .B(n3724), .Z(n3328) );
  NAND U3745 ( .A(n3329), .B(n3328), .Z(n3332) );
  NAND U3746 ( .A(n3333), .B(n3332), .Z(n3335) );
  XOR U3747 ( .A(n3331), .B(n3330), .Z(n3728) );
  XOR U3748 ( .A(n3333), .B(n3332), .Z(n3727) );
  NAND U3749 ( .A(n3728), .B(n3727), .Z(n3334) );
  NAND U3750 ( .A(n3335), .B(n3334), .Z(n3336) );
  NAND U3751 ( .A(n3337), .B(n3336), .Z(n3339) );
  XOR U3752 ( .A(n3337), .B(n3336), .Z(n3736) );
  AND U3753 ( .A(\stack[1][5] ), .B(o[21]), .Z(n3735) );
  NAND U3754 ( .A(n3736), .B(n3735), .Z(n3338) );
  NAND U3755 ( .A(n3339), .B(n3338), .Z(n3342) );
  NAND U3756 ( .A(n3343), .B(n3342), .Z(n3345) );
  XOR U3757 ( .A(n3341), .B(n3340), .Z(n3740) );
  XOR U3758 ( .A(n3343), .B(n3342), .Z(n3739) );
  NAND U3759 ( .A(n3740), .B(n3739), .Z(n3344) );
  NAND U3760 ( .A(n3345), .B(n3344), .Z(n3346) );
  NAND U3761 ( .A(n3347), .B(n3346), .Z(n3349) );
  XOR U3762 ( .A(n3347), .B(n3346), .Z(n3746) );
  AND U3763 ( .A(\stack[1][5] ), .B(o[23]), .Z(n3745) );
  NAND U3764 ( .A(n3746), .B(n3745), .Z(n3348) );
  NAND U3765 ( .A(n3349), .B(n3348), .Z(n3352) );
  NAND U3766 ( .A(n3353), .B(n3352), .Z(n3355) );
  XOR U3767 ( .A(n3353), .B(n3352), .Z(n3608) );
  NAND U3768 ( .A(n3609), .B(n3608), .Z(n3354) );
  NAND U3769 ( .A(n3355), .B(n3354), .Z(n3356) );
  XOR U3770 ( .A(n3357), .B(n3356), .Z(n3607) );
  AND U3771 ( .A(\stack[1][5] ), .B(o[25]), .Z(n3606) );
  NAND U3772 ( .A(n3607), .B(n3606), .Z(n3359) );
  NAND U3773 ( .A(n3357), .B(n3356), .Z(n3358) );
  AND U3774 ( .A(n3359), .B(n3358), .Z(n4430) );
  NAND U3775 ( .A(n3361), .B(n3360), .Z(n3365) );
  NAND U3776 ( .A(n3363), .B(n3362), .Z(n3364) );
  AND U3777 ( .A(n3365), .B(n3364), .Z(n3921) );
  NAND U3778 ( .A(n3367), .B(n3366), .Z(n3371) );
  NAND U3779 ( .A(n3369), .B(n3368), .Z(n3370) );
  AND U3780 ( .A(n3371), .B(n3370), .Z(n3605) );
  NAND U3781 ( .A(n3373), .B(n3372), .Z(n3377) );
  NAND U3782 ( .A(n3375), .B(n3374), .Z(n3376) );
  AND U3783 ( .A(n3377), .B(n3376), .Z(n3587) );
  NAND U3784 ( .A(n3379), .B(n3378), .Z(n3383) );
  NAND U3785 ( .A(n3381), .B(n3380), .Z(n3382) );
  AND U3786 ( .A(n3383), .B(n3382), .Z(n3569) );
  NAND U3787 ( .A(n3385), .B(n3384), .Z(n3389) );
  NAND U3788 ( .A(n3387), .B(n3386), .Z(n3388) );
  AND U3789 ( .A(n3389), .B(n3388), .Z(n3551) );
  NAND U3790 ( .A(n3391), .B(n3390), .Z(n3395) );
  NAND U3791 ( .A(n3393), .B(n3392), .Z(n3394) );
  AND U3792 ( .A(n3395), .B(n3394), .Z(n3534) );
  NAND U3793 ( .A(n3397), .B(n3396), .Z(n3401) );
  NAND U3794 ( .A(n3399), .B(n3398), .Z(n3400) );
  AND U3795 ( .A(n3401), .B(n3400), .Z(n3516) );
  NAND U3796 ( .A(n3403), .B(n3402), .Z(n3407) );
  NAND U3797 ( .A(n3405), .B(n3404), .Z(n3406) );
  AND U3798 ( .A(n3407), .B(n3406), .Z(n3498) );
  AND U3799 ( .A(o[28]), .B(\stack[1][3] ), .Z(n3409) );
  NAND U3800 ( .A(o[26]), .B(\stack[1][5] ), .Z(n3408) );
  XNOR U3801 ( .A(n3409), .B(n3408), .Z(n3413) );
  AND U3802 ( .A(o[30]), .B(\stack[1][1] ), .Z(n3411) );
  NAND U3803 ( .A(o[24]), .B(\stack[1][7] ), .Z(n3410) );
  XNOR U3804 ( .A(n3411), .B(n3410), .Z(n3412) );
  XOR U3805 ( .A(n3413), .B(n3412), .Z(n3421) );
  AND U3806 ( .A(o[16]), .B(\stack[1][15] ), .Z(n3415) );
  NAND U3807 ( .A(o[20]), .B(\stack[1][11] ), .Z(n3414) );
  XNOR U3808 ( .A(n3415), .B(n3414), .Z(n3419) );
  AND U3809 ( .A(o[15]), .B(\stack[1][16] ), .Z(n3417) );
  NAND U3810 ( .A(\stack[1][25] ), .B(o[6]), .Z(n3416) );
  XNOR U3811 ( .A(n3417), .B(n3416), .Z(n3418) );
  XNOR U3812 ( .A(n3419), .B(n3418), .Z(n3420) );
  XNOR U3813 ( .A(n3421), .B(n3420), .Z(n3462) );
  NAND U3814 ( .A(n3423), .B(n3422), .Z(n3428) );
  AND U3815 ( .A(o[0]), .B(\stack[1][28] ), .Z(n3425) );
  AND U3816 ( .A(n3425), .B(n3424), .Z(n3426) );
  NAND U3817 ( .A(o[2]), .B(n3426), .Z(n3427) );
  AND U3818 ( .A(n3428), .B(n3427), .Z(n3460) );
  AND U3819 ( .A(\stack[1][24] ), .B(o[7]), .Z(n3430) );
  NAND U3820 ( .A(\stack[1][27] ), .B(o[4]), .Z(n3429) );
  XNOR U3821 ( .A(n3430), .B(n3429), .Z(n3434) );
  AND U3822 ( .A(\stack[1][26] ), .B(o[5]), .Z(n3432) );
  NAND U3823 ( .A(\stack[1][28] ), .B(o[3]), .Z(n3431) );
  XNOR U3824 ( .A(n3432), .B(n3431), .Z(n3433) );
  XOR U3825 ( .A(n3434), .B(n3433), .Z(n3442) );
  AND U3826 ( .A(\stack[1][22] ), .B(o[9]), .Z(n3436) );
  NAND U3827 ( .A(o[0]), .B(\stack[1][31] ), .Z(n3435) );
  XNOR U3828 ( .A(n3436), .B(n3435), .Z(n3440) );
  AND U3829 ( .A(\stack[1][23] ), .B(o[8]), .Z(n3438) );
  NAND U3830 ( .A(\stack[1][21] ), .B(o[10]), .Z(n3437) );
  XNOR U3831 ( .A(n3438), .B(n3437), .Z(n3439) );
  XNOR U3832 ( .A(n3440), .B(n3439), .Z(n3441) );
  XNOR U3833 ( .A(n3442), .B(n3441), .Z(n3458) );
  AND U3834 ( .A(\stack[1][18] ), .B(o[13]), .Z(n3444) );
  NAND U3835 ( .A(\stack[1][20] ), .B(o[11]), .Z(n3443) );
  XNOR U3836 ( .A(n3444), .B(n3443), .Z(n3448) );
  AND U3837 ( .A(\stack[1][19] ), .B(o[12]), .Z(n3446) );
  NAND U3838 ( .A(o[18]), .B(\stack[1][13] ), .Z(n3445) );
  XNOR U3839 ( .A(n3446), .B(n3445), .Z(n3447) );
  XOR U3840 ( .A(n3448), .B(n3447), .Z(n3456) );
  AND U3841 ( .A(\stack[1][17] ), .B(o[14]), .Z(n3450) );
  NAND U3842 ( .A(o[17]), .B(\stack[1][14] ), .Z(n3449) );
  XNOR U3843 ( .A(n3450), .B(n3449), .Z(n3454) );
  AND U3844 ( .A(o[19]), .B(\stack[1][12] ), .Z(n3452) );
  NAND U3845 ( .A(o[22]), .B(\stack[1][9] ), .Z(n3451) );
  XNOR U3846 ( .A(n3452), .B(n3451), .Z(n3453) );
  XNOR U3847 ( .A(n3454), .B(n3453), .Z(n3455) );
  XNOR U3848 ( .A(n3456), .B(n3455), .Z(n3457) );
  XNOR U3849 ( .A(n3458), .B(n3457), .Z(n3459) );
  XNOR U3850 ( .A(n3460), .B(n3459), .Z(n3461) );
  XOR U3851 ( .A(n3462), .B(n3461), .Z(n3480) );
  AND U3852 ( .A(o[1]), .B(\stack[1][30] ), .Z(n3470) );
  NAND U3853 ( .A(n3470), .B(o[0]), .Z(n3463) );
  XNOR U3854 ( .A(o[2]), .B(n3463), .Z(n3464) );
  AND U3855 ( .A(\stack[1][29] ), .B(n3464), .Z(n3478) );
  AND U3856 ( .A(o[25]), .B(\stack[1][6] ), .Z(n3476) );
  AND U3857 ( .A(o[27]), .B(\stack[1][4] ), .Z(n3466) );
  NAND U3858 ( .A(o[29]), .B(\stack[1][2] ), .Z(n3465) );
  XNOR U3859 ( .A(n3466), .B(n3465), .Z(n3474) );
  AND U3860 ( .A(\stack[1][0] ), .B(o[31]), .Z(n3472) );
  AND U3861 ( .A(o[21]), .B(\stack[1][10] ), .Z(n3468) );
  NAND U3862 ( .A(o[23]), .B(\stack[1][8] ), .Z(n3467) );
  XNOR U3863 ( .A(n3468), .B(n3467), .Z(n3469) );
  XNOR U3864 ( .A(n3470), .B(n3469), .Z(n3471) );
  XNOR U3865 ( .A(n3472), .B(n3471), .Z(n3473) );
  XNOR U3866 ( .A(n3474), .B(n3473), .Z(n3475) );
  XNOR U3867 ( .A(n3476), .B(n3475), .Z(n3477) );
  XNOR U3868 ( .A(n3478), .B(n3477), .Z(n3479) );
  XNOR U3869 ( .A(n3480), .B(n3479), .Z(n3496) );
  NAND U3870 ( .A(n3482), .B(n3481), .Z(n3486) );
  NAND U3871 ( .A(n3484), .B(n3483), .Z(n3485) );
  AND U3872 ( .A(n3486), .B(n3485), .Z(n3494) );
  NAND U3873 ( .A(n3488), .B(n3487), .Z(n3492) );
  NAND U3874 ( .A(n3490), .B(n3489), .Z(n3491) );
  NAND U3875 ( .A(n3492), .B(n3491), .Z(n3493) );
  XNOR U3876 ( .A(n3494), .B(n3493), .Z(n3495) );
  XNOR U3877 ( .A(n3496), .B(n3495), .Z(n3497) );
  XNOR U3878 ( .A(n3498), .B(n3497), .Z(n3514) );
  NAND U3879 ( .A(n3500), .B(n3499), .Z(n3504) );
  NAND U3880 ( .A(n3502), .B(n3501), .Z(n3503) );
  AND U3881 ( .A(n3504), .B(n3503), .Z(n3512) );
  NAND U3882 ( .A(n3506), .B(n3505), .Z(n3510) );
  NAND U3883 ( .A(n3508), .B(n3507), .Z(n3509) );
  NAND U3884 ( .A(n3510), .B(n3509), .Z(n3511) );
  XNOR U3885 ( .A(n3512), .B(n3511), .Z(n3513) );
  XNOR U3886 ( .A(n3514), .B(n3513), .Z(n3515) );
  XNOR U3887 ( .A(n3516), .B(n3515), .Z(n3532) );
  NAND U3888 ( .A(n3518), .B(n3517), .Z(n3522) );
  AND U3889 ( .A(n3520), .B(n3519), .Z(n3521) );
  ANDN U3890 ( .B(n3522), .A(n3521), .Z(n3530) );
  AND U3891 ( .A(n3524), .B(n3523), .Z(n3528) );
  AND U3892 ( .A(n3526), .B(n3525), .Z(n3527) );
  OR U3893 ( .A(n3528), .B(n3527), .Z(n3529) );
  XNOR U3894 ( .A(n3530), .B(n3529), .Z(n3531) );
  XNOR U3895 ( .A(n3532), .B(n3531), .Z(n3533) );
  XNOR U3896 ( .A(n3534), .B(n3533), .Z(n3549) );
  NAND U3897 ( .A(n5047), .B(n3535), .Z(n3539) );
  NAND U3898 ( .A(n3537), .B(n3536), .Z(n3538) );
  AND U3899 ( .A(n3539), .B(n3538), .Z(n3547) );
  NAND U3900 ( .A(n3541), .B(n3540), .Z(n3545) );
  NAND U3901 ( .A(n3543), .B(n3542), .Z(n3544) );
  NAND U3902 ( .A(n3545), .B(n3544), .Z(n3546) );
  XNOR U3903 ( .A(n3547), .B(n3546), .Z(n3548) );
  XNOR U3904 ( .A(n3549), .B(n3548), .Z(n3550) );
  XNOR U3905 ( .A(n3551), .B(n3550), .Z(n3567) );
  NAND U3906 ( .A(n3553), .B(n3552), .Z(n3557) );
  NAND U3907 ( .A(n3555), .B(n3554), .Z(n3556) );
  AND U3908 ( .A(n3557), .B(n3556), .Z(n3565) );
  NAND U3909 ( .A(n3559), .B(n3558), .Z(n3563) );
  NAND U3910 ( .A(n3561), .B(n3560), .Z(n3562) );
  NAND U3911 ( .A(n3563), .B(n3562), .Z(n3564) );
  XNOR U3912 ( .A(n3565), .B(n3564), .Z(n3566) );
  XNOR U3913 ( .A(n3567), .B(n3566), .Z(n3568) );
  XNOR U3914 ( .A(n3569), .B(n3568), .Z(n3585) );
  NAND U3915 ( .A(n3571), .B(n3570), .Z(n3575) );
  NAND U3916 ( .A(n3573), .B(n3572), .Z(n3574) );
  AND U3917 ( .A(n3575), .B(n3574), .Z(n3583) );
  NAND U3918 ( .A(n3577), .B(n3576), .Z(n3581) );
  NAND U3919 ( .A(n3579), .B(n3578), .Z(n3580) );
  NAND U3920 ( .A(n3581), .B(n3580), .Z(n3582) );
  XNOR U3921 ( .A(n3583), .B(n3582), .Z(n3584) );
  XNOR U3922 ( .A(n3585), .B(n3584), .Z(n3586) );
  XNOR U3923 ( .A(n3587), .B(n3586), .Z(n3603) );
  NAND U3924 ( .A(n3589), .B(n3588), .Z(n3593) );
  NAND U3925 ( .A(n3591), .B(n3590), .Z(n3592) );
  AND U3926 ( .A(n3593), .B(n3592), .Z(n3601) );
  NAND U3927 ( .A(n3595), .B(n3594), .Z(n3599) );
  NAND U3928 ( .A(n3597), .B(n3596), .Z(n3598) );
  NAND U3929 ( .A(n3599), .B(n3598), .Z(n3600) );
  XNOR U3930 ( .A(n3601), .B(n3600), .Z(n3602) );
  XNOR U3931 ( .A(n3603), .B(n3602), .Z(n3604) );
  XNOR U3932 ( .A(n3605), .B(n3604), .Z(n3919) );
  XOR U3933 ( .A(n3607), .B(n3606), .Z(n3910) );
  XOR U3934 ( .A(n3609), .B(n3608), .Z(n3751) );
  NAND U3935 ( .A(\stack[1][4] ), .B(o[22]), .Z(n3733) );
  NAND U3936 ( .A(\stack[1][4] ), .B(o[18]), .Z(n3710) );
  NAND U3937 ( .A(\stack[1][4] ), .B(o[12]), .Z(n3672) );
  AND U3938 ( .A(o[10]), .B(\stack[1][4] ), .Z(n3662) );
  XNOR U3939 ( .A(n3611), .B(n3610), .Z(n3656) );
  AND U3940 ( .A(\stack[1][4] ), .B(o[5]), .Z(n3634) );
  XOR U3941 ( .A(n3613), .B(n3612), .Z(n3635) );
  NAND U3942 ( .A(n3634), .B(n3635), .Z(n3637) );
  AND U3943 ( .A(\stack[1][5] ), .B(o[1]), .Z(n3619) );
  AND U3944 ( .A(o[0]), .B(\stack[1][4] ), .Z(n3614) );
  AND U3945 ( .A(n3619), .B(n3614), .Z(n3615) );
  NAND U3946 ( .A(n3615), .B(o[2]), .Z(n3621) );
  NAND U3947 ( .A(n3619), .B(o[0]), .Z(n3616) );
  XNOR U3948 ( .A(o[2]), .B(n3616), .Z(n3617) );
  AND U3949 ( .A(\stack[1][4] ), .B(n3617), .Z(n3768) );
  NAND U3950 ( .A(\stack[1][6] ), .B(o[0]), .Z(n3618) );
  XNOR U3951 ( .A(n3619), .B(n3618), .Z(n3769) );
  NAND U3952 ( .A(n3768), .B(n3769), .Z(n3620) );
  NAND U3953 ( .A(n3621), .B(n3620), .Z(n3624) );
  NAND U3954 ( .A(n3624), .B(n3625), .Z(n3627) );
  AND U3955 ( .A(\stack[1][4] ), .B(o[3]), .Z(n3776) );
  NAND U3956 ( .A(n3776), .B(n3777), .Z(n3626) );
  NAND U3957 ( .A(n3627), .B(n3626), .Z(n3630) );
  AND U3958 ( .A(\stack[1][4] ), .B(o[4]), .Z(n3631) );
  NAND U3959 ( .A(n3630), .B(n3631), .Z(n3633) );
  XOR U3960 ( .A(n3629), .B(n3628), .Z(n3781) );
  NAND U3961 ( .A(n3781), .B(n3780), .Z(n3632) );
  NAND U3962 ( .A(n3633), .B(n3632), .Z(n3786) );
  NAND U3963 ( .A(n3786), .B(n3787), .Z(n3636) );
  NAND U3964 ( .A(n3637), .B(n3636), .Z(n3640) );
  XOR U3965 ( .A(n3639), .B(n3638), .Z(n3641) );
  NAND U3966 ( .A(n3640), .B(n3641), .Z(n3643) );
  AND U3967 ( .A(\stack[1][4] ), .B(o[6]), .Z(n3792) );
  NAND U3968 ( .A(n3792), .B(n3793), .Z(n3642) );
  NAND U3969 ( .A(n3643), .B(n3642), .Z(n3646) );
  XOR U3970 ( .A(n3645), .B(n3644), .Z(n3647) );
  NAND U3971 ( .A(n3646), .B(n3647), .Z(n3649) );
  AND U3972 ( .A(\stack[1][4] ), .B(o[7]), .Z(n3799) );
  NAND U3973 ( .A(n3799), .B(n3798), .Z(n3648) );
  NAND U3974 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U3975 ( .A(\stack[1][4] ), .B(o[8]), .Z(n3651) );
  NAND U3976 ( .A(n3650), .B(n3651), .Z(n3655) );
  NAND U3977 ( .A(n3805), .B(n3804), .Z(n3654) );
  AND U3978 ( .A(n3655), .B(n3654), .Z(n3657) );
  NAND U3979 ( .A(n3656), .B(n3657), .Z(n3659) );
  NAND U3980 ( .A(\stack[1][4] ), .B(o[9]), .Z(n3810) );
  NAND U3981 ( .A(n3811), .B(n3810), .Z(n3658) );
  AND U3982 ( .A(n3659), .B(n3658), .Z(n3663) );
  NAND U3983 ( .A(n3662), .B(n3663), .Z(n3665) );
  NAND U3984 ( .A(n3760), .B(n3759), .Z(n3664) );
  NAND U3985 ( .A(n3665), .B(n3664), .Z(n3668) );
  NAND U3986 ( .A(n3668), .B(n3669), .Z(n3671) );
  AND U3987 ( .A(\stack[1][4] ), .B(o[11]), .Z(n3820) );
  NAND U3988 ( .A(n3820), .B(n3821), .Z(n3670) );
  AND U3989 ( .A(n3671), .B(n3670), .Z(n3673) );
  NAND U3990 ( .A(n3672), .B(n3673), .Z(n3677) );
  NAND U3991 ( .A(n3758), .B(n3757), .Z(n3676) );
  NAND U3992 ( .A(n3677), .B(n3676), .Z(n3680) );
  XNOR U3993 ( .A(n3679), .B(n3678), .Z(n3681) );
  NAND U3994 ( .A(n3680), .B(n3681), .Z(n3683) );
  NAND U3995 ( .A(\stack[1][4] ), .B(o[13]), .Z(n3830) );
  NAND U3996 ( .A(n3831), .B(n3830), .Z(n3682) );
  NAND U3997 ( .A(n3683), .B(n3682), .Z(n3684) );
  NAND U3998 ( .A(\stack[1][4] ), .B(o[14]), .Z(n3685) );
  NAND U3999 ( .A(n3684), .B(n3685), .Z(n3689) );
  XNOR U4000 ( .A(n3687), .B(n3686), .Z(n3836) );
  NAND U4001 ( .A(n3837), .B(n3836), .Z(n3688) );
  AND U4002 ( .A(n3689), .B(n3688), .Z(n3693) );
  XOR U4003 ( .A(n3691), .B(n3690), .Z(n3692) );
  NAND U4004 ( .A(n3693), .B(n3692), .Z(n3695) );
  AND U4005 ( .A(\stack[1][4] ), .B(o[15]), .Z(n3843) );
  XOR U4006 ( .A(n3693), .B(n3692), .Z(n3842) );
  NAND U4007 ( .A(n3843), .B(n3842), .Z(n3694) );
  NAND U4008 ( .A(n3695), .B(n3694), .Z(n3698) );
  AND U4009 ( .A(\stack[1][4] ), .B(o[16]), .Z(n3699) );
  NAND U4010 ( .A(n3698), .B(n3699), .Z(n3701) );
  NAND U4011 ( .A(n3849), .B(n3848), .Z(n3700) );
  NAND U4012 ( .A(n3701), .B(n3700), .Z(n3704) );
  XOR U4013 ( .A(n3703), .B(n3702), .Z(n3705) );
  NAND U4014 ( .A(n3704), .B(n3705), .Z(n3707) );
  AND U4015 ( .A(\stack[1][4] ), .B(o[17]), .Z(n3855) );
  NAND U4016 ( .A(n3855), .B(n3854), .Z(n3706) );
  AND U4017 ( .A(n3707), .B(n3706), .Z(n3711) );
  NAND U4018 ( .A(n3710), .B(n3711), .Z(n3713) );
  XNOR U4019 ( .A(n3709), .B(n3708), .Z(n3755) );
  NAND U4020 ( .A(n3755), .B(n3756), .Z(n3712) );
  AND U4021 ( .A(n3713), .B(n3712), .Z(n3717) );
  XOR U4022 ( .A(n3715), .B(n3714), .Z(n3716) );
  NAND U4023 ( .A(n3717), .B(n3716), .Z(n3719) );
  AND U4024 ( .A(\stack[1][4] ), .B(o[19]), .Z(n3865) );
  XOR U4025 ( .A(n3717), .B(n3716), .Z(n3864) );
  NAND U4026 ( .A(n3865), .B(n3864), .Z(n3718) );
  NAND U4027 ( .A(n3719), .B(n3718), .Z(n3720) );
  AND U4028 ( .A(\stack[1][4] ), .B(o[20]), .Z(n3721) );
  NAND U4029 ( .A(n3720), .B(n3721), .Z(n3726) );
  IV U4030 ( .A(n3722), .Z(n3723) );
  XNOR U4031 ( .A(n3724), .B(n3723), .Z(n3870) );
  NAND U4032 ( .A(n3871), .B(n3870), .Z(n3725) );
  NAND U4033 ( .A(n3726), .B(n3725), .Z(n3729) );
  XOR U4034 ( .A(n3728), .B(n3727), .Z(n3730) );
  NAND U4035 ( .A(n3729), .B(n3730), .Z(n3732) );
  AND U4036 ( .A(\stack[1][4] ), .B(o[21]), .Z(n3876) );
  NAND U4037 ( .A(n3876), .B(n3877), .Z(n3731) );
  AND U4038 ( .A(n3732), .B(n3731), .Z(n3734) );
  NAND U4039 ( .A(n3733), .B(n3734), .Z(n3738) );
  XNOR U4040 ( .A(n3736), .B(n3735), .Z(n3882) );
  NAND U4041 ( .A(n3883), .B(n3882), .Z(n3737) );
  AND U4042 ( .A(n3738), .B(n3737), .Z(n3742) );
  XOR U4043 ( .A(n3740), .B(n3739), .Z(n3741) );
  NAND U4044 ( .A(n3742), .B(n3741), .Z(n3744) );
  AND U4045 ( .A(\stack[1][4] ), .B(o[23]), .Z(n3888) );
  XOR U4046 ( .A(n3742), .B(n3741), .Z(n3889) );
  NAND U4047 ( .A(n3888), .B(n3889), .Z(n3743) );
  NAND U4048 ( .A(n3744), .B(n3743), .Z(n3747) );
  AND U4049 ( .A(\stack[1][4] ), .B(o[24]), .Z(n3748) );
  NAND U4050 ( .A(n3747), .B(n3748), .Z(n3750) );
  XOR U4051 ( .A(n3746), .B(n3745), .Z(n3895) );
  NAND U4052 ( .A(n3895), .B(n3894), .Z(n3749) );
  NAND U4053 ( .A(n3750), .B(n3749), .Z(n3752) );
  NAND U4054 ( .A(n3751), .B(n3752), .Z(n3754) );
  XOR U4055 ( .A(n3752), .B(n3751), .Z(n3901) );
  AND U4056 ( .A(\stack[1][4] ), .B(o[25]), .Z(n3900) );
  NAND U4057 ( .A(n3901), .B(n3900), .Z(n3753) );
  NAND U4058 ( .A(n3754), .B(n3753), .Z(n3912) );
  AND U4059 ( .A(\stack[1][4] ), .B(o[26]), .Z(n3913) );
  XOR U4060 ( .A(n3912), .B(n3913), .Z(n3911) );
  AND U4061 ( .A(\stack[1][3] ), .B(o[26]), .Z(n3903) );
  XNOR U4062 ( .A(n3758), .B(n3757), .Z(n3826) );
  XNOR U4063 ( .A(n3760), .B(n3759), .Z(n3816) );
  AND U4064 ( .A(o[0]), .B(\stack[1][3] ), .Z(n4087) );
  AND U4065 ( .A(o[1]), .B(\stack[1][4] ), .Z(n3765) );
  AND U4066 ( .A(n4087), .B(n3765), .Z(n3761) );
  NAND U4067 ( .A(o[2]), .B(n3761), .Z(n3767) );
  NAND U4068 ( .A(n3765), .B(o[0]), .Z(n3762) );
  XNOR U4069 ( .A(o[2]), .B(n3762), .Z(n3763) );
  AND U4070 ( .A(\stack[1][3] ), .B(n3763), .Z(n3933) );
  NAND U4071 ( .A(\stack[1][5] ), .B(o[0]), .Z(n3764) );
  XNOR U4072 ( .A(n3765), .B(n3764), .Z(n3934) );
  NAND U4073 ( .A(n3933), .B(n3934), .Z(n3766) );
  NAND U4074 ( .A(n3767), .B(n3766), .Z(n3770) );
  NAND U4075 ( .A(n3770), .B(n3771), .Z(n3773) );
  AND U4076 ( .A(\stack[1][3] ), .B(o[3]), .Z(n3940) );
  NAND U4077 ( .A(n3940), .B(n3939), .Z(n3772) );
  NAND U4078 ( .A(n3773), .B(n3772), .Z(n3774) );
  AND U4079 ( .A(\stack[1][3] ), .B(o[4]), .Z(n3775) );
  NAND U4080 ( .A(n3774), .B(n3775), .Z(n3779) );
  NAND U4081 ( .A(n3925), .B(n3924), .Z(n3778) );
  NAND U4082 ( .A(n3779), .B(n3778), .Z(n3782) );
  XOR U4083 ( .A(n3781), .B(n3780), .Z(n3783) );
  NAND U4084 ( .A(n3782), .B(n3783), .Z(n3785) );
  AND U4085 ( .A(\stack[1][3] ), .B(o[5]), .Z(n3949) );
  NAND U4086 ( .A(n3949), .B(n3950), .Z(n3784) );
  NAND U4087 ( .A(n3785), .B(n3784), .Z(n3788) );
  NAND U4088 ( .A(n3788), .B(n3789), .Z(n3791) );
  AND U4089 ( .A(\stack[1][3] ), .B(o[6]), .Z(n3956) );
  NAND U4090 ( .A(n3956), .B(n3955), .Z(n3790) );
  NAND U4091 ( .A(n3791), .B(n3790), .Z(n3794) );
  NAND U4092 ( .A(n3794), .B(n3795), .Z(n3797) );
  AND U4093 ( .A(\stack[1][3] ), .B(o[7]), .Z(n3963) );
  NAND U4094 ( .A(n3963), .B(n3964), .Z(n3796) );
  NAND U4095 ( .A(n3797), .B(n3796), .Z(n3800) );
  AND U4096 ( .A(\stack[1][3] ), .B(o[8]), .Z(n3801) );
  NAND U4097 ( .A(n3800), .B(n3801), .Z(n3803) );
  XOR U4098 ( .A(n3799), .B(n3798), .Z(n3923) );
  NAND U4099 ( .A(n3923), .B(n3922), .Z(n3802) );
  NAND U4100 ( .A(n3803), .B(n3802), .Z(n3806) );
  XOR U4101 ( .A(n3805), .B(n3804), .Z(n3807) );
  NAND U4102 ( .A(n3806), .B(n3807), .Z(n3809) );
  AND U4103 ( .A(\stack[1][3] ), .B(o[9]), .Z(n3971) );
  NAND U4104 ( .A(n3971), .B(n3972), .Z(n3808) );
  NAND U4105 ( .A(n3809), .B(n3808), .Z(n3812) );
  AND U4106 ( .A(o[10]), .B(\stack[1][3] ), .Z(n3813) );
  NAND U4107 ( .A(n3812), .B(n3813), .Z(n3815) );
  XNOR U4108 ( .A(n3811), .B(n3810), .Z(n3977) );
  NAND U4109 ( .A(n3977), .B(n3978), .Z(n3814) );
  AND U4110 ( .A(n3815), .B(n3814), .Z(n3817) );
  NAND U4111 ( .A(n3816), .B(n3817), .Z(n3819) );
  NAND U4112 ( .A(\stack[1][3] ), .B(o[11]), .Z(n3983) );
  NAND U4113 ( .A(n3983), .B(n3984), .Z(n3818) );
  AND U4114 ( .A(n3819), .B(n3818), .Z(n3822) );
  AND U4115 ( .A(\stack[1][3] ), .B(o[12]), .Z(n3823) );
  NAND U4116 ( .A(n3822), .B(n3823), .Z(n3825) );
  NAND U4117 ( .A(n3990), .B(n3989), .Z(n3824) );
  NAND U4118 ( .A(n3825), .B(n3824), .Z(n3827) );
  NAND U4119 ( .A(n3826), .B(n3827), .Z(n3829) );
  AND U4120 ( .A(\stack[1][3] ), .B(o[13]), .Z(n3997) );
  NAND U4121 ( .A(n3997), .B(n3998), .Z(n3828) );
  NAND U4122 ( .A(n3829), .B(n3828), .Z(n3832) );
  AND U4123 ( .A(\stack[1][3] ), .B(o[14]), .Z(n3833) );
  NAND U4124 ( .A(n3832), .B(n3833), .Z(n3835) );
  XNOR U4125 ( .A(n3831), .B(n3830), .Z(n4001) );
  NAND U4126 ( .A(n4001), .B(n4002), .Z(n3834) );
  NAND U4127 ( .A(n3835), .B(n3834), .Z(n3838) );
  XNOR U4128 ( .A(n3837), .B(n3836), .Z(n3839) );
  NAND U4129 ( .A(n3838), .B(n3839), .Z(n3841) );
  AND U4130 ( .A(\stack[1][3] ), .B(o[15]), .Z(n4009) );
  NAND U4131 ( .A(n4010), .B(n4009), .Z(n3840) );
  NAND U4132 ( .A(n3841), .B(n3840), .Z(n3844) );
  AND U4133 ( .A(\stack[1][3] ), .B(o[16]), .Z(n3845) );
  NAND U4134 ( .A(n3844), .B(n3845), .Z(n3847) );
  XOR U4135 ( .A(n3843), .B(n3842), .Z(n4014) );
  NAND U4136 ( .A(n4014), .B(n4013), .Z(n3846) );
  NAND U4137 ( .A(n3847), .B(n3846), .Z(n3850) );
  XOR U4138 ( .A(n3849), .B(n3848), .Z(n3851) );
  NAND U4139 ( .A(n3850), .B(n3851), .Z(n3853) );
  AND U4140 ( .A(\stack[1][3] ), .B(o[17]), .Z(n4019) );
  NAND U4141 ( .A(n4019), .B(n4020), .Z(n3852) );
  NAND U4142 ( .A(n3853), .B(n3852), .Z(n3856) );
  AND U4143 ( .A(\stack[1][3] ), .B(o[18]), .Z(n3857) );
  NAND U4144 ( .A(n3856), .B(n3857), .Z(n3859) );
  XOR U4145 ( .A(n3855), .B(n3854), .Z(n4026) );
  NAND U4146 ( .A(n4026), .B(n4025), .Z(n3858) );
  NAND U4147 ( .A(n3859), .B(n3858), .Z(n3860) );
  NAND U4148 ( .A(n3861), .B(n3860), .Z(n3863) );
  AND U4149 ( .A(\stack[1][3] ), .B(o[19]), .Z(n4033) );
  XOR U4150 ( .A(n3861), .B(n3860), .Z(n4034) );
  NAND U4151 ( .A(n4033), .B(n4034), .Z(n3862) );
  NAND U4152 ( .A(n3863), .B(n3862), .Z(n3866) );
  AND U4153 ( .A(\stack[1][3] ), .B(o[20]), .Z(n3867) );
  NAND U4154 ( .A(n3866), .B(n3867), .Z(n3869) );
  XOR U4155 ( .A(n3865), .B(n3864), .Z(n4038) );
  NAND U4156 ( .A(n4038), .B(n4037), .Z(n3868) );
  NAND U4157 ( .A(n3869), .B(n3868), .Z(n3872) );
  XOR U4158 ( .A(n3871), .B(n3870), .Z(n3873) );
  NAND U4159 ( .A(n3872), .B(n3873), .Z(n3875) );
  AND U4160 ( .A(\stack[1][3] ), .B(o[21]), .Z(n4045) );
  NAND U4161 ( .A(n4045), .B(n4046), .Z(n3874) );
  NAND U4162 ( .A(n3875), .B(n3874), .Z(n3878) );
  AND U4163 ( .A(\stack[1][3] ), .B(o[22]), .Z(n3879) );
  NAND U4164 ( .A(n3878), .B(n3879), .Z(n3881) );
  NAND U4165 ( .A(n4050), .B(n4049), .Z(n3880) );
  NAND U4166 ( .A(n3881), .B(n3880), .Z(n3884) );
  XNOR U4167 ( .A(n3883), .B(n3882), .Z(n3885) );
  NAND U4168 ( .A(n3884), .B(n3885), .Z(n3887) );
  AND U4169 ( .A(\stack[1][3] ), .B(o[23]), .Z(n4057) );
  NAND U4170 ( .A(n4058), .B(n4057), .Z(n3886) );
  NAND U4171 ( .A(n3887), .B(n3886), .Z(n3890) );
  AND U4172 ( .A(\stack[1][3] ), .B(o[24]), .Z(n3891) );
  NAND U4173 ( .A(n3890), .B(n3891), .Z(n3893) );
  NAND U4174 ( .A(n4062), .B(n4061), .Z(n3892) );
  NAND U4175 ( .A(n3893), .B(n3892), .Z(n3896) );
  XOR U4176 ( .A(n3895), .B(n3894), .Z(n3897) );
  NAND U4177 ( .A(n3896), .B(n3897), .Z(n3899) );
  AND U4178 ( .A(\stack[1][3] ), .B(o[25]), .Z(n4067) );
  NAND U4179 ( .A(n4067), .B(n4068), .Z(n3898) );
  NAND U4180 ( .A(n3899), .B(n3898), .Z(n3902) );
  NAND U4181 ( .A(n3903), .B(n3902), .Z(n3905) );
  XOR U4182 ( .A(n3901), .B(n3900), .Z(n4074) );
  XOR U4183 ( .A(n3903), .B(n3902), .Z(n4073) );
  NAND U4184 ( .A(n4074), .B(n4073), .Z(n3904) );
  NAND U4185 ( .A(n3905), .B(n3904), .Z(n3906) );
  XOR U4186 ( .A(n3907), .B(n3906), .Z(n4080) );
  AND U4187 ( .A(\stack[1][3] ), .B(o[27]), .Z(n4079) );
  NAND U4188 ( .A(n4080), .B(n4079), .Z(n3909) );
  NAND U4189 ( .A(n3907), .B(n3906), .Z(n3908) );
  AND U4190 ( .A(n3909), .B(n3908), .Z(n3917) );
  NAND U4191 ( .A(n3911), .B(n3910), .Z(n3915) );
  NAND U4192 ( .A(n3913), .B(n3912), .Z(n3914) );
  NAND U4193 ( .A(n3915), .B(n3914), .Z(n3916) );
  XNOR U4194 ( .A(n3917), .B(n3916), .Z(n3918) );
  XNOR U4195 ( .A(n3919), .B(n3918), .Z(n3920) );
  XNOR U4196 ( .A(n3921), .B(n3920), .Z(n4428) );
  NAND U4197 ( .A(\stack[1][2] ), .B(o[24]), .Z(n4055) );
  NAND U4198 ( .A(\stack[1][2] ), .B(o[16]), .Z(n4007) );
  AND U4199 ( .A(\stack[1][2] ), .B(o[14]), .Z(n3995) );
  NAND U4200 ( .A(\stack[1][2] ), .B(o[12]), .Z(n3985) );
  XNOR U4201 ( .A(n3923), .B(n3922), .Z(n3967) );
  AND U4202 ( .A(\stack[1][2] ), .B(o[5]), .Z(n3945) );
  XOR U4203 ( .A(n3925), .B(n3924), .Z(n3946) );
  NAND U4204 ( .A(n3945), .B(n3946), .Z(n3948) );
  AND U4205 ( .A(\stack[1][2] ), .B(o[0]), .Z(n4271) );
  AND U4206 ( .A(\stack[1][3] ), .B(o[1]), .Z(n3928) );
  AND U4207 ( .A(n4271), .B(n3928), .Z(n3926) );
  NAND U4208 ( .A(o[2]), .B(n3926), .Z(n3932) );
  NAND U4209 ( .A(\stack[1][4] ), .B(o[0]), .Z(n3927) );
  XNOR U4210 ( .A(n3928), .B(n3927), .Z(n4093) );
  NAND U4211 ( .A(o[0]), .B(n3928), .Z(n3929) );
  XNOR U4212 ( .A(o[2]), .B(n3929), .Z(n3930) );
  AND U4213 ( .A(\stack[1][2] ), .B(n3930), .Z(n4094) );
  NAND U4214 ( .A(n4093), .B(n4094), .Z(n3931) );
  NAND U4215 ( .A(n3932), .B(n3931), .Z(n3935) );
  NAND U4216 ( .A(n3935), .B(n3936), .Z(n3938) );
  AND U4217 ( .A(\stack[1][2] ), .B(o[3]), .Z(n4100) );
  NAND U4218 ( .A(n4100), .B(n4099), .Z(n3937) );
  NAND U4219 ( .A(n3938), .B(n3937), .Z(n3941) );
  AND U4220 ( .A(\stack[1][2] ), .B(o[4]), .Z(n3942) );
  NAND U4221 ( .A(n3941), .B(n3942), .Z(n3944) );
  XOR U4222 ( .A(n3940), .B(n3939), .Z(n4106) );
  NAND U4223 ( .A(n4106), .B(n4105), .Z(n3943) );
  NAND U4224 ( .A(n3944), .B(n3943), .Z(n4111) );
  NAND U4225 ( .A(n4111), .B(n4112), .Z(n3947) );
  NAND U4226 ( .A(n3948), .B(n3947), .Z(n3951) );
  NAND U4227 ( .A(n3951), .B(n3952), .Z(n3954) );
  AND U4228 ( .A(\stack[1][2] ), .B(o[6]), .Z(n4117) );
  NAND U4229 ( .A(n4117), .B(n4118), .Z(n3953) );
  NAND U4230 ( .A(n3954), .B(n3953), .Z(n3957) );
  XOR U4231 ( .A(n3956), .B(n3955), .Z(n3958) );
  NAND U4232 ( .A(n3957), .B(n3958), .Z(n3960) );
  AND U4233 ( .A(\stack[1][2] ), .B(o[7]), .Z(n4123) );
  NAND U4234 ( .A(n4123), .B(n4124), .Z(n3959) );
  NAND U4235 ( .A(n3960), .B(n3959), .Z(n3961) );
  AND U4236 ( .A(\stack[1][2] ), .B(o[8]), .Z(n3962) );
  NAND U4237 ( .A(n3961), .B(n3962), .Z(n3966) );
  NAND U4238 ( .A(n4130), .B(n4129), .Z(n3965) );
  AND U4239 ( .A(n3966), .B(n3965), .Z(n3968) );
  NAND U4240 ( .A(n3967), .B(n3968), .Z(n3970) );
  NAND U4241 ( .A(\stack[1][2] ), .B(o[9]), .Z(n4135) );
  NAND U4242 ( .A(n4136), .B(n4135), .Z(n3969) );
  AND U4243 ( .A(n3970), .B(n3969), .Z(n3973) );
  AND U4244 ( .A(\stack[1][2] ), .B(o[10]), .Z(n3974) );
  NAND U4245 ( .A(n3973), .B(n3974), .Z(n3976) );
  NAND U4246 ( .A(n4084), .B(n4083), .Z(n3975) );
  NAND U4247 ( .A(n3976), .B(n3975), .Z(n3979) );
  NAND U4248 ( .A(n3979), .B(n3980), .Z(n3982) );
  AND U4249 ( .A(\stack[1][2] ), .B(o[11]), .Z(n4146) );
  NAND U4250 ( .A(n4146), .B(n4145), .Z(n3981) );
  AND U4251 ( .A(n3982), .B(n3981), .Z(n3986) );
  NAND U4252 ( .A(n3985), .B(n3986), .Z(n3988) );
  NAND U4253 ( .A(n4082), .B(n4081), .Z(n3987) );
  NAND U4254 ( .A(n3988), .B(n3987), .Z(n3991) );
  XNOR U4255 ( .A(n3990), .B(n3989), .Z(n3992) );
  NAND U4256 ( .A(n3991), .B(n3992), .Z(n3994) );
  NAND U4257 ( .A(\stack[1][2] ), .B(o[13]), .Z(n4155) );
  NAND U4258 ( .A(n4156), .B(n4155), .Z(n3993) );
  AND U4259 ( .A(n3994), .B(n3993), .Z(n3996) );
  NAND U4260 ( .A(n3995), .B(n3996), .Z(n4000) );
  NAND U4261 ( .A(n4162), .B(n4161), .Z(n3999) );
  NAND U4262 ( .A(n4000), .B(n3999), .Z(n4003) );
  NAND U4263 ( .A(n4003), .B(n4004), .Z(n4006) );
  AND U4264 ( .A(\stack[1][2] ), .B(o[15]), .Z(n4168) );
  NAND U4265 ( .A(n4168), .B(n4167), .Z(n4005) );
  AND U4266 ( .A(n4006), .B(n4005), .Z(n4008) );
  NAND U4267 ( .A(n4007), .B(n4008), .Z(n4012) );
  XNOR U4268 ( .A(n4010), .B(n4009), .Z(n4173) );
  NAND U4269 ( .A(n4174), .B(n4173), .Z(n4011) );
  AND U4270 ( .A(n4012), .B(n4011), .Z(n4016) );
  XOR U4271 ( .A(n4014), .B(n4013), .Z(n4015) );
  NAND U4272 ( .A(n4016), .B(n4015), .Z(n4018) );
  AND U4273 ( .A(\stack[1][2] ), .B(o[17]), .Z(n4179) );
  XOR U4274 ( .A(n4016), .B(n4015), .Z(n4180) );
  NAND U4275 ( .A(n4179), .B(n4180), .Z(n4017) );
  NAND U4276 ( .A(n4018), .B(n4017), .Z(n4021) );
  AND U4277 ( .A(\stack[1][2] ), .B(o[18]), .Z(n4022) );
  NAND U4278 ( .A(n4021), .B(n4022), .Z(n4024) );
  NAND U4279 ( .A(n4186), .B(n4185), .Z(n4023) );
  NAND U4280 ( .A(n4024), .B(n4023), .Z(n4027) );
  XOR U4281 ( .A(n4026), .B(n4025), .Z(n4028) );
  NAND U4282 ( .A(n4027), .B(n4028), .Z(n4030) );
  AND U4283 ( .A(\stack[1][2] ), .B(o[19]), .Z(n4191) );
  NAND U4284 ( .A(n4191), .B(n4192), .Z(n4029) );
  NAND U4285 ( .A(n4030), .B(n4029), .Z(n4031) );
  AND U4286 ( .A(\stack[1][2] ), .B(o[20]), .Z(n4032) );
  NAND U4287 ( .A(n4031), .B(n4032), .Z(n4036) );
  NAND U4288 ( .A(n4198), .B(n4197), .Z(n4035) );
  NAND U4289 ( .A(n4036), .B(n4035), .Z(n4039) );
  XOR U4290 ( .A(n4038), .B(n4037), .Z(n4040) );
  NAND U4291 ( .A(n4039), .B(n4040), .Z(n4042) );
  AND U4292 ( .A(\stack[1][2] ), .B(o[21]), .Z(n4204) );
  NAND U4293 ( .A(n4204), .B(n4203), .Z(n4041) );
  NAND U4294 ( .A(n4042), .B(n4041), .Z(n4043) );
  AND U4295 ( .A(\stack[1][2] ), .B(o[22]), .Z(n4044) );
  NAND U4296 ( .A(n4043), .B(n4044), .Z(n4048) );
  NAND U4297 ( .A(n4210), .B(n4209), .Z(n4047) );
  NAND U4298 ( .A(n4048), .B(n4047), .Z(n4051) );
  XOR U4299 ( .A(n4050), .B(n4049), .Z(n4052) );
  NAND U4300 ( .A(n4051), .B(n4052), .Z(n4054) );
  AND U4301 ( .A(\stack[1][2] ), .B(o[23]), .Z(n4215) );
  NAND U4302 ( .A(n4215), .B(n4216), .Z(n4053) );
  AND U4303 ( .A(n4054), .B(n4053), .Z(n4056) );
  NAND U4304 ( .A(n4055), .B(n4056), .Z(n4060) );
  XNOR U4305 ( .A(n4058), .B(n4057), .Z(n4221) );
  NAND U4306 ( .A(n4222), .B(n4221), .Z(n4059) );
  AND U4307 ( .A(n4060), .B(n4059), .Z(n4064) );
  XOR U4308 ( .A(n4062), .B(n4061), .Z(n4063) );
  NAND U4309 ( .A(n4064), .B(n4063), .Z(n4066) );
  AND U4310 ( .A(\stack[1][2] ), .B(o[25]), .Z(n4228) );
  XOR U4311 ( .A(n4064), .B(n4063), .Z(n4227) );
  NAND U4312 ( .A(n4228), .B(n4227), .Z(n4065) );
  NAND U4313 ( .A(n4066), .B(n4065), .Z(n4069) );
  AND U4314 ( .A(\stack[1][2] ), .B(o[26]), .Z(n4070) );
  NAND U4315 ( .A(n4069), .B(n4070), .Z(n4072) );
  NAND U4316 ( .A(n4234), .B(n4233), .Z(n4071) );
  NAND U4317 ( .A(n4072), .B(n4071), .Z(n4075) );
  XOR U4318 ( .A(n4074), .B(n4073), .Z(n4076) );
  NAND U4319 ( .A(n4075), .B(n4076), .Z(n4078) );
  AND U4320 ( .A(\stack[1][2] ), .B(o[27]), .Z(n4239) );
  NAND U4321 ( .A(n4239), .B(n4240), .Z(n4077) );
  NAND U4322 ( .A(n4078), .B(n4077), .Z(n4431) );
  AND U4323 ( .A(\stack[1][2] ), .B(o[28]), .Z(n4432) );
  XOR U4324 ( .A(n4431), .B(n4432), .Z(n4434) );
  XOR U4325 ( .A(n4080), .B(n4079), .Z(n4433) );
  XOR U4326 ( .A(n4434), .B(n4433), .Z(n4421) );
  XNOR U4327 ( .A(n4082), .B(n4081), .Z(n4151) );
  XNOR U4328 ( .A(n4084), .B(n4083), .Z(n4141) );
  AND U4329 ( .A(o[0]), .B(\stack[1][1] ), .Z(n5576) );
  AND U4330 ( .A(\stack[1][2] ), .B(o[1]), .Z(n4088) );
  AND U4331 ( .A(n5576), .B(n4088), .Z(n4085) );
  NAND U4332 ( .A(o[2]), .B(n4085), .Z(n4092) );
  NAND U4333 ( .A(o[1]), .B(\stack[1][2] ), .Z(n4086) );
  XNOR U4334 ( .A(n4087), .B(n4086), .Z(n4278) );
  NAND U4335 ( .A(n4088), .B(o[0]), .Z(n4089) );
  XNOR U4336 ( .A(o[2]), .B(n4089), .Z(n4090) );
  AND U4337 ( .A(\stack[1][1] ), .B(n4090), .Z(n4277) );
  NAND U4338 ( .A(n4278), .B(n4277), .Z(n4091) );
  NAND U4339 ( .A(n4092), .B(n4091), .Z(n4095) );
  NAND U4340 ( .A(n4095), .B(n4096), .Z(n4098) );
  AND U4341 ( .A(o[3]), .B(\stack[1][1] ), .Z(n4265) );
  NAND U4342 ( .A(n4266), .B(n4265), .Z(n4097) );
  NAND U4343 ( .A(n4098), .B(n4097), .Z(n4101) );
  AND U4344 ( .A(o[4]), .B(\stack[1][1] ), .Z(n4102) );
  NAND U4345 ( .A(n4101), .B(n4102), .Z(n4104) );
  XOR U4346 ( .A(n4100), .B(n4099), .Z(n4288) );
  NAND U4347 ( .A(n4288), .B(n4287), .Z(n4103) );
  NAND U4348 ( .A(n4104), .B(n4103), .Z(n4107) );
  XOR U4349 ( .A(n4106), .B(n4105), .Z(n4108) );
  NAND U4350 ( .A(n4107), .B(n4108), .Z(n4110) );
  AND U4351 ( .A(o[5]), .B(\stack[1][1] ), .Z(n4263) );
  NAND U4352 ( .A(n4264), .B(n4263), .Z(n4109) );
  NAND U4353 ( .A(n4110), .B(n4109), .Z(n4113) );
  NAND U4354 ( .A(n4113), .B(n4114), .Z(n4116) );
  AND U4355 ( .A(o[6]), .B(\stack[1][1] ), .Z(n4298) );
  NAND U4356 ( .A(n4298), .B(n4297), .Z(n4115) );
  NAND U4357 ( .A(n4116), .B(n4115), .Z(n4119) );
  NAND U4358 ( .A(n4119), .B(n4120), .Z(n4122) );
  AND U4359 ( .A(o[7]), .B(\stack[1][1] ), .Z(n4302) );
  NAND U4360 ( .A(n4302), .B(n4301), .Z(n4121) );
  NAND U4361 ( .A(n4122), .B(n4121), .Z(n4125) );
  AND U4362 ( .A(o[8]), .B(\stack[1][1] ), .Z(n4126) );
  NAND U4363 ( .A(n4125), .B(n4126), .Z(n4128) );
  NAND U4364 ( .A(n4310), .B(n4309), .Z(n4127) );
  NAND U4365 ( .A(n4128), .B(n4127), .Z(n4131) );
  XOR U4366 ( .A(n4130), .B(n4129), .Z(n4132) );
  NAND U4367 ( .A(n4131), .B(n4132), .Z(n4134) );
  AND U4368 ( .A(o[9]), .B(\stack[1][1] ), .Z(n4261) );
  NAND U4369 ( .A(n4262), .B(n4261), .Z(n4133) );
  NAND U4370 ( .A(n4134), .B(n4133), .Z(n4137) );
  AND U4371 ( .A(o[10]), .B(\stack[1][1] ), .Z(n4138) );
  NAND U4372 ( .A(n4137), .B(n4138), .Z(n4140) );
  XOR U4373 ( .A(n4136), .B(n4135), .Z(n4320) );
  NANDN U4374 ( .A(n4320), .B(n4319), .Z(n4139) );
  AND U4375 ( .A(n4140), .B(n4139), .Z(n4142) );
  NAND U4376 ( .A(n4141), .B(n4142), .Z(n4144) );
  NAND U4377 ( .A(o[11]), .B(\stack[1][1] ), .Z(n4323) );
  NAND U4378 ( .A(n4323), .B(n4324), .Z(n4143) );
  AND U4379 ( .A(n4144), .B(n4143), .Z(n4147) );
  AND U4380 ( .A(o[12]), .B(\stack[1][1] ), .Z(n4148) );
  NAND U4381 ( .A(n4147), .B(n4148), .Z(n4150) );
  XOR U4382 ( .A(n4146), .B(n4145), .Z(n4332) );
  NAND U4383 ( .A(n4332), .B(n4331), .Z(n4149) );
  NAND U4384 ( .A(n4150), .B(n4149), .Z(n4152) );
  NAND U4385 ( .A(n4151), .B(n4152), .Z(n4154) );
  AND U4386 ( .A(o[13]), .B(\stack[1][1] ), .Z(n4259) );
  NAND U4387 ( .A(n4260), .B(n4259), .Z(n4153) );
  NAND U4388 ( .A(n4154), .B(n4153), .Z(n4157) );
  AND U4389 ( .A(o[14]), .B(\stack[1][1] ), .Z(n4158) );
  NAND U4390 ( .A(n4157), .B(n4158), .Z(n4160) );
  XOR U4391 ( .A(n4156), .B(n4155), .Z(n4342) );
  NANDN U4392 ( .A(n4342), .B(n4341), .Z(n4159) );
  NAND U4393 ( .A(n4160), .B(n4159), .Z(n4163) );
  XOR U4394 ( .A(n4162), .B(n4161), .Z(n4164) );
  NAND U4395 ( .A(n4163), .B(n4164), .Z(n4166) );
  AND U4396 ( .A(o[15]), .B(\stack[1][1] ), .Z(n4257) );
  NAND U4397 ( .A(n4258), .B(n4257), .Z(n4165) );
  NAND U4398 ( .A(n4166), .B(n4165), .Z(n4169) );
  AND U4399 ( .A(o[16]), .B(\stack[1][1] ), .Z(n4170) );
  NAND U4400 ( .A(n4169), .B(n4170), .Z(n4172) );
  XOR U4401 ( .A(n4168), .B(n4167), .Z(n4352) );
  NAND U4402 ( .A(n4352), .B(n4351), .Z(n4171) );
  NAND U4403 ( .A(n4172), .B(n4171), .Z(n4175) );
  XNOR U4404 ( .A(n4174), .B(n4173), .Z(n4176) );
  NAND U4405 ( .A(n4175), .B(n4176), .Z(n4178) );
  AND U4406 ( .A(o[17]), .B(\stack[1][1] ), .Z(n4255) );
  NAND U4407 ( .A(n4256), .B(n4255), .Z(n4177) );
  NAND U4408 ( .A(n4178), .B(n4177), .Z(n4181) );
  AND U4409 ( .A(o[18]), .B(\stack[1][1] ), .Z(n4182) );
  NAND U4410 ( .A(n4181), .B(n4182), .Z(n4184) );
  NAND U4411 ( .A(n4362), .B(n4361), .Z(n4183) );
  NAND U4412 ( .A(n4184), .B(n4183), .Z(n4187) );
  XOR U4413 ( .A(n4186), .B(n4185), .Z(n4188) );
  NAND U4414 ( .A(n4187), .B(n4188), .Z(n4190) );
  AND U4415 ( .A(o[19]), .B(\stack[1][1] ), .Z(n4253) );
  NAND U4416 ( .A(n4254), .B(n4253), .Z(n4189) );
  NAND U4417 ( .A(n4190), .B(n4189), .Z(n4193) );
  AND U4418 ( .A(o[20]), .B(\stack[1][1] ), .Z(n4194) );
  NAND U4419 ( .A(n4193), .B(n4194), .Z(n4196) );
  NAND U4420 ( .A(n4372), .B(n4371), .Z(n4195) );
  NAND U4421 ( .A(n4196), .B(n4195), .Z(n4199) );
  XOR U4422 ( .A(n4198), .B(n4197), .Z(n4200) );
  NAND U4423 ( .A(n4199), .B(n4200), .Z(n4202) );
  AND U4424 ( .A(o[21]), .B(\stack[1][1] ), .Z(n4251) );
  NAND U4425 ( .A(n4252), .B(n4251), .Z(n4201) );
  NAND U4426 ( .A(n4202), .B(n4201), .Z(n4205) );
  AND U4427 ( .A(o[22]), .B(\stack[1][1] ), .Z(n4206) );
  NAND U4428 ( .A(n4205), .B(n4206), .Z(n4208) );
  XOR U4429 ( .A(n4204), .B(n4203), .Z(n4382) );
  NAND U4430 ( .A(n4382), .B(n4381), .Z(n4207) );
  NAND U4431 ( .A(n4208), .B(n4207), .Z(n4211) );
  XOR U4432 ( .A(n4210), .B(n4209), .Z(n4212) );
  NAND U4433 ( .A(n4211), .B(n4212), .Z(n4214) );
  AND U4434 ( .A(o[23]), .B(\stack[1][1] ), .Z(n4249) );
  NAND U4435 ( .A(n4250), .B(n4249), .Z(n4213) );
  NAND U4436 ( .A(n4214), .B(n4213), .Z(n4217) );
  AND U4437 ( .A(o[24]), .B(\stack[1][1] ), .Z(n4218) );
  NAND U4438 ( .A(n4217), .B(n4218), .Z(n4220) );
  NAND U4439 ( .A(n4392), .B(n4391), .Z(n4219) );
  NAND U4440 ( .A(n4220), .B(n4219), .Z(n4223) );
  XNOR U4441 ( .A(n4222), .B(n4221), .Z(n4224) );
  NAND U4442 ( .A(n4223), .B(n4224), .Z(n4226) );
  AND U4443 ( .A(o[25]), .B(\stack[1][1] ), .Z(n4247) );
  NAND U4444 ( .A(n4248), .B(n4247), .Z(n4225) );
  NAND U4445 ( .A(n4226), .B(n4225), .Z(n4229) );
  AND U4446 ( .A(o[26]), .B(\stack[1][1] ), .Z(n4230) );
  NAND U4447 ( .A(n4229), .B(n4230), .Z(n4232) );
  XOR U4448 ( .A(n4228), .B(n4227), .Z(n4402) );
  NAND U4449 ( .A(n4402), .B(n4401), .Z(n4231) );
  NAND U4450 ( .A(n4232), .B(n4231), .Z(n4235) );
  XOR U4451 ( .A(n4234), .B(n4233), .Z(n4236) );
  NAND U4452 ( .A(n4235), .B(n4236), .Z(n4238) );
  AND U4453 ( .A(o[27]), .B(\stack[1][1] ), .Z(n4245) );
  NAND U4454 ( .A(n4246), .B(n4245), .Z(n4237) );
  NAND U4455 ( .A(n4238), .B(n4237), .Z(n4241) );
  AND U4456 ( .A(o[28]), .B(\stack[1][1] ), .Z(n4242) );
  NAND U4457 ( .A(n4241), .B(n4242), .Z(n4244) );
  NAND U4458 ( .A(n4412), .B(n4411), .Z(n4243) );
  NAND U4459 ( .A(n4244), .B(n4243), .Z(n4422) );
  AND U4460 ( .A(\stack[1][1] ), .B(o[29]), .Z(n4419) );
  XNOR U4461 ( .A(n4420), .B(n4419), .Z(n4416) );
  NAND U4462 ( .A(o[29]), .B(\stack[1][0] ), .Z(n4409) );
  XNOR U4463 ( .A(n4246), .B(n4245), .Z(n4405) );
  NAND U4464 ( .A(o[27]), .B(\stack[1][0] ), .Z(n4399) );
  XNOR U4465 ( .A(n4248), .B(n4247), .Z(n4395) );
  NAND U4466 ( .A(o[25]), .B(\stack[1][0] ), .Z(n4389) );
  XNOR U4467 ( .A(n4250), .B(n4249), .Z(n4385) );
  NAND U4468 ( .A(o[23]), .B(\stack[1][0] ), .Z(n4379) );
  XNOR U4469 ( .A(n4252), .B(n4251), .Z(n4375) );
  NAND U4470 ( .A(o[21]), .B(\stack[1][0] ), .Z(n4369) );
  XNOR U4471 ( .A(n4254), .B(n4253), .Z(n4365) );
  NAND U4472 ( .A(o[19]), .B(\stack[1][0] ), .Z(n4359) );
  XNOR U4473 ( .A(n4256), .B(n4255), .Z(n4355) );
  NAND U4474 ( .A(o[17]), .B(\stack[1][0] ), .Z(n4349) );
  XNOR U4475 ( .A(n4258), .B(n4257), .Z(n4345) );
  NAND U4476 ( .A(o[15]), .B(\stack[1][0] ), .Z(n4339) );
  XNOR U4477 ( .A(n4260), .B(n4259), .Z(n4335) );
  NAND U4478 ( .A(o[13]), .B(\stack[1][0] ), .Z(n4329) );
  NAND U4479 ( .A(o[11]), .B(\stack[1][0] ), .Z(n4317) );
  XNOR U4480 ( .A(n4262), .B(n4261), .Z(n4313) );
  NAND U4481 ( .A(o[9]), .B(\stack[1][0] ), .Z(n4307) );
  NAND U4482 ( .A(o[7]), .B(\stack[1][0] ), .Z(n4295) );
  XNOR U4483 ( .A(n4264), .B(n4263), .Z(n4291) );
  NAND U4484 ( .A(o[5]), .B(\stack[1][0] ), .Z(n4285) );
  XNOR U4485 ( .A(n4266), .B(n4265), .Z(n4281) );
  NAND U4486 ( .A(o[3]), .B(\stack[1][0] ), .Z(n4275) );
  AND U4487 ( .A(o[1]), .B(\stack[1][0] ), .Z(n5575) );
  NAND U4488 ( .A(n5576), .B(n5575), .Z(n4268) );
  NAND U4489 ( .A(o[2]), .B(\stack[1][0] ), .Z(n4267) );
  AND U4490 ( .A(n4268), .B(n4267), .Z(n4274) );
  NAND U4491 ( .A(n5576), .B(o[1]), .Z(n4269) );
  XNOR U4492 ( .A(o[2]), .B(n4269), .Z(n4270) );
  AND U4493 ( .A(\stack[1][0] ), .B(n4270), .Z(n5546) );
  AND U4494 ( .A(\stack[1][1] ), .B(o[1]), .Z(n4272) );
  XNOR U4495 ( .A(n4272), .B(n4271), .Z(n5547) );
  NAND U4496 ( .A(n5546), .B(n5547), .Z(n4273) );
  NANDN U4497 ( .A(n4274), .B(n4273), .Z(n4276) );
  NAND U4498 ( .A(n4275), .B(n4276), .Z(n4280) );
  XNOR U4499 ( .A(n4278), .B(n4277), .Z(n5512) );
  NAND U4500 ( .A(n5511), .B(n5512), .Z(n4279) );
  NAND U4501 ( .A(n4280), .B(n4279), .Z(n4282) );
  NAND U4502 ( .A(n4281), .B(n4282), .Z(n4284) );
  NAND U4503 ( .A(o[4]), .B(\stack[1][0] ), .Z(n5474) );
  NAND U4504 ( .A(n5473), .B(n5474), .Z(n4283) );
  NAND U4505 ( .A(n4284), .B(n4283), .Z(n4286) );
  NAND U4506 ( .A(n4285), .B(n4286), .Z(n4290) );
  XNOR U4507 ( .A(n4288), .B(n4287), .Z(n5436) );
  NAND U4508 ( .A(n5435), .B(n5436), .Z(n4289) );
  NAND U4509 ( .A(n4290), .B(n4289), .Z(n4292) );
  NAND U4510 ( .A(n4291), .B(n4292), .Z(n4294) );
  NAND U4511 ( .A(o[6]), .B(\stack[1][0] ), .Z(n5398) );
  NAND U4512 ( .A(n5397), .B(n5398), .Z(n4293) );
  NAND U4513 ( .A(n4294), .B(n4293), .Z(n4296) );
  NAND U4514 ( .A(n4295), .B(n4296), .Z(n4300) );
  XNOR U4515 ( .A(n4298), .B(n4297), .Z(n5359) );
  NAND U4516 ( .A(n5358), .B(n5359), .Z(n4299) );
  NAND U4517 ( .A(n4300), .B(n4299), .Z(n4303) );
  XNOR U4518 ( .A(n4302), .B(n4301), .Z(n4304) );
  NAND U4519 ( .A(n4303), .B(n4304), .Z(n4306) );
  NAND U4520 ( .A(o[8]), .B(\stack[1][0] ), .Z(n5320) );
  NAND U4521 ( .A(n5319), .B(n5320), .Z(n4305) );
  NAND U4522 ( .A(n4306), .B(n4305), .Z(n4308) );
  NAND U4523 ( .A(n4307), .B(n4308), .Z(n4312) );
  XNOR U4524 ( .A(n4310), .B(n4309), .Z(n5281) );
  NAND U4525 ( .A(n5280), .B(n5281), .Z(n4311) );
  NAND U4526 ( .A(n4312), .B(n4311), .Z(n4314) );
  NAND U4527 ( .A(n4313), .B(n4314), .Z(n4316) );
  NAND U4528 ( .A(o[10]), .B(\stack[1][0] ), .Z(n5243) );
  NAND U4529 ( .A(n5242), .B(n5243), .Z(n4315) );
  NAND U4530 ( .A(n4316), .B(n4315), .Z(n4318) );
  NAND U4531 ( .A(n4317), .B(n4318), .Z(n4322) );
  XOR U4532 ( .A(n4320), .B(n4319), .Z(n5205) );
  NAND U4533 ( .A(n5204), .B(n5205), .Z(n4321) );
  NAND U4534 ( .A(n4322), .B(n4321), .Z(n4325) );
  NAND U4535 ( .A(n4325), .B(n4326), .Z(n4328) );
  NAND U4536 ( .A(o[12]), .B(\stack[1][0] ), .Z(n5167) );
  NAND U4537 ( .A(n5166), .B(n5167), .Z(n4327) );
  NAND U4538 ( .A(n4328), .B(n4327), .Z(n4330) );
  NAND U4539 ( .A(n4329), .B(n4330), .Z(n4334) );
  XNOR U4540 ( .A(n4332), .B(n4331), .Z(n5129) );
  NAND U4541 ( .A(n5128), .B(n5129), .Z(n4333) );
  NAND U4542 ( .A(n4334), .B(n4333), .Z(n4336) );
  NAND U4543 ( .A(n4335), .B(n4336), .Z(n4338) );
  NAND U4544 ( .A(o[14]), .B(\stack[1][0] ), .Z(n5091) );
  NAND U4545 ( .A(n5090), .B(n5091), .Z(n4337) );
  NAND U4546 ( .A(n4338), .B(n4337), .Z(n4340) );
  NAND U4547 ( .A(n4339), .B(n4340), .Z(n4344) );
  XOR U4548 ( .A(n4342), .B(n4341), .Z(n5051) );
  NAND U4549 ( .A(n5050), .B(n5051), .Z(n4343) );
  NAND U4550 ( .A(n4344), .B(n4343), .Z(n4346) );
  NAND U4551 ( .A(n4345), .B(n4346), .Z(n4348) );
  NAND U4552 ( .A(o[16]), .B(\stack[1][0] ), .Z(n5013) );
  NAND U4553 ( .A(n5012), .B(n5013), .Z(n4347) );
  NAND U4554 ( .A(n4348), .B(n4347), .Z(n4350) );
  NAND U4555 ( .A(n4349), .B(n4350), .Z(n4354) );
  XNOR U4556 ( .A(n4352), .B(n4351), .Z(n4974) );
  NAND U4557 ( .A(n4973), .B(n4974), .Z(n4353) );
  NAND U4558 ( .A(n4354), .B(n4353), .Z(n4356) );
  NAND U4559 ( .A(n4355), .B(n4356), .Z(n4358) );
  NAND U4560 ( .A(o[18]), .B(\stack[1][0] ), .Z(n4937) );
  NAND U4561 ( .A(n4936), .B(n4937), .Z(n4357) );
  NAND U4562 ( .A(n4358), .B(n4357), .Z(n4360) );
  NAND U4563 ( .A(n4359), .B(n4360), .Z(n4364) );
  XNOR U4564 ( .A(n4362), .B(n4361), .Z(n4898) );
  NAND U4565 ( .A(n4897), .B(n4898), .Z(n4363) );
  NAND U4566 ( .A(n4364), .B(n4363), .Z(n4366) );
  NAND U4567 ( .A(n4365), .B(n4366), .Z(n4368) );
  NAND U4568 ( .A(o[20]), .B(\stack[1][0] ), .Z(n4861) );
  NAND U4569 ( .A(n4860), .B(n4861), .Z(n4367) );
  NAND U4570 ( .A(n4368), .B(n4367), .Z(n4370) );
  NAND U4571 ( .A(n4369), .B(n4370), .Z(n4374) );
  XNOR U4572 ( .A(n4372), .B(n4371), .Z(n4822) );
  NAND U4573 ( .A(n4821), .B(n4822), .Z(n4373) );
  NAND U4574 ( .A(n4374), .B(n4373), .Z(n4376) );
  NAND U4575 ( .A(n4375), .B(n4376), .Z(n4378) );
  NAND U4576 ( .A(o[22]), .B(\stack[1][0] ), .Z(n4785) );
  NAND U4577 ( .A(n4784), .B(n4785), .Z(n4377) );
  NAND U4578 ( .A(n4378), .B(n4377), .Z(n4380) );
  NAND U4579 ( .A(n4379), .B(n4380), .Z(n4384) );
  XNOR U4580 ( .A(n4382), .B(n4381), .Z(n4746) );
  NAND U4581 ( .A(n4745), .B(n4746), .Z(n4383) );
  NAND U4582 ( .A(n4384), .B(n4383), .Z(n4386) );
  NAND U4583 ( .A(n4385), .B(n4386), .Z(n4388) );
  NAND U4584 ( .A(o[24]), .B(\stack[1][0] ), .Z(n4709) );
  NAND U4585 ( .A(n4708), .B(n4709), .Z(n4387) );
  NAND U4586 ( .A(n4388), .B(n4387), .Z(n4390) );
  NAND U4587 ( .A(n4389), .B(n4390), .Z(n4394) );
  XNOR U4588 ( .A(n4392), .B(n4391), .Z(n4670) );
  NAND U4589 ( .A(n4669), .B(n4670), .Z(n4393) );
  NAND U4590 ( .A(n4394), .B(n4393), .Z(n4396) );
  NAND U4591 ( .A(n4395), .B(n4396), .Z(n4398) );
  NAND U4592 ( .A(o[26]), .B(\stack[1][0] ), .Z(n4633) );
  NAND U4593 ( .A(n4632), .B(n4633), .Z(n4397) );
  NAND U4594 ( .A(n4398), .B(n4397), .Z(n4400) );
  NAND U4595 ( .A(n4399), .B(n4400), .Z(n4404) );
  XNOR U4596 ( .A(n4402), .B(n4401), .Z(n4594) );
  NAND U4597 ( .A(n4593), .B(n4594), .Z(n4403) );
  NAND U4598 ( .A(n4404), .B(n4403), .Z(n4406) );
  NAND U4599 ( .A(n4405), .B(n4406), .Z(n4408) );
  NAND U4600 ( .A(o[28]), .B(\stack[1][0] ), .Z(n4557) );
  NAND U4601 ( .A(n4556), .B(n4557), .Z(n4407) );
  NAND U4602 ( .A(n4408), .B(n4407), .Z(n4410) );
  NAND U4603 ( .A(n4409), .B(n4410), .Z(n4414) );
  XNOR U4604 ( .A(n4412), .B(n4411), .Z(n4518) );
  NAND U4605 ( .A(n4517), .B(n4518), .Z(n4413) );
  NAND U4606 ( .A(n4414), .B(n4413), .Z(n4415) );
  NAND U4607 ( .A(\stack[1][0] ), .B(o[30]), .Z(n4481) );
  NAND U4608 ( .A(n4480), .B(n4481), .Z(n4418) );
  NAND U4609 ( .A(n4416), .B(n4415), .Z(n4417) );
  AND U4610 ( .A(n4418), .B(n4417), .Z(n4426) );
  NAND U4611 ( .A(n4420), .B(n4419), .Z(n4424) );
  NAND U4612 ( .A(n4422), .B(n4421), .Z(n4423) );
  NAND U4613 ( .A(n4424), .B(n4423), .Z(n4425) );
  XNOR U4614 ( .A(n4426), .B(n4425), .Z(n4427) );
  XNOR U4615 ( .A(n4428), .B(n4427), .Z(n4429) );
  XNOR U4616 ( .A(n4430), .B(n4429), .Z(n4438) );
  NAND U4617 ( .A(n4432), .B(n4431), .Z(n4436) );
  NAND U4618 ( .A(n4434), .B(n4433), .Z(n4435) );
  NAND U4619 ( .A(n4436), .B(n4435), .Z(n4437) );
  XNOR U4620 ( .A(n4438), .B(n4437), .Z(n4439) );
  AND U4621 ( .A(n5578), .B(n4439), .Z(n4443) );
  AND U4622 ( .A(opcode[2]), .B(n5595), .Z(n5598) );
  NAND U4623 ( .A(\stack[1][31] ), .B(n5598), .Z(n4441) );
  AND U4624 ( .A(n5603), .B(x[31]), .Z(n4440) );
  ANDN U4625 ( .B(n4441), .A(n4440), .Z(n4442) );
  NANDN U4626 ( .A(n4443), .B(n4442), .Z(n4450) );
  XNOR U4627 ( .A(opcode[0]), .B(opcode[2]), .Z(n4445) );
  XNOR U4628 ( .A(opcode[2]), .B(opcode[1]), .Z(n4444) );
  NAND U4629 ( .A(n4445), .B(n4444), .Z(n5597) );
  AND U4630 ( .A(opcode[2]), .B(n1603), .Z(n5594) );
  NAND U4631 ( .A(\stack[1][31] ), .B(n5594), .Z(n4446) );
  NAND U4632 ( .A(n5597), .B(n4446), .Z(n4447) );
  AND U4633 ( .A(o[31]), .B(n4447), .Z(n4448) );
  NANDN U4634 ( .A(n4450), .B(n4449), .Z(n1076) );
  NAND U4635 ( .A(\stack[6][30] ), .B(n5603), .Z(n4452) );
  NANDN U4636 ( .A(n5603), .B(\stack[7][30] ), .Z(n4451) );
  NAND U4637 ( .A(n4452), .B(n4451), .Z(n1077) );
  NAND U4638 ( .A(\stack[5][30] ), .B(n5603), .Z(n4454) );
  NANDN U4639 ( .A(n5588), .B(\stack[7][30] ), .Z(n4453) );
  AND U4640 ( .A(n4454), .B(n4453), .Z(n4456) );
  NAND U4641 ( .A(n5591), .B(\stack[6][30] ), .Z(n4455) );
  NAND U4642 ( .A(n4456), .B(n4455), .Z(n1078) );
  NAND U4643 ( .A(\stack[4][30] ), .B(n5603), .Z(n4458) );
  NANDN U4644 ( .A(n5588), .B(\stack[6][30] ), .Z(n4457) );
  AND U4645 ( .A(n4458), .B(n4457), .Z(n4460) );
  NAND U4646 ( .A(n5591), .B(\stack[5][30] ), .Z(n4459) );
  NAND U4647 ( .A(n4460), .B(n4459), .Z(n1079) );
  NAND U4648 ( .A(\stack[3][30] ), .B(n5603), .Z(n4462) );
  NANDN U4649 ( .A(n5588), .B(\stack[5][30] ), .Z(n4461) );
  AND U4650 ( .A(n4462), .B(n4461), .Z(n4464) );
  NAND U4651 ( .A(n5591), .B(\stack[4][30] ), .Z(n4463) );
  NAND U4652 ( .A(n4464), .B(n4463), .Z(n1080) );
  NAND U4653 ( .A(\stack[2][30] ), .B(n5603), .Z(n4466) );
  NANDN U4654 ( .A(n5588), .B(\stack[4][30] ), .Z(n4465) );
  AND U4655 ( .A(n4466), .B(n4465), .Z(n4468) );
  NAND U4656 ( .A(n5591), .B(\stack[3][30] ), .Z(n4467) );
  NAND U4657 ( .A(n4468), .B(n4467), .Z(n1081) );
  NAND U4658 ( .A(n5603), .B(\stack[1][30] ), .Z(n4470) );
  NANDN U4659 ( .A(n5588), .B(\stack[3][30] ), .Z(n4469) );
  AND U4660 ( .A(n4470), .B(n4469), .Z(n4472) );
  NAND U4661 ( .A(n5591), .B(\stack[2][30] ), .Z(n4471) );
  NAND U4662 ( .A(n4472), .B(n4471), .Z(n1082) );
  NAND U4663 ( .A(n5603), .B(o[30]), .Z(n4474) );
  NANDN U4664 ( .A(n5588), .B(\stack[2][30] ), .Z(n4473) );
  AND U4665 ( .A(n4474), .B(n4473), .Z(n4476) );
  NAND U4666 ( .A(\stack[1][30] ), .B(n5591), .Z(n4475) );
  NAND U4667 ( .A(n4476), .B(n4475), .Z(n1083) );
  NAND U4668 ( .A(o[30]), .B(n5594), .Z(n4477) );
  NANDN U4669 ( .A(n5598), .B(n4477), .Z(n4478) );
  AND U4670 ( .A(\stack[1][30] ), .B(n4478), .Z(n4486) );
  NAND U4671 ( .A(x[30]), .B(n5603), .Z(n4479) );
  XNOR U4672 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U4673 ( .A(n5578), .B(n4482), .Z(n4483) );
  NAND U4674 ( .A(n4484), .B(n4483), .Z(n4485) );
  NOR U4675 ( .A(n4486), .B(n4485), .Z(n4488) );
  NANDN U4676 ( .A(n5597), .B(o[30]), .Z(n4487) );
  NAND U4677 ( .A(n4488), .B(n4487), .Z(n1084) );
  NAND U4678 ( .A(\stack[6][29] ), .B(n5603), .Z(n4490) );
  NANDN U4679 ( .A(n5603), .B(\stack[7][29] ), .Z(n4489) );
  NAND U4680 ( .A(n4490), .B(n4489), .Z(n1085) );
  NAND U4681 ( .A(\stack[5][29] ), .B(n5603), .Z(n4492) );
  NANDN U4682 ( .A(n5588), .B(\stack[7][29] ), .Z(n4491) );
  AND U4683 ( .A(n4492), .B(n4491), .Z(n4494) );
  NAND U4684 ( .A(n5591), .B(\stack[6][29] ), .Z(n4493) );
  NAND U4685 ( .A(n4494), .B(n4493), .Z(n1086) );
  NAND U4686 ( .A(\stack[4][29] ), .B(n5603), .Z(n4496) );
  NANDN U4687 ( .A(n5588), .B(\stack[6][29] ), .Z(n4495) );
  AND U4688 ( .A(n4496), .B(n4495), .Z(n4498) );
  NAND U4689 ( .A(n5591), .B(\stack[5][29] ), .Z(n4497) );
  NAND U4690 ( .A(n4498), .B(n4497), .Z(n1087) );
  NAND U4691 ( .A(\stack[3][29] ), .B(n5603), .Z(n4500) );
  NANDN U4692 ( .A(n5588), .B(\stack[5][29] ), .Z(n4499) );
  AND U4693 ( .A(n4500), .B(n4499), .Z(n4502) );
  NAND U4694 ( .A(n5591), .B(\stack[4][29] ), .Z(n4501) );
  NAND U4695 ( .A(n4502), .B(n4501), .Z(n1088) );
  NAND U4696 ( .A(\stack[2][29] ), .B(n5603), .Z(n4504) );
  NANDN U4697 ( .A(n5588), .B(\stack[4][29] ), .Z(n4503) );
  AND U4698 ( .A(n4504), .B(n4503), .Z(n4506) );
  NAND U4699 ( .A(n5591), .B(\stack[3][29] ), .Z(n4505) );
  NAND U4700 ( .A(n4506), .B(n4505), .Z(n1089) );
  NAND U4701 ( .A(n5603), .B(\stack[1][29] ), .Z(n4508) );
  NANDN U4702 ( .A(n5588), .B(\stack[3][29] ), .Z(n4507) );
  AND U4703 ( .A(n4508), .B(n4507), .Z(n4510) );
  NAND U4704 ( .A(n5591), .B(\stack[2][29] ), .Z(n4509) );
  NAND U4705 ( .A(n4510), .B(n4509), .Z(n1090) );
  NAND U4706 ( .A(n5603), .B(o[29]), .Z(n4512) );
  NANDN U4707 ( .A(n5588), .B(\stack[2][29] ), .Z(n4511) );
  AND U4708 ( .A(n4512), .B(n4511), .Z(n4514) );
  NAND U4709 ( .A(\stack[1][29] ), .B(n5591), .Z(n4513) );
  NAND U4710 ( .A(n4514), .B(n4513), .Z(n1091) );
  NAND U4711 ( .A(x[29]), .B(n5603), .Z(n4516) );
  NAND U4712 ( .A(\stack[1][29] ), .B(n5598), .Z(n4515) );
  AND U4713 ( .A(n4516), .B(n4515), .Z(n4521) );
  XNOR U4714 ( .A(n4518), .B(n4517), .Z(n4519) );
  NAND U4715 ( .A(n5578), .B(n4519), .Z(n4520) );
  NAND U4716 ( .A(n4521), .B(n4520), .Z(n4526) );
  NAND U4717 ( .A(\stack[1][29] ), .B(n5594), .Z(n4522) );
  NAND U4718 ( .A(n5597), .B(n4522), .Z(n4523) );
  AND U4719 ( .A(o[29]), .B(n4523), .Z(n4524) );
  NANDN U4720 ( .A(n4526), .B(n4525), .Z(n1092) );
  NAND U4721 ( .A(\stack[6][28] ), .B(n5603), .Z(n4528) );
  NANDN U4722 ( .A(n5603), .B(\stack[7][28] ), .Z(n4527) );
  NAND U4723 ( .A(n4528), .B(n4527), .Z(n1093) );
  NAND U4724 ( .A(\stack[5][28] ), .B(n5603), .Z(n4530) );
  NANDN U4725 ( .A(n5588), .B(\stack[7][28] ), .Z(n4529) );
  AND U4726 ( .A(n4530), .B(n4529), .Z(n4532) );
  NAND U4727 ( .A(n5591), .B(\stack[6][28] ), .Z(n4531) );
  NAND U4728 ( .A(n4532), .B(n4531), .Z(n1094) );
  NAND U4729 ( .A(\stack[4][28] ), .B(n5603), .Z(n4534) );
  NANDN U4730 ( .A(n5588), .B(\stack[6][28] ), .Z(n4533) );
  AND U4731 ( .A(n4534), .B(n4533), .Z(n4536) );
  NAND U4732 ( .A(n5591), .B(\stack[5][28] ), .Z(n4535) );
  NAND U4733 ( .A(n4536), .B(n4535), .Z(n1095) );
  NAND U4734 ( .A(\stack[3][28] ), .B(n5603), .Z(n4538) );
  NANDN U4735 ( .A(n5588), .B(\stack[5][28] ), .Z(n4537) );
  AND U4736 ( .A(n4538), .B(n4537), .Z(n4540) );
  NAND U4737 ( .A(n5591), .B(\stack[4][28] ), .Z(n4539) );
  NAND U4738 ( .A(n4540), .B(n4539), .Z(n1096) );
  NAND U4739 ( .A(\stack[2][28] ), .B(n5603), .Z(n4542) );
  NANDN U4740 ( .A(n5588), .B(\stack[4][28] ), .Z(n4541) );
  AND U4741 ( .A(n4542), .B(n4541), .Z(n4544) );
  NAND U4742 ( .A(n5591), .B(\stack[3][28] ), .Z(n4543) );
  NAND U4743 ( .A(n4544), .B(n4543), .Z(n1097) );
  NAND U4744 ( .A(n5603), .B(\stack[1][28] ), .Z(n4546) );
  NANDN U4745 ( .A(n5588), .B(\stack[3][28] ), .Z(n4545) );
  AND U4746 ( .A(n4546), .B(n4545), .Z(n4548) );
  NAND U4747 ( .A(n5591), .B(\stack[2][28] ), .Z(n4547) );
  NAND U4748 ( .A(n4548), .B(n4547), .Z(n1098) );
  NAND U4749 ( .A(n5603), .B(o[28]), .Z(n4550) );
  NANDN U4750 ( .A(n5588), .B(\stack[2][28] ), .Z(n4549) );
  AND U4751 ( .A(n4550), .B(n4549), .Z(n4552) );
  NAND U4752 ( .A(\stack[1][28] ), .B(n5591), .Z(n4551) );
  NAND U4753 ( .A(n4552), .B(n4551), .Z(n1099) );
  NAND U4754 ( .A(o[28]), .B(n5594), .Z(n4553) );
  NANDN U4755 ( .A(n5598), .B(n4553), .Z(n4554) );
  AND U4756 ( .A(\stack[1][28] ), .B(n4554), .Z(n4562) );
  NAND U4757 ( .A(x[28]), .B(n5603), .Z(n4555) );
  XNOR U4758 ( .A(n4557), .B(n4556), .Z(n4558) );
  NAND U4759 ( .A(n5578), .B(n4558), .Z(n4559) );
  NAND U4760 ( .A(n4560), .B(n4559), .Z(n4561) );
  NOR U4761 ( .A(n4562), .B(n4561), .Z(n4564) );
  NANDN U4762 ( .A(n5597), .B(o[28]), .Z(n4563) );
  NAND U4763 ( .A(n4564), .B(n4563), .Z(n1100) );
  NAND U4764 ( .A(\stack[6][27] ), .B(n5603), .Z(n4566) );
  NANDN U4765 ( .A(n5603), .B(\stack[7][27] ), .Z(n4565) );
  NAND U4766 ( .A(n4566), .B(n4565), .Z(n1101) );
  NAND U4767 ( .A(\stack[5][27] ), .B(n5603), .Z(n4568) );
  NANDN U4768 ( .A(n5588), .B(\stack[7][27] ), .Z(n4567) );
  AND U4769 ( .A(n4568), .B(n4567), .Z(n4570) );
  NAND U4770 ( .A(n5591), .B(\stack[6][27] ), .Z(n4569) );
  NAND U4771 ( .A(n4570), .B(n4569), .Z(n1102) );
  NAND U4772 ( .A(\stack[4][27] ), .B(n5603), .Z(n4572) );
  NANDN U4773 ( .A(n5588), .B(\stack[6][27] ), .Z(n4571) );
  AND U4774 ( .A(n4572), .B(n4571), .Z(n4574) );
  NAND U4775 ( .A(n5591), .B(\stack[5][27] ), .Z(n4573) );
  NAND U4776 ( .A(n4574), .B(n4573), .Z(n1103) );
  NAND U4777 ( .A(\stack[3][27] ), .B(n5603), .Z(n4576) );
  NANDN U4778 ( .A(n5588), .B(\stack[5][27] ), .Z(n4575) );
  AND U4779 ( .A(n4576), .B(n4575), .Z(n4578) );
  NAND U4780 ( .A(n5591), .B(\stack[4][27] ), .Z(n4577) );
  NAND U4781 ( .A(n4578), .B(n4577), .Z(n1104) );
  NAND U4782 ( .A(\stack[2][27] ), .B(n5603), .Z(n4580) );
  NANDN U4783 ( .A(n5588), .B(\stack[4][27] ), .Z(n4579) );
  AND U4784 ( .A(n4580), .B(n4579), .Z(n4582) );
  NAND U4785 ( .A(n5591), .B(\stack[3][27] ), .Z(n4581) );
  NAND U4786 ( .A(n4582), .B(n4581), .Z(n1105) );
  NAND U4787 ( .A(n5603), .B(\stack[1][27] ), .Z(n4584) );
  NANDN U4788 ( .A(n5588), .B(\stack[3][27] ), .Z(n4583) );
  AND U4789 ( .A(n4584), .B(n4583), .Z(n4586) );
  NAND U4790 ( .A(n5591), .B(\stack[2][27] ), .Z(n4585) );
  NAND U4791 ( .A(n4586), .B(n4585), .Z(n1106) );
  NAND U4792 ( .A(n5603), .B(o[27]), .Z(n4588) );
  NANDN U4793 ( .A(n5588), .B(\stack[2][27] ), .Z(n4587) );
  AND U4794 ( .A(n4588), .B(n4587), .Z(n4590) );
  NAND U4795 ( .A(\stack[1][27] ), .B(n5591), .Z(n4589) );
  NAND U4796 ( .A(n4590), .B(n4589), .Z(n1107) );
  NAND U4797 ( .A(x[27]), .B(n5603), .Z(n4592) );
  NAND U4798 ( .A(\stack[1][27] ), .B(n5598), .Z(n4591) );
  AND U4799 ( .A(n4592), .B(n4591), .Z(n4597) );
  XNOR U4800 ( .A(n4594), .B(n4593), .Z(n4595) );
  NAND U4801 ( .A(n5578), .B(n4595), .Z(n4596) );
  NAND U4802 ( .A(n4597), .B(n4596), .Z(n4602) );
  NAND U4803 ( .A(\stack[1][27] ), .B(n5594), .Z(n4598) );
  NAND U4804 ( .A(n5597), .B(n4598), .Z(n4599) );
  AND U4805 ( .A(o[27]), .B(n4599), .Z(n4600) );
  NANDN U4806 ( .A(n4602), .B(n4601), .Z(n1108) );
  NAND U4807 ( .A(\stack[6][26] ), .B(n5603), .Z(n4604) );
  NANDN U4808 ( .A(n5603), .B(\stack[7][26] ), .Z(n4603) );
  NAND U4809 ( .A(n4604), .B(n4603), .Z(n1109) );
  NAND U4810 ( .A(\stack[5][26] ), .B(n5603), .Z(n4606) );
  NANDN U4811 ( .A(n5588), .B(\stack[7][26] ), .Z(n4605) );
  AND U4812 ( .A(n4606), .B(n4605), .Z(n4608) );
  NAND U4813 ( .A(n5591), .B(\stack[6][26] ), .Z(n4607) );
  NAND U4814 ( .A(n4608), .B(n4607), .Z(n1110) );
  NAND U4815 ( .A(\stack[4][26] ), .B(n5603), .Z(n4610) );
  NANDN U4816 ( .A(n5588), .B(\stack[6][26] ), .Z(n4609) );
  AND U4817 ( .A(n4610), .B(n4609), .Z(n4612) );
  NAND U4818 ( .A(n5591), .B(\stack[5][26] ), .Z(n4611) );
  NAND U4819 ( .A(n4612), .B(n4611), .Z(n1111) );
  NAND U4820 ( .A(\stack[3][26] ), .B(n5603), .Z(n4614) );
  NANDN U4821 ( .A(n5588), .B(\stack[5][26] ), .Z(n4613) );
  AND U4822 ( .A(n4614), .B(n4613), .Z(n4616) );
  NAND U4823 ( .A(n5591), .B(\stack[4][26] ), .Z(n4615) );
  NAND U4824 ( .A(n4616), .B(n4615), .Z(n1112) );
  NAND U4825 ( .A(\stack[2][26] ), .B(n5603), .Z(n4618) );
  NANDN U4826 ( .A(n5588), .B(\stack[4][26] ), .Z(n4617) );
  AND U4827 ( .A(n4618), .B(n4617), .Z(n4620) );
  NAND U4828 ( .A(n5591), .B(\stack[3][26] ), .Z(n4619) );
  NAND U4829 ( .A(n4620), .B(n4619), .Z(n1113) );
  NAND U4830 ( .A(n5603), .B(\stack[1][26] ), .Z(n4622) );
  NANDN U4831 ( .A(n5588), .B(\stack[3][26] ), .Z(n4621) );
  AND U4832 ( .A(n4622), .B(n4621), .Z(n4624) );
  NAND U4833 ( .A(n5591), .B(\stack[2][26] ), .Z(n4623) );
  NAND U4834 ( .A(n4624), .B(n4623), .Z(n1114) );
  NAND U4835 ( .A(n5603), .B(o[26]), .Z(n4626) );
  NANDN U4836 ( .A(n5588), .B(\stack[2][26] ), .Z(n4625) );
  AND U4837 ( .A(n4626), .B(n4625), .Z(n4628) );
  NAND U4838 ( .A(\stack[1][26] ), .B(n5591), .Z(n4627) );
  NAND U4839 ( .A(n4628), .B(n4627), .Z(n1115) );
  NAND U4840 ( .A(o[26]), .B(n5594), .Z(n4629) );
  NANDN U4841 ( .A(n5598), .B(n4629), .Z(n4630) );
  AND U4842 ( .A(\stack[1][26] ), .B(n4630), .Z(n4638) );
  NAND U4843 ( .A(x[26]), .B(n5603), .Z(n4631) );
  XNOR U4844 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U4845 ( .A(n5578), .B(n4634), .Z(n4635) );
  NAND U4846 ( .A(n4636), .B(n4635), .Z(n4637) );
  NOR U4847 ( .A(n4638), .B(n4637), .Z(n4640) );
  NANDN U4848 ( .A(n5597), .B(o[26]), .Z(n4639) );
  NAND U4849 ( .A(n4640), .B(n4639), .Z(n1116) );
  NAND U4850 ( .A(\stack[6][25] ), .B(n5603), .Z(n4642) );
  NANDN U4851 ( .A(n5603), .B(\stack[7][25] ), .Z(n4641) );
  NAND U4852 ( .A(n4642), .B(n4641), .Z(n1117) );
  NAND U4853 ( .A(\stack[5][25] ), .B(n5603), .Z(n4644) );
  NANDN U4854 ( .A(n5588), .B(\stack[7][25] ), .Z(n4643) );
  AND U4855 ( .A(n4644), .B(n4643), .Z(n4646) );
  NAND U4856 ( .A(n5591), .B(\stack[6][25] ), .Z(n4645) );
  NAND U4857 ( .A(n4646), .B(n4645), .Z(n1118) );
  NAND U4858 ( .A(\stack[4][25] ), .B(n5603), .Z(n4648) );
  NANDN U4859 ( .A(n5588), .B(\stack[6][25] ), .Z(n4647) );
  AND U4860 ( .A(n4648), .B(n4647), .Z(n4650) );
  NAND U4861 ( .A(n5591), .B(\stack[5][25] ), .Z(n4649) );
  NAND U4862 ( .A(n4650), .B(n4649), .Z(n1119) );
  NAND U4863 ( .A(\stack[3][25] ), .B(n5603), .Z(n4652) );
  NANDN U4864 ( .A(n5588), .B(\stack[5][25] ), .Z(n4651) );
  AND U4865 ( .A(n4652), .B(n4651), .Z(n4654) );
  NAND U4866 ( .A(n5591), .B(\stack[4][25] ), .Z(n4653) );
  NAND U4867 ( .A(n4654), .B(n4653), .Z(n1120) );
  NAND U4868 ( .A(\stack[2][25] ), .B(n5603), .Z(n4656) );
  NANDN U4869 ( .A(n5588), .B(\stack[4][25] ), .Z(n4655) );
  AND U4870 ( .A(n4656), .B(n4655), .Z(n4658) );
  NAND U4871 ( .A(n5591), .B(\stack[3][25] ), .Z(n4657) );
  NAND U4872 ( .A(n4658), .B(n4657), .Z(n1121) );
  NAND U4873 ( .A(n5603), .B(\stack[1][25] ), .Z(n4660) );
  NANDN U4874 ( .A(n5588), .B(\stack[3][25] ), .Z(n4659) );
  AND U4875 ( .A(n4660), .B(n4659), .Z(n4662) );
  NAND U4876 ( .A(n5591), .B(\stack[2][25] ), .Z(n4661) );
  NAND U4877 ( .A(n4662), .B(n4661), .Z(n1122) );
  NAND U4878 ( .A(n5603), .B(o[25]), .Z(n4664) );
  NANDN U4879 ( .A(n5588), .B(\stack[2][25] ), .Z(n4663) );
  AND U4880 ( .A(n4664), .B(n4663), .Z(n4666) );
  NAND U4881 ( .A(\stack[1][25] ), .B(n5591), .Z(n4665) );
  NAND U4882 ( .A(n4666), .B(n4665), .Z(n1123) );
  NAND U4883 ( .A(x[25]), .B(n5603), .Z(n4668) );
  NAND U4884 ( .A(\stack[1][25] ), .B(n5598), .Z(n4667) );
  AND U4885 ( .A(n4668), .B(n4667), .Z(n4673) );
  XNOR U4886 ( .A(n4670), .B(n4669), .Z(n4671) );
  NAND U4887 ( .A(n5578), .B(n4671), .Z(n4672) );
  NAND U4888 ( .A(n4673), .B(n4672), .Z(n4678) );
  NAND U4889 ( .A(\stack[1][25] ), .B(n5594), .Z(n4674) );
  NAND U4890 ( .A(n5597), .B(n4674), .Z(n4675) );
  AND U4891 ( .A(o[25]), .B(n4675), .Z(n4676) );
  NANDN U4892 ( .A(n4678), .B(n4677), .Z(n1124) );
  NAND U4893 ( .A(\stack[6][24] ), .B(n5603), .Z(n4680) );
  NANDN U4894 ( .A(n5603), .B(\stack[7][24] ), .Z(n4679) );
  NAND U4895 ( .A(n4680), .B(n4679), .Z(n1125) );
  NAND U4896 ( .A(\stack[5][24] ), .B(n5603), .Z(n4682) );
  NANDN U4897 ( .A(n5588), .B(\stack[7][24] ), .Z(n4681) );
  AND U4898 ( .A(n4682), .B(n4681), .Z(n4684) );
  NAND U4899 ( .A(n5591), .B(\stack[6][24] ), .Z(n4683) );
  NAND U4900 ( .A(n4684), .B(n4683), .Z(n1126) );
  NAND U4901 ( .A(\stack[4][24] ), .B(n5603), .Z(n4686) );
  NANDN U4902 ( .A(n5588), .B(\stack[6][24] ), .Z(n4685) );
  AND U4903 ( .A(n4686), .B(n4685), .Z(n4688) );
  NAND U4904 ( .A(n5591), .B(\stack[5][24] ), .Z(n4687) );
  NAND U4905 ( .A(n4688), .B(n4687), .Z(n1127) );
  NAND U4906 ( .A(\stack[3][24] ), .B(n5603), .Z(n4690) );
  NANDN U4907 ( .A(n5588), .B(\stack[5][24] ), .Z(n4689) );
  AND U4908 ( .A(n4690), .B(n4689), .Z(n4692) );
  NAND U4909 ( .A(n5591), .B(\stack[4][24] ), .Z(n4691) );
  NAND U4910 ( .A(n4692), .B(n4691), .Z(n1128) );
  NAND U4911 ( .A(\stack[2][24] ), .B(n5603), .Z(n4694) );
  NANDN U4912 ( .A(n5588), .B(\stack[4][24] ), .Z(n4693) );
  AND U4913 ( .A(n4694), .B(n4693), .Z(n4696) );
  NAND U4914 ( .A(n5591), .B(\stack[3][24] ), .Z(n4695) );
  NAND U4915 ( .A(n4696), .B(n4695), .Z(n1129) );
  NAND U4916 ( .A(n5603), .B(\stack[1][24] ), .Z(n4698) );
  NANDN U4917 ( .A(n5588), .B(\stack[3][24] ), .Z(n4697) );
  AND U4918 ( .A(n4698), .B(n4697), .Z(n4700) );
  NAND U4919 ( .A(n5591), .B(\stack[2][24] ), .Z(n4699) );
  NAND U4920 ( .A(n4700), .B(n4699), .Z(n1130) );
  NAND U4921 ( .A(n5603), .B(o[24]), .Z(n4702) );
  NANDN U4922 ( .A(n5588), .B(\stack[2][24] ), .Z(n4701) );
  AND U4923 ( .A(n4702), .B(n4701), .Z(n4704) );
  NAND U4924 ( .A(\stack[1][24] ), .B(n5591), .Z(n4703) );
  NAND U4925 ( .A(n4704), .B(n4703), .Z(n1131) );
  NAND U4926 ( .A(o[24]), .B(n5594), .Z(n4705) );
  NANDN U4927 ( .A(n5598), .B(n4705), .Z(n4706) );
  AND U4928 ( .A(\stack[1][24] ), .B(n4706), .Z(n4714) );
  NAND U4929 ( .A(x[24]), .B(n5603), .Z(n4707) );
  XNOR U4930 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U4931 ( .A(n5578), .B(n4710), .Z(n4711) );
  NAND U4932 ( .A(n4712), .B(n4711), .Z(n4713) );
  NOR U4933 ( .A(n4714), .B(n4713), .Z(n4716) );
  NANDN U4934 ( .A(n5597), .B(o[24]), .Z(n4715) );
  NAND U4935 ( .A(n4716), .B(n4715), .Z(n1132) );
  NAND U4936 ( .A(\stack[6][23] ), .B(n5603), .Z(n4718) );
  NANDN U4937 ( .A(n5603), .B(\stack[7][23] ), .Z(n4717) );
  NAND U4938 ( .A(n4718), .B(n4717), .Z(n1133) );
  NAND U4939 ( .A(\stack[5][23] ), .B(n5603), .Z(n4720) );
  NANDN U4940 ( .A(n5588), .B(\stack[7][23] ), .Z(n4719) );
  AND U4941 ( .A(n4720), .B(n4719), .Z(n4722) );
  NAND U4942 ( .A(n5591), .B(\stack[6][23] ), .Z(n4721) );
  NAND U4943 ( .A(n4722), .B(n4721), .Z(n1134) );
  NAND U4944 ( .A(\stack[4][23] ), .B(n5603), .Z(n4724) );
  NANDN U4945 ( .A(n5588), .B(\stack[6][23] ), .Z(n4723) );
  AND U4946 ( .A(n4724), .B(n4723), .Z(n4726) );
  NAND U4947 ( .A(n5591), .B(\stack[5][23] ), .Z(n4725) );
  NAND U4948 ( .A(n4726), .B(n4725), .Z(n1135) );
  NAND U4949 ( .A(\stack[3][23] ), .B(n5603), .Z(n4728) );
  NANDN U4950 ( .A(n5588), .B(\stack[5][23] ), .Z(n4727) );
  AND U4951 ( .A(n4728), .B(n4727), .Z(n4730) );
  NAND U4952 ( .A(n5591), .B(\stack[4][23] ), .Z(n4729) );
  NAND U4953 ( .A(n4730), .B(n4729), .Z(n1136) );
  NAND U4954 ( .A(\stack[2][23] ), .B(n5603), .Z(n4732) );
  NANDN U4955 ( .A(n5588), .B(\stack[4][23] ), .Z(n4731) );
  AND U4956 ( .A(n4732), .B(n4731), .Z(n4734) );
  NAND U4957 ( .A(n5591), .B(\stack[3][23] ), .Z(n4733) );
  NAND U4958 ( .A(n4734), .B(n4733), .Z(n1137) );
  NAND U4959 ( .A(n5603), .B(\stack[1][23] ), .Z(n4736) );
  NANDN U4960 ( .A(n5588), .B(\stack[3][23] ), .Z(n4735) );
  AND U4961 ( .A(n4736), .B(n4735), .Z(n4738) );
  NAND U4962 ( .A(n5591), .B(\stack[2][23] ), .Z(n4737) );
  NAND U4963 ( .A(n4738), .B(n4737), .Z(n1138) );
  NAND U4964 ( .A(n5603), .B(o[23]), .Z(n4740) );
  NANDN U4965 ( .A(n5588), .B(\stack[2][23] ), .Z(n4739) );
  AND U4966 ( .A(n4740), .B(n4739), .Z(n4742) );
  NAND U4967 ( .A(\stack[1][23] ), .B(n5591), .Z(n4741) );
  NAND U4968 ( .A(n4742), .B(n4741), .Z(n1139) );
  NAND U4969 ( .A(x[23]), .B(n5603), .Z(n4744) );
  NAND U4970 ( .A(\stack[1][23] ), .B(n5598), .Z(n4743) );
  AND U4971 ( .A(n4744), .B(n4743), .Z(n4749) );
  XNOR U4972 ( .A(n4746), .B(n4745), .Z(n4747) );
  NAND U4973 ( .A(n5578), .B(n4747), .Z(n4748) );
  NAND U4974 ( .A(n4749), .B(n4748), .Z(n4754) );
  NAND U4975 ( .A(\stack[1][23] ), .B(n5594), .Z(n4750) );
  NAND U4976 ( .A(n5597), .B(n4750), .Z(n4751) );
  AND U4977 ( .A(o[23]), .B(n4751), .Z(n4752) );
  NANDN U4978 ( .A(n4754), .B(n4753), .Z(n1140) );
  NAND U4979 ( .A(\stack[6][22] ), .B(n5603), .Z(n4756) );
  NANDN U4980 ( .A(n5603), .B(\stack[7][22] ), .Z(n4755) );
  NAND U4981 ( .A(n4756), .B(n4755), .Z(n1141) );
  NAND U4982 ( .A(\stack[5][22] ), .B(n5603), .Z(n4758) );
  NANDN U4983 ( .A(n5588), .B(\stack[7][22] ), .Z(n4757) );
  AND U4984 ( .A(n4758), .B(n4757), .Z(n4760) );
  NAND U4985 ( .A(n5591), .B(\stack[6][22] ), .Z(n4759) );
  NAND U4986 ( .A(n4760), .B(n4759), .Z(n1142) );
  NAND U4987 ( .A(\stack[4][22] ), .B(n5603), .Z(n4762) );
  NANDN U4988 ( .A(n5588), .B(\stack[6][22] ), .Z(n4761) );
  AND U4989 ( .A(n4762), .B(n4761), .Z(n4764) );
  NAND U4990 ( .A(n5591), .B(\stack[5][22] ), .Z(n4763) );
  NAND U4991 ( .A(n4764), .B(n4763), .Z(n1143) );
  NAND U4992 ( .A(\stack[3][22] ), .B(n5603), .Z(n4766) );
  NANDN U4993 ( .A(n5588), .B(\stack[5][22] ), .Z(n4765) );
  AND U4994 ( .A(n4766), .B(n4765), .Z(n4768) );
  NAND U4995 ( .A(n5591), .B(\stack[4][22] ), .Z(n4767) );
  NAND U4996 ( .A(n4768), .B(n4767), .Z(n1144) );
  NAND U4997 ( .A(\stack[2][22] ), .B(n5603), .Z(n4770) );
  NANDN U4998 ( .A(n5588), .B(\stack[4][22] ), .Z(n4769) );
  AND U4999 ( .A(n4770), .B(n4769), .Z(n4772) );
  NAND U5000 ( .A(n5591), .B(\stack[3][22] ), .Z(n4771) );
  NAND U5001 ( .A(n4772), .B(n4771), .Z(n1145) );
  NAND U5002 ( .A(n5603), .B(\stack[1][22] ), .Z(n4774) );
  NANDN U5003 ( .A(n5588), .B(\stack[3][22] ), .Z(n4773) );
  AND U5004 ( .A(n4774), .B(n4773), .Z(n4776) );
  NAND U5005 ( .A(n5591), .B(\stack[2][22] ), .Z(n4775) );
  NAND U5006 ( .A(n4776), .B(n4775), .Z(n1146) );
  NAND U5007 ( .A(n5603), .B(o[22]), .Z(n4778) );
  NANDN U5008 ( .A(n5588), .B(\stack[2][22] ), .Z(n4777) );
  AND U5009 ( .A(n4778), .B(n4777), .Z(n4780) );
  NAND U5010 ( .A(\stack[1][22] ), .B(n5591), .Z(n4779) );
  NAND U5011 ( .A(n4780), .B(n4779), .Z(n1147) );
  NAND U5012 ( .A(o[22]), .B(n5594), .Z(n4781) );
  NANDN U5013 ( .A(n5598), .B(n4781), .Z(n4782) );
  AND U5014 ( .A(\stack[1][22] ), .B(n4782), .Z(n4790) );
  NAND U5015 ( .A(x[22]), .B(n5603), .Z(n4783) );
  XNOR U5016 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U5017 ( .A(n5578), .B(n4786), .Z(n4787) );
  NAND U5018 ( .A(n4788), .B(n4787), .Z(n4789) );
  NOR U5019 ( .A(n4790), .B(n4789), .Z(n4792) );
  NANDN U5020 ( .A(n5597), .B(o[22]), .Z(n4791) );
  NAND U5021 ( .A(n4792), .B(n4791), .Z(n1148) );
  NAND U5022 ( .A(\stack[6][21] ), .B(n5603), .Z(n4794) );
  NANDN U5023 ( .A(n5603), .B(\stack[7][21] ), .Z(n4793) );
  NAND U5024 ( .A(n4794), .B(n4793), .Z(n1149) );
  NAND U5025 ( .A(\stack[5][21] ), .B(n5603), .Z(n4796) );
  NANDN U5026 ( .A(n5588), .B(\stack[7][21] ), .Z(n4795) );
  AND U5027 ( .A(n4796), .B(n4795), .Z(n4798) );
  NAND U5028 ( .A(n5591), .B(\stack[6][21] ), .Z(n4797) );
  NAND U5029 ( .A(n4798), .B(n4797), .Z(n1150) );
  NAND U5030 ( .A(\stack[4][21] ), .B(n5603), .Z(n4800) );
  NANDN U5031 ( .A(n5588), .B(\stack[6][21] ), .Z(n4799) );
  AND U5032 ( .A(n4800), .B(n4799), .Z(n4802) );
  NAND U5033 ( .A(n5591), .B(\stack[5][21] ), .Z(n4801) );
  NAND U5034 ( .A(n4802), .B(n4801), .Z(n1151) );
  NAND U5035 ( .A(\stack[3][21] ), .B(n5603), .Z(n4804) );
  NANDN U5036 ( .A(n5588), .B(\stack[5][21] ), .Z(n4803) );
  AND U5037 ( .A(n4804), .B(n4803), .Z(n4806) );
  NAND U5038 ( .A(n5591), .B(\stack[4][21] ), .Z(n4805) );
  NAND U5039 ( .A(n4806), .B(n4805), .Z(n1152) );
  NAND U5040 ( .A(\stack[2][21] ), .B(n5603), .Z(n4808) );
  NANDN U5041 ( .A(n5588), .B(\stack[4][21] ), .Z(n4807) );
  AND U5042 ( .A(n4808), .B(n4807), .Z(n4810) );
  NAND U5043 ( .A(n5591), .B(\stack[3][21] ), .Z(n4809) );
  NAND U5044 ( .A(n4810), .B(n4809), .Z(n1153) );
  NAND U5045 ( .A(n5603), .B(\stack[1][21] ), .Z(n4812) );
  NANDN U5046 ( .A(n5588), .B(\stack[3][21] ), .Z(n4811) );
  AND U5047 ( .A(n4812), .B(n4811), .Z(n4814) );
  NAND U5048 ( .A(n5591), .B(\stack[2][21] ), .Z(n4813) );
  NAND U5049 ( .A(n4814), .B(n4813), .Z(n1154) );
  NAND U5050 ( .A(n5603), .B(o[21]), .Z(n4816) );
  NANDN U5051 ( .A(n5588), .B(\stack[2][21] ), .Z(n4815) );
  AND U5052 ( .A(n4816), .B(n4815), .Z(n4818) );
  NAND U5053 ( .A(\stack[1][21] ), .B(n5591), .Z(n4817) );
  NAND U5054 ( .A(n4818), .B(n4817), .Z(n1155) );
  NAND U5055 ( .A(x[21]), .B(n5603), .Z(n4820) );
  NAND U5056 ( .A(\stack[1][21] ), .B(n5598), .Z(n4819) );
  AND U5057 ( .A(n4820), .B(n4819), .Z(n4825) );
  XNOR U5058 ( .A(n4822), .B(n4821), .Z(n4823) );
  NAND U5059 ( .A(n5578), .B(n4823), .Z(n4824) );
  NAND U5060 ( .A(n4825), .B(n4824), .Z(n4830) );
  NAND U5061 ( .A(\stack[1][21] ), .B(n5594), .Z(n4826) );
  NAND U5062 ( .A(n5597), .B(n4826), .Z(n4827) );
  AND U5063 ( .A(o[21]), .B(n4827), .Z(n4828) );
  NANDN U5064 ( .A(n4830), .B(n4829), .Z(n1156) );
  NAND U5065 ( .A(\stack[6][20] ), .B(n5603), .Z(n4832) );
  NANDN U5066 ( .A(n5603), .B(\stack[7][20] ), .Z(n4831) );
  NAND U5067 ( .A(n4832), .B(n4831), .Z(n1157) );
  NAND U5068 ( .A(\stack[5][20] ), .B(n5603), .Z(n4834) );
  NANDN U5069 ( .A(n5588), .B(\stack[7][20] ), .Z(n4833) );
  AND U5070 ( .A(n4834), .B(n4833), .Z(n4836) );
  NAND U5071 ( .A(n5591), .B(\stack[6][20] ), .Z(n4835) );
  NAND U5072 ( .A(n4836), .B(n4835), .Z(n1158) );
  NAND U5073 ( .A(\stack[4][20] ), .B(n5603), .Z(n4838) );
  NANDN U5074 ( .A(n5588), .B(\stack[6][20] ), .Z(n4837) );
  AND U5075 ( .A(n4838), .B(n4837), .Z(n4840) );
  NAND U5076 ( .A(n5591), .B(\stack[5][20] ), .Z(n4839) );
  NAND U5077 ( .A(n4840), .B(n4839), .Z(n1159) );
  NAND U5078 ( .A(\stack[3][20] ), .B(n5603), .Z(n4842) );
  NANDN U5079 ( .A(n5588), .B(\stack[5][20] ), .Z(n4841) );
  AND U5080 ( .A(n4842), .B(n4841), .Z(n4844) );
  NAND U5081 ( .A(n5591), .B(\stack[4][20] ), .Z(n4843) );
  NAND U5082 ( .A(n4844), .B(n4843), .Z(n1160) );
  NAND U5083 ( .A(\stack[2][20] ), .B(n5603), .Z(n4846) );
  NANDN U5084 ( .A(n5588), .B(\stack[4][20] ), .Z(n4845) );
  AND U5085 ( .A(n4846), .B(n4845), .Z(n4848) );
  NAND U5086 ( .A(n5591), .B(\stack[3][20] ), .Z(n4847) );
  NAND U5087 ( .A(n4848), .B(n4847), .Z(n1161) );
  NAND U5088 ( .A(n5603), .B(\stack[1][20] ), .Z(n4850) );
  NANDN U5089 ( .A(n5588), .B(\stack[3][20] ), .Z(n4849) );
  AND U5090 ( .A(n4850), .B(n4849), .Z(n4852) );
  NAND U5091 ( .A(n5591), .B(\stack[2][20] ), .Z(n4851) );
  NAND U5092 ( .A(n4852), .B(n4851), .Z(n1162) );
  NAND U5093 ( .A(n5603), .B(o[20]), .Z(n4854) );
  NANDN U5094 ( .A(n5588), .B(\stack[2][20] ), .Z(n4853) );
  AND U5095 ( .A(n4854), .B(n4853), .Z(n4856) );
  NAND U5096 ( .A(\stack[1][20] ), .B(n5591), .Z(n4855) );
  NAND U5097 ( .A(n4856), .B(n4855), .Z(n1163) );
  NAND U5098 ( .A(o[20]), .B(n5594), .Z(n4857) );
  NANDN U5099 ( .A(n5598), .B(n4857), .Z(n4858) );
  AND U5100 ( .A(\stack[1][20] ), .B(n4858), .Z(n4866) );
  NAND U5101 ( .A(x[20]), .B(n5603), .Z(n4859) );
  XNOR U5102 ( .A(n4861), .B(n4860), .Z(n4862) );
  NAND U5103 ( .A(n5578), .B(n4862), .Z(n4863) );
  NAND U5104 ( .A(n4864), .B(n4863), .Z(n4865) );
  NOR U5105 ( .A(n4866), .B(n4865), .Z(n4868) );
  NANDN U5106 ( .A(n5597), .B(o[20]), .Z(n4867) );
  NAND U5107 ( .A(n4868), .B(n4867), .Z(n1164) );
  NAND U5108 ( .A(\stack[6][19] ), .B(n5603), .Z(n4870) );
  NANDN U5109 ( .A(n5603), .B(\stack[7][19] ), .Z(n4869) );
  NAND U5110 ( .A(n4870), .B(n4869), .Z(n1165) );
  NAND U5111 ( .A(\stack[5][19] ), .B(n5603), .Z(n4872) );
  NANDN U5112 ( .A(n5588), .B(\stack[7][19] ), .Z(n4871) );
  AND U5113 ( .A(n4872), .B(n4871), .Z(n4874) );
  NAND U5114 ( .A(n5591), .B(\stack[6][19] ), .Z(n4873) );
  NAND U5115 ( .A(n4874), .B(n4873), .Z(n1166) );
  NAND U5116 ( .A(\stack[4][19] ), .B(n5603), .Z(n4876) );
  NANDN U5117 ( .A(n5588), .B(\stack[6][19] ), .Z(n4875) );
  AND U5118 ( .A(n4876), .B(n4875), .Z(n4878) );
  NAND U5119 ( .A(n5591), .B(\stack[5][19] ), .Z(n4877) );
  NAND U5120 ( .A(n4878), .B(n4877), .Z(n1167) );
  NAND U5121 ( .A(\stack[3][19] ), .B(n5603), .Z(n4880) );
  NANDN U5122 ( .A(n5588), .B(\stack[5][19] ), .Z(n4879) );
  AND U5123 ( .A(n4880), .B(n4879), .Z(n4882) );
  NAND U5124 ( .A(n5591), .B(\stack[4][19] ), .Z(n4881) );
  NAND U5125 ( .A(n4882), .B(n4881), .Z(n1168) );
  NAND U5126 ( .A(\stack[2][19] ), .B(n5603), .Z(n4884) );
  NANDN U5127 ( .A(n5588), .B(\stack[4][19] ), .Z(n4883) );
  AND U5128 ( .A(n4884), .B(n4883), .Z(n4886) );
  NAND U5129 ( .A(n5591), .B(\stack[3][19] ), .Z(n4885) );
  NAND U5130 ( .A(n4886), .B(n4885), .Z(n1169) );
  NAND U5131 ( .A(n5603), .B(\stack[1][19] ), .Z(n4888) );
  NANDN U5132 ( .A(n5588), .B(\stack[3][19] ), .Z(n4887) );
  AND U5133 ( .A(n4888), .B(n4887), .Z(n4890) );
  NAND U5134 ( .A(n5591), .B(\stack[2][19] ), .Z(n4889) );
  NAND U5135 ( .A(n4890), .B(n4889), .Z(n1170) );
  NAND U5136 ( .A(n5603), .B(o[19]), .Z(n4892) );
  NANDN U5137 ( .A(n5588), .B(\stack[2][19] ), .Z(n4891) );
  AND U5138 ( .A(n4892), .B(n4891), .Z(n4894) );
  NAND U5139 ( .A(\stack[1][19] ), .B(n5591), .Z(n4893) );
  NAND U5140 ( .A(n4894), .B(n4893), .Z(n1171) );
  NAND U5141 ( .A(x[19]), .B(n5603), .Z(n4896) );
  NAND U5142 ( .A(\stack[1][19] ), .B(n5598), .Z(n4895) );
  AND U5143 ( .A(n4896), .B(n4895), .Z(n4901) );
  XNOR U5144 ( .A(n4898), .B(n4897), .Z(n4899) );
  NAND U5145 ( .A(n5578), .B(n4899), .Z(n4900) );
  NAND U5146 ( .A(n4901), .B(n4900), .Z(n4906) );
  NAND U5147 ( .A(\stack[1][19] ), .B(n5594), .Z(n4902) );
  NAND U5148 ( .A(n5597), .B(n4902), .Z(n4903) );
  AND U5149 ( .A(o[19]), .B(n4903), .Z(n4904) );
  NANDN U5150 ( .A(n4906), .B(n4905), .Z(n1172) );
  NAND U5151 ( .A(\stack[6][18] ), .B(n5603), .Z(n4908) );
  NANDN U5152 ( .A(n5603), .B(\stack[7][18] ), .Z(n4907) );
  NAND U5153 ( .A(n4908), .B(n4907), .Z(n1173) );
  NAND U5154 ( .A(\stack[5][18] ), .B(n5603), .Z(n4910) );
  NANDN U5155 ( .A(n5588), .B(\stack[7][18] ), .Z(n4909) );
  AND U5156 ( .A(n4910), .B(n4909), .Z(n4912) );
  NAND U5157 ( .A(n5591), .B(\stack[6][18] ), .Z(n4911) );
  NAND U5158 ( .A(n4912), .B(n4911), .Z(n1174) );
  NAND U5159 ( .A(\stack[4][18] ), .B(n5603), .Z(n4914) );
  NANDN U5160 ( .A(n5588), .B(\stack[6][18] ), .Z(n4913) );
  AND U5161 ( .A(n4914), .B(n4913), .Z(n4916) );
  NAND U5162 ( .A(n5591), .B(\stack[5][18] ), .Z(n4915) );
  NAND U5163 ( .A(n4916), .B(n4915), .Z(n1175) );
  NAND U5164 ( .A(\stack[3][18] ), .B(n5603), .Z(n4918) );
  NANDN U5165 ( .A(n5588), .B(\stack[5][18] ), .Z(n4917) );
  AND U5166 ( .A(n4918), .B(n4917), .Z(n4920) );
  NAND U5167 ( .A(n5591), .B(\stack[4][18] ), .Z(n4919) );
  NAND U5168 ( .A(n4920), .B(n4919), .Z(n1176) );
  NAND U5169 ( .A(\stack[2][18] ), .B(n5603), .Z(n4922) );
  NANDN U5170 ( .A(n5588), .B(\stack[4][18] ), .Z(n4921) );
  AND U5171 ( .A(n4922), .B(n4921), .Z(n4924) );
  NAND U5172 ( .A(n5591), .B(\stack[3][18] ), .Z(n4923) );
  NAND U5173 ( .A(n4924), .B(n4923), .Z(n1177) );
  NAND U5174 ( .A(n5603), .B(\stack[1][18] ), .Z(n4926) );
  NANDN U5175 ( .A(n5588), .B(\stack[3][18] ), .Z(n4925) );
  AND U5176 ( .A(n4926), .B(n4925), .Z(n4928) );
  NAND U5177 ( .A(n5591), .B(\stack[2][18] ), .Z(n4927) );
  NAND U5178 ( .A(n4928), .B(n4927), .Z(n1178) );
  NAND U5179 ( .A(n5603), .B(o[18]), .Z(n4930) );
  NANDN U5180 ( .A(n5588), .B(\stack[2][18] ), .Z(n4929) );
  AND U5181 ( .A(n4930), .B(n4929), .Z(n4932) );
  NAND U5182 ( .A(\stack[1][18] ), .B(n5591), .Z(n4931) );
  NAND U5183 ( .A(n4932), .B(n4931), .Z(n1179) );
  NAND U5184 ( .A(o[18]), .B(n5594), .Z(n4933) );
  NANDN U5185 ( .A(n5598), .B(n4933), .Z(n4934) );
  AND U5186 ( .A(\stack[1][18] ), .B(n4934), .Z(n4942) );
  NAND U5187 ( .A(x[18]), .B(n5603), .Z(n4935) );
  XNOR U5188 ( .A(n4937), .B(n4936), .Z(n4938) );
  NAND U5189 ( .A(n5578), .B(n4938), .Z(n4939) );
  NAND U5190 ( .A(n4940), .B(n4939), .Z(n4941) );
  NOR U5191 ( .A(n4942), .B(n4941), .Z(n4944) );
  NANDN U5192 ( .A(n5597), .B(o[18]), .Z(n4943) );
  NAND U5193 ( .A(n4944), .B(n4943), .Z(n1180) );
  NAND U5194 ( .A(\stack[6][17] ), .B(n5603), .Z(n4946) );
  NANDN U5195 ( .A(n5603), .B(\stack[7][17] ), .Z(n4945) );
  NAND U5196 ( .A(n4946), .B(n4945), .Z(n1181) );
  NAND U5197 ( .A(\stack[5][17] ), .B(n5603), .Z(n4948) );
  NANDN U5198 ( .A(n5588), .B(\stack[7][17] ), .Z(n4947) );
  AND U5199 ( .A(n4948), .B(n4947), .Z(n4950) );
  NAND U5200 ( .A(n5591), .B(\stack[6][17] ), .Z(n4949) );
  NAND U5201 ( .A(n4950), .B(n4949), .Z(n1182) );
  NAND U5202 ( .A(\stack[4][17] ), .B(n5603), .Z(n4952) );
  NANDN U5203 ( .A(n5588), .B(\stack[6][17] ), .Z(n4951) );
  AND U5204 ( .A(n4952), .B(n4951), .Z(n4954) );
  NAND U5205 ( .A(n5591), .B(\stack[5][17] ), .Z(n4953) );
  NAND U5206 ( .A(n4954), .B(n4953), .Z(n1183) );
  NAND U5207 ( .A(\stack[3][17] ), .B(n5603), .Z(n4956) );
  NANDN U5208 ( .A(n5588), .B(\stack[5][17] ), .Z(n4955) );
  AND U5209 ( .A(n4956), .B(n4955), .Z(n4958) );
  NAND U5210 ( .A(n5591), .B(\stack[4][17] ), .Z(n4957) );
  NAND U5211 ( .A(n4958), .B(n4957), .Z(n1184) );
  NAND U5212 ( .A(\stack[2][17] ), .B(n5603), .Z(n4960) );
  NANDN U5213 ( .A(n5588), .B(\stack[4][17] ), .Z(n4959) );
  AND U5214 ( .A(n4960), .B(n4959), .Z(n4962) );
  NAND U5215 ( .A(n5591), .B(\stack[3][17] ), .Z(n4961) );
  NAND U5216 ( .A(n4962), .B(n4961), .Z(n1185) );
  NAND U5217 ( .A(n5603), .B(\stack[1][17] ), .Z(n4964) );
  NANDN U5218 ( .A(n5588), .B(\stack[3][17] ), .Z(n4963) );
  AND U5219 ( .A(n4964), .B(n4963), .Z(n4966) );
  NAND U5220 ( .A(n5591), .B(\stack[2][17] ), .Z(n4965) );
  NAND U5221 ( .A(n4966), .B(n4965), .Z(n1186) );
  NAND U5222 ( .A(n5603), .B(o[17]), .Z(n4968) );
  NANDN U5223 ( .A(n5588), .B(\stack[2][17] ), .Z(n4967) );
  AND U5224 ( .A(n4968), .B(n4967), .Z(n4970) );
  NAND U5225 ( .A(\stack[1][17] ), .B(n5591), .Z(n4969) );
  NAND U5226 ( .A(n4970), .B(n4969), .Z(n1187) );
  NAND U5227 ( .A(x[17]), .B(n5603), .Z(n4972) );
  NAND U5228 ( .A(\stack[1][17] ), .B(n5598), .Z(n4971) );
  AND U5229 ( .A(n4972), .B(n4971), .Z(n4977) );
  XNOR U5230 ( .A(n4974), .B(n4973), .Z(n4975) );
  NAND U5231 ( .A(n5578), .B(n4975), .Z(n4976) );
  NAND U5232 ( .A(n4977), .B(n4976), .Z(n4982) );
  NAND U5233 ( .A(\stack[1][17] ), .B(n5594), .Z(n4978) );
  NAND U5234 ( .A(n5597), .B(n4978), .Z(n4979) );
  AND U5235 ( .A(o[17]), .B(n4979), .Z(n4980) );
  NANDN U5236 ( .A(n4982), .B(n4981), .Z(n1188) );
  NAND U5237 ( .A(\stack[6][16] ), .B(n5603), .Z(n4984) );
  NANDN U5238 ( .A(n5603), .B(\stack[7][16] ), .Z(n4983) );
  NAND U5239 ( .A(n4984), .B(n4983), .Z(n1189) );
  NAND U5240 ( .A(\stack[5][16] ), .B(n5603), .Z(n4986) );
  NANDN U5241 ( .A(n5588), .B(\stack[7][16] ), .Z(n4985) );
  AND U5242 ( .A(n4986), .B(n4985), .Z(n4988) );
  NAND U5243 ( .A(n5591), .B(\stack[6][16] ), .Z(n4987) );
  NAND U5244 ( .A(n4988), .B(n4987), .Z(n1190) );
  NAND U5245 ( .A(\stack[4][16] ), .B(n5603), .Z(n4990) );
  NANDN U5246 ( .A(n5588), .B(\stack[6][16] ), .Z(n4989) );
  AND U5247 ( .A(n4990), .B(n4989), .Z(n4992) );
  NAND U5248 ( .A(n5591), .B(\stack[5][16] ), .Z(n4991) );
  NAND U5249 ( .A(n4992), .B(n4991), .Z(n1191) );
  NAND U5250 ( .A(\stack[3][16] ), .B(n5603), .Z(n4994) );
  NANDN U5251 ( .A(n5588), .B(\stack[5][16] ), .Z(n4993) );
  AND U5252 ( .A(n4994), .B(n4993), .Z(n4996) );
  NAND U5253 ( .A(n5591), .B(\stack[4][16] ), .Z(n4995) );
  NAND U5254 ( .A(n4996), .B(n4995), .Z(n1192) );
  NAND U5255 ( .A(\stack[2][16] ), .B(n5603), .Z(n4998) );
  NANDN U5256 ( .A(n5588), .B(\stack[4][16] ), .Z(n4997) );
  AND U5257 ( .A(n4998), .B(n4997), .Z(n5000) );
  NAND U5258 ( .A(n5591), .B(\stack[3][16] ), .Z(n4999) );
  NAND U5259 ( .A(n5000), .B(n4999), .Z(n1193) );
  NAND U5260 ( .A(n5603), .B(\stack[1][16] ), .Z(n5002) );
  NANDN U5261 ( .A(n5588), .B(\stack[3][16] ), .Z(n5001) );
  AND U5262 ( .A(n5002), .B(n5001), .Z(n5004) );
  NAND U5263 ( .A(n5591), .B(\stack[2][16] ), .Z(n5003) );
  NAND U5264 ( .A(n5004), .B(n5003), .Z(n1194) );
  NAND U5265 ( .A(n5603), .B(o[16]), .Z(n5006) );
  NANDN U5266 ( .A(n5588), .B(\stack[2][16] ), .Z(n5005) );
  AND U5267 ( .A(n5006), .B(n5005), .Z(n5008) );
  NAND U5268 ( .A(\stack[1][16] ), .B(n5591), .Z(n5007) );
  NAND U5269 ( .A(n5008), .B(n5007), .Z(n1195) );
  NAND U5270 ( .A(o[16]), .B(n5594), .Z(n5009) );
  NANDN U5271 ( .A(n5598), .B(n5009), .Z(n5010) );
  AND U5272 ( .A(\stack[1][16] ), .B(n5010), .Z(n5018) );
  NAND U5273 ( .A(x[16]), .B(n5603), .Z(n5011) );
  XNOR U5274 ( .A(n5013), .B(n5012), .Z(n5014) );
  NAND U5275 ( .A(n5578), .B(n5014), .Z(n5015) );
  NAND U5276 ( .A(n5016), .B(n5015), .Z(n5017) );
  NOR U5277 ( .A(n5018), .B(n5017), .Z(n5020) );
  NANDN U5278 ( .A(n5597), .B(o[16]), .Z(n5019) );
  NAND U5279 ( .A(n5020), .B(n5019), .Z(n1196) );
  NAND U5280 ( .A(\stack[6][15] ), .B(n5603), .Z(n5022) );
  NANDN U5281 ( .A(n5603), .B(\stack[7][15] ), .Z(n5021) );
  NAND U5282 ( .A(n5022), .B(n5021), .Z(n1197) );
  NAND U5283 ( .A(\stack[5][15] ), .B(n5603), .Z(n5024) );
  NANDN U5284 ( .A(n5588), .B(\stack[7][15] ), .Z(n5023) );
  AND U5285 ( .A(n5024), .B(n5023), .Z(n5026) );
  NAND U5286 ( .A(n5591), .B(\stack[6][15] ), .Z(n5025) );
  NAND U5287 ( .A(n5026), .B(n5025), .Z(n1198) );
  NAND U5288 ( .A(\stack[4][15] ), .B(n5603), .Z(n5028) );
  NANDN U5289 ( .A(n5588), .B(\stack[6][15] ), .Z(n5027) );
  AND U5290 ( .A(n5028), .B(n5027), .Z(n5030) );
  NAND U5291 ( .A(n5591), .B(\stack[5][15] ), .Z(n5029) );
  NAND U5292 ( .A(n5030), .B(n5029), .Z(n1199) );
  NAND U5293 ( .A(\stack[3][15] ), .B(n5603), .Z(n5032) );
  NANDN U5294 ( .A(n5588), .B(\stack[5][15] ), .Z(n5031) );
  AND U5295 ( .A(n5032), .B(n5031), .Z(n5034) );
  NAND U5296 ( .A(n5591), .B(\stack[4][15] ), .Z(n5033) );
  NAND U5297 ( .A(n5034), .B(n5033), .Z(n1200) );
  NAND U5298 ( .A(\stack[2][15] ), .B(n5603), .Z(n5036) );
  NANDN U5299 ( .A(n5588), .B(\stack[4][15] ), .Z(n5035) );
  AND U5300 ( .A(n5036), .B(n5035), .Z(n5038) );
  NAND U5301 ( .A(n5591), .B(\stack[3][15] ), .Z(n5037) );
  NAND U5302 ( .A(n5038), .B(n5037), .Z(n1201) );
  NAND U5303 ( .A(n5603), .B(\stack[1][15] ), .Z(n5040) );
  NANDN U5304 ( .A(n5588), .B(\stack[3][15] ), .Z(n5039) );
  AND U5305 ( .A(n5040), .B(n5039), .Z(n5042) );
  NAND U5306 ( .A(n5591), .B(\stack[2][15] ), .Z(n5041) );
  NAND U5307 ( .A(n5042), .B(n5041), .Z(n1202) );
  NAND U5308 ( .A(n5603), .B(o[15]), .Z(n5044) );
  NANDN U5309 ( .A(n5588), .B(\stack[2][15] ), .Z(n5043) );
  AND U5310 ( .A(n5044), .B(n5043), .Z(n5046) );
  NAND U5311 ( .A(\stack[1][15] ), .B(n5591), .Z(n5045) );
  NAND U5312 ( .A(n5046), .B(n5045), .Z(n1203) );
  NAND U5313 ( .A(x[15]), .B(n5603), .Z(n5049) );
  NAND U5314 ( .A(n5047), .B(n5594), .Z(n5048) );
  AND U5315 ( .A(n5049), .B(n5048), .Z(n5054) );
  XNOR U5316 ( .A(n5051), .B(n5050), .Z(n5052) );
  NAND U5317 ( .A(n5578), .B(n5052), .Z(n5053) );
  NAND U5318 ( .A(n5054), .B(n5053), .Z(n5059) );
  NAND U5319 ( .A(\stack[1][15] ), .B(n5598), .Z(n5055) );
  NANDN U5320 ( .A(o[15]), .B(n5055), .Z(n5056) );
  ANDN U5321 ( .B(n5056), .A(n5597), .Z(n5057) );
  NANDN U5322 ( .A(n5059), .B(n5058), .Z(n1204) );
  NAND U5323 ( .A(\stack[6][14] ), .B(n5603), .Z(n5061) );
  NANDN U5324 ( .A(n5603), .B(\stack[7][14] ), .Z(n5060) );
  NAND U5325 ( .A(n5061), .B(n5060), .Z(n1205) );
  NAND U5326 ( .A(\stack[5][14] ), .B(n5603), .Z(n5063) );
  NANDN U5327 ( .A(n5588), .B(\stack[7][14] ), .Z(n5062) );
  AND U5328 ( .A(n5063), .B(n5062), .Z(n5065) );
  NAND U5329 ( .A(n5591), .B(\stack[6][14] ), .Z(n5064) );
  NAND U5330 ( .A(n5065), .B(n5064), .Z(n1206) );
  NAND U5331 ( .A(\stack[4][14] ), .B(n5603), .Z(n5067) );
  NANDN U5332 ( .A(n5588), .B(\stack[6][14] ), .Z(n5066) );
  AND U5333 ( .A(n5067), .B(n5066), .Z(n5069) );
  NAND U5334 ( .A(n5591), .B(\stack[5][14] ), .Z(n5068) );
  NAND U5335 ( .A(n5069), .B(n5068), .Z(n1207) );
  NAND U5336 ( .A(\stack[3][14] ), .B(n5603), .Z(n5071) );
  NANDN U5337 ( .A(n5588), .B(\stack[5][14] ), .Z(n5070) );
  AND U5338 ( .A(n5071), .B(n5070), .Z(n5073) );
  NAND U5339 ( .A(n5591), .B(\stack[4][14] ), .Z(n5072) );
  NAND U5340 ( .A(n5073), .B(n5072), .Z(n1208) );
  NAND U5341 ( .A(\stack[2][14] ), .B(n5603), .Z(n5075) );
  NANDN U5342 ( .A(n5588), .B(\stack[4][14] ), .Z(n5074) );
  AND U5343 ( .A(n5075), .B(n5074), .Z(n5077) );
  NAND U5344 ( .A(n5591), .B(\stack[3][14] ), .Z(n5076) );
  NAND U5345 ( .A(n5077), .B(n5076), .Z(n1209) );
  NAND U5346 ( .A(n5603), .B(\stack[1][14] ), .Z(n5079) );
  NANDN U5347 ( .A(n5588), .B(\stack[3][14] ), .Z(n5078) );
  AND U5348 ( .A(n5079), .B(n5078), .Z(n5081) );
  NAND U5349 ( .A(n5591), .B(\stack[2][14] ), .Z(n5080) );
  NAND U5350 ( .A(n5081), .B(n5080), .Z(n1210) );
  NAND U5351 ( .A(n5603), .B(o[14]), .Z(n5083) );
  NANDN U5352 ( .A(n5588), .B(\stack[2][14] ), .Z(n5082) );
  AND U5353 ( .A(n5083), .B(n5082), .Z(n5085) );
  NAND U5354 ( .A(\stack[1][14] ), .B(n5591), .Z(n5084) );
  NAND U5355 ( .A(n5085), .B(n5084), .Z(n1211) );
  NAND U5356 ( .A(x[14]), .B(n5603), .Z(n5087) );
  NAND U5357 ( .A(\stack[1][14] ), .B(n5598), .Z(n5086) );
  NAND U5358 ( .A(n5087), .B(n5086), .Z(n5096) );
  NANDN U5359 ( .A(n5088), .B(n5594), .Z(n5089) );
  XNOR U5360 ( .A(n5091), .B(n5090), .Z(n5092) );
  NAND U5361 ( .A(n5578), .B(n5092), .Z(n5093) );
  NAND U5362 ( .A(n5094), .B(n5093), .Z(n5095) );
  NOR U5363 ( .A(n5096), .B(n5095), .Z(n5098) );
  NANDN U5364 ( .A(n5597), .B(o[14]), .Z(n5097) );
  NAND U5365 ( .A(n5098), .B(n5097), .Z(n1212) );
  NAND U5366 ( .A(\stack[6][13] ), .B(n5603), .Z(n5100) );
  NANDN U5367 ( .A(n5603), .B(\stack[7][13] ), .Z(n5099) );
  NAND U5368 ( .A(n5100), .B(n5099), .Z(n1213) );
  NAND U5369 ( .A(\stack[5][13] ), .B(n5603), .Z(n5102) );
  NANDN U5370 ( .A(n5588), .B(\stack[7][13] ), .Z(n5101) );
  AND U5371 ( .A(n5102), .B(n5101), .Z(n5104) );
  NAND U5372 ( .A(n5591), .B(\stack[6][13] ), .Z(n5103) );
  NAND U5373 ( .A(n5104), .B(n5103), .Z(n1214) );
  NAND U5374 ( .A(\stack[4][13] ), .B(n5603), .Z(n5106) );
  NANDN U5375 ( .A(n5588), .B(\stack[6][13] ), .Z(n5105) );
  AND U5376 ( .A(n5106), .B(n5105), .Z(n5108) );
  NAND U5377 ( .A(n5591), .B(\stack[5][13] ), .Z(n5107) );
  NAND U5378 ( .A(n5108), .B(n5107), .Z(n1215) );
  NAND U5379 ( .A(\stack[3][13] ), .B(n5603), .Z(n5110) );
  NANDN U5380 ( .A(n5588), .B(\stack[5][13] ), .Z(n5109) );
  AND U5381 ( .A(n5110), .B(n5109), .Z(n5112) );
  NAND U5382 ( .A(n5591), .B(\stack[4][13] ), .Z(n5111) );
  NAND U5383 ( .A(n5112), .B(n5111), .Z(n1216) );
  NAND U5384 ( .A(\stack[2][13] ), .B(n5603), .Z(n5114) );
  NANDN U5385 ( .A(n5588), .B(\stack[4][13] ), .Z(n5113) );
  AND U5386 ( .A(n5114), .B(n5113), .Z(n5116) );
  NAND U5387 ( .A(n5591), .B(\stack[3][13] ), .Z(n5115) );
  NAND U5388 ( .A(n5116), .B(n5115), .Z(n1217) );
  NAND U5389 ( .A(n5603), .B(\stack[1][13] ), .Z(n5118) );
  NANDN U5390 ( .A(n5588), .B(\stack[3][13] ), .Z(n5117) );
  AND U5391 ( .A(n5118), .B(n5117), .Z(n5120) );
  NAND U5392 ( .A(n5591), .B(\stack[2][13] ), .Z(n5119) );
  NAND U5393 ( .A(n5120), .B(n5119), .Z(n1218) );
  NAND U5394 ( .A(n5603), .B(o[13]), .Z(n5122) );
  NANDN U5395 ( .A(n5588), .B(\stack[2][13] ), .Z(n5121) );
  AND U5396 ( .A(n5122), .B(n5121), .Z(n5124) );
  NAND U5397 ( .A(\stack[1][13] ), .B(n5591), .Z(n5123) );
  NAND U5398 ( .A(n5124), .B(n5123), .Z(n1219) );
  NAND U5399 ( .A(o[13]), .B(n5594), .Z(n5125) );
  NANDN U5400 ( .A(n5598), .B(n5125), .Z(n5126) );
  AND U5401 ( .A(\stack[1][13] ), .B(n5126), .Z(n5134) );
  NAND U5402 ( .A(x[13]), .B(n5603), .Z(n5127) );
  XNOR U5403 ( .A(n5129), .B(n5128), .Z(n5130) );
  NAND U5404 ( .A(n5578), .B(n5130), .Z(n5131) );
  NAND U5405 ( .A(n5132), .B(n5131), .Z(n5133) );
  NOR U5406 ( .A(n5134), .B(n5133), .Z(n5136) );
  NANDN U5407 ( .A(n5597), .B(o[13]), .Z(n5135) );
  NAND U5408 ( .A(n5136), .B(n5135), .Z(n1220) );
  NAND U5409 ( .A(\stack[6][12] ), .B(n5603), .Z(n5138) );
  NANDN U5410 ( .A(n5603), .B(\stack[7][12] ), .Z(n5137) );
  NAND U5411 ( .A(n5138), .B(n5137), .Z(n1221) );
  NAND U5412 ( .A(\stack[5][12] ), .B(n5603), .Z(n5140) );
  NANDN U5413 ( .A(n5588), .B(\stack[7][12] ), .Z(n5139) );
  AND U5414 ( .A(n5140), .B(n5139), .Z(n5142) );
  NAND U5415 ( .A(n5591), .B(\stack[6][12] ), .Z(n5141) );
  NAND U5416 ( .A(n5142), .B(n5141), .Z(n1222) );
  NAND U5417 ( .A(\stack[4][12] ), .B(n5603), .Z(n5144) );
  NANDN U5418 ( .A(n5588), .B(\stack[6][12] ), .Z(n5143) );
  AND U5419 ( .A(n5144), .B(n5143), .Z(n5146) );
  NAND U5420 ( .A(n5591), .B(\stack[5][12] ), .Z(n5145) );
  NAND U5421 ( .A(n5146), .B(n5145), .Z(n1223) );
  NAND U5422 ( .A(\stack[3][12] ), .B(n5603), .Z(n5148) );
  NANDN U5423 ( .A(n5588), .B(\stack[5][12] ), .Z(n5147) );
  AND U5424 ( .A(n5148), .B(n5147), .Z(n5150) );
  NAND U5425 ( .A(n5591), .B(\stack[4][12] ), .Z(n5149) );
  NAND U5426 ( .A(n5150), .B(n5149), .Z(n1224) );
  NAND U5427 ( .A(\stack[2][12] ), .B(n5603), .Z(n5152) );
  NANDN U5428 ( .A(n5588), .B(\stack[4][12] ), .Z(n5151) );
  AND U5429 ( .A(n5152), .B(n5151), .Z(n5154) );
  NAND U5430 ( .A(n5591), .B(\stack[3][12] ), .Z(n5153) );
  NAND U5431 ( .A(n5154), .B(n5153), .Z(n1225) );
  NAND U5432 ( .A(n5603), .B(\stack[1][12] ), .Z(n5156) );
  NANDN U5433 ( .A(n5588), .B(\stack[3][12] ), .Z(n5155) );
  AND U5434 ( .A(n5156), .B(n5155), .Z(n5158) );
  NAND U5435 ( .A(n5591), .B(\stack[2][12] ), .Z(n5157) );
  NAND U5436 ( .A(n5158), .B(n5157), .Z(n1226) );
  NAND U5437 ( .A(n5603), .B(o[12]), .Z(n5160) );
  NANDN U5438 ( .A(n5588), .B(\stack[2][12] ), .Z(n5159) );
  AND U5439 ( .A(n5160), .B(n5159), .Z(n5162) );
  NAND U5440 ( .A(\stack[1][12] ), .B(n5591), .Z(n5161) );
  NAND U5441 ( .A(n5162), .B(n5161), .Z(n1227) );
  NAND U5442 ( .A(o[12]), .B(n5594), .Z(n5163) );
  NANDN U5443 ( .A(n5598), .B(n5163), .Z(n5164) );
  AND U5444 ( .A(\stack[1][12] ), .B(n5164), .Z(n5172) );
  NAND U5445 ( .A(x[12]), .B(n5603), .Z(n5165) );
  XNOR U5446 ( .A(n5167), .B(n5166), .Z(n5168) );
  NAND U5447 ( .A(n5578), .B(n5168), .Z(n5169) );
  NAND U5448 ( .A(n5170), .B(n5169), .Z(n5171) );
  NOR U5449 ( .A(n5172), .B(n5171), .Z(n5174) );
  NANDN U5450 ( .A(n5597), .B(o[12]), .Z(n5173) );
  NAND U5451 ( .A(n5174), .B(n5173), .Z(n1228) );
  NAND U5452 ( .A(\stack[6][11] ), .B(n5603), .Z(n5176) );
  NANDN U5453 ( .A(n5603), .B(\stack[7][11] ), .Z(n5175) );
  NAND U5454 ( .A(n5176), .B(n5175), .Z(n1229) );
  NAND U5455 ( .A(\stack[5][11] ), .B(n5603), .Z(n5178) );
  NANDN U5456 ( .A(n5588), .B(\stack[7][11] ), .Z(n5177) );
  AND U5457 ( .A(n5178), .B(n5177), .Z(n5180) );
  NAND U5458 ( .A(n5591), .B(\stack[6][11] ), .Z(n5179) );
  NAND U5459 ( .A(n5180), .B(n5179), .Z(n1230) );
  NAND U5460 ( .A(\stack[4][11] ), .B(n5603), .Z(n5182) );
  NANDN U5461 ( .A(n5588), .B(\stack[6][11] ), .Z(n5181) );
  AND U5462 ( .A(n5182), .B(n5181), .Z(n5184) );
  NAND U5463 ( .A(n5591), .B(\stack[5][11] ), .Z(n5183) );
  NAND U5464 ( .A(n5184), .B(n5183), .Z(n1231) );
  NAND U5465 ( .A(\stack[3][11] ), .B(n5603), .Z(n5186) );
  NANDN U5466 ( .A(n5588), .B(\stack[5][11] ), .Z(n5185) );
  AND U5467 ( .A(n5186), .B(n5185), .Z(n5188) );
  NAND U5468 ( .A(n5591), .B(\stack[4][11] ), .Z(n5187) );
  NAND U5469 ( .A(n5188), .B(n5187), .Z(n1232) );
  NAND U5470 ( .A(\stack[2][11] ), .B(n5603), .Z(n5190) );
  NANDN U5471 ( .A(n5588), .B(\stack[4][11] ), .Z(n5189) );
  AND U5472 ( .A(n5190), .B(n5189), .Z(n5192) );
  NAND U5473 ( .A(n5591), .B(\stack[3][11] ), .Z(n5191) );
  NAND U5474 ( .A(n5192), .B(n5191), .Z(n1233) );
  NAND U5475 ( .A(n5603), .B(\stack[1][11] ), .Z(n5194) );
  NANDN U5476 ( .A(n5588), .B(\stack[3][11] ), .Z(n5193) );
  AND U5477 ( .A(n5194), .B(n5193), .Z(n5196) );
  NAND U5478 ( .A(n5591), .B(\stack[2][11] ), .Z(n5195) );
  NAND U5479 ( .A(n5196), .B(n5195), .Z(n1234) );
  NAND U5480 ( .A(n5603), .B(o[11]), .Z(n5198) );
  NANDN U5481 ( .A(n5588), .B(\stack[2][11] ), .Z(n5197) );
  AND U5482 ( .A(n5198), .B(n5197), .Z(n5200) );
  NAND U5483 ( .A(\stack[1][11] ), .B(n5591), .Z(n5199) );
  NAND U5484 ( .A(n5200), .B(n5199), .Z(n1235) );
  NAND U5485 ( .A(n5594), .B(o[11]), .Z(n5201) );
  NANDN U5486 ( .A(n5598), .B(n5201), .Z(n5202) );
  AND U5487 ( .A(\stack[1][11] ), .B(n5202), .Z(n5210) );
  NAND U5488 ( .A(x[11]), .B(n5603), .Z(n5203) );
  XNOR U5489 ( .A(n5205), .B(n5204), .Z(n5206) );
  NAND U5490 ( .A(n5578), .B(n5206), .Z(n5207) );
  NAND U5491 ( .A(n5208), .B(n5207), .Z(n5209) );
  NOR U5492 ( .A(n5210), .B(n5209), .Z(n5212) );
  NANDN U5493 ( .A(n5597), .B(o[11]), .Z(n5211) );
  NAND U5494 ( .A(n5212), .B(n5211), .Z(n1236) );
  NAND U5495 ( .A(\stack[6][10] ), .B(n5603), .Z(n5214) );
  NANDN U5496 ( .A(n5603), .B(\stack[7][10] ), .Z(n5213) );
  NAND U5497 ( .A(n5214), .B(n5213), .Z(n1237) );
  NAND U5498 ( .A(\stack[5][10] ), .B(n5603), .Z(n5216) );
  NANDN U5499 ( .A(n5588), .B(\stack[7][10] ), .Z(n5215) );
  AND U5500 ( .A(n5216), .B(n5215), .Z(n5218) );
  NAND U5501 ( .A(n5591), .B(\stack[6][10] ), .Z(n5217) );
  NAND U5502 ( .A(n5218), .B(n5217), .Z(n1238) );
  NAND U5503 ( .A(\stack[4][10] ), .B(n5603), .Z(n5220) );
  NANDN U5504 ( .A(n5588), .B(\stack[6][10] ), .Z(n5219) );
  AND U5505 ( .A(n5220), .B(n5219), .Z(n5222) );
  NAND U5506 ( .A(n5591), .B(\stack[5][10] ), .Z(n5221) );
  NAND U5507 ( .A(n5222), .B(n5221), .Z(n1239) );
  NAND U5508 ( .A(\stack[3][10] ), .B(n5603), .Z(n5224) );
  NANDN U5509 ( .A(n5588), .B(\stack[5][10] ), .Z(n5223) );
  AND U5510 ( .A(n5224), .B(n5223), .Z(n5226) );
  NAND U5511 ( .A(n5591), .B(\stack[4][10] ), .Z(n5225) );
  NAND U5512 ( .A(n5226), .B(n5225), .Z(n1240) );
  NAND U5513 ( .A(\stack[2][10] ), .B(n5603), .Z(n5228) );
  NANDN U5514 ( .A(n5588), .B(\stack[4][10] ), .Z(n5227) );
  AND U5515 ( .A(n5228), .B(n5227), .Z(n5230) );
  NAND U5516 ( .A(n5591), .B(\stack[3][10] ), .Z(n5229) );
  NAND U5517 ( .A(n5230), .B(n5229), .Z(n1241) );
  NAND U5518 ( .A(n5603), .B(\stack[1][10] ), .Z(n5232) );
  NANDN U5519 ( .A(n5588), .B(\stack[3][10] ), .Z(n5231) );
  AND U5520 ( .A(n5232), .B(n5231), .Z(n5234) );
  NAND U5521 ( .A(n5591), .B(\stack[2][10] ), .Z(n5233) );
  NAND U5522 ( .A(n5234), .B(n5233), .Z(n1242) );
  NAND U5523 ( .A(n5603), .B(o[10]), .Z(n5236) );
  NANDN U5524 ( .A(n5588), .B(\stack[2][10] ), .Z(n5235) );
  AND U5525 ( .A(n5236), .B(n5235), .Z(n5238) );
  NAND U5526 ( .A(\stack[1][10] ), .B(n5591), .Z(n5237) );
  NAND U5527 ( .A(n5238), .B(n5237), .Z(n1243) );
  NAND U5528 ( .A(n5594), .B(o[10]), .Z(n5239) );
  NANDN U5529 ( .A(n5598), .B(n5239), .Z(n5240) );
  AND U5530 ( .A(\stack[1][10] ), .B(n5240), .Z(n5248) );
  NAND U5531 ( .A(x[10]), .B(n5603), .Z(n5241) );
  XNOR U5532 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5533 ( .A(n5578), .B(n5244), .Z(n5245) );
  NAND U5534 ( .A(n5246), .B(n5245), .Z(n5247) );
  NOR U5535 ( .A(n5248), .B(n5247), .Z(n5250) );
  NANDN U5536 ( .A(n5597), .B(o[10]), .Z(n5249) );
  NAND U5537 ( .A(n5250), .B(n5249), .Z(n1244) );
  NAND U5538 ( .A(\stack[6][9] ), .B(n5603), .Z(n5252) );
  NANDN U5539 ( .A(n5603), .B(\stack[7][9] ), .Z(n5251) );
  NAND U5540 ( .A(n5252), .B(n5251), .Z(n1245) );
  NAND U5541 ( .A(\stack[5][9] ), .B(n5603), .Z(n5254) );
  NANDN U5542 ( .A(n5588), .B(\stack[7][9] ), .Z(n5253) );
  AND U5543 ( .A(n5254), .B(n5253), .Z(n5256) );
  NAND U5544 ( .A(n5591), .B(\stack[6][9] ), .Z(n5255) );
  NAND U5545 ( .A(n5256), .B(n5255), .Z(n1246) );
  NAND U5546 ( .A(\stack[4][9] ), .B(n5603), .Z(n5258) );
  NANDN U5547 ( .A(n5588), .B(\stack[6][9] ), .Z(n5257) );
  AND U5548 ( .A(n5258), .B(n5257), .Z(n5260) );
  NAND U5549 ( .A(n5591), .B(\stack[5][9] ), .Z(n5259) );
  NAND U5550 ( .A(n5260), .B(n5259), .Z(n1247) );
  NAND U5551 ( .A(\stack[3][9] ), .B(n5603), .Z(n5262) );
  NANDN U5552 ( .A(n5588), .B(\stack[5][9] ), .Z(n5261) );
  AND U5553 ( .A(n5262), .B(n5261), .Z(n5264) );
  NAND U5554 ( .A(n5591), .B(\stack[4][9] ), .Z(n5263) );
  NAND U5555 ( .A(n5264), .B(n5263), .Z(n1248) );
  NAND U5556 ( .A(\stack[2][9] ), .B(n5603), .Z(n5266) );
  NANDN U5557 ( .A(n5588), .B(\stack[4][9] ), .Z(n5265) );
  AND U5558 ( .A(n5266), .B(n5265), .Z(n5268) );
  NAND U5559 ( .A(n5591), .B(\stack[3][9] ), .Z(n5267) );
  NAND U5560 ( .A(n5268), .B(n5267), .Z(n1249) );
  NAND U5561 ( .A(n5603), .B(\stack[1][9] ), .Z(n5270) );
  NANDN U5562 ( .A(n5588), .B(\stack[3][9] ), .Z(n5269) );
  AND U5563 ( .A(n5270), .B(n5269), .Z(n5272) );
  NAND U5564 ( .A(n5591), .B(\stack[2][9] ), .Z(n5271) );
  NAND U5565 ( .A(n5272), .B(n5271), .Z(n1250) );
  NAND U5566 ( .A(n5603), .B(o[9]), .Z(n5274) );
  NANDN U5567 ( .A(n5588), .B(\stack[2][9] ), .Z(n5273) );
  AND U5568 ( .A(n5274), .B(n5273), .Z(n5276) );
  NAND U5569 ( .A(\stack[1][9] ), .B(n5591), .Z(n5275) );
  NAND U5570 ( .A(n5276), .B(n5275), .Z(n1251) );
  NAND U5571 ( .A(o[9]), .B(n5594), .Z(n5277) );
  NANDN U5572 ( .A(n5598), .B(n5277), .Z(n5278) );
  AND U5573 ( .A(\stack[1][9] ), .B(n5278), .Z(n5286) );
  NAND U5574 ( .A(x[9]), .B(n5603), .Z(n5279) );
  XNOR U5575 ( .A(n5281), .B(n5280), .Z(n5282) );
  NAND U5576 ( .A(n5578), .B(n5282), .Z(n5283) );
  NAND U5577 ( .A(n5284), .B(n5283), .Z(n5285) );
  NOR U5578 ( .A(n5286), .B(n5285), .Z(n5288) );
  NANDN U5579 ( .A(n5597), .B(o[9]), .Z(n5287) );
  NAND U5580 ( .A(n5288), .B(n5287), .Z(n1252) );
  NAND U5581 ( .A(\stack[6][8] ), .B(n5603), .Z(n5290) );
  NANDN U5582 ( .A(n5603), .B(\stack[7][8] ), .Z(n5289) );
  NAND U5583 ( .A(n5290), .B(n5289), .Z(n1253) );
  NAND U5584 ( .A(\stack[5][8] ), .B(n5603), .Z(n5292) );
  NANDN U5585 ( .A(n5588), .B(\stack[7][8] ), .Z(n5291) );
  AND U5586 ( .A(n5292), .B(n5291), .Z(n5294) );
  NAND U5587 ( .A(n5591), .B(\stack[6][8] ), .Z(n5293) );
  NAND U5588 ( .A(n5294), .B(n5293), .Z(n1254) );
  NAND U5589 ( .A(\stack[4][8] ), .B(n5603), .Z(n5296) );
  NANDN U5590 ( .A(n5588), .B(\stack[6][8] ), .Z(n5295) );
  AND U5591 ( .A(n5296), .B(n5295), .Z(n5298) );
  NAND U5592 ( .A(n5591), .B(\stack[5][8] ), .Z(n5297) );
  NAND U5593 ( .A(n5298), .B(n5297), .Z(n1255) );
  NAND U5594 ( .A(\stack[3][8] ), .B(n5603), .Z(n5300) );
  NANDN U5595 ( .A(n5588), .B(\stack[5][8] ), .Z(n5299) );
  AND U5596 ( .A(n5300), .B(n5299), .Z(n5302) );
  NAND U5597 ( .A(n5591), .B(\stack[4][8] ), .Z(n5301) );
  NAND U5598 ( .A(n5302), .B(n5301), .Z(n1256) );
  NAND U5599 ( .A(\stack[2][8] ), .B(n5603), .Z(n5304) );
  NANDN U5600 ( .A(n5588), .B(\stack[4][8] ), .Z(n5303) );
  AND U5601 ( .A(n5304), .B(n5303), .Z(n5306) );
  NAND U5602 ( .A(n5591), .B(\stack[3][8] ), .Z(n5305) );
  NAND U5603 ( .A(n5306), .B(n5305), .Z(n1257) );
  NAND U5604 ( .A(n5603), .B(\stack[1][8] ), .Z(n5308) );
  NANDN U5605 ( .A(n5588), .B(\stack[3][8] ), .Z(n5307) );
  AND U5606 ( .A(n5308), .B(n5307), .Z(n5310) );
  NAND U5607 ( .A(n5591), .B(\stack[2][8] ), .Z(n5309) );
  NAND U5608 ( .A(n5310), .B(n5309), .Z(n1258) );
  NAND U5609 ( .A(n5603), .B(o[8]), .Z(n5312) );
  NANDN U5610 ( .A(n5588), .B(\stack[2][8] ), .Z(n5311) );
  AND U5611 ( .A(n5312), .B(n5311), .Z(n5314) );
  NAND U5612 ( .A(\stack[1][8] ), .B(n5591), .Z(n5313) );
  NAND U5613 ( .A(n5314), .B(n5313), .Z(n1259) );
  NAND U5614 ( .A(x[8]), .B(n5603), .Z(n5317) );
  NAND U5615 ( .A(n5315), .B(n5594), .Z(n5316) );
  NAND U5616 ( .A(n5317), .B(n5316), .Z(n5325) );
  NAND U5617 ( .A(n5598), .B(\stack[1][8] ), .Z(n5318) );
  XNOR U5618 ( .A(n5320), .B(n5319), .Z(n5321) );
  NAND U5619 ( .A(n5578), .B(n5321), .Z(n5322) );
  NAND U5620 ( .A(n5323), .B(n5322), .Z(n5324) );
  NOR U5621 ( .A(n5325), .B(n5324), .Z(n5327) );
  NANDN U5622 ( .A(n5597), .B(o[8]), .Z(n5326) );
  NAND U5623 ( .A(n5327), .B(n5326), .Z(n1260) );
  NAND U5624 ( .A(\stack[6][7] ), .B(n5603), .Z(n5329) );
  NANDN U5625 ( .A(n5603), .B(\stack[7][7] ), .Z(n5328) );
  NAND U5626 ( .A(n5329), .B(n5328), .Z(n1261) );
  NAND U5627 ( .A(\stack[5][7] ), .B(n5603), .Z(n5331) );
  NANDN U5628 ( .A(n5588), .B(\stack[7][7] ), .Z(n5330) );
  AND U5629 ( .A(n5331), .B(n5330), .Z(n5333) );
  NAND U5630 ( .A(n5591), .B(\stack[6][7] ), .Z(n5332) );
  NAND U5631 ( .A(n5333), .B(n5332), .Z(n1262) );
  NAND U5632 ( .A(\stack[4][7] ), .B(n5603), .Z(n5335) );
  NANDN U5633 ( .A(n5588), .B(\stack[6][7] ), .Z(n5334) );
  AND U5634 ( .A(n5335), .B(n5334), .Z(n5337) );
  NAND U5635 ( .A(n5591), .B(\stack[5][7] ), .Z(n5336) );
  NAND U5636 ( .A(n5337), .B(n5336), .Z(n1263) );
  NAND U5637 ( .A(\stack[3][7] ), .B(n5603), .Z(n5339) );
  NANDN U5638 ( .A(n5588), .B(\stack[5][7] ), .Z(n5338) );
  AND U5639 ( .A(n5339), .B(n5338), .Z(n5341) );
  NAND U5640 ( .A(n5591), .B(\stack[4][7] ), .Z(n5340) );
  NAND U5641 ( .A(n5341), .B(n5340), .Z(n1264) );
  NAND U5642 ( .A(\stack[2][7] ), .B(n5603), .Z(n5343) );
  NANDN U5643 ( .A(n5588), .B(\stack[4][7] ), .Z(n5342) );
  AND U5644 ( .A(n5343), .B(n5342), .Z(n5345) );
  NAND U5645 ( .A(n5591), .B(\stack[3][7] ), .Z(n5344) );
  NAND U5646 ( .A(n5345), .B(n5344), .Z(n1265) );
  NAND U5647 ( .A(n5603), .B(\stack[1][7] ), .Z(n5347) );
  NANDN U5648 ( .A(n5588), .B(\stack[3][7] ), .Z(n5346) );
  AND U5649 ( .A(n5347), .B(n5346), .Z(n5349) );
  NAND U5650 ( .A(n5591), .B(\stack[2][7] ), .Z(n5348) );
  NAND U5651 ( .A(n5349), .B(n5348), .Z(n1266) );
  NAND U5652 ( .A(n5603), .B(o[7]), .Z(n5351) );
  NANDN U5653 ( .A(n5588), .B(\stack[2][7] ), .Z(n5350) );
  AND U5654 ( .A(n5351), .B(n5350), .Z(n5353) );
  NAND U5655 ( .A(\stack[1][7] ), .B(n5591), .Z(n5352) );
  NAND U5656 ( .A(n5353), .B(n5352), .Z(n1267) );
  NAND U5657 ( .A(x[7]), .B(n5603), .Z(n5356) );
  NAND U5658 ( .A(n5354), .B(n5594), .Z(n5355) );
  NAND U5659 ( .A(n5356), .B(n5355), .Z(n5364) );
  NAND U5660 ( .A(n5598), .B(\stack[1][7] ), .Z(n5357) );
  XNOR U5661 ( .A(n5359), .B(n5358), .Z(n5360) );
  NAND U5662 ( .A(n5578), .B(n5360), .Z(n5361) );
  NAND U5663 ( .A(n5362), .B(n5361), .Z(n5363) );
  NOR U5664 ( .A(n5364), .B(n5363), .Z(n5366) );
  NANDN U5665 ( .A(n5597), .B(o[7]), .Z(n5365) );
  NAND U5666 ( .A(n5366), .B(n5365), .Z(n1268) );
  NAND U5667 ( .A(\stack[6][6] ), .B(n5603), .Z(n5368) );
  NANDN U5668 ( .A(n5603), .B(\stack[7][6] ), .Z(n5367) );
  NAND U5669 ( .A(n5368), .B(n5367), .Z(n1269) );
  NAND U5670 ( .A(\stack[5][6] ), .B(n5603), .Z(n5370) );
  NANDN U5671 ( .A(n5588), .B(\stack[7][6] ), .Z(n5369) );
  AND U5672 ( .A(n5370), .B(n5369), .Z(n5372) );
  NAND U5673 ( .A(n5591), .B(\stack[6][6] ), .Z(n5371) );
  NAND U5674 ( .A(n5372), .B(n5371), .Z(n1270) );
  NAND U5675 ( .A(\stack[4][6] ), .B(n5603), .Z(n5374) );
  NANDN U5676 ( .A(n5588), .B(\stack[6][6] ), .Z(n5373) );
  AND U5677 ( .A(n5374), .B(n5373), .Z(n5376) );
  NAND U5678 ( .A(n5591), .B(\stack[5][6] ), .Z(n5375) );
  NAND U5679 ( .A(n5376), .B(n5375), .Z(n1271) );
  NAND U5680 ( .A(\stack[3][6] ), .B(n5603), .Z(n5378) );
  NANDN U5681 ( .A(n5588), .B(\stack[5][6] ), .Z(n5377) );
  AND U5682 ( .A(n5378), .B(n5377), .Z(n5380) );
  NAND U5683 ( .A(n5591), .B(\stack[4][6] ), .Z(n5379) );
  NAND U5684 ( .A(n5380), .B(n5379), .Z(n1272) );
  NAND U5685 ( .A(\stack[2][6] ), .B(n5603), .Z(n5382) );
  NANDN U5686 ( .A(n5588), .B(\stack[4][6] ), .Z(n5381) );
  AND U5687 ( .A(n5382), .B(n5381), .Z(n5384) );
  NAND U5688 ( .A(n5591), .B(\stack[3][6] ), .Z(n5383) );
  NAND U5689 ( .A(n5384), .B(n5383), .Z(n1273) );
  NAND U5690 ( .A(n5603), .B(\stack[1][6] ), .Z(n5386) );
  NANDN U5691 ( .A(n5588), .B(\stack[3][6] ), .Z(n5385) );
  AND U5692 ( .A(n5386), .B(n5385), .Z(n5388) );
  NAND U5693 ( .A(n5591), .B(\stack[2][6] ), .Z(n5387) );
  NAND U5694 ( .A(n5388), .B(n5387), .Z(n1274) );
  NAND U5695 ( .A(n5603), .B(o[6]), .Z(n5390) );
  NANDN U5696 ( .A(n5588), .B(\stack[2][6] ), .Z(n5389) );
  AND U5697 ( .A(n5390), .B(n5389), .Z(n5392) );
  NAND U5698 ( .A(\stack[1][6] ), .B(n5591), .Z(n5391) );
  NAND U5699 ( .A(n5392), .B(n5391), .Z(n1275) );
  NAND U5700 ( .A(x[6]), .B(n5603), .Z(n5394) );
  NAND U5701 ( .A(\stack[1][6] ), .B(n5598), .Z(n5393) );
  NAND U5702 ( .A(n5394), .B(n5393), .Z(n5403) );
  NAND U5703 ( .A(n5594), .B(n5395), .Z(n5396) );
  XNOR U5704 ( .A(n5398), .B(n5397), .Z(n5399) );
  NAND U5705 ( .A(n5578), .B(n5399), .Z(n5400) );
  NAND U5706 ( .A(n5401), .B(n5400), .Z(n5402) );
  NOR U5707 ( .A(n5403), .B(n5402), .Z(n5405) );
  NANDN U5708 ( .A(n5597), .B(o[6]), .Z(n5404) );
  NAND U5709 ( .A(n5405), .B(n5404), .Z(n1276) );
  NAND U5710 ( .A(\stack[6][5] ), .B(n5603), .Z(n5407) );
  NANDN U5711 ( .A(n5603), .B(\stack[7][5] ), .Z(n5406) );
  NAND U5712 ( .A(n5407), .B(n5406), .Z(n1277) );
  NAND U5713 ( .A(\stack[5][5] ), .B(n5603), .Z(n5409) );
  NANDN U5714 ( .A(n5588), .B(\stack[7][5] ), .Z(n5408) );
  AND U5715 ( .A(n5409), .B(n5408), .Z(n5411) );
  NAND U5716 ( .A(n5591), .B(\stack[6][5] ), .Z(n5410) );
  NAND U5717 ( .A(n5411), .B(n5410), .Z(n1278) );
  NAND U5718 ( .A(\stack[4][5] ), .B(n5603), .Z(n5413) );
  NANDN U5719 ( .A(n5588), .B(\stack[6][5] ), .Z(n5412) );
  AND U5720 ( .A(n5413), .B(n5412), .Z(n5415) );
  NAND U5721 ( .A(n5591), .B(\stack[5][5] ), .Z(n5414) );
  NAND U5722 ( .A(n5415), .B(n5414), .Z(n1279) );
  NAND U5723 ( .A(\stack[3][5] ), .B(n5603), .Z(n5417) );
  NANDN U5724 ( .A(n5588), .B(\stack[5][5] ), .Z(n5416) );
  AND U5725 ( .A(n5417), .B(n5416), .Z(n5419) );
  NAND U5726 ( .A(n5591), .B(\stack[4][5] ), .Z(n5418) );
  NAND U5727 ( .A(n5419), .B(n5418), .Z(n1280) );
  NAND U5728 ( .A(\stack[2][5] ), .B(n5603), .Z(n5421) );
  NANDN U5729 ( .A(n5588), .B(\stack[4][5] ), .Z(n5420) );
  AND U5730 ( .A(n5421), .B(n5420), .Z(n5423) );
  NAND U5731 ( .A(n5591), .B(\stack[3][5] ), .Z(n5422) );
  NAND U5732 ( .A(n5423), .B(n5422), .Z(n1281) );
  NAND U5733 ( .A(n5603), .B(\stack[1][5] ), .Z(n5425) );
  NANDN U5734 ( .A(n5588), .B(\stack[3][5] ), .Z(n5424) );
  AND U5735 ( .A(n5425), .B(n5424), .Z(n5427) );
  NAND U5736 ( .A(n5591), .B(\stack[2][5] ), .Z(n5426) );
  NAND U5737 ( .A(n5427), .B(n5426), .Z(n1282) );
  NAND U5738 ( .A(n5603), .B(o[5]), .Z(n5429) );
  NANDN U5739 ( .A(n5588), .B(\stack[2][5] ), .Z(n5428) );
  AND U5740 ( .A(n5429), .B(n5428), .Z(n5431) );
  NAND U5741 ( .A(\stack[1][5] ), .B(n5591), .Z(n5430) );
  NAND U5742 ( .A(n5431), .B(n5430), .Z(n1283) );
  NAND U5743 ( .A(n5594), .B(o[5]), .Z(n5432) );
  NANDN U5744 ( .A(n5598), .B(n5432), .Z(n5433) );
  AND U5745 ( .A(\stack[1][5] ), .B(n5433), .Z(n5441) );
  NAND U5746 ( .A(x[5]), .B(n5603), .Z(n5434) );
  XNOR U5747 ( .A(n5436), .B(n5435), .Z(n5437) );
  NAND U5748 ( .A(n5578), .B(n5437), .Z(n5438) );
  NAND U5749 ( .A(n5439), .B(n5438), .Z(n5440) );
  NOR U5750 ( .A(n5441), .B(n5440), .Z(n5443) );
  NANDN U5751 ( .A(n5597), .B(o[5]), .Z(n5442) );
  NAND U5752 ( .A(n5443), .B(n5442), .Z(n1284) );
  NAND U5753 ( .A(\stack[6][4] ), .B(n5603), .Z(n5445) );
  NANDN U5754 ( .A(n5603), .B(\stack[7][4] ), .Z(n5444) );
  NAND U5755 ( .A(n5445), .B(n5444), .Z(n1285) );
  NAND U5756 ( .A(\stack[5][4] ), .B(n5603), .Z(n5447) );
  NANDN U5757 ( .A(n5588), .B(\stack[7][4] ), .Z(n5446) );
  AND U5758 ( .A(n5447), .B(n5446), .Z(n5449) );
  NAND U5759 ( .A(n5591), .B(\stack[6][4] ), .Z(n5448) );
  NAND U5760 ( .A(n5449), .B(n5448), .Z(n1286) );
  NAND U5761 ( .A(\stack[4][4] ), .B(n5603), .Z(n5451) );
  NANDN U5762 ( .A(n5588), .B(\stack[6][4] ), .Z(n5450) );
  AND U5763 ( .A(n5451), .B(n5450), .Z(n5453) );
  NAND U5764 ( .A(n5591), .B(\stack[5][4] ), .Z(n5452) );
  NAND U5765 ( .A(n5453), .B(n5452), .Z(n1287) );
  NAND U5766 ( .A(\stack[3][4] ), .B(n5603), .Z(n5455) );
  NANDN U5767 ( .A(n5588), .B(\stack[5][4] ), .Z(n5454) );
  AND U5768 ( .A(n5455), .B(n5454), .Z(n5457) );
  NAND U5769 ( .A(n5591), .B(\stack[4][4] ), .Z(n5456) );
  NAND U5770 ( .A(n5457), .B(n5456), .Z(n1288) );
  NAND U5771 ( .A(\stack[2][4] ), .B(n5603), .Z(n5459) );
  NANDN U5772 ( .A(n5588), .B(\stack[4][4] ), .Z(n5458) );
  AND U5773 ( .A(n5459), .B(n5458), .Z(n5461) );
  NAND U5774 ( .A(n5591), .B(\stack[3][4] ), .Z(n5460) );
  NAND U5775 ( .A(n5461), .B(n5460), .Z(n1289) );
  NAND U5776 ( .A(n5603), .B(\stack[1][4] ), .Z(n5463) );
  NANDN U5777 ( .A(n5588), .B(\stack[3][4] ), .Z(n5462) );
  AND U5778 ( .A(n5463), .B(n5462), .Z(n5465) );
  NAND U5779 ( .A(n5591), .B(\stack[2][4] ), .Z(n5464) );
  NAND U5780 ( .A(n5465), .B(n5464), .Z(n1290) );
  NAND U5781 ( .A(n5603), .B(o[4]), .Z(n5467) );
  NANDN U5782 ( .A(n5588), .B(\stack[2][4] ), .Z(n5466) );
  AND U5783 ( .A(n5467), .B(n5466), .Z(n5469) );
  NAND U5784 ( .A(\stack[1][4] ), .B(n5591), .Z(n5468) );
  NAND U5785 ( .A(n5469), .B(n5468), .Z(n1291) );
  NAND U5786 ( .A(n5594), .B(o[4]), .Z(n5470) );
  NANDN U5787 ( .A(n5598), .B(n5470), .Z(n5471) );
  AND U5788 ( .A(\stack[1][4] ), .B(n5471), .Z(n5479) );
  NAND U5789 ( .A(x[4]), .B(n5603), .Z(n5472) );
  XNOR U5790 ( .A(n5474), .B(n5473), .Z(n5475) );
  NAND U5791 ( .A(n5578), .B(n5475), .Z(n5476) );
  NAND U5792 ( .A(n5477), .B(n5476), .Z(n5478) );
  NOR U5793 ( .A(n5479), .B(n5478), .Z(n5481) );
  NANDN U5794 ( .A(n5597), .B(o[4]), .Z(n5480) );
  NAND U5795 ( .A(n5481), .B(n5480), .Z(n1292) );
  NAND U5796 ( .A(\stack[6][3] ), .B(n5603), .Z(n5483) );
  NANDN U5797 ( .A(n5603), .B(\stack[7][3] ), .Z(n5482) );
  NAND U5798 ( .A(n5483), .B(n5482), .Z(n1293) );
  NAND U5799 ( .A(\stack[5][3] ), .B(n5603), .Z(n5485) );
  NANDN U5800 ( .A(n5588), .B(\stack[7][3] ), .Z(n5484) );
  AND U5801 ( .A(n5485), .B(n5484), .Z(n5487) );
  NAND U5802 ( .A(n5591), .B(\stack[6][3] ), .Z(n5486) );
  NAND U5803 ( .A(n5487), .B(n5486), .Z(n1294) );
  NAND U5804 ( .A(\stack[4][3] ), .B(n5603), .Z(n5489) );
  NANDN U5805 ( .A(n5588), .B(\stack[6][3] ), .Z(n5488) );
  AND U5806 ( .A(n5489), .B(n5488), .Z(n5491) );
  NAND U5807 ( .A(n5591), .B(\stack[5][3] ), .Z(n5490) );
  NAND U5808 ( .A(n5491), .B(n5490), .Z(n1295) );
  NAND U5809 ( .A(\stack[3][3] ), .B(n5603), .Z(n5493) );
  NANDN U5810 ( .A(n5588), .B(\stack[5][3] ), .Z(n5492) );
  AND U5811 ( .A(n5493), .B(n5492), .Z(n5495) );
  NAND U5812 ( .A(n5591), .B(\stack[4][3] ), .Z(n5494) );
  NAND U5813 ( .A(n5495), .B(n5494), .Z(n1296) );
  NAND U5814 ( .A(\stack[2][3] ), .B(n5603), .Z(n5497) );
  NANDN U5815 ( .A(n5588), .B(\stack[4][3] ), .Z(n5496) );
  AND U5816 ( .A(n5497), .B(n5496), .Z(n5499) );
  NAND U5817 ( .A(n5591), .B(\stack[3][3] ), .Z(n5498) );
  NAND U5818 ( .A(n5499), .B(n5498), .Z(n1297) );
  NAND U5819 ( .A(n5603), .B(\stack[1][3] ), .Z(n5501) );
  NANDN U5820 ( .A(n5588), .B(\stack[3][3] ), .Z(n5500) );
  AND U5821 ( .A(n5501), .B(n5500), .Z(n5503) );
  NAND U5822 ( .A(n5591), .B(\stack[2][3] ), .Z(n5502) );
  NAND U5823 ( .A(n5503), .B(n5502), .Z(n1298) );
  NAND U5824 ( .A(n5603), .B(o[3]), .Z(n5505) );
  NANDN U5825 ( .A(n5588), .B(\stack[2][3] ), .Z(n5504) );
  AND U5826 ( .A(n5505), .B(n5504), .Z(n5507) );
  NAND U5827 ( .A(\stack[1][3] ), .B(n5591), .Z(n5506) );
  NAND U5828 ( .A(n5507), .B(n5506), .Z(n1299) );
  NAND U5829 ( .A(n5594), .B(o[3]), .Z(n5508) );
  NANDN U5830 ( .A(n5598), .B(n5508), .Z(n5509) );
  AND U5831 ( .A(\stack[1][3] ), .B(n5509), .Z(n5517) );
  NAND U5832 ( .A(x[3]), .B(n5603), .Z(n5510) );
  XNOR U5833 ( .A(n5512), .B(n5511), .Z(n5513) );
  NAND U5834 ( .A(n5578), .B(n5513), .Z(n5514) );
  NAND U5835 ( .A(n5515), .B(n5514), .Z(n5516) );
  NOR U5836 ( .A(n5517), .B(n5516), .Z(n5519) );
  NANDN U5837 ( .A(n5597), .B(o[3]), .Z(n5518) );
  NAND U5838 ( .A(n5519), .B(n5518), .Z(n1300) );
  NAND U5839 ( .A(\stack[6][2] ), .B(n5603), .Z(n5521) );
  NANDN U5840 ( .A(n5603), .B(\stack[7][2] ), .Z(n5520) );
  NAND U5841 ( .A(n5521), .B(n5520), .Z(n1301) );
  NAND U5842 ( .A(\stack[5][2] ), .B(n5603), .Z(n5523) );
  NANDN U5843 ( .A(n5588), .B(\stack[7][2] ), .Z(n5522) );
  AND U5844 ( .A(n5523), .B(n5522), .Z(n5525) );
  NAND U5845 ( .A(n5591), .B(\stack[6][2] ), .Z(n5524) );
  NAND U5846 ( .A(n5525), .B(n5524), .Z(n1302) );
  NAND U5847 ( .A(\stack[4][2] ), .B(n5603), .Z(n5527) );
  NANDN U5848 ( .A(n5588), .B(\stack[6][2] ), .Z(n5526) );
  AND U5849 ( .A(n5527), .B(n5526), .Z(n5529) );
  NAND U5850 ( .A(n5591), .B(\stack[5][2] ), .Z(n5528) );
  NAND U5851 ( .A(n5529), .B(n5528), .Z(n1303) );
  NAND U5852 ( .A(\stack[3][2] ), .B(n5603), .Z(n5531) );
  NANDN U5853 ( .A(n5588), .B(\stack[5][2] ), .Z(n5530) );
  AND U5854 ( .A(n5531), .B(n5530), .Z(n5533) );
  NAND U5855 ( .A(n5591), .B(\stack[4][2] ), .Z(n5532) );
  NAND U5856 ( .A(n5533), .B(n5532), .Z(n1304) );
  NAND U5857 ( .A(\stack[2][2] ), .B(n5603), .Z(n5535) );
  NANDN U5858 ( .A(n5588), .B(\stack[4][2] ), .Z(n5534) );
  AND U5859 ( .A(n5535), .B(n5534), .Z(n5537) );
  NAND U5860 ( .A(n5591), .B(\stack[3][2] ), .Z(n5536) );
  NAND U5861 ( .A(n5537), .B(n5536), .Z(n1305) );
  NAND U5862 ( .A(n5603), .B(\stack[1][2] ), .Z(n5539) );
  NANDN U5863 ( .A(n5588), .B(\stack[3][2] ), .Z(n5538) );
  AND U5864 ( .A(n5539), .B(n5538), .Z(n5541) );
  NAND U5865 ( .A(n5591), .B(\stack[2][2] ), .Z(n5540) );
  NAND U5866 ( .A(n5541), .B(n5540), .Z(n1306) );
  NAND U5867 ( .A(n5603), .B(o[2]), .Z(n5543) );
  NANDN U5868 ( .A(n5588), .B(\stack[2][2] ), .Z(n5542) );
  AND U5869 ( .A(n5543), .B(n5542), .Z(n5545) );
  NAND U5870 ( .A(\stack[1][2] ), .B(n5591), .Z(n5544) );
  NAND U5871 ( .A(n5545), .B(n5544), .Z(n1307) );
  NAND U5872 ( .A(\stack[6][1] ), .B(n5603), .Z(n5549) );
  NANDN U5873 ( .A(n5603), .B(\stack[7][1] ), .Z(n5548) );
  NAND U5874 ( .A(n5549), .B(n5548), .Z(n1309) );
  NAND U5875 ( .A(\stack[5][1] ), .B(n5603), .Z(n5551) );
  NANDN U5876 ( .A(n5588), .B(\stack[7][1] ), .Z(n5550) );
  AND U5877 ( .A(n5551), .B(n5550), .Z(n5553) );
  NAND U5878 ( .A(n5591), .B(\stack[6][1] ), .Z(n5552) );
  NAND U5879 ( .A(n5553), .B(n5552), .Z(n1310) );
  NAND U5880 ( .A(\stack[4][1] ), .B(n5603), .Z(n5555) );
  NANDN U5881 ( .A(n5588), .B(\stack[6][1] ), .Z(n5554) );
  AND U5882 ( .A(n5555), .B(n5554), .Z(n5557) );
  NAND U5883 ( .A(n5591), .B(\stack[5][1] ), .Z(n5556) );
  NAND U5884 ( .A(n5557), .B(n5556), .Z(n1311) );
  NAND U5885 ( .A(\stack[3][1] ), .B(n5603), .Z(n5559) );
  NANDN U5886 ( .A(n5588), .B(\stack[5][1] ), .Z(n5558) );
  AND U5887 ( .A(n5559), .B(n5558), .Z(n5561) );
  NAND U5888 ( .A(n5591), .B(\stack[4][1] ), .Z(n5560) );
  NAND U5889 ( .A(n5561), .B(n5560), .Z(n1312) );
  NAND U5890 ( .A(\stack[2][1] ), .B(n5603), .Z(n5563) );
  NANDN U5891 ( .A(n5588), .B(\stack[4][1] ), .Z(n5562) );
  AND U5892 ( .A(n5563), .B(n5562), .Z(n5565) );
  NAND U5893 ( .A(n5591), .B(\stack[3][1] ), .Z(n5564) );
  NAND U5894 ( .A(n5565), .B(n5564), .Z(n1313) );
  NAND U5895 ( .A(n5603), .B(\stack[1][1] ), .Z(n5567) );
  NANDN U5896 ( .A(n5588), .B(\stack[3][1] ), .Z(n5566) );
  AND U5897 ( .A(n5567), .B(n5566), .Z(n5569) );
  NAND U5898 ( .A(n5591), .B(\stack[2][1] ), .Z(n5568) );
  NAND U5899 ( .A(n5569), .B(n5568), .Z(n1314) );
  NAND U5900 ( .A(n5603), .B(o[1]), .Z(n5571) );
  NANDN U5901 ( .A(n5588), .B(\stack[2][1] ), .Z(n5570) );
  AND U5902 ( .A(n5571), .B(n5570), .Z(n5573) );
  NAND U5903 ( .A(\stack[1][1] ), .B(n5591), .Z(n5572) );
  NAND U5904 ( .A(n5573), .B(n5572), .Z(n1315) );
  NANDN U5905 ( .A(n5597), .B(o[1]), .Z(n5574) );
  XOR U5906 ( .A(n5576), .B(n5575), .Z(n5577) );
  NAND U5907 ( .A(n5578), .B(n5577), .Z(n5583) );
  NAND U5908 ( .A(x[1]), .B(n5603), .Z(n5581) );
  NAND U5909 ( .A(o[1]), .B(\stack[1][1] ), .Z(n5579) );
  NANDN U5910 ( .A(n5579), .B(n5594), .Z(n5580) );
  AND U5911 ( .A(n5581), .B(n5580), .Z(n5582) );
  AND U5912 ( .A(n5583), .B(n5582), .Z(n5585) );
  NAND U5913 ( .A(\stack[1][1] ), .B(n5598), .Z(n5584) );
  AND U5914 ( .A(n5585), .B(n5584), .Z(n5586) );
  NANDN U5915 ( .A(n5587), .B(n5586), .Z(n1316) );
  NAND U5916 ( .A(n5603), .B(o[0]), .Z(n5590) );
  NANDN U5917 ( .A(n5588), .B(\stack[2][0] ), .Z(n5589) );
  AND U5918 ( .A(n5590), .B(n5589), .Z(n5593) );
  NAND U5919 ( .A(\stack[1][0] ), .B(n5591), .Z(n5592) );
  NAND U5920 ( .A(n5593), .B(n5592), .Z(n1317) );
  OR U5921 ( .A(n5595), .B(n5594), .Z(n5596) );
  AND U5922 ( .A(\stack[1][0] ), .B(n5596), .Z(n5599) );
  NANDN U5923 ( .A(n5599), .B(n5597), .Z(n5602) );
  NAND U5924 ( .A(n5599), .B(n5598), .Z(n5600) );
  NANDN U5925 ( .A(o[0]), .B(n5600), .Z(n5601) );
  NAND U5926 ( .A(n5602), .B(n5601), .Z(n5606) );
  NAND U5927 ( .A(x[0]), .B(n5603), .Z(n5604) );
  NAND U5928 ( .A(n5606), .B(n5605), .Z(n1318) );
endmodule

