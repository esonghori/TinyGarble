
module aes_seq_CC10 ( clk, rst, e_init, g_input, o );
  input [127:0] e_init;
  input [127:0] g_input;
  output [127:0] o;
  input clk, rst;
  wire   \w1[0][127] , \w1[0][126] , \w1[0][125] , \w1[0][124] , \w1[0][123] ,
         \w1[0][122] , \w1[0][121] , \w1[0][120] , \w1[0][119] , \w1[0][118] ,
         \w1[0][117] , \w1[0][116] , \w1[0][115] , \w1[0][114] , \w1[0][113] ,
         \w1[0][112] , \w1[0][111] , \w1[0][110] , \w1[0][109] , \w1[0][108] ,
         \w1[0][107] , \w1[0][106] , \w1[0][105] , \w1[0][104] , \w1[0][103] ,
         \w1[0][102] , \w1[0][101] , \w1[0][100] , \w1[0][99] , \w1[0][98] ,
         \w1[0][97] , \w1[0][96] , \w1[0][95] , \w1[0][94] , \w1[0][93] ,
         \w1[0][92] , \w1[0][91] , \w1[0][90] , \w1[0][89] , \w1[0][88] ,
         \w1[0][87] , \w1[0][86] , \w1[0][85] , \w1[0][84] , \w1[0][83] ,
         \w1[0][82] , \w1[0][81] , \w1[0][80] , \w1[0][79] , \w1[0][78] ,
         \w1[0][77] , \w1[0][76] , \w1[0][75] , \w1[0][74] , \w1[0][73] ,
         \w1[0][72] , \w1[0][71] , \w1[0][70] , \w1[0][69] , \w1[0][68] ,
         \w1[0][67] , \w1[0][66] , \w1[0][65] , \w1[0][64] , \w1[0][63] ,
         \w1[0][62] , \w1[0][61] , \w1[0][60] , \w1[0][59] , \w1[0][58] ,
         \w1[0][57] , \w1[0][56] , \w1[0][55] , \w1[0][54] , \w1[0][53] ,
         \w1[0][52] , \w1[0][51] , \w1[0][50] , \w1[0][49] , \w1[0][48] ,
         \w1[0][47] , \w1[0][46] , \w1[0][45] , \w1[0][44] , \w1[0][43] ,
         \w1[0][42] , \w1[0][41] , \w1[0][40] , \w1[0][39] , \w1[0][38] ,
         \w1[0][37] , \w1[0][36] , \w1[0][35] , \w1[0][34] , \w1[0][33] ,
         \w1[0][32] , \w1[0][31] , \w1[0][30] , \w1[0][29] , \w1[0][28] ,
         \w1[0][27] , \w1[0][26] , \w1[0][25] , \w1[0][24] , \w1[0][23] ,
         \w1[0][22] , \w1[0][21] , \w1[0][20] , \w1[0][19] , \w1[0][18] ,
         \w1[0][17] , \w1[0][16] , \w1[0][15] , \w1[0][14] , \w1[0][13] ,
         \w1[0][12] , \w1[0][11] , \w1[0][10] , \w1[0][9] , \w1[0][8] ,
         \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , \w1[0][3] ,
         \w1[0][2] , \w1[0][1] , \w1[0][0] , \SUBBYTES[0].a/n1744 ,
         \SUBBYTES[0].a/n1743 , \SUBBYTES[0].a/n1742 , \SUBBYTES[0].a/n1741 ,
         \SUBBYTES[0].a/n1740 , \SUBBYTES[0].a/n1739 , \SUBBYTES[0].a/n1738 ,
         \SUBBYTES[0].a/n1737 , \SUBBYTES[0].a/n1736 , \SUBBYTES[0].a/n1735 ,
         \SUBBYTES[0].a/n1734 , \SUBBYTES[0].a/n1733 , \SUBBYTES[0].a/n1732 ,
         \SUBBYTES[0].a/n1731 , \SUBBYTES[0].a/n1730 , \SUBBYTES[0].a/n1729 ,
         \SUBBYTES[0].a/n1728 , \SUBBYTES[0].a/n1727 , \SUBBYTES[0].a/n1726 ,
         \SUBBYTES[0].a/n1725 , \SUBBYTES[0].a/n1724 , \SUBBYTES[0].a/n1723 ,
         \SUBBYTES[0].a/n1722 , \SUBBYTES[0].a/n1721 , \SUBBYTES[0].a/n1720 ,
         \SUBBYTES[0].a/n1719 , \SUBBYTES[0].a/n1718 , \SUBBYTES[0].a/n1717 ,
         \SUBBYTES[0].a/n1716 , \SUBBYTES[0].a/n1715 , \SUBBYTES[0].a/n1714 ,
         \SUBBYTES[0].a/n1713 , \SUBBYTES[0].a/n1712 , \SUBBYTES[0].a/n1711 ,
         \SUBBYTES[0].a/n1710 , \SUBBYTES[0].a/n1709 , \SUBBYTES[0].a/n1708 ,
         \SUBBYTES[0].a/n1707 , \SUBBYTES[0].a/n1706 , \SUBBYTES[0].a/n1705 ,
         \SUBBYTES[0].a/n1704 , \SUBBYTES[0].a/n1703 , \SUBBYTES[0].a/n1702 ,
         \SUBBYTES[0].a/n1701 , \SUBBYTES[0].a/n1700 , \SUBBYTES[0].a/n1699 ,
         \SUBBYTES[0].a/n1698 , \SUBBYTES[0].a/n1697 , \SUBBYTES[0].a/n1696 ,
         \SUBBYTES[0].a/n1695 , \SUBBYTES[0].a/n1694 , \SUBBYTES[0].a/n1693 ,
         \SUBBYTES[0].a/n1692 , \SUBBYTES[0].a/n1691 , \SUBBYTES[0].a/n1690 ,
         \SUBBYTES[0].a/n1689 , \SUBBYTES[0].a/n1688 , \SUBBYTES[0].a/n1687 ,
         \SUBBYTES[0].a/n1686 , \SUBBYTES[0].a/n1685 , \SUBBYTES[0].a/n1684 ,
         \SUBBYTES[0].a/n1683 , \SUBBYTES[0].a/n1682 , \SUBBYTES[0].a/n1681 ,
         \SUBBYTES[0].a/n1680 , \SUBBYTES[0].a/n1679 , \SUBBYTES[0].a/n1678 ,
         \SUBBYTES[0].a/n1677 , \SUBBYTES[0].a/n1676 , \SUBBYTES[0].a/n1675 ,
         \SUBBYTES[0].a/n1674 , \SUBBYTES[0].a/n1673 , \SUBBYTES[0].a/n1672 ,
         \SUBBYTES[0].a/n1671 , \SUBBYTES[0].a/n1670 , \SUBBYTES[0].a/n1669 ,
         \SUBBYTES[0].a/n1668 , \SUBBYTES[0].a/n1667 , \SUBBYTES[0].a/n1666 ,
         \SUBBYTES[0].a/n1665 , \SUBBYTES[0].a/n1664 , \SUBBYTES[0].a/n1663 ,
         \SUBBYTES[0].a/n1662 , \SUBBYTES[0].a/n1661 , \SUBBYTES[0].a/n1660 ,
         \SUBBYTES[0].a/n1659 , \SUBBYTES[0].a/n1658 , \SUBBYTES[0].a/n1657 ,
         \SUBBYTES[0].a/n1656 , \SUBBYTES[0].a/n1655 , \SUBBYTES[0].a/n1654 ,
         \SUBBYTES[0].a/n1653 , \SUBBYTES[0].a/n1652 , \SUBBYTES[0].a/n1651 ,
         \SUBBYTES[0].a/n1650 , \SUBBYTES[0].a/n1649 , \SUBBYTES[0].a/n1648 ,
         \SUBBYTES[0].a/n1647 , \SUBBYTES[0].a/n1646 , \SUBBYTES[0].a/n1645 ,
         \SUBBYTES[0].a/n1644 , \SUBBYTES[0].a/n1643 , \SUBBYTES[0].a/n1642 ,
         \SUBBYTES[0].a/n1641 , \SUBBYTES[0].a/n1640 , \SUBBYTES[0].a/n1639 ,
         \SUBBYTES[0].a/n1638 , \SUBBYTES[0].a/n1637 , \SUBBYTES[0].a/n1636 ,
         \SUBBYTES[0].a/n1635 , \SUBBYTES[0].a/n1634 , \SUBBYTES[0].a/n1633 ,
         \SUBBYTES[0].a/n1632 , \SUBBYTES[0].a/n1631 , \SUBBYTES[0].a/n1630 ,
         \SUBBYTES[0].a/n1629 , \SUBBYTES[0].a/n1628 , \SUBBYTES[0].a/n1627 ,
         \SUBBYTES[0].a/n1626 , \SUBBYTES[0].a/n1625 , \SUBBYTES[0].a/n1624 ,
         \SUBBYTES[0].a/n1623 , \SUBBYTES[0].a/n1622 , \SUBBYTES[0].a/n1621 ,
         \SUBBYTES[0].a/n1620 , \SUBBYTES[0].a/n1619 , \SUBBYTES[0].a/n1618 ,
         \SUBBYTES[0].a/n1617 , \SUBBYTES[0].a/n1616 , \SUBBYTES[0].a/n1615 ,
         \SUBBYTES[0].a/n1614 , \SUBBYTES[0].a/n1613 , \SUBBYTES[0].a/n1612 ,
         \SUBBYTES[0].a/n1611 , \SUBBYTES[0].a/n1610 , \SUBBYTES[0].a/n1609 ,
         \SUBBYTES[0].a/n1608 , \SUBBYTES[0].a/n1607 , \SUBBYTES[0].a/n1606 ,
         \SUBBYTES[0].a/n1605 , \SUBBYTES[0].a/n1604 , \SUBBYTES[0].a/n1603 ,
         \SUBBYTES[0].a/n1602 , \SUBBYTES[0].a/n1601 , \SUBBYTES[0].a/n1600 ,
         \SUBBYTES[0].a/n1599 , \SUBBYTES[0].a/n1598 , \SUBBYTES[0].a/n1597 ,
         \SUBBYTES[0].a/n1596 , \SUBBYTES[0].a/n1595 , \SUBBYTES[0].a/n1594 ,
         \SUBBYTES[0].a/n1593 , \SUBBYTES[0].a/n1592 , \SUBBYTES[0].a/n1591 ,
         \SUBBYTES[0].a/n1590 , \SUBBYTES[0].a/n1589 , \SUBBYTES[0].a/n1588 ,
         \SUBBYTES[0].a/n1587 , \SUBBYTES[0].a/n1586 , \SUBBYTES[0].a/n1585 ,
         \SUBBYTES[0].a/n1584 , \SUBBYTES[0].a/n1583 , \SUBBYTES[0].a/n1582 ,
         \SUBBYTES[0].a/n1581 , \SUBBYTES[0].a/n1580 , \SUBBYTES[0].a/n1579 ,
         \SUBBYTES[0].a/n1578 , \SUBBYTES[0].a/n1577 , \SUBBYTES[0].a/n1576 ,
         \SUBBYTES[0].a/n1575 , \SUBBYTES[0].a/n1574 , \SUBBYTES[0].a/n1573 ,
         \SUBBYTES[0].a/n1572 , \SUBBYTES[0].a/n1571 , \SUBBYTES[0].a/n1570 ,
         \SUBBYTES[0].a/n1569 , \SUBBYTES[0].a/n1568 , \SUBBYTES[0].a/n1567 ,
         \SUBBYTES[0].a/n1566 , \SUBBYTES[0].a/n1565 , \SUBBYTES[0].a/n1564 ,
         \SUBBYTES[0].a/n1563 , \SUBBYTES[0].a/n1562 , \SUBBYTES[0].a/n1561 ,
         \SUBBYTES[0].a/n1560 , \SUBBYTES[0].a/n1559 , \SUBBYTES[0].a/n1558 ,
         \SUBBYTES[0].a/n1557 , \SUBBYTES[0].a/n1556 , \SUBBYTES[0].a/n1555 ,
         \SUBBYTES[0].a/n1554 , \SUBBYTES[0].a/n1553 , \SUBBYTES[0].a/n1552 ,
         \SUBBYTES[0].a/n1551 , \SUBBYTES[0].a/n1550 , \SUBBYTES[0].a/n1549 ,
         \SUBBYTES[0].a/n1548 , \SUBBYTES[0].a/n1547 , \SUBBYTES[0].a/n1546 ,
         \SUBBYTES[0].a/n1545 , \SUBBYTES[0].a/n1544 , \SUBBYTES[0].a/n1543 ,
         \SUBBYTES[0].a/n1542 , \SUBBYTES[0].a/n1541 , \SUBBYTES[0].a/n1540 ,
         \SUBBYTES[0].a/n1539 , \SUBBYTES[0].a/n1538 , \SUBBYTES[0].a/n1537 ,
         \SUBBYTES[0].a/n1536 , \SUBBYTES[0].a/n1535 , \SUBBYTES[0].a/n1534 ,
         \SUBBYTES[0].a/n1533 , \SUBBYTES[0].a/n1532 , \SUBBYTES[0].a/n1531 ,
         \SUBBYTES[0].a/n1530 , \SUBBYTES[0].a/n1529 , \SUBBYTES[0].a/n1528 ,
         \SUBBYTES[0].a/n1527 , \SUBBYTES[0].a/n1526 , \SUBBYTES[0].a/n1525 ,
         \SUBBYTES[0].a/n1524 , \SUBBYTES[0].a/n1523 , \SUBBYTES[0].a/n1522 ,
         \SUBBYTES[0].a/n1521 , \SUBBYTES[0].a/n1520 , \SUBBYTES[0].a/n1519 ,
         \SUBBYTES[0].a/n1518 , \SUBBYTES[0].a/n1517 , \SUBBYTES[0].a/n1516 ,
         \SUBBYTES[0].a/n1515 , \SUBBYTES[0].a/n1514 , \SUBBYTES[0].a/n1513 ,
         \SUBBYTES[0].a/n1512 , \SUBBYTES[0].a/n1511 , \SUBBYTES[0].a/n1510 ,
         \SUBBYTES[0].a/n1509 , \SUBBYTES[0].a/n1508 , \SUBBYTES[0].a/n1507 ,
         \SUBBYTES[0].a/n1506 , \SUBBYTES[0].a/n1505 , \SUBBYTES[0].a/n1504 ,
         \SUBBYTES[0].a/n1503 , \SUBBYTES[0].a/n1502 , \SUBBYTES[0].a/n1501 ,
         \SUBBYTES[0].a/n1500 , \SUBBYTES[0].a/n1499 , \SUBBYTES[0].a/n1498 ,
         \SUBBYTES[0].a/n1497 , \SUBBYTES[0].a/n1496 , \SUBBYTES[0].a/n1495 ,
         \SUBBYTES[0].a/n1494 , \SUBBYTES[0].a/n1493 , \SUBBYTES[0].a/n1492 ,
         \SUBBYTES[0].a/n1491 , \SUBBYTES[0].a/n1490 , \SUBBYTES[0].a/n1489 ,
         \SUBBYTES[0].a/n1488 , \SUBBYTES[0].a/n1487 , \SUBBYTES[0].a/n1486 ,
         \SUBBYTES[0].a/n1485 , \SUBBYTES[0].a/n1484 , \SUBBYTES[0].a/n1483 ,
         \SUBBYTES[0].a/n1482 , \SUBBYTES[0].a/n1481 , \SUBBYTES[0].a/n1480 ,
         \SUBBYTES[0].a/n1479 , \SUBBYTES[0].a/n1478 , \SUBBYTES[0].a/n1477 ,
         \SUBBYTES[0].a/n1476 , \SUBBYTES[0].a/n1475 , \SUBBYTES[0].a/n1474 ,
         \SUBBYTES[0].a/n1473 , \SUBBYTES[0].a/n1472 , \SUBBYTES[0].a/n1471 ,
         \SUBBYTES[0].a/n1470 , \SUBBYTES[0].a/n1469 , \SUBBYTES[0].a/n1468 ,
         \SUBBYTES[0].a/n1467 , \SUBBYTES[0].a/n1466 , \SUBBYTES[0].a/n1465 ,
         \SUBBYTES[0].a/n1464 , \SUBBYTES[0].a/n1463 , \SUBBYTES[0].a/n1462 ,
         \SUBBYTES[0].a/n1461 , \SUBBYTES[0].a/n1460 , \SUBBYTES[0].a/n1459 ,
         \SUBBYTES[0].a/n1458 , \SUBBYTES[0].a/n1457 , \SUBBYTES[0].a/n1456 ,
         \SUBBYTES[0].a/n1455 , \SUBBYTES[0].a/n1454 , \SUBBYTES[0].a/n1453 ,
         \SUBBYTES[0].a/n1452 , \SUBBYTES[0].a/n1451 , \SUBBYTES[0].a/n1450 ,
         \SUBBYTES[0].a/n1449 , \SUBBYTES[0].a/n1448 , \SUBBYTES[0].a/n1447 ,
         \SUBBYTES[0].a/n1446 , \SUBBYTES[0].a/n1445 , \SUBBYTES[0].a/n1444 ,
         \SUBBYTES[0].a/n1443 , \SUBBYTES[0].a/n1442 , \SUBBYTES[0].a/n1441 ,
         \SUBBYTES[0].a/n1440 , \SUBBYTES[0].a/n1439 , \SUBBYTES[0].a/n1438 ,
         \SUBBYTES[0].a/n1437 , \SUBBYTES[0].a/n1436 , \SUBBYTES[0].a/n1435 ,
         \SUBBYTES[0].a/n1434 , \SUBBYTES[0].a/n1433 , \SUBBYTES[0].a/n1432 ,
         \SUBBYTES[0].a/n1431 , \SUBBYTES[0].a/n1430 , \SUBBYTES[0].a/n1429 ,
         \SUBBYTES[0].a/n1428 , \SUBBYTES[0].a/n1427 , \SUBBYTES[0].a/n1426 ,
         \SUBBYTES[0].a/n1425 , \SUBBYTES[0].a/n1424 , \SUBBYTES[0].a/n1423 ,
         \SUBBYTES[0].a/n1422 , \SUBBYTES[0].a/n1421 , \SUBBYTES[0].a/n1420 ,
         \SUBBYTES[0].a/n1419 , \SUBBYTES[0].a/n1418 , \SUBBYTES[0].a/n1417 ,
         \SUBBYTES[0].a/n1416 , \SUBBYTES[0].a/n1415 , \SUBBYTES[0].a/n1414 ,
         \SUBBYTES[0].a/n1413 , \SUBBYTES[0].a/n1412 , \SUBBYTES[0].a/n1411 ,
         \SUBBYTES[0].a/n1410 , \SUBBYTES[0].a/n1409 , \SUBBYTES[0].a/n1408 ,
         \SUBBYTES[0].a/n1407 , \SUBBYTES[0].a/n1406 , \SUBBYTES[0].a/n1405 ,
         \SUBBYTES[0].a/n1404 , \SUBBYTES[0].a/n1403 , \SUBBYTES[0].a/n1402 ,
         \SUBBYTES[0].a/n1401 , \SUBBYTES[0].a/n1400 , \SUBBYTES[0].a/n1399 ,
         \SUBBYTES[0].a/n1398 , \SUBBYTES[0].a/n1397 , \SUBBYTES[0].a/n1396 ,
         \SUBBYTES[0].a/n1395 , \SUBBYTES[0].a/n1394 , \SUBBYTES[0].a/n1393 ,
         \SUBBYTES[0].a/n1392 , \SUBBYTES[0].a/n1391 , \SUBBYTES[0].a/n1390 ,
         \SUBBYTES[0].a/n1389 , \SUBBYTES[0].a/n1388 , \SUBBYTES[0].a/n1387 ,
         \SUBBYTES[0].a/n1386 , \SUBBYTES[0].a/n1385 , \SUBBYTES[0].a/n1384 ,
         \SUBBYTES[0].a/n1383 , \SUBBYTES[0].a/n1382 , \SUBBYTES[0].a/n1381 ,
         \SUBBYTES[0].a/n1380 , \SUBBYTES[0].a/n1379 , \SUBBYTES[0].a/n1378 ,
         \SUBBYTES[0].a/n1377 , \SUBBYTES[0].a/n1376 , \SUBBYTES[0].a/n1375 ,
         \SUBBYTES[0].a/n1374 , \SUBBYTES[0].a/n1373 , \SUBBYTES[0].a/n1372 ,
         \SUBBYTES[0].a/n1371 , \SUBBYTES[0].a/n1370 , \SUBBYTES[0].a/n1369 ,
         \SUBBYTES[0].a/n1368 , \SUBBYTES[0].a/n1367 , \SUBBYTES[0].a/n1366 ,
         \SUBBYTES[0].a/n1365 , \SUBBYTES[0].a/n1364 , \SUBBYTES[0].a/n1363 ,
         \SUBBYTES[0].a/n1362 , \SUBBYTES[0].a/n1361 , \SUBBYTES[0].a/n1360 ,
         \SUBBYTES[0].a/n1359 , \SUBBYTES[0].a/n1358 , \SUBBYTES[0].a/n1357 ,
         \SUBBYTES[0].a/n1356 , \SUBBYTES[0].a/n1355 , \SUBBYTES[0].a/n1354 ,
         \SUBBYTES[0].a/n1353 , \SUBBYTES[0].a/n1352 , \SUBBYTES[0].a/n1351 ,
         \SUBBYTES[0].a/n1350 , \SUBBYTES[0].a/n1349 , \SUBBYTES[0].a/n1348 ,
         \SUBBYTES[0].a/n1347 , \SUBBYTES[0].a/n1346 , \SUBBYTES[0].a/n1345 ,
         \SUBBYTES[0].a/n1344 , \SUBBYTES[0].a/n1343 , \SUBBYTES[0].a/n1342 ,
         \SUBBYTES[0].a/n1341 , \SUBBYTES[0].a/n1340 , \SUBBYTES[0].a/n1339 ,
         \SUBBYTES[0].a/n1338 , \SUBBYTES[0].a/n1337 , \SUBBYTES[0].a/n1336 ,
         \SUBBYTES[0].a/n1335 , \SUBBYTES[0].a/n1334 , \SUBBYTES[0].a/n1333 ,
         \SUBBYTES[0].a/n1332 , \SUBBYTES[0].a/n1331 , \SUBBYTES[0].a/n1330 ,
         \SUBBYTES[0].a/n1329 , \SUBBYTES[0].a/n1328 , \SUBBYTES[0].a/n1327 ,
         \SUBBYTES[0].a/n1326 , \SUBBYTES[0].a/n1325 , \SUBBYTES[0].a/n1324 ,
         \SUBBYTES[0].a/n1323 , \SUBBYTES[0].a/n1322 , \SUBBYTES[0].a/n1321 ,
         \SUBBYTES[0].a/n1320 , \SUBBYTES[0].a/n1319 , \SUBBYTES[0].a/n1318 ,
         \SUBBYTES[0].a/n1317 , \SUBBYTES[0].a/n1316 , \SUBBYTES[0].a/n1315 ,
         \SUBBYTES[0].a/n1314 , \SUBBYTES[0].a/n1313 , \SUBBYTES[0].a/n1312 ,
         \SUBBYTES[0].a/n1311 , \SUBBYTES[0].a/n1310 , \SUBBYTES[0].a/n1309 ,
         \SUBBYTES[0].a/n1308 , \SUBBYTES[0].a/n1307 , \SUBBYTES[0].a/n1306 ,
         \SUBBYTES[0].a/n1305 , \SUBBYTES[0].a/n1304 , \SUBBYTES[0].a/n1303 ,
         \SUBBYTES[0].a/n1302 , \SUBBYTES[0].a/n1301 , \SUBBYTES[0].a/n1300 ,
         \SUBBYTES[0].a/n1299 , \SUBBYTES[0].a/n1298 , \SUBBYTES[0].a/n1297 ,
         \SUBBYTES[0].a/n1296 , \SUBBYTES[0].a/n1295 , \SUBBYTES[0].a/n1294 ,
         \SUBBYTES[0].a/n1293 , \SUBBYTES[0].a/n1292 , \SUBBYTES[0].a/n1291 ,
         \SUBBYTES[0].a/n1290 , \SUBBYTES[0].a/n1289 , \SUBBYTES[0].a/n1288 ,
         \SUBBYTES[0].a/n1287 , \SUBBYTES[0].a/n1286 , \SUBBYTES[0].a/n1285 ,
         \SUBBYTES[0].a/n1284 , \SUBBYTES[0].a/n1283 , \SUBBYTES[0].a/n1282 ,
         \SUBBYTES[0].a/n1281 , \SUBBYTES[0].a/n1280 , \SUBBYTES[0].a/n1279 ,
         \SUBBYTES[0].a/n1278 , \SUBBYTES[0].a/n1277 , \SUBBYTES[0].a/n1276 ,
         \SUBBYTES[0].a/n1275 , \SUBBYTES[0].a/n1274 , \SUBBYTES[0].a/n1273 ,
         \SUBBYTES[0].a/n1272 , \SUBBYTES[0].a/n1271 , \SUBBYTES[0].a/n1270 ,
         \SUBBYTES[0].a/n1269 , \SUBBYTES[0].a/n1268 , \SUBBYTES[0].a/n1267 ,
         \SUBBYTES[0].a/n1266 , \SUBBYTES[0].a/n1265 , \SUBBYTES[0].a/n1264 ,
         \SUBBYTES[0].a/n1263 , \SUBBYTES[0].a/n1262 , \SUBBYTES[0].a/n1261 ,
         \SUBBYTES[0].a/n1260 , \SUBBYTES[0].a/n1259 , \SUBBYTES[0].a/n1258 ,
         \SUBBYTES[0].a/n1257 , \SUBBYTES[0].a/n1256 , \SUBBYTES[0].a/n1255 ,
         \SUBBYTES[0].a/n1254 , \SUBBYTES[0].a/n1253 , \SUBBYTES[0].a/n1252 ,
         \SUBBYTES[0].a/n1251 , \SUBBYTES[0].a/n1250 , \SUBBYTES[0].a/n1249 ,
         \SUBBYTES[0].a/n1248 , \SUBBYTES[0].a/n1247 , \SUBBYTES[0].a/n1246 ,
         \SUBBYTES[0].a/n1245 , \SUBBYTES[0].a/n1244 , \SUBBYTES[0].a/n1243 ,
         \SUBBYTES[0].a/n1242 , \SUBBYTES[0].a/n1241 , \SUBBYTES[0].a/n1240 ,
         \SUBBYTES[0].a/n1239 , \SUBBYTES[0].a/n1238 , \SUBBYTES[0].a/n1237 ,
         \SUBBYTES[0].a/n1236 , \SUBBYTES[0].a/n1235 , \SUBBYTES[0].a/n1234 ,
         \SUBBYTES[0].a/n1233 , \SUBBYTES[0].a/n1232 , \SUBBYTES[0].a/n1231 ,
         \SUBBYTES[0].a/n1230 , \SUBBYTES[0].a/n1229 , \SUBBYTES[0].a/n1228 ,
         \SUBBYTES[0].a/n1227 , \SUBBYTES[0].a/n1226 , \SUBBYTES[0].a/n1225 ,
         \SUBBYTES[0].a/n1224 , \SUBBYTES[0].a/n1223 , \SUBBYTES[0].a/n1222 ,
         \SUBBYTES[0].a/n1221 , \SUBBYTES[0].a/n1220 , \SUBBYTES[0].a/n1219 ,
         \SUBBYTES[0].a/n1218 , \SUBBYTES[0].a/n1217 , \SUBBYTES[0].a/n1216 ,
         \SUBBYTES[0].a/n1215 , \SUBBYTES[0].a/n1214 , \SUBBYTES[0].a/n1213 ,
         \SUBBYTES[0].a/n1212 , \SUBBYTES[0].a/n1211 , \SUBBYTES[0].a/n1210 ,
         \SUBBYTES[0].a/n1209 , \SUBBYTES[0].a/n1208 , \SUBBYTES[0].a/n1207 ,
         \SUBBYTES[0].a/n1206 , \SUBBYTES[0].a/n1205 , \SUBBYTES[0].a/n1204 ,
         \SUBBYTES[0].a/n1203 , \SUBBYTES[0].a/n1202 , \SUBBYTES[0].a/n1201 ,
         \SUBBYTES[0].a/n1200 , \SUBBYTES[0].a/n1199 , \SUBBYTES[0].a/n1198 ,
         \SUBBYTES[0].a/n1197 , \SUBBYTES[0].a/n1196 , \SUBBYTES[0].a/n1195 ,
         \SUBBYTES[0].a/n1194 , \SUBBYTES[0].a/n1193 , \SUBBYTES[0].a/n1192 ,
         \SUBBYTES[0].a/n1191 , \SUBBYTES[0].a/n1190 , \SUBBYTES[0].a/n1189 ,
         \SUBBYTES[0].a/n1188 , \SUBBYTES[0].a/n1187 , \SUBBYTES[0].a/n1186 ,
         \SUBBYTES[0].a/n1185 , \SUBBYTES[0].a/n1184 , \SUBBYTES[0].a/n1183 ,
         \SUBBYTES[0].a/n1182 , \SUBBYTES[0].a/n1181 , \SUBBYTES[0].a/n1180 ,
         \SUBBYTES[0].a/n1179 , \SUBBYTES[0].a/n1178 , \SUBBYTES[0].a/n1177 ,
         \SUBBYTES[0].a/n1176 , \SUBBYTES[0].a/n1175 , \SUBBYTES[0].a/n1174 ,
         \SUBBYTES[0].a/n1173 , \SUBBYTES[0].a/n1172 , \SUBBYTES[0].a/n1171 ,
         \SUBBYTES[0].a/n1170 , \SUBBYTES[0].a/n1169 , \SUBBYTES[0].a/n1168 ,
         \SUBBYTES[0].a/n1167 , \SUBBYTES[0].a/n1166 , \SUBBYTES[0].a/n1165 ,
         \SUBBYTES[0].a/n1164 , \SUBBYTES[0].a/n1163 , \SUBBYTES[0].a/n1162 ,
         \SUBBYTES[0].a/n1161 , \SUBBYTES[0].a/n1160 , \SUBBYTES[0].a/n1159 ,
         \SUBBYTES[0].a/n1158 , \SUBBYTES[0].a/n1157 , \SUBBYTES[0].a/n1156 ,
         \SUBBYTES[0].a/n1155 , \SUBBYTES[0].a/n1154 , \SUBBYTES[0].a/n1153 ,
         \SUBBYTES[0].a/n1152 , \SUBBYTES[0].a/n1151 , \SUBBYTES[0].a/n1150 ,
         \SUBBYTES[0].a/n1149 , \SUBBYTES[0].a/n1148 , \SUBBYTES[0].a/n1147 ,
         \SUBBYTES[0].a/n1146 , \SUBBYTES[0].a/n1145 , \SUBBYTES[0].a/n1144 ,
         \SUBBYTES[0].a/n1143 , \SUBBYTES[0].a/n1142 , \SUBBYTES[0].a/n1141 ,
         \SUBBYTES[0].a/n1140 , \SUBBYTES[0].a/n1139 , \SUBBYTES[0].a/n1138 ,
         \SUBBYTES[0].a/n1137 , \SUBBYTES[0].a/n1136 , \SUBBYTES[0].a/n1135 ,
         \SUBBYTES[0].a/n1134 , \SUBBYTES[0].a/n1133 , \SUBBYTES[0].a/n1132 ,
         \SUBBYTES[0].a/n1131 , \SUBBYTES[0].a/n1130 , \SUBBYTES[0].a/n1129 ,
         \SUBBYTES[0].a/n1128 , \SUBBYTES[0].a/n1127 , \SUBBYTES[0].a/n1126 ,
         \SUBBYTES[0].a/n1125 , \SUBBYTES[0].a/n1124 , \SUBBYTES[0].a/n1123 ,
         \SUBBYTES[0].a/n1122 , \SUBBYTES[0].a/n1121 , \SUBBYTES[0].a/n1120 ,
         \SUBBYTES[0].a/n1119 , \SUBBYTES[0].a/n1118 , \SUBBYTES[0].a/n1117 ,
         \SUBBYTES[0].a/n1116 , \SUBBYTES[0].a/n1115 , \SUBBYTES[0].a/n1114 ,
         \SUBBYTES[0].a/n1113 , \SUBBYTES[0].a/n1112 , \SUBBYTES[0].a/n1111 ,
         \SUBBYTES[0].a/n1110 , \SUBBYTES[0].a/n1109 , \SUBBYTES[0].a/n1108 ,
         \SUBBYTES[0].a/n1107 , \SUBBYTES[0].a/n1106 , \SUBBYTES[0].a/n1105 ,
         \SUBBYTES[0].a/n1104 , \SUBBYTES[0].a/n1103 , \SUBBYTES[0].a/n1102 ,
         \SUBBYTES[0].a/n1101 , \SUBBYTES[0].a/n1100 , \SUBBYTES[0].a/n1099 ,
         \SUBBYTES[0].a/n1098 , \SUBBYTES[0].a/n1097 , \SUBBYTES[0].a/n1096 ,
         \SUBBYTES[0].a/n1095 , \SUBBYTES[0].a/n1094 , \SUBBYTES[0].a/n1093 ,
         \SUBBYTES[0].a/n1092 , \SUBBYTES[0].a/n1091 , \SUBBYTES[0].a/n1090 ,
         \SUBBYTES[0].a/n1089 , \SUBBYTES[0].a/n1088 , \SUBBYTES[0].a/n1087 ,
         \SUBBYTES[0].a/n1086 , \SUBBYTES[0].a/n1085 , \SUBBYTES[0].a/n1084 ,
         \SUBBYTES[0].a/n1083 , \SUBBYTES[0].a/n1082 , \SUBBYTES[0].a/n1081 ,
         \SUBBYTES[0].a/n1080 , \SUBBYTES[0].a/n1079 , \SUBBYTES[0].a/n1078 ,
         \SUBBYTES[0].a/n1077 , \SUBBYTES[0].a/n1076 , \SUBBYTES[0].a/n1075 ,
         \SUBBYTES[0].a/n1074 , \SUBBYTES[0].a/n1073 , \SUBBYTES[0].a/n1072 ,
         \SUBBYTES[0].a/n1071 , \SUBBYTES[0].a/n1070 , \SUBBYTES[0].a/n1069 ,
         \SUBBYTES[0].a/n1068 , \SUBBYTES[0].a/n1067 , \SUBBYTES[0].a/n1066 ,
         \SUBBYTES[0].a/n1065 , \SUBBYTES[0].a/n1064 , \SUBBYTES[0].a/n1063 ,
         \SUBBYTES[0].a/n1062 , \SUBBYTES[0].a/n1061 , \SUBBYTES[0].a/n1060 ,
         \SUBBYTES[0].a/n1059 , \SUBBYTES[0].a/n1058 , \SUBBYTES[0].a/n1057 ,
         \SUBBYTES[0].a/n1056 , \SUBBYTES[0].a/n1055 , \SUBBYTES[0].a/n1054 ,
         \SUBBYTES[0].a/n1053 , \SUBBYTES[0].a/n1052 , \SUBBYTES[0].a/n1051 ,
         \SUBBYTES[0].a/n1050 , \SUBBYTES[0].a/n1049 , \SUBBYTES[0].a/n1048 ,
         \SUBBYTES[0].a/n1047 , \SUBBYTES[0].a/n1046 , \SUBBYTES[0].a/n1045 ,
         \SUBBYTES[0].a/n1044 , \SUBBYTES[0].a/n1043 , \SUBBYTES[0].a/n1042 ,
         \SUBBYTES[0].a/n1041 , \SUBBYTES[0].a/n1040 , \SUBBYTES[0].a/n1039 ,
         \SUBBYTES[0].a/n1038 , \SUBBYTES[0].a/n1037 , \SUBBYTES[0].a/n1036 ,
         \SUBBYTES[0].a/n1035 , \SUBBYTES[0].a/n1034 , \SUBBYTES[0].a/n1033 ,
         \SUBBYTES[0].a/n1032 , \SUBBYTES[0].a/n1031 , \SUBBYTES[0].a/n1030 ,
         \SUBBYTES[0].a/n1029 , \SUBBYTES[0].a/n1028 , \SUBBYTES[0].a/n1027 ,
         \SUBBYTES[0].a/n1026 , \SUBBYTES[0].a/n1025 , \SUBBYTES[0].a/n1024 ,
         \SUBBYTES[0].a/n1023 , \SUBBYTES[0].a/n1022 , \SUBBYTES[0].a/n1021 ,
         \SUBBYTES[0].a/n1020 , \SUBBYTES[0].a/n1019 , \SUBBYTES[0].a/n1018 ,
         \SUBBYTES[0].a/n1017 , \SUBBYTES[0].a/n1016 , \SUBBYTES[0].a/n1015 ,
         \SUBBYTES[0].a/n1014 , \SUBBYTES[0].a/n1013 , \SUBBYTES[0].a/n1012 ,
         \SUBBYTES[0].a/n1011 , \SUBBYTES[0].a/n1010 , \SUBBYTES[0].a/n1009 ,
         \SUBBYTES[0].a/n1008 , \SUBBYTES[0].a/n1007 , \SUBBYTES[0].a/n1006 ,
         \SUBBYTES[0].a/n1005 , \SUBBYTES[0].a/n1004 , \SUBBYTES[0].a/n1003 ,
         \SUBBYTES[0].a/n1002 , \SUBBYTES[0].a/n1001 , \SUBBYTES[0].a/n1000 ,
         \SUBBYTES[0].a/n999 , \SUBBYTES[0].a/n998 , \SUBBYTES[0].a/n997 ,
         \SUBBYTES[0].a/n996 , \SUBBYTES[0].a/n995 , \SUBBYTES[0].a/n994 ,
         \SUBBYTES[0].a/n993 , \SUBBYTES[0].a/n992 , \SUBBYTES[0].a/n991 ,
         \SUBBYTES[0].a/n990 , \SUBBYTES[0].a/n989 , \SUBBYTES[0].a/n988 ,
         \SUBBYTES[0].a/n987 , \SUBBYTES[0].a/n986 , \SUBBYTES[0].a/n985 ,
         \SUBBYTES[0].a/n984 , \SUBBYTES[0].a/n983 , \SUBBYTES[0].a/n982 ,
         \SUBBYTES[0].a/n981 , \SUBBYTES[0].a/n980 , \SUBBYTES[0].a/n979 ,
         \SUBBYTES[0].a/n978 , \SUBBYTES[0].a/n977 , \SUBBYTES[0].a/n976 ,
         \SUBBYTES[0].a/n975 , \SUBBYTES[0].a/n974 , \SUBBYTES[0].a/n973 ,
         \SUBBYTES[0].a/n972 , \SUBBYTES[0].a/n971 , \SUBBYTES[0].a/n970 ,
         \SUBBYTES[0].a/n969 , \SUBBYTES[0].a/n968 , \SUBBYTES[0].a/n967 ,
         \SUBBYTES[0].a/n966 , \SUBBYTES[0].a/n965 , \SUBBYTES[0].a/n964 ,
         \SUBBYTES[0].a/n963 , \SUBBYTES[0].a/n962 , \SUBBYTES[0].a/n961 ,
         \SUBBYTES[0].a/n960 , \SUBBYTES[0].a/n959 , \SUBBYTES[0].a/n958 ,
         \SUBBYTES[0].a/n957 , \SUBBYTES[0].a/n956 , \SUBBYTES[0].a/n955 ,
         \SUBBYTES[0].a/n954 , \SUBBYTES[0].a/n953 , \SUBBYTES[0].a/n952 ,
         \SUBBYTES[0].a/n951 , \SUBBYTES[0].a/n950 , \SUBBYTES[0].a/n949 ,
         \SUBBYTES[0].a/n948 , \SUBBYTES[0].a/n947 , \SUBBYTES[0].a/n946 ,
         \SUBBYTES[0].a/n945 , \SUBBYTES[0].a/n944 , \SUBBYTES[0].a/n943 ,
         \SUBBYTES[0].a/n942 , \SUBBYTES[0].a/n941 , \SUBBYTES[0].a/n940 ,
         \SUBBYTES[0].a/n939 , \SUBBYTES[0].a/n938 , \SUBBYTES[0].a/n937 ,
         \SUBBYTES[0].a/n936 , \SUBBYTES[0].a/n935 , \SUBBYTES[0].a/n934 ,
         \SUBBYTES[0].a/n933 , \SUBBYTES[0].a/n932 , \SUBBYTES[0].a/n931 ,
         \SUBBYTES[0].a/n930 , \SUBBYTES[0].a/n929 , \SUBBYTES[0].a/n928 ,
         \SUBBYTES[0].a/n927 , \SUBBYTES[0].a/n926 , \SUBBYTES[0].a/n925 ,
         \SUBBYTES[0].a/n924 , \SUBBYTES[0].a/n923 , \SUBBYTES[0].a/n922 ,
         \SUBBYTES[0].a/n921 , \SUBBYTES[0].a/n920 , \SUBBYTES[0].a/n919 ,
         \SUBBYTES[0].a/n918 , \SUBBYTES[0].a/n917 , \SUBBYTES[0].a/n916 ,
         \SUBBYTES[0].a/n915 , \SUBBYTES[0].a/n914 , \SUBBYTES[0].a/n913 ,
         \SUBBYTES[0].a/n912 , \SUBBYTES[0].a/n911 , \SUBBYTES[0].a/n910 ,
         \SUBBYTES[0].a/n909 , \SUBBYTES[0].a/n908 , \SUBBYTES[0].a/n907 ,
         \SUBBYTES[0].a/n906 , \SUBBYTES[0].a/n905 , \SUBBYTES[0].a/n904 ,
         \SUBBYTES[0].a/n903 , \SUBBYTES[0].a/n902 , \SUBBYTES[0].a/n901 ,
         \SUBBYTES[0].a/n900 , \SUBBYTES[0].a/n899 , \SUBBYTES[0].a/n898 ,
         \SUBBYTES[0].a/n897 , \SUBBYTES[0].a/n896 , \SUBBYTES[0].a/n895 ,
         \SUBBYTES[0].a/n894 , \SUBBYTES[0].a/n893 , \SUBBYTES[0].a/n892 ,
         \SUBBYTES[0].a/n891 , \SUBBYTES[0].a/n890 , \SUBBYTES[0].a/n889 ,
         \SUBBYTES[0].a/n888 , \SUBBYTES[0].a/n887 , \SUBBYTES[0].a/n886 ,
         \SUBBYTES[0].a/n885 , \SUBBYTES[0].a/n884 , \SUBBYTES[0].a/n883 ,
         \SUBBYTES[0].a/n882 , \SUBBYTES[0].a/n881 , \SUBBYTES[0].a/n880 ,
         \SUBBYTES[0].a/n879 , \SUBBYTES[0].a/n878 , \SUBBYTES[0].a/n877 ,
         \SUBBYTES[0].a/n876 , \SUBBYTES[0].a/n875 , \SUBBYTES[0].a/n874 ,
         \SUBBYTES[0].a/n873 , \SUBBYTES[0].a/n872 , \SUBBYTES[0].a/n871 ,
         \SUBBYTES[0].a/n870 , \SUBBYTES[0].a/n869 , \SUBBYTES[0].a/n868 ,
         \SUBBYTES[0].a/n867 , \SUBBYTES[0].a/n866 , \SUBBYTES[0].a/n865 ,
         \SUBBYTES[0].a/n864 , \SUBBYTES[0].a/n863 , \SUBBYTES[0].a/n862 ,
         \SUBBYTES[0].a/n861 , \SUBBYTES[0].a/n860 , \SUBBYTES[0].a/n859 ,
         \SUBBYTES[0].a/n858 , \SUBBYTES[0].a/n857 , \SUBBYTES[0].a/n856 ,
         \SUBBYTES[0].a/n855 , \SUBBYTES[0].a/n854 , \SUBBYTES[0].a/n853 ,
         \SUBBYTES[0].a/n852 , \SUBBYTES[0].a/n851 , \SUBBYTES[0].a/n850 ,
         \SUBBYTES[0].a/n849 , \SUBBYTES[0].a/n848 , \SUBBYTES[0].a/n847 ,
         \SUBBYTES[0].a/n846 , \SUBBYTES[0].a/n845 , \SUBBYTES[0].a/n844 ,
         \SUBBYTES[0].a/n843 , \SUBBYTES[0].a/n842 , \SUBBYTES[0].a/n841 ,
         \SUBBYTES[0].a/n840 , \SUBBYTES[0].a/n839 , \SUBBYTES[0].a/n838 ,
         \SUBBYTES[0].a/n837 , \SUBBYTES[0].a/n836 , \SUBBYTES[0].a/n835 ,
         \SUBBYTES[0].a/n834 , \SUBBYTES[0].a/n833 , \SUBBYTES[0].a/n832 ,
         \SUBBYTES[0].a/n831 , \SUBBYTES[0].a/n830 , \SUBBYTES[0].a/n829 ,
         \SUBBYTES[0].a/n828 , \SUBBYTES[0].a/n827 , \SUBBYTES[0].a/n826 ,
         \SUBBYTES[0].a/n825 , \SUBBYTES[0].a/n824 , \SUBBYTES[0].a/n823 ,
         \SUBBYTES[0].a/n822 , \SUBBYTES[0].a/n821 , \SUBBYTES[0].a/n820 ,
         \SUBBYTES[0].a/n819 , \SUBBYTES[0].a/n818 , \SUBBYTES[0].a/n817 ,
         \SUBBYTES[0].a/n816 , \SUBBYTES[0].a/n815 , \SUBBYTES[0].a/n814 ,
         \SUBBYTES[0].a/n813 , \SUBBYTES[0].a/n812 , \SUBBYTES[0].a/n811 ,
         \SUBBYTES[0].a/n810 , \SUBBYTES[0].a/n809 , \SUBBYTES[0].a/n808 ,
         \SUBBYTES[0].a/n807 , \SUBBYTES[0].a/n806 , \SUBBYTES[0].a/n805 ,
         \SUBBYTES[0].a/n804 , \SUBBYTES[0].a/n803 , \SUBBYTES[0].a/n802 ,
         \SUBBYTES[0].a/n801 , \SUBBYTES[0].a/n800 , \SUBBYTES[0].a/n799 ,
         \SUBBYTES[0].a/n798 , \SUBBYTES[0].a/n797 , \SUBBYTES[0].a/n796 ,
         \SUBBYTES[0].a/n795 , \SUBBYTES[0].a/n794 , \SUBBYTES[0].a/n793 ,
         \SUBBYTES[0].a/n792 , \SUBBYTES[0].a/n791 , \SUBBYTES[0].a/n790 ,
         \SUBBYTES[0].a/n789 , \SUBBYTES[0].a/n788 , \SUBBYTES[0].a/n787 ,
         \SUBBYTES[0].a/n786 , \SUBBYTES[0].a/n785 , \SUBBYTES[0].a/n784 ,
         \SUBBYTES[0].a/n783 , \SUBBYTES[0].a/n782 , \SUBBYTES[0].a/n781 ,
         \SUBBYTES[0].a/n780 , \SUBBYTES[0].a/n779 , \SUBBYTES[0].a/n778 ,
         \SUBBYTES[0].a/n777 , \SUBBYTES[0].a/n776 , \SUBBYTES[0].a/n775 ,
         \SUBBYTES[0].a/n774 , \SUBBYTES[0].a/n773 , \SUBBYTES[0].a/n772 ,
         \SUBBYTES[0].a/n771 , \SUBBYTES[0].a/n770 , \SUBBYTES[0].a/n769 ,
         \SUBBYTES[0].a/n768 , \SUBBYTES[0].a/n767 , \SUBBYTES[0].a/n766 ,
         \SUBBYTES[0].a/n765 , \SUBBYTES[0].a/n764 , \SUBBYTES[0].a/n763 ,
         \SUBBYTES[0].a/n762 , \SUBBYTES[0].a/n761 , \SUBBYTES[0].a/n760 ,
         \SUBBYTES[0].a/n759 , \SUBBYTES[0].a/n758 , \SUBBYTES[0].a/n757 ,
         \SUBBYTES[0].a/n756 , \SUBBYTES[0].a/n755 , \SUBBYTES[0].a/n754 ,
         \SUBBYTES[0].a/n753 , \SUBBYTES[0].a/n752 , \SUBBYTES[0].a/n751 ,
         \SUBBYTES[0].a/n750 , \SUBBYTES[0].a/n749 , \SUBBYTES[0].a/n748 ,
         \SUBBYTES[0].a/n747 , \SUBBYTES[0].a/n746 , \SUBBYTES[0].a/n745 ,
         \SUBBYTES[0].a/n744 , \SUBBYTES[0].a/n743 , \SUBBYTES[0].a/n742 ,
         \SUBBYTES[0].a/n741 , \SUBBYTES[0].a/n740 , \SUBBYTES[0].a/n739 ,
         \SUBBYTES[0].a/n738 , \SUBBYTES[0].a/n737 , \SUBBYTES[0].a/n736 ,
         \SUBBYTES[0].a/n735 , \SUBBYTES[0].a/n734 , \SUBBYTES[0].a/n733 ,
         \SUBBYTES[0].a/n732 , \SUBBYTES[0].a/n731 , \SUBBYTES[0].a/n730 ,
         \SUBBYTES[0].a/n729 , \SUBBYTES[0].a/n728 , \SUBBYTES[0].a/n727 ,
         \SUBBYTES[0].a/n726 , \SUBBYTES[0].a/n725 , \SUBBYTES[0].a/n724 ,
         \SUBBYTES[0].a/n723 , \SUBBYTES[0].a/n722 , \SUBBYTES[0].a/n721 ,
         \SUBBYTES[0].a/n720 , \SUBBYTES[0].a/n719 , \SUBBYTES[0].a/n718 ,
         \SUBBYTES[0].a/n717 , \SUBBYTES[0].a/n716 , \SUBBYTES[0].a/n715 ,
         \SUBBYTES[0].a/n714 , \SUBBYTES[0].a/n713 , \SUBBYTES[0].a/n712 ,
         \SUBBYTES[0].a/n711 , \SUBBYTES[0].a/n710 , \SUBBYTES[0].a/n709 ,
         \SUBBYTES[0].a/n708 , \SUBBYTES[0].a/n707 , \SUBBYTES[0].a/n706 ,
         \SUBBYTES[0].a/n705 , \SUBBYTES[0].a/n704 , \SUBBYTES[0].a/n703 ,
         \SUBBYTES[0].a/n702 , \SUBBYTES[0].a/n701 , \SUBBYTES[0].a/n700 ,
         \SUBBYTES[0].a/n699 , \SUBBYTES[0].a/n698 , \SUBBYTES[0].a/n697 ,
         \SUBBYTES[0].a/n696 , \SUBBYTES[0].a/n695 , \SUBBYTES[0].a/n694 ,
         \SUBBYTES[0].a/n693 , \SUBBYTES[0].a/n692 , \SUBBYTES[0].a/n691 ,
         \SUBBYTES[0].a/n690 , \SUBBYTES[0].a/n689 , \SUBBYTES[0].a/n688 ,
         \SUBBYTES[0].a/n687 , \SUBBYTES[0].a/n686 , \SUBBYTES[0].a/n685 ,
         \SUBBYTES[0].a/n684 , \SUBBYTES[0].a/n683 , \SUBBYTES[0].a/n682 ,
         \SUBBYTES[0].a/n681 , \SUBBYTES[0].a/n680 , \SUBBYTES[0].a/n679 ,
         \SUBBYTES[0].a/n678 , \SUBBYTES[0].a/n677 , \SUBBYTES[0].a/n676 ,
         \SUBBYTES[0].a/n675 , \SUBBYTES[0].a/n674 , \SUBBYTES[0].a/n673 ,
         \SUBBYTES[0].a/n672 , \SUBBYTES[0].a/n671 , \SUBBYTES[0].a/n670 ,
         \SUBBYTES[0].a/n669 , \SUBBYTES[0].a/n668 , \SUBBYTES[0].a/n667 ,
         \SUBBYTES[0].a/n666 , \SUBBYTES[0].a/n665 , \SUBBYTES[0].a/n664 ,
         \SUBBYTES[0].a/n663 , \SUBBYTES[0].a/n662 , \SUBBYTES[0].a/n661 ,
         \SUBBYTES[0].a/n660 , \SUBBYTES[0].a/n659 , \SUBBYTES[0].a/n658 ,
         \SUBBYTES[0].a/n657 , \SUBBYTES[0].a/n656 , \SUBBYTES[0].a/n655 ,
         \SUBBYTES[0].a/n654 , \SUBBYTES[0].a/n653 , \SUBBYTES[0].a/n652 ,
         \SUBBYTES[0].a/n651 , \SUBBYTES[0].a/n650 , \SUBBYTES[0].a/n649 ,
         \SUBBYTES[0].a/n648 , \SUBBYTES[0].a/n647 , \SUBBYTES[0].a/n646 ,
         \SUBBYTES[0].a/n645 , \SUBBYTES[0].a/n644 , \SUBBYTES[0].a/n643 ,
         \SUBBYTES[0].a/n642 , \SUBBYTES[0].a/n641 , \SUBBYTES[0].a/n640 ,
         \SUBBYTES[0].a/n639 , \SUBBYTES[0].a/n638 , \SUBBYTES[0].a/n637 ,
         \SUBBYTES[0].a/n636 , \SUBBYTES[0].a/n635 , \SUBBYTES[0].a/n634 ,
         \SUBBYTES[0].a/n633 , \SUBBYTES[0].a/n632 , \SUBBYTES[0].a/n631 ,
         \SUBBYTES[0].a/n630 , \SUBBYTES[0].a/n629 , \SUBBYTES[0].a/n628 ,
         \SUBBYTES[0].a/n627 , \SUBBYTES[0].a/n626 , \SUBBYTES[0].a/n625 ,
         \SUBBYTES[0].a/n624 , \SUBBYTES[0].a/n623 , \SUBBYTES[0].a/n622 ,
         \SUBBYTES[0].a/n621 , \SUBBYTES[0].a/n620 , \SUBBYTES[0].a/n619 ,
         \SUBBYTES[0].a/n618 , \SUBBYTES[0].a/n617 , \SUBBYTES[0].a/n616 ,
         \SUBBYTES[0].a/n615 , \SUBBYTES[0].a/n614 , \SUBBYTES[0].a/n613 ,
         \SUBBYTES[0].a/n612 , \SUBBYTES[0].a/n611 , \SUBBYTES[0].a/n610 ,
         \SUBBYTES[0].a/n609 , \SUBBYTES[0].a/n608 , \SUBBYTES[0].a/n607 ,
         \SUBBYTES[0].a/n606 , \SUBBYTES[0].a/n605 , \SUBBYTES[0].a/n604 ,
         \SUBBYTES[0].a/n603 , \SUBBYTES[0].a/n602 , \SUBBYTES[0].a/n601 ,
         \SUBBYTES[0].a/n600 , \SUBBYTES[0].a/n599 , \SUBBYTES[0].a/n598 ,
         \SUBBYTES[0].a/n597 , \SUBBYTES[0].a/n596 , \SUBBYTES[0].a/n595 ,
         \SUBBYTES[0].a/n594 , \SUBBYTES[0].a/n593 , \SUBBYTES[0].a/n592 ,
         \SUBBYTES[0].a/n591 , \SUBBYTES[0].a/n590 , \SUBBYTES[0].a/n589 ,
         \SUBBYTES[0].a/n588 , \SUBBYTES[0].a/n587 , \SUBBYTES[0].a/n586 ,
         \SUBBYTES[0].a/n585 , \SUBBYTES[0].a/n584 , \SUBBYTES[0].a/n583 ,
         \SUBBYTES[0].a/n582 , \SUBBYTES[0].a/n581 , \SUBBYTES[0].a/n580 ,
         \SUBBYTES[0].a/n579 , \SUBBYTES[0].a/n578 , \SUBBYTES[0].a/n577 ,
         \SUBBYTES[0].a/n576 , \SUBBYTES[0].a/n575 , \SUBBYTES[0].a/n574 ,
         \SUBBYTES[0].a/n573 , \SUBBYTES[0].a/n572 , \SUBBYTES[0].a/n571 ,
         \SUBBYTES[0].a/n570 , \SUBBYTES[0].a/n569 , \SUBBYTES[0].a/n568 ,
         \SUBBYTES[0].a/n567 , \SUBBYTES[0].a/n566 , \SUBBYTES[0].a/n565 ,
         \SUBBYTES[0].a/n564 , \SUBBYTES[0].a/n563 , \SUBBYTES[0].a/n562 ,
         \SUBBYTES[0].a/n561 , \SUBBYTES[0].a/n560 , \SUBBYTES[0].a/n559 ,
         \SUBBYTES[0].a/n558 , \SUBBYTES[0].a/n557 , \SUBBYTES[0].a/n556 ,
         \SUBBYTES[0].a/n555 , \SUBBYTES[0].a/n554 , \SUBBYTES[0].a/n553 ,
         \SUBBYTES[0].a/n552 , \SUBBYTES[0].a/n551 , \SUBBYTES[0].a/n550 ,
         \SUBBYTES[0].a/n549 , \SUBBYTES[0].a/n548 , \SUBBYTES[0].a/n547 ,
         \SUBBYTES[0].a/n546 , \SUBBYTES[0].a/n545 , \SUBBYTES[0].a/n544 ,
         \SUBBYTES[0].a/n543 , \SUBBYTES[0].a/n542 , \SUBBYTES[0].a/n541 ,
         \SUBBYTES[0].a/n540 , \SUBBYTES[0].a/n539 , \SUBBYTES[0].a/n538 ,
         \SUBBYTES[0].a/n537 , \SUBBYTES[0].a/n536 , \SUBBYTES[0].a/n535 ,
         \SUBBYTES[0].a/n534 , \SUBBYTES[0].a/n533 , \SUBBYTES[0].a/n532 ,
         \SUBBYTES[0].a/n531 , \SUBBYTES[0].a/n530 , \SUBBYTES[0].a/n529 ,
         \SUBBYTES[0].a/n528 , \SUBBYTES[0].a/n527 , \SUBBYTES[0].a/n526 ,
         \SUBBYTES[0].a/n525 , \SUBBYTES[0].a/n524 , \SUBBYTES[0].a/n523 ,
         \SUBBYTES[0].a/n522 , \SUBBYTES[0].a/n521 , \SUBBYTES[0].a/n520 ,
         \SUBBYTES[0].a/n519 , \SUBBYTES[0].a/n518 , \SUBBYTES[0].a/n517 ,
         \SUBBYTES[0].a/n516 , \SUBBYTES[0].a/n515 , \SUBBYTES[0].a/n514 ,
         \SUBBYTES[0].a/n513 , \SUBBYTES[0].a/n512 , \SUBBYTES[0].a/n511 ,
         \SUBBYTES[0].a/n510 , \SUBBYTES[0].a/n509 , \SUBBYTES[0].a/n508 ,
         \SUBBYTES[0].a/n507 , \SUBBYTES[0].a/n506 , \SUBBYTES[0].a/n505 ,
         \SUBBYTES[0].a/n504 , \SUBBYTES[0].a/n503 , \SUBBYTES[0].a/n502 ,
         \SUBBYTES[0].a/n501 , \SUBBYTES[0].a/n500 , \SUBBYTES[0].a/n499 ,
         \SUBBYTES[0].a/n498 , \SUBBYTES[0].a/n497 , \SUBBYTES[0].a/n496 ,
         \SUBBYTES[0].a/n495 , \SUBBYTES[0].a/n494 , \SUBBYTES[0].a/n493 ,
         \SUBBYTES[0].a/n492 , \SUBBYTES[0].a/n491 , \SUBBYTES[0].a/n490 ,
         \SUBBYTES[0].a/n489 , \SUBBYTES[0].a/n488 , \SUBBYTES[0].a/n487 ,
         \SUBBYTES[0].a/n486 , \SUBBYTES[0].a/n485 , \SUBBYTES[0].a/n484 ,
         \SUBBYTES[0].a/n483 , \SUBBYTES[0].a/n482 , \SUBBYTES[0].a/n481 ,
         \SUBBYTES[0].a/n480 , \SUBBYTES[0].a/n479 , \SUBBYTES[0].a/n478 ,
         \SUBBYTES[0].a/n477 , \SUBBYTES[0].a/n476 , \SUBBYTES[0].a/n475 ,
         \SUBBYTES[0].a/n474 , \SUBBYTES[0].a/n473 , \SUBBYTES[0].a/n472 ,
         \SUBBYTES[0].a/n471 , \SUBBYTES[0].a/n470 , \SUBBYTES[0].a/n469 ,
         \SUBBYTES[0].a/n468 , \SUBBYTES[0].a/n467 , \SUBBYTES[0].a/n466 ,
         \SUBBYTES[0].a/n465 , \SUBBYTES[0].a/n464 , \SUBBYTES[0].a/n463 ,
         \SUBBYTES[0].a/n462 , \SUBBYTES[0].a/n461 , \SUBBYTES[0].a/n460 ,
         \SUBBYTES[0].a/n459 , \SUBBYTES[0].a/n458 , \SUBBYTES[0].a/n457 ,
         \SUBBYTES[0].a/n456 , \SUBBYTES[0].a/n455 , \SUBBYTES[0].a/n454 ,
         \SUBBYTES[0].a/n453 , \SUBBYTES[0].a/n452 , \SUBBYTES[0].a/n451 ,
         \SUBBYTES[0].a/n450 , \SUBBYTES[0].a/n449 , \SUBBYTES[0].a/n448 ,
         \SUBBYTES[0].a/n447 , \SUBBYTES[0].a/n446 , \SUBBYTES[0].a/n445 ,
         \SUBBYTES[0].a/n444 , \SUBBYTES[0].a/n443 , \SUBBYTES[0].a/n442 ,
         \SUBBYTES[0].a/n441 , \SUBBYTES[0].a/n440 , \SUBBYTES[0].a/n439 ,
         \SUBBYTES[0].a/n438 , \SUBBYTES[0].a/n437 , \SUBBYTES[0].a/n436 ,
         \SUBBYTES[0].a/n435 , \SUBBYTES[0].a/n434 , \SUBBYTES[0].a/n433 ,
         \SUBBYTES[0].a/n432 , \SUBBYTES[0].a/n431 , \SUBBYTES[0].a/n430 ,
         \SUBBYTES[0].a/n429 , \SUBBYTES[0].a/n428 , \SUBBYTES[0].a/n427 ,
         \SUBBYTES[0].a/n426 , \SUBBYTES[0].a/n425 , \SUBBYTES[0].a/n424 ,
         \SUBBYTES[0].a/n423 , \SUBBYTES[0].a/n422 , \SUBBYTES[0].a/n421 ,
         \SUBBYTES[0].a/n420 , \SUBBYTES[0].a/n419 , \SUBBYTES[0].a/n418 ,
         \SUBBYTES[0].a/n417 , \SUBBYTES[0].a/n416 , \SUBBYTES[0].a/n415 ,
         \SUBBYTES[0].a/n414 , \SUBBYTES[0].a/n413 , \SUBBYTES[0].a/n412 ,
         \SUBBYTES[0].a/n411 , \SUBBYTES[0].a/n410 , \SUBBYTES[0].a/n409 ,
         \SUBBYTES[0].a/n408 , \SUBBYTES[0].a/n407 , \SUBBYTES[0].a/n406 ,
         \SUBBYTES[0].a/n405 , \SUBBYTES[0].a/n404 , \SUBBYTES[0].a/n403 ,
         \SUBBYTES[0].a/n402 , \SUBBYTES[0].a/n401 , \SUBBYTES[0].a/n400 ,
         \SUBBYTES[0].a/n399 , \SUBBYTES[0].a/n398 , \SUBBYTES[0].a/n397 ,
         \SUBBYTES[0].a/n396 , \SUBBYTES[0].a/n395 , \SUBBYTES[0].a/n394 ,
         \SUBBYTES[0].a/n393 , \SUBBYTES[0].a/n392 , \SUBBYTES[0].a/n391 ,
         \SUBBYTES[0].a/n390 , \SUBBYTES[0].a/n389 , \SUBBYTES[0].a/n388 ,
         \SUBBYTES[0].a/n387 , \SUBBYTES[0].a/n386 , \SUBBYTES[0].a/n385 ,
         \SUBBYTES[0].a/n160 , \SUBBYTES[0].a/n159 , \SUBBYTES[0].a/n150 ,
         \SUBBYTES[0].a/n149 , \SUBBYTES[0].a/n140 , \SUBBYTES[0].a/n139 ,
         \SUBBYTES[0].a/n130 , \SUBBYTES[0].a/n129 , \SUBBYTES[0].a/n120 ,
         \SUBBYTES[0].a/n119 , \SUBBYTES[0].a/n110 , \SUBBYTES[0].a/n109 ,
         \SUBBYTES[0].a/n100 , \SUBBYTES[0].a/n99 , \SUBBYTES[0].a/n90 ,
         \SUBBYTES[0].a/n89 , \SUBBYTES[0].a/n80 , \SUBBYTES[0].a/n79 ,
         \SUBBYTES[0].a/n70 , \SUBBYTES[0].a/n69 , \SUBBYTES[0].a/n60 ,
         \SUBBYTES[0].a/n59 , \SUBBYTES[0].a/n50 , \SUBBYTES[0].a/n49 ,
         \SUBBYTES[0].a/n40 , \SUBBYTES[0].a/n39 , \SUBBYTES[0].a/n30 ,
         \SUBBYTES[0].a/n29 , \SUBBYTES[0].a/n20 , \SUBBYTES[0].a/n19 ,
         \SUBBYTES[0].a/n10 , \SUBBYTES[0].a/n9 , \SUBBYTES[0].a/w3400 ,
         \SUBBYTES[0].a/w3398 , \SUBBYTES[0].a/w3397 , \SUBBYTES[0].a/w3396 ,
         \SUBBYTES[0].a/w3393 , \SUBBYTES[0].a/w3391 , \SUBBYTES[0].a/w3390 ,
         \SUBBYTES[0].a/w3389 , \SUBBYTES[0].a/w3385 , \SUBBYTES[0].a/w3383 ,
         \SUBBYTES[0].a/w3382 , \SUBBYTES[0].a/w3381 , \SUBBYTES[0].a/w3380 ,
         \SUBBYTES[0].a/w3379 , \SUBBYTES[0].a/w3378 , \SUBBYTES[0].a/w3377 ,
         \SUBBYTES[0].a/w3376 , \SUBBYTES[0].a/w3368 , \SUBBYTES[0].a/w3366 ,
         \SUBBYTES[0].a/w3365 , \SUBBYTES[0].a/w3361 , \SUBBYTES[0].a/w3359 ,
         \SUBBYTES[0].a/w3358 , \SUBBYTES[0].a/w3357 , \SUBBYTES[0].a/w3353 ,
         \SUBBYTES[0].a/w3351 , \SUBBYTES[0].a/w3350 , \SUBBYTES[0].a/w3337 ,
         \SUBBYTES[0].a/w3336 , \SUBBYTES[0].a/w3335 , \SUBBYTES[0].a/w3333 ,
         \SUBBYTES[0].a/w3330 , \SUBBYTES[0].a/w3329 , \SUBBYTES[0].a/w3327 ,
         \SUBBYTES[0].a/w3326 , \SUBBYTES[0].a/w3324 , \SUBBYTES[0].a/w3322 ,
         \SUBBYTES[0].a/w3321 , \SUBBYTES[0].a/w3315 , \SUBBYTES[0].a/w3314 ,
         \SUBBYTES[0].a/w3313 , \SUBBYTES[0].a/w3312 , \SUBBYTES[0].a/w3306 ,
         \SUBBYTES[0].a/w3304 , \SUBBYTES[0].a/w3303 , \SUBBYTES[0].a/w3299 ,
         \SUBBYTES[0].a/w3297 , \SUBBYTES[0].a/w3296 , \SUBBYTES[0].a/w3291 ,
         \SUBBYTES[0].a/w3289 , \SUBBYTES[0].a/w3288 , \SUBBYTES[0].a/w3272 ,
         \SUBBYTES[0].a/w3271 , \SUBBYTES[0].a/w3270 , \SUBBYTES[0].a/w3269 ,
         \SUBBYTES[0].a/w3268 , \SUBBYTES[0].a/w3266 , \SUBBYTES[0].a/w3265 ,
         \SUBBYTES[0].a/w3193 , \SUBBYTES[0].a/w3191 , \SUBBYTES[0].a/w3190 ,
         \SUBBYTES[0].a/w3189 , \SUBBYTES[0].a/w3186 , \SUBBYTES[0].a/w3184 ,
         \SUBBYTES[0].a/w3183 , \SUBBYTES[0].a/w3182 , \SUBBYTES[0].a/w3178 ,
         \SUBBYTES[0].a/w3176 , \SUBBYTES[0].a/w3175 , \SUBBYTES[0].a/w3174 ,
         \SUBBYTES[0].a/w3173 , \SUBBYTES[0].a/w3172 , \SUBBYTES[0].a/w3171 ,
         \SUBBYTES[0].a/w3170 , \SUBBYTES[0].a/w3169 , \SUBBYTES[0].a/w3161 ,
         \SUBBYTES[0].a/w3159 , \SUBBYTES[0].a/w3158 , \SUBBYTES[0].a/w3154 ,
         \SUBBYTES[0].a/w3152 , \SUBBYTES[0].a/w3151 , \SUBBYTES[0].a/w3150 ,
         \SUBBYTES[0].a/w3146 , \SUBBYTES[0].a/w3144 , \SUBBYTES[0].a/w3143 ,
         \SUBBYTES[0].a/w3130 , \SUBBYTES[0].a/w3129 , \SUBBYTES[0].a/w3128 ,
         \SUBBYTES[0].a/w3126 , \SUBBYTES[0].a/w3123 , \SUBBYTES[0].a/w3122 ,
         \SUBBYTES[0].a/w3120 , \SUBBYTES[0].a/w3119 , \SUBBYTES[0].a/w3117 ,
         \SUBBYTES[0].a/w3115 , \SUBBYTES[0].a/w3114 , \SUBBYTES[0].a/w3108 ,
         \SUBBYTES[0].a/w3107 , \SUBBYTES[0].a/w3106 , \SUBBYTES[0].a/w3105 ,
         \SUBBYTES[0].a/w3099 , \SUBBYTES[0].a/w3097 , \SUBBYTES[0].a/w3096 ,
         \SUBBYTES[0].a/w3092 , \SUBBYTES[0].a/w3090 , \SUBBYTES[0].a/w3089 ,
         \SUBBYTES[0].a/w3084 , \SUBBYTES[0].a/w3082 , \SUBBYTES[0].a/w3081 ,
         \SUBBYTES[0].a/w3065 , \SUBBYTES[0].a/w3064 , \SUBBYTES[0].a/w3063 ,
         \SUBBYTES[0].a/w3062 , \SUBBYTES[0].a/w3061 , \SUBBYTES[0].a/w3059 ,
         \SUBBYTES[0].a/w3058 , \SUBBYTES[0].a/w2986 , \SUBBYTES[0].a/w2984 ,
         \SUBBYTES[0].a/w2983 , \SUBBYTES[0].a/w2982 , \SUBBYTES[0].a/w2979 ,
         \SUBBYTES[0].a/w2977 , \SUBBYTES[0].a/w2976 , \SUBBYTES[0].a/w2975 ,
         \SUBBYTES[0].a/w2971 , \SUBBYTES[0].a/w2969 , \SUBBYTES[0].a/w2968 ,
         \SUBBYTES[0].a/w2967 , \SUBBYTES[0].a/w2966 , \SUBBYTES[0].a/w2965 ,
         \SUBBYTES[0].a/w2964 , \SUBBYTES[0].a/w2963 , \SUBBYTES[0].a/w2962 ,
         \SUBBYTES[0].a/w2954 , \SUBBYTES[0].a/w2952 , \SUBBYTES[0].a/w2951 ,
         \SUBBYTES[0].a/w2947 , \SUBBYTES[0].a/w2945 , \SUBBYTES[0].a/w2944 ,
         \SUBBYTES[0].a/w2943 , \SUBBYTES[0].a/w2939 , \SUBBYTES[0].a/w2937 ,
         \SUBBYTES[0].a/w2936 , \SUBBYTES[0].a/w2923 , \SUBBYTES[0].a/w2922 ,
         \SUBBYTES[0].a/w2921 , \SUBBYTES[0].a/w2919 , \SUBBYTES[0].a/w2916 ,
         \SUBBYTES[0].a/w2915 , \SUBBYTES[0].a/w2913 , \SUBBYTES[0].a/w2912 ,
         \SUBBYTES[0].a/w2910 , \SUBBYTES[0].a/w2908 , \SUBBYTES[0].a/w2907 ,
         \SUBBYTES[0].a/w2901 , \SUBBYTES[0].a/w2900 , \SUBBYTES[0].a/w2899 ,
         \SUBBYTES[0].a/w2898 , \SUBBYTES[0].a/w2892 , \SUBBYTES[0].a/w2890 ,
         \SUBBYTES[0].a/w2889 , \SUBBYTES[0].a/w2885 , \SUBBYTES[0].a/w2883 ,
         \SUBBYTES[0].a/w2882 , \SUBBYTES[0].a/w2877 , \SUBBYTES[0].a/w2875 ,
         \SUBBYTES[0].a/w2874 , \SUBBYTES[0].a/w2858 , \SUBBYTES[0].a/w2857 ,
         \SUBBYTES[0].a/w2856 , \SUBBYTES[0].a/w2855 , \SUBBYTES[0].a/w2854 ,
         \SUBBYTES[0].a/w2852 , \SUBBYTES[0].a/w2851 , \SUBBYTES[0].a/w2779 ,
         \SUBBYTES[0].a/w2777 , \SUBBYTES[0].a/w2776 , \SUBBYTES[0].a/w2775 ,
         \SUBBYTES[0].a/w2772 , \SUBBYTES[0].a/w2770 , \SUBBYTES[0].a/w2769 ,
         \SUBBYTES[0].a/w2768 , \SUBBYTES[0].a/w2764 , \SUBBYTES[0].a/w2762 ,
         \SUBBYTES[0].a/w2761 , \SUBBYTES[0].a/w2760 , \SUBBYTES[0].a/w2759 ,
         \SUBBYTES[0].a/w2758 , \SUBBYTES[0].a/w2757 , \SUBBYTES[0].a/w2756 ,
         \SUBBYTES[0].a/w2755 , \SUBBYTES[0].a/w2747 , \SUBBYTES[0].a/w2745 ,
         \SUBBYTES[0].a/w2744 , \SUBBYTES[0].a/w2740 , \SUBBYTES[0].a/w2738 ,
         \SUBBYTES[0].a/w2737 , \SUBBYTES[0].a/w2736 , \SUBBYTES[0].a/w2732 ,
         \SUBBYTES[0].a/w2730 , \SUBBYTES[0].a/w2729 , \SUBBYTES[0].a/w2716 ,
         \SUBBYTES[0].a/w2715 , \SUBBYTES[0].a/w2714 , \SUBBYTES[0].a/w2712 ,
         \SUBBYTES[0].a/w2709 , \SUBBYTES[0].a/w2708 , \SUBBYTES[0].a/w2706 ,
         \SUBBYTES[0].a/w2705 , \SUBBYTES[0].a/w2703 , \SUBBYTES[0].a/w2701 ,
         \SUBBYTES[0].a/w2700 , \SUBBYTES[0].a/w2694 , \SUBBYTES[0].a/w2693 ,
         \SUBBYTES[0].a/w2692 , \SUBBYTES[0].a/w2691 , \SUBBYTES[0].a/w2685 ,
         \SUBBYTES[0].a/w2683 , \SUBBYTES[0].a/w2682 , \SUBBYTES[0].a/w2678 ,
         \SUBBYTES[0].a/w2676 , \SUBBYTES[0].a/w2675 , \SUBBYTES[0].a/w2670 ,
         \SUBBYTES[0].a/w2668 , \SUBBYTES[0].a/w2667 , \SUBBYTES[0].a/w2651 ,
         \SUBBYTES[0].a/w2650 , \SUBBYTES[0].a/w2649 , \SUBBYTES[0].a/w2648 ,
         \SUBBYTES[0].a/w2647 , \SUBBYTES[0].a/w2645 , \SUBBYTES[0].a/w2644 ,
         \SUBBYTES[0].a/w2572 , \SUBBYTES[0].a/w2570 , \SUBBYTES[0].a/w2569 ,
         \SUBBYTES[0].a/w2568 , \SUBBYTES[0].a/w2565 , \SUBBYTES[0].a/w2563 ,
         \SUBBYTES[0].a/w2562 , \SUBBYTES[0].a/w2561 , \SUBBYTES[0].a/w2557 ,
         \SUBBYTES[0].a/w2555 , \SUBBYTES[0].a/w2554 , \SUBBYTES[0].a/w2553 ,
         \SUBBYTES[0].a/w2552 , \SUBBYTES[0].a/w2551 , \SUBBYTES[0].a/w2550 ,
         \SUBBYTES[0].a/w2549 , \SUBBYTES[0].a/w2548 , \SUBBYTES[0].a/w2540 ,
         \SUBBYTES[0].a/w2538 , \SUBBYTES[0].a/w2537 , \SUBBYTES[0].a/w2533 ,
         \SUBBYTES[0].a/w2531 , \SUBBYTES[0].a/w2530 , \SUBBYTES[0].a/w2529 ,
         \SUBBYTES[0].a/w2525 , \SUBBYTES[0].a/w2523 , \SUBBYTES[0].a/w2522 ,
         \SUBBYTES[0].a/w2509 , \SUBBYTES[0].a/w2508 , \SUBBYTES[0].a/w2507 ,
         \SUBBYTES[0].a/w2505 , \SUBBYTES[0].a/w2502 , \SUBBYTES[0].a/w2501 ,
         \SUBBYTES[0].a/w2499 , \SUBBYTES[0].a/w2498 , \SUBBYTES[0].a/w2496 ,
         \SUBBYTES[0].a/w2494 , \SUBBYTES[0].a/w2493 , \SUBBYTES[0].a/w2487 ,
         \SUBBYTES[0].a/w2486 , \SUBBYTES[0].a/w2485 , \SUBBYTES[0].a/w2484 ,
         \SUBBYTES[0].a/w2478 , \SUBBYTES[0].a/w2476 , \SUBBYTES[0].a/w2475 ,
         \SUBBYTES[0].a/w2471 , \SUBBYTES[0].a/w2469 , \SUBBYTES[0].a/w2468 ,
         \SUBBYTES[0].a/w2463 , \SUBBYTES[0].a/w2461 , \SUBBYTES[0].a/w2460 ,
         \SUBBYTES[0].a/w2444 , \SUBBYTES[0].a/w2443 , \SUBBYTES[0].a/w2442 ,
         \SUBBYTES[0].a/w2441 , \SUBBYTES[0].a/w2440 , \SUBBYTES[0].a/w2438 ,
         \SUBBYTES[0].a/w2437 , \SUBBYTES[0].a/w2365 , \SUBBYTES[0].a/w2363 ,
         \SUBBYTES[0].a/w2362 , \SUBBYTES[0].a/w2361 , \SUBBYTES[0].a/w2358 ,
         \SUBBYTES[0].a/w2356 , \SUBBYTES[0].a/w2355 , \SUBBYTES[0].a/w2354 ,
         \SUBBYTES[0].a/w2350 , \SUBBYTES[0].a/w2348 , \SUBBYTES[0].a/w2347 ,
         \SUBBYTES[0].a/w2346 , \SUBBYTES[0].a/w2345 , \SUBBYTES[0].a/w2344 ,
         \SUBBYTES[0].a/w2343 , \SUBBYTES[0].a/w2342 , \SUBBYTES[0].a/w2341 ,
         \SUBBYTES[0].a/w2333 , \SUBBYTES[0].a/w2331 , \SUBBYTES[0].a/w2330 ,
         \SUBBYTES[0].a/w2326 , \SUBBYTES[0].a/w2324 , \SUBBYTES[0].a/w2323 ,
         \SUBBYTES[0].a/w2322 , \SUBBYTES[0].a/w2318 , \SUBBYTES[0].a/w2316 ,
         \SUBBYTES[0].a/w2315 , \SUBBYTES[0].a/w2302 , \SUBBYTES[0].a/w2301 ,
         \SUBBYTES[0].a/w2300 , \SUBBYTES[0].a/w2298 , \SUBBYTES[0].a/w2295 ,
         \SUBBYTES[0].a/w2294 , \SUBBYTES[0].a/w2292 , \SUBBYTES[0].a/w2291 ,
         \SUBBYTES[0].a/w2289 , \SUBBYTES[0].a/w2287 , \SUBBYTES[0].a/w2286 ,
         \SUBBYTES[0].a/w2280 , \SUBBYTES[0].a/w2279 , \SUBBYTES[0].a/w2278 ,
         \SUBBYTES[0].a/w2277 , \SUBBYTES[0].a/w2271 , \SUBBYTES[0].a/w2269 ,
         \SUBBYTES[0].a/w2268 , \SUBBYTES[0].a/w2264 , \SUBBYTES[0].a/w2262 ,
         \SUBBYTES[0].a/w2261 , \SUBBYTES[0].a/w2256 , \SUBBYTES[0].a/w2254 ,
         \SUBBYTES[0].a/w2253 , \SUBBYTES[0].a/w2237 , \SUBBYTES[0].a/w2236 ,
         \SUBBYTES[0].a/w2235 , \SUBBYTES[0].a/w2234 , \SUBBYTES[0].a/w2233 ,
         \SUBBYTES[0].a/w2231 , \SUBBYTES[0].a/w2230 , \SUBBYTES[0].a/w2158 ,
         \SUBBYTES[0].a/w2156 , \SUBBYTES[0].a/w2155 , \SUBBYTES[0].a/w2154 ,
         \SUBBYTES[0].a/w2151 , \SUBBYTES[0].a/w2149 , \SUBBYTES[0].a/w2148 ,
         \SUBBYTES[0].a/w2147 , \SUBBYTES[0].a/w2143 , \SUBBYTES[0].a/w2141 ,
         \SUBBYTES[0].a/w2140 , \SUBBYTES[0].a/w2139 , \SUBBYTES[0].a/w2138 ,
         \SUBBYTES[0].a/w2137 , \SUBBYTES[0].a/w2136 , \SUBBYTES[0].a/w2135 ,
         \SUBBYTES[0].a/w2134 , \SUBBYTES[0].a/w2126 , \SUBBYTES[0].a/w2124 ,
         \SUBBYTES[0].a/w2123 , \SUBBYTES[0].a/w2119 , \SUBBYTES[0].a/w2117 ,
         \SUBBYTES[0].a/w2116 , \SUBBYTES[0].a/w2115 , \SUBBYTES[0].a/w2111 ,
         \SUBBYTES[0].a/w2109 , \SUBBYTES[0].a/w2108 , \SUBBYTES[0].a/w2095 ,
         \SUBBYTES[0].a/w2094 , \SUBBYTES[0].a/w2093 , \SUBBYTES[0].a/w2091 ,
         \SUBBYTES[0].a/w2088 , \SUBBYTES[0].a/w2087 , \SUBBYTES[0].a/w2085 ,
         \SUBBYTES[0].a/w2084 , \SUBBYTES[0].a/w2082 , \SUBBYTES[0].a/w2080 ,
         \SUBBYTES[0].a/w2079 , \SUBBYTES[0].a/w2073 , \SUBBYTES[0].a/w2072 ,
         \SUBBYTES[0].a/w2071 , \SUBBYTES[0].a/w2070 , \SUBBYTES[0].a/w2064 ,
         \SUBBYTES[0].a/w2062 , \SUBBYTES[0].a/w2061 , \SUBBYTES[0].a/w2057 ,
         \SUBBYTES[0].a/w2055 , \SUBBYTES[0].a/w2054 , \SUBBYTES[0].a/w2049 ,
         \SUBBYTES[0].a/w2047 , \SUBBYTES[0].a/w2046 , \SUBBYTES[0].a/w2030 ,
         \SUBBYTES[0].a/w2029 , \SUBBYTES[0].a/w2028 , \SUBBYTES[0].a/w2027 ,
         \SUBBYTES[0].a/w2026 , \SUBBYTES[0].a/w2024 , \SUBBYTES[0].a/w2023 ,
         \SUBBYTES[0].a/w1951 , \SUBBYTES[0].a/w1949 , \SUBBYTES[0].a/w1948 ,
         \SUBBYTES[0].a/w1947 , \SUBBYTES[0].a/w1944 , \SUBBYTES[0].a/w1942 ,
         \SUBBYTES[0].a/w1941 , \SUBBYTES[0].a/w1940 , \SUBBYTES[0].a/w1936 ,
         \SUBBYTES[0].a/w1934 , \SUBBYTES[0].a/w1933 , \SUBBYTES[0].a/w1932 ,
         \SUBBYTES[0].a/w1931 , \SUBBYTES[0].a/w1930 , \SUBBYTES[0].a/w1929 ,
         \SUBBYTES[0].a/w1928 , \SUBBYTES[0].a/w1927 , \SUBBYTES[0].a/w1919 ,
         \SUBBYTES[0].a/w1917 , \SUBBYTES[0].a/w1916 , \SUBBYTES[0].a/w1912 ,
         \SUBBYTES[0].a/w1910 , \SUBBYTES[0].a/w1909 , \SUBBYTES[0].a/w1908 ,
         \SUBBYTES[0].a/w1904 , \SUBBYTES[0].a/w1902 , \SUBBYTES[0].a/w1901 ,
         \SUBBYTES[0].a/w1888 , \SUBBYTES[0].a/w1887 , \SUBBYTES[0].a/w1886 ,
         \SUBBYTES[0].a/w1884 , \SUBBYTES[0].a/w1881 , \SUBBYTES[0].a/w1880 ,
         \SUBBYTES[0].a/w1878 , \SUBBYTES[0].a/w1877 , \SUBBYTES[0].a/w1875 ,
         \SUBBYTES[0].a/w1873 , \SUBBYTES[0].a/w1872 , \SUBBYTES[0].a/w1866 ,
         \SUBBYTES[0].a/w1865 , \SUBBYTES[0].a/w1864 , \SUBBYTES[0].a/w1863 ,
         \SUBBYTES[0].a/w1857 , \SUBBYTES[0].a/w1855 , \SUBBYTES[0].a/w1854 ,
         \SUBBYTES[0].a/w1850 , \SUBBYTES[0].a/w1848 , \SUBBYTES[0].a/w1847 ,
         \SUBBYTES[0].a/w1842 , \SUBBYTES[0].a/w1840 , \SUBBYTES[0].a/w1839 ,
         \SUBBYTES[0].a/w1823 , \SUBBYTES[0].a/w1822 , \SUBBYTES[0].a/w1821 ,
         \SUBBYTES[0].a/w1820 , \SUBBYTES[0].a/w1819 , \SUBBYTES[0].a/w1817 ,
         \SUBBYTES[0].a/w1816 , \SUBBYTES[0].a/w1744 , \SUBBYTES[0].a/w1742 ,
         \SUBBYTES[0].a/w1741 , \SUBBYTES[0].a/w1740 , \SUBBYTES[0].a/w1737 ,
         \SUBBYTES[0].a/w1735 , \SUBBYTES[0].a/w1734 , \SUBBYTES[0].a/w1733 ,
         \SUBBYTES[0].a/w1729 , \SUBBYTES[0].a/w1727 , \SUBBYTES[0].a/w1726 ,
         \SUBBYTES[0].a/w1725 , \SUBBYTES[0].a/w1724 , \SUBBYTES[0].a/w1723 ,
         \SUBBYTES[0].a/w1722 , \SUBBYTES[0].a/w1721 , \SUBBYTES[0].a/w1720 ,
         \SUBBYTES[0].a/w1712 , \SUBBYTES[0].a/w1710 , \SUBBYTES[0].a/w1709 ,
         \SUBBYTES[0].a/w1705 , \SUBBYTES[0].a/w1703 , \SUBBYTES[0].a/w1702 ,
         \SUBBYTES[0].a/w1701 , \SUBBYTES[0].a/w1697 , \SUBBYTES[0].a/w1695 ,
         \SUBBYTES[0].a/w1694 , \SUBBYTES[0].a/w1681 , \SUBBYTES[0].a/w1680 ,
         \SUBBYTES[0].a/w1679 , \SUBBYTES[0].a/w1677 , \SUBBYTES[0].a/w1674 ,
         \SUBBYTES[0].a/w1673 , \SUBBYTES[0].a/w1671 , \SUBBYTES[0].a/w1670 ,
         \SUBBYTES[0].a/w1668 , \SUBBYTES[0].a/w1666 , \SUBBYTES[0].a/w1665 ,
         \SUBBYTES[0].a/w1659 , \SUBBYTES[0].a/w1658 , \SUBBYTES[0].a/w1657 ,
         \SUBBYTES[0].a/w1656 , \SUBBYTES[0].a/w1650 , \SUBBYTES[0].a/w1648 ,
         \SUBBYTES[0].a/w1647 , \SUBBYTES[0].a/w1643 , \SUBBYTES[0].a/w1641 ,
         \SUBBYTES[0].a/w1640 , \SUBBYTES[0].a/w1635 , \SUBBYTES[0].a/w1633 ,
         \SUBBYTES[0].a/w1632 , \SUBBYTES[0].a/w1616 , \SUBBYTES[0].a/w1615 ,
         \SUBBYTES[0].a/w1614 , \SUBBYTES[0].a/w1613 , \SUBBYTES[0].a/w1612 ,
         \SUBBYTES[0].a/w1610 , \SUBBYTES[0].a/w1609 , \SUBBYTES[0].a/w1537 ,
         \SUBBYTES[0].a/w1535 , \SUBBYTES[0].a/w1534 , \SUBBYTES[0].a/w1533 ,
         \SUBBYTES[0].a/w1530 , \SUBBYTES[0].a/w1528 , \SUBBYTES[0].a/w1527 ,
         \SUBBYTES[0].a/w1526 , \SUBBYTES[0].a/w1522 , \SUBBYTES[0].a/w1520 ,
         \SUBBYTES[0].a/w1519 , \SUBBYTES[0].a/w1518 , \SUBBYTES[0].a/w1517 ,
         \SUBBYTES[0].a/w1516 , \SUBBYTES[0].a/w1515 , \SUBBYTES[0].a/w1514 ,
         \SUBBYTES[0].a/w1513 , \SUBBYTES[0].a/w1505 , \SUBBYTES[0].a/w1503 ,
         \SUBBYTES[0].a/w1502 , \SUBBYTES[0].a/w1498 , \SUBBYTES[0].a/w1496 ,
         \SUBBYTES[0].a/w1495 , \SUBBYTES[0].a/w1494 , \SUBBYTES[0].a/w1490 ,
         \SUBBYTES[0].a/w1488 , \SUBBYTES[0].a/w1487 , \SUBBYTES[0].a/w1474 ,
         \SUBBYTES[0].a/w1473 , \SUBBYTES[0].a/w1472 , \SUBBYTES[0].a/w1470 ,
         \SUBBYTES[0].a/w1467 , \SUBBYTES[0].a/w1466 , \SUBBYTES[0].a/w1464 ,
         \SUBBYTES[0].a/w1463 , \SUBBYTES[0].a/w1461 , \SUBBYTES[0].a/w1459 ,
         \SUBBYTES[0].a/w1458 , \SUBBYTES[0].a/w1452 , \SUBBYTES[0].a/w1451 ,
         \SUBBYTES[0].a/w1450 , \SUBBYTES[0].a/w1449 , \SUBBYTES[0].a/w1443 ,
         \SUBBYTES[0].a/w1441 , \SUBBYTES[0].a/w1440 , \SUBBYTES[0].a/w1436 ,
         \SUBBYTES[0].a/w1434 , \SUBBYTES[0].a/w1433 , \SUBBYTES[0].a/w1428 ,
         \SUBBYTES[0].a/w1426 , \SUBBYTES[0].a/w1425 , \SUBBYTES[0].a/w1409 ,
         \SUBBYTES[0].a/w1408 , \SUBBYTES[0].a/w1407 , \SUBBYTES[0].a/w1406 ,
         \SUBBYTES[0].a/w1405 , \SUBBYTES[0].a/w1403 , \SUBBYTES[0].a/w1402 ,
         \SUBBYTES[0].a/w1330 , \SUBBYTES[0].a/w1328 , \SUBBYTES[0].a/w1327 ,
         \SUBBYTES[0].a/w1326 , \SUBBYTES[0].a/w1323 , \SUBBYTES[0].a/w1321 ,
         \SUBBYTES[0].a/w1320 , \SUBBYTES[0].a/w1319 , \SUBBYTES[0].a/w1315 ,
         \SUBBYTES[0].a/w1313 , \SUBBYTES[0].a/w1312 , \SUBBYTES[0].a/w1311 ,
         \SUBBYTES[0].a/w1310 , \SUBBYTES[0].a/w1309 , \SUBBYTES[0].a/w1308 ,
         \SUBBYTES[0].a/w1307 , \SUBBYTES[0].a/w1306 , \SUBBYTES[0].a/w1298 ,
         \SUBBYTES[0].a/w1296 , \SUBBYTES[0].a/w1295 , \SUBBYTES[0].a/w1291 ,
         \SUBBYTES[0].a/w1289 , \SUBBYTES[0].a/w1288 , \SUBBYTES[0].a/w1287 ,
         \SUBBYTES[0].a/w1283 , \SUBBYTES[0].a/w1281 , \SUBBYTES[0].a/w1280 ,
         \SUBBYTES[0].a/w1267 , \SUBBYTES[0].a/w1266 , \SUBBYTES[0].a/w1265 ,
         \SUBBYTES[0].a/w1263 , \SUBBYTES[0].a/w1260 , \SUBBYTES[0].a/w1259 ,
         \SUBBYTES[0].a/w1257 , \SUBBYTES[0].a/w1256 , \SUBBYTES[0].a/w1254 ,
         \SUBBYTES[0].a/w1252 , \SUBBYTES[0].a/w1251 , \SUBBYTES[0].a/w1245 ,
         \SUBBYTES[0].a/w1244 , \SUBBYTES[0].a/w1243 , \SUBBYTES[0].a/w1242 ,
         \SUBBYTES[0].a/w1236 , \SUBBYTES[0].a/w1234 , \SUBBYTES[0].a/w1233 ,
         \SUBBYTES[0].a/w1229 , \SUBBYTES[0].a/w1227 , \SUBBYTES[0].a/w1226 ,
         \SUBBYTES[0].a/w1221 , \SUBBYTES[0].a/w1219 , \SUBBYTES[0].a/w1218 ,
         \SUBBYTES[0].a/w1202 , \SUBBYTES[0].a/w1201 , \SUBBYTES[0].a/w1200 ,
         \SUBBYTES[0].a/w1199 , \SUBBYTES[0].a/w1198 , \SUBBYTES[0].a/w1196 ,
         \SUBBYTES[0].a/w1195 , \SUBBYTES[0].a/w1123 , \SUBBYTES[0].a/w1121 ,
         \SUBBYTES[0].a/w1120 , \SUBBYTES[0].a/w1119 , \SUBBYTES[0].a/w1116 ,
         \SUBBYTES[0].a/w1114 , \SUBBYTES[0].a/w1113 , \SUBBYTES[0].a/w1112 ,
         \SUBBYTES[0].a/w1108 , \SUBBYTES[0].a/w1106 , \SUBBYTES[0].a/w1105 ,
         \SUBBYTES[0].a/w1104 , \SUBBYTES[0].a/w1103 , \SUBBYTES[0].a/w1102 ,
         \SUBBYTES[0].a/w1101 , \SUBBYTES[0].a/w1100 , \SUBBYTES[0].a/w1099 ,
         \SUBBYTES[0].a/w1091 , \SUBBYTES[0].a/w1089 , \SUBBYTES[0].a/w1088 ,
         \SUBBYTES[0].a/w1084 , \SUBBYTES[0].a/w1082 , \SUBBYTES[0].a/w1081 ,
         \SUBBYTES[0].a/w1080 , \SUBBYTES[0].a/w1076 , \SUBBYTES[0].a/w1074 ,
         \SUBBYTES[0].a/w1073 , \SUBBYTES[0].a/w1060 , \SUBBYTES[0].a/w1059 ,
         \SUBBYTES[0].a/w1058 , \SUBBYTES[0].a/w1056 , \SUBBYTES[0].a/w1053 ,
         \SUBBYTES[0].a/w1052 , \SUBBYTES[0].a/w1050 , \SUBBYTES[0].a/w1049 ,
         \SUBBYTES[0].a/w1047 , \SUBBYTES[0].a/w1045 , \SUBBYTES[0].a/w1044 ,
         \SUBBYTES[0].a/w1038 , \SUBBYTES[0].a/w1037 , \SUBBYTES[0].a/w1036 ,
         \SUBBYTES[0].a/w1035 , \SUBBYTES[0].a/w1029 , \SUBBYTES[0].a/w1027 ,
         \SUBBYTES[0].a/w1026 , \SUBBYTES[0].a/w1022 , \SUBBYTES[0].a/w1020 ,
         \SUBBYTES[0].a/w1019 , \SUBBYTES[0].a/w1014 , \SUBBYTES[0].a/w1012 ,
         \SUBBYTES[0].a/w1011 , \SUBBYTES[0].a/w995 , \SUBBYTES[0].a/w994 ,
         \SUBBYTES[0].a/w993 , \SUBBYTES[0].a/w992 , \SUBBYTES[0].a/w991 ,
         \SUBBYTES[0].a/w989 , \SUBBYTES[0].a/w988 , \SUBBYTES[0].a/w916 ,
         \SUBBYTES[0].a/w914 , \SUBBYTES[0].a/w913 , \SUBBYTES[0].a/w912 ,
         \SUBBYTES[0].a/w909 , \SUBBYTES[0].a/w907 , \SUBBYTES[0].a/w906 ,
         \SUBBYTES[0].a/w905 , \SUBBYTES[0].a/w901 , \SUBBYTES[0].a/w899 ,
         \SUBBYTES[0].a/w898 , \SUBBYTES[0].a/w897 , \SUBBYTES[0].a/w896 ,
         \SUBBYTES[0].a/w895 , \SUBBYTES[0].a/w894 , \SUBBYTES[0].a/w893 ,
         \SUBBYTES[0].a/w892 , \SUBBYTES[0].a/w884 , \SUBBYTES[0].a/w882 ,
         \SUBBYTES[0].a/w881 , \SUBBYTES[0].a/w877 , \SUBBYTES[0].a/w875 ,
         \SUBBYTES[0].a/w874 , \SUBBYTES[0].a/w873 , \SUBBYTES[0].a/w869 ,
         \SUBBYTES[0].a/w867 , \SUBBYTES[0].a/w866 , \SUBBYTES[0].a/w853 ,
         \SUBBYTES[0].a/w852 , \SUBBYTES[0].a/w851 , \SUBBYTES[0].a/w849 ,
         \SUBBYTES[0].a/w846 , \SUBBYTES[0].a/w845 , \SUBBYTES[0].a/w843 ,
         \SUBBYTES[0].a/w842 , \SUBBYTES[0].a/w840 , \SUBBYTES[0].a/w838 ,
         \SUBBYTES[0].a/w837 , \SUBBYTES[0].a/w831 , \SUBBYTES[0].a/w830 ,
         \SUBBYTES[0].a/w829 , \SUBBYTES[0].a/w828 , \SUBBYTES[0].a/w822 ,
         \SUBBYTES[0].a/w820 , \SUBBYTES[0].a/w819 , \SUBBYTES[0].a/w815 ,
         \SUBBYTES[0].a/w813 , \SUBBYTES[0].a/w812 , \SUBBYTES[0].a/w807 ,
         \SUBBYTES[0].a/w805 , \SUBBYTES[0].a/w804 , \SUBBYTES[0].a/w788 ,
         \SUBBYTES[0].a/w787 , \SUBBYTES[0].a/w786 , \SUBBYTES[0].a/w785 ,
         \SUBBYTES[0].a/w784 , \SUBBYTES[0].a/w782 , \SUBBYTES[0].a/w781 ,
         \SUBBYTES[0].a/w709 , \SUBBYTES[0].a/w707 , \SUBBYTES[0].a/w706 ,
         \SUBBYTES[0].a/w705 , \SUBBYTES[0].a/w702 , \SUBBYTES[0].a/w700 ,
         \SUBBYTES[0].a/w699 , \SUBBYTES[0].a/w698 , \SUBBYTES[0].a/w694 ,
         \SUBBYTES[0].a/w692 , \SUBBYTES[0].a/w691 , \SUBBYTES[0].a/w690 ,
         \SUBBYTES[0].a/w689 , \SUBBYTES[0].a/w688 , \SUBBYTES[0].a/w687 ,
         \SUBBYTES[0].a/w686 , \SUBBYTES[0].a/w685 , \SUBBYTES[0].a/w677 ,
         \SUBBYTES[0].a/w675 , \SUBBYTES[0].a/w674 , \SUBBYTES[0].a/w670 ,
         \SUBBYTES[0].a/w668 , \SUBBYTES[0].a/w667 , \SUBBYTES[0].a/w666 ,
         \SUBBYTES[0].a/w662 , \SUBBYTES[0].a/w660 , \SUBBYTES[0].a/w659 ,
         \SUBBYTES[0].a/w646 , \SUBBYTES[0].a/w645 , \SUBBYTES[0].a/w644 ,
         \SUBBYTES[0].a/w642 , \SUBBYTES[0].a/w639 , \SUBBYTES[0].a/w638 ,
         \SUBBYTES[0].a/w636 , \SUBBYTES[0].a/w635 , \SUBBYTES[0].a/w633 ,
         \SUBBYTES[0].a/w631 , \SUBBYTES[0].a/w630 , \SUBBYTES[0].a/w624 ,
         \SUBBYTES[0].a/w623 , \SUBBYTES[0].a/w622 , \SUBBYTES[0].a/w621 ,
         \SUBBYTES[0].a/w615 , \SUBBYTES[0].a/w613 , \SUBBYTES[0].a/w612 ,
         \SUBBYTES[0].a/w608 , \SUBBYTES[0].a/w606 , \SUBBYTES[0].a/w605 ,
         \SUBBYTES[0].a/w600 , \SUBBYTES[0].a/w598 , \SUBBYTES[0].a/w597 ,
         \SUBBYTES[0].a/w581 , \SUBBYTES[0].a/w580 , \SUBBYTES[0].a/w579 ,
         \SUBBYTES[0].a/w578 , \SUBBYTES[0].a/w577 , \SUBBYTES[0].a/w575 ,
         \SUBBYTES[0].a/w574 , \SUBBYTES[0].a/w502 , \SUBBYTES[0].a/w500 ,
         \SUBBYTES[0].a/w499 , \SUBBYTES[0].a/w498 , \SUBBYTES[0].a/w495 ,
         \SUBBYTES[0].a/w493 , \SUBBYTES[0].a/w492 , \SUBBYTES[0].a/w491 ,
         \SUBBYTES[0].a/w487 , \SUBBYTES[0].a/w485 , \SUBBYTES[0].a/w484 ,
         \SUBBYTES[0].a/w483 , \SUBBYTES[0].a/w482 , \SUBBYTES[0].a/w481 ,
         \SUBBYTES[0].a/w480 , \SUBBYTES[0].a/w479 , \SUBBYTES[0].a/w478 ,
         \SUBBYTES[0].a/w470 , \SUBBYTES[0].a/w468 , \SUBBYTES[0].a/w467 ,
         \SUBBYTES[0].a/w463 , \SUBBYTES[0].a/w461 , \SUBBYTES[0].a/w460 ,
         \SUBBYTES[0].a/w459 , \SUBBYTES[0].a/w455 , \SUBBYTES[0].a/w453 ,
         \SUBBYTES[0].a/w452 , \SUBBYTES[0].a/w439 , \SUBBYTES[0].a/w438 ,
         \SUBBYTES[0].a/w437 , \SUBBYTES[0].a/w435 , \SUBBYTES[0].a/w432 ,
         \SUBBYTES[0].a/w431 , \SUBBYTES[0].a/w429 , \SUBBYTES[0].a/w428 ,
         \SUBBYTES[0].a/w426 , \SUBBYTES[0].a/w424 , \SUBBYTES[0].a/w423 ,
         \SUBBYTES[0].a/w417 , \SUBBYTES[0].a/w416 , \SUBBYTES[0].a/w415 ,
         \SUBBYTES[0].a/w414 , \SUBBYTES[0].a/w408 , \SUBBYTES[0].a/w406 ,
         \SUBBYTES[0].a/w405 , \SUBBYTES[0].a/w401 , \SUBBYTES[0].a/w399 ,
         \SUBBYTES[0].a/w398 , \SUBBYTES[0].a/w393 , \SUBBYTES[0].a/w391 ,
         \SUBBYTES[0].a/w390 , \SUBBYTES[0].a/w374 , \SUBBYTES[0].a/w373 ,
         \SUBBYTES[0].a/w372 , \SUBBYTES[0].a/w371 , \SUBBYTES[0].a/w370 ,
         \SUBBYTES[0].a/w368 , \SUBBYTES[0].a/w367 , \SUBBYTES[0].a/w295 ,
         \SUBBYTES[0].a/w293 , \SUBBYTES[0].a/w292 , \SUBBYTES[0].a/w291 ,
         \SUBBYTES[0].a/w288 , \SUBBYTES[0].a/w286 , \SUBBYTES[0].a/w285 ,
         \SUBBYTES[0].a/w284 , \SUBBYTES[0].a/w280 , \SUBBYTES[0].a/w278 ,
         \SUBBYTES[0].a/w277 , \SUBBYTES[0].a/w276 , \SUBBYTES[0].a/w275 ,
         \SUBBYTES[0].a/w274 , \SUBBYTES[0].a/w273 , \SUBBYTES[0].a/w272 ,
         \SUBBYTES[0].a/w271 , \SUBBYTES[0].a/w263 , \SUBBYTES[0].a/w261 ,
         \SUBBYTES[0].a/w260 , \SUBBYTES[0].a/w256 , \SUBBYTES[0].a/w254 ,
         \SUBBYTES[0].a/w253 , \SUBBYTES[0].a/w252 , \SUBBYTES[0].a/w248 ,
         \SUBBYTES[0].a/w246 , \SUBBYTES[0].a/w245 , \SUBBYTES[0].a/w232 ,
         \SUBBYTES[0].a/w231 , \SUBBYTES[0].a/w230 , \SUBBYTES[0].a/w228 ,
         \SUBBYTES[0].a/w225 , \SUBBYTES[0].a/w224 , \SUBBYTES[0].a/w222 ,
         \SUBBYTES[0].a/w221 , \SUBBYTES[0].a/w219 , \SUBBYTES[0].a/w217 ,
         \SUBBYTES[0].a/w216 , \SUBBYTES[0].a/w210 , \SUBBYTES[0].a/w209 ,
         \SUBBYTES[0].a/w208 , \SUBBYTES[0].a/w207 , \SUBBYTES[0].a/w201 ,
         \SUBBYTES[0].a/w199 , \SUBBYTES[0].a/w198 , \SUBBYTES[0].a/w194 ,
         \SUBBYTES[0].a/w192 , \SUBBYTES[0].a/w191 , \SUBBYTES[0].a/w186 ,
         \SUBBYTES[0].a/w184 , \SUBBYTES[0].a/w183 , \SUBBYTES[0].a/w167 ,
         \SUBBYTES[0].a/w166 , \SUBBYTES[0].a/w165 , \SUBBYTES[0].a/w164 ,
         \SUBBYTES[0].a/w163 , \SUBBYTES[0].a/w161 , \SUBBYTES[0].a/w160 , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240;
  wire   [127:0] state;

  DFF \state_reg[127]  ( .D(state[127]), .CLK(clk), .RST(rst), .I(e_init[127]), 
        .Q(state[127]) );
  DFF \state_reg[126]  ( .D(state[126]), .CLK(clk), .RST(rst), .I(e_init[126]), 
        .Q(state[126]) );
  DFF \state_reg[125]  ( .D(state[125]), .CLK(clk), .RST(rst), .I(e_init[125]), 
        .Q(state[125]) );
  DFF \state_reg[124]  ( .D(state[124]), .CLK(clk), .RST(rst), .I(e_init[124]), 
        .Q(state[124]) );
  DFF \state_reg[123]  ( .D(state[123]), .CLK(clk), .RST(rst), .I(e_init[123]), 
        .Q(state[123]) );
  DFF \state_reg[122]  ( .D(state[122]), .CLK(clk), .RST(rst), .I(e_init[122]), 
        .Q(state[122]) );
  DFF \state_reg[121]  ( .D(state[121]), .CLK(clk), .RST(rst), .I(e_init[121]), 
        .Q(state[121]) );
  DFF \state_reg[120]  ( .D(state[120]), .CLK(clk), .RST(rst), .I(e_init[120]), 
        .Q(state[120]) );
  DFF \state_reg[119]  ( .D(state[119]), .CLK(clk), .RST(rst), .I(e_init[119]), 
        .Q(state[119]) );
  DFF \state_reg[118]  ( .D(state[118]), .CLK(clk), .RST(rst), .I(e_init[118]), 
        .Q(state[118]) );
  DFF \state_reg[117]  ( .D(state[117]), .CLK(clk), .RST(rst), .I(e_init[117]), 
        .Q(state[117]) );
  DFF \state_reg[116]  ( .D(state[116]), .CLK(clk), .RST(rst), .I(e_init[116]), 
        .Q(state[116]) );
  DFF \state_reg[115]  ( .D(state[115]), .CLK(clk), .RST(rst), .I(e_init[115]), 
        .Q(state[115]) );
  DFF \state_reg[114]  ( .D(state[114]), .CLK(clk), .RST(rst), .I(e_init[114]), 
        .Q(state[114]) );
  DFF \state_reg[113]  ( .D(state[113]), .CLK(clk), .RST(rst), .I(e_init[113]), 
        .Q(state[113]) );
  DFF \state_reg[112]  ( .D(state[112]), .CLK(clk), .RST(rst), .I(e_init[112]), 
        .Q(state[112]) );
  DFF \state_reg[111]  ( .D(state[111]), .CLK(clk), .RST(rst), .I(e_init[111]), 
        .Q(state[111]) );
  DFF \state_reg[110]  ( .D(state[110]), .CLK(clk), .RST(rst), .I(e_init[110]), 
        .Q(state[110]) );
  DFF \state_reg[109]  ( .D(state[109]), .CLK(clk), .RST(rst), .I(e_init[109]), 
        .Q(state[109]) );
  DFF \state_reg[108]  ( .D(state[108]), .CLK(clk), .RST(rst), .I(e_init[108]), 
        .Q(state[108]) );
  DFF \state_reg[107]  ( .D(state[107]), .CLK(clk), .RST(rst), .I(e_init[107]), 
        .Q(state[107]) );
  DFF \state_reg[106]  ( .D(state[106]), .CLK(clk), .RST(rst), .I(e_init[106]), 
        .Q(state[106]) );
  DFF \state_reg[105]  ( .D(state[105]), .CLK(clk), .RST(rst), .I(e_init[105]), 
        .Q(state[105]) );
  DFF \state_reg[104]  ( .D(state[104]), .CLK(clk), .RST(rst), .I(e_init[104]), 
        .Q(state[104]) );
  DFF \state_reg[103]  ( .D(state[103]), .CLK(clk), .RST(rst), .I(e_init[103]), 
        .Q(state[103]) );
  DFF \state_reg[102]  ( .D(state[102]), .CLK(clk), .RST(rst), .I(e_init[102]), 
        .Q(state[102]) );
  DFF \state_reg[101]  ( .D(state[101]), .CLK(clk), .RST(rst), .I(e_init[101]), 
        .Q(state[101]) );
  DFF \state_reg[100]  ( .D(state[100]), .CLK(clk), .RST(rst), .I(e_init[100]), 
        .Q(state[100]) );
  DFF \state_reg[99]  ( .D(state[99]), .CLK(clk), .RST(rst), .I(e_init[99]), 
        .Q(state[99]) );
  DFF \state_reg[98]  ( .D(state[98]), .CLK(clk), .RST(rst), .I(e_init[98]), 
        .Q(state[98]) );
  DFF \state_reg[97]  ( .D(state[97]), .CLK(clk), .RST(rst), .I(e_init[97]), 
        .Q(state[97]) );
  DFF \state_reg[96]  ( .D(state[96]), .CLK(clk), .RST(rst), .I(e_init[96]), 
        .Q(state[96]) );
  DFF \state_reg[95]  ( .D(state[95]), .CLK(clk), .RST(rst), .I(e_init[95]), 
        .Q(state[95]) );
  DFF \state_reg[94]  ( .D(state[94]), .CLK(clk), .RST(rst), .I(e_init[94]), 
        .Q(state[94]) );
  DFF \state_reg[93]  ( .D(state[93]), .CLK(clk), .RST(rst), .I(e_init[93]), 
        .Q(state[93]) );
  DFF \state_reg[92]  ( .D(state[92]), .CLK(clk), .RST(rst), .I(e_init[92]), 
        .Q(state[92]) );
  DFF \state_reg[91]  ( .D(state[91]), .CLK(clk), .RST(rst), .I(e_init[91]), 
        .Q(state[91]) );
  DFF \state_reg[90]  ( .D(state[90]), .CLK(clk), .RST(rst), .I(e_init[90]), 
        .Q(state[90]) );
  DFF \state_reg[89]  ( .D(state[89]), .CLK(clk), .RST(rst), .I(e_init[89]), 
        .Q(state[89]) );
  DFF \state_reg[88]  ( .D(state[88]), .CLK(clk), .RST(rst), .I(e_init[88]), 
        .Q(state[88]) );
  DFF \state_reg[87]  ( .D(state[87]), .CLK(clk), .RST(rst), .I(e_init[87]), 
        .Q(state[87]) );
  DFF \state_reg[86]  ( .D(state[86]), .CLK(clk), .RST(rst), .I(e_init[86]), 
        .Q(state[86]) );
  DFF \state_reg[85]  ( .D(state[85]), .CLK(clk), .RST(rst), .I(e_init[85]), 
        .Q(state[85]) );
  DFF \state_reg[84]  ( .D(state[84]), .CLK(clk), .RST(rst), .I(e_init[84]), 
        .Q(state[84]) );
  DFF \state_reg[83]  ( .D(state[83]), .CLK(clk), .RST(rst), .I(e_init[83]), 
        .Q(state[83]) );
  DFF \state_reg[82]  ( .D(state[82]), .CLK(clk), .RST(rst), .I(e_init[82]), 
        .Q(state[82]) );
  DFF \state_reg[81]  ( .D(state[81]), .CLK(clk), .RST(rst), .I(e_init[81]), 
        .Q(state[81]) );
  DFF \state_reg[80]  ( .D(state[80]), .CLK(clk), .RST(rst), .I(e_init[80]), 
        .Q(state[80]) );
  DFF \state_reg[79]  ( .D(state[79]), .CLK(clk), .RST(rst), .I(e_init[79]), 
        .Q(state[79]) );
  DFF \state_reg[78]  ( .D(state[78]), .CLK(clk), .RST(rst), .I(e_init[78]), 
        .Q(state[78]) );
  DFF \state_reg[77]  ( .D(state[77]), .CLK(clk), .RST(rst), .I(e_init[77]), 
        .Q(state[77]) );
  DFF \state_reg[76]  ( .D(state[76]), .CLK(clk), .RST(rst), .I(e_init[76]), 
        .Q(state[76]) );
  DFF \state_reg[75]  ( .D(state[75]), .CLK(clk), .RST(rst), .I(e_init[75]), 
        .Q(state[75]) );
  DFF \state_reg[74]  ( .D(state[74]), .CLK(clk), .RST(rst), .I(e_init[74]), 
        .Q(state[74]) );
  DFF \state_reg[73]  ( .D(state[73]), .CLK(clk), .RST(rst), .I(e_init[73]), 
        .Q(state[73]) );
  DFF \state_reg[72]  ( .D(state[72]), .CLK(clk), .RST(rst), .I(e_init[72]), 
        .Q(state[72]) );
  DFF \state_reg[71]  ( .D(state[71]), .CLK(clk), .RST(rst), .I(e_init[71]), 
        .Q(state[71]) );
  DFF \state_reg[70]  ( .D(state[70]), .CLK(clk), .RST(rst), .I(e_init[70]), 
        .Q(state[70]) );
  DFF \state_reg[69]  ( .D(state[69]), .CLK(clk), .RST(rst), .I(e_init[69]), 
        .Q(state[69]) );
  DFF \state_reg[68]  ( .D(state[68]), .CLK(clk), .RST(rst), .I(e_init[68]), 
        .Q(state[68]) );
  DFF \state_reg[67]  ( .D(state[67]), .CLK(clk), .RST(rst), .I(e_init[67]), 
        .Q(state[67]) );
  DFF \state_reg[66]  ( .D(state[66]), .CLK(clk), .RST(rst), .I(e_init[66]), 
        .Q(state[66]) );
  DFF \state_reg[65]  ( .D(state[65]), .CLK(clk), .RST(rst), .I(e_init[65]), 
        .Q(state[65]) );
  DFF \state_reg[64]  ( .D(state[64]), .CLK(clk), .RST(rst), .I(e_init[64]), 
        .Q(state[64]) );
  DFF \state_reg[63]  ( .D(state[63]), .CLK(clk), .RST(rst), .I(e_init[63]), 
        .Q(state[63]) );
  DFF \state_reg[62]  ( .D(state[62]), .CLK(clk), .RST(rst), .I(e_init[62]), 
        .Q(state[62]) );
  DFF \state_reg[61]  ( .D(state[61]), .CLK(clk), .RST(rst), .I(e_init[61]), 
        .Q(state[61]) );
  DFF \state_reg[60]  ( .D(state[60]), .CLK(clk), .RST(rst), .I(e_init[60]), 
        .Q(state[60]) );
  DFF \state_reg[59]  ( .D(state[59]), .CLK(clk), .RST(rst), .I(e_init[59]), 
        .Q(state[59]) );
  DFF \state_reg[58]  ( .D(state[58]), .CLK(clk), .RST(rst), .I(e_init[58]), 
        .Q(state[58]) );
  DFF \state_reg[57]  ( .D(state[57]), .CLK(clk), .RST(rst), .I(e_init[57]), 
        .Q(state[57]) );
  DFF \state_reg[56]  ( .D(state[56]), .CLK(clk), .RST(rst), .I(e_init[56]), 
        .Q(state[56]) );
  DFF \state_reg[55]  ( .D(state[55]), .CLK(clk), .RST(rst), .I(e_init[55]), 
        .Q(state[55]) );
  DFF \state_reg[54]  ( .D(state[54]), .CLK(clk), .RST(rst), .I(e_init[54]), 
        .Q(state[54]) );
  DFF \state_reg[53]  ( .D(state[53]), .CLK(clk), .RST(rst), .I(e_init[53]), 
        .Q(state[53]) );
  DFF \state_reg[52]  ( .D(state[52]), .CLK(clk), .RST(rst), .I(e_init[52]), 
        .Q(state[52]) );
  DFF \state_reg[51]  ( .D(state[51]), .CLK(clk), .RST(rst), .I(e_init[51]), 
        .Q(state[51]) );
  DFF \state_reg[50]  ( .D(state[50]), .CLK(clk), .RST(rst), .I(e_init[50]), 
        .Q(state[50]) );
  DFF \state_reg[49]  ( .D(state[49]), .CLK(clk), .RST(rst), .I(e_init[49]), 
        .Q(state[49]) );
  DFF \state_reg[48]  ( .D(state[48]), .CLK(clk), .RST(rst), .I(e_init[48]), 
        .Q(state[48]) );
  DFF \state_reg[47]  ( .D(state[47]), .CLK(clk), .RST(rst), .I(e_init[47]), 
        .Q(state[47]) );
  DFF \state_reg[46]  ( .D(state[46]), .CLK(clk), .RST(rst), .I(e_init[46]), 
        .Q(state[46]) );
  DFF \state_reg[45]  ( .D(state[45]), .CLK(clk), .RST(rst), .I(e_init[45]), 
        .Q(state[45]) );
  DFF \state_reg[44]  ( .D(state[44]), .CLK(clk), .RST(rst), .I(e_init[44]), 
        .Q(state[44]) );
  DFF \state_reg[43]  ( .D(state[43]), .CLK(clk), .RST(rst), .I(e_init[43]), 
        .Q(state[43]) );
  DFF \state_reg[42]  ( .D(state[42]), .CLK(clk), .RST(rst), .I(e_init[42]), 
        .Q(state[42]) );
  DFF \state_reg[41]  ( .D(state[41]), .CLK(clk), .RST(rst), .I(e_init[41]), 
        .Q(state[41]) );
  DFF \state_reg[40]  ( .D(state[40]), .CLK(clk), .RST(rst), .I(e_init[40]), 
        .Q(state[40]) );
  DFF \state_reg[39]  ( .D(state[39]), .CLK(clk), .RST(rst), .I(e_init[39]), 
        .Q(state[39]) );
  DFF \state_reg[38]  ( .D(state[38]), .CLK(clk), .RST(rst), .I(e_init[38]), 
        .Q(state[38]) );
  DFF \state_reg[37]  ( .D(state[37]), .CLK(clk), .RST(rst), .I(e_init[37]), 
        .Q(state[37]) );
  DFF \state_reg[36]  ( .D(state[36]), .CLK(clk), .RST(rst), .I(e_init[36]), 
        .Q(state[36]) );
  DFF \state_reg[35]  ( .D(state[35]), .CLK(clk), .RST(rst), .I(e_init[35]), 
        .Q(state[35]) );
  DFF \state_reg[34]  ( .D(state[34]), .CLK(clk), .RST(rst), .I(e_init[34]), 
        .Q(state[34]) );
  DFF \state_reg[33]  ( .D(state[33]), .CLK(clk), .RST(rst), .I(e_init[33]), 
        .Q(state[33]) );
  DFF \state_reg[32]  ( .D(state[32]), .CLK(clk), .RST(rst), .I(e_init[32]), 
        .Q(state[32]) );
  DFF \state_reg[31]  ( .D(state[31]), .CLK(clk), .RST(rst), .I(e_init[31]), 
        .Q(state[31]) );
  DFF \state_reg[30]  ( .D(state[30]), .CLK(clk), .RST(rst), .I(e_init[30]), 
        .Q(state[30]) );
  DFF \state_reg[29]  ( .D(state[29]), .CLK(clk), .RST(rst), .I(e_init[29]), 
        .Q(state[29]) );
  DFF \state_reg[28]  ( .D(state[28]), .CLK(clk), .RST(rst), .I(e_init[28]), 
        .Q(state[28]) );
  DFF \state_reg[27]  ( .D(state[27]), .CLK(clk), .RST(rst), .I(e_init[27]), 
        .Q(state[27]) );
  DFF \state_reg[26]  ( .D(state[26]), .CLK(clk), .RST(rst), .I(e_init[26]), 
        .Q(state[26]) );
  DFF \state_reg[25]  ( .D(state[25]), .CLK(clk), .RST(rst), .I(e_init[25]), 
        .Q(state[25]) );
  DFF \state_reg[24]  ( .D(state[24]), .CLK(clk), .RST(rst), .I(e_init[24]), 
        .Q(state[24]) );
  DFF \state_reg[23]  ( .D(state[23]), .CLK(clk), .RST(rst), .I(e_init[23]), 
        .Q(state[23]) );
  DFF \state_reg[22]  ( .D(state[22]), .CLK(clk), .RST(rst), .I(e_init[22]), 
        .Q(state[22]) );
  DFF \state_reg[21]  ( .D(state[21]), .CLK(clk), .RST(rst), .I(e_init[21]), 
        .Q(state[21]) );
  DFF \state_reg[20]  ( .D(state[20]), .CLK(clk), .RST(rst), .I(e_init[20]), 
        .Q(state[20]) );
  DFF \state_reg[19]  ( .D(state[19]), .CLK(clk), .RST(rst), .I(e_init[19]), 
        .Q(state[19]) );
  DFF \state_reg[18]  ( .D(state[18]), .CLK(clk), .RST(rst), .I(e_init[18]), 
        .Q(state[18]) );
  DFF \state_reg[17]  ( .D(state[17]), .CLK(clk), .RST(rst), .I(e_init[17]), 
        .Q(state[17]) );
  DFF \state_reg[16]  ( .D(state[16]), .CLK(clk), .RST(rst), .I(e_init[16]), 
        .Q(state[16]) );
  DFF \state_reg[15]  ( .D(state[15]), .CLK(clk), .RST(rst), .I(e_init[15]), 
        .Q(state[15]) );
  DFF \state_reg[14]  ( .D(state[14]), .CLK(clk), .RST(rst), .I(e_init[14]), 
        .Q(state[14]) );
  DFF \state_reg[13]  ( .D(state[13]), .CLK(clk), .RST(rst), .I(e_init[13]), 
        .Q(state[13]) );
  DFF \state_reg[12]  ( .D(state[12]), .CLK(clk), .RST(rst), .I(e_init[12]), 
        .Q(state[12]) );
  DFF \state_reg[11]  ( .D(state[11]), .CLK(clk), .RST(rst), .I(e_init[11]), 
        .Q(state[11]) );
  DFF \state_reg[10]  ( .D(state[10]), .CLK(clk), .RST(rst), .I(e_init[10]), 
        .Q(state[10]) );
  DFF \state_reg[9]  ( .D(state[9]), .CLK(clk), .RST(rst), .I(e_init[9]), .Q(
        state[9]) );
  DFF \state_reg[8]  ( .D(state[8]), .CLK(clk), .RST(rst), .I(e_init[8]), .Q(
        state[8]) );
  DFF \state_reg[7]  ( .D(state[7]), .CLK(clk), .RST(rst), .I(e_init[7]), .Q(
        state[7]) );
  DFF \state_reg[6]  ( .D(state[6]), .CLK(clk), .RST(rst), .I(e_init[6]), .Q(
        state[6]) );
  DFF \state_reg[5]  ( .D(state[5]), .CLK(clk), .RST(rst), .I(e_init[5]), .Q(
        state[5]) );
  DFF \state_reg[4]  ( .D(state[4]), .CLK(clk), .RST(rst), .I(e_init[4]), .Q(
        state[4]) );
  DFF \state_reg[3]  ( .D(state[3]), .CLK(clk), .RST(rst), .I(e_init[3]), .Q(
        state[3]) );
  DFF \state_reg[2]  ( .D(state[2]), .CLK(clk), .RST(rst), .I(e_init[2]), .Q(
        state[2]) );
  DFF \state_reg[1]  ( .D(state[1]), .CLK(clk), .RST(rst), .I(e_init[1]), .Q(
        state[1]) );
  DFF \state_reg[0]  ( .D(state[0]), .CLK(clk), .RST(rst), .I(e_init[0]), .Q(
        state[0]) );
  XOR \SUBBYTES[0].a/U5649  ( .A(\SUBBYTES[0].a/w3390 ), .B(
        \SUBBYTES[0].a/w3391 ), .Z(\SUBBYTES[0].a/n1426 ) );
  XOR \SUBBYTES[0].a/U5648  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n385 ), .Z(\SUBBYTES[0].a/n1425 ) );
  XOR \SUBBYTES[0].a/U5647  ( .A(\SUBBYTES[0].a/w3383 ), .B(
        \SUBBYTES[0].a/w3400 ), .Z(\SUBBYTES[0].a/n385 ) );
  XOR \SUBBYTES[0].a/U5646  ( .A(\SUBBYTES[0].a/n1425 ), .B(
        \SUBBYTES[0].a/n386 ), .Z(\SUBBYTES[0].a/n1617 ) );
  XOR \SUBBYTES[0].a/U5645  ( .A(\SUBBYTES[0].a/w3382 ), .B(
        \SUBBYTES[0].a/w3397 ), .Z(\SUBBYTES[0].a/n386 ) );
  XOR \SUBBYTES[0].a/U5644  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n387 ), .Z(\SUBBYTES[0].a/n1619 ) );
  XOR \SUBBYTES[0].a/U5643  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n387 ) );
  XOR \SUBBYTES[0].a/U5642  ( .A(\SUBBYTES[0].a/w3359 ), .B(
        \SUBBYTES[0].a/n388 ), .Z(\SUBBYTES[0].a/n1428 ) );
  XOR \SUBBYTES[0].a/U5641  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3351 ), .Z(\SUBBYTES[0].a/n388 ) );
  XOR \SUBBYTES[0].a/U5640  ( .A(\SUBBYTES[0].a/n1428 ), .B(
        \SUBBYTES[0].a/n389 ), .Z(\SUBBYTES[0].a/n1618 ) );
  XOR \SUBBYTES[0].a/U5639  ( .A(\SUBBYTES[0].a/w3361 ), .B(
        \SUBBYTES[0].a/n1619 ), .Z(\SUBBYTES[0].a/n389 ) );
  XOR \SUBBYTES[0].a/U5638  ( .A(\SUBBYTES[0].a/n391 ), .B(
        \SUBBYTES[0].a/n390 ), .Z(\SUBBYTES[0].a/n1429 ) );
  XOR \SUBBYTES[0].a/U5637  ( .A(\SUBBYTES[0].a/n393 ), .B(
        \SUBBYTES[0].a/n392 ), .Z(\SUBBYTES[0].a/n390 ) );
  XOR \SUBBYTES[0].a/U5636  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n391 ) );
  XOR \SUBBYTES[0].a/U5635  ( .A(\SUBBYTES[0].a/w3361 ), .B(
        \SUBBYTES[0].a/w3385 ), .Z(\SUBBYTES[0].a/n392 ) );
  XOR \SUBBYTES[0].a/U5634  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3359 ), .Z(\SUBBYTES[0].a/n393 ) );
  XOR \SUBBYTES[0].a/U5633  ( .A(\SUBBYTES[0].a/w3382 ), .B(
        \SUBBYTES[0].a/n394 ), .Z(\SUBBYTES[0].a/n1427 ) );
  XOR \SUBBYTES[0].a/U5632  ( .A(\SUBBYTES[0].a/w3365 ), .B(
        \SUBBYTES[0].a/w3368 ), .Z(\SUBBYTES[0].a/n394 ) );
  XOR \SUBBYTES[0].a/U5631  ( .A(\SUBBYTES[0].a/n1427 ), .B(
        \SUBBYTES[0].a/n395 ), .Z(\SUBBYTES[0].a/n1620 ) );
  XOR \SUBBYTES[0].a/U5630  ( .A(\SUBBYTES[0].a/w3353 ), .B(
        \SUBBYTES[0].a/n1429 ), .Z(\SUBBYTES[0].a/n395 ) );
  XOR \SUBBYTES[0].a/U5629  ( .A(\SUBBYTES[0].a/n1425 ), .B(
        \SUBBYTES[0].a/n396 ), .Z(\SUBBYTES[0].a/n1621 ) );
  XOR \SUBBYTES[0].a/U5628  ( .A(\SUBBYTES[0].a/w3385 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n396 ) );
  XOR \SUBBYTES[0].a/U5627  ( .A(\SUBBYTES[0].a/n398 ), .B(
        \SUBBYTES[0].a/n397 ), .Z(\SUBBYTES[0].a/n1622 ) );
  XOR \SUBBYTES[0].a/U5626  ( .A(\SUBBYTES[0].a/n400 ), .B(
        \SUBBYTES[0].a/n399 ), .Z(\SUBBYTES[0].a/n397 ) );
  XOR \SUBBYTES[0].a/U5625  ( .A(\SUBBYTES[0].a/n402 ), .B(
        \SUBBYTES[0].a/n401 ), .Z(\SUBBYTES[0].a/n398 ) );
  XOR \SUBBYTES[0].a/U5624  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3400 ), .Z(\SUBBYTES[0].a/n399 ) );
  XOR \SUBBYTES[0].a/U5623  ( .A(\SUBBYTES[0].a/w3390 ), .B(
        \SUBBYTES[0].a/w3393 ), .Z(\SUBBYTES[0].a/n400 ) );
  XOR \SUBBYTES[0].a/U5622  ( .A(\SUBBYTES[0].a/w3365 ), .B(
        \SUBBYTES[0].a/w3366 ), .Z(\SUBBYTES[0].a/n401 ) );
  XOR \SUBBYTES[0].a/U5621  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3353 ), .Z(\SUBBYTES[0].a/n402 ) );
  XOR \SUBBYTES[0].a/U5620  ( .A(\SUBBYTES[0].a/n404 ), .B(
        \SUBBYTES[0].a/n403 ), .Z(\SUBBYTES[0].a/n1623 ) );
  XOR \SUBBYTES[0].a/U5619  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n405 ), .Z(\SUBBYTES[0].a/n403 ) );
  XOR \SUBBYTES[0].a/U5618  ( .A(\SUBBYTES[0].a/n1428 ), .B(
        \SUBBYTES[0].a/n1427 ), .Z(\SUBBYTES[0].a/n404 ) );
  XOR \SUBBYTES[0].a/U5617  ( .A(\SUBBYTES[0].a/w3358 ), .B(
        \SUBBYTES[0].a/w3385 ), .Z(\SUBBYTES[0].a/n405 ) );
  XOR \SUBBYTES[0].a/U5616  ( .A(\SUBBYTES[0].a/n407 ), .B(
        \SUBBYTES[0].a/n406 ), .Z(\SUBBYTES[0].a/n1624 ) );
  XOR \SUBBYTES[0].a/U5615  ( .A(\SUBBYTES[0].a/n1429 ), .B(
        \SUBBYTES[0].a/n408 ), .Z(\SUBBYTES[0].a/n406 ) );
  XOR \SUBBYTES[0].a/U5614  ( .A(\SUBBYTES[0].a/w3391 ), .B(
        \SUBBYTES[0].a/w3393 ), .Z(\SUBBYTES[0].a/n407 ) );
  XOR \SUBBYTES[0].a/U5613  ( .A(\SUBBYTES[0].a/w3351 ), .B(
        \SUBBYTES[0].a/w3383 ), .Z(\SUBBYTES[0].a/n408 ) );
  XOR \SUBBYTES[0].a/U5612  ( .A(\SUBBYTES[0].a/w3183 ), .B(
        \SUBBYTES[0].a/w3184 ), .Z(\SUBBYTES[0].a/n1431 ) );
  XOR \SUBBYTES[0].a/U5611  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n409 ), .Z(\SUBBYTES[0].a/n1430 ) );
  XOR \SUBBYTES[0].a/U5610  ( .A(\SUBBYTES[0].a/w3176 ), .B(
        \SUBBYTES[0].a/w3193 ), .Z(\SUBBYTES[0].a/n409 ) );
  XOR \SUBBYTES[0].a/U5609  ( .A(\SUBBYTES[0].a/n1430 ), .B(
        \SUBBYTES[0].a/n410 ), .Z(\SUBBYTES[0].a/n1625 ) );
  XOR \SUBBYTES[0].a/U5608  ( .A(\SUBBYTES[0].a/w3175 ), .B(
        \SUBBYTES[0].a/w3190 ), .Z(\SUBBYTES[0].a/n410 ) );
  XOR \SUBBYTES[0].a/U5607  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n411 ), .Z(\SUBBYTES[0].a/n1627 ) );
  XOR \SUBBYTES[0].a/U5606  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n411 ) );
  XOR \SUBBYTES[0].a/U5605  ( .A(\SUBBYTES[0].a/w3152 ), .B(
        \SUBBYTES[0].a/n412 ), .Z(\SUBBYTES[0].a/n1433 ) );
  XOR \SUBBYTES[0].a/U5604  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3144 ), .Z(\SUBBYTES[0].a/n412 ) );
  XOR \SUBBYTES[0].a/U5603  ( .A(\SUBBYTES[0].a/n1433 ), .B(
        \SUBBYTES[0].a/n413 ), .Z(\SUBBYTES[0].a/n1626 ) );
  XOR \SUBBYTES[0].a/U5602  ( .A(\SUBBYTES[0].a/w3154 ), .B(
        \SUBBYTES[0].a/n1627 ), .Z(\SUBBYTES[0].a/n413 ) );
  XOR \SUBBYTES[0].a/U5601  ( .A(\SUBBYTES[0].a/n415 ), .B(
        \SUBBYTES[0].a/n414 ), .Z(\SUBBYTES[0].a/n1434 ) );
  XOR \SUBBYTES[0].a/U5600  ( .A(\SUBBYTES[0].a/n417 ), .B(
        \SUBBYTES[0].a/n416 ), .Z(\SUBBYTES[0].a/n414 ) );
  XOR \SUBBYTES[0].a/U5599  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n415 ) );
  XOR \SUBBYTES[0].a/U5598  ( .A(\SUBBYTES[0].a/w3154 ), .B(
        \SUBBYTES[0].a/w3178 ), .Z(\SUBBYTES[0].a/n416 ) );
  XOR \SUBBYTES[0].a/U5597  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3152 ), .Z(\SUBBYTES[0].a/n417 ) );
  XOR \SUBBYTES[0].a/U5596  ( .A(\SUBBYTES[0].a/w3175 ), .B(
        \SUBBYTES[0].a/n418 ), .Z(\SUBBYTES[0].a/n1432 ) );
  XOR \SUBBYTES[0].a/U5595  ( .A(\SUBBYTES[0].a/w3158 ), .B(
        \SUBBYTES[0].a/w3161 ), .Z(\SUBBYTES[0].a/n418 ) );
  XOR \SUBBYTES[0].a/U5594  ( .A(\SUBBYTES[0].a/n1432 ), .B(
        \SUBBYTES[0].a/n419 ), .Z(\SUBBYTES[0].a/n1628 ) );
  XOR \SUBBYTES[0].a/U5593  ( .A(\SUBBYTES[0].a/w3146 ), .B(
        \SUBBYTES[0].a/n1434 ), .Z(\SUBBYTES[0].a/n419 ) );
  XOR \SUBBYTES[0].a/U5592  ( .A(\SUBBYTES[0].a/n1430 ), .B(
        \SUBBYTES[0].a/n420 ), .Z(\SUBBYTES[0].a/n1629 ) );
  XOR \SUBBYTES[0].a/U5591  ( .A(\SUBBYTES[0].a/w3178 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n420 ) );
  XOR \SUBBYTES[0].a/U5590  ( .A(\SUBBYTES[0].a/n422 ), .B(
        \SUBBYTES[0].a/n421 ), .Z(\SUBBYTES[0].a/n1630 ) );
  XOR \SUBBYTES[0].a/U5589  ( .A(\SUBBYTES[0].a/n424 ), .B(
        \SUBBYTES[0].a/n423 ), .Z(\SUBBYTES[0].a/n421 ) );
  XOR \SUBBYTES[0].a/U5588  ( .A(\SUBBYTES[0].a/n426 ), .B(
        \SUBBYTES[0].a/n425 ), .Z(\SUBBYTES[0].a/n422 ) );
  XOR \SUBBYTES[0].a/U5587  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3193 ), .Z(\SUBBYTES[0].a/n423 ) );
  XOR \SUBBYTES[0].a/U5586  ( .A(\SUBBYTES[0].a/w3183 ), .B(
        \SUBBYTES[0].a/w3186 ), .Z(\SUBBYTES[0].a/n424 ) );
  XOR \SUBBYTES[0].a/U5585  ( .A(\SUBBYTES[0].a/w3158 ), .B(
        \SUBBYTES[0].a/w3159 ), .Z(\SUBBYTES[0].a/n425 ) );
  XOR \SUBBYTES[0].a/U5584  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3146 ), .Z(\SUBBYTES[0].a/n426 ) );
  XOR \SUBBYTES[0].a/U5583  ( .A(\SUBBYTES[0].a/n428 ), .B(
        \SUBBYTES[0].a/n427 ), .Z(\SUBBYTES[0].a/n1631 ) );
  XOR \SUBBYTES[0].a/U5582  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n429 ), .Z(\SUBBYTES[0].a/n427 ) );
  XOR \SUBBYTES[0].a/U5581  ( .A(\SUBBYTES[0].a/n1433 ), .B(
        \SUBBYTES[0].a/n1432 ), .Z(\SUBBYTES[0].a/n428 ) );
  XOR \SUBBYTES[0].a/U5580  ( .A(\SUBBYTES[0].a/w3151 ), .B(
        \SUBBYTES[0].a/w3178 ), .Z(\SUBBYTES[0].a/n429 ) );
  XOR \SUBBYTES[0].a/U5579  ( .A(\SUBBYTES[0].a/n431 ), .B(
        \SUBBYTES[0].a/n430 ), .Z(\SUBBYTES[0].a/n1632 ) );
  XOR \SUBBYTES[0].a/U5578  ( .A(\SUBBYTES[0].a/n1434 ), .B(
        \SUBBYTES[0].a/n432 ), .Z(\SUBBYTES[0].a/n430 ) );
  XOR \SUBBYTES[0].a/U5577  ( .A(\SUBBYTES[0].a/w3184 ), .B(
        \SUBBYTES[0].a/w3186 ), .Z(\SUBBYTES[0].a/n431 ) );
  XOR \SUBBYTES[0].a/U5576  ( .A(\SUBBYTES[0].a/w3144 ), .B(
        \SUBBYTES[0].a/w3176 ), .Z(\SUBBYTES[0].a/n432 ) );
  XOR \SUBBYTES[0].a/U5575  ( .A(\SUBBYTES[0].a/w2976 ), .B(
        \SUBBYTES[0].a/w2977 ), .Z(\SUBBYTES[0].a/n1436 ) );
  XOR \SUBBYTES[0].a/U5574  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n433 ), .Z(\SUBBYTES[0].a/n1435 ) );
  XOR \SUBBYTES[0].a/U5573  ( .A(\SUBBYTES[0].a/w2969 ), .B(
        \SUBBYTES[0].a/w2986 ), .Z(\SUBBYTES[0].a/n433 ) );
  XOR \SUBBYTES[0].a/U5572  ( .A(\SUBBYTES[0].a/n1435 ), .B(
        \SUBBYTES[0].a/n434 ), .Z(\SUBBYTES[0].a/n1633 ) );
  XOR \SUBBYTES[0].a/U5571  ( .A(\SUBBYTES[0].a/w2968 ), .B(
        \SUBBYTES[0].a/w2983 ), .Z(\SUBBYTES[0].a/n434 ) );
  XOR \SUBBYTES[0].a/U5570  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n435 ), .Z(\SUBBYTES[0].a/n1635 ) );
  XOR \SUBBYTES[0].a/U5569  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n435 ) );
  XOR \SUBBYTES[0].a/U5568  ( .A(\SUBBYTES[0].a/w2945 ), .B(
        \SUBBYTES[0].a/n436 ), .Z(\SUBBYTES[0].a/n1438 ) );
  XOR \SUBBYTES[0].a/U5567  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2937 ), .Z(\SUBBYTES[0].a/n436 ) );
  XOR \SUBBYTES[0].a/U5566  ( .A(\SUBBYTES[0].a/n1438 ), .B(
        \SUBBYTES[0].a/n437 ), .Z(\SUBBYTES[0].a/n1634 ) );
  XOR \SUBBYTES[0].a/U5565  ( .A(\SUBBYTES[0].a/w2947 ), .B(
        \SUBBYTES[0].a/n1635 ), .Z(\SUBBYTES[0].a/n437 ) );
  XOR \SUBBYTES[0].a/U5564  ( .A(\SUBBYTES[0].a/n439 ), .B(
        \SUBBYTES[0].a/n438 ), .Z(\SUBBYTES[0].a/n1439 ) );
  XOR \SUBBYTES[0].a/U5563  ( .A(\SUBBYTES[0].a/n441 ), .B(
        \SUBBYTES[0].a/n440 ), .Z(\SUBBYTES[0].a/n438 ) );
  XOR \SUBBYTES[0].a/U5562  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n439 ) );
  XOR \SUBBYTES[0].a/U5561  ( .A(\SUBBYTES[0].a/w2947 ), .B(
        \SUBBYTES[0].a/w2971 ), .Z(\SUBBYTES[0].a/n440 ) );
  XOR \SUBBYTES[0].a/U5560  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2945 ), .Z(\SUBBYTES[0].a/n441 ) );
  XOR \SUBBYTES[0].a/U5559  ( .A(\SUBBYTES[0].a/w2968 ), .B(
        \SUBBYTES[0].a/n442 ), .Z(\SUBBYTES[0].a/n1437 ) );
  XOR \SUBBYTES[0].a/U5558  ( .A(\SUBBYTES[0].a/w2951 ), .B(
        \SUBBYTES[0].a/w2954 ), .Z(\SUBBYTES[0].a/n442 ) );
  XOR \SUBBYTES[0].a/U5557  ( .A(\SUBBYTES[0].a/n1437 ), .B(
        \SUBBYTES[0].a/n443 ), .Z(\SUBBYTES[0].a/n1636 ) );
  XOR \SUBBYTES[0].a/U5556  ( .A(\SUBBYTES[0].a/w2939 ), .B(
        \SUBBYTES[0].a/n1439 ), .Z(\SUBBYTES[0].a/n443 ) );
  XOR \SUBBYTES[0].a/U5555  ( .A(\SUBBYTES[0].a/n1435 ), .B(
        \SUBBYTES[0].a/n444 ), .Z(\SUBBYTES[0].a/n1637 ) );
  XOR \SUBBYTES[0].a/U5554  ( .A(\SUBBYTES[0].a/w2971 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n444 ) );
  XOR \SUBBYTES[0].a/U5553  ( .A(\SUBBYTES[0].a/n446 ), .B(
        \SUBBYTES[0].a/n445 ), .Z(\SUBBYTES[0].a/n1638 ) );
  XOR \SUBBYTES[0].a/U5552  ( .A(\SUBBYTES[0].a/n448 ), .B(
        \SUBBYTES[0].a/n447 ), .Z(\SUBBYTES[0].a/n445 ) );
  XOR \SUBBYTES[0].a/U5551  ( .A(\SUBBYTES[0].a/n450 ), .B(
        \SUBBYTES[0].a/n449 ), .Z(\SUBBYTES[0].a/n446 ) );
  XOR \SUBBYTES[0].a/U5550  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2986 ), .Z(\SUBBYTES[0].a/n447 ) );
  XOR \SUBBYTES[0].a/U5549  ( .A(\SUBBYTES[0].a/w2976 ), .B(
        \SUBBYTES[0].a/w2979 ), .Z(\SUBBYTES[0].a/n448 ) );
  XOR \SUBBYTES[0].a/U5548  ( .A(\SUBBYTES[0].a/w2951 ), .B(
        \SUBBYTES[0].a/w2952 ), .Z(\SUBBYTES[0].a/n449 ) );
  XOR \SUBBYTES[0].a/U5547  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2939 ), .Z(\SUBBYTES[0].a/n450 ) );
  XOR \SUBBYTES[0].a/U5546  ( .A(\SUBBYTES[0].a/n452 ), .B(
        \SUBBYTES[0].a/n451 ), .Z(\SUBBYTES[0].a/n1639 ) );
  XOR \SUBBYTES[0].a/U5545  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n453 ), .Z(\SUBBYTES[0].a/n451 ) );
  XOR \SUBBYTES[0].a/U5544  ( .A(\SUBBYTES[0].a/n1438 ), .B(
        \SUBBYTES[0].a/n1437 ), .Z(\SUBBYTES[0].a/n452 ) );
  XOR \SUBBYTES[0].a/U5543  ( .A(\SUBBYTES[0].a/w2944 ), .B(
        \SUBBYTES[0].a/w2971 ), .Z(\SUBBYTES[0].a/n453 ) );
  XOR \SUBBYTES[0].a/U5542  ( .A(\SUBBYTES[0].a/n455 ), .B(
        \SUBBYTES[0].a/n454 ), .Z(\SUBBYTES[0].a/n1640 ) );
  XOR \SUBBYTES[0].a/U5541  ( .A(\SUBBYTES[0].a/n1439 ), .B(
        \SUBBYTES[0].a/n456 ), .Z(\SUBBYTES[0].a/n454 ) );
  XOR \SUBBYTES[0].a/U5540  ( .A(\SUBBYTES[0].a/w2977 ), .B(
        \SUBBYTES[0].a/w2979 ), .Z(\SUBBYTES[0].a/n455 ) );
  XOR \SUBBYTES[0].a/U5539  ( .A(\SUBBYTES[0].a/w2937 ), .B(
        \SUBBYTES[0].a/w2969 ), .Z(\SUBBYTES[0].a/n456 ) );
  XOR \SUBBYTES[0].a/U5538  ( .A(\SUBBYTES[0].a/w2769 ), .B(
        \SUBBYTES[0].a/w2770 ), .Z(\SUBBYTES[0].a/n1441 ) );
  XOR \SUBBYTES[0].a/U5537  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n457 ), .Z(\SUBBYTES[0].a/n1440 ) );
  XOR \SUBBYTES[0].a/U5536  ( .A(\SUBBYTES[0].a/w2762 ), .B(
        \SUBBYTES[0].a/w2779 ), .Z(\SUBBYTES[0].a/n457 ) );
  XOR \SUBBYTES[0].a/U5535  ( .A(\SUBBYTES[0].a/n1440 ), .B(
        \SUBBYTES[0].a/n458 ), .Z(\SUBBYTES[0].a/n1641 ) );
  XOR \SUBBYTES[0].a/U5534  ( .A(\SUBBYTES[0].a/w2761 ), .B(
        \SUBBYTES[0].a/w2776 ), .Z(\SUBBYTES[0].a/n458 ) );
  XOR \SUBBYTES[0].a/U5533  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n459 ), .Z(\SUBBYTES[0].a/n1643 ) );
  XOR \SUBBYTES[0].a/U5532  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n459 ) );
  XOR \SUBBYTES[0].a/U5531  ( .A(\SUBBYTES[0].a/w2738 ), .B(
        \SUBBYTES[0].a/n460 ), .Z(\SUBBYTES[0].a/n1443 ) );
  XOR \SUBBYTES[0].a/U5530  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2730 ), .Z(\SUBBYTES[0].a/n460 ) );
  XOR \SUBBYTES[0].a/U5529  ( .A(\SUBBYTES[0].a/n1443 ), .B(
        \SUBBYTES[0].a/n461 ), .Z(\SUBBYTES[0].a/n1642 ) );
  XOR \SUBBYTES[0].a/U5528  ( .A(\SUBBYTES[0].a/w2740 ), .B(
        \SUBBYTES[0].a/n1643 ), .Z(\SUBBYTES[0].a/n461 ) );
  XOR \SUBBYTES[0].a/U5527  ( .A(\SUBBYTES[0].a/n463 ), .B(
        \SUBBYTES[0].a/n462 ), .Z(\SUBBYTES[0].a/n1444 ) );
  XOR \SUBBYTES[0].a/U5526  ( .A(\SUBBYTES[0].a/n465 ), .B(
        \SUBBYTES[0].a/n464 ), .Z(\SUBBYTES[0].a/n462 ) );
  XOR \SUBBYTES[0].a/U5525  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n463 ) );
  XOR \SUBBYTES[0].a/U5524  ( .A(\SUBBYTES[0].a/w2740 ), .B(
        \SUBBYTES[0].a/w2764 ), .Z(\SUBBYTES[0].a/n464 ) );
  XOR \SUBBYTES[0].a/U5523  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2738 ), .Z(\SUBBYTES[0].a/n465 ) );
  XOR \SUBBYTES[0].a/U5522  ( .A(\SUBBYTES[0].a/w2761 ), .B(
        \SUBBYTES[0].a/n466 ), .Z(\SUBBYTES[0].a/n1442 ) );
  XOR \SUBBYTES[0].a/U5521  ( .A(\SUBBYTES[0].a/w2744 ), .B(
        \SUBBYTES[0].a/w2747 ), .Z(\SUBBYTES[0].a/n466 ) );
  XOR \SUBBYTES[0].a/U5520  ( .A(\SUBBYTES[0].a/n1442 ), .B(
        \SUBBYTES[0].a/n467 ), .Z(\SUBBYTES[0].a/n1644 ) );
  XOR \SUBBYTES[0].a/U5519  ( .A(\SUBBYTES[0].a/w2732 ), .B(
        \SUBBYTES[0].a/n1444 ), .Z(\SUBBYTES[0].a/n467 ) );
  XOR \SUBBYTES[0].a/U5518  ( .A(\SUBBYTES[0].a/n1440 ), .B(
        \SUBBYTES[0].a/n468 ), .Z(\SUBBYTES[0].a/n1645 ) );
  XOR \SUBBYTES[0].a/U5517  ( .A(\SUBBYTES[0].a/w2764 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n468 ) );
  XOR \SUBBYTES[0].a/U5516  ( .A(\SUBBYTES[0].a/n470 ), .B(
        \SUBBYTES[0].a/n469 ), .Z(\SUBBYTES[0].a/n1646 ) );
  XOR \SUBBYTES[0].a/U5515  ( .A(\SUBBYTES[0].a/n472 ), .B(
        \SUBBYTES[0].a/n471 ), .Z(\SUBBYTES[0].a/n469 ) );
  XOR \SUBBYTES[0].a/U5514  ( .A(\SUBBYTES[0].a/n474 ), .B(
        \SUBBYTES[0].a/n473 ), .Z(\SUBBYTES[0].a/n470 ) );
  XOR \SUBBYTES[0].a/U5513  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2779 ), .Z(\SUBBYTES[0].a/n471 ) );
  XOR \SUBBYTES[0].a/U5512  ( .A(\SUBBYTES[0].a/w2769 ), .B(
        \SUBBYTES[0].a/w2772 ), .Z(\SUBBYTES[0].a/n472 ) );
  XOR \SUBBYTES[0].a/U5511  ( .A(\SUBBYTES[0].a/w2744 ), .B(
        \SUBBYTES[0].a/w2745 ), .Z(\SUBBYTES[0].a/n473 ) );
  XOR \SUBBYTES[0].a/U5510  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2732 ), .Z(\SUBBYTES[0].a/n474 ) );
  XOR \SUBBYTES[0].a/U5509  ( .A(\SUBBYTES[0].a/n476 ), .B(
        \SUBBYTES[0].a/n475 ), .Z(\SUBBYTES[0].a/n1647 ) );
  XOR \SUBBYTES[0].a/U5508  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n477 ), .Z(\SUBBYTES[0].a/n475 ) );
  XOR \SUBBYTES[0].a/U5507  ( .A(\SUBBYTES[0].a/n1443 ), .B(
        \SUBBYTES[0].a/n1442 ), .Z(\SUBBYTES[0].a/n476 ) );
  XOR \SUBBYTES[0].a/U5506  ( .A(\SUBBYTES[0].a/w2737 ), .B(
        \SUBBYTES[0].a/w2764 ), .Z(\SUBBYTES[0].a/n477 ) );
  XOR \SUBBYTES[0].a/U5505  ( .A(\SUBBYTES[0].a/n479 ), .B(
        \SUBBYTES[0].a/n478 ), .Z(\SUBBYTES[0].a/n1648 ) );
  XOR \SUBBYTES[0].a/U5504  ( .A(\SUBBYTES[0].a/n1444 ), .B(
        \SUBBYTES[0].a/n480 ), .Z(\SUBBYTES[0].a/n478 ) );
  XOR \SUBBYTES[0].a/U5503  ( .A(\SUBBYTES[0].a/w2770 ), .B(
        \SUBBYTES[0].a/w2772 ), .Z(\SUBBYTES[0].a/n479 ) );
  XOR \SUBBYTES[0].a/U5502  ( .A(\SUBBYTES[0].a/w2730 ), .B(
        \SUBBYTES[0].a/w2762 ), .Z(\SUBBYTES[0].a/n480 ) );
  XOR \SUBBYTES[0].a/U5501  ( .A(\SUBBYTES[0].a/w2562 ), .B(
        \SUBBYTES[0].a/w2563 ), .Z(\SUBBYTES[0].a/n1446 ) );
  XOR \SUBBYTES[0].a/U5500  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n481 ), .Z(\SUBBYTES[0].a/n1445 ) );
  XOR \SUBBYTES[0].a/U5499  ( .A(\SUBBYTES[0].a/w2555 ), .B(
        \SUBBYTES[0].a/w2572 ), .Z(\SUBBYTES[0].a/n481 ) );
  XOR \SUBBYTES[0].a/U5498  ( .A(\SUBBYTES[0].a/n1445 ), .B(
        \SUBBYTES[0].a/n482 ), .Z(\SUBBYTES[0].a/n1649 ) );
  XOR \SUBBYTES[0].a/U5497  ( .A(\SUBBYTES[0].a/w2554 ), .B(
        \SUBBYTES[0].a/w2569 ), .Z(\SUBBYTES[0].a/n482 ) );
  XOR \SUBBYTES[0].a/U5496  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n483 ), .Z(\SUBBYTES[0].a/n1651 ) );
  XOR \SUBBYTES[0].a/U5495  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n483 ) );
  XOR \SUBBYTES[0].a/U5494  ( .A(\SUBBYTES[0].a/w2531 ), .B(
        \SUBBYTES[0].a/n484 ), .Z(\SUBBYTES[0].a/n1448 ) );
  XOR \SUBBYTES[0].a/U5493  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2523 ), .Z(\SUBBYTES[0].a/n484 ) );
  XOR \SUBBYTES[0].a/U5492  ( .A(\SUBBYTES[0].a/n1448 ), .B(
        \SUBBYTES[0].a/n485 ), .Z(\SUBBYTES[0].a/n1650 ) );
  XOR \SUBBYTES[0].a/U5491  ( .A(\SUBBYTES[0].a/w2533 ), .B(
        \SUBBYTES[0].a/n1651 ), .Z(\SUBBYTES[0].a/n485 ) );
  XOR \SUBBYTES[0].a/U5490  ( .A(\SUBBYTES[0].a/n487 ), .B(
        \SUBBYTES[0].a/n486 ), .Z(\SUBBYTES[0].a/n1449 ) );
  XOR \SUBBYTES[0].a/U5489  ( .A(\SUBBYTES[0].a/n489 ), .B(
        \SUBBYTES[0].a/n488 ), .Z(\SUBBYTES[0].a/n486 ) );
  XOR \SUBBYTES[0].a/U5488  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n487 ) );
  XOR \SUBBYTES[0].a/U5487  ( .A(\SUBBYTES[0].a/w2533 ), .B(
        \SUBBYTES[0].a/w2557 ), .Z(\SUBBYTES[0].a/n488 ) );
  XOR \SUBBYTES[0].a/U5486  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2531 ), .Z(\SUBBYTES[0].a/n489 ) );
  XOR \SUBBYTES[0].a/U5485  ( .A(\SUBBYTES[0].a/w2554 ), .B(
        \SUBBYTES[0].a/n490 ), .Z(\SUBBYTES[0].a/n1447 ) );
  XOR \SUBBYTES[0].a/U5484  ( .A(\SUBBYTES[0].a/w2537 ), .B(
        \SUBBYTES[0].a/w2540 ), .Z(\SUBBYTES[0].a/n490 ) );
  XOR \SUBBYTES[0].a/U5483  ( .A(\SUBBYTES[0].a/n1447 ), .B(
        \SUBBYTES[0].a/n491 ), .Z(\SUBBYTES[0].a/n1652 ) );
  XOR \SUBBYTES[0].a/U5482  ( .A(\SUBBYTES[0].a/w2525 ), .B(
        \SUBBYTES[0].a/n1449 ), .Z(\SUBBYTES[0].a/n491 ) );
  XOR \SUBBYTES[0].a/U5481  ( .A(\SUBBYTES[0].a/n1445 ), .B(
        \SUBBYTES[0].a/n492 ), .Z(\SUBBYTES[0].a/n1653 ) );
  XOR \SUBBYTES[0].a/U5480  ( .A(\SUBBYTES[0].a/w2557 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n492 ) );
  XOR \SUBBYTES[0].a/U5479  ( .A(\SUBBYTES[0].a/n494 ), .B(
        \SUBBYTES[0].a/n493 ), .Z(\SUBBYTES[0].a/n1654 ) );
  XOR \SUBBYTES[0].a/U5478  ( .A(\SUBBYTES[0].a/n496 ), .B(
        \SUBBYTES[0].a/n495 ), .Z(\SUBBYTES[0].a/n493 ) );
  XOR \SUBBYTES[0].a/U5477  ( .A(\SUBBYTES[0].a/n498 ), .B(
        \SUBBYTES[0].a/n497 ), .Z(\SUBBYTES[0].a/n494 ) );
  XOR \SUBBYTES[0].a/U5476  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2572 ), .Z(\SUBBYTES[0].a/n495 ) );
  XOR \SUBBYTES[0].a/U5475  ( .A(\SUBBYTES[0].a/w2562 ), .B(
        \SUBBYTES[0].a/w2565 ), .Z(\SUBBYTES[0].a/n496 ) );
  XOR \SUBBYTES[0].a/U5474  ( .A(\SUBBYTES[0].a/w2537 ), .B(
        \SUBBYTES[0].a/w2538 ), .Z(\SUBBYTES[0].a/n497 ) );
  XOR \SUBBYTES[0].a/U5473  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2525 ), .Z(\SUBBYTES[0].a/n498 ) );
  XOR \SUBBYTES[0].a/U5472  ( .A(\SUBBYTES[0].a/n500 ), .B(
        \SUBBYTES[0].a/n499 ), .Z(\SUBBYTES[0].a/n1655 ) );
  XOR \SUBBYTES[0].a/U5471  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n501 ), .Z(\SUBBYTES[0].a/n499 ) );
  XOR \SUBBYTES[0].a/U5470  ( .A(\SUBBYTES[0].a/n1448 ), .B(
        \SUBBYTES[0].a/n1447 ), .Z(\SUBBYTES[0].a/n500 ) );
  XOR \SUBBYTES[0].a/U5469  ( .A(\SUBBYTES[0].a/w2530 ), .B(
        \SUBBYTES[0].a/w2557 ), .Z(\SUBBYTES[0].a/n501 ) );
  XOR \SUBBYTES[0].a/U5468  ( .A(\SUBBYTES[0].a/n503 ), .B(
        \SUBBYTES[0].a/n502 ), .Z(\SUBBYTES[0].a/n1656 ) );
  XOR \SUBBYTES[0].a/U5467  ( .A(\SUBBYTES[0].a/n1449 ), .B(
        \SUBBYTES[0].a/n504 ), .Z(\SUBBYTES[0].a/n502 ) );
  XOR \SUBBYTES[0].a/U5466  ( .A(\SUBBYTES[0].a/w2563 ), .B(
        \SUBBYTES[0].a/w2565 ), .Z(\SUBBYTES[0].a/n503 ) );
  XOR \SUBBYTES[0].a/U5465  ( .A(\SUBBYTES[0].a/w2523 ), .B(
        \SUBBYTES[0].a/w2555 ), .Z(\SUBBYTES[0].a/n504 ) );
  XOR \SUBBYTES[0].a/U5464  ( .A(\SUBBYTES[0].a/w2355 ), .B(
        \SUBBYTES[0].a/w2356 ), .Z(\SUBBYTES[0].a/n1451 ) );
  XOR \SUBBYTES[0].a/U5463  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n505 ), .Z(\SUBBYTES[0].a/n1450 ) );
  XOR \SUBBYTES[0].a/U5462  ( .A(\SUBBYTES[0].a/w2348 ), .B(
        \SUBBYTES[0].a/w2365 ), .Z(\SUBBYTES[0].a/n505 ) );
  XOR \SUBBYTES[0].a/U5461  ( .A(\SUBBYTES[0].a/n1450 ), .B(
        \SUBBYTES[0].a/n506 ), .Z(\SUBBYTES[0].a/n1657 ) );
  XOR \SUBBYTES[0].a/U5460  ( .A(\SUBBYTES[0].a/w2347 ), .B(
        \SUBBYTES[0].a/w2362 ), .Z(\SUBBYTES[0].a/n506 ) );
  XOR \SUBBYTES[0].a/U5459  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n507 ), .Z(\SUBBYTES[0].a/n1659 ) );
  XOR \SUBBYTES[0].a/U5458  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n507 ) );
  XOR \SUBBYTES[0].a/U5457  ( .A(\SUBBYTES[0].a/w2324 ), .B(
        \SUBBYTES[0].a/n508 ), .Z(\SUBBYTES[0].a/n1453 ) );
  XOR \SUBBYTES[0].a/U5456  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2316 ), .Z(\SUBBYTES[0].a/n508 ) );
  XOR \SUBBYTES[0].a/U5455  ( .A(\SUBBYTES[0].a/n1453 ), .B(
        \SUBBYTES[0].a/n509 ), .Z(\SUBBYTES[0].a/n1658 ) );
  XOR \SUBBYTES[0].a/U5454  ( .A(\SUBBYTES[0].a/w2326 ), .B(
        \SUBBYTES[0].a/n1659 ), .Z(\SUBBYTES[0].a/n509 ) );
  XOR \SUBBYTES[0].a/U5453  ( .A(\SUBBYTES[0].a/n511 ), .B(
        \SUBBYTES[0].a/n510 ), .Z(\SUBBYTES[0].a/n1454 ) );
  XOR \SUBBYTES[0].a/U5452  ( .A(\SUBBYTES[0].a/n513 ), .B(
        \SUBBYTES[0].a/n512 ), .Z(\SUBBYTES[0].a/n510 ) );
  XOR \SUBBYTES[0].a/U5451  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n511 ) );
  XOR \SUBBYTES[0].a/U5450  ( .A(\SUBBYTES[0].a/w2326 ), .B(
        \SUBBYTES[0].a/w2350 ), .Z(\SUBBYTES[0].a/n512 ) );
  XOR \SUBBYTES[0].a/U5449  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2324 ), .Z(\SUBBYTES[0].a/n513 ) );
  XOR \SUBBYTES[0].a/U5448  ( .A(\SUBBYTES[0].a/w2347 ), .B(
        \SUBBYTES[0].a/n514 ), .Z(\SUBBYTES[0].a/n1452 ) );
  XOR \SUBBYTES[0].a/U5447  ( .A(\SUBBYTES[0].a/w2330 ), .B(
        \SUBBYTES[0].a/w2333 ), .Z(\SUBBYTES[0].a/n514 ) );
  XOR \SUBBYTES[0].a/U5446  ( .A(\SUBBYTES[0].a/n1452 ), .B(
        \SUBBYTES[0].a/n515 ), .Z(\SUBBYTES[0].a/n1660 ) );
  XOR \SUBBYTES[0].a/U5445  ( .A(\SUBBYTES[0].a/w2318 ), .B(
        \SUBBYTES[0].a/n1454 ), .Z(\SUBBYTES[0].a/n515 ) );
  XOR \SUBBYTES[0].a/U5444  ( .A(\SUBBYTES[0].a/n1450 ), .B(
        \SUBBYTES[0].a/n516 ), .Z(\SUBBYTES[0].a/n1661 ) );
  XOR \SUBBYTES[0].a/U5443  ( .A(\SUBBYTES[0].a/w2350 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n516 ) );
  XOR \SUBBYTES[0].a/U5442  ( .A(\SUBBYTES[0].a/n518 ), .B(
        \SUBBYTES[0].a/n517 ), .Z(\SUBBYTES[0].a/n1662 ) );
  XOR \SUBBYTES[0].a/U5441  ( .A(\SUBBYTES[0].a/n520 ), .B(
        \SUBBYTES[0].a/n519 ), .Z(\SUBBYTES[0].a/n517 ) );
  XOR \SUBBYTES[0].a/U5440  ( .A(\SUBBYTES[0].a/n522 ), .B(
        \SUBBYTES[0].a/n521 ), .Z(\SUBBYTES[0].a/n518 ) );
  XOR \SUBBYTES[0].a/U5439  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2365 ), .Z(\SUBBYTES[0].a/n519 ) );
  XOR \SUBBYTES[0].a/U5438  ( .A(\SUBBYTES[0].a/w2355 ), .B(
        \SUBBYTES[0].a/w2358 ), .Z(\SUBBYTES[0].a/n520 ) );
  XOR \SUBBYTES[0].a/U5437  ( .A(\SUBBYTES[0].a/w2330 ), .B(
        \SUBBYTES[0].a/w2331 ), .Z(\SUBBYTES[0].a/n521 ) );
  XOR \SUBBYTES[0].a/U5436  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2318 ), .Z(\SUBBYTES[0].a/n522 ) );
  XOR \SUBBYTES[0].a/U5435  ( .A(\SUBBYTES[0].a/n524 ), .B(
        \SUBBYTES[0].a/n523 ), .Z(\SUBBYTES[0].a/n1663 ) );
  XOR \SUBBYTES[0].a/U5434  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n525 ), .Z(\SUBBYTES[0].a/n523 ) );
  XOR \SUBBYTES[0].a/U5433  ( .A(\SUBBYTES[0].a/n1453 ), .B(
        \SUBBYTES[0].a/n1452 ), .Z(\SUBBYTES[0].a/n524 ) );
  XOR \SUBBYTES[0].a/U5432  ( .A(\SUBBYTES[0].a/w2323 ), .B(
        \SUBBYTES[0].a/w2350 ), .Z(\SUBBYTES[0].a/n525 ) );
  XOR \SUBBYTES[0].a/U5431  ( .A(\SUBBYTES[0].a/n527 ), .B(
        \SUBBYTES[0].a/n526 ), .Z(\SUBBYTES[0].a/n1664 ) );
  XOR \SUBBYTES[0].a/U5430  ( .A(\SUBBYTES[0].a/n1454 ), .B(
        \SUBBYTES[0].a/n528 ), .Z(\SUBBYTES[0].a/n526 ) );
  XOR \SUBBYTES[0].a/U5429  ( .A(\SUBBYTES[0].a/w2356 ), .B(
        \SUBBYTES[0].a/w2358 ), .Z(\SUBBYTES[0].a/n527 ) );
  XOR \SUBBYTES[0].a/U5428  ( .A(\SUBBYTES[0].a/w2316 ), .B(
        \SUBBYTES[0].a/w2348 ), .Z(\SUBBYTES[0].a/n528 ) );
  XOR \SUBBYTES[0].a/U5427  ( .A(\SUBBYTES[0].a/w2148 ), .B(
        \SUBBYTES[0].a/w2149 ), .Z(\SUBBYTES[0].a/n1456 ) );
  XOR \SUBBYTES[0].a/U5426  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n529 ), .Z(\SUBBYTES[0].a/n1455 ) );
  XOR \SUBBYTES[0].a/U5425  ( .A(\SUBBYTES[0].a/w2141 ), .B(
        \SUBBYTES[0].a/w2158 ), .Z(\SUBBYTES[0].a/n529 ) );
  XOR \SUBBYTES[0].a/U5424  ( .A(\SUBBYTES[0].a/n1455 ), .B(
        \SUBBYTES[0].a/n530 ), .Z(\SUBBYTES[0].a/n1665 ) );
  XOR \SUBBYTES[0].a/U5423  ( .A(\SUBBYTES[0].a/w2140 ), .B(
        \SUBBYTES[0].a/w2155 ), .Z(\SUBBYTES[0].a/n530 ) );
  XOR \SUBBYTES[0].a/U5422  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n531 ), .Z(\SUBBYTES[0].a/n1667 ) );
  XOR \SUBBYTES[0].a/U5421  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n531 ) );
  XOR \SUBBYTES[0].a/U5420  ( .A(\SUBBYTES[0].a/w2117 ), .B(
        \SUBBYTES[0].a/n532 ), .Z(\SUBBYTES[0].a/n1458 ) );
  XOR \SUBBYTES[0].a/U5419  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2109 ), .Z(\SUBBYTES[0].a/n532 ) );
  XOR \SUBBYTES[0].a/U5418  ( .A(\SUBBYTES[0].a/n1458 ), .B(
        \SUBBYTES[0].a/n533 ), .Z(\SUBBYTES[0].a/n1666 ) );
  XOR \SUBBYTES[0].a/U5417  ( .A(\SUBBYTES[0].a/w2119 ), .B(
        \SUBBYTES[0].a/n1667 ), .Z(\SUBBYTES[0].a/n533 ) );
  XOR \SUBBYTES[0].a/U5416  ( .A(\SUBBYTES[0].a/n535 ), .B(
        \SUBBYTES[0].a/n534 ), .Z(\SUBBYTES[0].a/n1459 ) );
  XOR \SUBBYTES[0].a/U5415  ( .A(\SUBBYTES[0].a/n537 ), .B(
        \SUBBYTES[0].a/n536 ), .Z(\SUBBYTES[0].a/n534 ) );
  XOR \SUBBYTES[0].a/U5414  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n535 ) );
  XOR \SUBBYTES[0].a/U5413  ( .A(\SUBBYTES[0].a/w2119 ), .B(
        \SUBBYTES[0].a/w2143 ), .Z(\SUBBYTES[0].a/n536 ) );
  XOR \SUBBYTES[0].a/U5412  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2117 ), .Z(\SUBBYTES[0].a/n537 ) );
  XOR \SUBBYTES[0].a/U5411  ( .A(\SUBBYTES[0].a/w2140 ), .B(
        \SUBBYTES[0].a/n538 ), .Z(\SUBBYTES[0].a/n1457 ) );
  XOR \SUBBYTES[0].a/U5410  ( .A(\SUBBYTES[0].a/w2123 ), .B(
        \SUBBYTES[0].a/w2126 ), .Z(\SUBBYTES[0].a/n538 ) );
  XOR \SUBBYTES[0].a/U5409  ( .A(\SUBBYTES[0].a/n1457 ), .B(
        \SUBBYTES[0].a/n539 ), .Z(\SUBBYTES[0].a/n1668 ) );
  XOR \SUBBYTES[0].a/U5408  ( .A(\SUBBYTES[0].a/w2111 ), .B(
        \SUBBYTES[0].a/n1459 ), .Z(\SUBBYTES[0].a/n539 ) );
  XOR \SUBBYTES[0].a/U5407  ( .A(\SUBBYTES[0].a/n1455 ), .B(
        \SUBBYTES[0].a/n540 ), .Z(\SUBBYTES[0].a/n1669 ) );
  XOR \SUBBYTES[0].a/U5406  ( .A(\SUBBYTES[0].a/w2143 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n540 ) );
  XOR \SUBBYTES[0].a/U5405  ( .A(\SUBBYTES[0].a/n542 ), .B(
        \SUBBYTES[0].a/n541 ), .Z(\SUBBYTES[0].a/n1670 ) );
  XOR \SUBBYTES[0].a/U5404  ( .A(\SUBBYTES[0].a/n544 ), .B(
        \SUBBYTES[0].a/n543 ), .Z(\SUBBYTES[0].a/n541 ) );
  XOR \SUBBYTES[0].a/U5403  ( .A(\SUBBYTES[0].a/n546 ), .B(
        \SUBBYTES[0].a/n545 ), .Z(\SUBBYTES[0].a/n542 ) );
  XOR \SUBBYTES[0].a/U5402  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2158 ), .Z(\SUBBYTES[0].a/n543 ) );
  XOR \SUBBYTES[0].a/U5401  ( .A(\SUBBYTES[0].a/w2148 ), .B(
        \SUBBYTES[0].a/w2151 ), .Z(\SUBBYTES[0].a/n544 ) );
  XOR \SUBBYTES[0].a/U5400  ( .A(\SUBBYTES[0].a/w2123 ), .B(
        \SUBBYTES[0].a/w2124 ), .Z(\SUBBYTES[0].a/n545 ) );
  XOR \SUBBYTES[0].a/U5399  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2111 ), .Z(\SUBBYTES[0].a/n546 ) );
  XOR \SUBBYTES[0].a/U5398  ( .A(\SUBBYTES[0].a/n548 ), .B(
        \SUBBYTES[0].a/n547 ), .Z(\SUBBYTES[0].a/n1671 ) );
  XOR \SUBBYTES[0].a/U5397  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n549 ), .Z(\SUBBYTES[0].a/n547 ) );
  XOR \SUBBYTES[0].a/U5396  ( .A(\SUBBYTES[0].a/n1458 ), .B(
        \SUBBYTES[0].a/n1457 ), .Z(\SUBBYTES[0].a/n548 ) );
  XOR \SUBBYTES[0].a/U5395  ( .A(\SUBBYTES[0].a/w2116 ), .B(
        \SUBBYTES[0].a/w2143 ), .Z(\SUBBYTES[0].a/n549 ) );
  XOR \SUBBYTES[0].a/U5394  ( .A(\SUBBYTES[0].a/n551 ), .B(
        \SUBBYTES[0].a/n550 ), .Z(\SUBBYTES[0].a/n1672 ) );
  XOR \SUBBYTES[0].a/U5393  ( .A(\SUBBYTES[0].a/n1459 ), .B(
        \SUBBYTES[0].a/n552 ), .Z(\SUBBYTES[0].a/n550 ) );
  XOR \SUBBYTES[0].a/U5392  ( .A(\SUBBYTES[0].a/w2149 ), .B(
        \SUBBYTES[0].a/w2151 ), .Z(\SUBBYTES[0].a/n551 ) );
  XOR \SUBBYTES[0].a/U5391  ( .A(\SUBBYTES[0].a/w2109 ), .B(
        \SUBBYTES[0].a/w2141 ), .Z(\SUBBYTES[0].a/n552 ) );
  XOR \SUBBYTES[0].a/U5390  ( .A(\SUBBYTES[0].a/w1941 ), .B(
        \SUBBYTES[0].a/w1942 ), .Z(\SUBBYTES[0].a/n1461 ) );
  XOR \SUBBYTES[0].a/U5389  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n553 ), .Z(\SUBBYTES[0].a/n1460 ) );
  XOR \SUBBYTES[0].a/U5388  ( .A(\SUBBYTES[0].a/w1934 ), .B(
        \SUBBYTES[0].a/w1951 ), .Z(\SUBBYTES[0].a/n553 ) );
  XOR \SUBBYTES[0].a/U5387  ( .A(\SUBBYTES[0].a/n1460 ), .B(
        \SUBBYTES[0].a/n554 ), .Z(\SUBBYTES[0].a/n1673 ) );
  XOR \SUBBYTES[0].a/U5386  ( .A(\SUBBYTES[0].a/w1933 ), .B(
        \SUBBYTES[0].a/w1948 ), .Z(\SUBBYTES[0].a/n554 ) );
  XOR \SUBBYTES[0].a/U5385  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n555 ), .Z(\SUBBYTES[0].a/n1675 ) );
  XOR \SUBBYTES[0].a/U5384  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n555 ) );
  XOR \SUBBYTES[0].a/U5383  ( .A(\SUBBYTES[0].a/w1910 ), .B(
        \SUBBYTES[0].a/n556 ), .Z(\SUBBYTES[0].a/n1463 ) );
  XOR \SUBBYTES[0].a/U5382  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1902 ), .Z(\SUBBYTES[0].a/n556 ) );
  XOR \SUBBYTES[0].a/U5381  ( .A(\SUBBYTES[0].a/n1463 ), .B(
        \SUBBYTES[0].a/n557 ), .Z(\SUBBYTES[0].a/n1674 ) );
  XOR \SUBBYTES[0].a/U5380  ( .A(\SUBBYTES[0].a/w1912 ), .B(
        \SUBBYTES[0].a/n1675 ), .Z(\SUBBYTES[0].a/n557 ) );
  XOR \SUBBYTES[0].a/U5379  ( .A(\SUBBYTES[0].a/n559 ), .B(
        \SUBBYTES[0].a/n558 ), .Z(\SUBBYTES[0].a/n1464 ) );
  XOR \SUBBYTES[0].a/U5378  ( .A(\SUBBYTES[0].a/n561 ), .B(
        \SUBBYTES[0].a/n560 ), .Z(\SUBBYTES[0].a/n558 ) );
  XOR \SUBBYTES[0].a/U5377  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n559 ) );
  XOR \SUBBYTES[0].a/U5376  ( .A(\SUBBYTES[0].a/w1912 ), .B(
        \SUBBYTES[0].a/w1936 ), .Z(\SUBBYTES[0].a/n560 ) );
  XOR \SUBBYTES[0].a/U5375  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1910 ), .Z(\SUBBYTES[0].a/n561 ) );
  XOR \SUBBYTES[0].a/U5374  ( .A(\SUBBYTES[0].a/w1933 ), .B(
        \SUBBYTES[0].a/n562 ), .Z(\SUBBYTES[0].a/n1462 ) );
  XOR \SUBBYTES[0].a/U5373  ( .A(\SUBBYTES[0].a/w1916 ), .B(
        \SUBBYTES[0].a/w1919 ), .Z(\SUBBYTES[0].a/n562 ) );
  XOR \SUBBYTES[0].a/U5372  ( .A(\SUBBYTES[0].a/n1462 ), .B(
        \SUBBYTES[0].a/n563 ), .Z(\SUBBYTES[0].a/n1676 ) );
  XOR \SUBBYTES[0].a/U5371  ( .A(\SUBBYTES[0].a/w1904 ), .B(
        \SUBBYTES[0].a/n1464 ), .Z(\SUBBYTES[0].a/n563 ) );
  XOR \SUBBYTES[0].a/U5370  ( .A(\SUBBYTES[0].a/n1460 ), .B(
        \SUBBYTES[0].a/n564 ), .Z(\SUBBYTES[0].a/n1677 ) );
  XOR \SUBBYTES[0].a/U5369  ( .A(\SUBBYTES[0].a/w1936 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n564 ) );
  XOR \SUBBYTES[0].a/U5368  ( .A(\SUBBYTES[0].a/n566 ), .B(
        \SUBBYTES[0].a/n565 ), .Z(\SUBBYTES[0].a/n1678 ) );
  XOR \SUBBYTES[0].a/U5367  ( .A(\SUBBYTES[0].a/n568 ), .B(
        \SUBBYTES[0].a/n567 ), .Z(\SUBBYTES[0].a/n565 ) );
  XOR \SUBBYTES[0].a/U5366  ( .A(\SUBBYTES[0].a/n570 ), .B(
        \SUBBYTES[0].a/n569 ), .Z(\SUBBYTES[0].a/n566 ) );
  XOR \SUBBYTES[0].a/U5365  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1951 ), .Z(\SUBBYTES[0].a/n567 ) );
  XOR \SUBBYTES[0].a/U5364  ( .A(\SUBBYTES[0].a/w1941 ), .B(
        \SUBBYTES[0].a/w1944 ), .Z(\SUBBYTES[0].a/n568 ) );
  XOR \SUBBYTES[0].a/U5363  ( .A(\SUBBYTES[0].a/w1916 ), .B(
        \SUBBYTES[0].a/w1917 ), .Z(\SUBBYTES[0].a/n569 ) );
  XOR \SUBBYTES[0].a/U5362  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1904 ), .Z(\SUBBYTES[0].a/n570 ) );
  XOR \SUBBYTES[0].a/U5361  ( .A(\SUBBYTES[0].a/n572 ), .B(
        \SUBBYTES[0].a/n571 ), .Z(\SUBBYTES[0].a/n1679 ) );
  XOR \SUBBYTES[0].a/U5360  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n573 ), .Z(\SUBBYTES[0].a/n571 ) );
  XOR \SUBBYTES[0].a/U5359  ( .A(\SUBBYTES[0].a/n1463 ), .B(
        \SUBBYTES[0].a/n1462 ), .Z(\SUBBYTES[0].a/n572 ) );
  XOR \SUBBYTES[0].a/U5358  ( .A(\SUBBYTES[0].a/w1909 ), .B(
        \SUBBYTES[0].a/w1936 ), .Z(\SUBBYTES[0].a/n573 ) );
  XOR \SUBBYTES[0].a/U5357  ( .A(\SUBBYTES[0].a/n575 ), .B(
        \SUBBYTES[0].a/n574 ), .Z(\SUBBYTES[0].a/n1680 ) );
  XOR \SUBBYTES[0].a/U5356  ( .A(\SUBBYTES[0].a/n1464 ), .B(
        \SUBBYTES[0].a/n576 ), .Z(\SUBBYTES[0].a/n574 ) );
  XOR \SUBBYTES[0].a/U5355  ( .A(\SUBBYTES[0].a/w1942 ), .B(
        \SUBBYTES[0].a/w1944 ), .Z(\SUBBYTES[0].a/n575 ) );
  XOR \SUBBYTES[0].a/U5354  ( .A(\SUBBYTES[0].a/w1902 ), .B(
        \SUBBYTES[0].a/w1934 ), .Z(\SUBBYTES[0].a/n576 ) );
  XOR \SUBBYTES[0].a/U5353  ( .A(\SUBBYTES[0].a/w1734 ), .B(
        \SUBBYTES[0].a/w1735 ), .Z(\SUBBYTES[0].a/n1466 ) );
  XOR \SUBBYTES[0].a/U5352  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n577 ), .Z(\SUBBYTES[0].a/n1465 ) );
  XOR \SUBBYTES[0].a/U5351  ( .A(\SUBBYTES[0].a/w1727 ), .B(
        \SUBBYTES[0].a/w1744 ), .Z(\SUBBYTES[0].a/n577 ) );
  XOR \SUBBYTES[0].a/U5350  ( .A(\SUBBYTES[0].a/n1465 ), .B(
        \SUBBYTES[0].a/n578 ), .Z(\SUBBYTES[0].a/n1681 ) );
  XOR \SUBBYTES[0].a/U5349  ( .A(\SUBBYTES[0].a/w1726 ), .B(
        \SUBBYTES[0].a/w1741 ), .Z(\SUBBYTES[0].a/n578 ) );
  XOR \SUBBYTES[0].a/U5348  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n579 ), .Z(\SUBBYTES[0].a/n1683 ) );
  XOR \SUBBYTES[0].a/U5347  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n579 ) );
  XOR \SUBBYTES[0].a/U5346  ( .A(\SUBBYTES[0].a/w1703 ), .B(
        \SUBBYTES[0].a/n580 ), .Z(\SUBBYTES[0].a/n1468 ) );
  XOR \SUBBYTES[0].a/U5345  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1695 ), .Z(\SUBBYTES[0].a/n580 ) );
  XOR \SUBBYTES[0].a/U5344  ( .A(\SUBBYTES[0].a/n1468 ), .B(
        \SUBBYTES[0].a/n581 ), .Z(\SUBBYTES[0].a/n1682 ) );
  XOR \SUBBYTES[0].a/U5343  ( .A(\SUBBYTES[0].a/w1705 ), .B(
        \SUBBYTES[0].a/n1683 ), .Z(\SUBBYTES[0].a/n581 ) );
  XOR \SUBBYTES[0].a/U5342  ( .A(\SUBBYTES[0].a/n583 ), .B(
        \SUBBYTES[0].a/n582 ), .Z(\SUBBYTES[0].a/n1469 ) );
  XOR \SUBBYTES[0].a/U5341  ( .A(\SUBBYTES[0].a/n585 ), .B(
        \SUBBYTES[0].a/n584 ), .Z(\SUBBYTES[0].a/n582 ) );
  XOR \SUBBYTES[0].a/U5340  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n583 ) );
  XOR \SUBBYTES[0].a/U5339  ( .A(\SUBBYTES[0].a/w1705 ), .B(
        \SUBBYTES[0].a/w1729 ), .Z(\SUBBYTES[0].a/n584 ) );
  XOR \SUBBYTES[0].a/U5338  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1703 ), .Z(\SUBBYTES[0].a/n585 ) );
  XOR \SUBBYTES[0].a/U5337  ( .A(\SUBBYTES[0].a/w1726 ), .B(
        \SUBBYTES[0].a/n586 ), .Z(\SUBBYTES[0].a/n1467 ) );
  XOR \SUBBYTES[0].a/U5336  ( .A(\SUBBYTES[0].a/w1709 ), .B(
        \SUBBYTES[0].a/w1712 ), .Z(\SUBBYTES[0].a/n586 ) );
  XOR \SUBBYTES[0].a/U5335  ( .A(\SUBBYTES[0].a/n1467 ), .B(
        \SUBBYTES[0].a/n587 ), .Z(\SUBBYTES[0].a/n1684 ) );
  XOR \SUBBYTES[0].a/U5334  ( .A(\SUBBYTES[0].a/w1697 ), .B(
        \SUBBYTES[0].a/n1469 ), .Z(\SUBBYTES[0].a/n587 ) );
  XOR \SUBBYTES[0].a/U5333  ( .A(\SUBBYTES[0].a/n1465 ), .B(
        \SUBBYTES[0].a/n588 ), .Z(\SUBBYTES[0].a/n1685 ) );
  XOR \SUBBYTES[0].a/U5332  ( .A(\SUBBYTES[0].a/w1729 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n588 ) );
  XOR \SUBBYTES[0].a/U5331  ( .A(\SUBBYTES[0].a/n590 ), .B(
        \SUBBYTES[0].a/n589 ), .Z(\SUBBYTES[0].a/n1686 ) );
  XOR \SUBBYTES[0].a/U5330  ( .A(\SUBBYTES[0].a/n592 ), .B(
        \SUBBYTES[0].a/n591 ), .Z(\SUBBYTES[0].a/n589 ) );
  XOR \SUBBYTES[0].a/U5329  ( .A(\SUBBYTES[0].a/n594 ), .B(
        \SUBBYTES[0].a/n593 ), .Z(\SUBBYTES[0].a/n590 ) );
  XOR \SUBBYTES[0].a/U5328  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1744 ), .Z(\SUBBYTES[0].a/n591 ) );
  XOR \SUBBYTES[0].a/U5327  ( .A(\SUBBYTES[0].a/w1734 ), .B(
        \SUBBYTES[0].a/w1737 ), .Z(\SUBBYTES[0].a/n592 ) );
  XOR \SUBBYTES[0].a/U5326  ( .A(\SUBBYTES[0].a/w1709 ), .B(
        \SUBBYTES[0].a/w1710 ), .Z(\SUBBYTES[0].a/n593 ) );
  XOR \SUBBYTES[0].a/U5325  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1697 ), .Z(\SUBBYTES[0].a/n594 ) );
  XOR \SUBBYTES[0].a/U5324  ( .A(\SUBBYTES[0].a/n596 ), .B(
        \SUBBYTES[0].a/n595 ), .Z(\SUBBYTES[0].a/n1687 ) );
  XOR \SUBBYTES[0].a/U5323  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n597 ), .Z(\SUBBYTES[0].a/n595 ) );
  XOR \SUBBYTES[0].a/U5322  ( .A(\SUBBYTES[0].a/n1468 ), .B(
        \SUBBYTES[0].a/n1467 ), .Z(\SUBBYTES[0].a/n596 ) );
  XOR \SUBBYTES[0].a/U5321  ( .A(\SUBBYTES[0].a/w1702 ), .B(
        \SUBBYTES[0].a/w1729 ), .Z(\SUBBYTES[0].a/n597 ) );
  XOR \SUBBYTES[0].a/U5320  ( .A(\SUBBYTES[0].a/n599 ), .B(
        \SUBBYTES[0].a/n598 ), .Z(\SUBBYTES[0].a/n1688 ) );
  XOR \SUBBYTES[0].a/U5319  ( .A(\SUBBYTES[0].a/n1469 ), .B(
        \SUBBYTES[0].a/n600 ), .Z(\SUBBYTES[0].a/n598 ) );
  XOR \SUBBYTES[0].a/U5318  ( .A(\SUBBYTES[0].a/w1735 ), .B(
        \SUBBYTES[0].a/w1737 ), .Z(\SUBBYTES[0].a/n599 ) );
  XOR \SUBBYTES[0].a/U5317  ( .A(\SUBBYTES[0].a/w1695 ), .B(
        \SUBBYTES[0].a/w1727 ), .Z(\SUBBYTES[0].a/n600 ) );
  XOR \SUBBYTES[0].a/U5316  ( .A(\SUBBYTES[0].a/w1527 ), .B(
        \SUBBYTES[0].a/w1528 ), .Z(\SUBBYTES[0].a/n1471 ) );
  XOR \SUBBYTES[0].a/U5315  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n601 ), .Z(\SUBBYTES[0].a/n1470 ) );
  XOR \SUBBYTES[0].a/U5314  ( .A(\SUBBYTES[0].a/w1520 ), .B(
        \SUBBYTES[0].a/w1537 ), .Z(\SUBBYTES[0].a/n601 ) );
  XOR \SUBBYTES[0].a/U5313  ( .A(\SUBBYTES[0].a/n1470 ), .B(
        \SUBBYTES[0].a/n602 ), .Z(\SUBBYTES[0].a/n1689 ) );
  XOR \SUBBYTES[0].a/U5312  ( .A(\SUBBYTES[0].a/w1519 ), .B(
        \SUBBYTES[0].a/w1534 ), .Z(\SUBBYTES[0].a/n602 ) );
  XOR \SUBBYTES[0].a/U5311  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n603 ), .Z(\SUBBYTES[0].a/n1691 ) );
  XOR \SUBBYTES[0].a/U5310  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n603 ) );
  XOR \SUBBYTES[0].a/U5309  ( .A(\SUBBYTES[0].a/w1496 ), .B(
        \SUBBYTES[0].a/n604 ), .Z(\SUBBYTES[0].a/n1473 ) );
  XOR \SUBBYTES[0].a/U5308  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1488 ), .Z(\SUBBYTES[0].a/n604 ) );
  XOR \SUBBYTES[0].a/U5307  ( .A(\SUBBYTES[0].a/n1473 ), .B(
        \SUBBYTES[0].a/n605 ), .Z(\SUBBYTES[0].a/n1690 ) );
  XOR \SUBBYTES[0].a/U5306  ( .A(\SUBBYTES[0].a/w1498 ), .B(
        \SUBBYTES[0].a/n1691 ), .Z(\SUBBYTES[0].a/n605 ) );
  XOR \SUBBYTES[0].a/U5305  ( .A(\SUBBYTES[0].a/n607 ), .B(
        \SUBBYTES[0].a/n606 ), .Z(\SUBBYTES[0].a/n1474 ) );
  XOR \SUBBYTES[0].a/U5304  ( .A(\SUBBYTES[0].a/n609 ), .B(
        \SUBBYTES[0].a/n608 ), .Z(\SUBBYTES[0].a/n606 ) );
  XOR \SUBBYTES[0].a/U5303  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n607 ) );
  XOR \SUBBYTES[0].a/U5302  ( .A(\SUBBYTES[0].a/w1498 ), .B(
        \SUBBYTES[0].a/w1522 ), .Z(\SUBBYTES[0].a/n608 ) );
  XOR \SUBBYTES[0].a/U5301  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1496 ), .Z(\SUBBYTES[0].a/n609 ) );
  XOR \SUBBYTES[0].a/U5300  ( .A(\SUBBYTES[0].a/w1519 ), .B(
        \SUBBYTES[0].a/n610 ), .Z(\SUBBYTES[0].a/n1472 ) );
  XOR \SUBBYTES[0].a/U5299  ( .A(\SUBBYTES[0].a/w1502 ), .B(
        \SUBBYTES[0].a/w1505 ), .Z(\SUBBYTES[0].a/n610 ) );
  XOR \SUBBYTES[0].a/U5298  ( .A(\SUBBYTES[0].a/n1472 ), .B(
        \SUBBYTES[0].a/n611 ), .Z(\SUBBYTES[0].a/n1692 ) );
  XOR \SUBBYTES[0].a/U5297  ( .A(\SUBBYTES[0].a/w1490 ), .B(
        \SUBBYTES[0].a/n1474 ), .Z(\SUBBYTES[0].a/n611 ) );
  XOR \SUBBYTES[0].a/U5296  ( .A(\SUBBYTES[0].a/n1470 ), .B(
        \SUBBYTES[0].a/n612 ), .Z(\SUBBYTES[0].a/n1693 ) );
  XOR \SUBBYTES[0].a/U5295  ( .A(\SUBBYTES[0].a/w1522 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n612 ) );
  XOR \SUBBYTES[0].a/U5294  ( .A(\SUBBYTES[0].a/n614 ), .B(
        \SUBBYTES[0].a/n613 ), .Z(\SUBBYTES[0].a/n1694 ) );
  XOR \SUBBYTES[0].a/U5293  ( .A(\SUBBYTES[0].a/n616 ), .B(
        \SUBBYTES[0].a/n615 ), .Z(\SUBBYTES[0].a/n613 ) );
  XOR \SUBBYTES[0].a/U5292  ( .A(\SUBBYTES[0].a/n618 ), .B(
        \SUBBYTES[0].a/n617 ), .Z(\SUBBYTES[0].a/n614 ) );
  XOR \SUBBYTES[0].a/U5291  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1537 ), .Z(\SUBBYTES[0].a/n615 ) );
  XOR \SUBBYTES[0].a/U5290  ( .A(\SUBBYTES[0].a/w1527 ), .B(
        \SUBBYTES[0].a/w1530 ), .Z(\SUBBYTES[0].a/n616 ) );
  XOR \SUBBYTES[0].a/U5289  ( .A(\SUBBYTES[0].a/w1502 ), .B(
        \SUBBYTES[0].a/w1503 ), .Z(\SUBBYTES[0].a/n617 ) );
  XOR \SUBBYTES[0].a/U5288  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1490 ), .Z(\SUBBYTES[0].a/n618 ) );
  XOR \SUBBYTES[0].a/U5287  ( .A(\SUBBYTES[0].a/n620 ), .B(
        \SUBBYTES[0].a/n619 ), .Z(\SUBBYTES[0].a/n1695 ) );
  XOR \SUBBYTES[0].a/U5286  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n621 ), .Z(\SUBBYTES[0].a/n619 ) );
  XOR \SUBBYTES[0].a/U5285  ( .A(\SUBBYTES[0].a/n1473 ), .B(
        \SUBBYTES[0].a/n1472 ), .Z(\SUBBYTES[0].a/n620 ) );
  XOR \SUBBYTES[0].a/U5284  ( .A(\SUBBYTES[0].a/w1495 ), .B(
        \SUBBYTES[0].a/w1522 ), .Z(\SUBBYTES[0].a/n621 ) );
  XOR \SUBBYTES[0].a/U5283  ( .A(\SUBBYTES[0].a/n623 ), .B(
        \SUBBYTES[0].a/n622 ), .Z(\SUBBYTES[0].a/n1696 ) );
  XOR \SUBBYTES[0].a/U5282  ( .A(\SUBBYTES[0].a/n1474 ), .B(
        \SUBBYTES[0].a/n624 ), .Z(\SUBBYTES[0].a/n622 ) );
  XOR \SUBBYTES[0].a/U5281  ( .A(\SUBBYTES[0].a/w1528 ), .B(
        \SUBBYTES[0].a/w1530 ), .Z(\SUBBYTES[0].a/n623 ) );
  XOR \SUBBYTES[0].a/U5280  ( .A(\SUBBYTES[0].a/w1488 ), .B(
        \SUBBYTES[0].a/w1520 ), .Z(\SUBBYTES[0].a/n624 ) );
  XOR \SUBBYTES[0].a/U5279  ( .A(\SUBBYTES[0].a/w1320 ), .B(
        \SUBBYTES[0].a/w1321 ), .Z(\SUBBYTES[0].a/n1476 ) );
  XOR \SUBBYTES[0].a/U5278  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n625 ), .Z(\SUBBYTES[0].a/n1475 ) );
  XOR \SUBBYTES[0].a/U5277  ( .A(\SUBBYTES[0].a/w1313 ), .B(
        \SUBBYTES[0].a/w1330 ), .Z(\SUBBYTES[0].a/n625 ) );
  XOR \SUBBYTES[0].a/U5276  ( .A(\SUBBYTES[0].a/n1475 ), .B(
        \SUBBYTES[0].a/n626 ), .Z(\SUBBYTES[0].a/n1697 ) );
  XOR \SUBBYTES[0].a/U5275  ( .A(\SUBBYTES[0].a/w1312 ), .B(
        \SUBBYTES[0].a/w1327 ), .Z(\SUBBYTES[0].a/n626 ) );
  XOR \SUBBYTES[0].a/U5274  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n627 ), .Z(\SUBBYTES[0].a/n1699 ) );
  XOR \SUBBYTES[0].a/U5273  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n627 ) );
  XOR \SUBBYTES[0].a/U5272  ( .A(\SUBBYTES[0].a/w1289 ), .B(
        \SUBBYTES[0].a/n628 ), .Z(\SUBBYTES[0].a/n1478 ) );
  XOR \SUBBYTES[0].a/U5271  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1281 ), .Z(\SUBBYTES[0].a/n628 ) );
  XOR \SUBBYTES[0].a/U5270  ( .A(\SUBBYTES[0].a/n1478 ), .B(
        \SUBBYTES[0].a/n629 ), .Z(\SUBBYTES[0].a/n1698 ) );
  XOR \SUBBYTES[0].a/U5269  ( .A(\SUBBYTES[0].a/w1291 ), .B(
        \SUBBYTES[0].a/n1699 ), .Z(\SUBBYTES[0].a/n629 ) );
  XOR \SUBBYTES[0].a/U5268  ( .A(\SUBBYTES[0].a/n631 ), .B(
        \SUBBYTES[0].a/n630 ), .Z(\SUBBYTES[0].a/n1479 ) );
  XOR \SUBBYTES[0].a/U5267  ( .A(\SUBBYTES[0].a/n633 ), .B(
        \SUBBYTES[0].a/n632 ), .Z(\SUBBYTES[0].a/n630 ) );
  XOR \SUBBYTES[0].a/U5266  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n631 ) );
  XOR \SUBBYTES[0].a/U5265  ( .A(\SUBBYTES[0].a/w1291 ), .B(
        \SUBBYTES[0].a/w1315 ), .Z(\SUBBYTES[0].a/n632 ) );
  XOR \SUBBYTES[0].a/U5264  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1289 ), .Z(\SUBBYTES[0].a/n633 ) );
  XOR \SUBBYTES[0].a/U5263  ( .A(\SUBBYTES[0].a/w1312 ), .B(
        \SUBBYTES[0].a/n634 ), .Z(\SUBBYTES[0].a/n1477 ) );
  XOR \SUBBYTES[0].a/U5262  ( .A(\SUBBYTES[0].a/w1295 ), .B(
        \SUBBYTES[0].a/w1298 ), .Z(\SUBBYTES[0].a/n634 ) );
  XOR \SUBBYTES[0].a/U5261  ( .A(\SUBBYTES[0].a/n1477 ), .B(
        \SUBBYTES[0].a/n635 ), .Z(\SUBBYTES[0].a/n1700 ) );
  XOR \SUBBYTES[0].a/U5260  ( .A(\SUBBYTES[0].a/w1283 ), .B(
        \SUBBYTES[0].a/n1479 ), .Z(\SUBBYTES[0].a/n635 ) );
  XOR \SUBBYTES[0].a/U5259  ( .A(\SUBBYTES[0].a/n1475 ), .B(
        \SUBBYTES[0].a/n636 ), .Z(\SUBBYTES[0].a/n1701 ) );
  XOR \SUBBYTES[0].a/U5258  ( .A(\SUBBYTES[0].a/w1315 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n636 ) );
  XOR \SUBBYTES[0].a/U5257  ( .A(\SUBBYTES[0].a/n638 ), .B(
        \SUBBYTES[0].a/n637 ), .Z(\SUBBYTES[0].a/n1702 ) );
  XOR \SUBBYTES[0].a/U5256  ( .A(\SUBBYTES[0].a/n640 ), .B(
        \SUBBYTES[0].a/n639 ), .Z(\SUBBYTES[0].a/n637 ) );
  XOR \SUBBYTES[0].a/U5255  ( .A(\SUBBYTES[0].a/n642 ), .B(
        \SUBBYTES[0].a/n641 ), .Z(\SUBBYTES[0].a/n638 ) );
  XOR \SUBBYTES[0].a/U5254  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1330 ), .Z(\SUBBYTES[0].a/n639 ) );
  XOR \SUBBYTES[0].a/U5253  ( .A(\SUBBYTES[0].a/w1320 ), .B(
        \SUBBYTES[0].a/w1323 ), .Z(\SUBBYTES[0].a/n640 ) );
  XOR \SUBBYTES[0].a/U5252  ( .A(\SUBBYTES[0].a/w1295 ), .B(
        \SUBBYTES[0].a/w1296 ), .Z(\SUBBYTES[0].a/n641 ) );
  XOR \SUBBYTES[0].a/U5251  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1283 ), .Z(\SUBBYTES[0].a/n642 ) );
  XOR \SUBBYTES[0].a/U5250  ( .A(\SUBBYTES[0].a/n644 ), .B(
        \SUBBYTES[0].a/n643 ), .Z(\SUBBYTES[0].a/n1703 ) );
  XOR \SUBBYTES[0].a/U5249  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n645 ), .Z(\SUBBYTES[0].a/n643 ) );
  XOR \SUBBYTES[0].a/U5248  ( .A(\SUBBYTES[0].a/n1478 ), .B(
        \SUBBYTES[0].a/n1477 ), .Z(\SUBBYTES[0].a/n644 ) );
  XOR \SUBBYTES[0].a/U5247  ( .A(\SUBBYTES[0].a/w1288 ), .B(
        \SUBBYTES[0].a/w1315 ), .Z(\SUBBYTES[0].a/n645 ) );
  XOR \SUBBYTES[0].a/U5246  ( .A(\SUBBYTES[0].a/n647 ), .B(
        \SUBBYTES[0].a/n646 ), .Z(\SUBBYTES[0].a/n1704 ) );
  XOR \SUBBYTES[0].a/U5245  ( .A(\SUBBYTES[0].a/n1479 ), .B(
        \SUBBYTES[0].a/n648 ), .Z(\SUBBYTES[0].a/n646 ) );
  XOR \SUBBYTES[0].a/U5244  ( .A(\SUBBYTES[0].a/w1321 ), .B(
        \SUBBYTES[0].a/w1323 ), .Z(\SUBBYTES[0].a/n647 ) );
  XOR \SUBBYTES[0].a/U5243  ( .A(\SUBBYTES[0].a/w1281 ), .B(
        \SUBBYTES[0].a/w1313 ), .Z(\SUBBYTES[0].a/n648 ) );
  XOR \SUBBYTES[0].a/U5242  ( .A(\SUBBYTES[0].a/w1113 ), .B(
        \SUBBYTES[0].a/w1114 ), .Z(\SUBBYTES[0].a/n1481 ) );
  XOR \SUBBYTES[0].a/U5241  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n649 ), .Z(\SUBBYTES[0].a/n1480 ) );
  XOR \SUBBYTES[0].a/U5240  ( .A(\SUBBYTES[0].a/w1106 ), .B(
        \SUBBYTES[0].a/w1123 ), .Z(\SUBBYTES[0].a/n649 ) );
  XOR \SUBBYTES[0].a/U5239  ( .A(\SUBBYTES[0].a/n1480 ), .B(
        \SUBBYTES[0].a/n650 ), .Z(\SUBBYTES[0].a/n1705 ) );
  XOR \SUBBYTES[0].a/U5238  ( .A(\SUBBYTES[0].a/w1105 ), .B(
        \SUBBYTES[0].a/w1120 ), .Z(\SUBBYTES[0].a/n650 ) );
  XOR \SUBBYTES[0].a/U5237  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n651 ), .Z(\SUBBYTES[0].a/n1707 ) );
  XOR \SUBBYTES[0].a/U5236  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n651 ) );
  XOR \SUBBYTES[0].a/U5235  ( .A(\SUBBYTES[0].a/w1082 ), .B(
        \SUBBYTES[0].a/n652 ), .Z(\SUBBYTES[0].a/n1483 ) );
  XOR \SUBBYTES[0].a/U5234  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1074 ), .Z(\SUBBYTES[0].a/n652 ) );
  XOR \SUBBYTES[0].a/U5233  ( .A(\SUBBYTES[0].a/n1483 ), .B(
        \SUBBYTES[0].a/n653 ), .Z(\SUBBYTES[0].a/n1706 ) );
  XOR \SUBBYTES[0].a/U5232  ( .A(\SUBBYTES[0].a/w1084 ), .B(
        \SUBBYTES[0].a/n1707 ), .Z(\SUBBYTES[0].a/n653 ) );
  XOR \SUBBYTES[0].a/U5231  ( .A(\SUBBYTES[0].a/n655 ), .B(
        \SUBBYTES[0].a/n654 ), .Z(\SUBBYTES[0].a/n1484 ) );
  XOR \SUBBYTES[0].a/U5230  ( .A(\SUBBYTES[0].a/n657 ), .B(
        \SUBBYTES[0].a/n656 ), .Z(\SUBBYTES[0].a/n654 ) );
  XOR \SUBBYTES[0].a/U5229  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n655 ) );
  XOR \SUBBYTES[0].a/U5228  ( .A(\SUBBYTES[0].a/w1084 ), .B(
        \SUBBYTES[0].a/w1108 ), .Z(\SUBBYTES[0].a/n656 ) );
  XOR \SUBBYTES[0].a/U5227  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1082 ), .Z(\SUBBYTES[0].a/n657 ) );
  XOR \SUBBYTES[0].a/U5226  ( .A(\SUBBYTES[0].a/w1105 ), .B(
        \SUBBYTES[0].a/n658 ), .Z(\SUBBYTES[0].a/n1482 ) );
  XOR \SUBBYTES[0].a/U5225  ( .A(\SUBBYTES[0].a/w1088 ), .B(
        \SUBBYTES[0].a/w1091 ), .Z(\SUBBYTES[0].a/n658 ) );
  XOR \SUBBYTES[0].a/U5224  ( .A(\SUBBYTES[0].a/n1482 ), .B(
        \SUBBYTES[0].a/n659 ), .Z(\SUBBYTES[0].a/n1708 ) );
  XOR \SUBBYTES[0].a/U5223  ( .A(\SUBBYTES[0].a/w1076 ), .B(
        \SUBBYTES[0].a/n1484 ), .Z(\SUBBYTES[0].a/n659 ) );
  XOR \SUBBYTES[0].a/U5222  ( .A(\SUBBYTES[0].a/n1480 ), .B(
        \SUBBYTES[0].a/n660 ), .Z(\SUBBYTES[0].a/n1709 ) );
  XOR \SUBBYTES[0].a/U5221  ( .A(\SUBBYTES[0].a/w1108 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n660 ) );
  XOR \SUBBYTES[0].a/U5220  ( .A(\SUBBYTES[0].a/n662 ), .B(
        \SUBBYTES[0].a/n661 ), .Z(\SUBBYTES[0].a/n1710 ) );
  XOR \SUBBYTES[0].a/U5219  ( .A(\SUBBYTES[0].a/n664 ), .B(
        \SUBBYTES[0].a/n663 ), .Z(\SUBBYTES[0].a/n661 ) );
  XOR \SUBBYTES[0].a/U5218  ( .A(\SUBBYTES[0].a/n666 ), .B(
        \SUBBYTES[0].a/n665 ), .Z(\SUBBYTES[0].a/n662 ) );
  XOR \SUBBYTES[0].a/U5217  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1123 ), .Z(\SUBBYTES[0].a/n663 ) );
  XOR \SUBBYTES[0].a/U5216  ( .A(\SUBBYTES[0].a/w1113 ), .B(
        \SUBBYTES[0].a/w1116 ), .Z(\SUBBYTES[0].a/n664 ) );
  XOR \SUBBYTES[0].a/U5215  ( .A(\SUBBYTES[0].a/w1088 ), .B(
        \SUBBYTES[0].a/w1089 ), .Z(\SUBBYTES[0].a/n665 ) );
  XOR \SUBBYTES[0].a/U5214  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1076 ), .Z(\SUBBYTES[0].a/n666 ) );
  XOR \SUBBYTES[0].a/U5213  ( .A(\SUBBYTES[0].a/n668 ), .B(
        \SUBBYTES[0].a/n667 ), .Z(\SUBBYTES[0].a/n1711 ) );
  XOR \SUBBYTES[0].a/U5212  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n669 ), .Z(\SUBBYTES[0].a/n667 ) );
  XOR \SUBBYTES[0].a/U5211  ( .A(\SUBBYTES[0].a/n1483 ), .B(
        \SUBBYTES[0].a/n1482 ), .Z(\SUBBYTES[0].a/n668 ) );
  XOR \SUBBYTES[0].a/U5210  ( .A(\SUBBYTES[0].a/w1081 ), .B(
        \SUBBYTES[0].a/w1108 ), .Z(\SUBBYTES[0].a/n669 ) );
  XOR \SUBBYTES[0].a/U5209  ( .A(\SUBBYTES[0].a/n671 ), .B(
        \SUBBYTES[0].a/n670 ), .Z(\SUBBYTES[0].a/n1712 ) );
  XOR \SUBBYTES[0].a/U5208  ( .A(\SUBBYTES[0].a/n1484 ), .B(
        \SUBBYTES[0].a/n672 ), .Z(\SUBBYTES[0].a/n670 ) );
  XOR \SUBBYTES[0].a/U5207  ( .A(\SUBBYTES[0].a/w1114 ), .B(
        \SUBBYTES[0].a/w1116 ), .Z(\SUBBYTES[0].a/n671 ) );
  XOR \SUBBYTES[0].a/U5206  ( .A(\SUBBYTES[0].a/w1074 ), .B(
        \SUBBYTES[0].a/w1106 ), .Z(\SUBBYTES[0].a/n672 ) );
  XOR \SUBBYTES[0].a/U5205  ( .A(\SUBBYTES[0].a/w906 ), .B(
        \SUBBYTES[0].a/w907 ), .Z(\SUBBYTES[0].a/n1486 ) );
  XOR \SUBBYTES[0].a/U5204  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n673 ), .Z(\SUBBYTES[0].a/n1485 ) );
  XOR \SUBBYTES[0].a/U5203  ( .A(\SUBBYTES[0].a/w899 ), .B(
        \SUBBYTES[0].a/w916 ), .Z(\SUBBYTES[0].a/n673 ) );
  XOR \SUBBYTES[0].a/U5202  ( .A(\SUBBYTES[0].a/n1485 ), .B(
        \SUBBYTES[0].a/n674 ), .Z(\SUBBYTES[0].a/n1713 ) );
  XOR \SUBBYTES[0].a/U5201  ( .A(\SUBBYTES[0].a/w898 ), .B(
        \SUBBYTES[0].a/w913 ), .Z(\SUBBYTES[0].a/n674 ) );
  XOR \SUBBYTES[0].a/U5200  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n675 ), .Z(\SUBBYTES[0].a/n1715 ) );
  XOR \SUBBYTES[0].a/U5199  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n675 ) );
  XOR \SUBBYTES[0].a/U5198  ( .A(\SUBBYTES[0].a/w875 ), .B(
        \SUBBYTES[0].a/n676 ), .Z(\SUBBYTES[0].a/n1488 ) );
  XOR \SUBBYTES[0].a/U5197  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w867 ), .Z(\SUBBYTES[0].a/n676 ) );
  XOR \SUBBYTES[0].a/U5196  ( .A(\SUBBYTES[0].a/n1488 ), .B(
        \SUBBYTES[0].a/n677 ), .Z(\SUBBYTES[0].a/n1714 ) );
  XOR \SUBBYTES[0].a/U5195  ( .A(\SUBBYTES[0].a/w877 ), .B(
        \SUBBYTES[0].a/n1715 ), .Z(\SUBBYTES[0].a/n677 ) );
  XOR \SUBBYTES[0].a/U5194  ( .A(\SUBBYTES[0].a/n679 ), .B(
        \SUBBYTES[0].a/n678 ), .Z(\SUBBYTES[0].a/n1489 ) );
  XOR \SUBBYTES[0].a/U5193  ( .A(\SUBBYTES[0].a/n681 ), .B(
        \SUBBYTES[0].a/n680 ), .Z(\SUBBYTES[0].a/n678 ) );
  XOR \SUBBYTES[0].a/U5192  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n679 ) );
  XOR \SUBBYTES[0].a/U5191  ( .A(\SUBBYTES[0].a/w877 ), .B(
        \SUBBYTES[0].a/w901 ), .Z(\SUBBYTES[0].a/n680 ) );
  XOR \SUBBYTES[0].a/U5190  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w875 ), .Z(\SUBBYTES[0].a/n681 ) );
  XOR \SUBBYTES[0].a/U5189  ( .A(\SUBBYTES[0].a/w898 ), .B(
        \SUBBYTES[0].a/n682 ), .Z(\SUBBYTES[0].a/n1487 ) );
  XOR \SUBBYTES[0].a/U5188  ( .A(\SUBBYTES[0].a/w881 ), .B(
        \SUBBYTES[0].a/w884 ), .Z(\SUBBYTES[0].a/n682 ) );
  XOR \SUBBYTES[0].a/U5187  ( .A(\SUBBYTES[0].a/n1487 ), .B(
        \SUBBYTES[0].a/n683 ), .Z(\SUBBYTES[0].a/n1716 ) );
  XOR \SUBBYTES[0].a/U5186  ( .A(\SUBBYTES[0].a/w869 ), .B(
        \SUBBYTES[0].a/n1489 ), .Z(\SUBBYTES[0].a/n683 ) );
  XOR \SUBBYTES[0].a/U5185  ( .A(\SUBBYTES[0].a/n1485 ), .B(
        \SUBBYTES[0].a/n684 ), .Z(\SUBBYTES[0].a/n1717 ) );
  XOR \SUBBYTES[0].a/U5184  ( .A(\SUBBYTES[0].a/w901 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n684 ) );
  XOR \SUBBYTES[0].a/U5183  ( .A(\SUBBYTES[0].a/n686 ), .B(
        \SUBBYTES[0].a/n685 ), .Z(\SUBBYTES[0].a/n1718 ) );
  XOR \SUBBYTES[0].a/U5182  ( .A(\SUBBYTES[0].a/n688 ), .B(
        \SUBBYTES[0].a/n687 ), .Z(\SUBBYTES[0].a/n685 ) );
  XOR \SUBBYTES[0].a/U5181  ( .A(\SUBBYTES[0].a/n690 ), .B(
        \SUBBYTES[0].a/n689 ), .Z(\SUBBYTES[0].a/n686 ) );
  XOR \SUBBYTES[0].a/U5180  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w916 ), .Z(\SUBBYTES[0].a/n687 ) );
  XOR \SUBBYTES[0].a/U5179  ( .A(\SUBBYTES[0].a/w906 ), .B(
        \SUBBYTES[0].a/w909 ), .Z(\SUBBYTES[0].a/n688 ) );
  XOR \SUBBYTES[0].a/U5178  ( .A(\SUBBYTES[0].a/w881 ), .B(
        \SUBBYTES[0].a/w882 ), .Z(\SUBBYTES[0].a/n689 ) );
  XOR \SUBBYTES[0].a/U5177  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w869 ), .Z(\SUBBYTES[0].a/n690 ) );
  XOR \SUBBYTES[0].a/U5176  ( .A(\SUBBYTES[0].a/n692 ), .B(
        \SUBBYTES[0].a/n691 ), .Z(\SUBBYTES[0].a/n1719 ) );
  XOR \SUBBYTES[0].a/U5175  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n693 ), .Z(\SUBBYTES[0].a/n691 ) );
  XOR \SUBBYTES[0].a/U5174  ( .A(\SUBBYTES[0].a/n1488 ), .B(
        \SUBBYTES[0].a/n1487 ), .Z(\SUBBYTES[0].a/n692 ) );
  XOR \SUBBYTES[0].a/U5173  ( .A(\SUBBYTES[0].a/w874 ), .B(
        \SUBBYTES[0].a/w901 ), .Z(\SUBBYTES[0].a/n693 ) );
  XOR \SUBBYTES[0].a/U5172  ( .A(\SUBBYTES[0].a/n695 ), .B(
        \SUBBYTES[0].a/n694 ), .Z(\SUBBYTES[0].a/n1720 ) );
  XOR \SUBBYTES[0].a/U5171  ( .A(\SUBBYTES[0].a/n1489 ), .B(
        \SUBBYTES[0].a/n696 ), .Z(\SUBBYTES[0].a/n694 ) );
  XOR \SUBBYTES[0].a/U5170  ( .A(\SUBBYTES[0].a/w907 ), .B(
        \SUBBYTES[0].a/w909 ), .Z(\SUBBYTES[0].a/n695 ) );
  XOR \SUBBYTES[0].a/U5169  ( .A(\SUBBYTES[0].a/w867 ), .B(
        \SUBBYTES[0].a/w899 ), .Z(\SUBBYTES[0].a/n696 ) );
  XOR \SUBBYTES[0].a/U5168  ( .A(\SUBBYTES[0].a/w699 ), .B(
        \SUBBYTES[0].a/w700 ), .Z(\SUBBYTES[0].a/n1491 ) );
  XOR \SUBBYTES[0].a/U5167  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n697 ), .Z(\SUBBYTES[0].a/n1490 ) );
  XOR \SUBBYTES[0].a/U5166  ( .A(\SUBBYTES[0].a/w692 ), .B(
        \SUBBYTES[0].a/w709 ), .Z(\SUBBYTES[0].a/n697 ) );
  XOR \SUBBYTES[0].a/U5165  ( .A(\SUBBYTES[0].a/n1490 ), .B(
        \SUBBYTES[0].a/n698 ), .Z(\SUBBYTES[0].a/n1721 ) );
  XOR \SUBBYTES[0].a/U5164  ( .A(\SUBBYTES[0].a/w691 ), .B(
        \SUBBYTES[0].a/w706 ), .Z(\SUBBYTES[0].a/n698 ) );
  XOR \SUBBYTES[0].a/U5163  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n699 ), .Z(\SUBBYTES[0].a/n1723 ) );
  XOR \SUBBYTES[0].a/U5162  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n699 ) );
  XOR \SUBBYTES[0].a/U5161  ( .A(\SUBBYTES[0].a/w668 ), .B(
        \SUBBYTES[0].a/n700 ), .Z(\SUBBYTES[0].a/n1493 ) );
  XOR \SUBBYTES[0].a/U5160  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w660 ), .Z(\SUBBYTES[0].a/n700 ) );
  XOR \SUBBYTES[0].a/U5159  ( .A(\SUBBYTES[0].a/n1493 ), .B(
        \SUBBYTES[0].a/n701 ), .Z(\SUBBYTES[0].a/n1722 ) );
  XOR \SUBBYTES[0].a/U5158  ( .A(\SUBBYTES[0].a/w670 ), .B(
        \SUBBYTES[0].a/n1723 ), .Z(\SUBBYTES[0].a/n701 ) );
  XOR \SUBBYTES[0].a/U5157  ( .A(\SUBBYTES[0].a/n703 ), .B(
        \SUBBYTES[0].a/n702 ), .Z(\SUBBYTES[0].a/n1494 ) );
  XOR \SUBBYTES[0].a/U5156  ( .A(\SUBBYTES[0].a/n705 ), .B(
        \SUBBYTES[0].a/n704 ), .Z(\SUBBYTES[0].a/n702 ) );
  XOR \SUBBYTES[0].a/U5155  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n703 ) );
  XOR \SUBBYTES[0].a/U5154  ( .A(\SUBBYTES[0].a/w670 ), .B(
        \SUBBYTES[0].a/w694 ), .Z(\SUBBYTES[0].a/n704 ) );
  XOR \SUBBYTES[0].a/U5153  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w668 ), .Z(\SUBBYTES[0].a/n705 ) );
  XOR \SUBBYTES[0].a/U5152  ( .A(\SUBBYTES[0].a/w691 ), .B(
        \SUBBYTES[0].a/n706 ), .Z(\SUBBYTES[0].a/n1492 ) );
  XOR \SUBBYTES[0].a/U5151  ( .A(\SUBBYTES[0].a/w674 ), .B(
        \SUBBYTES[0].a/w677 ), .Z(\SUBBYTES[0].a/n706 ) );
  XOR \SUBBYTES[0].a/U5150  ( .A(\SUBBYTES[0].a/n1492 ), .B(
        \SUBBYTES[0].a/n707 ), .Z(\SUBBYTES[0].a/n1724 ) );
  XOR \SUBBYTES[0].a/U5149  ( .A(\SUBBYTES[0].a/w662 ), .B(
        \SUBBYTES[0].a/n1494 ), .Z(\SUBBYTES[0].a/n707 ) );
  XOR \SUBBYTES[0].a/U5148  ( .A(\SUBBYTES[0].a/n1490 ), .B(
        \SUBBYTES[0].a/n708 ), .Z(\SUBBYTES[0].a/n1725 ) );
  XOR \SUBBYTES[0].a/U5147  ( .A(\SUBBYTES[0].a/w694 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n708 ) );
  XOR \SUBBYTES[0].a/U5146  ( .A(\SUBBYTES[0].a/n710 ), .B(
        \SUBBYTES[0].a/n709 ), .Z(\SUBBYTES[0].a/n1726 ) );
  XOR \SUBBYTES[0].a/U5145  ( .A(\SUBBYTES[0].a/n712 ), .B(
        \SUBBYTES[0].a/n711 ), .Z(\SUBBYTES[0].a/n709 ) );
  XOR \SUBBYTES[0].a/U5144  ( .A(\SUBBYTES[0].a/n714 ), .B(
        \SUBBYTES[0].a/n713 ), .Z(\SUBBYTES[0].a/n710 ) );
  XOR \SUBBYTES[0].a/U5143  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w709 ), .Z(\SUBBYTES[0].a/n711 ) );
  XOR \SUBBYTES[0].a/U5142  ( .A(\SUBBYTES[0].a/w699 ), .B(
        \SUBBYTES[0].a/w702 ), .Z(\SUBBYTES[0].a/n712 ) );
  XOR \SUBBYTES[0].a/U5141  ( .A(\SUBBYTES[0].a/w674 ), .B(
        \SUBBYTES[0].a/w675 ), .Z(\SUBBYTES[0].a/n713 ) );
  XOR \SUBBYTES[0].a/U5140  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w662 ), .Z(\SUBBYTES[0].a/n714 ) );
  XOR \SUBBYTES[0].a/U5139  ( .A(\SUBBYTES[0].a/n716 ), .B(
        \SUBBYTES[0].a/n715 ), .Z(\SUBBYTES[0].a/n1727 ) );
  XOR \SUBBYTES[0].a/U5138  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n717 ), .Z(\SUBBYTES[0].a/n715 ) );
  XOR \SUBBYTES[0].a/U5137  ( .A(\SUBBYTES[0].a/n1493 ), .B(
        \SUBBYTES[0].a/n1492 ), .Z(\SUBBYTES[0].a/n716 ) );
  XOR \SUBBYTES[0].a/U5136  ( .A(\SUBBYTES[0].a/w667 ), .B(
        \SUBBYTES[0].a/w694 ), .Z(\SUBBYTES[0].a/n717 ) );
  XOR \SUBBYTES[0].a/U5135  ( .A(\SUBBYTES[0].a/n719 ), .B(
        \SUBBYTES[0].a/n718 ), .Z(\SUBBYTES[0].a/n1728 ) );
  XOR \SUBBYTES[0].a/U5134  ( .A(\SUBBYTES[0].a/n1494 ), .B(
        \SUBBYTES[0].a/n720 ), .Z(\SUBBYTES[0].a/n718 ) );
  XOR \SUBBYTES[0].a/U5133  ( .A(\SUBBYTES[0].a/w700 ), .B(
        \SUBBYTES[0].a/w702 ), .Z(\SUBBYTES[0].a/n719 ) );
  XOR \SUBBYTES[0].a/U5132  ( .A(\SUBBYTES[0].a/w660 ), .B(
        \SUBBYTES[0].a/w692 ), .Z(\SUBBYTES[0].a/n720 ) );
  XOR \SUBBYTES[0].a/U5131  ( .A(\SUBBYTES[0].a/w492 ), .B(
        \SUBBYTES[0].a/w493 ), .Z(\SUBBYTES[0].a/n1496 ) );
  XOR \SUBBYTES[0].a/U5130  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n721 ), .Z(\SUBBYTES[0].a/n1495 ) );
  XOR \SUBBYTES[0].a/U5129  ( .A(\SUBBYTES[0].a/w485 ), .B(
        \SUBBYTES[0].a/w502 ), .Z(\SUBBYTES[0].a/n721 ) );
  XOR \SUBBYTES[0].a/U5128  ( .A(\SUBBYTES[0].a/n1495 ), .B(
        \SUBBYTES[0].a/n722 ), .Z(\SUBBYTES[0].a/n1729 ) );
  XOR \SUBBYTES[0].a/U5127  ( .A(\SUBBYTES[0].a/w484 ), .B(
        \SUBBYTES[0].a/w499 ), .Z(\SUBBYTES[0].a/n722 ) );
  XOR \SUBBYTES[0].a/U5126  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n723 ), .Z(\SUBBYTES[0].a/n1731 ) );
  XOR \SUBBYTES[0].a/U5125  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n723 ) );
  XOR \SUBBYTES[0].a/U5124  ( .A(\SUBBYTES[0].a/w461 ), .B(
        \SUBBYTES[0].a/n724 ), .Z(\SUBBYTES[0].a/n1498 ) );
  XOR \SUBBYTES[0].a/U5123  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w453 ), .Z(\SUBBYTES[0].a/n724 ) );
  XOR \SUBBYTES[0].a/U5122  ( .A(\SUBBYTES[0].a/n1498 ), .B(
        \SUBBYTES[0].a/n725 ), .Z(\SUBBYTES[0].a/n1730 ) );
  XOR \SUBBYTES[0].a/U5121  ( .A(\SUBBYTES[0].a/w463 ), .B(
        \SUBBYTES[0].a/n1731 ), .Z(\SUBBYTES[0].a/n725 ) );
  XOR \SUBBYTES[0].a/U5120  ( .A(\SUBBYTES[0].a/n727 ), .B(
        \SUBBYTES[0].a/n726 ), .Z(\SUBBYTES[0].a/n1499 ) );
  XOR \SUBBYTES[0].a/U5119  ( .A(\SUBBYTES[0].a/n729 ), .B(
        \SUBBYTES[0].a/n728 ), .Z(\SUBBYTES[0].a/n726 ) );
  XOR \SUBBYTES[0].a/U5118  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n727 ) );
  XOR \SUBBYTES[0].a/U5117  ( .A(\SUBBYTES[0].a/w463 ), .B(
        \SUBBYTES[0].a/w487 ), .Z(\SUBBYTES[0].a/n728 ) );
  XOR \SUBBYTES[0].a/U5116  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w461 ), .Z(\SUBBYTES[0].a/n729 ) );
  XOR \SUBBYTES[0].a/U5115  ( .A(\SUBBYTES[0].a/w484 ), .B(
        \SUBBYTES[0].a/n730 ), .Z(\SUBBYTES[0].a/n1497 ) );
  XOR \SUBBYTES[0].a/U5114  ( .A(\SUBBYTES[0].a/w467 ), .B(
        \SUBBYTES[0].a/w470 ), .Z(\SUBBYTES[0].a/n730 ) );
  XOR \SUBBYTES[0].a/U5113  ( .A(\SUBBYTES[0].a/n1497 ), .B(
        \SUBBYTES[0].a/n731 ), .Z(\SUBBYTES[0].a/n1732 ) );
  XOR \SUBBYTES[0].a/U5112  ( .A(\SUBBYTES[0].a/w455 ), .B(
        \SUBBYTES[0].a/n1499 ), .Z(\SUBBYTES[0].a/n731 ) );
  XOR \SUBBYTES[0].a/U5111  ( .A(\SUBBYTES[0].a/n1495 ), .B(
        \SUBBYTES[0].a/n732 ), .Z(\SUBBYTES[0].a/n1733 ) );
  XOR \SUBBYTES[0].a/U5110  ( .A(\SUBBYTES[0].a/w487 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n732 ) );
  XOR \SUBBYTES[0].a/U5109  ( .A(\SUBBYTES[0].a/n734 ), .B(
        \SUBBYTES[0].a/n733 ), .Z(\SUBBYTES[0].a/n1734 ) );
  XOR \SUBBYTES[0].a/U5108  ( .A(\SUBBYTES[0].a/n736 ), .B(
        \SUBBYTES[0].a/n735 ), .Z(\SUBBYTES[0].a/n733 ) );
  XOR \SUBBYTES[0].a/U5107  ( .A(\SUBBYTES[0].a/n738 ), .B(
        \SUBBYTES[0].a/n737 ), .Z(\SUBBYTES[0].a/n734 ) );
  XOR \SUBBYTES[0].a/U5106  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w502 ), .Z(\SUBBYTES[0].a/n735 ) );
  XOR \SUBBYTES[0].a/U5105  ( .A(\SUBBYTES[0].a/w492 ), .B(
        \SUBBYTES[0].a/w495 ), .Z(\SUBBYTES[0].a/n736 ) );
  XOR \SUBBYTES[0].a/U5104  ( .A(\SUBBYTES[0].a/w467 ), .B(
        \SUBBYTES[0].a/w468 ), .Z(\SUBBYTES[0].a/n737 ) );
  XOR \SUBBYTES[0].a/U5103  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w455 ), .Z(\SUBBYTES[0].a/n738 ) );
  XOR \SUBBYTES[0].a/U5102  ( .A(\SUBBYTES[0].a/n740 ), .B(
        \SUBBYTES[0].a/n739 ), .Z(\SUBBYTES[0].a/n1735 ) );
  XOR \SUBBYTES[0].a/U5101  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n741 ), .Z(\SUBBYTES[0].a/n739 ) );
  XOR \SUBBYTES[0].a/U5100  ( .A(\SUBBYTES[0].a/n1498 ), .B(
        \SUBBYTES[0].a/n1497 ), .Z(\SUBBYTES[0].a/n740 ) );
  XOR \SUBBYTES[0].a/U5099  ( .A(\SUBBYTES[0].a/w460 ), .B(
        \SUBBYTES[0].a/w487 ), .Z(\SUBBYTES[0].a/n741 ) );
  XOR \SUBBYTES[0].a/U5098  ( .A(\SUBBYTES[0].a/n743 ), .B(
        \SUBBYTES[0].a/n742 ), .Z(\SUBBYTES[0].a/n1736 ) );
  XOR \SUBBYTES[0].a/U5097  ( .A(\SUBBYTES[0].a/n1499 ), .B(
        \SUBBYTES[0].a/n744 ), .Z(\SUBBYTES[0].a/n742 ) );
  XOR \SUBBYTES[0].a/U5096  ( .A(\SUBBYTES[0].a/w493 ), .B(
        \SUBBYTES[0].a/w495 ), .Z(\SUBBYTES[0].a/n743 ) );
  XOR \SUBBYTES[0].a/U5095  ( .A(\SUBBYTES[0].a/w453 ), .B(
        \SUBBYTES[0].a/w485 ), .Z(\SUBBYTES[0].a/n744 ) );
  XOR \SUBBYTES[0].a/U5094  ( .A(\SUBBYTES[0].a/w285 ), .B(
        \SUBBYTES[0].a/w286 ), .Z(\SUBBYTES[0].a/n1501 ) );
  XOR \SUBBYTES[0].a/U5093  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n745 ), .Z(\SUBBYTES[0].a/n1500 ) );
  XOR \SUBBYTES[0].a/U5092  ( .A(\SUBBYTES[0].a/w278 ), .B(
        \SUBBYTES[0].a/w295 ), .Z(\SUBBYTES[0].a/n745 ) );
  XOR \SUBBYTES[0].a/U5091  ( .A(\SUBBYTES[0].a/n1500 ), .B(
        \SUBBYTES[0].a/n746 ), .Z(\SUBBYTES[0].a/n1737 ) );
  XOR \SUBBYTES[0].a/U5090  ( .A(\SUBBYTES[0].a/w277 ), .B(
        \SUBBYTES[0].a/w292 ), .Z(\SUBBYTES[0].a/n746 ) );
  XOR \SUBBYTES[0].a/U5089  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n747 ), .Z(\SUBBYTES[0].a/n1739 ) );
  XOR \SUBBYTES[0].a/U5088  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n747 ) );
  XOR \SUBBYTES[0].a/U5087  ( .A(\SUBBYTES[0].a/w254 ), .B(
        \SUBBYTES[0].a/n748 ), .Z(\SUBBYTES[0].a/n1503 ) );
  XOR \SUBBYTES[0].a/U5086  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w246 ), .Z(\SUBBYTES[0].a/n748 ) );
  XOR \SUBBYTES[0].a/U5085  ( .A(\SUBBYTES[0].a/n1503 ), .B(
        \SUBBYTES[0].a/n749 ), .Z(\SUBBYTES[0].a/n1738 ) );
  XOR \SUBBYTES[0].a/U5084  ( .A(\SUBBYTES[0].a/w256 ), .B(
        \SUBBYTES[0].a/n1739 ), .Z(\SUBBYTES[0].a/n749 ) );
  XOR \SUBBYTES[0].a/U5083  ( .A(\SUBBYTES[0].a/n751 ), .B(
        \SUBBYTES[0].a/n750 ), .Z(\SUBBYTES[0].a/n1504 ) );
  XOR \SUBBYTES[0].a/U5082  ( .A(\SUBBYTES[0].a/n753 ), .B(
        \SUBBYTES[0].a/n752 ), .Z(\SUBBYTES[0].a/n750 ) );
  XOR \SUBBYTES[0].a/U5081  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n751 ) );
  XOR \SUBBYTES[0].a/U5080  ( .A(\SUBBYTES[0].a/w256 ), .B(
        \SUBBYTES[0].a/w280 ), .Z(\SUBBYTES[0].a/n752 ) );
  XOR \SUBBYTES[0].a/U5079  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w254 ), .Z(\SUBBYTES[0].a/n753 ) );
  XOR \SUBBYTES[0].a/U5078  ( .A(\SUBBYTES[0].a/w277 ), .B(
        \SUBBYTES[0].a/n754 ), .Z(\SUBBYTES[0].a/n1502 ) );
  XOR \SUBBYTES[0].a/U5077  ( .A(\SUBBYTES[0].a/w260 ), .B(
        \SUBBYTES[0].a/w263 ), .Z(\SUBBYTES[0].a/n754 ) );
  XOR \SUBBYTES[0].a/U5076  ( .A(\SUBBYTES[0].a/n1502 ), .B(
        \SUBBYTES[0].a/n755 ), .Z(\SUBBYTES[0].a/n1740 ) );
  XOR \SUBBYTES[0].a/U5075  ( .A(\SUBBYTES[0].a/w248 ), .B(
        \SUBBYTES[0].a/n1504 ), .Z(\SUBBYTES[0].a/n755 ) );
  XOR \SUBBYTES[0].a/U5074  ( .A(\SUBBYTES[0].a/n1500 ), .B(
        \SUBBYTES[0].a/n756 ), .Z(\SUBBYTES[0].a/n1741 ) );
  XOR \SUBBYTES[0].a/U5073  ( .A(\SUBBYTES[0].a/w280 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n756 ) );
  XOR \SUBBYTES[0].a/U5072  ( .A(\SUBBYTES[0].a/n758 ), .B(
        \SUBBYTES[0].a/n757 ), .Z(\SUBBYTES[0].a/n1742 ) );
  XOR \SUBBYTES[0].a/U5071  ( .A(\SUBBYTES[0].a/n760 ), .B(
        \SUBBYTES[0].a/n759 ), .Z(\SUBBYTES[0].a/n757 ) );
  XOR \SUBBYTES[0].a/U5070  ( .A(\SUBBYTES[0].a/n762 ), .B(
        \SUBBYTES[0].a/n761 ), .Z(\SUBBYTES[0].a/n758 ) );
  XOR \SUBBYTES[0].a/U5069  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w295 ), .Z(\SUBBYTES[0].a/n759 ) );
  XOR \SUBBYTES[0].a/U5068  ( .A(\SUBBYTES[0].a/w285 ), .B(
        \SUBBYTES[0].a/w288 ), .Z(\SUBBYTES[0].a/n760 ) );
  XOR \SUBBYTES[0].a/U5067  ( .A(\SUBBYTES[0].a/w260 ), .B(
        \SUBBYTES[0].a/w261 ), .Z(\SUBBYTES[0].a/n761 ) );
  XOR \SUBBYTES[0].a/U5066  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w248 ), .Z(\SUBBYTES[0].a/n762 ) );
  XOR \SUBBYTES[0].a/U5065  ( .A(\SUBBYTES[0].a/n764 ), .B(
        \SUBBYTES[0].a/n763 ), .Z(\SUBBYTES[0].a/n1743 ) );
  XOR \SUBBYTES[0].a/U5064  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n765 ), .Z(\SUBBYTES[0].a/n763 ) );
  XOR \SUBBYTES[0].a/U5063  ( .A(\SUBBYTES[0].a/n1503 ), .B(
        \SUBBYTES[0].a/n1502 ), .Z(\SUBBYTES[0].a/n764 ) );
  XOR \SUBBYTES[0].a/U5062  ( .A(\SUBBYTES[0].a/w253 ), .B(
        \SUBBYTES[0].a/w280 ), .Z(\SUBBYTES[0].a/n765 ) );
  XOR \SUBBYTES[0].a/U5061  ( .A(\SUBBYTES[0].a/n767 ), .B(
        \SUBBYTES[0].a/n766 ), .Z(\SUBBYTES[0].a/n1744 ) );
  XOR \SUBBYTES[0].a/U5060  ( .A(\SUBBYTES[0].a/n1504 ), .B(
        \SUBBYTES[0].a/n768 ), .Z(\SUBBYTES[0].a/n766 ) );
  XOR \SUBBYTES[0].a/U5059  ( .A(\SUBBYTES[0].a/w286 ), .B(
        \SUBBYTES[0].a/w288 ), .Z(\SUBBYTES[0].a/n767 ) );
  XOR \SUBBYTES[0].a/U5058  ( .A(\SUBBYTES[0].a/w246 ), .B(
        \SUBBYTES[0].a/w278 ), .Z(\SUBBYTES[0].a/n768 ) );
  XOR \SUBBYTES[0].a/U5057  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n769 ), .Z(
        \SUBBYTES[0].a/n1505 ) );
  XOR \SUBBYTES[0].a/U5056  ( .A(\w1[0][3] ), .B(\w1[0][2] ), .Z(
        \SUBBYTES[0].a/n769 ) );
  XOR \SUBBYTES[0].a/U5055  ( .A(\w1[0][6] ), .B(\SUBBYTES[0].a/n1505 ), .Z(
        \SUBBYTES[0].a/w3378 ) );
  XOR \SUBBYTES[0].a/U5054  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/w3265 ) );
  XOR \SUBBYTES[0].a/U5053  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/n770 ), .Z(
        \SUBBYTES[0].a/w3266 ) );
  XOR \SUBBYTES[0].a/U5052  ( .A(\w1[0][6] ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n770 ) );
  XOR \SUBBYTES[0].a/U5051  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n1505 ), .Z(
        \SUBBYTES[0].a/w3396 ) );
  XOR \SUBBYTES[0].a/U5050  ( .A(\SUBBYTES[0].a/n772 ), .B(
        \SUBBYTES[0].a/n771 ), .Z(\SUBBYTES[0].a/w3389 ) );
  XOR \SUBBYTES[0].a/U5049  ( .A(\w1[0][3] ), .B(\w1[0][1] ), .Z(
        \SUBBYTES[0].a/n771 ) );
  XOR \SUBBYTES[0].a/U5048  ( .A(\w1[0][7] ), .B(\w1[0][4] ), .Z(
        \SUBBYTES[0].a/n772 ) );
  XOR \SUBBYTES[0].a/U5047  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3389 ), .Z(
        \SUBBYTES[0].a/w3268 ) );
  XOR \SUBBYTES[0].a/U5046  ( .A(\SUBBYTES[0].a/n774 ), .B(
        \SUBBYTES[0].a/n773 ), .Z(\SUBBYTES[0].a/w3376 ) );
  XOR \SUBBYTES[0].a/U5045  ( .A(\SUBBYTES[0].a/w3337 ), .B(n16), .Z(
        \SUBBYTES[0].a/n773 ) );
  XOR \SUBBYTES[0].a/U5044  ( .A(\SUBBYTES[0].a/w3330 ), .B(
        \SUBBYTES[0].a/w3333 ), .Z(\SUBBYTES[0].a/n774 ) );
  XOR \SUBBYTES[0].a/U5043  ( .A(\SUBBYTES[0].a/n776 ), .B(
        \SUBBYTES[0].a/n775 ), .Z(\SUBBYTES[0].a/w3377 ) );
  XOR \SUBBYTES[0].a/U5042  ( .A(\SUBBYTES[0].a/w3337 ), .B(
        \SUBBYTES[0].a/n160 ), .Z(\SUBBYTES[0].a/n775 ) );
  XOR \SUBBYTES[0].a/U5041  ( .A(\SUBBYTES[0].a/w3330 ), .B(
        \SUBBYTES[0].a/n159 ), .Z(\SUBBYTES[0].a/n776 ) );
  XOR \SUBBYTES[0].a/U5040  ( .A(\SUBBYTES[0].a/w3389 ), .B(
        \SUBBYTES[0].a/n777 ), .Z(\SUBBYTES[0].a/w3379 ) );
  XOR \SUBBYTES[0].a/U5039  ( .A(\w1[0][6] ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n777 ) );
  XOR \SUBBYTES[0].a/U5038  ( .A(\SUBBYTES[0].a/n779 ), .B(
        \SUBBYTES[0].a/n778 ), .Z(\SUBBYTES[0].a/w3380 ) );
  XOR \SUBBYTES[0].a/U5037  ( .A(\SUBBYTES[0].a/n160 ), .B(n16), .Z(
        \SUBBYTES[0].a/n778 ) );
  XOR \SUBBYTES[0].a/U5036  ( .A(\SUBBYTES[0].a/n159 ), .B(
        \SUBBYTES[0].a/w3333 ), .Z(\SUBBYTES[0].a/n779 ) );
  XOR \SUBBYTES[0].a/U5035  ( .A(\w1[0][7] ), .B(\w1[0][2] ), .Z(
        \SUBBYTES[0].a/n1511 ) );
  XOR \SUBBYTES[0].a/U5034  ( .A(\SUBBYTES[0].a/n1511 ), .B(
        \SUBBYTES[0].a/n780 ), .Z(\SUBBYTES[0].a/w3381 ) );
  XOR \SUBBYTES[0].a/U5033  ( .A(\w1[0][5] ), .B(\w1[0][4] ), .Z(
        \SUBBYTES[0].a/n780 ) );
  XOR \SUBBYTES[0].a/U5032  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3269 ) );
  XOR \SUBBYTES[0].a/U5031  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3270 ) );
  XOR \SUBBYTES[0].a/U5030  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3271 ) );
  XOR \SUBBYTES[0].a/U5029  ( .A(\SUBBYTES[0].a/w3270 ), .B(
        \SUBBYTES[0].a/n1511 ), .Z(\SUBBYTES[0].a/w3272 ) );
  XOR \SUBBYTES[0].a/U5028  ( .A(\SUBBYTES[0].a/n1511 ), .B(
        \SUBBYTES[0].a/n781 ), .Z(\SUBBYTES[0].a/w3357 ) );
  XOR \SUBBYTES[0].a/U5027  ( .A(\w1[0][4] ), .B(\w1[0][1] ), .Z(
        \SUBBYTES[0].a/n781 ) );
  XOR \SUBBYTES[0].a/U5026  ( .A(\SUBBYTES[0].a/n783 ), .B(
        \SUBBYTES[0].a/n782 ), .Z(\SUBBYTES[0].a/n1508 ) );
  XOR \SUBBYTES[0].a/U5025  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/n784 ), .Z(
        \SUBBYTES[0].a/n782 ) );
  XOR \SUBBYTES[0].a/U5024  ( .A(\SUBBYTES[0].a/w3322 ), .B(\w1[0][6] ), .Z(
        \SUBBYTES[0].a/n783 ) );
  XOR \SUBBYTES[0].a/U5023  ( .A(\SUBBYTES[0].a/w3296 ), .B(
        \SUBBYTES[0].a/w3303 ), .Z(\SUBBYTES[0].a/n784 ) );
  XOR \SUBBYTES[0].a/U5022  ( .A(\SUBBYTES[0].a/n786 ), .B(
        \SUBBYTES[0].a/n785 ), .Z(\SUBBYTES[0].a/n1506 ) );
  XOR \SUBBYTES[0].a/U5021  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n787 ), .Z(
        \SUBBYTES[0].a/n785 ) );
  XOR \SUBBYTES[0].a/U5020  ( .A(\SUBBYTES[0].a/w3321 ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n786 ) );
  XOR \SUBBYTES[0].a/U5019  ( .A(\SUBBYTES[0].a/w3297 ), .B(
        \SUBBYTES[0].a/w3304 ), .Z(\SUBBYTES[0].a/n787 ) );
  XOR \SUBBYTES[0].a/U5018  ( .A(\SUBBYTES[0].a/n1508 ), .B(
        \SUBBYTES[0].a/n1506 ), .Z(\SUBBYTES[0].a/w3327 ) );
  XOR \SUBBYTES[0].a/U5017  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n788 ), .Z(
        \SUBBYTES[0].a/n1509 ) );
  XOR \SUBBYTES[0].a/U5016  ( .A(\SUBBYTES[0].a/w3289 ), .B(
        \SUBBYTES[0].a/w3299 ), .Z(\SUBBYTES[0].a/n788 ) );
  XOR \SUBBYTES[0].a/U5015  ( .A(\SUBBYTES[0].a/n790 ), .B(
        \SUBBYTES[0].a/n789 ), .Z(\SUBBYTES[0].a/w3314 ) );
  XOR \SUBBYTES[0].a/U5014  ( .A(\SUBBYTES[0].a/n1509 ), .B(
        \SUBBYTES[0].a/n791 ), .Z(\SUBBYTES[0].a/n789 ) );
  XOR \SUBBYTES[0].a/U5013  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/n790 ) );
  XOR \SUBBYTES[0].a/U5012  ( .A(\SUBBYTES[0].a/w3291 ), .B(
        \SUBBYTES[0].a/w3296 ), .Z(\SUBBYTES[0].a/n791 ) );
  XOR \SUBBYTES[0].a/U5011  ( .A(\SUBBYTES[0].a/n793 ), .B(
        \SUBBYTES[0].a/n792 ), .Z(\SUBBYTES[0].a/n1507 ) );
  XOR \SUBBYTES[0].a/U5010  ( .A(\SUBBYTES[0].a/w3324 ), .B(\w1[0][7] ), .Z(
        \SUBBYTES[0].a/n792 ) );
  XOR \SUBBYTES[0].a/U5009  ( .A(\SUBBYTES[0].a/w3299 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n793 ) );
  XOR \SUBBYTES[0].a/U5008  ( .A(\SUBBYTES[0].a/n1506 ), .B(
        \SUBBYTES[0].a/n1507 ), .Z(\SUBBYTES[0].a/w3326 ) );
  XOR \SUBBYTES[0].a/U5007  ( .A(\w1[0][3] ), .B(\SUBBYTES[0].a/n794 ), .Z(
        \SUBBYTES[0].a/n1510 ) );
  XOR \SUBBYTES[0].a/U5006  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3291 ), .Z(\SUBBYTES[0].a/n794 ) );
  XOR \SUBBYTES[0].a/U5005  ( .A(\SUBBYTES[0].a/n796 ), .B(
        \SUBBYTES[0].a/n795 ), .Z(\SUBBYTES[0].a/w3315 ) );
  XOR \SUBBYTES[0].a/U5004  ( .A(\SUBBYTES[0].a/n1510 ), .B(
        \SUBBYTES[0].a/n797 ), .Z(\SUBBYTES[0].a/n795 ) );
  XOR \SUBBYTES[0].a/U5003  ( .A(\w1[0][6] ), .B(\SUBBYTES[0].a/w3357 ), .Z(
        \SUBBYTES[0].a/n796 ) );
  XOR \SUBBYTES[0].a/U5002  ( .A(\SUBBYTES[0].a/w3296 ), .B(
        \SUBBYTES[0].a/w3297 ), .Z(\SUBBYTES[0].a/n797 ) );
  XOR \SUBBYTES[0].a/U5001  ( .A(\SUBBYTES[0].a/n1508 ), .B(
        \SUBBYTES[0].a/n1507 ), .Z(\SUBBYTES[0].a/w3335 ) );
  XOR \SUBBYTES[0].a/U5000  ( .A(\SUBBYTES[0].a/n799 ), .B(
        \SUBBYTES[0].a/n798 ), .Z(\SUBBYTES[0].a/w3336 ) );
  XOR \SUBBYTES[0].a/U4999  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/n1509 ), .Z(
        \SUBBYTES[0].a/n798 ) );
  XOR \SUBBYTES[0].a/U4998  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3297 ), .Z(\SUBBYTES[0].a/n799 ) );
  XOR \SUBBYTES[0].a/U4997  ( .A(\SUBBYTES[0].a/n801 ), .B(
        \SUBBYTES[0].a/n800 ), .Z(\SUBBYTES[0].a/w3312 ) );
  XOR \SUBBYTES[0].a/U4996  ( .A(\SUBBYTES[0].a/n803 ), .B(
        \SUBBYTES[0].a/n802 ), .Z(\SUBBYTES[0].a/n800 ) );
  XOR \SUBBYTES[0].a/U4995  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/w3396 ), .Z(
        \SUBBYTES[0].a/n801 ) );
  XOR \SUBBYTES[0].a/U4994  ( .A(\SUBBYTES[0].a/w3303 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n802 ) );
  XOR \SUBBYTES[0].a/U4993  ( .A(\SUBBYTES[0].a/w3289 ), .B(
        \SUBBYTES[0].a/w3291 ), .Z(\SUBBYTES[0].a/n803 ) );
  XOR \SUBBYTES[0].a/U4992  ( .A(\SUBBYTES[0].a/n805 ), .B(
        \SUBBYTES[0].a/n804 ), .Z(\SUBBYTES[0].a/w3313 ) );
  XOR \SUBBYTES[0].a/U4991  ( .A(\SUBBYTES[0].a/n1510 ), .B(
        \SUBBYTES[0].a/n806 ), .Z(\SUBBYTES[0].a/n804 ) );
  XOR \SUBBYTES[0].a/U4990  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n1511 ), .Z(
        \SUBBYTES[0].a/n805 ) );
  XOR \SUBBYTES[0].a/U4989  ( .A(\SUBBYTES[0].a/w3303 ), .B(
        \SUBBYTES[0].a/w3304 ), .Z(\SUBBYTES[0].a/n806 ) );
  XOR \SUBBYTES[0].a/U4988  ( .A(\SUBBYTES[0].a/n808 ), .B(
        \SUBBYTES[0].a/n807 ), .Z(\SUBBYTES[0].a/w3329 ) );
  XOR \SUBBYTES[0].a/U4987  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n809 ), .Z(
        \SUBBYTES[0].a/n807 ) );
  XOR \SUBBYTES[0].a/U4986  ( .A(\SUBBYTES[0].a/w3304 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n808 ) );
  XOR \SUBBYTES[0].a/U4985  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3289 ), .Z(\SUBBYTES[0].a/n809 ) );
  XOR \SUBBYTES[0].a/U4984  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n810 ), .Z(
        \SUBBYTES[0].a/n1512 ) );
  XOR \SUBBYTES[0].a/U4983  ( .A(\w1[0][11] ), .B(\w1[0][10] ), .Z(
        \SUBBYTES[0].a/n810 ) );
  XOR \SUBBYTES[0].a/U4982  ( .A(\w1[0][14] ), .B(\SUBBYTES[0].a/n1512 ), .Z(
        \SUBBYTES[0].a/w3171 ) );
  XOR \SUBBYTES[0].a/U4981  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/w3058 ) );
  XOR \SUBBYTES[0].a/U4980  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/n811 ), .Z(
        \SUBBYTES[0].a/w3059 ) );
  XOR \SUBBYTES[0].a/U4979  ( .A(\w1[0][14] ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n811 ) );
  XOR \SUBBYTES[0].a/U4978  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n1512 ), .Z(
        \SUBBYTES[0].a/w3189 ) );
  XOR \SUBBYTES[0].a/U4977  ( .A(\SUBBYTES[0].a/n813 ), .B(
        \SUBBYTES[0].a/n812 ), .Z(\SUBBYTES[0].a/w3182 ) );
  XOR \SUBBYTES[0].a/U4976  ( .A(\w1[0][11] ), .B(\w1[0][9] ), .Z(
        \SUBBYTES[0].a/n812 ) );
  XOR \SUBBYTES[0].a/U4975  ( .A(\w1[0][15] ), .B(\w1[0][12] ), .Z(
        \SUBBYTES[0].a/n813 ) );
  XOR \SUBBYTES[0].a/U4974  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3182 ), .Z(
        \SUBBYTES[0].a/w3061 ) );
  XOR \SUBBYTES[0].a/U4973  ( .A(\SUBBYTES[0].a/n815 ), .B(
        \SUBBYTES[0].a/n814 ), .Z(\SUBBYTES[0].a/w3169 ) );
  XOR \SUBBYTES[0].a/U4972  ( .A(\SUBBYTES[0].a/w3130 ), .B(n15), .Z(
        \SUBBYTES[0].a/n814 ) );
  XOR \SUBBYTES[0].a/U4971  ( .A(\SUBBYTES[0].a/w3123 ), .B(
        \SUBBYTES[0].a/w3126 ), .Z(\SUBBYTES[0].a/n815 ) );
  XOR \SUBBYTES[0].a/U4970  ( .A(\SUBBYTES[0].a/n817 ), .B(
        \SUBBYTES[0].a/n816 ), .Z(\SUBBYTES[0].a/w3170 ) );
  XOR \SUBBYTES[0].a/U4969  ( .A(\SUBBYTES[0].a/w3130 ), .B(
        \SUBBYTES[0].a/n150 ), .Z(\SUBBYTES[0].a/n816 ) );
  XOR \SUBBYTES[0].a/U4968  ( .A(\SUBBYTES[0].a/w3123 ), .B(
        \SUBBYTES[0].a/n149 ), .Z(\SUBBYTES[0].a/n817 ) );
  XOR \SUBBYTES[0].a/U4967  ( .A(\SUBBYTES[0].a/w3182 ), .B(
        \SUBBYTES[0].a/n818 ), .Z(\SUBBYTES[0].a/w3172 ) );
  XOR \SUBBYTES[0].a/U4966  ( .A(\w1[0][14] ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n818 ) );
  XOR \SUBBYTES[0].a/U4965  ( .A(\SUBBYTES[0].a/n820 ), .B(
        \SUBBYTES[0].a/n819 ), .Z(\SUBBYTES[0].a/w3173 ) );
  XOR \SUBBYTES[0].a/U4964  ( .A(\SUBBYTES[0].a/n150 ), .B(n15), .Z(
        \SUBBYTES[0].a/n819 ) );
  XOR \SUBBYTES[0].a/U4963  ( .A(\SUBBYTES[0].a/n149 ), .B(
        \SUBBYTES[0].a/w3126 ), .Z(\SUBBYTES[0].a/n820 ) );
  XOR \SUBBYTES[0].a/U4962  ( .A(\w1[0][15] ), .B(\w1[0][10] ), .Z(
        \SUBBYTES[0].a/n1518 ) );
  XOR \SUBBYTES[0].a/U4961  ( .A(\SUBBYTES[0].a/n1518 ), .B(
        \SUBBYTES[0].a/n821 ), .Z(\SUBBYTES[0].a/w3174 ) );
  XOR \SUBBYTES[0].a/U4960  ( .A(\w1[0][13] ), .B(\w1[0][12] ), .Z(
        \SUBBYTES[0].a/n821 ) );
  XOR \SUBBYTES[0].a/U4959  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3062 ) );
  XOR \SUBBYTES[0].a/U4958  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3063 ) );
  XOR \SUBBYTES[0].a/U4957  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3064 ) );
  XOR \SUBBYTES[0].a/U4956  ( .A(\SUBBYTES[0].a/w3063 ), .B(
        \SUBBYTES[0].a/n1518 ), .Z(\SUBBYTES[0].a/w3065 ) );
  XOR \SUBBYTES[0].a/U4955  ( .A(\SUBBYTES[0].a/n1518 ), .B(
        \SUBBYTES[0].a/n822 ), .Z(\SUBBYTES[0].a/w3150 ) );
  XOR \SUBBYTES[0].a/U4954  ( .A(\w1[0][12] ), .B(\w1[0][9] ), .Z(
        \SUBBYTES[0].a/n822 ) );
  XOR \SUBBYTES[0].a/U4953  ( .A(\SUBBYTES[0].a/n824 ), .B(
        \SUBBYTES[0].a/n823 ), .Z(\SUBBYTES[0].a/n1515 ) );
  XOR \SUBBYTES[0].a/U4952  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/n825 ), .Z(
        \SUBBYTES[0].a/n823 ) );
  XOR \SUBBYTES[0].a/U4951  ( .A(\SUBBYTES[0].a/w3115 ), .B(\w1[0][14] ), .Z(
        \SUBBYTES[0].a/n824 ) );
  XOR \SUBBYTES[0].a/U4950  ( .A(\SUBBYTES[0].a/w3089 ), .B(
        \SUBBYTES[0].a/w3096 ), .Z(\SUBBYTES[0].a/n825 ) );
  XOR \SUBBYTES[0].a/U4949  ( .A(\SUBBYTES[0].a/n827 ), .B(
        \SUBBYTES[0].a/n826 ), .Z(\SUBBYTES[0].a/n1513 ) );
  XOR \SUBBYTES[0].a/U4948  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n828 ), .Z(
        \SUBBYTES[0].a/n826 ) );
  XOR \SUBBYTES[0].a/U4947  ( .A(\SUBBYTES[0].a/w3114 ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n827 ) );
  XOR \SUBBYTES[0].a/U4946  ( .A(\SUBBYTES[0].a/w3090 ), .B(
        \SUBBYTES[0].a/w3097 ), .Z(\SUBBYTES[0].a/n828 ) );
  XOR \SUBBYTES[0].a/U4945  ( .A(\SUBBYTES[0].a/n1515 ), .B(
        \SUBBYTES[0].a/n1513 ), .Z(\SUBBYTES[0].a/w3120 ) );
  XOR \SUBBYTES[0].a/U4944  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n829 ), .Z(
        \SUBBYTES[0].a/n1516 ) );
  XOR \SUBBYTES[0].a/U4943  ( .A(\SUBBYTES[0].a/w3082 ), .B(
        \SUBBYTES[0].a/w3092 ), .Z(\SUBBYTES[0].a/n829 ) );
  XOR \SUBBYTES[0].a/U4942  ( .A(\SUBBYTES[0].a/n831 ), .B(
        \SUBBYTES[0].a/n830 ), .Z(\SUBBYTES[0].a/w3107 ) );
  XOR \SUBBYTES[0].a/U4941  ( .A(\SUBBYTES[0].a/n1516 ), .B(
        \SUBBYTES[0].a/n832 ), .Z(\SUBBYTES[0].a/n830 ) );
  XOR \SUBBYTES[0].a/U4940  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/n831 ) );
  XOR \SUBBYTES[0].a/U4939  ( .A(\SUBBYTES[0].a/w3084 ), .B(
        \SUBBYTES[0].a/w3089 ), .Z(\SUBBYTES[0].a/n832 ) );
  XOR \SUBBYTES[0].a/U4938  ( .A(\SUBBYTES[0].a/n834 ), .B(
        \SUBBYTES[0].a/n833 ), .Z(\SUBBYTES[0].a/n1514 ) );
  XOR \SUBBYTES[0].a/U4937  ( .A(\SUBBYTES[0].a/w3117 ), .B(\w1[0][15] ), .Z(
        \SUBBYTES[0].a/n833 ) );
  XOR \SUBBYTES[0].a/U4936  ( .A(\SUBBYTES[0].a/w3092 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n834 ) );
  XOR \SUBBYTES[0].a/U4935  ( .A(\SUBBYTES[0].a/n1513 ), .B(
        \SUBBYTES[0].a/n1514 ), .Z(\SUBBYTES[0].a/w3119 ) );
  XOR \SUBBYTES[0].a/U4934  ( .A(\w1[0][11] ), .B(\SUBBYTES[0].a/n835 ), .Z(
        \SUBBYTES[0].a/n1517 ) );
  XOR \SUBBYTES[0].a/U4933  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3084 ), .Z(\SUBBYTES[0].a/n835 ) );
  XOR \SUBBYTES[0].a/U4932  ( .A(\SUBBYTES[0].a/n837 ), .B(
        \SUBBYTES[0].a/n836 ), .Z(\SUBBYTES[0].a/w3108 ) );
  XOR \SUBBYTES[0].a/U4931  ( .A(\SUBBYTES[0].a/n1517 ), .B(
        \SUBBYTES[0].a/n838 ), .Z(\SUBBYTES[0].a/n836 ) );
  XOR \SUBBYTES[0].a/U4930  ( .A(\w1[0][14] ), .B(\SUBBYTES[0].a/w3150 ), .Z(
        \SUBBYTES[0].a/n837 ) );
  XOR \SUBBYTES[0].a/U4929  ( .A(\SUBBYTES[0].a/w3089 ), .B(
        \SUBBYTES[0].a/w3090 ), .Z(\SUBBYTES[0].a/n838 ) );
  XOR \SUBBYTES[0].a/U4928  ( .A(\SUBBYTES[0].a/n1515 ), .B(
        \SUBBYTES[0].a/n1514 ), .Z(\SUBBYTES[0].a/w3128 ) );
  XOR \SUBBYTES[0].a/U4927  ( .A(\SUBBYTES[0].a/n840 ), .B(
        \SUBBYTES[0].a/n839 ), .Z(\SUBBYTES[0].a/w3129 ) );
  XOR \SUBBYTES[0].a/U4926  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/n1516 ), .Z(
        \SUBBYTES[0].a/n839 ) );
  XOR \SUBBYTES[0].a/U4925  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3090 ), .Z(\SUBBYTES[0].a/n840 ) );
  XOR \SUBBYTES[0].a/U4924  ( .A(\SUBBYTES[0].a/n842 ), .B(
        \SUBBYTES[0].a/n841 ), .Z(\SUBBYTES[0].a/w3105 ) );
  XOR \SUBBYTES[0].a/U4923  ( .A(\SUBBYTES[0].a/n844 ), .B(
        \SUBBYTES[0].a/n843 ), .Z(\SUBBYTES[0].a/n841 ) );
  XOR \SUBBYTES[0].a/U4922  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/w3189 ), .Z(
        \SUBBYTES[0].a/n842 ) );
  XOR \SUBBYTES[0].a/U4921  ( .A(\SUBBYTES[0].a/w3096 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n843 ) );
  XOR \SUBBYTES[0].a/U4920  ( .A(\SUBBYTES[0].a/w3082 ), .B(
        \SUBBYTES[0].a/w3084 ), .Z(\SUBBYTES[0].a/n844 ) );
  XOR \SUBBYTES[0].a/U4919  ( .A(\SUBBYTES[0].a/n846 ), .B(
        \SUBBYTES[0].a/n845 ), .Z(\SUBBYTES[0].a/w3106 ) );
  XOR \SUBBYTES[0].a/U4918  ( .A(\SUBBYTES[0].a/n1517 ), .B(
        \SUBBYTES[0].a/n847 ), .Z(\SUBBYTES[0].a/n845 ) );
  XOR \SUBBYTES[0].a/U4917  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n1518 ), .Z(
        \SUBBYTES[0].a/n846 ) );
  XOR \SUBBYTES[0].a/U4916  ( .A(\SUBBYTES[0].a/w3096 ), .B(
        \SUBBYTES[0].a/w3097 ), .Z(\SUBBYTES[0].a/n847 ) );
  XOR \SUBBYTES[0].a/U4915  ( .A(\SUBBYTES[0].a/n849 ), .B(
        \SUBBYTES[0].a/n848 ), .Z(\SUBBYTES[0].a/w3122 ) );
  XOR \SUBBYTES[0].a/U4914  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n850 ), .Z(
        \SUBBYTES[0].a/n848 ) );
  XOR \SUBBYTES[0].a/U4913  ( .A(\SUBBYTES[0].a/w3097 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n849 ) );
  XOR \SUBBYTES[0].a/U4912  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3082 ), .Z(\SUBBYTES[0].a/n850 ) );
  XOR \SUBBYTES[0].a/U4911  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n851 ), .Z(
        \SUBBYTES[0].a/n1519 ) );
  XOR \SUBBYTES[0].a/U4910  ( .A(\w1[0][19] ), .B(\w1[0][18] ), .Z(
        \SUBBYTES[0].a/n851 ) );
  XOR \SUBBYTES[0].a/U4909  ( .A(\w1[0][22] ), .B(\SUBBYTES[0].a/n1519 ), .Z(
        \SUBBYTES[0].a/w2964 ) );
  XOR \SUBBYTES[0].a/U4908  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/w2851 ) );
  XOR \SUBBYTES[0].a/U4907  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/n852 ), .Z(
        \SUBBYTES[0].a/w2852 ) );
  XOR \SUBBYTES[0].a/U4906  ( .A(\w1[0][22] ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n852 ) );
  XOR \SUBBYTES[0].a/U4905  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n1519 ), .Z(
        \SUBBYTES[0].a/w2982 ) );
  XOR \SUBBYTES[0].a/U4904  ( .A(\SUBBYTES[0].a/n854 ), .B(
        \SUBBYTES[0].a/n853 ), .Z(\SUBBYTES[0].a/w2975 ) );
  XOR \SUBBYTES[0].a/U4903  ( .A(\w1[0][19] ), .B(\w1[0][17] ), .Z(
        \SUBBYTES[0].a/n853 ) );
  XOR \SUBBYTES[0].a/U4902  ( .A(\w1[0][23] ), .B(\w1[0][20] ), .Z(
        \SUBBYTES[0].a/n854 ) );
  XOR \SUBBYTES[0].a/U4901  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2975 ), .Z(
        \SUBBYTES[0].a/w2854 ) );
  XOR \SUBBYTES[0].a/U4900  ( .A(\SUBBYTES[0].a/n856 ), .B(
        \SUBBYTES[0].a/n855 ), .Z(\SUBBYTES[0].a/w2962 ) );
  XOR \SUBBYTES[0].a/U4899  ( .A(\SUBBYTES[0].a/w2923 ), .B(n14), .Z(
        \SUBBYTES[0].a/n855 ) );
  XOR \SUBBYTES[0].a/U4898  ( .A(\SUBBYTES[0].a/w2916 ), .B(
        \SUBBYTES[0].a/w2919 ), .Z(\SUBBYTES[0].a/n856 ) );
  XOR \SUBBYTES[0].a/U4897  ( .A(\SUBBYTES[0].a/n858 ), .B(
        \SUBBYTES[0].a/n857 ), .Z(\SUBBYTES[0].a/w2963 ) );
  XOR \SUBBYTES[0].a/U4896  ( .A(\SUBBYTES[0].a/w2923 ), .B(
        \SUBBYTES[0].a/n140 ), .Z(\SUBBYTES[0].a/n857 ) );
  XOR \SUBBYTES[0].a/U4895  ( .A(\SUBBYTES[0].a/w2916 ), .B(
        \SUBBYTES[0].a/n139 ), .Z(\SUBBYTES[0].a/n858 ) );
  XOR \SUBBYTES[0].a/U4894  ( .A(\SUBBYTES[0].a/w2975 ), .B(
        \SUBBYTES[0].a/n859 ), .Z(\SUBBYTES[0].a/w2965 ) );
  XOR \SUBBYTES[0].a/U4893  ( .A(\w1[0][22] ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n859 ) );
  XOR \SUBBYTES[0].a/U4892  ( .A(\SUBBYTES[0].a/n861 ), .B(
        \SUBBYTES[0].a/n860 ), .Z(\SUBBYTES[0].a/w2966 ) );
  XOR \SUBBYTES[0].a/U4891  ( .A(\SUBBYTES[0].a/n140 ), .B(n14), .Z(
        \SUBBYTES[0].a/n860 ) );
  XOR \SUBBYTES[0].a/U4890  ( .A(\SUBBYTES[0].a/n139 ), .B(
        \SUBBYTES[0].a/w2919 ), .Z(\SUBBYTES[0].a/n861 ) );
  XOR \SUBBYTES[0].a/U4889  ( .A(\w1[0][23] ), .B(\w1[0][18] ), .Z(
        \SUBBYTES[0].a/n1525 ) );
  XOR \SUBBYTES[0].a/U4888  ( .A(\SUBBYTES[0].a/n1525 ), .B(
        \SUBBYTES[0].a/n862 ), .Z(\SUBBYTES[0].a/w2967 ) );
  XOR \SUBBYTES[0].a/U4887  ( .A(\w1[0][21] ), .B(\w1[0][20] ), .Z(
        \SUBBYTES[0].a/n862 ) );
  XOR \SUBBYTES[0].a/U4886  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2855 ) );
  XOR \SUBBYTES[0].a/U4885  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2856 ) );
  XOR \SUBBYTES[0].a/U4884  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2857 ) );
  XOR \SUBBYTES[0].a/U4883  ( .A(\SUBBYTES[0].a/w2856 ), .B(
        \SUBBYTES[0].a/n1525 ), .Z(\SUBBYTES[0].a/w2858 ) );
  XOR \SUBBYTES[0].a/U4882  ( .A(\SUBBYTES[0].a/n1525 ), .B(
        \SUBBYTES[0].a/n863 ), .Z(\SUBBYTES[0].a/w2943 ) );
  XOR \SUBBYTES[0].a/U4881  ( .A(\w1[0][20] ), .B(\w1[0][17] ), .Z(
        \SUBBYTES[0].a/n863 ) );
  XOR \SUBBYTES[0].a/U4880  ( .A(\SUBBYTES[0].a/n865 ), .B(
        \SUBBYTES[0].a/n864 ), .Z(\SUBBYTES[0].a/n1522 ) );
  XOR \SUBBYTES[0].a/U4879  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/n866 ), .Z(
        \SUBBYTES[0].a/n864 ) );
  XOR \SUBBYTES[0].a/U4878  ( .A(\SUBBYTES[0].a/w2908 ), .B(\w1[0][22] ), .Z(
        \SUBBYTES[0].a/n865 ) );
  XOR \SUBBYTES[0].a/U4877  ( .A(\SUBBYTES[0].a/w2882 ), .B(
        \SUBBYTES[0].a/w2889 ), .Z(\SUBBYTES[0].a/n866 ) );
  XOR \SUBBYTES[0].a/U4876  ( .A(\SUBBYTES[0].a/n868 ), .B(
        \SUBBYTES[0].a/n867 ), .Z(\SUBBYTES[0].a/n1520 ) );
  XOR \SUBBYTES[0].a/U4875  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n869 ), .Z(
        \SUBBYTES[0].a/n867 ) );
  XOR \SUBBYTES[0].a/U4874  ( .A(\SUBBYTES[0].a/w2907 ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n868 ) );
  XOR \SUBBYTES[0].a/U4873  ( .A(\SUBBYTES[0].a/w2883 ), .B(
        \SUBBYTES[0].a/w2890 ), .Z(\SUBBYTES[0].a/n869 ) );
  XOR \SUBBYTES[0].a/U4872  ( .A(\SUBBYTES[0].a/n1522 ), .B(
        \SUBBYTES[0].a/n1520 ), .Z(\SUBBYTES[0].a/w2913 ) );
  XOR \SUBBYTES[0].a/U4871  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n870 ), .Z(
        \SUBBYTES[0].a/n1523 ) );
  XOR \SUBBYTES[0].a/U4870  ( .A(\SUBBYTES[0].a/w2875 ), .B(
        \SUBBYTES[0].a/w2885 ), .Z(\SUBBYTES[0].a/n870 ) );
  XOR \SUBBYTES[0].a/U4869  ( .A(\SUBBYTES[0].a/n872 ), .B(
        \SUBBYTES[0].a/n871 ), .Z(\SUBBYTES[0].a/w2900 ) );
  XOR \SUBBYTES[0].a/U4868  ( .A(\SUBBYTES[0].a/n1523 ), .B(
        \SUBBYTES[0].a/n873 ), .Z(\SUBBYTES[0].a/n871 ) );
  XOR \SUBBYTES[0].a/U4867  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/n872 ) );
  XOR \SUBBYTES[0].a/U4866  ( .A(\SUBBYTES[0].a/w2877 ), .B(
        \SUBBYTES[0].a/w2882 ), .Z(\SUBBYTES[0].a/n873 ) );
  XOR \SUBBYTES[0].a/U4865  ( .A(\SUBBYTES[0].a/n875 ), .B(
        \SUBBYTES[0].a/n874 ), .Z(\SUBBYTES[0].a/n1521 ) );
  XOR \SUBBYTES[0].a/U4864  ( .A(\SUBBYTES[0].a/w2910 ), .B(\w1[0][23] ), .Z(
        \SUBBYTES[0].a/n874 ) );
  XOR \SUBBYTES[0].a/U4863  ( .A(\SUBBYTES[0].a/w2885 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n875 ) );
  XOR \SUBBYTES[0].a/U4862  ( .A(\SUBBYTES[0].a/n1520 ), .B(
        \SUBBYTES[0].a/n1521 ), .Z(\SUBBYTES[0].a/w2912 ) );
  XOR \SUBBYTES[0].a/U4861  ( .A(\w1[0][19] ), .B(\SUBBYTES[0].a/n876 ), .Z(
        \SUBBYTES[0].a/n1524 ) );
  XOR \SUBBYTES[0].a/U4860  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2877 ), .Z(\SUBBYTES[0].a/n876 ) );
  XOR \SUBBYTES[0].a/U4859  ( .A(\SUBBYTES[0].a/n878 ), .B(
        \SUBBYTES[0].a/n877 ), .Z(\SUBBYTES[0].a/w2901 ) );
  XOR \SUBBYTES[0].a/U4858  ( .A(\SUBBYTES[0].a/n1524 ), .B(
        \SUBBYTES[0].a/n879 ), .Z(\SUBBYTES[0].a/n877 ) );
  XOR \SUBBYTES[0].a/U4857  ( .A(\w1[0][22] ), .B(\SUBBYTES[0].a/w2943 ), .Z(
        \SUBBYTES[0].a/n878 ) );
  XOR \SUBBYTES[0].a/U4856  ( .A(\SUBBYTES[0].a/w2882 ), .B(
        \SUBBYTES[0].a/w2883 ), .Z(\SUBBYTES[0].a/n879 ) );
  XOR \SUBBYTES[0].a/U4855  ( .A(\SUBBYTES[0].a/n1522 ), .B(
        \SUBBYTES[0].a/n1521 ), .Z(\SUBBYTES[0].a/w2921 ) );
  XOR \SUBBYTES[0].a/U4854  ( .A(\SUBBYTES[0].a/n881 ), .B(
        \SUBBYTES[0].a/n880 ), .Z(\SUBBYTES[0].a/w2922 ) );
  XOR \SUBBYTES[0].a/U4853  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/n1523 ), .Z(
        \SUBBYTES[0].a/n880 ) );
  XOR \SUBBYTES[0].a/U4852  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2883 ), .Z(\SUBBYTES[0].a/n881 ) );
  XOR \SUBBYTES[0].a/U4851  ( .A(\SUBBYTES[0].a/n883 ), .B(
        \SUBBYTES[0].a/n882 ), .Z(\SUBBYTES[0].a/w2898 ) );
  XOR \SUBBYTES[0].a/U4850  ( .A(\SUBBYTES[0].a/n885 ), .B(
        \SUBBYTES[0].a/n884 ), .Z(\SUBBYTES[0].a/n882 ) );
  XOR \SUBBYTES[0].a/U4849  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/w2982 ), .Z(
        \SUBBYTES[0].a/n883 ) );
  XOR \SUBBYTES[0].a/U4848  ( .A(\SUBBYTES[0].a/w2889 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n884 ) );
  XOR \SUBBYTES[0].a/U4847  ( .A(\SUBBYTES[0].a/w2875 ), .B(
        \SUBBYTES[0].a/w2877 ), .Z(\SUBBYTES[0].a/n885 ) );
  XOR \SUBBYTES[0].a/U4846  ( .A(\SUBBYTES[0].a/n887 ), .B(
        \SUBBYTES[0].a/n886 ), .Z(\SUBBYTES[0].a/w2899 ) );
  XOR \SUBBYTES[0].a/U4845  ( .A(\SUBBYTES[0].a/n1524 ), .B(
        \SUBBYTES[0].a/n888 ), .Z(\SUBBYTES[0].a/n886 ) );
  XOR \SUBBYTES[0].a/U4844  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n1525 ), .Z(
        \SUBBYTES[0].a/n887 ) );
  XOR \SUBBYTES[0].a/U4843  ( .A(\SUBBYTES[0].a/w2889 ), .B(
        \SUBBYTES[0].a/w2890 ), .Z(\SUBBYTES[0].a/n888 ) );
  XOR \SUBBYTES[0].a/U4842  ( .A(\SUBBYTES[0].a/n890 ), .B(
        \SUBBYTES[0].a/n889 ), .Z(\SUBBYTES[0].a/w2915 ) );
  XOR \SUBBYTES[0].a/U4841  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n891 ), .Z(
        \SUBBYTES[0].a/n889 ) );
  XOR \SUBBYTES[0].a/U4840  ( .A(\SUBBYTES[0].a/w2890 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n890 ) );
  XOR \SUBBYTES[0].a/U4839  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2875 ), .Z(\SUBBYTES[0].a/n891 ) );
  XOR \SUBBYTES[0].a/U4838  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n892 ), .Z(
        \SUBBYTES[0].a/n1526 ) );
  XOR \SUBBYTES[0].a/U4837  ( .A(\w1[0][27] ), .B(\w1[0][26] ), .Z(
        \SUBBYTES[0].a/n892 ) );
  XOR \SUBBYTES[0].a/U4836  ( .A(\w1[0][30] ), .B(\SUBBYTES[0].a/n1526 ), .Z(
        \SUBBYTES[0].a/w2757 ) );
  XOR \SUBBYTES[0].a/U4835  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/w2644 ) );
  XOR \SUBBYTES[0].a/U4834  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/n893 ), .Z(
        \SUBBYTES[0].a/w2645 ) );
  XOR \SUBBYTES[0].a/U4833  ( .A(\w1[0][30] ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n893 ) );
  XOR \SUBBYTES[0].a/U4832  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n1526 ), .Z(
        \SUBBYTES[0].a/w2775 ) );
  XOR \SUBBYTES[0].a/U4831  ( .A(\SUBBYTES[0].a/n895 ), .B(
        \SUBBYTES[0].a/n894 ), .Z(\SUBBYTES[0].a/w2768 ) );
  XOR \SUBBYTES[0].a/U4830  ( .A(\w1[0][27] ), .B(\w1[0][25] ), .Z(
        \SUBBYTES[0].a/n894 ) );
  XOR \SUBBYTES[0].a/U4829  ( .A(\w1[0][31] ), .B(\w1[0][28] ), .Z(
        \SUBBYTES[0].a/n895 ) );
  XOR \SUBBYTES[0].a/U4828  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2768 ), .Z(
        \SUBBYTES[0].a/w2647 ) );
  XOR \SUBBYTES[0].a/U4827  ( .A(\SUBBYTES[0].a/n897 ), .B(
        \SUBBYTES[0].a/n896 ), .Z(\SUBBYTES[0].a/w2755 ) );
  XOR \SUBBYTES[0].a/U4826  ( .A(\SUBBYTES[0].a/w2716 ), .B(n13), .Z(
        \SUBBYTES[0].a/n896 ) );
  XOR \SUBBYTES[0].a/U4825  ( .A(\SUBBYTES[0].a/w2709 ), .B(
        \SUBBYTES[0].a/w2712 ), .Z(\SUBBYTES[0].a/n897 ) );
  XOR \SUBBYTES[0].a/U4824  ( .A(\SUBBYTES[0].a/n899 ), .B(
        \SUBBYTES[0].a/n898 ), .Z(\SUBBYTES[0].a/w2756 ) );
  XOR \SUBBYTES[0].a/U4823  ( .A(\SUBBYTES[0].a/w2716 ), .B(
        \SUBBYTES[0].a/n130 ), .Z(\SUBBYTES[0].a/n898 ) );
  XOR \SUBBYTES[0].a/U4822  ( .A(\SUBBYTES[0].a/w2709 ), .B(
        \SUBBYTES[0].a/n129 ), .Z(\SUBBYTES[0].a/n899 ) );
  XOR \SUBBYTES[0].a/U4821  ( .A(\SUBBYTES[0].a/w2768 ), .B(
        \SUBBYTES[0].a/n900 ), .Z(\SUBBYTES[0].a/w2758 ) );
  XOR \SUBBYTES[0].a/U4820  ( .A(\w1[0][30] ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n900 ) );
  XOR \SUBBYTES[0].a/U4819  ( .A(\SUBBYTES[0].a/n902 ), .B(
        \SUBBYTES[0].a/n901 ), .Z(\SUBBYTES[0].a/w2759 ) );
  XOR \SUBBYTES[0].a/U4818  ( .A(\SUBBYTES[0].a/n130 ), .B(n13), .Z(
        \SUBBYTES[0].a/n901 ) );
  XOR \SUBBYTES[0].a/U4817  ( .A(\SUBBYTES[0].a/n129 ), .B(
        \SUBBYTES[0].a/w2712 ), .Z(\SUBBYTES[0].a/n902 ) );
  XOR \SUBBYTES[0].a/U4816  ( .A(\w1[0][31] ), .B(\w1[0][26] ), .Z(
        \SUBBYTES[0].a/n1532 ) );
  XOR \SUBBYTES[0].a/U4815  ( .A(\SUBBYTES[0].a/n1532 ), .B(
        \SUBBYTES[0].a/n903 ), .Z(\SUBBYTES[0].a/w2760 ) );
  XOR \SUBBYTES[0].a/U4814  ( .A(\w1[0][29] ), .B(\w1[0][28] ), .Z(
        \SUBBYTES[0].a/n903 ) );
  XOR \SUBBYTES[0].a/U4813  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2648 ) );
  XOR \SUBBYTES[0].a/U4812  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2649 ) );
  XOR \SUBBYTES[0].a/U4811  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2650 ) );
  XOR \SUBBYTES[0].a/U4810  ( .A(\SUBBYTES[0].a/w2649 ), .B(
        \SUBBYTES[0].a/n1532 ), .Z(\SUBBYTES[0].a/w2651 ) );
  XOR \SUBBYTES[0].a/U4809  ( .A(\SUBBYTES[0].a/n1532 ), .B(
        \SUBBYTES[0].a/n904 ), .Z(\SUBBYTES[0].a/w2736 ) );
  XOR \SUBBYTES[0].a/U4808  ( .A(\w1[0][28] ), .B(\w1[0][25] ), .Z(
        \SUBBYTES[0].a/n904 ) );
  XOR \SUBBYTES[0].a/U4807  ( .A(\SUBBYTES[0].a/n906 ), .B(
        \SUBBYTES[0].a/n905 ), .Z(\SUBBYTES[0].a/n1529 ) );
  XOR \SUBBYTES[0].a/U4806  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/n907 ), .Z(
        \SUBBYTES[0].a/n905 ) );
  XOR \SUBBYTES[0].a/U4805  ( .A(\SUBBYTES[0].a/w2701 ), .B(\w1[0][30] ), .Z(
        \SUBBYTES[0].a/n906 ) );
  XOR \SUBBYTES[0].a/U4804  ( .A(\SUBBYTES[0].a/w2675 ), .B(
        \SUBBYTES[0].a/w2682 ), .Z(\SUBBYTES[0].a/n907 ) );
  XOR \SUBBYTES[0].a/U4803  ( .A(\SUBBYTES[0].a/n909 ), .B(
        \SUBBYTES[0].a/n908 ), .Z(\SUBBYTES[0].a/n1527 ) );
  XOR \SUBBYTES[0].a/U4802  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n910 ), .Z(
        \SUBBYTES[0].a/n908 ) );
  XOR \SUBBYTES[0].a/U4801  ( .A(\SUBBYTES[0].a/w2700 ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n909 ) );
  XOR \SUBBYTES[0].a/U4800  ( .A(\SUBBYTES[0].a/w2676 ), .B(
        \SUBBYTES[0].a/w2683 ), .Z(\SUBBYTES[0].a/n910 ) );
  XOR \SUBBYTES[0].a/U4799  ( .A(\SUBBYTES[0].a/n1529 ), .B(
        \SUBBYTES[0].a/n1527 ), .Z(\SUBBYTES[0].a/w2706 ) );
  XOR \SUBBYTES[0].a/U4798  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n911 ), .Z(
        \SUBBYTES[0].a/n1530 ) );
  XOR \SUBBYTES[0].a/U4797  ( .A(\SUBBYTES[0].a/w2668 ), .B(
        \SUBBYTES[0].a/w2678 ), .Z(\SUBBYTES[0].a/n911 ) );
  XOR \SUBBYTES[0].a/U4796  ( .A(\SUBBYTES[0].a/n913 ), .B(
        \SUBBYTES[0].a/n912 ), .Z(\SUBBYTES[0].a/w2693 ) );
  XOR \SUBBYTES[0].a/U4795  ( .A(\SUBBYTES[0].a/n1530 ), .B(
        \SUBBYTES[0].a/n914 ), .Z(\SUBBYTES[0].a/n912 ) );
  XOR \SUBBYTES[0].a/U4794  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/n913 ) );
  XOR \SUBBYTES[0].a/U4793  ( .A(\SUBBYTES[0].a/w2670 ), .B(
        \SUBBYTES[0].a/w2675 ), .Z(\SUBBYTES[0].a/n914 ) );
  XOR \SUBBYTES[0].a/U4792  ( .A(\SUBBYTES[0].a/n916 ), .B(
        \SUBBYTES[0].a/n915 ), .Z(\SUBBYTES[0].a/n1528 ) );
  XOR \SUBBYTES[0].a/U4791  ( .A(\SUBBYTES[0].a/w2703 ), .B(\w1[0][31] ), .Z(
        \SUBBYTES[0].a/n915 ) );
  XOR \SUBBYTES[0].a/U4790  ( .A(\SUBBYTES[0].a/w2678 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n916 ) );
  XOR \SUBBYTES[0].a/U4789  ( .A(\SUBBYTES[0].a/n1527 ), .B(
        \SUBBYTES[0].a/n1528 ), .Z(\SUBBYTES[0].a/w2705 ) );
  XOR \SUBBYTES[0].a/U4788  ( .A(\w1[0][27] ), .B(\SUBBYTES[0].a/n917 ), .Z(
        \SUBBYTES[0].a/n1531 ) );
  XOR \SUBBYTES[0].a/U4787  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2670 ), .Z(\SUBBYTES[0].a/n917 ) );
  XOR \SUBBYTES[0].a/U4786  ( .A(\SUBBYTES[0].a/n919 ), .B(
        \SUBBYTES[0].a/n918 ), .Z(\SUBBYTES[0].a/w2694 ) );
  XOR \SUBBYTES[0].a/U4785  ( .A(\SUBBYTES[0].a/n1531 ), .B(
        \SUBBYTES[0].a/n920 ), .Z(\SUBBYTES[0].a/n918 ) );
  XOR \SUBBYTES[0].a/U4784  ( .A(\w1[0][30] ), .B(\SUBBYTES[0].a/w2736 ), .Z(
        \SUBBYTES[0].a/n919 ) );
  XOR \SUBBYTES[0].a/U4783  ( .A(\SUBBYTES[0].a/w2675 ), .B(
        \SUBBYTES[0].a/w2676 ), .Z(\SUBBYTES[0].a/n920 ) );
  XOR \SUBBYTES[0].a/U4782  ( .A(\SUBBYTES[0].a/n1529 ), .B(
        \SUBBYTES[0].a/n1528 ), .Z(\SUBBYTES[0].a/w2714 ) );
  XOR \SUBBYTES[0].a/U4781  ( .A(\SUBBYTES[0].a/n922 ), .B(
        \SUBBYTES[0].a/n921 ), .Z(\SUBBYTES[0].a/w2715 ) );
  XOR \SUBBYTES[0].a/U4780  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/n1530 ), .Z(
        \SUBBYTES[0].a/n921 ) );
  XOR \SUBBYTES[0].a/U4779  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2676 ), .Z(\SUBBYTES[0].a/n922 ) );
  XOR \SUBBYTES[0].a/U4778  ( .A(\SUBBYTES[0].a/n924 ), .B(
        \SUBBYTES[0].a/n923 ), .Z(\SUBBYTES[0].a/w2691 ) );
  XOR \SUBBYTES[0].a/U4777  ( .A(\SUBBYTES[0].a/n926 ), .B(
        \SUBBYTES[0].a/n925 ), .Z(\SUBBYTES[0].a/n923 ) );
  XOR \SUBBYTES[0].a/U4776  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/w2775 ), .Z(
        \SUBBYTES[0].a/n924 ) );
  XOR \SUBBYTES[0].a/U4775  ( .A(\SUBBYTES[0].a/w2682 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n925 ) );
  XOR \SUBBYTES[0].a/U4774  ( .A(\SUBBYTES[0].a/w2668 ), .B(
        \SUBBYTES[0].a/w2670 ), .Z(\SUBBYTES[0].a/n926 ) );
  XOR \SUBBYTES[0].a/U4773  ( .A(\SUBBYTES[0].a/n928 ), .B(
        \SUBBYTES[0].a/n927 ), .Z(\SUBBYTES[0].a/w2692 ) );
  XOR \SUBBYTES[0].a/U4772  ( .A(\SUBBYTES[0].a/n1531 ), .B(
        \SUBBYTES[0].a/n929 ), .Z(\SUBBYTES[0].a/n927 ) );
  XOR \SUBBYTES[0].a/U4771  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n1532 ), .Z(
        \SUBBYTES[0].a/n928 ) );
  XOR \SUBBYTES[0].a/U4770  ( .A(\SUBBYTES[0].a/w2682 ), .B(
        \SUBBYTES[0].a/w2683 ), .Z(\SUBBYTES[0].a/n929 ) );
  XOR \SUBBYTES[0].a/U4769  ( .A(\SUBBYTES[0].a/n931 ), .B(
        \SUBBYTES[0].a/n930 ), .Z(\SUBBYTES[0].a/w2708 ) );
  XOR \SUBBYTES[0].a/U4768  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n932 ), .Z(
        \SUBBYTES[0].a/n930 ) );
  XOR \SUBBYTES[0].a/U4767  ( .A(\SUBBYTES[0].a/w2683 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n931 ) );
  XOR \SUBBYTES[0].a/U4766  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2668 ), .Z(\SUBBYTES[0].a/n932 ) );
  XOR \SUBBYTES[0].a/U4765  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n933 ), .Z(
        \SUBBYTES[0].a/n1533 ) );
  XOR \SUBBYTES[0].a/U4764  ( .A(\w1[0][35] ), .B(\w1[0][34] ), .Z(
        \SUBBYTES[0].a/n933 ) );
  XOR \SUBBYTES[0].a/U4763  ( .A(\w1[0][38] ), .B(\SUBBYTES[0].a/n1533 ), .Z(
        \SUBBYTES[0].a/w2550 ) );
  XOR \SUBBYTES[0].a/U4762  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/w2437 ) );
  XOR \SUBBYTES[0].a/U4761  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/n934 ), .Z(
        \SUBBYTES[0].a/w2438 ) );
  XOR \SUBBYTES[0].a/U4760  ( .A(\w1[0][38] ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n934 ) );
  XOR \SUBBYTES[0].a/U4759  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n1533 ), .Z(
        \SUBBYTES[0].a/w2568 ) );
  XOR \SUBBYTES[0].a/U4758  ( .A(\SUBBYTES[0].a/n936 ), .B(
        \SUBBYTES[0].a/n935 ), .Z(\SUBBYTES[0].a/w2561 ) );
  XOR \SUBBYTES[0].a/U4757  ( .A(\w1[0][35] ), .B(\w1[0][33] ), .Z(
        \SUBBYTES[0].a/n935 ) );
  XOR \SUBBYTES[0].a/U4756  ( .A(\w1[0][39] ), .B(\w1[0][36] ), .Z(
        \SUBBYTES[0].a/n936 ) );
  XOR \SUBBYTES[0].a/U4755  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2561 ), .Z(
        \SUBBYTES[0].a/w2440 ) );
  XOR \SUBBYTES[0].a/U4754  ( .A(\SUBBYTES[0].a/n938 ), .B(
        \SUBBYTES[0].a/n937 ), .Z(\SUBBYTES[0].a/w2548 ) );
  XOR \SUBBYTES[0].a/U4753  ( .A(\SUBBYTES[0].a/w2509 ), .B(n12), .Z(
        \SUBBYTES[0].a/n937 ) );
  XOR \SUBBYTES[0].a/U4752  ( .A(\SUBBYTES[0].a/w2502 ), .B(
        \SUBBYTES[0].a/w2505 ), .Z(\SUBBYTES[0].a/n938 ) );
  XOR \SUBBYTES[0].a/U4751  ( .A(\SUBBYTES[0].a/n940 ), .B(
        \SUBBYTES[0].a/n939 ), .Z(\SUBBYTES[0].a/w2549 ) );
  XOR \SUBBYTES[0].a/U4750  ( .A(\SUBBYTES[0].a/w2509 ), .B(
        \SUBBYTES[0].a/n120 ), .Z(\SUBBYTES[0].a/n939 ) );
  XOR \SUBBYTES[0].a/U4749  ( .A(\SUBBYTES[0].a/w2502 ), .B(
        \SUBBYTES[0].a/n119 ), .Z(\SUBBYTES[0].a/n940 ) );
  XOR \SUBBYTES[0].a/U4748  ( .A(\SUBBYTES[0].a/w2561 ), .B(
        \SUBBYTES[0].a/n941 ), .Z(\SUBBYTES[0].a/w2551 ) );
  XOR \SUBBYTES[0].a/U4747  ( .A(\w1[0][38] ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n941 ) );
  XOR \SUBBYTES[0].a/U4746  ( .A(\SUBBYTES[0].a/n943 ), .B(
        \SUBBYTES[0].a/n942 ), .Z(\SUBBYTES[0].a/w2552 ) );
  XOR \SUBBYTES[0].a/U4745  ( .A(\SUBBYTES[0].a/n120 ), .B(n12), .Z(
        \SUBBYTES[0].a/n942 ) );
  XOR \SUBBYTES[0].a/U4744  ( .A(\SUBBYTES[0].a/n119 ), .B(
        \SUBBYTES[0].a/w2505 ), .Z(\SUBBYTES[0].a/n943 ) );
  XOR \SUBBYTES[0].a/U4743  ( .A(\w1[0][39] ), .B(\w1[0][34] ), .Z(
        \SUBBYTES[0].a/n1539 ) );
  XOR \SUBBYTES[0].a/U4742  ( .A(\SUBBYTES[0].a/n1539 ), .B(
        \SUBBYTES[0].a/n944 ), .Z(\SUBBYTES[0].a/w2553 ) );
  XOR \SUBBYTES[0].a/U4741  ( .A(\w1[0][37] ), .B(\w1[0][36] ), .Z(
        \SUBBYTES[0].a/n944 ) );
  XOR \SUBBYTES[0].a/U4740  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2441 ) );
  XOR \SUBBYTES[0].a/U4739  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2442 ) );
  XOR \SUBBYTES[0].a/U4738  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2443 ) );
  XOR \SUBBYTES[0].a/U4737  ( .A(\SUBBYTES[0].a/w2442 ), .B(
        \SUBBYTES[0].a/n1539 ), .Z(\SUBBYTES[0].a/w2444 ) );
  XOR \SUBBYTES[0].a/U4736  ( .A(\SUBBYTES[0].a/n1539 ), .B(
        \SUBBYTES[0].a/n945 ), .Z(\SUBBYTES[0].a/w2529 ) );
  XOR \SUBBYTES[0].a/U4735  ( .A(\w1[0][36] ), .B(\w1[0][33] ), .Z(
        \SUBBYTES[0].a/n945 ) );
  XOR \SUBBYTES[0].a/U4734  ( .A(\SUBBYTES[0].a/n947 ), .B(
        \SUBBYTES[0].a/n946 ), .Z(\SUBBYTES[0].a/n1536 ) );
  XOR \SUBBYTES[0].a/U4733  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/n948 ), .Z(
        \SUBBYTES[0].a/n946 ) );
  XOR \SUBBYTES[0].a/U4732  ( .A(\SUBBYTES[0].a/w2494 ), .B(\w1[0][38] ), .Z(
        \SUBBYTES[0].a/n947 ) );
  XOR \SUBBYTES[0].a/U4731  ( .A(\SUBBYTES[0].a/w2468 ), .B(
        \SUBBYTES[0].a/w2475 ), .Z(\SUBBYTES[0].a/n948 ) );
  XOR \SUBBYTES[0].a/U4730  ( .A(\SUBBYTES[0].a/n950 ), .B(
        \SUBBYTES[0].a/n949 ), .Z(\SUBBYTES[0].a/n1534 ) );
  XOR \SUBBYTES[0].a/U4729  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n951 ), .Z(
        \SUBBYTES[0].a/n949 ) );
  XOR \SUBBYTES[0].a/U4728  ( .A(\SUBBYTES[0].a/w2493 ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n950 ) );
  XOR \SUBBYTES[0].a/U4727  ( .A(\SUBBYTES[0].a/w2469 ), .B(
        \SUBBYTES[0].a/w2476 ), .Z(\SUBBYTES[0].a/n951 ) );
  XOR \SUBBYTES[0].a/U4726  ( .A(\SUBBYTES[0].a/n1536 ), .B(
        \SUBBYTES[0].a/n1534 ), .Z(\SUBBYTES[0].a/w2499 ) );
  XOR \SUBBYTES[0].a/U4725  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n952 ), .Z(
        \SUBBYTES[0].a/n1537 ) );
  XOR \SUBBYTES[0].a/U4724  ( .A(\SUBBYTES[0].a/w2461 ), .B(
        \SUBBYTES[0].a/w2471 ), .Z(\SUBBYTES[0].a/n952 ) );
  XOR \SUBBYTES[0].a/U4723  ( .A(\SUBBYTES[0].a/n954 ), .B(
        \SUBBYTES[0].a/n953 ), .Z(\SUBBYTES[0].a/w2486 ) );
  XOR \SUBBYTES[0].a/U4722  ( .A(\SUBBYTES[0].a/n1537 ), .B(
        \SUBBYTES[0].a/n955 ), .Z(\SUBBYTES[0].a/n953 ) );
  XOR \SUBBYTES[0].a/U4721  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/n954 ) );
  XOR \SUBBYTES[0].a/U4720  ( .A(\SUBBYTES[0].a/w2463 ), .B(
        \SUBBYTES[0].a/w2468 ), .Z(\SUBBYTES[0].a/n955 ) );
  XOR \SUBBYTES[0].a/U4719  ( .A(\SUBBYTES[0].a/n957 ), .B(
        \SUBBYTES[0].a/n956 ), .Z(\SUBBYTES[0].a/n1535 ) );
  XOR \SUBBYTES[0].a/U4718  ( .A(\SUBBYTES[0].a/w2496 ), .B(\w1[0][39] ), .Z(
        \SUBBYTES[0].a/n956 ) );
  XOR \SUBBYTES[0].a/U4717  ( .A(\SUBBYTES[0].a/w2471 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n957 ) );
  XOR \SUBBYTES[0].a/U4716  ( .A(\SUBBYTES[0].a/n1534 ), .B(
        \SUBBYTES[0].a/n1535 ), .Z(\SUBBYTES[0].a/w2498 ) );
  XOR \SUBBYTES[0].a/U4715  ( .A(\w1[0][35] ), .B(\SUBBYTES[0].a/n958 ), .Z(
        \SUBBYTES[0].a/n1538 ) );
  XOR \SUBBYTES[0].a/U4714  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2463 ), .Z(\SUBBYTES[0].a/n958 ) );
  XOR \SUBBYTES[0].a/U4713  ( .A(\SUBBYTES[0].a/n960 ), .B(
        \SUBBYTES[0].a/n959 ), .Z(\SUBBYTES[0].a/w2487 ) );
  XOR \SUBBYTES[0].a/U4712  ( .A(\SUBBYTES[0].a/n1538 ), .B(
        \SUBBYTES[0].a/n961 ), .Z(\SUBBYTES[0].a/n959 ) );
  XOR \SUBBYTES[0].a/U4711  ( .A(\w1[0][38] ), .B(\SUBBYTES[0].a/w2529 ), .Z(
        \SUBBYTES[0].a/n960 ) );
  XOR \SUBBYTES[0].a/U4710  ( .A(\SUBBYTES[0].a/w2468 ), .B(
        \SUBBYTES[0].a/w2469 ), .Z(\SUBBYTES[0].a/n961 ) );
  XOR \SUBBYTES[0].a/U4709  ( .A(\SUBBYTES[0].a/n1536 ), .B(
        \SUBBYTES[0].a/n1535 ), .Z(\SUBBYTES[0].a/w2507 ) );
  XOR \SUBBYTES[0].a/U4708  ( .A(\SUBBYTES[0].a/n963 ), .B(
        \SUBBYTES[0].a/n962 ), .Z(\SUBBYTES[0].a/w2508 ) );
  XOR \SUBBYTES[0].a/U4707  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/n1537 ), .Z(
        \SUBBYTES[0].a/n962 ) );
  XOR \SUBBYTES[0].a/U4706  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2469 ), .Z(\SUBBYTES[0].a/n963 ) );
  XOR \SUBBYTES[0].a/U4705  ( .A(\SUBBYTES[0].a/n965 ), .B(
        \SUBBYTES[0].a/n964 ), .Z(\SUBBYTES[0].a/w2484 ) );
  XOR \SUBBYTES[0].a/U4704  ( .A(\SUBBYTES[0].a/n967 ), .B(
        \SUBBYTES[0].a/n966 ), .Z(\SUBBYTES[0].a/n964 ) );
  XOR \SUBBYTES[0].a/U4703  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/w2568 ), .Z(
        \SUBBYTES[0].a/n965 ) );
  XOR \SUBBYTES[0].a/U4702  ( .A(\SUBBYTES[0].a/w2475 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n966 ) );
  XOR \SUBBYTES[0].a/U4701  ( .A(\SUBBYTES[0].a/w2461 ), .B(
        \SUBBYTES[0].a/w2463 ), .Z(\SUBBYTES[0].a/n967 ) );
  XOR \SUBBYTES[0].a/U4700  ( .A(\SUBBYTES[0].a/n969 ), .B(
        \SUBBYTES[0].a/n968 ), .Z(\SUBBYTES[0].a/w2485 ) );
  XOR \SUBBYTES[0].a/U4699  ( .A(\SUBBYTES[0].a/n1538 ), .B(
        \SUBBYTES[0].a/n970 ), .Z(\SUBBYTES[0].a/n968 ) );
  XOR \SUBBYTES[0].a/U4698  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n1539 ), .Z(
        \SUBBYTES[0].a/n969 ) );
  XOR \SUBBYTES[0].a/U4697  ( .A(\SUBBYTES[0].a/w2475 ), .B(
        \SUBBYTES[0].a/w2476 ), .Z(\SUBBYTES[0].a/n970 ) );
  XOR \SUBBYTES[0].a/U4696  ( .A(\SUBBYTES[0].a/n972 ), .B(
        \SUBBYTES[0].a/n971 ), .Z(\SUBBYTES[0].a/w2501 ) );
  XOR \SUBBYTES[0].a/U4695  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n973 ), .Z(
        \SUBBYTES[0].a/n971 ) );
  XOR \SUBBYTES[0].a/U4694  ( .A(\SUBBYTES[0].a/w2476 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n972 ) );
  XOR \SUBBYTES[0].a/U4693  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2461 ), .Z(\SUBBYTES[0].a/n973 ) );
  XOR \SUBBYTES[0].a/U4692  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n974 ), .Z(
        \SUBBYTES[0].a/n1540 ) );
  XOR \SUBBYTES[0].a/U4691  ( .A(\w1[0][43] ), .B(\w1[0][42] ), .Z(
        \SUBBYTES[0].a/n974 ) );
  XOR \SUBBYTES[0].a/U4690  ( .A(\w1[0][46] ), .B(\SUBBYTES[0].a/n1540 ), .Z(
        \SUBBYTES[0].a/w2343 ) );
  XOR \SUBBYTES[0].a/U4689  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/w2230 ) );
  XOR \SUBBYTES[0].a/U4688  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/n975 ), .Z(
        \SUBBYTES[0].a/w2231 ) );
  XOR \SUBBYTES[0].a/U4687  ( .A(\w1[0][46] ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n975 ) );
  XOR \SUBBYTES[0].a/U4686  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n1540 ), .Z(
        \SUBBYTES[0].a/w2361 ) );
  XOR \SUBBYTES[0].a/U4685  ( .A(\SUBBYTES[0].a/n977 ), .B(
        \SUBBYTES[0].a/n976 ), .Z(\SUBBYTES[0].a/w2354 ) );
  XOR \SUBBYTES[0].a/U4684  ( .A(\w1[0][43] ), .B(\w1[0][41] ), .Z(
        \SUBBYTES[0].a/n976 ) );
  XOR \SUBBYTES[0].a/U4683  ( .A(\w1[0][47] ), .B(\w1[0][44] ), .Z(
        \SUBBYTES[0].a/n977 ) );
  XOR \SUBBYTES[0].a/U4682  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2354 ), .Z(
        \SUBBYTES[0].a/w2233 ) );
  XOR \SUBBYTES[0].a/U4681  ( .A(\SUBBYTES[0].a/n979 ), .B(
        \SUBBYTES[0].a/n978 ), .Z(\SUBBYTES[0].a/w2341 ) );
  XOR \SUBBYTES[0].a/U4680  ( .A(\SUBBYTES[0].a/w2302 ), .B(n11), .Z(
        \SUBBYTES[0].a/n978 ) );
  XOR \SUBBYTES[0].a/U4679  ( .A(\SUBBYTES[0].a/w2295 ), .B(
        \SUBBYTES[0].a/w2298 ), .Z(\SUBBYTES[0].a/n979 ) );
  XOR \SUBBYTES[0].a/U4678  ( .A(\SUBBYTES[0].a/n981 ), .B(
        \SUBBYTES[0].a/n980 ), .Z(\SUBBYTES[0].a/w2342 ) );
  XOR \SUBBYTES[0].a/U4677  ( .A(\SUBBYTES[0].a/w2302 ), .B(
        \SUBBYTES[0].a/n110 ), .Z(\SUBBYTES[0].a/n980 ) );
  XOR \SUBBYTES[0].a/U4676  ( .A(\SUBBYTES[0].a/w2295 ), .B(
        \SUBBYTES[0].a/n109 ), .Z(\SUBBYTES[0].a/n981 ) );
  XOR \SUBBYTES[0].a/U4675  ( .A(\SUBBYTES[0].a/w2354 ), .B(
        \SUBBYTES[0].a/n982 ), .Z(\SUBBYTES[0].a/w2344 ) );
  XOR \SUBBYTES[0].a/U4674  ( .A(\w1[0][46] ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n982 ) );
  XOR \SUBBYTES[0].a/U4673  ( .A(\SUBBYTES[0].a/n984 ), .B(
        \SUBBYTES[0].a/n983 ), .Z(\SUBBYTES[0].a/w2345 ) );
  XOR \SUBBYTES[0].a/U4672  ( .A(\SUBBYTES[0].a/n110 ), .B(n11), .Z(
        \SUBBYTES[0].a/n983 ) );
  XOR \SUBBYTES[0].a/U4671  ( .A(\SUBBYTES[0].a/n109 ), .B(
        \SUBBYTES[0].a/w2298 ), .Z(\SUBBYTES[0].a/n984 ) );
  XOR \SUBBYTES[0].a/U4670  ( .A(\w1[0][47] ), .B(\w1[0][42] ), .Z(
        \SUBBYTES[0].a/n1546 ) );
  XOR \SUBBYTES[0].a/U4669  ( .A(\SUBBYTES[0].a/n1546 ), .B(
        \SUBBYTES[0].a/n985 ), .Z(\SUBBYTES[0].a/w2346 ) );
  XOR \SUBBYTES[0].a/U4668  ( .A(\w1[0][45] ), .B(\w1[0][44] ), .Z(
        \SUBBYTES[0].a/n985 ) );
  XOR \SUBBYTES[0].a/U4667  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2234 ) );
  XOR \SUBBYTES[0].a/U4666  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2235 ) );
  XOR \SUBBYTES[0].a/U4665  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2236 ) );
  XOR \SUBBYTES[0].a/U4664  ( .A(\SUBBYTES[0].a/w2235 ), .B(
        \SUBBYTES[0].a/n1546 ), .Z(\SUBBYTES[0].a/w2237 ) );
  XOR \SUBBYTES[0].a/U4663  ( .A(\SUBBYTES[0].a/n1546 ), .B(
        \SUBBYTES[0].a/n986 ), .Z(\SUBBYTES[0].a/w2322 ) );
  XOR \SUBBYTES[0].a/U4662  ( .A(\w1[0][44] ), .B(\w1[0][41] ), .Z(
        \SUBBYTES[0].a/n986 ) );
  XOR \SUBBYTES[0].a/U4661  ( .A(\SUBBYTES[0].a/n988 ), .B(
        \SUBBYTES[0].a/n987 ), .Z(\SUBBYTES[0].a/n1543 ) );
  XOR \SUBBYTES[0].a/U4660  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/n989 ), .Z(
        \SUBBYTES[0].a/n987 ) );
  XOR \SUBBYTES[0].a/U4659  ( .A(\SUBBYTES[0].a/w2287 ), .B(\w1[0][46] ), .Z(
        \SUBBYTES[0].a/n988 ) );
  XOR \SUBBYTES[0].a/U4658  ( .A(\SUBBYTES[0].a/w2261 ), .B(
        \SUBBYTES[0].a/w2268 ), .Z(\SUBBYTES[0].a/n989 ) );
  XOR \SUBBYTES[0].a/U4657  ( .A(\SUBBYTES[0].a/n991 ), .B(
        \SUBBYTES[0].a/n990 ), .Z(\SUBBYTES[0].a/n1541 ) );
  XOR \SUBBYTES[0].a/U4656  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n992 ), .Z(
        \SUBBYTES[0].a/n990 ) );
  XOR \SUBBYTES[0].a/U4655  ( .A(\SUBBYTES[0].a/w2286 ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n991 ) );
  XOR \SUBBYTES[0].a/U4654  ( .A(\SUBBYTES[0].a/w2262 ), .B(
        \SUBBYTES[0].a/w2269 ), .Z(\SUBBYTES[0].a/n992 ) );
  XOR \SUBBYTES[0].a/U4653  ( .A(\SUBBYTES[0].a/n1543 ), .B(
        \SUBBYTES[0].a/n1541 ), .Z(\SUBBYTES[0].a/w2292 ) );
  XOR \SUBBYTES[0].a/U4652  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n993 ), .Z(
        \SUBBYTES[0].a/n1544 ) );
  XOR \SUBBYTES[0].a/U4651  ( .A(\SUBBYTES[0].a/w2254 ), .B(
        \SUBBYTES[0].a/w2264 ), .Z(\SUBBYTES[0].a/n993 ) );
  XOR \SUBBYTES[0].a/U4650  ( .A(\SUBBYTES[0].a/n995 ), .B(
        \SUBBYTES[0].a/n994 ), .Z(\SUBBYTES[0].a/w2279 ) );
  XOR \SUBBYTES[0].a/U4649  ( .A(\SUBBYTES[0].a/n1544 ), .B(
        \SUBBYTES[0].a/n996 ), .Z(\SUBBYTES[0].a/n994 ) );
  XOR \SUBBYTES[0].a/U4648  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/n995 ) );
  XOR \SUBBYTES[0].a/U4647  ( .A(\SUBBYTES[0].a/w2256 ), .B(
        \SUBBYTES[0].a/w2261 ), .Z(\SUBBYTES[0].a/n996 ) );
  XOR \SUBBYTES[0].a/U4646  ( .A(\SUBBYTES[0].a/n998 ), .B(
        \SUBBYTES[0].a/n997 ), .Z(\SUBBYTES[0].a/n1542 ) );
  XOR \SUBBYTES[0].a/U4645  ( .A(\SUBBYTES[0].a/w2289 ), .B(\w1[0][47] ), .Z(
        \SUBBYTES[0].a/n997 ) );
  XOR \SUBBYTES[0].a/U4644  ( .A(\SUBBYTES[0].a/w2264 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n998 ) );
  XOR \SUBBYTES[0].a/U4643  ( .A(\SUBBYTES[0].a/n1541 ), .B(
        \SUBBYTES[0].a/n1542 ), .Z(\SUBBYTES[0].a/w2291 ) );
  XOR \SUBBYTES[0].a/U4642  ( .A(\w1[0][43] ), .B(\SUBBYTES[0].a/n999 ), .Z(
        \SUBBYTES[0].a/n1545 ) );
  XOR \SUBBYTES[0].a/U4641  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2256 ), .Z(\SUBBYTES[0].a/n999 ) );
  XOR \SUBBYTES[0].a/U4640  ( .A(\SUBBYTES[0].a/n1001 ), .B(
        \SUBBYTES[0].a/n1000 ), .Z(\SUBBYTES[0].a/w2280 ) );
  XOR \SUBBYTES[0].a/U4639  ( .A(\SUBBYTES[0].a/n1545 ), .B(
        \SUBBYTES[0].a/n1002 ), .Z(\SUBBYTES[0].a/n1000 ) );
  XOR \SUBBYTES[0].a/U4638  ( .A(\w1[0][46] ), .B(\SUBBYTES[0].a/w2322 ), .Z(
        \SUBBYTES[0].a/n1001 ) );
  XOR \SUBBYTES[0].a/U4637  ( .A(\SUBBYTES[0].a/w2261 ), .B(
        \SUBBYTES[0].a/w2262 ), .Z(\SUBBYTES[0].a/n1002 ) );
  XOR \SUBBYTES[0].a/U4636  ( .A(\SUBBYTES[0].a/n1543 ), .B(
        \SUBBYTES[0].a/n1542 ), .Z(\SUBBYTES[0].a/w2300 ) );
  XOR \SUBBYTES[0].a/U4635  ( .A(\SUBBYTES[0].a/n1004 ), .B(
        \SUBBYTES[0].a/n1003 ), .Z(\SUBBYTES[0].a/w2301 ) );
  XOR \SUBBYTES[0].a/U4634  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/n1544 ), .Z(
        \SUBBYTES[0].a/n1003 ) );
  XOR \SUBBYTES[0].a/U4633  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2262 ), .Z(\SUBBYTES[0].a/n1004 ) );
  XOR \SUBBYTES[0].a/U4632  ( .A(\SUBBYTES[0].a/n1006 ), .B(
        \SUBBYTES[0].a/n1005 ), .Z(\SUBBYTES[0].a/w2277 ) );
  XOR \SUBBYTES[0].a/U4631  ( .A(\SUBBYTES[0].a/n1008 ), .B(
        \SUBBYTES[0].a/n1007 ), .Z(\SUBBYTES[0].a/n1005 ) );
  XOR \SUBBYTES[0].a/U4630  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/w2361 ), .Z(
        \SUBBYTES[0].a/n1006 ) );
  XOR \SUBBYTES[0].a/U4629  ( .A(\SUBBYTES[0].a/w2268 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n1007 ) );
  XOR \SUBBYTES[0].a/U4628  ( .A(\SUBBYTES[0].a/w2254 ), .B(
        \SUBBYTES[0].a/w2256 ), .Z(\SUBBYTES[0].a/n1008 ) );
  XOR \SUBBYTES[0].a/U4627  ( .A(\SUBBYTES[0].a/n1010 ), .B(
        \SUBBYTES[0].a/n1009 ), .Z(\SUBBYTES[0].a/w2278 ) );
  XOR \SUBBYTES[0].a/U4626  ( .A(\SUBBYTES[0].a/n1545 ), .B(
        \SUBBYTES[0].a/n1011 ), .Z(\SUBBYTES[0].a/n1009 ) );
  XOR \SUBBYTES[0].a/U4625  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n1546 ), .Z(
        \SUBBYTES[0].a/n1010 ) );
  XOR \SUBBYTES[0].a/U4624  ( .A(\SUBBYTES[0].a/w2268 ), .B(
        \SUBBYTES[0].a/w2269 ), .Z(\SUBBYTES[0].a/n1011 ) );
  XOR \SUBBYTES[0].a/U4623  ( .A(\SUBBYTES[0].a/n1013 ), .B(
        \SUBBYTES[0].a/n1012 ), .Z(\SUBBYTES[0].a/w2294 ) );
  XOR \SUBBYTES[0].a/U4622  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n1014 ), .Z(
        \SUBBYTES[0].a/n1012 ) );
  XOR \SUBBYTES[0].a/U4621  ( .A(\SUBBYTES[0].a/w2269 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n1013 ) );
  XOR \SUBBYTES[0].a/U4620  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2254 ), .Z(\SUBBYTES[0].a/n1014 ) );
  XOR \SUBBYTES[0].a/U4619  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1015 ), .Z(
        \SUBBYTES[0].a/n1547 ) );
  XOR \SUBBYTES[0].a/U4618  ( .A(\w1[0][51] ), .B(\w1[0][50] ), .Z(
        \SUBBYTES[0].a/n1015 ) );
  XOR \SUBBYTES[0].a/U4617  ( .A(\w1[0][54] ), .B(\SUBBYTES[0].a/n1547 ), .Z(
        \SUBBYTES[0].a/w2136 ) );
  XOR \SUBBYTES[0].a/U4616  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/w2023 ) );
  XOR \SUBBYTES[0].a/U4615  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/n1016 ), .Z(
        \SUBBYTES[0].a/w2024 ) );
  XOR \SUBBYTES[0].a/U4614  ( .A(\w1[0][54] ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1016 ) );
  XOR \SUBBYTES[0].a/U4613  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1547 ), .Z(
        \SUBBYTES[0].a/w2154 ) );
  XOR \SUBBYTES[0].a/U4612  ( .A(\SUBBYTES[0].a/n1018 ), .B(
        \SUBBYTES[0].a/n1017 ), .Z(\SUBBYTES[0].a/w2147 ) );
  XOR \SUBBYTES[0].a/U4611  ( .A(\w1[0][51] ), .B(\w1[0][49] ), .Z(
        \SUBBYTES[0].a/n1017 ) );
  XOR \SUBBYTES[0].a/U4610  ( .A(\w1[0][55] ), .B(\w1[0][52] ), .Z(
        \SUBBYTES[0].a/n1018 ) );
  XOR \SUBBYTES[0].a/U4609  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2147 ), .Z(
        \SUBBYTES[0].a/w2026 ) );
  XOR \SUBBYTES[0].a/U4608  ( .A(\SUBBYTES[0].a/n1020 ), .B(
        \SUBBYTES[0].a/n1019 ), .Z(\SUBBYTES[0].a/w2134 ) );
  XOR \SUBBYTES[0].a/U4607  ( .A(\SUBBYTES[0].a/w2095 ), .B(n10), .Z(
        \SUBBYTES[0].a/n1019 ) );
  XOR \SUBBYTES[0].a/U4606  ( .A(\SUBBYTES[0].a/w2088 ), .B(
        \SUBBYTES[0].a/w2091 ), .Z(\SUBBYTES[0].a/n1020 ) );
  XOR \SUBBYTES[0].a/U4605  ( .A(\SUBBYTES[0].a/n1022 ), .B(
        \SUBBYTES[0].a/n1021 ), .Z(\SUBBYTES[0].a/w2135 ) );
  XOR \SUBBYTES[0].a/U4604  ( .A(\SUBBYTES[0].a/w2095 ), .B(
        \SUBBYTES[0].a/n100 ), .Z(\SUBBYTES[0].a/n1021 ) );
  XOR \SUBBYTES[0].a/U4603  ( .A(\SUBBYTES[0].a/w2088 ), .B(
        \SUBBYTES[0].a/n99 ), .Z(\SUBBYTES[0].a/n1022 ) );
  XOR \SUBBYTES[0].a/U4602  ( .A(\SUBBYTES[0].a/w2147 ), .B(
        \SUBBYTES[0].a/n1023 ), .Z(\SUBBYTES[0].a/w2137 ) );
  XOR \SUBBYTES[0].a/U4601  ( .A(\w1[0][54] ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1023 ) );
  XOR \SUBBYTES[0].a/U4600  ( .A(\SUBBYTES[0].a/n1025 ), .B(
        \SUBBYTES[0].a/n1024 ), .Z(\SUBBYTES[0].a/w2138 ) );
  XOR \SUBBYTES[0].a/U4599  ( .A(\SUBBYTES[0].a/n100 ), .B(n10), .Z(
        \SUBBYTES[0].a/n1024 ) );
  XOR \SUBBYTES[0].a/U4598  ( .A(\SUBBYTES[0].a/n99 ), .B(
        \SUBBYTES[0].a/w2091 ), .Z(\SUBBYTES[0].a/n1025 ) );
  XOR \SUBBYTES[0].a/U4597  ( .A(\w1[0][55] ), .B(\w1[0][50] ), .Z(
        \SUBBYTES[0].a/n1553 ) );
  XOR \SUBBYTES[0].a/U4596  ( .A(\SUBBYTES[0].a/n1553 ), .B(
        \SUBBYTES[0].a/n1026 ), .Z(\SUBBYTES[0].a/w2139 ) );
  XOR \SUBBYTES[0].a/U4595  ( .A(\w1[0][53] ), .B(\w1[0][52] ), .Z(
        \SUBBYTES[0].a/n1026 ) );
  XOR \SUBBYTES[0].a/U4594  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2027 ) );
  XOR \SUBBYTES[0].a/U4593  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2028 ) );
  XOR \SUBBYTES[0].a/U4592  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2029 ) );
  XOR \SUBBYTES[0].a/U4591  ( .A(\SUBBYTES[0].a/w2028 ), .B(
        \SUBBYTES[0].a/n1553 ), .Z(\SUBBYTES[0].a/w2030 ) );
  XOR \SUBBYTES[0].a/U4590  ( .A(\SUBBYTES[0].a/n1553 ), .B(
        \SUBBYTES[0].a/n1027 ), .Z(\SUBBYTES[0].a/w2115 ) );
  XOR \SUBBYTES[0].a/U4589  ( .A(\w1[0][52] ), .B(\w1[0][49] ), .Z(
        \SUBBYTES[0].a/n1027 ) );
  XOR \SUBBYTES[0].a/U4588  ( .A(\SUBBYTES[0].a/n1029 ), .B(
        \SUBBYTES[0].a/n1028 ), .Z(\SUBBYTES[0].a/n1550 ) );
  XOR \SUBBYTES[0].a/U4587  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/n1030 ), .Z(
        \SUBBYTES[0].a/n1028 ) );
  XOR \SUBBYTES[0].a/U4586  ( .A(\SUBBYTES[0].a/w2080 ), .B(\w1[0][54] ), .Z(
        \SUBBYTES[0].a/n1029 ) );
  XOR \SUBBYTES[0].a/U4585  ( .A(\SUBBYTES[0].a/w2054 ), .B(
        \SUBBYTES[0].a/w2061 ), .Z(\SUBBYTES[0].a/n1030 ) );
  XOR \SUBBYTES[0].a/U4584  ( .A(\SUBBYTES[0].a/n1032 ), .B(
        \SUBBYTES[0].a/n1031 ), .Z(\SUBBYTES[0].a/n1548 ) );
  XOR \SUBBYTES[0].a/U4583  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1033 ), .Z(
        \SUBBYTES[0].a/n1031 ) );
  XOR \SUBBYTES[0].a/U4582  ( .A(\SUBBYTES[0].a/w2079 ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1032 ) );
  XOR \SUBBYTES[0].a/U4581  ( .A(\SUBBYTES[0].a/w2055 ), .B(
        \SUBBYTES[0].a/w2062 ), .Z(\SUBBYTES[0].a/n1033 ) );
  XOR \SUBBYTES[0].a/U4580  ( .A(\SUBBYTES[0].a/n1550 ), .B(
        \SUBBYTES[0].a/n1548 ), .Z(\SUBBYTES[0].a/w2085 ) );
  XOR \SUBBYTES[0].a/U4579  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1034 ), .Z(
        \SUBBYTES[0].a/n1551 ) );
  XOR \SUBBYTES[0].a/U4578  ( .A(\SUBBYTES[0].a/w2047 ), .B(
        \SUBBYTES[0].a/w2057 ), .Z(\SUBBYTES[0].a/n1034 ) );
  XOR \SUBBYTES[0].a/U4577  ( .A(\SUBBYTES[0].a/n1036 ), .B(
        \SUBBYTES[0].a/n1035 ), .Z(\SUBBYTES[0].a/w2072 ) );
  XOR \SUBBYTES[0].a/U4576  ( .A(\SUBBYTES[0].a/n1551 ), .B(
        \SUBBYTES[0].a/n1037 ), .Z(\SUBBYTES[0].a/n1035 ) );
  XOR \SUBBYTES[0].a/U4575  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/n1036 ) );
  XOR \SUBBYTES[0].a/U4574  ( .A(\SUBBYTES[0].a/w2049 ), .B(
        \SUBBYTES[0].a/w2054 ), .Z(\SUBBYTES[0].a/n1037 ) );
  XOR \SUBBYTES[0].a/U4573  ( .A(\SUBBYTES[0].a/n1039 ), .B(
        \SUBBYTES[0].a/n1038 ), .Z(\SUBBYTES[0].a/n1549 ) );
  XOR \SUBBYTES[0].a/U4572  ( .A(\SUBBYTES[0].a/w2082 ), .B(\w1[0][55] ), .Z(
        \SUBBYTES[0].a/n1038 ) );
  XOR \SUBBYTES[0].a/U4571  ( .A(\SUBBYTES[0].a/w2057 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1039 ) );
  XOR \SUBBYTES[0].a/U4570  ( .A(\SUBBYTES[0].a/n1548 ), .B(
        \SUBBYTES[0].a/n1549 ), .Z(\SUBBYTES[0].a/w2084 ) );
  XOR \SUBBYTES[0].a/U4569  ( .A(\w1[0][51] ), .B(\SUBBYTES[0].a/n1040 ), .Z(
        \SUBBYTES[0].a/n1552 ) );
  XOR \SUBBYTES[0].a/U4568  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2049 ), .Z(\SUBBYTES[0].a/n1040 ) );
  XOR \SUBBYTES[0].a/U4567  ( .A(\SUBBYTES[0].a/n1042 ), .B(
        \SUBBYTES[0].a/n1041 ), .Z(\SUBBYTES[0].a/w2073 ) );
  XOR \SUBBYTES[0].a/U4566  ( .A(\SUBBYTES[0].a/n1552 ), .B(
        \SUBBYTES[0].a/n1043 ), .Z(\SUBBYTES[0].a/n1041 ) );
  XOR \SUBBYTES[0].a/U4565  ( .A(\w1[0][54] ), .B(\SUBBYTES[0].a/w2115 ), .Z(
        \SUBBYTES[0].a/n1042 ) );
  XOR \SUBBYTES[0].a/U4564  ( .A(\SUBBYTES[0].a/w2054 ), .B(
        \SUBBYTES[0].a/w2055 ), .Z(\SUBBYTES[0].a/n1043 ) );
  XOR \SUBBYTES[0].a/U4563  ( .A(\SUBBYTES[0].a/n1550 ), .B(
        \SUBBYTES[0].a/n1549 ), .Z(\SUBBYTES[0].a/w2093 ) );
  XOR \SUBBYTES[0].a/U4562  ( .A(\SUBBYTES[0].a/n1045 ), .B(
        \SUBBYTES[0].a/n1044 ), .Z(\SUBBYTES[0].a/w2094 ) );
  XOR \SUBBYTES[0].a/U4561  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/n1551 ), .Z(
        \SUBBYTES[0].a/n1044 ) );
  XOR \SUBBYTES[0].a/U4560  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2055 ), .Z(\SUBBYTES[0].a/n1045 ) );
  XOR \SUBBYTES[0].a/U4559  ( .A(\SUBBYTES[0].a/n1047 ), .B(
        \SUBBYTES[0].a/n1046 ), .Z(\SUBBYTES[0].a/w2070 ) );
  XOR \SUBBYTES[0].a/U4558  ( .A(\SUBBYTES[0].a/n1049 ), .B(
        \SUBBYTES[0].a/n1048 ), .Z(\SUBBYTES[0].a/n1046 ) );
  XOR \SUBBYTES[0].a/U4557  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/w2154 ), .Z(
        \SUBBYTES[0].a/n1047 ) );
  XOR \SUBBYTES[0].a/U4556  ( .A(\SUBBYTES[0].a/w2061 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1048 ) );
  XOR \SUBBYTES[0].a/U4555  ( .A(\SUBBYTES[0].a/w2047 ), .B(
        \SUBBYTES[0].a/w2049 ), .Z(\SUBBYTES[0].a/n1049 ) );
  XOR \SUBBYTES[0].a/U4554  ( .A(\SUBBYTES[0].a/n1051 ), .B(
        \SUBBYTES[0].a/n1050 ), .Z(\SUBBYTES[0].a/w2071 ) );
  XOR \SUBBYTES[0].a/U4553  ( .A(\SUBBYTES[0].a/n1552 ), .B(
        \SUBBYTES[0].a/n1052 ), .Z(\SUBBYTES[0].a/n1050 ) );
  XOR \SUBBYTES[0].a/U4552  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1553 ), .Z(
        \SUBBYTES[0].a/n1051 ) );
  XOR \SUBBYTES[0].a/U4551  ( .A(\SUBBYTES[0].a/w2061 ), .B(
        \SUBBYTES[0].a/w2062 ), .Z(\SUBBYTES[0].a/n1052 ) );
  XOR \SUBBYTES[0].a/U4550  ( .A(\SUBBYTES[0].a/n1054 ), .B(
        \SUBBYTES[0].a/n1053 ), .Z(\SUBBYTES[0].a/w2087 ) );
  XOR \SUBBYTES[0].a/U4549  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1055 ), .Z(
        \SUBBYTES[0].a/n1053 ) );
  XOR \SUBBYTES[0].a/U4548  ( .A(\SUBBYTES[0].a/w2062 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1054 ) );
  XOR \SUBBYTES[0].a/U4547  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2047 ), .Z(\SUBBYTES[0].a/n1055 ) );
  XOR \SUBBYTES[0].a/U4546  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1056 ), .Z(
        \SUBBYTES[0].a/n1554 ) );
  XOR \SUBBYTES[0].a/U4545  ( .A(\w1[0][59] ), .B(\w1[0][58] ), .Z(
        \SUBBYTES[0].a/n1056 ) );
  XOR \SUBBYTES[0].a/U4544  ( .A(\w1[0][62] ), .B(\SUBBYTES[0].a/n1554 ), .Z(
        \SUBBYTES[0].a/w1929 ) );
  XOR \SUBBYTES[0].a/U4543  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/w1816 ) );
  XOR \SUBBYTES[0].a/U4542  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/n1057 ), .Z(
        \SUBBYTES[0].a/w1817 ) );
  XOR \SUBBYTES[0].a/U4541  ( .A(\w1[0][62] ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1057 ) );
  XOR \SUBBYTES[0].a/U4540  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1554 ), .Z(
        \SUBBYTES[0].a/w1947 ) );
  XOR \SUBBYTES[0].a/U4539  ( .A(\SUBBYTES[0].a/n1059 ), .B(
        \SUBBYTES[0].a/n1058 ), .Z(\SUBBYTES[0].a/w1940 ) );
  XOR \SUBBYTES[0].a/U4538  ( .A(\w1[0][59] ), .B(\w1[0][57] ), .Z(
        \SUBBYTES[0].a/n1058 ) );
  XOR \SUBBYTES[0].a/U4537  ( .A(\w1[0][63] ), .B(\w1[0][60] ), .Z(
        \SUBBYTES[0].a/n1059 ) );
  XOR \SUBBYTES[0].a/U4536  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1940 ), .Z(
        \SUBBYTES[0].a/w1819 ) );
  XOR \SUBBYTES[0].a/U4535  ( .A(\SUBBYTES[0].a/n1061 ), .B(
        \SUBBYTES[0].a/n1060 ), .Z(\SUBBYTES[0].a/w1927 ) );
  XOR \SUBBYTES[0].a/U4534  ( .A(\SUBBYTES[0].a/w1888 ), .B(n9), .Z(
        \SUBBYTES[0].a/n1060 ) );
  XOR \SUBBYTES[0].a/U4533  ( .A(\SUBBYTES[0].a/w1881 ), .B(
        \SUBBYTES[0].a/w1884 ), .Z(\SUBBYTES[0].a/n1061 ) );
  XOR \SUBBYTES[0].a/U4532  ( .A(\SUBBYTES[0].a/n1063 ), .B(
        \SUBBYTES[0].a/n1062 ), .Z(\SUBBYTES[0].a/w1928 ) );
  XOR \SUBBYTES[0].a/U4531  ( .A(\SUBBYTES[0].a/w1888 ), .B(
        \SUBBYTES[0].a/n90 ), .Z(\SUBBYTES[0].a/n1062 ) );
  XOR \SUBBYTES[0].a/U4530  ( .A(\SUBBYTES[0].a/w1881 ), .B(
        \SUBBYTES[0].a/n89 ), .Z(\SUBBYTES[0].a/n1063 ) );
  XOR \SUBBYTES[0].a/U4529  ( .A(\SUBBYTES[0].a/w1940 ), .B(
        \SUBBYTES[0].a/n1064 ), .Z(\SUBBYTES[0].a/w1930 ) );
  XOR \SUBBYTES[0].a/U4528  ( .A(\w1[0][62] ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1064 ) );
  XOR \SUBBYTES[0].a/U4527  ( .A(\SUBBYTES[0].a/n1066 ), .B(
        \SUBBYTES[0].a/n1065 ), .Z(\SUBBYTES[0].a/w1931 ) );
  XOR \SUBBYTES[0].a/U4526  ( .A(\SUBBYTES[0].a/n90 ), .B(n9), .Z(
        \SUBBYTES[0].a/n1065 ) );
  XOR \SUBBYTES[0].a/U4525  ( .A(\SUBBYTES[0].a/n89 ), .B(
        \SUBBYTES[0].a/w1884 ), .Z(\SUBBYTES[0].a/n1066 ) );
  XOR \SUBBYTES[0].a/U4524  ( .A(\w1[0][63] ), .B(\w1[0][58] ), .Z(
        \SUBBYTES[0].a/n1560 ) );
  XOR \SUBBYTES[0].a/U4523  ( .A(\SUBBYTES[0].a/n1560 ), .B(
        \SUBBYTES[0].a/n1067 ), .Z(\SUBBYTES[0].a/w1932 ) );
  XOR \SUBBYTES[0].a/U4522  ( .A(\w1[0][61] ), .B(\w1[0][60] ), .Z(
        \SUBBYTES[0].a/n1067 ) );
  XOR \SUBBYTES[0].a/U4521  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1820 ) );
  XOR \SUBBYTES[0].a/U4520  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1821 ) );
  XOR \SUBBYTES[0].a/U4519  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1822 ) );
  XOR \SUBBYTES[0].a/U4518  ( .A(\SUBBYTES[0].a/w1821 ), .B(
        \SUBBYTES[0].a/n1560 ), .Z(\SUBBYTES[0].a/w1823 ) );
  XOR \SUBBYTES[0].a/U4517  ( .A(\SUBBYTES[0].a/n1560 ), .B(
        \SUBBYTES[0].a/n1068 ), .Z(\SUBBYTES[0].a/w1908 ) );
  XOR \SUBBYTES[0].a/U4516  ( .A(\w1[0][60] ), .B(\w1[0][57] ), .Z(
        \SUBBYTES[0].a/n1068 ) );
  XOR \SUBBYTES[0].a/U4515  ( .A(\SUBBYTES[0].a/n1070 ), .B(
        \SUBBYTES[0].a/n1069 ), .Z(\SUBBYTES[0].a/n1557 ) );
  XOR \SUBBYTES[0].a/U4514  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/n1071 ), .Z(
        \SUBBYTES[0].a/n1069 ) );
  XOR \SUBBYTES[0].a/U4513  ( .A(\SUBBYTES[0].a/w1873 ), .B(\w1[0][62] ), .Z(
        \SUBBYTES[0].a/n1070 ) );
  XOR \SUBBYTES[0].a/U4512  ( .A(\SUBBYTES[0].a/w1847 ), .B(
        \SUBBYTES[0].a/w1854 ), .Z(\SUBBYTES[0].a/n1071 ) );
  XOR \SUBBYTES[0].a/U4511  ( .A(\SUBBYTES[0].a/n1073 ), .B(
        \SUBBYTES[0].a/n1072 ), .Z(\SUBBYTES[0].a/n1555 ) );
  XOR \SUBBYTES[0].a/U4510  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1074 ), .Z(
        \SUBBYTES[0].a/n1072 ) );
  XOR \SUBBYTES[0].a/U4509  ( .A(\SUBBYTES[0].a/w1872 ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1073 ) );
  XOR \SUBBYTES[0].a/U4508  ( .A(\SUBBYTES[0].a/w1848 ), .B(
        \SUBBYTES[0].a/w1855 ), .Z(\SUBBYTES[0].a/n1074 ) );
  XOR \SUBBYTES[0].a/U4507  ( .A(\SUBBYTES[0].a/n1557 ), .B(
        \SUBBYTES[0].a/n1555 ), .Z(\SUBBYTES[0].a/w1878 ) );
  XOR \SUBBYTES[0].a/U4506  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1075 ), .Z(
        \SUBBYTES[0].a/n1558 ) );
  XOR \SUBBYTES[0].a/U4505  ( .A(\SUBBYTES[0].a/w1840 ), .B(
        \SUBBYTES[0].a/w1850 ), .Z(\SUBBYTES[0].a/n1075 ) );
  XOR \SUBBYTES[0].a/U4504  ( .A(\SUBBYTES[0].a/n1077 ), .B(
        \SUBBYTES[0].a/n1076 ), .Z(\SUBBYTES[0].a/w1865 ) );
  XOR \SUBBYTES[0].a/U4503  ( .A(\SUBBYTES[0].a/n1558 ), .B(
        \SUBBYTES[0].a/n1078 ), .Z(\SUBBYTES[0].a/n1076 ) );
  XOR \SUBBYTES[0].a/U4502  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/n1077 ) );
  XOR \SUBBYTES[0].a/U4501  ( .A(\SUBBYTES[0].a/w1842 ), .B(
        \SUBBYTES[0].a/w1847 ), .Z(\SUBBYTES[0].a/n1078 ) );
  XOR \SUBBYTES[0].a/U4500  ( .A(\SUBBYTES[0].a/n1080 ), .B(
        \SUBBYTES[0].a/n1079 ), .Z(\SUBBYTES[0].a/n1556 ) );
  XOR \SUBBYTES[0].a/U4499  ( .A(\SUBBYTES[0].a/w1875 ), .B(\w1[0][63] ), .Z(
        \SUBBYTES[0].a/n1079 ) );
  XOR \SUBBYTES[0].a/U4498  ( .A(\SUBBYTES[0].a/w1850 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1080 ) );
  XOR \SUBBYTES[0].a/U4497  ( .A(\SUBBYTES[0].a/n1555 ), .B(
        \SUBBYTES[0].a/n1556 ), .Z(\SUBBYTES[0].a/w1877 ) );
  XOR \SUBBYTES[0].a/U4496  ( .A(\w1[0][59] ), .B(\SUBBYTES[0].a/n1081 ), .Z(
        \SUBBYTES[0].a/n1559 ) );
  XOR \SUBBYTES[0].a/U4495  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1842 ), .Z(\SUBBYTES[0].a/n1081 ) );
  XOR \SUBBYTES[0].a/U4494  ( .A(\SUBBYTES[0].a/n1083 ), .B(
        \SUBBYTES[0].a/n1082 ), .Z(\SUBBYTES[0].a/w1866 ) );
  XOR \SUBBYTES[0].a/U4493  ( .A(\SUBBYTES[0].a/n1559 ), .B(
        \SUBBYTES[0].a/n1084 ), .Z(\SUBBYTES[0].a/n1082 ) );
  XOR \SUBBYTES[0].a/U4492  ( .A(\w1[0][62] ), .B(\SUBBYTES[0].a/w1908 ), .Z(
        \SUBBYTES[0].a/n1083 ) );
  XOR \SUBBYTES[0].a/U4491  ( .A(\SUBBYTES[0].a/w1847 ), .B(
        \SUBBYTES[0].a/w1848 ), .Z(\SUBBYTES[0].a/n1084 ) );
  XOR \SUBBYTES[0].a/U4490  ( .A(\SUBBYTES[0].a/n1557 ), .B(
        \SUBBYTES[0].a/n1556 ), .Z(\SUBBYTES[0].a/w1886 ) );
  XOR \SUBBYTES[0].a/U4489  ( .A(\SUBBYTES[0].a/n1086 ), .B(
        \SUBBYTES[0].a/n1085 ), .Z(\SUBBYTES[0].a/w1887 ) );
  XOR \SUBBYTES[0].a/U4488  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/n1558 ), .Z(
        \SUBBYTES[0].a/n1085 ) );
  XOR \SUBBYTES[0].a/U4487  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1848 ), .Z(\SUBBYTES[0].a/n1086 ) );
  XOR \SUBBYTES[0].a/U4486  ( .A(\SUBBYTES[0].a/n1088 ), .B(
        \SUBBYTES[0].a/n1087 ), .Z(\SUBBYTES[0].a/w1863 ) );
  XOR \SUBBYTES[0].a/U4485  ( .A(\SUBBYTES[0].a/n1090 ), .B(
        \SUBBYTES[0].a/n1089 ), .Z(\SUBBYTES[0].a/n1087 ) );
  XOR \SUBBYTES[0].a/U4484  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/w1947 ), .Z(
        \SUBBYTES[0].a/n1088 ) );
  XOR \SUBBYTES[0].a/U4483  ( .A(\SUBBYTES[0].a/w1854 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1089 ) );
  XOR \SUBBYTES[0].a/U4482  ( .A(\SUBBYTES[0].a/w1840 ), .B(
        \SUBBYTES[0].a/w1842 ), .Z(\SUBBYTES[0].a/n1090 ) );
  XOR \SUBBYTES[0].a/U4481  ( .A(\SUBBYTES[0].a/n1092 ), .B(
        \SUBBYTES[0].a/n1091 ), .Z(\SUBBYTES[0].a/w1864 ) );
  XOR \SUBBYTES[0].a/U4480  ( .A(\SUBBYTES[0].a/n1559 ), .B(
        \SUBBYTES[0].a/n1093 ), .Z(\SUBBYTES[0].a/n1091 ) );
  XOR \SUBBYTES[0].a/U4479  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1560 ), .Z(
        \SUBBYTES[0].a/n1092 ) );
  XOR \SUBBYTES[0].a/U4478  ( .A(\SUBBYTES[0].a/w1854 ), .B(
        \SUBBYTES[0].a/w1855 ), .Z(\SUBBYTES[0].a/n1093 ) );
  XOR \SUBBYTES[0].a/U4477  ( .A(\SUBBYTES[0].a/n1095 ), .B(
        \SUBBYTES[0].a/n1094 ), .Z(\SUBBYTES[0].a/w1880 ) );
  XOR \SUBBYTES[0].a/U4476  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1096 ), .Z(
        \SUBBYTES[0].a/n1094 ) );
  XOR \SUBBYTES[0].a/U4475  ( .A(\SUBBYTES[0].a/w1855 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1095 ) );
  XOR \SUBBYTES[0].a/U4474  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1840 ), .Z(\SUBBYTES[0].a/n1096 ) );
  XOR \SUBBYTES[0].a/U4473  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1097 ), .Z(
        \SUBBYTES[0].a/n1561 ) );
  XOR \SUBBYTES[0].a/U4472  ( .A(\w1[0][67] ), .B(\w1[0][66] ), .Z(
        \SUBBYTES[0].a/n1097 ) );
  XOR \SUBBYTES[0].a/U4471  ( .A(\w1[0][70] ), .B(\SUBBYTES[0].a/n1561 ), .Z(
        \SUBBYTES[0].a/w1722 ) );
  XOR \SUBBYTES[0].a/U4470  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/w1609 ) );
  XOR \SUBBYTES[0].a/U4469  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/n1098 ), .Z(
        \SUBBYTES[0].a/w1610 ) );
  XOR \SUBBYTES[0].a/U4468  ( .A(\w1[0][70] ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1098 ) );
  XOR \SUBBYTES[0].a/U4467  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1561 ), .Z(
        \SUBBYTES[0].a/w1740 ) );
  XOR \SUBBYTES[0].a/U4466  ( .A(\SUBBYTES[0].a/n1100 ), .B(
        \SUBBYTES[0].a/n1099 ), .Z(\SUBBYTES[0].a/w1733 ) );
  XOR \SUBBYTES[0].a/U4465  ( .A(\w1[0][67] ), .B(\w1[0][65] ), .Z(
        \SUBBYTES[0].a/n1099 ) );
  XOR \SUBBYTES[0].a/U4464  ( .A(\w1[0][71] ), .B(\w1[0][68] ), .Z(
        \SUBBYTES[0].a/n1100 ) );
  XOR \SUBBYTES[0].a/U4463  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1733 ), .Z(
        \SUBBYTES[0].a/w1612 ) );
  XOR \SUBBYTES[0].a/U4462  ( .A(\SUBBYTES[0].a/n1102 ), .B(
        \SUBBYTES[0].a/n1101 ), .Z(\SUBBYTES[0].a/w1720 ) );
  XOR \SUBBYTES[0].a/U4461  ( .A(\SUBBYTES[0].a/w1681 ), .B(n8), .Z(
        \SUBBYTES[0].a/n1101 ) );
  XOR \SUBBYTES[0].a/U4460  ( .A(\SUBBYTES[0].a/w1674 ), .B(
        \SUBBYTES[0].a/w1677 ), .Z(\SUBBYTES[0].a/n1102 ) );
  XOR \SUBBYTES[0].a/U4459  ( .A(\SUBBYTES[0].a/n1104 ), .B(
        \SUBBYTES[0].a/n1103 ), .Z(\SUBBYTES[0].a/w1721 ) );
  XOR \SUBBYTES[0].a/U4458  ( .A(\SUBBYTES[0].a/w1681 ), .B(
        \SUBBYTES[0].a/n80 ), .Z(\SUBBYTES[0].a/n1103 ) );
  XOR \SUBBYTES[0].a/U4457  ( .A(\SUBBYTES[0].a/w1674 ), .B(
        \SUBBYTES[0].a/n79 ), .Z(\SUBBYTES[0].a/n1104 ) );
  XOR \SUBBYTES[0].a/U4456  ( .A(\SUBBYTES[0].a/w1733 ), .B(
        \SUBBYTES[0].a/n1105 ), .Z(\SUBBYTES[0].a/w1723 ) );
  XOR \SUBBYTES[0].a/U4455  ( .A(\w1[0][70] ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1105 ) );
  XOR \SUBBYTES[0].a/U4454  ( .A(\SUBBYTES[0].a/n1107 ), .B(
        \SUBBYTES[0].a/n1106 ), .Z(\SUBBYTES[0].a/w1724 ) );
  XOR \SUBBYTES[0].a/U4453  ( .A(\SUBBYTES[0].a/n80 ), .B(n8), .Z(
        \SUBBYTES[0].a/n1106 ) );
  XOR \SUBBYTES[0].a/U4452  ( .A(\SUBBYTES[0].a/n79 ), .B(
        \SUBBYTES[0].a/w1677 ), .Z(\SUBBYTES[0].a/n1107 ) );
  XOR \SUBBYTES[0].a/U4451  ( .A(\w1[0][71] ), .B(\w1[0][66] ), .Z(
        \SUBBYTES[0].a/n1567 ) );
  XOR \SUBBYTES[0].a/U4450  ( .A(\SUBBYTES[0].a/n1567 ), .B(
        \SUBBYTES[0].a/n1108 ), .Z(\SUBBYTES[0].a/w1725 ) );
  XOR \SUBBYTES[0].a/U4449  ( .A(\w1[0][69] ), .B(\w1[0][68] ), .Z(
        \SUBBYTES[0].a/n1108 ) );
  XOR \SUBBYTES[0].a/U4448  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1613 ) );
  XOR \SUBBYTES[0].a/U4447  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1614 ) );
  XOR \SUBBYTES[0].a/U4446  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1615 ) );
  XOR \SUBBYTES[0].a/U4445  ( .A(\SUBBYTES[0].a/w1614 ), .B(
        \SUBBYTES[0].a/n1567 ), .Z(\SUBBYTES[0].a/w1616 ) );
  XOR \SUBBYTES[0].a/U4444  ( .A(\SUBBYTES[0].a/n1567 ), .B(
        \SUBBYTES[0].a/n1109 ), .Z(\SUBBYTES[0].a/w1701 ) );
  XOR \SUBBYTES[0].a/U4443  ( .A(\w1[0][68] ), .B(\w1[0][65] ), .Z(
        \SUBBYTES[0].a/n1109 ) );
  XOR \SUBBYTES[0].a/U4442  ( .A(\SUBBYTES[0].a/n1111 ), .B(
        \SUBBYTES[0].a/n1110 ), .Z(\SUBBYTES[0].a/n1564 ) );
  XOR \SUBBYTES[0].a/U4441  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/n1112 ), .Z(
        \SUBBYTES[0].a/n1110 ) );
  XOR \SUBBYTES[0].a/U4440  ( .A(\SUBBYTES[0].a/w1666 ), .B(\w1[0][70] ), .Z(
        \SUBBYTES[0].a/n1111 ) );
  XOR \SUBBYTES[0].a/U4439  ( .A(\SUBBYTES[0].a/w1640 ), .B(
        \SUBBYTES[0].a/w1647 ), .Z(\SUBBYTES[0].a/n1112 ) );
  XOR \SUBBYTES[0].a/U4438  ( .A(\SUBBYTES[0].a/n1114 ), .B(
        \SUBBYTES[0].a/n1113 ), .Z(\SUBBYTES[0].a/n1562 ) );
  XOR \SUBBYTES[0].a/U4437  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1115 ), .Z(
        \SUBBYTES[0].a/n1113 ) );
  XOR \SUBBYTES[0].a/U4436  ( .A(\SUBBYTES[0].a/w1665 ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1114 ) );
  XOR \SUBBYTES[0].a/U4435  ( .A(\SUBBYTES[0].a/w1641 ), .B(
        \SUBBYTES[0].a/w1648 ), .Z(\SUBBYTES[0].a/n1115 ) );
  XOR \SUBBYTES[0].a/U4434  ( .A(\SUBBYTES[0].a/n1564 ), .B(
        \SUBBYTES[0].a/n1562 ), .Z(\SUBBYTES[0].a/w1671 ) );
  XOR \SUBBYTES[0].a/U4433  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1116 ), .Z(
        \SUBBYTES[0].a/n1565 ) );
  XOR \SUBBYTES[0].a/U4432  ( .A(\SUBBYTES[0].a/w1633 ), .B(
        \SUBBYTES[0].a/w1643 ), .Z(\SUBBYTES[0].a/n1116 ) );
  XOR \SUBBYTES[0].a/U4431  ( .A(\SUBBYTES[0].a/n1118 ), .B(
        \SUBBYTES[0].a/n1117 ), .Z(\SUBBYTES[0].a/w1658 ) );
  XOR \SUBBYTES[0].a/U4430  ( .A(\SUBBYTES[0].a/n1565 ), .B(
        \SUBBYTES[0].a/n1119 ), .Z(\SUBBYTES[0].a/n1117 ) );
  XOR \SUBBYTES[0].a/U4429  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/n1118 ) );
  XOR \SUBBYTES[0].a/U4428  ( .A(\SUBBYTES[0].a/w1635 ), .B(
        \SUBBYTES[0].a/w1640 ), .Z(\SUBBYTES[0].a/n1119 ) );
  XOR \SUBBYTES[0].a/U4427  ( .A(\SUBBYTES[0].a/n1121 ), .B(
        \SUBBYTES[0].a/n1120 ), .Z(\SUBBYTES[0].a/n1563 ) );
  XOR \SUBBYTES[0].a/U4426  ( .A(\SUBBYTES[0].a/w1668 ), .B(\w1[0][71] ), .Z(
        \SUBBYTES[0].a/n1120 ) );
  XOR \SUBBYTES[0].a/U4425  ( .A(\SUBBYTES[0].a/w1643 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1121 ) );
  XOR \SUBBYTES[0].a/U4424  ( .A(\SUBBYTES[0].a/n1562 ), .B(
        \SUBBYTES[0].a/n1563 ), .Z(\SUBBYTES[0].a/w1670 ) );
  XOR \SUBBYTES[0].a/U4423  ( .A(\w1[0][67] ), .B(\SUBBYTES[0].a/n1122 ), .Z(
        \SUBBYTES[0].a/n1566 ) );
  XOR \SUBBYTES[0].a/U4422  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1635 ), .Z(\SUBBYTES[0].a/n1122 ) );
  XOR \SUBBYTES[0].a/U4421  ( .A(\SUBBYTES[0].a/n1124 ), .B(
        \SUBBYTES[0].a/n1123 ), .Z(\SUBBYTES[0].a/w1659 ) );
  XOR \SUBBYTES[0].a/U4420  ( .A(\SUBBYTES[0].a/n1566 ), .B(
        \SUBBYTES[0].a/n1125 ), .Z(\SUBBYTES[0].a/n1123 ) );
  XOR \SUBBYTES[0].a/U4419  ( .A(\w1[0][70] ), .B(\SUBBYTES[0].a/w1701 ), .Z(
        \SUBBYTES[0].a/n1124 ) );
  XOR \SUBBYTES[0].a/U4418  ( .A(\SUBBYTES[0].a/w1640 ), .B(
        \SUBBYTES[0].a/w1641 ), .Z(\SUBBYTES[0].a/n1125 ) );
  XOR \SUBBYTES[0].a/U4417  ( .A(\SUBBYTES[0].a/n1564 ), .B(
        \SUBBYTES[0].a/n1563 ), .Z(\SUBBYTES[0].a/w1679 ) );
  XOR \SUBBYTES[0].a/U4416  ( .A(\SUBBYTES[0].a/n1127 ), .B(
        \SUBBYTES[0].a/n1126 ), .Z(\SUBBYTES[0].a/w1680 ) );
  XOR \SUBBYTES[0].a/U4415  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/n1565 ), .Z(
        \SUBBYTES[0].a/n1126 ) );
  XOR \SUBBYTES[0].a/U4414  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1641 ), .Z(\SUBBYTES[0].a/n1127 ) );
  XOR \SUBBYTES[0].a/U4413  ( .A(\SUBBYTES[0].a/n1129 ), .B(
        \SUBBYTES[0].a/n1128 ), .Z(\SUBBYTES[0].a/w1656 ) );
  XOR \SUBBYTES[0].a/U4412  ( .A(\SUBBYTES[0].a/n1131 ), .B(
        \SUBBYTES[0].a/n1130 ), .Z(\SUBBYTES[0].a/n1128 ) );
  XOR \SUBBYTES[0].a/U4411  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/w1740 ), .Z(
        \SUBBYTES[0].a/n1129 ) );
  XOR \SUBBYTES[0].a/U4410  ( .A(\SUBBYTES[0].a/w1647 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1130 ) );
  XOR \SUBBYTES[0].a/U4409  ( .A(\SUBBYTES[0].a/w1633 ), .B(
        \SUBBYTES[0].a/w1635 ), .Z(\SUBBYTES[0].a/n1131 ) );
  XOR \SUBBYTES[0].a/U4408  ( .A(\SUBBYTES[0].a/n1133 ), .B(
        \SUBBYTES[0].a/n1132 ), .Z(\SUBBYTES[0].a/w1657 ) );
  XOR \SUBBYTES[0].a/U4407  ( .A(\SUBBYTES[0].a/n1566 ), .B(
        \SUBBYTES[0].a/n1134 ), .Z(\SUBBYTES[0].a/n1132 ) );
  XOR \SUBBYTES[0].a/U4406  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1567 ), .Z(
        \SUBBYTES[0].a/n1133 ) );
  XOR \SUBBYTES[0].a/U4405  ( .A(\SUBBYTES[0].a/w1647 ), .B(
        \SUBBYTES[0].a/w1648 ), .Z(\SUBBYTES[0].a/n1134 ) );
  XOR \SUBBYTES[0].a/U4404  ( .A(\SUBBYTES[0].a/n1136 ), .B(
        \SUBBYTES[0].a/n1135 ), .Z(\SUBBYTES[0].a/w1673 ) );
  XOR \SUBBYTES[0].a/U4403  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1137 ), .Z(
        \SUBBYTES[0].a/n1135 ) );
  XOR \SUBBYTES[0].a/U4402  ( .A(\SUBBYTES[0].a/w1648 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1136 ) );
  XOR \SUBBYTES[0].a/U4401  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1633 ), .Z(\SUBBYTES[0].a/n1137 ) );
  XOR \SUBBYTES[0].a/U4400  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1138 ), .Z(
        \SUBBYTES[0].a/n1568 ) );
  XOR \SUBBYTES[0].a/U4399  ( .A(\w1[0][75] ), .B(\w1[0][74] ), .Z(
        \SUBBYTES[0].a/n1138 ) );
  XOR \SUBBYTES[0].a/U4398  ( .A(\w1[0][78] ), .B(\SUBBYTES[0].a/n1568 ), .Z(
        \SUBBYTES[0].a/w1515 ) );
  XOR \SUBBYTES[0].a/U4397  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/w1402 ) );
  XOR \SUBBYTES[0].a/U4396  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/n1139 ), .Z(
        \SUBBYTES[0].a/w1403 ) );
  XOR \SUBBYTES[0].a/U4395  ( .A(\w1[0][78] ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1139 ) );
  XOR \SUBBYTES[0].a/U4394  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1568 ), .Z(
        \SUBBYTES[0].a/w1533 ) );
  XOR \SUBBYTES[0].a/U4393  ( .A(\SUBBYTES[0].a/n1141 ), .B(
        \SUBBYTES[0].a/n1140 ), .Z(\SUBBYTES[0].a/w1526 ) );
  XOR \SUBBYTES[0].a/U4392  ( .A(\w1[0][75] ), .B(\w1[0][73] ), .Z(
        \SUBBYTES[0].a/n1140 ) );
  XOR \SUBBYTES[0].a/U4391  ( .A(\w1[0][79] ), .B(\w1[0][76] ), .Z(
        \SUBBYTES[0].a/n1141 ) );
  XOR \SUBBYTES[0].a/U4390  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1526 ), .Z(
        \SUBBYTES[0].a/w1405 ) );
  XOR \SUBBYTES[0].a/U4389  ( .A(\SUBBYTES[0].a/n1143 ), .B(
        \SUBBYTES[0].a/n1142 ), .Z(\SUBBYTES[0].a/w1513 ) );
  XOR \SUBBYTES[0].a/U4388  ( .A(\SUBBYTES[0].a/w1474 ), .B(n7), .Z(
        \SUBBYTES[0].a/n1142 ) );
  XOR \SUBBYTES[0].a/U4387  ( .A(\SUBBYTES[0].a/w1467 ), .B(
        \SUBBYTES[0].a/w1470 ), .Z(\SUBBYTES[0].a/n1143 ) );
  XOR \SUBBYTES[0].a/U4386  ( .A(\SUBBYTES[0].a/n1145 ), .B(
        \SUBBYTES[0].a/n1144 ), .Z(\SUBBYTES[0].a/w1514 ) );
  XOR \SUBBYTES[0].a/U4385  ( .A(\SUBBYTES[0].a/w1474 ), .B(
        \SUBBYTES[0].a/n70 ), .Z(\SUBBYTES[0].a/n1144 ) );
  XOR \SUBBYTES[0].a/U4384  ( .A(\SUBBYTES[0].a/w1467 ), .B(
        \SUBBYTES[0].a/n69 ), .Z(\SUBBYTES[0].a/n1145 ) );
  XOR \SUBBYTES[0].a/U4383  ( .A(\SUBBYTES[0].a/w1526 ), .B(
        \SUBBYTES[0].a/n1146 ), .Z(\SUBBYTES[0].a/w1516 ) );
  XOR \SUBBYTES[0].a/U4382  ( .A(\w1[0][78] ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1146 ) );
  XOR \SUBBYTES[0].a/U4381  ( .A(\SUBBYTES[0].a/n1148 ), .B(
        \SUBBYTES[0].a/n1147 ), .Z(\SUBBYTES[0].a/w1517 ) );
  XOR \SUBBYTES[0].a/U4380  ( .A(\SUBBYTES[0].a/n70 ), .B(n7), .Z(
        \SUBBYTES[0].a/n1147 ) );
  XOR \SUBBYTES[0].a/U4379  ( .A(\SUBBYTES[0].a/n69 ), .B(
        \SUBBYTES[0].a/w1470 ), .Z(\SUBBYTES[0].a/n1148 ) );
  XOR \SUBBYTES[0].a/U4378  ( .A(\w1[0][79] ), .B(\w1[0][74] ), .Z(
        \SUBBYTES[0].a/n1574 ) );
  XOR \SUBBYTES[0].a/U4377  ( .A(\SUBBYTES[0].a/n1574 ), .B(
        \SUBBYTES[0].a/n1149 ), .Z(\SUBBYTES[0].a/w1518 ) );
  XOR \SUBBYTES[0].a/U4376  ( .A(\w1[0][77] ), .B(\w1[0][76] ), .Z(
        \SUBBYTES[0].a/n1149 ) );
  XOR \SUBBYTES[0].a/U4375  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1406 ) );
  XOR \SUBBYTES[0].a/U4374  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1407 ) );
  XOR \SUBBYTES[0].a/U4373  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1408 ) );
  XOR \SUBBYTES[0].a/U4372  ( .A(\SUBBYTES[0].a/w1407 ), .B(
        \SUBBYTES[0].a/n1574 ), .Z(\SUBBYTES[0].a/w1409 ) );
  XOR \SUBBYTES[0].a/U4371  ( .A(\SUBBYTES[0].a/n1574 ), .B(
        \SUBBYTES[0].a/n1150 ), .Z(\SUBBYTES[0].a/w1494 ) );
  XOR \SUBBYTES[0].a/U4370  ( .A(\w1[0][76] ), .B(\w1[0][73] ), .Z(
        \SUBBYTES[0].a/n1150 ) );
  XOR \SUBBYTES[0].a/U4369  ( .A(\SUBBYTES[0].a/n1152 ), .B(
        \SUBBYTES[0].a/n1151 ), .Z(\SUBBYTES[0].a/n1571 ) );
  XOR \SUBBYTES[0].a/U4368  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/n1153 ), .Z(
        \SUBBYTES[0].a/n1151 ) );
  XOR \SUBBYTES[0].a/U4367  ( .A(\SUBBYTES[0].a/w1459 ), .B(\w1[0][78] ), .Z(
        \SUBBYTES[0].a/n1152 ) );
  XOR \SUBBYTES[0].a/U4366  ( .A(\SUBBYTES[0].a/w1433 ), .B(
        \SUBBYTES[0].a/w1440 ), .Z(\SUBBYTES[0].a/n1153 ) );
  XOR \SUBBYTES[0].a/U4365  ( .A(\SUBBYTES[0].a/n1155 ), .B(
        \SUBBYTES[0].a/n1154 ), .Z(\SUBBYTES[0].a/n1569 ) );
  XOR \SUBBYTES[0].a/U4364  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1156 ), .Z(
        \SUBBYTES[0].a/n1154 ) );
  XOR \SUBBYTES[0].a/U4363  ( .A(\SUBBYTES[0].a/w1458 ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1155 ) );
  XOR \SUBBYTES[0].a/U4362  ( .A(\SUBBYTES[0].a/w1434 ), .B(
        \SUBBYTES[0].a/w1441 ), .Z(\SUBBYTES[0].a/n1156 ) );
  XOR \SUBBYTES[0].a/U4361  ( .A(\SUBBYTES[0].a/n1571 ), .B(
        \SUBBYTES[0].a/n1569 ), .Z(\SUBBYTES[0].a/w1464 ) );
  XOR \SUBBYTES[0].a/U4360  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1157 ), .Z(
        \SUBBYTES[0].a/n1572 ) );
  XOR \SUBBYTES[0].a/U4359  ( .A(\SUBBYTES[0].a/w1426 ), .B(
        \SUBBYTES[0].a/w1436 ), .Z(\SUBBYTES[0].a/n1157 ) );
  XOR \SUBBYTES[0].a/U4358  ( .A(\SUBBYTES[0].a/n1159 ), .B(
        \SUBBYTES[0].a/n1158 ), .Z(\SUBBYTES[0].a/w1451 ) );
  XOR \SUBBYTES[0].a/U4357  ( .A(\SUBBYTES[0].a/n1572 ), .B(
        \SUBBYTES[0].a/n1160 ), .Z(\SUBBYTES[0].a/n1158 ) );
  XOR \SUBBYTES[0].a/U4356  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/n1159 ) );
  XOR \SUBBYTES[0].a/U4355  ( .A(\SUBBYTES[0].a/w1428 ), .B(
        \SUBBYTES[0].a/w1433 ), .Z(\SUBBYTES[0].a/n1160 ) );
  XOR \SUBBYTES[0].a/U4354  ( .A(\SUBBYTES[0].a/n1162 ), .B(
        \SUBBYTES[0].a/n1161 ), .Z(\SUBBYTES[0].a/n1570 ) );
  XOR \SUBBYTES[0].a/U4353  ( .A(\SUBBYTES[0].a/w1461 ), .B(\w1[0][79] ), .Z(
        \SUBBYTES[0].a/n1161 ) );
  XOR \SUBBYTES[0].a/U4352  ( .A(\SUBBYTES[0].a/w1436 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1162 ) );
  XOR \SUBBYTES[0].a/U4351  ( .A(\SUBBYTES[0].a/n1569 ), .B(
        \SUBBYTES[0].a/n1570 ), .Z(\SUBBYTES[0].a/w1463 ) );
  XOR \SUBBYTES[0].a/U4350  ( .A(\w1[0][75] ), .B(\SUBBYTES[0].a/n1163 ), .Z(
        \SUBBYTES[0].a/n1573 ) );
  XOR \SUBBYTES[0].a/U4349  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1428 ), .Z(\SUBBYTES[0].a/n1163 ) );
  XOR \SUBBYTES[0].a/U4348  ( .A(\SUBBYTES[0].a/n1165 ), .B(
        \SUBBYTES[0].a/n1164 ), .Z(\SUBBYTES[0].a/w1452 ) );
  XOR \SUBBYTES[0].a/U4347  ( .A(\SUBBYTES[0].a/n1573 ), .B(
        \SUBBYTES[0].a/n1166 ), .Z(\SUBBYTES[0].a/n1164 ) );
  XOR \SUBBYTES[0].a/U4346  ( .A(\w1[0][78] ), .B(\SUBBYTES[0].a/w1494 ), .Z(
        \SUBBYTES[0].a/n1165 ) );
  XOR \SUBBYTES[0].a/U4345  ( .A(\SUBBYTES[0].a/w1433 ), .B(
        \SUBBYTES[0].a/w1434 ), .Z(\SUBBYTES[0].a/n1166 ) );
  XOR \SUBBYTES[0].a/U4344  ( .A(\SUBBYTES[0].a/n1571 ), .B(
        \SUBBYTES[0].a/n1570 ), .Z(\SUBBYTES[0].a/w1472 ) );
  XOR \SUBBYTES[0].a/U4343  ( .A(\SUBBYTES[0].a/n1168 ), .B(
        \SUBBYTES[0].a/n1167 ), .Z(\SUBBYTES[0].a/w1473 ) );
  XOR \SUBBYTES[0].a/U4342  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/n1572 ), .Z(
        \SUBBYTES[0].a/n1167 ) );
  XOR \SUBBYTES[0].a/U4341  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1434 ), .Z(\SUBBYTES[0].a/n1168 ) );
  XOR \SUBBYTES[0].a/U4340  ( .A(\SUBBYTES[0].a/n1170 ), .B(
        \SUBBYTES[0].a/n1169 ), .Z(\SUBBYTES[0].a/w1449 ) );
  XOR \SUBBYTES[0].a/U4339  ( .A(\SUBBYTES[0].a/n1172 ), .B(
        \SUBBYTES[0].a/n1171 ), .Z(\SUBBYTES[0].a/n1169 ) );
  XOR \SUBBYTES[0].a/U4338  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/w1533 ), .Z(
        \SUBBYTES[0].a/n1170 ) );
  XOR \SUBBYTES[0].a/U4337  ( .A(\SUBBYTES[0].a/w1440 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1171 ) );
  XOR \SUBBYTES[0].a/U4336  ( .A(\SUBBYTES[0].a/w1426 ), .B(
        \SUBBYTES[0].a/w1428 ), .Z(\SUBBYTES[0].a/n1172 ) );
  XOR \SUBBYTES[0].a/U4335  ( .A(\SUBBYTES[0].a/n1174 ), .B(
        \SUBBYTES[0].a/n1173 ), .Z(\SUBBYTES[0].a/w1450 ) );
  XOR \SUBBYTES[0].a/U4334  ( .A(\SUBBYTES[0].a/n1573 ), .B(
        \SUBBYTES[0].a/n1175 ), .Z(\SUBBYTES[0].a/n1173 ) );
  XOR \SUBBYTES[0].a/U4333  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1574 ), .Z(
        \SUBBYTES[0].a/n1174 ) );
  XOR \SUBBYTES[0].a/U4332  ( .A(\SUBBYTES[0].a/w1440 ), .B(
        \SUBBYTES[0].a/w1441 ), .Z(\SUBBYTES[0].a/n1175 ) );
  XOR \SUBBYTES[0].a/U4331  ( .A(\SUBBYTES[0].a/n1177 ), .B(
        \SUBBYTES[0].a/n1176 ), .Z(\SUBBYTES[0].a/w1466 ) );
  XOR \SUBBYTES[0].a/U4330  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1178 ), .Z(
        \SUBBYTES[0].a/n1176 ) );
  XOR \SUBBYTES[0].a/U4329  ( .A(\SUBBYTES[0].a/w1441 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1177 ) );
  XOR \SUBBYTES[0].a/U4328  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1426 ), .Z(\SUBBYTES[0].a/n1178 ) );
  XOR \SUBBYTES[0].a/U4327  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1179 ), .Z(
        \SUBBYTES[0].a/n1575 ) );
  XOR \SUBBYTES[0].a/U4326  ( .A(\w1[0][83] ), .B(\w1[0][82] ), .Z(
        \SUBBYTES[0].a/n1179 ) );
  XOR \SUBBYTES[0].a/U4325  ( .A(\w1[0][86] ), .B(\SUBBYTES[0].a/n1575 ), .Z(
        \SUBBYTES[0].a/w1308 ) );
  XOR \SUBBYTES[0].a/U4324  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/w1195 ) );
  XOR \SUBBYTES[0].a/U4323  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/n1180 ), .Z(
        \SUBBYTES[0].a/w1196 ) );
  XOR \SUBBYTES[0].a/U4322  ( .A(\w1[0][86] ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1180 ) );
  XOR \SUBBYTES[0].a/U4321  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1575 ), .Z(
        \SUBBYTES[0].a/w1326 ) );
  XOR \SUBBYTES[0].a/U4320  ( .A(\SUBBYTES[0].a/n1182 ), .B(
        \SUBBYTES[0].a/n1181 ), .Z(\SUBBYTES[0].a/w1319 ) );
  XOR \SUBBYTES[0].a/U4319  ( .A(\w1[0][83] ), .B(\w1[0][81] ), .Z(
        \SUBBYTES[0].a/n1181 ) );
  XOR \SUBBYTES[0].a/U4318  ( .A(\w1[0][87] ), .B(\w1[0][84] ), .Z(
        \SUBBYTES[0].a/n1182 ) );
  XOR \SUBBYTES[0].a/U4317  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1319 ), .Z(
        \SUBBYTES[0].a/w1198 ) );
  XOR \SUBBYTES[0].a/U4316  ( .A(\SUBBYTES[0].a/n1184 ), .B(
        \SUBBYTES[0].a/n1183 ), .Z(\SUBBYTES[0].a/w1306 ) );
  XOR \SUBBYTES[0].a/U4315  ( .A(\SUBBYTES[0].a/w1267 ), .B(n6), .Z(
        \SUBBYTES[0].a/n1183 ) );
  XOR \SUBBYTES[0].a/U4314  ( .A(\SUBBYTES[0].a/w1260 ), .B(
        \SUBBYTES[0].a/w1263 ), .Z(\SUBBYTES[0].a/n1184 ) );
  XOR \SUBBYTES[0].a/U4313  ( .A(\SUBBYTES[0].a/n1186 ), .B(
        \SUBBYTES[0].a/n1185 ), .Z(\SUBBYTES[0].a/w1307 ) );
  XOR \SUBBYTES[0].a/U4312  ( .A(\SUBBYTES[0].a/w1267 ), .B(
        \SUBBYTES[0].a/n60 ), .Z(\SUBBYTES[0].a/n1185 ) );
  XOR \SUBBYTES[0].a/U4311  ( .A(\SUBBYTES[0].a/w1260 ), .B(
        \SUBBYTES[0].a/n59 ), .Z(\SUBBYTES[0].a/n1186 ) );
  XOR \SUBBYTES[0].a/U4310  ( .A(\SUBBYTES[0].a/w1319 ), .B(
        \SUBBYTES[0].a/n1187 ), .Z(\SUBBYTES[0].a/w1309 ) );
  XOR \SUBBYTES[0].a/U4309  ( .A(\w1[0][86] ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1187 ) );
  XOR \SUBBYTES[0].a/U4308  ( .A(\SUBBYTES[0].a/n1189 ), .B(
        \SUBBYTES[0].a/n1188 ), .Z(\SUBBYTES[0].a/w1310 ) );
  XOR \SUBBYTES[0].a/U4307  ( .A(\SUBBYTES[0].a/n60 ), .B(n6), .Z(
        \SUBBYTES[0].a/n1188 ) );
  XOR \SUBBYTES[0].a/U4306  ( .A(\SUBBYTES[0].a/n59 ), .B(
        \SUBBYTES[0].a/w1263 ), .Z(\SUBBYTES[0].a/n1189 ) );
  XOR \SUBBYTES[0].a/U4305  ( .A(\w1[0][87] ), .B(\w1[0][82] ), .Z(
        \SUBBYTES[0].a/n1581 ) );
  XOR \SUBBYTES[0].a/U4304  ( .A(\SUBBYTES[0].a/n1581 ), .B(
        \SUBBYTES[0].a/n1190 ), .Z(\SUBBYTES[0].a/w1311 ) );
  XOR \SUBBYTES[0].a/U4303  ( .A(\w1[0][85] ), .B(\w1[0][84] ), .Z(
        \SUBBYTES[0].a/n1190 ) );
  XOR \SUBBYTES[0].a/U4302  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1199 ) );
  XOR \SUBBYTES[0].a/U4301  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1200 ) );
  XOR \SUBBYTES[0].a/U4300  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1201 ) );
  XOR \SUBBYTES[0].a/U4299  ( .A(\SUBBYTES[0].a/w1200 ), .B(
        \SUBBYTES[0].a/n1581 ), .Z(\SUBBYTES[0].a/w1202 ) );
  XOR \SUBBYTES[0].a/U4298  ( .A(\SUBBYTES[0].a/n1581 ), .B(
        \SUBBYTES[0].a/n1191 ), .Z(\SUBBYTES[0].a/w1287 ) );
  XOR \SUBBYTES[0].a/U4297  ( .A(\w1[0][84] ), .B(\w1[0][81] ), .Z(
        \SUBBYTES[0].a/n1191 ) );
  XOR \SUBBYTES[0].a/U4296  ( .A(\SUBBYTES[0].a/n1193 ), .B(
        \SUBBYTES[0].a/n1192 ), .Z(\SUBBYTES[0].a/n1578 ) );
  XOR \SUBBYTES[0].a/U4295  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/n1194 ), .Z(
        \SUBBYTES[0].a/n1192 ) );
  XOR \SUBBYTES[0].a/U4294  ( .A(\SUBBYTES[0].a/w1252 ), .B(\w1[0][86] ), .Z(
        \SUBBYTES[0].a/n1193 ) );
  XOR \SUBBYTES[0].a/U4293  ( .A(\SUBBYTES[0].a/w1226 ), .B(
        \SUBBYTES[0].a/w1233 ), .Z(\SUBBYTES[0].a/n1194 ) );
  XOR \SUBBYTES[0].a/U4292  ( .A(\SUBBYTES[0].a/n1196 ), .B(
        \SUBBYTES[0].a/n1195 ), .Z(\SUBBYTES[0].a/n1576 ) );
  XOR \SUBBYTES[0].a/U4291  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1197 ), .Z(
        \SUBBYTES[0].a/n1195 ) );
  XOR \SUBBYTES[0].a/U4290  ( .A(\SUBBYTES[0].a/w1251 ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1196 ) );
  XOR \SUBBYTES[0].a/U4289  ( .A(\SUBBYTES[0].a/w1227 ), .B(
        \SUBBYTES[0].a/w1234 ), .Z(\SUBBYTES[0].a/n1197 ) );
  XOR \SUBBYTES[0].a/U4288  ( .A(\SUBBYTES[0].a/n1578 ), .B(
        \SUBBYTES[0].a/n1576 ), .Z(\SUBBYTES[0].a/w1257 ) );
  XOR \SUBBYTES[0].a/U4287  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1198 ), .Z(
        \SUBBYTES[0].a/n1579 ) );
  XOR \SUBBYTES[0].a/U4286  ( .A(\SUBBYTES[0].a/w1219 ), .B(
        \SUBBYTES[0].a/w1229 ), .Z(\SUBBYTES[0].a/n1198 ) );
  XOR \SUBBYTES[0].a/U4285  ( .A(\SUBBYTES[0].a/n1200 ), .B(
        \SUBBYTES[0].a/n1199 ), .Z(\SUBBYTES[0].a/w1244 ) );
  XOR \SUBBYTES[0].a/U4284  ( .A(\SUBBYTES[0].a/n1579 ), .B(
        \SUBBYTES[0].a/n1201 ), .Z(\SUBBYTES[0].a/n1199 ) );
  XOR \SUBBYTES[0].a/U4283  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/n1200 ) );
  XOR \SUBBYTES[0].a/U4282  ( .A(\SUBBYTES[0].a/w1221 ), .B(
        \SUBBYTES[0].a/w1226 ), .Z(\SUBBYTES[0].a/n1201 ) );
  XOR \SUBBYTES[0].a/U4281  ( .A(\SUBBYTES[0].a/n1203 ), .B(
        \SUBBYTES[0].a/n1202 ), .Z(\SUBBYTES[0].a/n1577 ) );
  XOR \SUBBYTES[0].a/U4280  ( .A(\SUBBYTES[0].a/w1254 ), .B(\w1[0][87] ), .Z(
        \SUBBYTES[0].a/n1202 ) );
  XOR \SUBBYTES[0].a/U4279  ( .A(\SUBBYTES[0].a/w1229 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1203 ) );
  XOR \SUBBYTES[0].a/U4278  ( .A(\SUBBYTES[0].a/n1576 ), .B(
        \SUBBYTES[0].a/n1577 ), .Z(\SUBBYTES[0].a/w1256 ) );
  XOR \SUBBYTES[0].a/U4277  ( .A(\w1[0][83] ), .B(\SUBBYTES[0].a/n1204 ), .Z(
        \SUBBYTES[0].a/n1580 ) );
  XOR \SUBBYTES[0].a/U4276  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1221 ), .Z(\SUBBYTES[0].a/n1204 ) );
  XOR \SUBBYTES[0].a/U4275  ( .A(\SUBBYTES[0].a/n1206 ), .B(
        \SUBBYTES[0].a/n1205 ), .Z(\SUBBYTES[0].a/w1245 ) );
  XOR \SUBBYTES[0].a/U4274  ( .A(\SUBBYTES[0].a/n1580 ), .B(
        \SUBBYTES[0].a/n1207 ), .Z(\SUBBYTES[0].a/n1205 ) );
  XOR \SUBBYTES[0].a/U4273  ( .A(\w1[0][86] ), .B(\SUBBYTES[0].a/w1287 ), .Z(
        \SUBBYTES[0].a/n1206 ) );
  XOR \SUBBYTES[0].a/U4272  ( .A(\SUBBYTES[0].a/w1226 ), .B(
        \SUBBYTES[0].a/w1227 ), .Z(\SUBBYTES[0].a/n1207 ) );
  XOR \SUBBYTES[0].a/U4271  ( .A(\SUBBYTES[0].a/n1578 ), .B(
        \SUBBYTES[0].a/n1577 ), .Z(\SUBBYTES[0].a/w1265 ) );
  XOR \SUBBYTES[0].a/U4270  ( .A(\SUBBYTES[0].a/n1209 ), .B(
        \SUBBYTES[0].a/n1208 ), .Z(\SUBBYTES[0].a/w1266 ) );
  XOR \SUBBYTES[0].a/U4269  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/n1579 ), .Z(
        \SUBBYTES[0].a/n1208 ) );
  XOR \SUBBYTES[0].a/U4268  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1227 ), .Z(\SUBBYTES[0].a/n1209 ) );
  XOR \SUBBYTES[0].a/U4267  ( .A(\SUBBYTES[0].a/n1211 ), .B(
        \SUBBYTES[0].a/n1210 ), .Z(\SUBBYTES[0].a/w1242 ) );
  XOR \SUBBYTES[0].a/U4266  ( .A(\SUBBYTES[0].a/n1213 ), .B(
        \SUBBYTES[0].a/n1212 ), .Z(\SUBBYTES[0].a/n1210 ) );
  XOR \SUBBYTES[0].a/U4265  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/w1326 ), .Z(
        \SUBBYTES[0].a/n1211 ) );
  XOR \SUBBYTES[0].a/U4264  ( .A(\SUBBYTES[0].a/w1233 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1212 ) );
  XOR \SUBBYTES[0].a/U4263  ( .A(\SUBBYTES[0].a/w1219 ), .B(
        \SUBBYTES[0].a/w1221 ), .Z(\SUBBYTES[0].a/n1213 ) );
  XOR \SUBBYTES[0].a/U4262  ( .A(\SUBBYTES[0].a/n1215 ), .B(
        \SUBBYTES[0].a/n1214 ), .Z(\SUBBYTES[0].a/w1243 ) );
  XOR \SUBBYTES[0].a/U4261  ( .A(\SUBBYTES[0].a/n1580 ), .B(
        \SUBBYTES[0].a/n1216 ), .Z(\SUBBYTES[0].a/n1214 ) );
  XOR \SUBBYTES[0].a/U4260  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1581 ), .Z(
        \SUBBYTES[0].a/n1215 ) );
  XOR \SUBBYTES[0].a/U4259  ( .A(\SUBBYTES[0].a/w1233 ), .B(
        \SUBBYTES[0].a/w1234 ), .Z(\SUBBYTES[0].a/n1216 ) );
  XOR \SUBBYTES[0].a/U4258  ( .A(\SUBBYTES[0].a/n1218 ), .B(
        \SUBBYTES[0].a/n1217 ), .Z(\SUBBYTES[0].a/w1259 ) );
  XOR \SUBBYTES[0].a/U4257  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1219 ), .Z(
        \SUBBYTES[0].a/n1217 ) );
  XOR \SUBBYTES[0].a/U4256  ( .A(\SUBBYTES[0].a/w1234 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1218 ) );
  XOR \SUBBYTES[0].a/U4255  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1219 ), .Z(\SUBBYTES[0].a/n1219 ) );
  XOR \SUBBYTES[0].a/U4254  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1220 ), .Z(
        \SUBBYTES[0].a/n1582 ) );
  XOR \SUBBYTES[0].a/U4253  ( .A(\w1[0][91] ), .B(\w1[0][90] ), .Z(
        \SUBBYTES[0].a/n1220 ) );
  XOR \SUBBYTES[0].a/U4252  ( .A(\w1[0][94] ), .B(\SUBBYTES[0].a/n1582 ), .Z(
        \SUBBYTES[0].a/w1101 ) );
  XOR \SUBBYTES[0].a/U4251  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/w988 ) );
  XOR \SUBBYTES[0].a/U4250  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/n1221 ), .Z(
        \SUBBYTES[0].a/w989 ) );
  XOR \SUBBYTES[0].a/U4249  ( .A(\w1[0][94] ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1221 ) );
  XOR \SUBBYTES[0].a/U4248  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1582 ), .Z(
        \SUBBYTES[0].a/w1119 ) );
  XOR \SUBBYTES[0].a/U4247  ( .A(\SUBBYTES[0].a/n1223 ), .B(
        \SUBBYTES[0].a/n1222 ), .Z(\SUBBYTES[0].a/w1112 ) );
  XOR \SUBBYTES[0].a/U4246  ( .A(\w1[0][91] ), .B(\w1[0][89] ), .Z(
        \SUBBYTES[0].a/n1222 ) );
  XOR \SUBBYTES[0].a/U4245  ( .A(\w1[0][95] ), .B(\w1[0][92] ), .Z(
        \SUBBYTES[0].a/n1223 ) );
  XOR \SUBBYTES[0].a/U4244  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w1112 ), .Z(
        \SUBBYTES[0].a/w991 ) );
  XOR \SUBBYTES[0].a/U4243  ( .A(\SUBBYTES[0].a/n1225 ), .B(
        \SUBBYTES[0].a/n1224 ), .Z(\SUBBYTES[0].a/w1099 ) );
  XOR \SUBBYTES[0].a/U4242  ( .A(\SUBBYTES[0].a/w1060 ), .B(n5), .Z(
        \SUBBYTES[0].a/n1224 ) );
  XOR \SUBBYTES[0].a/U4241  ( .A(\SUBBYTES[0].a/w1053 ), .B(
        \SUBBYTES[0].a/w1056 ), .Z(\SUBBYTES[0].a/n1225 ) );
  XOR \SUBBYTES[0].a/U4240  ( .A(\SUBBYTES[0].a/n1227 ), .B(
        \SUBBYTES[0].a/n1226 ), .Z(\SUBBYTES[0].a/w1100 ) );
  XOR \SUBBYTES[0].a/U4239  ( .A(\SUBBYTES[0].a/w1060 ), .B(
        \SUBBYTES[0].a/n50 ), .Z(\SUBBYTES[0].a/n1226 ) );
  XOR \SUBBYTES[0].a/U4238  ( .A(\SUBBYTES[0].a/w1053 ), .B(
        \SUBBYTES[0].a/n49 ), .Z(\SUBBYTES[0].a/n1227 ) );
  XOR \SUBBYTES[0].a/U4237  ( .A(\SUBBYTES[0].a/w1112 ), .B(
        \SUBBYTES[0].a/n1228 ), .Z(\SUBBYTES[0].a/w1102 ) );
  XOR \SUBBYTES[0].a/U4236  ( .A(\w1[0][94] ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1228 ) );
  XOR \SUBBYTES[0].a/U4235  ( .A(\SUBBYTES[0].a/n1230 ), .B(
        \SUBBYTES[0].a/n1229 ), .Z(\SUBBYTES[0].a/w1103 ) );
  XOR \SUBBYTES[0].a/U4234  ( .A(\SUBBYTES[0].a/n50 ), .B(n5), .Z(
        \SUBBYTES[0].a/n1229 ) );
  XOR \SUBBYTES[0].a/U4233  ( .A(\SUBBYTES[0].a/n49 ), .B(
        \SUBBYTES[0].a/w1056 ), .Z(\SUBBYTES[0].a/n1230 ) );
  XOR \SUBBYTES[0].a/U4232  ( .A(\w1[0][95] ), .B(\w1[0][90] ), .Z(
        \SUBBYTES[0].a/n1588 ) );
  XOR \SUBBYTES[0].a/U4231  ( .A(\SUBBYTES[0].a/n1588 ), .B(
        \SUBBYTES[0].a/n1231 ), .Z(\SUBBYTES[0].a/w1104 ) );
  XOR \SUBBYTES[0].a/U4230  ( .A(\w1[0][93] ), .B(\w1[0][92] ), .Z(
        \SUBBYTES[0].a/n1231 ) );
  XOR \SUBBYTES[0].a/U4229  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w992 ) );
  XOR \SUBBYTES[0].a/U4228  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w993 ) );
  XOR \SUBBYTES[0].a/U4227  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w994 ) );
  XOR \SUBBYTES[0].a/U4226  ( .A(\SUBBYTES[0].a/w993 ), .B(
        \SUBBYTES[0].a/n1588 ), .Z(\SUBBYTES[0].a/w995 ) );
  XOR \SUBBYTES[0].a/U4225  ( .A(\SUBBYTES[0].a/n1588 ), .B(
        \SUBBYTES[0].a/n1232 ), .Z(\SUBBYTES[0].a/w1080 ) );
  XOR \SUBBYTES[0].a/U4224  ( .A(\w1[0][92] ), .B(\w1[0][89] ), .Z(
        \SUBBYTES[0].a/n1232 ) );
  XOR \SUBBYTES[0].a/U4223  ( .A(\SUBBYTES[0].a/n1234 ), .B(
        \SUBBYTES[0].a/n1233 ), .Z(\SUBBYTES[0].a/n1585 ) );
  XOR \SUBBYTES[0].a/U4222  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/n1235 ), .Z(
        \SUBBYTES[0].a/n1233 ) );
  XOR \SUBBYTES[0].a/U4221  ( .A(\SUBBYTES[0].a/w1045 ), .B(\w1[0][94] ), .Z(
        \SUBBYTES[0].a/n1234 ) );
  XOR \SUBBYTES[0].a/U4220  ( .A(\SUBBYTES[0].a/w1019 ), .B(
        \SUBBYTES[0].a/w1026 ), .Z(\SUBBYTES[0].a/n1235 ) );
  XOR \SUBBYTES[0].a/U4219  ( .A(\SUBBYTES[0].a/n1237 ), .B(
        \SUBBYTES[0].a/n1236 ), .Z(\SUBBYTES[0].a/n1583 ) );
  XOR \SUBBYTES[0].a/U4218  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1238 ), .Z(
        \SUBBYTES[0].a/n1236 ) );
  XOR \SUBBYTES[0].a/U4217  ( .A(\SUBBYTES[0].a/w1044 ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1237 ) );
  XOR \SUBBYTES[0].a/U4216  ( .A(\SUBBYTES[0].a/w1020 ), .B(
        \SUBBYTES[0].a/w1027 ), .Z(\SUBBYTES[0].a/n1238 ) );
  XOR \SUBBYTES[0].a/U4215  ( .A(\SUBBYTES[0].a/n1585 ), .B(
        \SUBBYTES[0].a/n1583 ), .Z(\SUBBYTES[0].a/w1050 ) );
  XOR \SUBBYTES[0].a/U4214  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1239 ), .Z(
        \SUBBYTES[0].a/n1586 ) );
  XOR \SUBBYTES[0].a/U4213  ( .A(\SUBBYTES[0].a/w1012 ), .B(
        \SUBBYTES[0].a/w1022 ), .Z(\SUBBYTES[0].a/n1239 ) );
  XOR \SUBBYTES[0].a/U4212  ( .A(\SUBBYTES[0].a/n1241 ), .B(
        \SUBBYTES[0].a/n1240 ), .Z(\SUBBYTES[0].a/w1037 ) );
  XOR \SUBBYTES[0].a/U4211  ( .A(\SUBBYTES[0].a/n1586 ), .B(
        \SUBBYTES[0].a/n1242 ), .Z(\SUBBYTES[0].a/n1240 ) );
  XOR \SUBBYTES[0].a/U4210  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/n1241 ) );
  XOR \SUBBYTES[0].a/U4209  ( .A(\SUBBYTES[0].a/w1014 ), .B(
        \SUBBYTES[0].a/w1019 ), .Z(\SUBBYTES[0].a/n1242 ) );
  XOR \SUBBYTES[0].a/U4208  ( .A(\SUBBYTES[0].a/n1244 ), .B(
        \SUBBYTES[0].a/n1243 ), .Z(\SUBBYTES[0].a/n1584 ) );
  XOR \SUBBYTES[0].a/U4207  ( .A(\SUBBYTES[0].a/w1047 ), .B(\w1[0][95] ), .Z(
        \SUBBYTES[0].a/n1243 ) );
  XOR \SUBBYTES[0].a/U4206  ( .A(\SUBBYTES[0].a/w1022 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1244 ) );
  XOR \SUBBYTES[0].a/U4205  ( .A(\SUBBYTES[0].a/n1583 ), .B(
        \SUBBYTES[0].a/n1584 ), .Z(\SUBBYTES[0].a/w1049 ) );
  XOR \SUBBYTES[0].a/U4204  ( .A(\w1[0][91] ), .B(\SUBBYTES[0].a/n1245 ), .Z(
        \SUBBYTES[0].a/n1587 ) );
  XOR \SUBBYTES[0].a/U4203  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1014 ), .Z(\SUBBYTES[0].a/n1245 ) );
  XOR \SUBBYTES[0].a/U4202  ( .A(\SUBBYTES[0].a/n1247 ), .B(
        \SUBBYTES[0].a/n1246 ), .Z(\SUBBYTES[0].a/w1038 ) );
  XOR \SUBBYTES[0].a/U4201  ( .A(\SUBBYTES[0].a/n1587 ), .B(
        \SUBBYTES[0].a/n1248 ), .Z(\SUBBYTES[0].a/n1246 ) );
  XOR \SUBBYTES[0].a/U4200  ( .A(\w1[0][94] ), .B(\SUBBYTES[0].a/w1080 ), .Z(
        \SUBBYTES[0].a/n1247 ) );
  XOR \SUBBYTES[0].a/U4199  ( .A(\SUBBYTES[0].a/w1019 ), .B(
        \SUBBYTES[0].a/w1020 ), .Z(\SUBBYTES[0].a/n1248 ) );
  XOR \SUBBYTES[0].a/U4198  ( .A(\SUBBYTES[0].a/n1585 ), .B(
        \SUBBYTES[0].a/n1584 ), .Z(\SUBBYTES[0].a/w1058 ) );
  XOR \SUBBYTES[0].a/U4197  ( .A(\SUBBYTES[0].a/n1250 ), .B(
        \SUBBYTES[0].a/n1249 ), .Z(\SUBBYTES[0].a/w1059 ) );
  XOR \SUBBYTES[0].a/U4196  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/n1586 ), .Z(
        \SUBBYTES[0].a/n1249 ) );
  XOR \SUBBYTES[0].a/U4195  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1020 ), .Z(\SUBBYTES[0].a/n1250 ) );
  XOR \SUBBYTES[0].a/U4194  ( .A(\SUBBYTES[0].a/n1252 ), .B(
        \SUBBYTES[0].a/n1251 ), .Z(\SUBBYTES[0].a/w1035 ) );
  XOR \SUBBYTES[0].a/U4193  ( .A(\SUBBYTES[0].a/n1254 ), .B(
        \SUBBYTES[0].a/n1253 ), .Z(\SUBBYTES[0].a/n1251 ) );
  XOR \SUBBYTES[0].a/U4192  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/w1119 ), .Z(
        \SUBBYTES[0].a/n1252 ) );
  XOR \SUBBYTES[0].a/U4191  ( .A(\SUBBYTES[0].a/w1026 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1253 ) );
  XOR \SUBBYTES[0].a/U4190  ( .A(\SUBBYTES[0].a/w1012 ), .B(
        \SUBBYTES[0].a/w1014 ), .Z(\SUBBYTES[0].a/n1254 ) );
  XOR \SUBBYTES[0].a/U4189  ( .A(\SUBBYTES[0].a/n1256 ), .B(
        \SUBBYTES[0].a/n1255 ), .Z(\SUBBYTES[0].a/w1036 ) );
  XOR \SUBBYTES[0].a/U4188  ( .A(\SUBBYTES[0].a/n1587 ), .B(
        \SUBBYTES[0].a/n1257 ), .Z(\SUBBYTES[0].a/n1255 ) );
  XOR \SUBBYTES[0].a/U4187  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1588 ), .Z(
        \SUBBYTES[0].a/n1256 ) );
  XOR \SUBBYTES[0].a/U4186  ( .A(\SUBBYTES[0].a/w1026 ), .B(
        \SUBBYTES[0].a/w1027 ), .Z(\SUBBYTES[0].a/n1257 ) );
  XOR \SUBBYTES[0].a/U4185  ( .A(\SUBBYTES[0].a/n1259 ), .B(
        \SUBBYTES[0].a/n1258 ), .Z(\SUBBYTES[0].a/w1052 ) );
  XOR \SUBBYTES[0].a/U4184  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1260 ), .Z(
        \SUBBYTES[0].a/n1258 ) );
  XOR \SUBBYTES[0].a/U4183  ( .A(\SUBBYTES[0].a/w1027 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1259 ) );
  XOR \SUBBYTES[0].a/U4182  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1012 ), .Z(\SUBBYTES[0].a/n1260 ) );
  XOR \SUBBYTES[0].a/U4181  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1261 ), .Z(
        \SUBBYTES[0].a/n1589 ) );
  XOR \SUBBYTES[0].a/U4180  ( .A(\w1[0][99] ), .B(\w1[0][98] ), .Z(
        \SUBBYTES[0].a/n1261 ) );
  XOR \SUBBYTES[0].a/U4179  ( .A(\w1[0][102] ), .B(\SUBBYTES[0].a/n1589 ), .Z(
        \SUBBYTES[0].a/w894 ) );
  XOR \SUBBYTES[0].a/U4178  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/w781 ) );
  XOR \SUBBYTES[0].a/U4177  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/n1262 ), .Z(
        \SUBBYTES[0].a/w782 ) );
  XOR \SUBBYTES[0].a/U4176  ( .A(\w1[0][102] ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1262 ) );
  XOR \SUBBYTES[0].a/U4175  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1589 ), .Z(
        \SUBBYTES[0].a/w912 ) );
  XOR \SUBBYTES[0].a/U4174  ( .A(\SUBBYTES[0].a/n1264 ), .B(
        \SUBBYTES[0].a/n1263 ), .Z(\SUBBYTES[0].a/w905 ) );
  XOR \SUBBYTES[0].a/U4173  ( .A(\w1[0][99] ), .B(\w1[0][97] ), .Z(
        \SUBBYTES[0].a/n1263 ) );
  XOR \SUBBYTES[0].a/U4172  ( .A(\w1[0][103] ), .B(\w1[0][100] ), .Z(
        \SUBBYTES[0].a/n1264 ) );
  XOR \SUBBYTES[0].a/U4171  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w905 ), .Z(
        \SUBBYTES[0].a/w784 ) );
  XOR \SUBBYTES[0].a/U4170  ( .A(\SUBBYTES[0].a/n1266 ), .B(
        \SUBBYTES[0].a/n1265 ), .Z(\SUBBYTES[0].a/w892 ) );
  XOR \SUBBYTES[0].a/U4169  ( .A(\SUBBYTES[0].a/w853 ), .B(n4), .Z(
        \SUBBYTES[0].a/n1265 ) );
  XOR \SUBBYTES[0].a/U4168  ( .A(\SUBBYTES[0].a/w846 ), .B(
        \SUBBYTES[0].a/w849 ), .Z(\SUBBYTES[0].a/n1266 ) );
  XOR \SUBBYTES[0].a/U4167  ( .A(\SUBBYTES[0].a/n1268 ), .B(
        \SUBBYTES[0].a/n1267 ), .Z(\SUBBYTES[0].a/w893 ) );
  XOR \SUBBYTES[0].a/U4166  ( .A(\SUBBYTES[0].a/w853 ), .B(\SUBBYTES[0].a/n40 ), .Z(\SUBBYTES[0].a/n1267 ) );
  XOR \SUBBYTES[0].a/U4165  ( .A(\SUBBYTES[0].a/w846 ), .B(\SUBBYTES[0].a/n39 ), .Z(\SUBBYTES[0].a/n1268 ) );
  XOR \SUBBYTES[0].a/U4164  ( .A(\SUBBYTES[0].a/w905 ), .B(
        \SUBBYTES[0].a/n1269 ), .Z(\SUBBYTES[0].a/w895 ) );
  XOR \SUBBYTES[0].a/U4163  ( .A(\w1[0][102] ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1269 ) );
  XOR \SUBBYTES[0].a/U4162  ( .A(\SUBBYTES[0].a/n1271 ), .B(
        \SUBBYTES[0].a/n1270 ), .Z(\SUBBYTES[0].a/w896 ) );
  XOR \SUBBYTES[0].a/U4161  ( .A(\SUBBYTES[0].a/n40 ), .B(n4), .Z(
        \SUBBYTES[0].a/n1270 ) );
  XOR \SUBBYTES[0].a/U4160  ( .A(\SUBBYTES[0].a/n39 ), .B(\SUBBYTES[0].a/w849 ), .Z(\SUBBYTES[0].a/n1271 ) );
  XOR \SUBBYTES[0].a/U4159  ( .A(\w1[0][103] ), .B(\w1[0][98] ), .Z(
        \SUBBYTES[0].a/n1595 ) );
  XOR \SUBBYTES[0].a/U4158  ( .A(\SUBBYTES[0].a/n1595 ), .B(
        \SUBBYTES[0].a/n1272 ), .Z(\SUBBYTES[0].a/w897 ) );
  XOR \SUBBYTES[0].a/U4157  ( .A(\w1[0][101] ), .B(\w1[0][100] ), .Z(
        \SUBBYTES[0].a/n1272 ) );
  XOR \SUBBYTES[0].a/U4156  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w785 ) );
  XOR \SUBBYTES[0].a/U4155  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w786 ) );
  XOR \SUBBYTES[0].a/U4154  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w787 ) );
  XOR \SUBBYTES[0].a/U4153  ( .A(\SUBBYTES[0].a/w786 ), .B(
        \SUBBYTES[0].a/n1595 ), .Z(\SUBBYTES[0].a/w788 ) );
  XOR \SUBBYTES[0].a/U4152  ( .A(\SUBBYTES[0].a/n1595 ), .B(
        \SUBBYTES[0].a/n1273 ), .Z(\SUBBYTES[0].a/w873 ) );
  XOR \SUBBYTES[0].a/U4151  ( .A(\w1[0][100] ), .B(\w1[0][97] ), .Z(
        \SUBBYTES[0].a/n1273 ) );
  XOR \SUBBYTES[0].a/U4150  ( .A(\SUBBYTES[0].a/n1275 ), .B(
        \SUBBYTES[0].a/n1274 ), .Z(\SUBBYTES[0].a/n1592 ) );
  XOR \SUBBYTES[0].a/U4149  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/n1276 ), .Z(
        \SUBBYTES[0].a/n1274 ) );
  XOR \SUBBYTES[0].a/U4148  ( .A(\SUBBYTES[0].a/w838 ), .B(\w1[0][102] ), .Z(
        \SUBBYTES[0].a/n1275 ) );
  XOR \SUBBYTES[0].a/U4147  ( .A(\SUBBYTES[0].a/w812 ), .B(
        \SUBBYTES[0].a/w819 ), .Z(\SUBBYTES[0].a/n1276 ) );
  XOR \SUBBYTES[0].a/U4146  ( .A(\SUBBYTES[0].a/n1278 ), .B(
        \SUBBYTES[0].a/n1277 ), .Z(\SUBBYTES[0].a/n1590 ) );
  XOR \SUBBYTES[0].a/U4145  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1279 ), .Z(
        \SUBBYTES[0].a/n1277 ) );
  XOR \SUBBYTES[0].a/U4144  ( .A(\SUBBYTES[0].a/w837 ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1278 ) );
  XOR \SUBBYTES[0].a/U4143  ( .A(\SUBBYTES[0].a/w813 ), .B(
        \SUBBYTES[0].a/w820 ), .Z(\SUBBYTES[0].a/n1279 ) );
  XOR \SUBBYTES[0].a/U4142  ( .A(\SUBBYTES[0].a/n1592 ), .B(
        \SUBBYTES[0].a/n1590 ), .Z(\SUBBYTES[0].a/w843 ) );
  XOR \SUBBYTES[0].a/U4141  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1280 ), .Z(
        \SUBBYTES[0].a/n1593 ) );
  XOR \SUBBYTES[0].a/U4140  ( .A(\SUBBYTES[0].a/w805 ), .B(
        \SUBBYTES[0].a/w815 ), .Z(\SUBBYTES[0].a/n1280 ) );
  XOR \SUBBYTES[0].a/U4139  ( .A(\SUBBYTES[0].a/n1282 ), .B(
        \SUBBYTES[0].a/n1281 ), .Z(\SUBBYTES[0].a/w830 ) );
  XOR \SUBBYTES[0].a/U4138  ( .A(\SUBBYTES[0].a/n1593 ), .B(
        \SUBBYTES[0].a/n1283 ), .Z(\SUBBYTES[0].a/n1281 ) );
  XOR \SUBBYTES[0].a/U4137  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/n1282 ) );
  XOR \SUBBYTES[0].a/U4136  ( .A(\SUBBYTES[0].a/w807 ), .B(
        \SUBBYTES[0].a/w812 ), .Z(\SUBBYTES[0].a/n1283 ) );
  XOR \SUBBYTES[0].a/U4135  ( .A(\SUBBYTES[0].a/n1285 ), .B(
        \SUBBYTES[0].a/n1284 ), .Z(\SUBBYTES[0].a/n1591 ) );
  XOR \SUBBYTES[0].a/U4134  ( .A(\SUBBYTES[0].a/w840 ), .B(\w1[0][103] ), .Z(
        \SUBBYTES[0].a/n1284 ) );
  XOR \SUBBYTES[0].a/U4133  ( .A(\SUBBYTES[0].a/w815 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1285 ) );
  XOR \SUBBYTES[0].a/U4132  ( .A(\SUBBYTES[0].a/n1590 ), .B(
        \SUBBYTES[0].a/n1591 ), .Z(\SUBBYTES[0].a/w842 ) );
  XOR \SUBBYTES[0].a/U4131  ( .A(\w1[0][99] ), .B(\SUBBYTES[0].a/n1286 ), .Z(
        \SUBBYTES[0].a/n1594 ) );
  XOR \SUBBYTES[0].a/U4130  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w807 ), .Z(\SUBBYTES[0].a/n1286 ) );
  XOR \SUBBYTES[0].a/U4129  ( .A(\SUBBYTES[0].a/n1288 ), .B(
        \SUBBYTES[0].a/n1287 ), .Z(\SUBBYTES[0].a/w831 ) );
  XOR \SUBBYTES[0].a/U4128  ( .A(\SUBBYTES[0].a/n1594 ), .B(
        \SUBBYTES[0].a/n1289 ), .Z(\SUBBYTES[0].a/n1287 ) );
  XOR \SUBBYTES[0].a/U4127  ( .A(\w1[0][102] ), .B(\SUBBYTES[0].a/w873 ), .Z(
        \SUBBYTES[0].a/n1288 ) );
  XOR \SUBBYTES[0].a/U4126  ( .A(\SUBBYTES[0].a/w812 ), .B(
        \SUBBYTES[0].a/w813 ), .Z(\SUBBYTES[0].a/n1289 ) );
  XOR \SUBBYTES[0].a/U4125  ( .A(\SUBBYTES[0].a/n1592 ), .B(
        \SUBBYTES[0].a/n1591 ), .Z(\SUBBYTES[0].a/w851 ) );
  XOR \SUBBYTES[0].a/U4124  ( .A(\SUBBYTES[0].a/n1291 ), .B(
        \SUBBYTES[0].a/n1290 ), .Z(\SUBBYTES[0].a/w852 ) );
  XOR \SUBBYTES[0].a/U4123  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/n1593 ), .Z(
        \SUBBYTES[0].a/n1290 ) );
  XOR \SUBBYTES[0].a/U4122  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w813 ), .Z(\SUBBYTES[0].a/n1291 ) );
  XOR \SUBBYTES[0].a/U4121  ( .A(\SUBBYTES[0].a/n1293 ), .B(
        \SUBBYTES[0].a/n1292 ), .Z(\SUBBYTES[0].a/w828 ) );
  XOR \SUBBYTES[0].a/U4120  ( .A(\SUBBYTES[0].a/n1295 ), .B(
        \SUBBYTES[0].a/n1294 ), .Z(\SUBBYTES[0].a/n1292 ) );
  XOR \SUBBYTES[0].a/U4119  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/w912 ), .Z(
        \SUBBYTES[0].a/n1293 ) );
  XOR \SUBBYTES[0].a/U4118  ( .A(\SUBBYTES[0].a/w819 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1294 ) );
  XOR \SUBBYTES[0].a/U4117  ( .A(\SUBBYTES[0].a/w805 ), .B(
        \SUBBYTES[0].a/w807 ), .Z(\SUBBYTES[0].a/n1295 ) );
  XOR \SUBBYTES[0].a/U4116  ( .A(\SUBBYTES[0].a/n1297 ), .B(
        \SUBBYTES[0].a/n1296 ), .Z(\SUBBYTES[0].a/w829 ) );
  XOR \SUBBYTES[0].a/U4115  ( .A(\SUBBYTES[0].a/n1594 ), .B(
        \SUBBYTES[0].a/n1298 ), .Z(\SUBBYTES[0].a/n1296 ) );
  XOR \SUBBYTES[0].a/U4114  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1595 ), .Z(
        \SUBBYTES[0].a/n1297 ) );
  XOR \SUBBYTES[0].a/U4113  ( .A(\SUBBYTES[0].a/w819 ), .B(
        \SUBBYTES[0].a/w820 ), .Z(\SUBBYTES[0].a/n1298 ) );
  XOR \SUBBYTES[0].a/U4112  ( .A(\SUBBYTES[0].a/n1300 ), .B(
        \SUBBYTES[0].a/n1299 ), .Z(\SUBBYTES[0].a/w845 ) );
  XOR \SUBBYTES[0].a/U4111  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1301 ), .Z(
        \SUBBYTES[0].a/n1299 ) );
  XOR \SUBBYTES[0].a/U4110  ( .A(\SUBBYTES[0].a/w820 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1300 ) );
  XOR \SUBBYTES[0].a/U4109  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w805 ), .Z(\SUBBYTES[0].a/n1301 ) );
  XOR \SUBBYTES[0].a/U4108  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1302 ), .Z(
        \SUBBYTES[0].a/n1596 ) );
  XOR \SUBBYTES[0].a/U4107  ( .A(\w1[0][107] ), .B(\w1[0][106] ), .Z(
        \SUBBYTES[0].a/n1302 ) );
  XOR \SUBBYTES[0].a/U4106  ( .A(\w1[0][110] ), .B(\SUBBYTES[0].a/n1596 ), .Z(
        \SUBBYTES[0].a/w687 ) );
  XOR \SUBBYTES[0].a/U4105  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/w574 ) );
  XOR \SUBBYTES[0].a/U4104  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/n1303 ), .Z(
        \SUBBYTES[0].a/w575 ) );
  XOR \SUBBYTES[0].a/U4103  ( .A(\w1[0][110] ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1303 ) );
  XOR \SUBBYTES[0].a/U4102  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1596 ), .Z(
        \SUBBYTES[0].a/w705 ) );
  XOR \SUBBYTES[0].a/U4101  ( .A(\SUBBYTES[0].a/n1305 ), .B(
        \SUBBYTES[0].a/n1304 ), .Z(\SUBBYTES[0].a/w698 ) );
  XOR \SUBBYTES[0].a/U4100  ( .A(\w1[0][107] ), .B(\w1[0][105] ), .Z(
        \SUBBYTES[0].a/n1304 ) );
  XOR \SUBBYTES[0].a/U4099  ( .A(\w1[0][111] ), .B(\w1[0][108] ), .Z(
        \SUBBYTES[0].a/n1305 ) );
  XOR \SUBBYTES[0].a/U4098  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w698 ), .Z(
        \SUBBYTES[0].a/w577 ) );
  XOR \SUBBYTES[0].a/U4097  ( .A(\SUBBYTES[0].a/n1307 ), .B(
        \SUBBYTES[0].a/n1306 ), .Z(\SUBBYTES[0].a/w685 ) );
  XOR \SUBBYTES[0].a/U4096  ( .A(\SUBBYTES[0].a/w646 ), .B(n3), .Z(
        \SUBBYTES[0].a/n1306 ) );
  XOR \SUBBYTES[0].a/U4095  ( .A(\SUBBYTES[0].a/w639 ), .B(
        \SUBBYTES[0].a/w642 ), .Z(\SUBBYTES[0].a/n1307 ) );
  XOR \SUBBYTES[0].a/U4094  ( .A(\SUBBYTES[0].a/n1309 ), .B(
        \SUBBYTES[0].a/n1308 ), .Z(\SUBBYTES[0].a/w686 ) );
  XOR \SUBBYTES[0].a/U4093  ( .A(\SUBBYTES[0].a/w646 ), .B(\SUBBYTES[0].a/n30 ), .Z(\SUBBYTES[0].a/n1308 ) );
  XOR \SUBBYTES[0].a/U4092  ( .A(\SUBBYTES[0].a/w639 ), .B(\SUBBYTES[0].a/n29 ), .Z(\SUBBYTES[0].a/n1309 ) );
  XOR \SUBBYTES[0].a/U4091  ( .A(\SUBBYTES[0].a/w698 ), .B(
        \SUBBYTES[0].a/n1310 ), .Z(\SUBBYTES[0].a/w688 ) );
  XOR \SUBBYTES[0].a/U4090  ( .A(\w1[0][110] ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1310 ) );
  XOR \SUBBYTES[0].a/U4089  ( .A(\SUBBYTES[0].a/n1312 ), .B(
        \SUBBYTES[0].a/n1311 ), .Z(\SUBBYTES[0].a/w689 ) );
  XOR \SUBBYTES[0].a/U4088  ( .A(\SUBBYTES[0].a/n30 ), .B(n3), .Z(
        \SUBBYTES[0].a/n1311 ) );
  XOR \SUBBYTES[0].a/U4087  ( .A(\SUBBYTES[0].a/n29 ), .B(\SUBBYTES[0].a/w642 ), .Z(\SUBBYTES[0].a/n1312 ) );
  XOR \SUBBYTES[0].a/U4086  ( .A(\w1[0][111] ), .B(\w1[0][106] ), .Z(
        \SUBBYTES[0].a/n1602 ) );
  XOR \SUBBYTES[0].a/U4085  ( .A(\SUBBYTES[0].a/n1602 ), .B(
        \SUBBYTES[0].a/n1313 ), .Z(\SUBBYTES[0].a/w690 ) );
  XOR \SUBBYTES[0].a/U4084  ( .A(\w1[0][109] ), .B(\w1[0][108] ), .Z(
        \SUBBYTES[0].a/n1313 ) );
  XOR \SUBBYTES[0].a/U4083  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w578 ) );
  XOR \SUBBYTES[0].a/U4082  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w579 ) );
  XOR \SUBBYTES[0].a/U4081  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w580 ) );
  XOR \SUBBYTES[0].a/U4080  ( .A(\SUBBYTES[0].a/w579 ), .B(
        \SUBBYTES[0].a/n1602 ), .Z(\SUBBYTES[0].a/w581 ) );
  XOR \SUBBYTES[0].a/U4079  ( .A(\SUBBYTES[0].a/n1602 ), .B(
        \SUBBYTES[0].a/n1314 ), .Z(\SUBBYTES[0].a/w666 ) );
  XOR \SUBBYTES[0].a/U4078  ( .A(\w1[0][108] ), .B(\w1[0][105] ), .Z(
        \SUBBYTES[0].a/n1314 ) );
  XOR \SUBBYTES[0].a/U4077  ( .A(\SUBBYTES[0].a/n1316 ), .B(
        \SUBBYTES[0].a/n1315 ), .Z(\SUBBYTES[0].a/n1599 ) );
  XOR \SUBBYTES[0].a/U4076  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/n1317 ), .Z(
        \SUBBYTES[0].a/n1315 ) );
  XOR \SUBBYTES[0].a/U4075  ( .A(\SUBBYTES[0].a/w631 ), .B(\w1[0][110] ), .Z(
        \SUBBYTES[0].a/n1316 ) );
  XOR \SUBBYTES[0].a/U4074  ( .A(\SUBBYTES[0].a/w605 ), .B(
        \SUBBYTES[0].a/w612 ), .Z(\SUBBYTES[0].a/n1317 ) );
  XOR \SUBBYTES[0].a/U4073  ( .A(\SUBBYTES[0].a/n1319 ), .B(
        \SUBBYTES[0].a/n1318 ), .Z(\SUBBYTES[0].a/n1597 ) );
  XOR \SUBBYTES[0].a/U4072  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1320 ), .Z(
        \SUBBYTES[0].a/n1318 ) );
  XOR \SUBBYTES[0].a/U4071  ( .A(\SUBBYTES[0].a/w630 ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1319 ) );
  XOR \SUBBYTES[0].a/U4070  ( .A(\SUBBYTES[0].a/w606 ), .B(
        \SUBBYTES[0].a/w613 ), .Z(\SUBBYTES[0].a/n1320 ) );
  XOR \SUBBYTES[0].a/U4069  ( .A(\SUBBYTES[0].a/n1599 ), .B(
        \SUBBYTES[0].a/n1597 ), .Z(\SUBBYTES[0].a/w636 ) );
  XOR \SUBBYTES[0].a/U4068  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1321 ), .Z(
        \SUBBYTES[0].a/n1600 ) );
  XOR \SUBBYTES[0].a/U4067  ( .A(\SUBBYTES[0].a/w598 ), .B(
        \SUBBYTES[0].a/w608 ), .Z(\SUBBYTES[0].a/n1321 ) );
  XOR \SUBBYTES[0].a/U4066  ( .A(\SUBBYTES[0].a/n1323 ), .B(
        \SUBBYTES[0].a/n1322 ), .Z(\SUBBYTES[0].a/w623 ) );
  XOR \SUBBYTES[0].a/U4065  ( .A(\SUBBYTES[0].a/n1600 ), .B(
        \SUBBYTES[0].a/n1324 ), .Z(\SUBBYTES[0].a/n1322 ) );
  XOR \SUBBYTES[0].a/U4064  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/n1323 ) );
  XOR \SUBBYTES[0].a/U4063  ( .A(\SUBBYTES[0].a/w600 ), .B(
        \SUBBYTES[0].a/w605 ), .Z(\SUBBYTES[0].a/n1324 ) );
  XOR \SUBBYTES[0].a/U4062  ( .A(\SUBBYTES[0].a/n1326 ), .B(
        \SUBBYTES[0].a/n1325 ), .Z(\SUBBYTES[0].a/n1598 ) );
  XOR \SUBBYTES[0].a/U4061  ( .A(\SUBBYTES[0].a/w633 ), .B(\w1[0][111] ), .Z(
        \SUBBYTES[0].a/n1325 ) );
  XOR \SUBBYTES[0].a/U4060  ( .A(\SUBBYTES[0].a/w608 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1326 ) );
  XOR \SUBBYTES[0].a/U4059  ( .A(\SUBBYTES[0].a/n1597 ), .B(
        \SUBBYTES[0].a/n1598 ), .Z(\SUBBYTES[0].a/w635 ) );
  XOR \SUBBYTES[0].a/U4058  ( .A(\w1[0][107] ), .B(\SUBBYTES[0].a/n1327 ), .Z(
        \SUBBYTES[0].a/n1601 ) );
  XOR \SUBBYTES[0].a/U4057  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w600 ), .Z(\SUBBYTES[0].a/n1327 ) );
  XOR \SUBBYTES[0].a/U4056  ( .A(\SUBBYTES[0].a/n1329 ), .B(
        \SUBBYTES[0].a/n1328 ), .Z(\SUBBYTES[0].a/w624 ) );
  XOR \SUBBYTES[0].a/U4055  ( .A(\SUBBYTES[0].a/n1601 ), .B(
        \SUBBYTES[0].a/n1330 ), .Z(\SUBBYTES[0].a/n1328 ) );
  XOR \SUBBYTES[0].a/U4054  ( .A(\w1[0][110] ), .B(\SUBBYTES[0].a/w666 ), .Z(
        \SUBBYTES[0].a/n1329 ) );
  XOR \SUBBYTES[0].a/U4053  ( .A(\SUBBYTES[0].a/w605 ), .B(
        \SUBBYTES[0].a/w606 ), .Z(\SUBBYTES[0].a/n1330 ) );
  XOR \SUBBYTES[0].a/U4052  ( .A(\SUBBYTES[0].a/n1599 ), .B(
        \SUBBYTES[0].a/n1598 ), .Z(\SUBBYTES[0].a/w644 ) );
  XOR \SUBBYTES[0].a/U4051  ( .A(\SUBBYTES[0].a/n1332 ), .B(
        \SUBBYTES[0].a/n1331 ), .Z(\SUBBYTES[0].a/w645 ) );
  XOR \SUBBYTES[0].a/U4050  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/n1600 ), .Z(
        \SUBBYTES[0].a/n1331 ) );
  XOR \SUBBYTES[0].a/U4049  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w606 ), .Z(\SUBBYTES[0].a/n1332 ) );
  XOR \SUBBYTES[0].a/U4048  ( .A(\SUBBYTES[0].a/n1334 ), .B(
        \SUBBYTES[0].a/n1333 ), .Z(\SUBBYTES[0].a/w621 ) );
  XOR \SUBBYTES[0].a/U4047  ( .A(\SUBBYTES[0].a/n1336 ), .B(
        \SUBBYTES[0].a/n1335 ), .Z(\SUBBYTES[0].a/n1333 ) );
  XOR \SUBBYTES[0].a/U4046  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/w705 ), .Z(
        \SUBBYTES[0].a/n1334 ) );
  XOR \SUBBYTES[0].a/U4045  ( .A(\SUBBYTES[0].a/w612 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1335 ) );
  XOR \SUBBYTES[0].a/U4044  ( .A(\SUBBYTES[0].a/w598 ), .B(
        \SUBBYTES[0].a/w600 ), .Z(\SUBBYTES[0].a/n1336 ) );
  XOR \SUBBYTES[0].a/U4043  ( .A(\SUBBYTES[0].a/n1338 ), .B(
        \SUBBYTES[0].a/n1337 ), .Z(\SUBBYTES[0].a/w622 ) );
  XOR \SUBBYTES[0].a/U4042  ( .A(\SUBBYTES[0].a/n1601 ), .B(
        \SUBBYTES[0].a/n1339 ), .Z(\SUBBYTES[0].a/n1337 ) );
  XOR \SUBBYTES[0].a/U4041  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1602 ), .Z(
        \SUBBYTES[0].a/n1338 ) );
  XOR \SUBBYTES[0].a/U4040  ( .A(\SUBBYTES[0].a/w612 ), .B(
        \SUBBYTES[0].a/w613 ), .Z(\SUBBYTES[0].a/n1339 ) );
  XOR \SUBBYTES[0].a/U4039  ( .A(\SUBBYTES[0].a/n1341 ), .B(
        \SUBBYTES[0].a/n1340 ), .Z(\SUBBYTES[0].a/w638 ) );
  XOR \SUBBYTES[0].a/U4038  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1342 ), .Z(
        \SUBBYTES[0].a/n1340 ) );
  XOR \SUBBYTES[0].a/U4037  ( .A(\SUBBYTES[0].a/w613 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1341 ) );
  XOR \SUBBYTES[0].a/U4036  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w598 ), .Z(\SUBBYTES[0].a/n1342 ) );
  XOR \SUBBYTES[0].a/U4035  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1343 ), .Z(
        \SUBBYTES[0].a/n1603 ) );
  XOR \SUBBYTES[0].a/U4034  ( .A(\w1[0][115] ), .B(\w1[0][114] ), .Z(
        \SUBBYTES[0].a/n1343 ) );
  XOR \SUBBYTES[0].a/U4033  ( .A(\w1[0][118] ), .B(\SUBBYTES[0].a/n1603 ), .Z(
        \SUBBYTES[0].a/w480 ) );
  XOR \SUBBYTES[0].a/U4032  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/w367 ) );
  XOR \SUBBYTES[0].a/U4031  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/n1344 ), .Z(
        \SUBBYTES[0].a/w368 ) );
  XOR \SUBBYTES[0].a/U4030  ( .A(\w1[0][118] ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1344 ) );
  XOR \SUBBYTES[0].a/U4029  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1603 ), .Z(
        \SUBBYTES[0].a/w498 ) );
  XOR \SUBBYTES[0].a/U4028  ( .A(\SUBBYTES[0].a/n1346 ), .B(
        \SUBBYTES[0].a/n1345 ), .Z(\SUBBYTES[0].a/w491 ) );
  XOR \SUBBYTES[0].a/U4027  ( .A(\w1[0][115] ), .B(\w1[0][113] ), .Z(
        \SUBBYTES[0].a/n1345 ) );
  XOR \SUBBYTES[0].a/U4026  ( .A(\w1[0][119] ), .B(\w1[0][116] ), .Z(
        \SUBBYTES[0].a/n1346 ) );
  XOR \SUBBYTES[0].a/U4025  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w491 ), .Z(
        \SUBBYTES[0].a/w370 ) );
  XOR \SUBBYTES[0].a/U4024  ( .A(\SUBBYTES[0].a/n1348 ), .B(
        \SUBBYTES[0].a/n1347 ), .Z(\SUBBYTES[0].a/w478 ) );
  XOR \SUBBYTES[0].a/U4023  ( .A(\SUBBYTES[0].a/w439 ), .B(n2), .Z(
        \SUBBYTES[0].a/n1347 ) );
  XOR \SUBBYTES[0].a/U4022  ( .A(\SUBBYTES[0].a/w432 ), .B(
        \SUBBYTES[0].a/w435 ), .Z(\SUBBYTES[0].a/n1348 ) );
  XOR \SUBBYTES[0].a/U4021  ( .A(\SUBBYTES[0].a/n1350 ), .B(
        \SUBBYTES[0].a/n1349 ), .Z(\SUBBYTES[0].a/w479 ) );
  XOR \SUBBYTES[0].a/U4020  ( .A(\SUBBYTES[0].a/w439 ), .B(\SUBBYTES[0].a/n20 ), .Z(\SUBBYTES[0].a/n1349 ) );
  XOR \SUBBYTES[0].a/U4019  ( .A(\SUBBYTES[0].a/w432 ), .B(\SUBBYTES[0].a/n19 ), .Z(\SUBBYTES[0].a/n1350 ) );
  XOR \SUBBYTES[0].a/U4018  ( .A(\SUBBYTES[0].a/w491 ), .B(
        \SUBBYTES[0].a/n1351 ), .Z(\SUBBYTES[0].a/w481 ) );
  XOR \SUBBYTES[0].a/U4017  ( .A(\w1[0][118] ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1351 ) );
  XOR \SUBBYTES[0].a/U4016  ( .A(\SUBBYTES[0].a/n1353 ), .B(
        \SUBBYTES[0].a/n1352 ), .Z(\SUBBYTES[0].a/w482 ) );
  XOR \SUBBYTES[0].a/U4015  ( .A(\SUBBYTES[0].a/n20 ), .B(n2), .Z(
        \SUBBYTES[0].a/n1352 ) );
  XOR \SUBBYTES[0].a/U4014  ( .A(\SUBBYTES[0].a/n19 ), .B(\SUBBYTES[0].a/w435 ), .Z(\SUBBYTES[0].a/n1353 ) );
  XOR \SUBBYTES[0].a/U4013  ( .A(\w1[0][119] ), .B(\w1[0][114] ), .Z(
        \SUBBYTES[0].a/n1609 ) );
  XOR \SUBBYTES[0].a/U4012  ( .A(\SUBBYTES[0].a/n1609 ), .B(
        \SUBBYTES[0].a/n1354 ), .Z(\SUBBYTES[0].a/w483 ) );
  XOR \SUBBYTES[0].a/U4011  ( .A(\w1[0][117] ), .B(\w1[0][116] ), .Z(
        \SUBBYTES[0].a/n1354 ) );
  XOR \SUBBYTES[0].a/U4010  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w371 ) );
  XOR \SUBBYTES[0].a/U4009  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w372 ) );
  XOR \SUBBYTES[0].a/U4008  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w373 ) );
  XOR \SUBBYTES[0].a/U4007  ( .A(\SUBBYTES[0].a/w372 ), .B(
        \SUBBYTES[0].a/n1609 ), .Z(\SUBBYTES[0].a/w374 ) );
  XOR \SUBBYTES[0].a/U4006  ( .A(\SUBBYTES[0].a/n1609 ), .B(
        \SUBBYTES[0].a/n1355 ), .Z(\SUBBYTES[0].a/w459 ) );
  XOR \SUBBYTES[0].a/U4005  ( .A(\w1[0][116] ), .B(\w1[0][113] ), .Z(
        \SUBBYTES[0].a/n1355 ) );
  XOR \SUBBYTES[0].a/U4004  ( .A(\SUBBYTES[0].a/n1357 ), .B(
        \SUBBYTES[0].a/n1356 ), .Z(\SUBBYTES[0].a/n1606 ) );
  XOR \SUBBYTES[0].a/U4003  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/n1358 ), .Z(
        \SUBBYTES[0].a/n1356 ) );
  XOR \SUBBYTES[0].a/U4002  ( .A(\SUBBYTES[0].a/w424 ), .B(\w1[0][118] ), .Z(
        \SUBBYTES[0].a/n1357 ) );
  XOR \SUBBYTES[0].a/U4001  ( .A(\SUBBYTES[0].a/w398 ), .B(
        \SUBBYTES[0].a/w405 ), .Z(\SUBBYTES[0].a/n1358 ) );
  XOR \SUBBYTES[0].a/U4000  ( .A(\SUBBYTES[0].a/n1360 ), .B(
        \SUBBYTES[0].a/n1359 ), .Z(\SUBBYTES[0].a/n1604 ) );
  XOR \SUBBYTES[0].a/U3999  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1361 ), .Z(
        \SUBBYTES[0].a/n1359 ) );
  XOR \SUBBYTES[0].a/U3998  ( .A(\SUBBYTES[0].a/w423 ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1360 ) );
  XOR \SUBBYTES[0].a/U3997  ( .A(\SUBBYTES[0].a/w399 ), .B(
        \SUBBYTES[0].a/w406 ), .Z(\SUBBYTES[0].a/n1361 ) );
  XOR \SUBBYTES[0].a/U3996  ( .A(\SUBBYTES[0].a/n1606 ), .B(
        \SUBBYTES[0].a/n1604 ), .Z(\SUBBYTES[0].a/w429 ) );
  XOR \SUBBYTES[0].a/U3995  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1362 ), .Z(
        \SUBBYTES[0].a/n1607 ) );
  XOR \SUBBYTES[0].a/U3994  ( .A(\SUBBYTES[0].a/w391 ), .B(
        \SUBBYTES[0].a/w401 ), .Z(\SUBBYTES[0].a/n1362 ) );
  XOR \SUBBYTES[0].a/U3993  ( .A(\SUBBYTES[0].a/n1364 ), .B(
        \SUBBYTES[0].a/n1363 ), .Z(\SUBBYTES[0].a/w416 ) );
  XOR \SUBBYTES[0].a/U3992  ( .A(\SUBBYTES[0].a/n1607 ), .B(
        \SUBBYTES[0].a/n1365 ), .Z(\SUBBYTES[0].a/n1363 ) );
  XOR \SUBBYTES[0].a/U3991  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/n1364 ) );
  XOR \SUBBYTES[0].a/U3990  ( .A(\SUBBYTES[0].a/w393 ), .B(
        \SUBBYTES[0].a/w398 ), .Z(\SUBBYTES[0].a/n1365 ) );
  XOR \SUBBYTES[0].a/U3989  ( .A(\SUBBYTES[0].a/n1367 ), .B(
        \SUBBYTES[0].a/n1366 ), .Z(\SUBBYTES[0].a/n1605 ) );
  XOR \SUBBYTES[0].a/U3988  ( .A(\SUBBYTES[0].a/w426 ), .B(\w1[0][119] ), .Z(
        \SUBBYTES[0].a/n1366 ) );
  XOR \SUBBYTES[0].a/U3987  ( .A(\SUBBYTES[0].a/w401 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1367 ) );
  XOR \SUBBYTES[0].a/U3986  ( .A(\SUBBYTES[0].a/n1604 ), .B(
        \SUBBYTES[0].a/n1605 ), .Z(\SUBBYTES[0].a/w428 ) );
  XOR \SUBBYTES[0].a/U3985  ( .A(\w1[0][115] ), .B(\SUBBYTES[0].a/n1368 ), .Z(
        \SUBBYTES[0].a/n1608 ) );
  XOR \SUBBYTES[0].a/U3984  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w393 ), .Z(\SUBBYTES[0].a/n1368 ) );
  XOR \SUBBYTES[0].a/U3983  ( .A(\SUBBYTES[0].a/n1370 ), .B(
        \SUBBYTES[0].a/n1369 ), .Z(\SUBBYTES[0].a/w417 ) );
  XOR \SUBBYTES[0].a/U3982  ( .A(\SUBBYTES[0].a/n1608 ), .B(
        \SUBBYTES[0].a/n1371 ), .Z(\SUBBYTES[0].a/n1369 ) );
  XOR \SUBBYTES[0].a/U3981  ( .A(\w1[0][118] ), .B(\SUBBYTES[0].a/w459 ), .Z(
        \SUBBYTES[0].a/n1370 ) );
  XOR \SUBBYTES[0].a/U3980  ( .A(\SUBBYTES[0].a/w398 ), .B(
        \SUBBYTES[0].a/w399 ), .Z(\SUBBYTES[0].a/n1371 ) );
  XOR \SUBBYTES[0].a/U3979  ( .A(\SUBBYTES[0].a/n1606 ), .B(
        \SUBBYTES[0].a/n1605 ), .Z(\SUBBYTES[0].a/w437 ) );
  XOR \SUBBYTES[0].a/U3978  ( .A(\SUBBYTES[0].a/n1373 ), .B(
        \SUBBYTES[0].a/n1372 ), .Z(\SUBBYTES[0].a/w438 ) );
  XOR \SUBBYTES[0].a/U3977  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/n1607 ), .Z(
        \SUBBYTES[0].a/n1372 ) );
  XOR \SUBBYTES[0].a/U3976  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w399 ), .Z(\SUBBYTES[0].a/n1373 ) );
  XOR \SUBBYTES[0].a/U3975  ( .A(\SUBBYTES[0].a/n1375 ), .B(
        \SUBBYTES[0].a/n1374 ), .Z(\SUBBYTES[0].a/w414 ) );
  XOR \SUBBYTES[0].a/U3974  ( .A(\SUBBYTES[0].a/n1377 ), .B(
        \SUBBYTES[0].a/n1376 ), .Z(\SUBBYTES[0].a/n1374 ) );
  XOR \SUBBYTES[0].a/U3973  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/w498 ), .Z(
        \SUBBYTES[0].a/n1375 ) );
  XOR \SUBBYTES[0].a/U3972  ( .A(\SUBBYTES[0].a/w405 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1376 ) );
  XOR \SUBBYTES[0].a/U3971  ( .A(\SUBBYTES[0].a/w391 ), .B(
        \SUBBYTES[0].a/w393 ), .Z(\SUBBYTES[0].a/n1377 ) );
  XOR \SUBBYTES[0].a/U3970  ( .A(\SUBBYTES[0].a/n1379 ), .B(
        \SUBBYTES[0].a/n1378 ), .Z(\SUBBYTES[0].a/w415 ) );
  XOR \SUBBYTES[0].a/U3969  ( .A(\SUBBYTES[0].a/n1608 ), .B(
        \SUBBYTES[0].a/n1380 ), .Z(\SUBBYTES[0].a/n1378 ) );
  XOR \SUBBYTES[0].a/U3968  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1609 ), .Z(
        \SUBBYTES[0].a/n1379 ) );
  XOR \SUBBYTES[0].a/U3967  ( .A(\SUBBYTES[0].a/w405 ), .B(
        \SUBBYTES[0].a/w406 ), .Z(\SUBBYTES[0].a/n1380 ) );
  XOR \SUBBYTES[0].a/U3966  ( .A(\SUBBYTES[0].a/n1382 ), .B(
        \SUBBYTES[0].a/n1381 ), .Z(\SUBBYTES[0].a/w431 ) );
  XOR \SUBBYTES[0].a/U3965  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1383 ), .Z(
        \SUBBYTES[0].a/n1381 ) );
  XOR \SUBBYTES[0].a/U3964  ( .A(\SUBBYTES[0].a/w406 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1382 ) );
  XOR \SUBBYTES[0].a/U3963  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w391 ), .Z(\SUBBYTES[0].a/n1383 ) );
  XOR \SUBBYTES[0].a/U3962  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1384 ), .Z(
        \SUBBYTES[0].a/n1610 ) );
  XOR \SUBBYTES[0].a/U3961  ( .A(\w1[0][123] ), .B(\w1[0][122] ), .Z(
        \SUBBYTES[0].a/n1384 ) );
  XOR \SUBBYTES[0].a/U3960  ( .A(\w1[0][126] ), .B(\SUBBYTES[0].a/n1610 ), .Z(
        \SUBBYTES[0].a/w273 ) );
  XOR \SUBBYTES[0].a/U3959  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/w160 ) );
  XOR \SUBBYTES[0].a/U3958  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/n1385 ), .Z(
        \SUBBYTES[0].a/w161 ) );
  XOR \SUBBYTES[0].a/U3957  ( .A(\w1[0][126] ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1385 ) );
  XOR \SUBBYTES[0].a/U3956  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1610 ), .Z(
        \SUBBYTES[0].a/w291 ) );
  XOR \SUBBYTES[0].a/U3955  ( .A(\SUBBYTES[0].a/n1387 ), .B(
        \SUBBYTES[0].a/n1386 ), .Z(\SUBBYTES[0].a/w284 ) );
  XOR \SUBBYTES[0].a/U3954  ( .A(\w1[0][123] ), .B(\w1[0][121] ), .Z(
        \SUBBYTES[0].a/n1386 ) );
  XOR \SUBBYTES[0].a/U3953  ( .A(\w1[0][127] ), .B(\w1[0][124] ), .Z(
        \SUBBYTES[0].a/n1387 ) );
  XOR \SUBBYTES[0].a/U3952  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w284 ), .Z(
        \SUBBYTES[0].a/w163 ) );
  XOR \SUBBYTES[0].a/U3951  ( .A(\SUBBYTES[0].a/n1389 ), .B(
        \SUBBYTES[0].a/n1388 ), .Z(\SUBBYTES[0].a/w271 ) );
  XOR \SUBBYTES[0].a/U3950  ( .A(\SUBBYTES[0].a/w232 ), .B(n1), .Z(
        \SUBBYTES[0].a/n1388 ) );
  XOR \SUBBYTES[0].a/U3949  ( .A(\SUBBYTES[0].a/w225 ), .B(
        \SUBBYTES[0].a/w228 ), .Z(\SUBBYTES[0].a/n1389 ) );
  XOR \SUBBYTES[0].a/U3948  ( .A(\SUBBYTES[0].a/n1391 ), .B(
        \SUBBYTES[0].a/n1390 ), .Z(\SUBBYTES[0].a/w272 ) );
  XOR \SUBBYTES[0].a/U3947  ( .A(\SUBBYTES[0].a/w232 ), .B(\SUBBYTES[0].a/n10 ), .Z(\SUBBYTES[0].a/n1390 ) );
  XOR \SUBBYTES[0].a/U3946  ( .A(\SUBBYTES[0].a/w225 ), .B(\SUBBYTES[0].a/n9 ), 
        .Z(\SUBBYTES[0].a/n1391 ) );
  XOR \SUBBYTES[0].a/U3945  ( .A(\SUBBYTES[0].a/w284 ), .B(
        \SUBBYTES[0].a/n1392 ), .Z(\SUBBYTES[0].a/w274 ) );
  XOR \SUBBYTES[0].a/U3944  ( .A(\w1[0][126] ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1392 ) );
  XOR \SUBBYTES[0].a/U3943  ( .A(\SUBBYTES[0].a/n1394 ), .B(
        \SUBBYTES[0].a/n1393 ), .Z(\SUBBYTES[0].a/w275 ) );
  XOR \SUBBYTES[0].a/U3942  ( .A(\SUBBYTES[0].a/n10 ), .B(n1), .Z(
        \SUBBYTES[0].a/n1393 ) );
  XOR \SUBBYTES[0].a/U3941  ( .A(\SUBBYTES[0].a/n9 ), .B(\SUBBYTES[0].a/w228 ), 
        .Z(\SUBBYTES[0].a/n1394 ) );
  XOR \SUBBYTES[0].a/U3940  ( .A(\w1[0][127] ), .B(\w1[0][122] ), .Z(
        \SUBBYTES[0].a/n1616 ) );
  XOR \SUBBYTES[0].a/U3939  ( .A(\SUBBYTES[0].a/n1616 ), .B(
        \SUBBYTES[0].a/n1395 ), .Z(\SUBBYTES[0].a/w276 ) );
  XOR \SUBBYTES[0].a/U3938  ( .A(\w1[0][125] ), .B(\w1[0][124] ), .Z(
        \SUBBYTES[0].a/n1395 ) );
  XOR \SUBBYTES[0].a/U3937  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w164 ) );
  XOR \SUBBYTES[0].a/U3936  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w165 ) );
  XOR \SUBBYTES[0].a/U3935  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w166 ) );
  XOR \SUBBYTES[0].a/U3934  ( .A(\SUBBYTES[0].a/w165 ), .B(
        \SUBBYTES[0].a/n1616 ), .Z(\SUBBYTES[0].a/w167 ) );
  XOR \SUBBYTES[0].a/U3933  ( .A(\SUBBYTES[0].a/n1616 ), .B(
        \SUBBYTES[0].a/n1396 ), .Z(\SUBBYTES[0].a/w252 ) );
  XOR \SUBBYTES[0].a/U3932  ( .A(\w1[0][124] ), .B(\w1[0][121] ), .Z(
        \SUBBYTES[0].a/n1396 ) );
  XOR \SUBBYTES[0].a/U3931  ( .A(\SUBBYTES[0].a/n1398 ), .B(
        \SUBBYTES[0].a/n1397 ), .Z(\SUBBYTES[0].a/n1613 ) );
  XOR \SUBBYTES[0].a/U3930  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/n1399 ), .Z(
        \SUBBYTES[0].a/n1397 ) );
  XOR \SUBBYTES[0].a/U3929  ( .A(\SUBBYTES[0].a/w217 ), .B(\w1[0][126] ), .Z(
        \SUBBYTES[0].a/n1398 ) );
  XOR \SUBBYTES[0].a/U3928  ( .A(\SUBBYTES[0].a/w191 ), .B(
        \SUBBYTES[0].a/w198 ), .Z(\SUBBYTES[0].a/n1399 ) );
  XOR \SUBBYTES[0].a/U3927  ( .A(\SUBBYTES[0].a/n1401 ), .B(
        \SUBBYTES[0].a/n1400 ), .Z(\SUBBYTES[0].a/n1611 ) );
  XOR \SUBBYTES[0].a/U3926  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1402 ), .Z(
        \SUBBYTES[0].a/n1400 ) );
  XOR \SUBBYTES[0].a/U3925  ( .A(\SUBBYTES[0].a/w216 ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1401 ) );
  XOR \SUBBYTES[0].a/U3924  ( .A(\SUBBYTES[0].a/w192 ), .B(
        \SUBBYTES[0].a/w199 ), .Z(\SUBBYTES[0].a/n1402 ) );
  XOR \SUBBYTES[0].a/U3923  ( .A(\SUBBYTES[0].a/n1613 ), .B(
        \SUBBYTES[0].a/n1611 ), .Z(\SUBBYTES[0].a/w222 ) );
  XOR \SUBBYTES[0].a/U3922  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1403 ), .Z(
        \SUBBYTES[0].a/n1614 ) );
  XOR \SUBBYTES[0].a/U3921  ( .A(\SUBBYTES[0].a/w184 ), .B(
        \SUBBYTES[0].a/w194 ), .Z(\SUBBYTES[0].a/n1403 ) );
  XOR \SUBBYTES[0].a/U3920  ( .A(\SUBBYTES[0].a/n1405 ), .B(
        \SUBBYTES[0].a/n1404 ), .Z(\SUBBYTES[0].a/w209 ) );
  XOR \SUBBYTES[0].a/U3919  ( .A(\SUBBYTES[0].a/n1614 ), .B(
        \SUBBYTES[0].a/n1406 ), .Z(\SUBBYTES[0].a/n1404 ) );
  XOR \SUBBYTES[0].a/U3918  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/n1405 ) );
  XOR \SUBBYTES[0].a/U3917  ( .A(\SUBBYTES[0].a/w186 ), .B(
        \SUBBYTES[0].a/w191 ), .Z(\SUBBYTES[0].a/n1406 ) );
  XOR \SUBBYTES[0].a/U3916  ( .A(\SUBBYTES[0].a/n1408 ), .B(
        \SUBBYTES[0].a/n1407 ), .Z(\SUBBYTES[0].a/n1612 ) );
  XOR \SUBBYTES[0].a/U3915  ( .A(\SUBBYTES[0].a/w219 ), .B(\w1[0][127] ), .Z(
        \SUBBYTES[0].a/n1407 ) );
  XOR \SUBBYTES[0].a/U3914  ( .A(\SUBBYTES[0].a/w194 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1408 ) );
  XOR \SUBBYTES[0].a/U3913  ( .A(\SUBBYTES[0].a/n1611 ), .B(
        \SUBBYTES[0].a/n1612 ), .Z(\SUBBYTES[0].a/w221 ) );
  XOR \SUBBYTES[0].a/U3912  ( .A(\w1[0][123] ), .B(\SUBBYTES[0].a/n1409 ), .Z(
        \SUBBYTES[0].a/n1615 ) );
  XOR \SUBBYTES[0].a/U3911  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w186 ), .Z(\SUBBYTES[0].a/n1409 ) );
  XOR \SUBBYTES[0].a/U3910  ( .A(\SUBBYTES[0].a/n1411 ), .B(
        \SUBBYTES[0].a/n1410 ), .Z(\SUBBYTES[0].a/w210 ) );
  XOR \SUBBYTES[0].a/U3909  ( .A(\SUBBYTES[0].a/n1615 ), .B(
        \SUBBYTES[0].a/n1412 ), .Z(\SUBBYTES[0].a/n1410 ) );
  XOR \SUBBYTES[0].a/U3908  ( .A(\w1[0][126] ), .B(\SUBBYTES[0].a/w252 ), .Z(
        \SUBBYTES[0].a/n1411 ) );
  XOR \SUBBYTES[0].a/U3907  ( .A(\SUBBYTES[0].a/w191 ), .B(
        \SUBBYTES[0].a/w192 ), .Z(\SUBBYTES[0].a/n1412 ) );
  XOR \SUBBYTES[0].a/U3906  ( .A(\SUBBYTES[0].a/n1613 ), .B(
        \SUBBYTES[0].a/n1612 ), .Z(\SUBBYTES[0].a/w230 ) );
  XOR \SUBBYTES[0].a/U3905  ( .A(\SUBBYTES[0].a/n1414 ), .B(
        \SUBBYTES[0].a/n1413 ), .Z(\SUBBYTES[0].a/w231 ) );
  XOR \SUBBYTES[0].a/U3904  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/n1614 ), .Z(
        \SUBBYTES[0].a/n1413 ) );
  XOR \SUBBYTES[0].a/U3903  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w192 ), .Z(\SUBBYTES[0].a/n1414 ) );
  XOR \SUBBYTES[0].a/U3902  ( .A(\SUBBYTES[0].a/n1416 ), .B(
        \SUBBYTES[0].a/n1415 ), .Z(\SUBBYTES[0].a/w207 ) );
  XOR \SUBBYTES[0].a/U3901  ( .A(\SUBBYTES[0].a/n1418 ), .B(
        \SUBBYTES[0].a/n1417 ), .Z(\SUBBYTES[0].a/n1415 ) );
  XOR \SUBBYTES[0].a/U3900  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/w291 ), .Z(
        \SUBBYTES[0].a/n1416 ) );
  XOR \SUBBYTES[0].a/U3899  ( .A(\SUBBYTES[0].a/w198 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1417 ) );
  XOR \SUBBYTES[0].a/U3898  ( .A(\SUBBYTES[0].a/w184 ), .B(
        \SUBBYTES[0].a/w186 ), .Z(\SUBBYTES[0].a/n1418 ) );
  XOR \SUBBYTES[0].a/U3897  ( .A(\SUBBYTES[0].a/n1420 ), .B(
        \SUBBYTES[0].a/n1419 ), .Z(\SUBBYTES[0].a/w208 ) );
  XOR \SUBBYTES[0].a/U3896  ( .A(\SUBBYTES[0].a/n1615 ), .B(
        \SUBBYTES[0].a/n1421 ), .Z(\SUBBYTES[0].a/n1419 ) );
  XOR \SUBBYTES[0].a/U3895  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1616 ), .Z(
        \SUBBYTES[0].a/n1420 ) );
  XOR \SUBBYTES[0].a/U3894  ( .A(\SUBBYTES[0].a/w198 ), .B(
        \SUBBYTES[0].a/w199 ), .Z(\SUBBYTES[0].a/n1421 ) );
  XOR \SUBBYTES[0].a/U3893  ( .A(\SUBBYTES[0].a/n1423 ), .B(
        \SUBBYTES[0].a/n1422 ), .Z(\SUBBYTES[0].a/w224 ) );
  XOR \SUBBYTES[0].a/U3892  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1424 ), .Z(
        \SUBBYTES[0].a/n1422 ) );
  XOR \SUBBYTES[0].a/U3891  ( .A(\SUBBYTES[0].a/w199 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1423 ) );
  XOR \SUBBYTES[0].a/U3890  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w184 ), .Z(\SUBBYTES[0].a/n1424 ) );
  AND U4 ( .A(\SUBBYTES[0].a/w209 ), .B(\SUBBYTES[0].a/w222 ), .Z(n1) );
  AND U5 ( .A(\SUBBYTES[0].a/w416 ), .B(\SUBBYTES[0].a/w429 ), .Z(n2) );
  AND U6 ( .A(\SUBBYTES[0].a/w623 ), .B(\SUBBYTES[0].a/w636 ), .Z(n3) );
  AND U7 ( .A(\SUBBYTES[0].a/w830 ), .B(\SUBBYTES[0].a/w843 ), .Z(n4) );
  AND U8 ( .A(\SUBBYTES[0].a/w1037 ), .B(\SUBBYTES[0].a/w1050 ), .Z(n5) );
  AND U9 ( .A(\SUBBYTES[0].a/w1244 ), .B(\SUBBYTES[0].a/w1257 ), .Z(n6) );
  AND U10 ( .A(\SUBBYTES[0].a/w1451 ), .B(\SUBBYTES[0].a/w1464 ), .Z(n7) );
  AND U11 ( .A(\SUBBYTES[0].a/w1658 ), .B(\SUBBYTES[0].a/w1671 ), .Z(n8) );
  AND U12 ( .A(\SUBBYTES[0].a/w1865 ), .B(\SUBBYTES[0].a/w1878 ), .Z(n9) );
  AND U13 ( .A(\SUBBYTES[0].a/w2072 ), .B(\SUBBYTES[0].a/w2085 ), .Z(n10) );
  AND U14 ( .A(\SUBBYTES[0].a/w2279 ), .B(\SUBBYTES[0].a/w2292 ), .Z(n11) );
  AND U15 ( .A(\SUBBYTES[0].a/w2486 ), .B(\SUBBYTES[0].a/w2499 ), .Z(n12) );
  AND U16 ( .A(\SUBBYTES[0].a/w2693 ), .B(\SUBBYTES[0].a/w2706 ), .Z(n13) );
  AND U17 ( .A(\SUBBYTES[0].a/w2900 ), .B(\SUBBYTES[0].a/w2913 ), .Z(n14) );
  AND U18 ( .A(\SUBBYTES[0].a/w3107 ), .B(\SUBBYTES[0].a/w3120 ), .Z(n15) );
  AND U19 ( .A(\SUBBYTES[0].a/w3314 ), .B(\SUBBYTES[0].a/w3327 ), .Z(n16) );
  XOR U20 ( .A(state[99]), .B(g_input[99]), .Z(\w1[0][99] ) );
  XOR U21 ( .A(state[94]), .B(g_input[94]), .Z(\w1[0][94] ) );
  XOR U22 ( .A(state[93]), .B(g_input[93]), .Z(\w1[0][93] ) );
  XOR U23 ( .A(state[91]), .B(g_input[91]), .Z(\w1[0][91] ) );
  XOR U24 ( .A(state[86]), .B(g_input[86]), .Z(\w1[0][86] ) );
  XOR U25 ( .A(state[85]), .B(g_input[85]), .Z(\w1[0][85] ) );
  XOR U26 ( .A(state[83]), .B(g_input[83]), .Z(\w1[0][83] ) );
  XOR U27 ( .A(state[78]), .B(g_input[78]), .Z(\w1[0][78] ) );
  XOR U28 ( .A(state[77]), .B(g_input[77]), .Z(\w1[0][77] ) );
  XOR U29 ( .A(state[75]), .B(g_input[75]), .Z(\w1[0][75] ) );
  XOR U30 ( .A(state[70]), .B(g_input[70]), .Z(\w1[0][70] ) );
  XOR U31 ( .A(state[6]), .B(g_input[6]), .Z(\w1[0][6] ) );
  XOR U32 ( .A(state[69]), .B(g_input[69]), .Z(\w1[0][69] ) );
  XOR U33 ( .A(state[67]), .B(g_input[67]), .Z(\w1[0][67] ) );
  XOR U34 ( .A(state[62]), .B(g_input[62]), .Z(\w1[0][62] ) );
  XOR U35 ( .A(state[61]), .B(g_input[61]), .Z(\w1[0][61] ) );
  XOR U36 ( .A(state[5]), .B(g_input[5]), .Z(\w1[0][5] ) );
  XOR U37 ( .A(state[59]), .B(g_input[59]), .Z(\w1[0][59] ) );
  XOR U38 ( .A(state[54]), .B(g_input[54]), .Z(\w1[0][54] ) );
  XOR U39 ( .A(state[53]), .B(g_input[53]), .Z(\w1[0][53] ) );
  XOR U40 ( .A(state[51]), .B(g_input[51]), .Z(\w1[0][51] ) );
  XOR U41 ( .A(state[46]), .B(g_input[46]), .Z(\w1[0][46] ) );
  XOR U42 ( .A(state[45]), .B(g_input[45]), .Z(\w1[0][45] ) );
  XOR U43 ( .A(state[43]), .B(g_input[43]), .Z(\w1[0][43] ) );
  XOR U44 ( .A(state[3]), .B(g_input[3]), .Z(\w1[0][3] ) );
  XOR U45 ( .A(state[38]), .B(g_input[38]), .Z(\w1[0][38] ) );
  XOR U46 ( .A(state[37]), .B(g_input[37]), .Z(\w1[0][37] ) );
  XOR U47 ( .A(state[35]), .B(g_input[35]), .Z(\w1[0][35] ) );
  XOR U48 ( .A(state[30]), .B(g_input[30]), .Z(\w1[0][30] ) );
  XOR U49 ( .A(state[29]), .B(g_input[29]), .Z(\w1[0][29] ) );
  XOR U50 ( .A(state[27]), .B(g_input[27]), .Z(\w1[0][27] ) );
  XOR U51 ( .A(state[22]), .B(g_input[22]), .Z(\w1[0][22] ) );
  XOR U52 ( .A(state[21]), .B(g_input[21]), .Z(\w1[0][21] ) );
  XOR U53 ( .A(state[19]), .B(g_input[19]), .Z(\w1[0][19] ) );
  XOR U54 ( .A(state[14]), .B(g_input[14]), .Z(\w1[0][14] ) );
  XOR U55 ( .A(state[13]), .B(g_input[13]), .Z(\w1[0][13] ) );
  XOR U56 ( .A(state[126]), .B(g_input[126]), .Z(\w1[0][126] ) );
  XOR U57 ( .A(state[125]), .B(g_input[125]), .Z(\w1[0][125] ) );
  XOR U58 ( .A(state[123]), .B(g_input[123]), .Z(\w1[0][123] ) );
  XOR U59 ( .A(state[11]), .B(g_input[11]), .Z(\w1[0][11] ) );
  XOR U60 ( .A(state[118]), .B(g_input[118]), .Z(\w1[0][118] ) );
  XOR U61 ( .A(state[117]), .B(g_input[117]), .Z(\w1[0][117] ) );
  XOR U62 ( .A(state[115]), .B(g_input[115]), .Z(\w1[0][115] ) );
  XOR U63 ( .A(state[110]), .B(g_input[110]), .Z(\w1[0][110] ) );
  XOR U64 ( .A(state[109]), .B(g_input[109]), .Z(\w1[0][109] ) );
  XOR U65 ( .A(state[107]), .B(g_input[107]), .Z(\w1[0][107] ) );
  XOR U66 ( .A(state[102]), .B(g_input[102]), .Z(\w1[0][102] ) );
  XOR U67 ( .A(state[101]), .B(g_input[101]), .Z(\w1[0][101] ) );
  XNOR U68 ( .A(g_input[9]), .B(\SUBBYTES[0].a/n1690 ), .Z(o[9]) );
  XNOR U69 ( .A(g_input[99]), .B(\SUBBYTES[0].a/n1620 ), .Z(o[99]) );
  XNOR U70 ( .A(g_input[98]), .B(\SUBBYTES[0].a/n1619 ), .Z(o[98]) );
  XNOR U71 ( .A(g_input[97]), .B(\SUBBYTES[0].a/n1618 ), .Z(o[97]) );
  XNOR U72 ( .A(g_input[96]), .B(\SUBBYTES[0].a/n1617 ), .Z(o[96]) );
  XNOR U73 ( .A(g_input[95]), .B(\SUBBYTES[0].a/n1712 ), .Z(o[95]) );
  XNOR U74 ( .A(g_input[94]), .B(\SUBBYTES[0].a/n1711 ), .Z(o[94]) );
  XNOR U75 ( .A(g_input[93]), .B(\SUBBYTES[0].a/n1710 ), .Z(o[93]) );
  XNOR U76 ( .A(g_input[92]), .B(\SUBBYTES[0].a/n1709 ), .Z(o[92]) );
  XNOR U77 ( .A(g_input[91]), .B(\SUBBYTES[0].a/n1708 ), .Z(o[91]) );
  XNOR U78 ( .A(g_input[90]), .B(\SUBBYTES[0].a/n1707 ), .Z(o[90]) );
  XNOR U79 ( .A(g_input[8]), .B(\SUBBYTES[0].a/n1689 ), .Z(o[8]) );
  XNOR U80 ( .A(g_input[89]), .B(\SUBBYTES[0].a/n1706 ), .Z(o[89]) );
  XNOR U81 ( .A(g_input[88]), .B(\SUBBYTES[0].a/n1705 ), .Z(o[88]) );
  XNOR U82 ( .A(g_input[87]), .B(\SUBBYTES[0].a/n1672 ), .Z(o[87]) );
  XNOR U83 ( .A(g_input[86]), .B(\SUBBYTES[0].a/n1671 ), .Z(o[86]) );
  XNOR U84 ( .A(g_input[85]), .B(\SUBBYTES[0].a/n1670 ), .Z(o[85]) );
  XNOR U85 ( .A(g_input[84]), .B(\SUBBYTES[0].a/n1669 ), .Z(o[84]) );
  XNOR U86 ( .A(g_input[83]), .B(\SUBBYTES[0].a/n1668 ), .Z(o[83]) );
  XNOR U87 ( .A(g_input[82]), .B(\SUBBYTES[0].a/n1667 ), .Z(o[82]) );
  XNOR U88 ( .A(g_input[81]), .B(\SUBBYTES[0].a/n1666 ), .Z(o[81]) );
  XNOR U89 ( .A(g_input[80]), .B(\SUBBYTES[0].a/n1665 ), .Z(o[80]) );
  XNOR U90 ( .A(g_input[7]), .B(\SUBBYTES[0].a/n1656 ), .Z(o[7]) );
  XNOR U91 ( .A(g_input[79]), .B(\SUBBYTES[0].a/n1632 ), .Z(o[79]) );
  XNOR U92 ( .A(g_input[78]), .B(\SUBBYTES[0].a/n1631 ), .Z(o[78]) );
  XNOR U93 ( .A(g_input[77]), .B(\SUBBYTES[0].a/n1630 ), .Z(o[77]) );
  XNOR U94 ( .A(g_input[76]), .B(\SUBBYTES[0].a/n1629 ), .Z(o[76]) );
  XNOR U95 ( .A(g_input[75]), .B(\SUBBYTES[0].a/n1628 ), .Z(o[75]) );
  XNOR U96 ( .A(g_input[74]), .B(\SUBBYTES[0].a/n1627 ), .Z(o[74]) );
  XNOR U97 ( .A(g_input[73]), .B(\SUBBYTES[0].a/n1626 ), .Z(o[73]) );
  XNOR U98 ( .A(g_input[72]), .B(\SUBBYTES[0].a/n1625 ), .Z(o[72]) );
  XNOR U99 ( .A(g_input[71]), .B(\SUBBYTES[0].a/n1720 ), .Z(o[71]) );
  XNOR U100 ( .A(g_input[70]), .B(\SUBBYTES[0].a/n1719 ), .Z(o[70]) );
  XNOR U101 ( .A(g_input[6]), .B(\SUBBYTES[0].a/n1655 ), .Z(o[6]) );
  XNOR U102 ( .A(g_input[69]), .B(\SUBBYTES[0].a/n1718 ), .Z(o[69]) );
  XNOR U103 ( .A(g_input[68]), .B(\SUBBYTES[0].a/n1717 ), .Z(o[68]) );
  XNOR U104 ( .A(g_input[67]), .B(\SUBBYTES[0].a/n1716 ), .Z(o[67]) );
  XNOR U105 ( .A(g_input[66]), .B(\SUBBYTES[0].a/n1715 ), .Z(o[66]) );
  XNOR U106 ( .A(g_input[65]), .B(\SUBBYTES[0].a/n1714 ), .Z(o[65]) );
  XNOR U107 ( .A(g_input[64]), .B(\SUBBYTES[0].a/n1713 ), .Z(o[64]) );
  XNOR U108 ( .A(g_input[63]), .B(\SUBBYTES[0].a/n1680 ), .Z(o[63]) );
  XNOR U109 ( .A(g_input[62]), .B(\SUBBYTES[0].a/n1679 ), .Z(o[62]) );
  XNOR U110 ( .A(g_input[61]), .B(\SUBBYTES[0].a/n1678 ), .Z(o[61]) );
  XNOR U111 ( .A(g_input[60]), .B(\SUBBYTES[0].a/n1677 ), .Z(o[60]) );
  XNOR U112 ( .A(g_input[5]), .B(\SUBBYTES[0].a/n1654 ), .Z(o[5]) );
  XNOR U113 ( .A(g_input[59]), .B(\SUBBYTES[0].a/n1676 ), .Z(o[59]) );
  XNOR U114 ( .A(g_input[58]), .B(\SUBBYTES[0].a/n1675 ), .Z(o[58]) );
  XNOR U115 ( .A(g_input[57]), .B(\SUBBYTES[0].a/n1674 ), .Z(o[57]) );
  XNOR U116 ( .A(g_input[56]), .B(\SUBBYTES[0].a/n1673 ), .Z(o[56]) );
  XNOR U117 ( .A(g_input[55]), .B(\SUBBYTES[0].a/n1640 ), .Z(o[55]) );
  XNOR U118 ( .A(g_input[54]), .B(\SUBBYTES[0].a/n1639 ), .Z(o[54]) );
  XNOR U119 ( .A(g_input[53]), .B(\SUBBYTES[0].a/n1638 ), .Z(o[53]) );
  XNOR U120 ( .A(g_input[52]), .B(\SUBBYTES[0].a/n1637 ), .Z(o[52]) );
  XNOR U121 ( .A(g_input[51]), .B(\SUBBYTES[0].a/n1636 ), .Z(o[51]) );
  XNOR U122 ( .A(g_input[50]), .B(\SUBBYTES[0].a/n1635 ), .Z(o[50]) );
  XNOR U123 ( .A(g_input[4]), .B(\SUBBYTES[0].a/n1653 ), .Z(o[4]) );
  XNOR U124 ( .A(g_input[49]), .B(\SUBBYTES[0].a/n1634 ), .Z(o[49]) );
  XNOR U125 ( .A(g_input[48]), .B(\SUBBYTES[0].a/n1633 ), .Z(o[48]) );
  XNOR U126 ( .A(g_input[47]), .B(\SUBBYTES[0].a/n1728 ), .Z(o[47]) );
  XNOR U127 ( .A(g_input[46]), .B(\SUBBYTES[0].a/n1727 ), .Z(o[46]) );
  XNOR U128 ( .A(g_input[45]), .B(\SUBBYTES[0].a/n1726 ), .Z(o[45]) );
  XNOR U129 ( .A(g_input[44]), .B(\SUBBYTES[0].a/n1725 ), .Z(o[44]) );
  XNOR U130 ( .A(g_input[43]), .B(\SUBBYTES[0].a/n1724 ), .Z(o[43]) );
  XNOR U131 ( .A(g_input[42]), .B(\SUBBYTES[0].a/n1723 ), .Z(o[42]) );
  XNOR U132 ( .A(g_input[41]), .B(\SUBBYTES[0].a/n1722 ), .Z(o[41]) );
  XNOR U133 ( .A(g_input[40]), .B(\SUBBYTES[0].a/n1721 ), .Z(o[40]) );
  XNOR U134 ( .A(g_input[3]), .B(\SUBBYTES[0].a/n1652 ), .Z(o[3]) );
  XNOR U135 ( .A(g_input[39]), .B(\SUBBYTES[0].a/n1688 ), .Z(o[39]) );
  XNOR U136 ( .A(g_input[38]), .B(\SUBBYTES[0].a/n1687 ), .Z(o[38]) );
  XNOR U137 ( .A(g_input[37]), .B(\SUBBYTES[0].a/n1686 ), .Z(o[37]) );
  XNOR U138 ( .A(g_input[36]), .B(\SUBBYTES[0].a/n1685 ), .Z(o[36]) );
  XNOR U139 ( .A(g_input[35]), .B(\SUBBYTES[0].a/n1684 ), .Z(o[35]) );
  XNOR U140 ( .A(g_input[34]), .B(\SUBBYTES[0].a/n1683 ), .Z(o[34]) );
  XNOR U141 ( .A(g_input[33]), .B(\SUBBYTES[0].a/n1682 ), .Z(o[33]) );
  XNOR U142 ( .A(g_input[32]), .B(\SUBBYTES[0].a/n1681 ), .Z(o[32]) );
  XNOR U143 ( .A(g_input[31]), .B(\SUBBYTES[0].a/n1648 ), .Z(o[31]) );
  XNOR U144 ( .A(g_input[30]), .B(\SUBBYTES[0].a/n1647 ), .Z(o[30]) );
  XNOR U145 ( .A(g_input[2]), .B(\SUBBYTES[0].a/n1651 ), .Z(o[2]) );
  XNOR U146 ( .A(g_input[29]), .B(\SUBBYTES[0].a/n1646 ), .Z(o[29]) );
  XNOR U147 ( .A(g_input[28]), .B(\SUBBYTES[0].a/n1645 ), .Z(o[28]) );
  XNOR U148 ( .A(g_input[27]), .B(\SUBBYTES[0].a/n1644 ), .Z(o[27]) );
  XNOR U149 ( .A(g_input[26]), .B(\SUBBYTES[0].a/n1643 ), .Z(o[26]) );
  XNOR U150 ( .A(g_input[25]), .B(\SUBBYTES[0].a/n1642 ), .Z(o[25]) );
  XNOR U151 ( .A(g_input[24]), .B(\SUBBYTES[0].a/n1641 ), .Z(o[24]) );
  XNOR U152 ( .A(g_input[23]), .B(\SUBBYTES[0].a/n1736 ), .Z(o[23]) );
  XNOR U153 ( .A(g_input[22]), .B(\SUBBYTES[0].a/n1735 ), .Z(o[22]) );
  XNOR U154 ( .A(g_input[21]), .B(\SUBBYTES[0].a/n1734 ), .Z(o[21]) );
  XNOR U155 ( .A(g_input[20]), .B(\SUBBYTES[0].a/n1733 ), .Z(o[20]) );
  XNOR U156 ( .A(g_input[1]), .B(\SUBBYTES[0].a/n1650 ), .Z(o[1]) );
  XNOR U157 ( .A(g_input[19]), .B(\SUBBYTES[0].a/n1732 ), .Z(o[19]) );
  XNOR U158 ( .A(g_input[18]), .B(\SUBBYTES[0].a/n1731 ), .Z(o[18]) );
  XNOR U159 ( .A(g_input[17]), .B(\SUBBYTES[0].a/n1730 ), .Z(o[17]) );
  XNOR U160 ( .A(g_input[16]), .B(\SUBBYTES[0].a/n1729 ), .Z(o[16]) );
  XNOR U161 ( .A(g_input[15]), .B(\SUBBYTES[0].a/n1696 ), .Z(o[15]) );
  XNOR U162 ( .A(g_input[14]), .B(\SUBBYTES[0].a/n1695 ), .Z(o[14]) );
  XNOR U163 ( .A(g_input[13]), .B(\SUBBYTES[0].a/n1694 ), .Z(o[13]) );
  XNOR U164 ( .A(g_input[12]), .B(\SUBBYTES[0].a/n1693 ), .Z(o[12]) );
  XNOR U165 ( .A(g_input[127]), .B(\SUBBYTES[0].a/n1744 ), .Z(o[127]) );
  XNOR U166 ( .A(g_input[126]), .B(\SUBBYTES[0].a/n1743 ), .Z(o[126]) );
  XNOR U167 ( .A(g_input[125]), .B(\SUBBYTES[0].a/n1742 ), .Z(o[125]) );
  XNOR U168 ( .A(g_input[124]), .B(\SUBBYTES[0].a/n1741 ), .Z(o[124]) );
  XNOR U169 ( .A(g_input[123]), .B(\SUBBYTES[0].a/n1740 ), .Z(o[123]) );
  XNOR U170 ( .A(g_input[122]), .B(\SUBBYTES[0].a/n1739 ), .Z(o[122]) );
  XNOR U171 ( .A(g_input[121]), .B(\SUBBYTES[0].a/n1738 ), .Z(o[121]) );
  XNOR U172 ( .A(g_input[120]), .B(\SUBBYTES[0].a/n1737 ), .Z(o[120]) );
  XNOR U173 ( .A(g_input[11]), .B(\SUBBYTES[0].a/n1692 ), .Z(o[11]) );
  XNOR U174 ( .A(g_input[119]), .B(\SUBBYTES[0].a/n1704 ), .Z(o[119]) );
  XNOR U175 ( .A(g_input[118]), .B(\SUBBYTES[0].a/n1703 ), .Z(o[118]) );
  XNOR U176 ( .A(g_input[117]), .B(\SUBBYTES[0].a/n1702 ), .Z(o[117]) );
  XNOR U177 ( .A(g_input[116]), .B(\SUBBYTES[0].a/n1701 ), .Z(o[116]) );
  XNOR U178 ( .A(g_input[115]), .B(\SUBBYTES[0].a/n1700 ), .Z(o[115]) );
  XNOR U179 ( .A(g_input[114]), .B(\SUBBYTES[0].a/n1699 ), .Z(o[114]) );
  XNOR U180 ( .A(g_input[113]), .B(\SUBBYTES[0].a/n1698 ), .Z(o[113]) );
  XNOR U181 ( .A(g_input[112]), .B(\SUBBYTES[0].a/n1697 ), .Z(o[112]) );
  XNOR U182 ( .A(g_input[111]), .B(\SUBBYTES[0].a/n1664 ), .Z(o[111]) );
  XNOR U183 ( .A(g_input[110]), .B(\SUBBYTES[0].a/n1663 ), .Z(o[110]) );
  XNOR U184 ( .A(g_input[10]), .B(\SUBBYTES[0].a/n1691 ), .Z(o[10]) );
  XNOR U185 ( .A(g_input[109]), .B(\SUBBYTES[0].a/n1662 ), .Z(o[109]) );
  XNOR U186 ( .A(g_input[108]), .B(\SUBBYTES[0].a/n1661 ), .Z(o[108]) );
  XNOR U187 ( .A(g_input[107]), .B(\SUBBYTES[0].a/n1660 ), .Z(o[107]) );
  XNOR U188 ( .A(g_input[106]), .B(\SUBBYTES[0].a/n1659 ), .Z(o[106]) );
  XNOR U189 ( .A(g_input[105]), .B(\SUBBYTES[0].a/n1658 ), .Z(o[105]) );
  XNOR U190 ( .A(g_input[104]), .B(\SUBBYTES[0].a/n1657 ), .Z(o[104]) );
  XNOR U191 ( .A(g_input[103]), .B(\SUBBYTES[0].a/n1624 ), .Z(o[103]) );
  XNOR U192 ( .A(g_input[102]), .B(\SUBBYTES[0].a/n1623 ), .Z(o[102]) );
  XNOR U193 ( .A(g_input[101]), .B(\SUBBYTES[0].a/n1622 ), .Z(o[101]) );
  XNOR U194 ( .A(g_input[100]), .B(\SUBBYTES[0].a/n1621 ), .Z(o[100]) );
  XNOR U195 ( .A(g_input[0]), .B(\SUBBYTES[0].a/n1649 ), .Z(o[0]) );
  AND U196 ( .A(n17), .B(\SUBBYTES[0].a/w781 ), .Z(\SUBBYTES[0].a/w916 ) );
  AND U197 ( .A(n18), .B(\SUBBYTES[0].a/w782 ), .Z(\SUBBYTES[0].a/w914 ) );
  AND U198 ( .A(\SUBBYTES[0].a/w912 ), .B(n19), .Z(\SUBBYTES[0].a/w913 ) );
  ANDN U199 ( .A(\w1[0][96] ), .B(n20), .Z(\SUBBYTES[0].a/w909 ) );
  AND U200 ( .A(n21), .B(\SUBBYTES[0].a/w784 ), .Z(\SUBBYTES[0].a/w907 ) );
  AND U201 ( .A(\SUBBYTES[0].a/w905 ), .B(n22), .Z(\SUBBYTES[0].a/w906 ) );
  XOR U202 ( .A(\SUBBYTES[0].a/w849 ), .B(\SUBBYTES[0].a/n39 ), .Z(n22) );
  AND U203 ( .A(\SUBBYTES[0].a/w892 ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/w901 ) );
  AND U204 ( .A(\SUBBYTES[0].a/w893 ), .B(\SUBBYTES[0].a/w895 ), .Z(
        \SUBBYTES[0].a/w899 ) );
  AND U205 ( .A(\SUBBYTES[0].a/w896 ), .B(\SUBBYTES[0].a/w897 ), .Z(
        \SUBBYTES[0].a/w898 ) );
  AND U206 ( .A(\SUBBYTES[0].a/w785 ), .B(n17), .Z(\SUBBYTES[0].a/w884 ) );
  XOR U207 ( .A(\SUBBYTES[0].a/w853 ), .B(n4), .Z(n17) );
  AND U208 ( .A(\SUBBYTES[0].a/w786 ), .B(n18), .Z(\SUBBYTES[0].a/w882 ) );
  XOR U209 ( .A(\SUBBYTES[0].a/n40 ), .B(\SUBBYTES[0].a/w853 ), .Z(n18) );
  ANDN U210 ( .A(n19), .B(n23), .Z(\SUBBYTES[0].a/w881 ) );
  XOR U211 ( .A(n4), .B(\SUBBYTES[0].a/n40 ), .Z(n19) );
  ANDN U212 ( .A(\SUBBYTES[0].a/w787 ), .B(n20), .Z(\SUBBYTES[0].a/w877 ) );
  XNOR U213 ( .A(\SUBBYTES[0].a/w846 ), .B(\SUBBYTES[0].a/w849 ), .Z(n20) );
  AND U214 ( .A(\SUBBYTES[0].a/w788 ), .B(n21), .Z(\SUBBYTES[0].a/w875 ) );
  XNOR U215 ( .A(n24), .B(\SUBBYTES[0].a/w846 ), .Z(n21) );
  AND U216 ( .A(\SUBBYTES[0].a/w873 ), .B(n25), .Z(\SUBBYTES[0].a/w874 ) );
  XOR U217 ( .A(n26), .B(n24), .Z(n25) );
  IV U218 ( .A(\SUBBYTES[0].a/n39 ), .Z(n24) );
  ANDN U219 ( .A(\SUBBYTES[0].a/w892 ), .B(n27), .Z(\SUBBYTES[0].a/w869 ) );
  ANDN U220 ( .A(\SUBBYTES[0].a/w893 ), .B(n28), .Z(\SUBBYTES[0].a/w867 ) );
  AND U221 ( .A(n29), .B(\SUBBYTES[0].a/w896 ), .Z(\SUBBYTES[0].a/w866 ) );
  AND U222 ( .A(\SUBBYTES[0].a/w852 ), .B(\SUBBYTES[0].a/w851 ), .Z(
        \SUBBYTES[0].a/w853 ) );
  IV U223 ( .A(n26), .Z(\SUBBYTES[0].a/w849 ) );
  NAND U224 ( .A(\SUBBYTES[0].a/w828 ), .B(\SUBBYTES[0].a/w843 ), .Z(n26) );
  AND U225 ( .A(\SUBBYTES[0].a/w845 ), .B(\SUBBYTES[0].a/w851 ), .Z(
        \SUBBYTES[0].a/w846 ) );
  AND U226 ( .A(\SUBBYTES[0].a/w830 ), .B(\SUBBYTES[0].a/w828 ), .Z(
        \SUBBYTES[0].a/w840 ) );
  AND U227 ( .A(\SUBBYTES[0].a/w831 ), .B(\SUBBYTES[0].a/w829 ), .Z(
        \SUBBYTES[0].a/w838 ) );
  AND U228 ( .A(\SUBBYTES[0].a/w845 ), .B(\SUBBYTES[0].a/w852 ), .Z(
        \SUBBYTES[0].a/w837 ) );
  AND U229 ( .A(\SUBBYTES[0].a/w785 ), .B(\SUBBYTES[0].a/w781 ), .Z(
        \SUBBYTES[0].a/w822 ) );
  AND U230 ( .A(\SUBBYTES[0].a/w786 ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w820 ) );
  ANDN U231 ( .A(\SUBBYTES[0].a/w912 ), .B(n23), .Z(\SUBBYTES[0].a/w819 ) );
  XNOR U232 ( .A(\w1[0][103] ), .B(\w1[0][97] ), .Z(n23) );
  XOR U233 ( .A(g_input[97]), .B(state[97]), .Z(\w1[0][97] ) );
  IV U234 ( .A(n30), .Z(\w1[0][103] ) );
  AND U235 ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w787 ), .Z(
        \SUBBYTES[0].a/w815 ) );
  XOR U236 ( .A(g_input[96]), .B(state[96]), .Z(\w1[0][96] ) );
  AND U237 ( .A(\SUBBYTES[0].a/w788 ), .B(\SUBBYTES[0].a/w784 ), .Z(
        \SUBBYTES[0].a/w813 ) );
  AND U238 ( .A(\SUBBYTES[0].a/w873 ), .B(\SUBBYTES[0].a/w905 ), .Z(
        \SUBBYTES[0].a/w812 ) );
  ANDN U239 ( .A(\SUBBYTES[0].a/w894 ), .B(n27), .Z(\SUBBYTES[0].a/w807 ) );
  XOR U240 ( .A(\w1[0][100] ), .B(n30), .Z(n27) );
  ANDN U241 ( .A(\SUBBYTES[0].a/w895 ), .B(n28), .Z(\SUBBYTES[0].a/w805 ) );
  XOR U242 ( .A(n30), .B(\w1[0][98] ), .Z(n28) );
  XNOR U243 ( .A(g_input[103]), .B(state[103]), .Z(n30) );
  AND U244 ( .A(\SUBBYTES[0].a/w897 ), .B(n29), .Z(\SUBBYTES[0].a/w804 ) );
  XOR U245 ( .A(\w1[0][100] ), .B(\w1[0][98] ), .Z(n29) );
  XOR U246 ( .A(g_input[98]), .B(state[98]), .Z(\w1[0][98] ) );
  XOR U247 ( .A(g_input[100]), .B(state[100]), .Z(\w1[0][100] ) );
  AND U248 ( .A(n31), .B(\SUBBYTES[0].a/w574 ), .Z(\SUBBYTES[0].a/w709 ) );
  AND U249 ( .A(n32), .B(\SUBBYTES[0].a/w575 ), .Z(\SUBBYTES[0].a/w707 ) );
  AND U250 ( .A(\SUBBYTES[0].a/w705 ), .B(n33), .Z(\SUBBYTES[0].a/w706 ) );
  ANDN U251 ( .A(\w1[0][104] ), .B(n34), .Z(\SUBBYTES[0].a/w702 ) );
  AND U252 ( .A(n35), .B(\SUBBYTES[0].a/w577 ), .Z(\SUBBYTES[0].a/w700 ) );
  AND U253 ( .A(\SUBBYTES[0].a/w698 ), .B(n36), .Z(\SUBBYTES[0].a/w699 ) );
  XOR U254 ( .A(\SUBBYTES[0].a/w642 ), .B(\SUBBYTES[0].a/n29 ), .Z(n36) );
  AND U255 ( .A(\SUBBYTES[0].a/w685 ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/w694 ) );
  AND U256 ( .A(\SUBBYTES[0].a/w686 ), .B(\SUBBYTES[0].a/w688 ), .Z(
        \SUBBYTES[0].a/w692 ) );
  AND U257 ( .A(\SUBBYTES[0].a/w689 ), .B(\SUBBYTES[0].a/w690 ), .Z(
        \SUBBYTES[0].a/w691 ) );
  AND U258 ( .A(\SUBBYTES[0].a/w578 ), .B(n31), .Z(\SUBBYTES[0].a/w677 ) );
  XOR U259 ( .A(\SUBBYTES[0].a/w646 ), .B(n3), .Z(n31) );
  AND U260 ( .A(\SUBBYTES[0].a/w579 ), .B(n32), .Z(\SUBBYTES[0].a/w675 ) );
  XOR U261 ( .A(\SUBBYTES[0].a/n30 ), .B(\SUBBYTES[0].a/w646 ), .Z(n32) );
  AND U262 ( .A(n37), .B(n33), .Z(\SUBBYTES[0].a/w674 ) );
  XOR U263 ( .A(n3), .B(\SUBBYTES[0].a/n30 ), .Z(n33) );
  ANDN U264 ( .A(\SUBBYTES[0].a/w580 ), .B(n34), .Z(\SUBBYTES[0].a/w670 ) );
  XNOR U265 ( .A(\SUBBYTES[0].a/w639 ), .B(\SUBBYTES[0].a/w642 ), .Z(n34) );
  AND U266 ( .A(\SUBBYTES[0].a/w581 ), .B(n35), .Z(\SUBBYTES[0].a/w668 ) );
  XNOR U267 ( .A(n38), .B(\SUBBYTES[0].a/w639 ), .Z(n35) );
  AND U268 ( .A(\SUBBYTES[0].a/w666 ), .B(n39), .Z(\SUBBYTES[0].a/w667 ) );
  XOR U269 ( .A(n40), .B(n38), .Z(n39) );
  IV U270 ( .A(\SUBBYTES[0].a/n29 ), .Z(n38) );
  AND U271 ( .A(n41), .B(\SUBBYTES[0].a/w685 ), .Z(\SUBBYTES[0].a/w662 ) );
  ANDN U272 ( .A(\SUBBYTES[0].a/w686 ), .B(n42), .Z(\SUBBYTES[0].a/w660 ) );
  AND U273 ( .A(n43), .B(\SUBBYTES[0].a/w689 ), .Z(\SUBBYTES[0].a/w659 ) );
  AND U274 ( .A(\SUBBYTES[0].a/w645 ), .B(\SUBBYTES[0].a/w644 ), .Z(
        \SUBBYTES[0].a/w646 ) );
  IV U275 ( .A(n40), .Z(\SUBBYTES[0].a/w642 ) );
  NAND U276 ( .A(\SUBBYTES[0].a/w621 ), .B(\SUBBYTES[0].a/w636 ), .Z(n40) );
  AND U277 ( .A(\SUBBYTES[0].a/w638 ), .B(\SUBBYTES[0].a/w644 ), .Z(
        \SUBBYTES[0].a/w639 ) );
  AND U278 ( .A(\SUBBYTES[0].a/w623 ), .B(\SUBBYTES[0].a/w621 ), .Z(
        \SUBBYTES[0].a/w633 ) );
  AND U279 ( .A(\SUBBYTES[0].a/w624 ), .B(\SUBBYTES[0].a/w622 ), .Z(
        \SUBBYTES[0].a/w631 ) );
  AND U280 ( .A(\SUBBYTES[0].a/w638 ), .B(\SUBBYTES[0].a/w645 ), .Z(
        \SUBBYTES[0].a/w630 ) );
  AND U281 ( .A(\SUBBYTES[0].a/w578 ), .B(\SUBBYTES[0].a/w574 ), .Z(
        \SUBBYTES[0].a/w615 ) );
  AND U282 ( .A(\SUBBYTES[0].a/w579 ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w613 ) );
  AND U283 ( .A(\SUBBYTES[0].a/w705 ), .B(n37), .Z(\SUBBYTES[0].a/w612 ) );
  XNOR U284 ( .A(\w1[0][105] ), .B(n44), .Z(n37) );
  XOR U285 ( .A(g_input[105]), .B(state[105]), .Z(\w1[0][105] ) );
  AND U286 ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w580 ), .Z(
        \SUBBYTES[0].a/w608 ) );
  XOR U287 ( .A(g_input[104]), .B(state[104]), .Z(\w1[0][104] ) );
  AND U288 ( .A(\SUBBYTES[0].a/w581 ), .B(\SUBBYTES[0].a/w577 ), .Z(
        \SUBBYTES[0].a/w606 ) );
  AND U289 ( .A(\SUBBYTES[0].a/w666 ), .B(\SUBBYTES[0].a/w698 ), .Z(
        \SUBBYTES[0].a/w605 ) );
  AND U290 ( .A(\SUBBYTES[0].a/w687 ), .B(n41), .Z(\SUBBYTES[0].a/w600 ) );
  XOR U291 ( .A(\w1[0][108] ), .B(\w1[0][111] ), .Z(n41) );
  ANDN U292 ( .A(\SUBBYTES[0].a/w688 ), .B(n42), .Z(\SUBBYTES[0].a/w598 ) );
  XNOR U293 ( .A(\w1[0][106] ), .B(\w1[0][111] ), .Z(n42) );
  IV U294 ( .A(n44), .Z(\w1[0][111] ) );
  XNOR U295 ( .A(g_input[111]), .B(state[111]), .Z(n44) );
  AND U296 ( .A(\SUBBYTES[0].a/w690 ), .B(n43), .Z(\SUBBYTES[0].a/w597 ) );
  XOR U297 ( .A(\w1[0][106] ), .B(\w1[0][108] ), .Z(n43) );
  XOR U298 ( .A(g_input[108]), .B(state[108]), .Z(\w1[0][108] ) );
  XOR U299 ( .A(g_input[106]), .B(state[106]), .Z(\w1[0][106] ) );
  AND U300 ( .A(n45), .B(\SUBBYTES[0].a/w367 ), .Z(\SUBBYTES[0].a/w502 ) );
  AND U301 ( .A(n46), .B(\SUBBYTES[0].a/w368 ), .Z(\SUBBYTES[0].a/w500 ) );
  AND U302 ( .A(\SUBBYTES[0].a/w498 ), .B(n47), .Z(\SUBBYTES[0].a/w499 ) );
  ANDN U303 ( .A(\w1[0][112] ), .B(n48), .Z(\SUBBYTES[0].a/w495 ) );
  AND U304 ( .A(n49), .B(\SUBBYTES[0].a/w370 ), .Z(\SUBBYTES[0].a/w493 ) );
  AND U305 ( .A(\SUBBYTES[0].a/w491 ), .B(n50), .Z(\SUBBYTES[0].a/w492 ) );
  XOR U306 ( .A(\SUBBYTES[0].a/w435 ), .B(\SUBBYTES[0].a/n19 ), .Z(n50) );
  AND U307 ( .A(\SUBBYTES[0].a/w478 ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/w487 ) );
  AND U308 ( .A(\SUBBYTES[0].a/w479 ), .B(\SUBBYTES[0].a/w481 ), .Z(
        \SUBBYTES[0].a/w485 ) );
  AND U309 ( .A(\SUBBYTES[0].a/w482 ), .B(\SUBBYTES[0].a/w483 ), .Z(
        \SUBBYTES[0].a/w484 ) );
  AND U310 ( .A(\SUBBYTES[0].a/w371 ), .B(n45), .Z(\SUBBYTES[0].a/w470 ) );
  XOR U311 ( .A(\SUBBYTES[0].a/w439 ), .B(n2), .Z(n45) );
  AND U312 ( .A(\SUBBYTES[0].a/w372 ), .B(n46), .Z(\SUBBYTES[0].a/w468 ) );
  XOR U313 ( .A(\SUBBYTES[0].a/n20 ), .B(\SUBBYTES[0].a/w439 ), .Z(n46) );
  AND U314 ( .A(n51), .B(n47), .Z(\SUBBYTES[0].a/w467 ) );
  XOR U315 ( .A(n2), .B(\SUBBYTES[0].a/n20 ), .Z(n47) );
  ANDN U316 ( .A(\SUBBYTES[0].a/w373 ), .B(n48), .Z(\SUBBYTES[0].a/w463 ) );
  XNOR U317 ( .A(\SUBBYTES[0].a/w432 ), .B(\SUBBYTES[0].a/w435 ), .Z(n48) );
  AND U318 ( .A(\SUBBYTES[0].a/w374 ), .B(n49), .Z(\SUBBYTES[0].a/w461 ) );
  XNOR U319 ( .A(n52), .B(\SUBBYTES[0].a/w432 ), .Z(n49) );
  AND U320 ( .A(\SUBBYTES[0].a/w459 ), .B(n53), .Z(\SUBBYTES[0].a/w460 ) );
  XOR U321 ( .A(n54), .B(n52), .Z(n53) );
  IV U322 ( .A(\SUBBYTES[0].a/n19 ), .Z(n52) );
  AND U323 ( .A(n55), .B(\SUBBYTES[0].a/w478 ), .Z(\SUBBYTES[0].a/w455 ) );
  ANDN U324 ( .A(\SUBBYTES[0].a/w479 ), .B(n56), .Z(\SUBBYTES[0].a/w453 ) );
  AND U325 ( .A(n57), .B(\SUBBYTES[0].a/w482 ), .Z(\SUBBYTES[0].a/w452 ) );
  AND U326 ( .A(\SUBBYTES[0].a/w438 ), .B(\SUBBYTES[0].a/w437 ), .Z(
        \SUBBYTES[0].a/w439 ) );
  IV U327 ( .A(n54), .Z(\SUBBYTES[0].a/w435 ) );
  NAND U328 ( .A(\SUBBYTES[0].a/w414 ), .B(\SUBBYTES[0].a/w429 ), .Z(n54) );
  AND U329 ( .A(\SUBBYTES[0].a/w431 ), .B(\SUBBYTES[0].a/w437 ), .Z(
        \SUBBYTES[0].a/w432 ) );
  AND U330 ( .A(\SUBBYTES[0].a/w416 ), .B(\SUBBYTES[0].a/w414 ), .Z(
        \SUBBYTES[0].a/w426 ) );
  AND U331 ( .A(\SUBBYTES[0].a/w417 ), .B(\SUBBYTES[0].a/w415 ), .Z(
        \SUBBYTES[0].a/w424 ) );
  AND U332 ( .A(\SUBBYTES[0].a/w431 ), .B(\SUBBYTES[0].a/w438 ), .Z(
        \SUBBYTES[0].a/w423 ) );
  AND U333 ( .A(\SUBBYTES[0].a/w371 ), .B(\SUBBYTES[0].a/w367 ), .Z(
        \SUBBYTES[0].a/w408 ) );
  AND U334 ( .A(\SUBBYTES[0].a/w372 ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w406 ) );
  AND U335 ( .A(\SUBBYTES[0].a/w498 ), .B(n51), .Z(\SUBBYTES[0].a/w405 ) );
  XNOR U336 ( .A(\w1[0][113] ), .B(n58), .Z(n51) );
  XOR U337 ( .A(g_input[113]), .B(state[113]), .Z(\w1[0][113] ) );
  AND U338 ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w373 ), .Z(
        \SUBBYTES[0].a/w401 ) );
  XOR U339 ( .A(g_input[112]), .B(state[112]), .Z(\w1[0][112] ) );
  AND U340 ( .A(\SUBBYTES[0].a/w374 ), .B(\SUBBYTES[0].a/w370 ), .Z(
        \SUBBYTES[0].a/w399 ) );
  AND U341 ( .A(\SUBBYTES[0].a/w459 ), .B(\SUBBYTES[0].a/w491 ), .Z(
        \SUBBYTES[0].a/w398 ) );
  AND U342 ( .A(\SUBBYTES[0].a/w480 ), .B(n55), .Z(\SUBBYTES[0].a/w393 ) );
  XOR U343 ( .A(\w1[0][116] ), .B(\w1[0][119] ), .Z(n55) );
  ANDN U344 ( .A(\SUBBYTES[0].a/w481 ), .B(n56), .Z(\SUBBYTES[0].a/w391 ) );
  XNOR U345 ( .A(\w1[0][114] ), .B(\w1[0][119] ), .Z(n56) );
  IV U346 ( .A(n58), .Z(\w1[0][119] ) );
  XNOR U347 ( .A(g_input[119]), .B(state[119]), .Z(n58) );
  AND U348 ( .A(\SUBBYTES[0].a/w483 ), .B(n57), .Z(\SUBBYTES[0].a/w390 ) );
  XOR U349 ( .A(\w1[0][114] ), .B(\w1[0][116] ), .Z(n57) );
  XOR U350 ( .A(g_input[116]), .B(state[116]), .Z(\w1[0][116] ) );
  XOR U351 ( .A(g_input[114]), .B(state[114]), .Z(\w1[0][114] ) );
  AND U352 ( .A(n59), .B(\SUBBYTES[0].a/w3265 ), .Z(\SUBBYTES[0].a/w3400 ) );
  AND U353 ( .A(n60), .B(\SUBBYTES[0].a/w3266 ), .Z(\SUBBYTES[0].a/w3398 ) );
  AND U354 ( .A(\SUBBYTES[0].a/w3396 ), .B(n61), .Z(\SUBBYTES[0].a/w3397 ) );
  ANDN U355 ( .A(\w1[0][0] ), .B(n62), .Z(\SUBBYTES[0].a/w3393 ) );
  AND U356 ( .A(n63), .B(\SUBBYTES[0].a/w3268 ), .Z(\SUBBYTES[0].a/w3391 ) );
  AND U357 ( .A(\SUBBYTES[0].a/w3389 ), .B(n64), .Z(\SUBBYTES[0].a/w3390 ) );
  XOR U358 ( .A(\SUBBYTES[0].a/w3333 ), .B(\SUBBYTES[0].a/n159 ), .Z(n64) );
  AND U359 ( .A(\SUBBYTES[0].a/w3376 ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/w3385 ) );
  AND U360 ( .A(\SUBBYTES[0].a/w3377 ), .B(\SUBBYTES[0].a/w3379 ), .Z(
        \SUBBYTES[0].a/w3383 ) );
  AND U361 ( .A(\SUBBYTES[0].a/w3380 ), .B(\SUBBYTES[0].a/w3381 ), .Z(
        \SUBBYTES[0].a/w3382 ) );
  AND U362 ( .A(\SUBBYTES[0].a/w3269 ), .B(n59), .Z(\SUBBYTES[0].a/w3368 ) );
  XOR U363 ( .A(\SUBBYTES[0].a/w3337 ), .B(n16), .Z(n59) );
  AND U364 ( .A(\SUBBYTES[0].a/w3270 ), .B(n60), .Z(\SUBBYTES[0].a/w3366 ) );
  XOR U365 ( .A(\SUBBYTES[0].a/n160 ), .B(\SUBBYTES[0].a/w3337 ), .Z(n60) );
  AND U366 ( .A(n65), .B(n61), .Z(\SUBBYTES[0].a/w3365 ) );
  XOR U367 ( .A(n16), .B(\SUBBYTES[0].a/n160 ), .Z(n61) );
  ANDN U368 ( .A(\SUBBYTES[0].a/w3271 ), .B(n62), .Z(\SUBBYTES[0].a/w3361 ) );
  XNOR U369 ( .A(\SUBBYTES[0].a/w3330 ), .B(\SUBBYTES[0].a/w3333 ), .Z(n62) );
  AND U370 ( .A(\SUBBYTES[0].a/w3272 ), .B(n63), .Z(\SUBBYTES[0].a/w3359 ) );
  XNOR U371 ( .A(n66), .B(\SUBBYTES[0].a/w3330 ), .Z(n63) );
  AND U372 ( .A(\SUBBYTES[0].a/w3357 ), .B(n67), .Z(\SUBBYTES[0].a/w3358 ) );
  XOR U373 ( .A(n68), .B(n66), .Z(n67) );
  IV U374 ( .A(\SUBBYTES[0].a/n159 ), .Z(n66) );
  AND U375 ( .A(n69), .B(\SUBBYTES[0].a/w3376 ), .Z(\SUBBYTES[0].a/w3353 ) );
  ANDN U376 ( .A(\SUBBYTES[0].a/w3377 ), .B(n70), .Z(\SUBBYTES[0].a/w3351 ) );
  AND U377 ( .A(n71), .B(\SUBBYTES[0].a/w3380 ), .Z(\SUBBYTES[0].a/w3350 ) );
  AND U378 ( .A(\SUBBYTES[0].a/w3336 ), .B(\SUBBYTES[0].a/w3335 ), .Z(
        \SUBBYTES[0].a/w3337 ) );
  IV U379 ( .A(n68), .Z(\SUBBYTES[0].a/w3333 ) );
  NAND U380 ( .A(\SUBBYTES[0].a/w3312 ), .B(\SUBBYTES[0].a/w3327 ), .Z(n68) );
  AND U381 ( .A(\SUBBYTES[0].a/w3329 ), .B(\SUBBYTES[0].a/w3335 ), .Z(
        \SUBBYTES[0].a/w3330 ) );
  AND U382 ( .A(\SUBBYTES[0].a/w3314 ), .B(\SUBBYTES[0].a/w3312 ), .Z(
        \SUBBYTES[0].a/w3324 ) );
  AND U383 ( .A(\SUBBYTES[0].a/w3315 ), .B(\SUBBYTES[0].a/w3313 ), .Z(
        \SUBBYTES[0].a/w3322 ) );
  AND U384 ( .A(\SUBBYTES[0].a/w3329 ), .B(\SUBBYTES[0].a/w3336 ), .Z(
        \SUBBYTES[0].a/w3321 ) );
  AND U385 ( .A(\SUBBYTES[0].a/w3269 ), .B(\SUBBYTES[0].a/w3265 ), .Z(
        \SUBBYTES[0].a/w3306 ) );
  AND U386 ( .A(\SUBBYTES[0].a/w3270 ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3304 ) );
  AND U387 ( .A(\SUBBYTES[0].a/w3396 ), .B(n65), .Z(\SUBBYTES[0].a/w3303 ) );
  XNOR U388 ( .A(\w1[0][1] ), .B(n72), .Z(n65) );
  XOR U389 ( .A(g_input[1]), .B(state[1]), .Z(\w1[0][1] ) );
  AND U390 ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3271 ), .Z(
        \SUBBYTES[0].a/w3299 ) );
  XOR U391 ( .A(g_input[0]), .B(state[0]), .Z(\w1[0][0] ) );
  AND U392 ( .A(\SUBBYTES[0].a/w3272 ), .B(\SUBBYTES[0].a/w3268 ), .Z(
        \SUBBYTES[0].a/w3297 ) );
  AND U393 ( .A(\SUBBYTES[0].a/w3357 ), .B(\SUBBYTES[0].a/w3389 ), .Z(
        \SUBBYTES[0].a/w3296 ) );
  AND U394 ( .A(\SUBBYTES[0].a/w3378 ), .B(n69), .Z(\SUBBYTES[0].a/w3291 ) );
  XOR U395 ( .A(\w1[0][4] ), .B(\w1[0][7] ), .Z(n69) );
  ANDN U396 ( .A(\SUBBYTES[0].a/w3379 ), .B(n70), .Z(\SUBBYTES[0].a/w3289 ) );
  XNOR U397 ( .A(\w1[0][2] ), .B(\w1[0][7] ), .Z(n70) );
  IV U398 ( .A(n72), .Z(\w1[0][7] ) );
  XNOR U399 ( .A(g_input[7]), .B(state[7]), .Z(n72) );
  AND U400 ( .A(\SUBBYTES[0].a/w3381 ), .B(n71), .Z(\SUBBYTES[0].a/w3288 ) );
  XOR U401 ( .A(\w1[0][2] ), .B(\w1[0][4] ), .Z(n71) );
  XOR U402 ( .A(g_input[4]), .B(state[4]), .Z(\w1[0][4] ) );
  XOR U403 ( .A(g_input[2]), .B(state[2]), .Z(\w1[0][2] ) );
  AND U404 ( .A(n73), .B(\SUBBYTES[0].a/w3058 ), .Z(\SUBBYTES[0].a/w3193 ) );
  AND U405 ( .A(n74), .B(\SUBBYTES[0].a/w3059 ), .Z(\SUBBYTES[0].a/w3191 ) );
  AND U406 ( .A(\SUBBYTES[0].a/w3189 ), .B(n75), .Z(\SUBBYTES[0].a/w3190 ) );
  ANDN U407 ( .A(\w1[0][8] ), .B(n76), .Z(\SUBBYTES[0].a/w3186 ) );
  AND U408 ( .A(n77), .B(\SUBBYTES[0].a/w3061 ), .Z(\SUBBYTES[0].a/w3184 ) );
  AND U409 ( .A(\SUBBYTES[0].a/w3182 ), .B(n78), .Z(\SUBBYTES[0].a/w3183 ) );
  XOR U410 ( .A(\SUBBYTES[0].a/w3126 ), .B(\SUBBYTES[0].a/n149 ), .Z(n78) );
  AND U411 ( .A(\SUBBYTES[0].a/w3169 ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/w3178 ) );
  AND U412 ( .A(\SUBBYTES[0].a/w3170 ), .B(\SUBBYTES[0].a/w3172 ), .Z(
        \SUBBYTES[0].a/w3176 ) );
  AND U413 ( .A(\SUBBYTES[0].a/w3173 ), .B(\SUBBYTES[0].a/w3174 ), .Z(
        \SUBBYTES[0].a/w3175 ) );
  AND U414 ( .A(\SUBBYTES[0].a/w3062 ), .B(n73), .Z(\SUBBYTES[0].a/w3161 ) );
  XOR U415 ( .A(\SUBBYTES[0].a/w3130 ), .B(n15), .Z(n73) );
  AND U416 ( .A(\SUBBYTES[0].a/w3063 ), .B(n74), .Z(\SUBBYTES[0].a/w3159 ) );
  XOR U417 ( .A(\SUBBYTES[0].a/n150 ), .B(\SUBBYTES[0].a/w3130 ), .Z(n74) );
  AND U418 ( .A(n79), .B(n75), .Z(\SUBBYTES[0].a/w3158 ) );
  XOR U419 ( .A(n15), .B(\SUBBYTES[0].a/n150 ), .Z(n75) );
  ANDN U420 ( .A(\SUBBYTES[0].a/w3064 ), .B(n76), .Z(\SUBBYTES[0].a/w3154 ) );
  XNOR U421 ( .A(\SUBBYTES[0].a/w3123 ), .B(\SUBBYTES[0].a/w3126 ), .Z(n76) );
  AND U422 ( .A(\SUBBYTES[0].a/w3065 ), .B(n77), .Z(\SUBBYTES[0].a/w3152 ) );
  XNOR U423 ( .A(n80), .B(\SUBBYTES[0].a/w3123 ), .Z(n77) );
  AND U424 ( .A(\SUBBYTES[0].a/w3150 ), .B(n81), .Z(\SUBBYTES[0].a/w3151 ) );
  XOR U425 ( .A(n82), .B(n80), .Z(n81) );
  IV U426 ( .A(\SUBBYTES[0].a/n149 ), .Z(n80) );
  AND U427 ( .A(n83), .B(\SUBBYTES[0].a/w3169 ), .Z(\SUBBYTES[0].a/w3146 ) );
  ANDN U428 ( .A(\SUBBYTES[0].a/w3170 ), .B(n84), .Z(\SUBBYTES[0].a/w3144 ) );
  AND U429 ( .A(n85), .B(\SUBBYTES[0].a/w3173 ), .Z(\SUBBYTES[0].a/w3143 ) );
  AND U430 ( .A(\SUBBYTES[0].a/w3129 ), .B(\SUBBYTES[0].a/w3128 ), .Z(
        \SUBBYTES[0].a/w3130 ) );
  IV U431 ( .A(n82), .Z(\SUBBYTES[0].a/w3126 ) );
  NAND U432 ( .A(\SUBBYTES[0].a/w3105 ), .B(\SUBBYTES[0].a/w3120 ), .Z(n82) );
  AND U433 ( .A(\SUBBYTES[0].a/w3122 ), .B(\SUBBYTES[0].a/w3128 ), .Z(
        \SUBBYTES[0].a/w3123 ) );
  AND U434 ( .A(\SUBBYTES[0].a/w3107 ), .B(\SUBBYTES[0].a/w3105 ), .Z(
        \SUBBYTES[0].a/w3117 ) );
  AND U435 ( .A(\SUBBYTES[0].a/w3108 ), .B(\SUBBYTES[0].a/w3106 ), .Z(
        \SUBBYTES[0].a/w3115 ) );
  AND U436 ( .A(\SUBBYTES[0].a/w3122 ), .B(\SUBBYTES[0].a/w3129 ), .Z(
        \SUBBYTES[0].a/w3114 ) );
  AND U437 ( .A(\SUBBYTES[0].a/w3062 ), .B(\SUBBYTES[0].a/w3058 ), .Z(
        \SUBBYTES[0].a/w3099 ) );
  AND U438 ( .A(\SUBBYTES[0].a/w3063 ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3097 ) );
  AND U439 ( .A(\SUBBYTES[0].a/w3189 ), .B(n79), .Z(\SUBBYTES[0].a/w3096 ) );
  XNOR U440 ( .A(n86), .B(\w1[0][9] ), .Z(n79) );
  XOR U441 ( .A(g_input[9]), .B(state[9]), .Z(\w1[0][9] ) );
  AND U442 ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3064 ), .Z(
        \SUBBYTES[0].a/w3092 ) );
  XOR U443 ( .A(g_input[8]), .B(state[8]), .Z(\w1[0][8] ) );
  AND U444 ( .A(\SUBBYTES[0].a/w3065 ), .B(\SUBBYTES[0].a/w3061 ), .Z(
        \SUBBYTES[0].a/w3090 ) );
  AND U445 ( .A(\SUBBYTES[0].a/w3150 ), .B(\SUBBYTES[0].a/w3182 ), .Z(
        \SUBBYTES[0].a/w3089 ) );
  AND U446 ( .A(\SUBBYTES[0].a/w3171 ), .B(n83), .Z(\SUBBYTES[0].a/w3084 ) );
  XOR U447 ( .A(\w1[0][12] ), .B(\w1[0][15] ), .Z(n83) );
  ANDN U448 ( .A(\SUBBYTES[0].a/w3172 ), .B(n84), .Z(\SUBBYTES[0].a/w3082 ) );
  XNOR U449 ( .A(\w1[0][10] ), .B(\w1[0][15] ), .Z(n84) );
  IV U450 ( .A(n86), .Z(\w1[0][15] ) );
  XNOR U451 ( .A(g_input[15]), .B(state[15]), .Z(n86) );
  AND U452 ( .A(\SUBBYTES[0].a/w3174 ), .B(n85), .Z(\SUBBYTES[0].a/w3081 ) );
  XOR U453 ( .A(\w1[0][10] ), .B(\w1[0][12] ), .Z(n85) );
  XOR U454 ( .A(g_input[12]), .B(state[12]), .Z(\w1[0][12] ) );
  XOR U455 ( .A(g_input[10]), .B(state[10]), .Z(\w1[0][10] ) );
  AND U456 ( .A(n87), .B(\SUBBYTES[0].a/w2851 ), .Z(\SUBBYTES[0].a/w2986 ) );
  AND U457 ( .A(n88), .B(\SUBBYTES[0].a/w2852 ), .Z(\SUBBYTES[0].a/w2984 ) );
  AND U458 ( .A(\SUBBYTES[0].a/w2982 ), .B(n89), .Z(\SUBBYTES[0].a/w2983 ) );
  ANDN U459 ( .A(\w1[0][16] ), .B(n90), .Z(\SUBBYTES[0].a/w2979 ) );
  AND U460 ( .A(n91), .B(\SUBBYTES[0].a/w2854 ), .Z(\SUBBYTES[0].a/w2977 ) );
  AND U461 ( .A(\SUBBYTES[0].a/w2975 ), .B(n92), .Z(\SUBBYTES[0].a/w2976 ) );
  XOR U462 ( .A(\SUBBYTES[0].a/w2919 ), .B(\SUBBYTES[0].a/n139 ), .Z(n92) );
  AND U463 ( .A(\SUBBYTES[0].a/w2962 ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/w2971 ) );
  AND U464 ( .A(\SUBBYTES[0].a/w2963 ), .B(\SUBBYTES[0].a/w2965 ), .Z(
        \SUBBYTES[0].a/w2969 ) );
  AND U465 ( .A(\SUBBYTES[0].a/w2966 ), .B(\SUBBYTES[0].a/w2967 ), .Z(
        \SUBBYTES[0].a/w2968 ) );
  AND U466 ( .A(\SUBBYTES[0].a/w2855 ), .B(n87), .Z(\SUBBYTES[0].a/w2954 ) );
  XOR U467 ( .A(\SUBBYTES[0].a/w2923 ), .B(n14), .Z(n87) );
  AND U468 ( .A(\SUBBYTES[0].a/w2856 ), .B(n88), .Z(\SUBBYTES[0].a/w2952 ) );
  XOR U469 ( .A(\SUBBYTES[0].a/n140 ), .B(\SUBBYTES[0].a/w2923 ), .Z(n88) );
  AND U470 ( .A(n93), .B(n89), .Z(\SUBBYTES[0].a/w2951 ) );
  XOR U471 ( .A(n14), .B(\SUBBYTES[0].a/n140 ), .Z(n89) );
  AND U472 ( .A(n94), .B(\SUBBYTES[0].a/w160 ), .Z(\SUBBYTES[0].a/w295 ) );
  ANDN U473 ( .A(\SUBBYTES[0].a/w2857 ), .B(n90), .Z(\SUBBYTES[0].a/w2947 ) );
  XNOR U474 ( .A(\SUBBYTES[0].a/w2916 ), .B(\SUBBYTES[0].a/w2919 ), .Z(n90) );
  AND U475 ( .A(\SUBBYTES[0].a/w2858 ), .B(n91), .Z(\SUBBYTES[0].a/w2945 ) );
  XNOR U476 ( .A(n95), .B(\SUBBYTES[0].a/w2916 ), .Z(n91) );
  AND U477 ( .A(\SUBBYTES[0].a/w2943 ), .B(n96), .Z(\SUBBYTES[0].a/w2944 ) );
  XOR U478 ( .A(n97), .B(n95), .Z(n96) );
  IV U479 ( .A(\SUBBYTES[0].a/n139 ), .Z(n95) );
  AND U480 ( .A(n98), .B(\SUBBYTES[0].a/w2962 ), .Z(\SUBBYTES[0].a/w2939 ) );
  ANDN U481 ( .A(\SUBBYTES[0].a/w2963 ), .B(n99), .Z(\SUBBYTES[0].a/w2937 ) );
  AND U482 ( .A(n100), .B(\SUBBYTES[0].a/w2966 ), .Z(\SUBBYTES[0].a/w2936 ) );
  AND U483 ( .A(n101), .B(\SUBBYTES[0].a/w161 ), .Z(\SUBBYTES[0].a/w293 ) );
  AND U484 ( .A(\SUBBYTES[0].a/w2922 ), .B(\SUBBYTES[0].a/w2921 ), .Z(
        \SUBBYTES[0].a/w2923 ) );
  AND U485 ( .A(\SUBBYTES[0].a/w291 ), .B(n102), .Z(\SUBBYTES[0].a/w292 ) );
  IV U486 ( .A(n97), .Z(\SUBBYTES[0].a/w2919 ) );
  NAND U487 ( .A(\SUBBYTES[0].a/w2898 ), .B(\SUBBYTES[0].a/w2913 ), .Z(n97) );
  AND U488 ( .A(\SUBBYTES[0].a/w2915 ), .B(\SUBBYTES[0].a/w2921 ), .Z(
        \SUBBYTES[0].a/w2916 ) );
  AND U489 ( .A(\SUBBYTES[0].a/w2900 ), .B(\SUBBYTES[0].a/w2898 ), .Z(
        \SUBBYTES[0].a/w2910 ) );
  AND U490 ( .A(\SUBBYTES[0].a/w2901 ), .B(\SUBBYTES[0].a/w2899 ), .Z(
        \SUBBYTES[0].a/w2908 ) );
  AND U491 ( .A(\SUBBYTES[0].a/w2915 ), .B(\SUBBYTES[0].a/w2922 ), .Z(
        \SUBBYTES[0].a/w2907 ) );
  AND U492 ( .A(\SUBBYTES[0].a/w2855 ), .B(\SUBBYTES[0].a/w2851 ), .Z(
        \SUBBYTES[0].a/w2892 ) );
  AND U493 ( .A(\SUBBYTES[0].a/w2856 ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2890 ) );
  AND U494 ( .A(\SUBBYTES[0].a/w2982 ), .B(n93), .Z(\SUBBYTES[0].a/w2889 ) );
  XNOR U495 ( .A(\w1[0][17] ), .B(n103), .Z(n93) );
  XOR U496 ( .A(g_input[17]), .B(state[17]), .Z(\w1[0][17] ) );
  AND U497 ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2857 ), .Z(
        \SUBBYTES[0].a/w2885 ) );
  XOR U498 ( .A(g_input[16]), .B(state[16]), .Z(\w1[0][16] ) );
  AND U499 ( .A(\SUBBYTES[0].a/w2858 ), .B(\SUBBYTES[0].a/w2854 ), .Z(
        \SUBBYTES[0].a/w2883 ) );
  AND U500 ( .A(\SUBBYTES[0].a/w2943 ), .B(\SUBBYTES[0].a/w2975 ), .Z(
        \SUBBYTES[0].a/w2882 ) );
  ANDN U501 ( .A(\w1[0][120] ), .B(n104), .Z(\SUBBYTES[0].a/w288 ) );
  AND U502 ( .A(\SUBBYTES[0].a/w2964 ), .B(n98), .Z(\SUBBYTES[0].a/w2877 ) );
  XOR U503 ( .A(\w1[0][20] ), .B(\w1[0][23] ), .Z(n98) );
  ANDN U504 ( .A(\SUBBYTES[0].a/w2965 ), .B(n99), .Z(\SUBBYTES[0].a/w2875 ) );
  XNOR U505 ( .A(\w1[0][18] ), .B(\w1[0][23] ), .Z(n99) );
  IV U506 ( .A(n103), .Z(\w1[0][23] ) );
  XNOR U507 ( .A(g_input[23]), .B(state[23]), .Z(n103) );
  AND U508 ( .A(\SUBBYTES[0].a/w2967 ), .B(n100), .Z(\SUBBYTES[0].a/w2874 ) );
  XOR U509 ( .A(\w1[0][18] ), .B(\w1[0][20] ), .Z(n100) );
  XOR U510 ( .A(g_input[20]), .B(state[20]), .Z(\w1[0][20] ) );
  XOR U511 ( .A(g_input[18]), .B(state[18]), .Z(\w1[0][18] ) );
  AND U512 ( .A(n105), .B(\SUBBYTES[0].a/w163 ), .Z(\SUBBYTES[0].a/w286 ) );
  AND U513 ( .A(\SUBBYTES[0].a/w284 ), .B(n106), .Z(\SUBBYTES[0].a/w285 ) );
  XOR U514 ( .A(\SUBBYTES[0].a/w228 ), .B(\SUBBYTES[0].a/n9 ), .Z(n106) );
  AND U515 ( .A(\SUBBYTES[0].a/w271 ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/w280 ) );
  AND U516 ( .A(\SUBBYTES[0].a/w272 ), .B(\SUBBYTES[0].a/w274 ), .Z(
        \SUBBYTES[0].a/w278 ) );
  AND U517 ( .A(n107), .B(\SUBBYTES[0].a/w2644 ), .Z(\SUBBYTES[0].a/w2779 ) );
  AND U518 ( .A(n108), .B(\SUBBYTES[0].a/w2645 ), .Z(\SUBBYTES[0].a/w2777 ) );
  AND U519 ( .A(\SUBBYTES[0].a/w2775 ), .B(n109), .Z(\SUBBYTES[0].a/w2776 ) );
  ANDN U520 ( .A(\w1[0][24] ), .B(n110), .Z(\SUBBYTES[0].a/w2772 ) );
  AND U521 ( .A(n111), .B(\SUBBYTES[0].a/w2647 ), .Z(\SUBBYTES[0].a/w2770 ) );
  AND U522 ( .A(\SUBBYTES[0].a/w275 ), .B(\SUBBYTES[0].a/w276 ), .Z(
        \SUBBYTES[0].a/w277 ) );
  AND U523 ( .A(\SUBBYTES[0].a/w2768 ), .B(n112), .Z(\SUBBYTES[0].a/w2769 ) );
  XOR U524 ( .A(\SUBBYTES[0].a/w2712 ), .B(\SUBBYTES[0].a/n129 ), .Z(n112) );
  AND U525 ( .A(\SUBBYTES[0].a/w2755 ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/w2764 ) );
  AND U526 ( .A(\SUBBYTES[0].a/w2756 ), .B(\SUBBYTES[0].a/w2758 ), .Z(
        \SUBBYTES[0].a/w2762 ) );
  AND U527 ( .A(\SUBBYTES[0].a/w2759 ), .B(\SUBBYTES[0].a/w2760 ), .Z(
        \SUBBYTES[0].a/w2761 ) );
  AND U528 ( .A(\SUBBYTES[0].a/w2648 ), .B(n107), .Z(\SUBBYTES[0].a/w2747 ) );
  XOR U529 ( .A(\SUBBYTES[0].a/w2716 ), .B(n13), .Z(n107) );
  AND U530 ( .A(\SUBBYTES[0].a/w2649 ), .B(n108), .Z(\SUBBYTES[0].a/w2745 ) );
  XOR U531 ( .A(\SUBBYTES[0].a/n130 ), .B(\SUBBYTES[0].a/w2716 ), .Z(n108) );
  AND U532 ( .A(n113), .B(n109), .Z(\SUBBYTES[0].a/w2744 ) );
  XOR U533 ( .A(n13), .B(\SUBBYTES[0].a/n130 ), .Z(n109) );
  ANDN U534 ( .A(\SUBBYTES[0].a/w2650 ), .B(n110), .Z(\SUBBYTES[0].a/w2740 )
         );
  XNOR U535 ( .A(\SUBBYTES[0].a/w2709 ), .B(\SUBBYTES[0].a/w2712 ), .Z(n110)
         );
  AND U536 ( .A(\SUBBYTES[0].a/w2651 ), .B(n111), .Z(\SUBBYTES[0].a/w2738 ) );
  XNOR U537 ( .A(n114), .B(\SUBBYTES[0].a/w2709 ), .Z(n111) );
  AND U538 ( .A(\SUBBYTES[0].a/w2736 ), .B(n115), .Z(\SUBBYTES[0].a/w2737 ) );
  XOR U539 ( .A(n116), .B(n114), .Z(n115) );
  IV U540 ( .A(\SUBBYTES[0].a/n129 ), .Z(n114) );
  AND U541 ( .A(n117), .B(\SUBBYTES[0].a/w2755 ), .Z(\SUBBYTES[0].a/w2732 ) );
  ANDN U542 ( .A(\SUBBYTES[0].a/w2756 ), .B(n118), .Z(\SUBBYTES[0].a/w2730 )
         );
  AND U543 ( .A(n119), .B(\SUBBYTES[0].a/w2759 ), .Z(\SUBBYTES[0].a/w2729 ) );
  AND U544 ( .A(\SUBBYTES[0].a/w2715 ), .B(\SUBBYTES[0].a/w2714 ), .Z(
        \SUBBYTES[0].a/w2716 ) );
  IV U545 ( .A(n116), .Z(\SUBBYTES[0].a/w2712 ) );
  NAND U546 ( .A(\SUBBYTES[0].a/w2691 ), .B(\SUBBYTES[0].a/w2706 ), .Z(n116)
         );
  AND U547 ( .A(\SUBBYTES[0].a/w2708 ), .B(\SUBBYTES[0].a/w2714 ), .Z(
        \SUBBYTES[0].a/w2709 ) );
  AND U548 ( .A(\SUBBYTES[0].a/w2693 ), .B(\SUBBYTES[0].a/w2691 ), .Z(
        \SUBBYTES[0].a/w2703 ) );
  AND U549 ( .A(\SUBBYTES[0].a/w2694 ), .B(\SUBBYTES[0].a/w2692 ), .Z(
        \SUBBYTES[0].a/w2701 ) );
  AND U550 ( .A(\SUBBYTES[0].a/w2708 ), .B(\SUBBYTES[0].a/w2715 ), .Z(
        \SUBBYTES[0].a/w2700 ) );
  AND U551 ( .A(\SUBBYTES[0].a/w2648 ), .B(\SUBBYTES[0].a/w2644 ), .Z(
        \SUBBYTES[0].a/w2685 ) );
  AND U552 ( .A(\SUBBYTES[0].a/w2649 ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2683 ) );
  AND U553 ( .A(\SUBBYTES[0].a/w2775 ), .B(n113), .Z(\SUBBYTES[0].a/w2682 ) );
  XNOR U554 ( .A(\w1[0][25] ), .B(n120), .Z(n113) );
  XOR U555 ( .A(g_input[25]), .B(state[25]), .Z(\w1[0][25] ) );
  AND U556 ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2650 ), .Z(
        \SUBBYTES[0].a/w2678 ) );
  XOR U557 ( .A(g_input[24]), .B(state[24]), .Z(\w1[0][24] ) );
  AND U558 ( .A(\SUBBYTES[0].a/w2651 ), .B(\SUBBYTES[0].a/w2647 ), .Z(
        \SUBBYTES[0].a/w2676 ) );
  AND U559 ( .A(\SUBBYTES[0].a/w2736 ), .B(\SUBBYTES[0].a/w2768 ), .Z(
        \SUBBYTES[0].a/w2675 ) );
  AND U560 ( .A(\SUBBYTES[0].a/w2757 ), .B(n117), .Z(\SUBBYTES[0].a/w2670 ) );
  XOR U561 ( .A(\w1[0][28] ), .B(\w1[0][31] ), .Z(n117) );
  ANDN U562 ( .A(\SUBBYTES[0].a/w2758 ), .B(n118), .Z(\SUBBYTES[0].a/w2668 )
         );
  XNOR U563 ( .A(\w1[0][26] ), .B(\w1[0][31] ), .Z(n118) );
  IV U564 ( .A(n120), .Z(\w1[0][31] ) );
  XNOR U565 ( .A(g_input[31]), .B(state[31]), .Z(n120) );
  AND U566 ( .A(\SUBBYTES[0].a/w2760 ), .B(n119), .Z(\SUBBYTES[0].a/w2667 ) );
  XOR U567 ( .A(\w1[0][26] ), .B(\w1[0][28] ), .Z(n119) );
  XOR U568 ( .A(g_input[28]), .B(state[28]), .Z(\w1[0][28] ) );
  XOR U569 ( .A(g_input[26]), .B(state[26]), .Z(\w1[0][26] ) );
  AND U570 ( .A(\SUBBYTES[0].a/w164 ), .B(n94), .Z(\SUBBYTES[0].a/w263 ) );
  XOR U571 ( .A(\SUBBYTES[0].a/w232 ), .B(n1), .Z(n94) );
  AND U572 ( .A(\SUBBYTES[0].a/w165 ), .B(n101), .Z(\SUBBYTES[0].a/w261 ) );
  XOR U573 ( .A(\SUBBYTES[0].a/n10 ), .B(\SUBBYTES[0].a/w232 ), .Z(n101) );
  AND U574 ( .A(n121), .B(n102), .Z(\SUBBYTES[0].a/w260 ) );
  XOR U575 ( .A(n1), .B(\SUBBYTES[0].a/n10 ), .Z(n102) );
  AND U576 ( .A(n122), .B(\SUBBYTES[0].a/w2437 ), .Z(\SUBBYTES[0].a/w2572 ) );
  AND U577 ( .A(n123), .B(\SUBBYTES[0].a/w2438 ), .Z(\SUBBYTES[0].a/w2570 ) );
  AND U578 ( .A(\SUBBYTES[0].a/w2568 ), .B(n124), .Z(\SUBBYTES[0].a/w2569 ) );
  ANDN U579 ( .A(\w1[0][32] ), .B(n125), .Z(\SUBBYTES[0].a/w2565 ) );
  AND U580 ( .A(n126), .B(\SUBBYTES[0].a/w2440 ), .Z(\SUBBYTES[0].a/w2563 ) );
  AND U581 ( .A(\SUBBYTES[0].a/w2561 ), .B(n127), .Z(\SUBBYTES[0].a/w2562 ) );
  XOR U582 ( .A(\SUBBYTES[0].a/w2505 ), .B(\SUBBYTES[0].a/n119 ), .Z(n127) );
  ANDN U583 ( .A(\SUBBYTES[0].a/w166 ), .B(n104), .Z(\SUBBYTES[0].a/w256 ) );
  XNOR U584 ( .A(\SUBBYTES[0].a/w225 ), .B(\SUBBYTES[0].a/w228 ), .Z(n104) );
  AND U585 ( .A(\SUBBYTES[0].a/w2548 ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/w2557 ) );
  AND U586 ( .A(\SUBBYTES[0].a/w2549 ), .B(\SUBBYTES[0].a/w2551 ), .Z(
        \SUBBYTES[0].a/w2555 ) );
  AND U587 ( .A(\SUBBYTES[0].a/w2552 ), .B(\SUBBYTES[0].a/w2553 ), .Z(
        \SUBBYTES[0].a/w2554 ) );
  AND U588 ( .A(\SUBBYTES[0].a/w2441 ), .B(n122), .Z(\SUBBYTES[0].a/w2540 ) );
  XOR U589 ( .A(\SUBBYTES[0].a/w2509 ), .B(n12), .Z(n122) );
  AND U590 ( .A(\SUBBYTES[0].a/w167 ), .B(n105), .Z(\SUBBYTES[0].a/w254 ) );
  XNOR U591 ( .A(n128), .B(\SUBBYTES[0].a/w225 ), .Z(n105) );
  AND U592 ( .A(\SUBBYTES[0].a/w2442 ), .B(n123), .Z(\SUBBYTES[0].a/w2538 ) );
  XOR U593 ( .A(\SUBBYTES[0].a/n120 ), .B(\SUBBYTES[0].a/w2509 ), .Z(n123) );
  AND U594 ( .A(n129), .B(n124), .Z(\SUBBYTES[0].a/w2537 ) );
  XOR U595 ( .A(n12), .B(\SUBBYTES[0].a/n120 ), .Z(n124) );
  ANDN U596 ( .A(\SUBBYTES[0].a/w2443 ), .B(n125), .Z(\SUBBYTES[0].a/w2533 )
         );
  XNOR U597 ( .A(\SUBBYTES[0].a/w2502 ), .B(\SUBBYTES[0].a/w2505 ), .Z(n125)
         );
  AND U598 ( .A(\SUBBYTES[0].a/w2444 ), .B(n126), .Z(\SUBBYTES[0].a/w2531 ) );
  XNOR U599 ( .A(n130), .B(\SUBBYTES[0].a/w2502 ), .Z(n126) );
  AND U600 ( .A(\SUBBYTES[0].a/w2529 ), .B(n131), .Z(\SUBBYTES[0].a/w2530 ) );
  XOR U601 ( .A(n132), .B(n130), .Z(n131) );
  IV U602 ( .A(\SUBBYTES[0].a/n119 ), .Z(n130) );
  AND U603 ( .A(\SUBBYTES[0].a/w252 ), .B(n133), .Z(\SUBBYTES[0].a/w253 ) );
  XOR U604 ( .A(n134), .B(n128), .Z(n133) );
  IV U605 ( .A(\SUBBYTES[0].a/n9 ), .Z(n128) );
  AND U606 ( .A(n135), .B(\SUBBYTES[0].a/w2548 ), .Z(\SUBBYTES[0].a/w2525 ) );
  ANDN U607 ( .A(\SUBBYTES[0].a/w2549 ), .B(n136), .Z(\SUBBYTES[0].a/w2523 )
         );
  AND U608 ( .A(n137), .B(\SUBBYTES[0].a/w2552 ), .Z(\SUBBYTES[0].a/w2522 ) );
  AND U609 ( .A(\SUBBYTES[0].a/w2508 ), .B(\SUBBYTES[0].a/w2507 ), .Z(
        \SUBBYTES[0].a/w2509 ) );
  IV U610 ( .A(n132), .Z(\SUBBYTES[0].a/w2505 ) );
  NAND U611 ( .A(\SUBBYTES[0].a/w2484 ), .B(\SUBBYTES[0].a/w2499 ), .Z(n132)
         );
  AND U612 ( .A(\SUBBYTES[0].a/w2501 ), .B(\SUBBYTES[0].a/w2507 ), .Z(
        \SUBBYTES[0].a/w2502 ) );
  AND U613 ( .A(\SUBBYTES[0].a/w2486 ), .B(\SUBBYTES[0].a/w2484 ), .Z(
        \SUBBYTES[0].a/w2496 ) );
  AND U614 ( .A(\SUBBYTES[0].a/w2487 ), .B(\SUBBYTES[0].a/w2485 ), .Z(
        \SUBBYTES[0].a/w2494 ) );
  AND U615 ( .A(\SUBBYTES[0].a/w2501 ), .B(\SUBBYTES[0].a/w2508 ), .Z(
        \SUBBYTES[0].a/w2493 ) );
  AND U616 ( .A(n138), .B(\SUBBYTES[0].a/w271 ), .Z(\SUBBYTES[0].a/w248 ) );
  AND U617 ( .A(\SUBBYTES[0].a/w2441 ), .B(\SUBBYTES[0].a/w2437 ), .Z(
        \SUBBYTES[0].a/w2478 ) );
  AND U618 ( .A(\SUBBYTES[0].a/w2442 ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2476 ) );
  AND U619 ( .A(\SUBBYTES[0].a/w2568 ), .B(n129), .Z(\SUBBYTES[0].a/w2475 ) );
  XNOR U620 ( .A(\w1[0][33] ), .B(n139), .Z(n129) );
  XOR U621 ( .A(g_input[33]), .B(state[33]), .Z(\w1[0][33] ) );
  AND U622 ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2443 ), .Z(
        \SUBBYTES[0].a/w2471 ) );
  XOR U623 ( .A(g_input[32]), .B(state[32]), .Z(\w1[0][32] ) );
  AND U624 ( .A(\SUBBYTES[0].a/w2444 ), .B(\SUBBYTES[0].a/w2440 ), .Z(
        \SUBBYTES[0].a/w2469 ) );
  AND U625 ( .A(\SUBBYTES[0].a/w2529 ), .B(\SUBBYTES[0].a/w2561 ), .Z(
        \SUBBYTES[0].a/w2468 ) );
  AND U626 ( .A(\SUBBYTES[0].a/w2550 ), .B(n135), .Z(\SUBBYTES[0].a/w2463 ) );
  XOR U627 ( .A(\w1[0][36] ), .B(\w1[0][39] ), .Z(n135) );
  ANDN U628 ( .A(\SUBBYTES[0].a/w2551 ), .B(n136), .Z(\SUBBYTES[0].a/w2461 )
         );
  XNOR U629 ( .A(\w1[0][34] ), .B(\w1[0][39] ), .Z(n136) );
  IV U630 ( .A(n139), .Z(\w1[0][39] ) );
  XNOR U631 ( .A(g_input[39]), .B(state[39]), .Z(n139) );
  AND U632 ( .A(\SUBBYTES[0].a/w2553 ), .B(n137), .Z(\SUBBYTES[0].a/w2460 ) );
  XOR U633 ( .A(\w1[0][34] ), .B(\w1[0][36] ), .Z(n137) );
  XOR U634 ( .A(g_input[36]), .B(state[36]), .Z(\w1[0][36] ) );
  XOR U635 ( .A(g_input[34]), .B(state[34]), .Z(\w1[0][34] ) );
  ANDN U636 ( .A(\SUBBYTES[0].a/w272 ), .B(n140), .Z(\SUBBYTES[0].a/w246 ) );
  AND U637 ( .A(n141), .B(\SUBBYTES[0].a/w275 ), .Z(\SUBBYTES[0].a/w245 ) );
  AND U638 ( .A(n142), .B(\SUBBYTES[0].a/w2230 ), .Z(\SUBBYTES[0].a/w2365 ) );
  AND U639 ( .A(n143), .B(\SUBBYTES[0].a/w2231 ), .Z(\SUBBYTES[0].a/w2363 ) );
  AND U640 ( .A(\SUBBYTES[0].a/w2361 ), .B(n144), .Z(\SUBBYTES[0].a/w2362 ) );
  ANDN U641 ( .A(\w1[0][40] ), .B(n145), .Z(\SUBBYTES[0].a/w2358 ) );
  AND U642 ( .A(n146), .B(\SUBBYTES[0].a/w2233 ), .Z(\SUBBYTES[0].a/w2356 ) );
  AND U643 ( .A(\SUBBYTES[0].a/w2354 ), .B(n147), .Z(\SUBBYTES[0].a/w2355 ) );
  XOR U644 ( .A(\SUBBYTES[0].a/w2298 ), .B(\SUBBYTES[0].a/n109 ), .Z(n147) );
  AND U645 ( .A(\SUBBYTES[0].a/w2341 ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/w2350 ) );
  AND U646 ( .A(\SUBBYTES[0].a/w2342 ), .B(\SUBBYTES[0].a/w2344 ), .Z(
        \SUBBYTES[0].a/w2348 ) );
  AND U647 ( .A(\SUBBYTES[0].a/w2345 ), .B(\SUBBYTES[0].a/w2346 ), .Z(
        \SUBBYTES[0].a/w2347 ) );
  AND U648 ( .A(\SUBBYTES[0].a/w2234 ), .B(n142), .Z(\SUBBYTES[0].a/w2333 ) );
  XOR U649 ( .A(\SUBBYTES[0].a/w2302 ), .B(n11), .Z(n142) );
  AND U650 ( .A(\SUBBYTES[0].a/w2235 ), .B(n143), .Z(\SUBBYTES[0].a/w2331 ) );
  XOR U651 ( .A(\SUBBYTES[0].a/n110 ), .B(\SUBBYTES[0].a/w2302 ), .Z(n143) );
  AND U652 ( .A(n148), .B(n144), .Z(\SUBBYTES[0].a/w2330 ) );
  XOR U653 ( .A(n11), .B(\SUBBYTES[0].a/n110 ), .Z(n144) );
  ANDN U654 ( .A(\SUBBYTES[0].a/w2236 ), .B(n145), .Z(\SUBBYTES[0].a/w2326 )
         );
  XNOR U655 ( .A(\SUBBYTES[0].a/w2295 ), .B(\SUBBYTES[0].a/w2298 ), .Z(n145)
         );
  AND U656 ( .A(\SUBBYTES[0].a/w2237 ), .B(n146), .Z(\SUBBYTES[0].a/w2324 ) );
  XNOR U657 ( .A(n149), .B(\SUBBYTES[0].a/w2295 ), .Z(n146) );
  AND U658 ( .A(\SUBBYTES[0].a/w2322 ), .B(n150), .Z(\SUBBYTES[0].a/w2323 ) );
  XOR U659 ( .A(n151), .B(n149), .Z(n150) );
  IV U660 ( .A(\SUBBYTES[0].a/n109 ), .Z(n149) );
  AND U661 ( .A(\SUBBYTES[0].a/w231 ), .B(\SUBBYTES[0].a/w230 ), .Z(
        \SUBBYTES[0].a/w232 ) );
  AND U662 ( .A(n152), .B(\SUBBYTES[0].a/w2341 ), .Z(\SUBBYTES[0].a/w2318 ) );
  ANDN U663 ( .A(\SUBBYTES[0].a/w2342 ), .B(n153), .Z(\SUBBYTES[0].a/w2316 )
         );
  AND U664 ( .A(n154), .B(\SUBBYTES[0].a/w2345 ), .Z(\SUBBYTES[0].a/w2315 ) );
  AND U665 ( .A(\SUBBYTES[0].a/w2301 ), .B(\SUBBYTES[0].a/w2300 ), .Z(
        \SUBBYTES[0].a/w2302 ) );
  IV U666 ( .A(n151), .Z(\SUBBYTES[0].a/w2298 ) );
  NAND U667 ( .A(\SUBBYTES[0].a/w2277 ), .B(\SUBBYTES[0].a/w2292 ), .Z(n151)
         );
  AND U668 ( .A(\SUBBYTES[0].a/w2294 ), .B(\SUBBYTES[0].a/w2300 ), .Z(
        \SUBBYTES[0].a/w2295 ) );
  AND U669 ( .A(\SUBBYTES[0].a/w2279 ), .B(\SUBBYTES[0].a/w2277 ), .Z(
        \SUBBYTES[0].a/w2289 ) );
  AND U670 ( .A(\SUBBYTES[0].a/w2280 ), .B(\SUBBYTES[0].a/w2278 ), .Z(
        \SUBBYTES[0].a/w2287 ) );
  AND U671 ( .A(\SUBBYTES[0].a/w2294 ), .B(\SUBBYTES[0].a/w2301 ), .Z(
        \SUBBYTES[0].a/w2286 ) );
  IV U672 ( .A(n134), .Z(\SUBBYTES[0].a/w228 ) );
  NAND U673 ( .A(\SUBBYTES[0].a/w207 ), .B(\SUBBYTES[0].a/w222 ), .Z(n134) );
  AND U674 ( .A(\SUBBYTES[0].a/w2234 ), .B(\SUBBYTES[0].a/w2230 ), .Z(
        \SUBBYTES[0].a/w2271 ) );
  AND U675 ( .A(\SUBBYTES[0].a/w2235 ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2269 ) );
  AND U676 ( .A(\SUBBYTES[0].a/w2361 ), .B(n148), .Z(\SUBBYTES[0].a/w2268 ) );
  XNOR U677 ( .A(\w1[0][41] ), .B(n155), .Z(n148) );
  XOR U678 ( .A(g_input[41]), .B(state[41]), .Z(\w1[0][41] ) );
  AND U679 ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2236 ), .Z(
        \SUBBYTES[0].a/w2264 ) );
  XOR U680 ( .A(g_input[40]), .B(state[40]), .Z(\w1[0][40] ) );
  AND U681 ( .A(\SUBBYTES[0].a/w2237 ), .B(\SUBBYTES[0].a/w2233 ), .Z(
        \SUBBYTES[0].a/w2262 ) );
  AND U682 ( .A(\SUBBYTES[0].a/w2322 ), .B(\SUBBYTES[0].a/w2354 ), .Z(
        \SUBBYTES[0].a/w2261 ) );
  AND U683 ( .A(\SUBBYTES[0].a/w2343 ), .B(n152), .Z(\SUBBYTES[0].a/w2256 ) );
  XOR U684 ( .A(\w1[0][44] ), .B(\w1[0][47] ), .Z(n152) );
  ANDN U685 ( .A(\SUBBYTES[0].a/w2344 ), .B(n153), .Z(\SUBBYTES[0].a/w2254 )
         );
  XNOR U686 ( .A(\w1[0][42] ), .B(\w1[0][47] ), .Z(n153) );
  IV U687 ( .A(n155), .Z(\w1[0][47] ) );
  XNOR U688 ( .A(g_input[47]), .B(state[47]), .Z(n155) );
  AND U689 ( .A(\SUBBYTES[0].a/w2346 ), .B(n154), .Z(\SUBBYTES[0].a/w2253 ) );
  XOR U690 ( .A(\w1[0][42] ), .B(\w1[0][44] ), .Z(n154) );
  XOR U691 ( .A(g_input[44]), .B(state[44]), .Z(\w1[0][44] ) );
  XOR U692 ( .A(g_input[42]), .B(state[42]), .Z(\w1[0][42] ) );
  AND U693 ( .A(\SUBBYTES[0].a/w224 ), .B(\SUBBYTES[0].a/w230 ), .Z(
        \SUBBYTES[0].a/w225 ) );
  AND U694 ( .A(\SUBBYTES[0].a/w209 ), .B(\SUBBYTES[0].a/w207 ), .Z(
        \SUBBYTES[0].a/w219 ) );
  AND U695 ( .A(\SUBBYTES[0].a/w210 ), .B(\SUBBYTES[0].a/w208 ), .Z(
        \SUBBYTES[0].a/w217 ) );
  AND U696 ( .A(\SUBBYTES[0].a/w224 ), .B(\SUBBYTES[0].a/w231 ), .Z(
        \SUBBYTES[0].a/w216 ) );
  AND U697 ( .A(n156), .B(\SUBBYTES[0].a/w2023 ), .Z(\SUBBYTES[0].a/w2158 ) );
  AND U698 ( .A(n157), .B(\SUBBYTES[0].a/w2024 ), .Z(\SUBBYTES[0].a/w2156 ) );
  AND U699 ( .A(\SUBBYTES[0].a/w2154 ), .B(n158), .Z(\SUBBYTES[0].a/w2155 ) );
  ANDN U700 ( .A(\w1[0][48] ), .B(n159), .Z(\SUBBYTES[0].a/w2151 ) );
  AND U701 ( .A(n160), .B(\SUBBYTES[0].a/w2026 ), .Z(\SUBBYTES[0].a/w2149 ) );
  AND U702 ( .A(\SUBBYTES[0].a/w2147 ), .B(n161), .Z(\SUBBYTES[0].a/w2148 ) );
  XOR U703 ( .A(\SUBBYTES[0].a/w2091 ), .B(\SUBBYTES[0].a/n99 ), .Z(n161) );
  AND U704 ( .A(\SUBBYTES[0].a/w2134 ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/w2143 ) );
  AND U705 ( .A(\SUBBYTES[0].a/w2135 ), .B(\SUBBYTES[0].a/w2137 ), .Z(
        \SUBBYTES[0].a/w2141 ) );
  AND U706 ( .A(\SUBBYTES[0].a/w2138 ), .B(\SUBBYTES[0].a/w2139 ), .Z(
        \SUBBYTES[0].a/w2140 ) );
  AND U707 ( .A(\SUBBYTES[0].a/w2027 ), .B(n156), .Z(\SUBBYTES[0].a/w2126 ) );
  XOR U708 ( .A(\SUBBYTES[0].a/w2095 ), .B(n10), .Z(n156) );
  AND U709 ( .A(\SUBBYTES[0].a/w2028 ), .B(n157), .Z(\SUBBYTES[0].a/w2124 ) );
  XOR U710 ( .A(\SUBBYTES[0].a/n100 ), .B(\SUBBYTES[0].a/w2095 ), .Z(n157) );
  AND U711 ( .A(n162), .B(n158), .Z(\SUBBYTES[0].a/w2123 ) );
  XOR U712 ( .A(n10), .B(\SUBBYTES[0].a/n100 ), .Z(n158) );
  ANDN U713 ( .A(\SUBBYTES[0].a/w2029 ), .B(n159), .Z(\SUBBYTES[0].a/w2119 )
         );
  XNOR U714 ( .A(\SUBBYTES[0].a/w2088 ), .B(\SUBBYTES[0].a/w2091 ), .Z(n159)
         );
  AND U715 ( .A(\SUBBYTES[0].a/w2030 ), .B(n160), .Z(\SUBBYTES[0].a/w2117 ) );
  XNOR U716 ( .A(n163), .B(\SUBBYTES[0].a/w2088 ), .Z(n160) );
  AND U717 ( .A(\SUBBYTES[0].a/w2115 ), .B(n164), .Z(\SUBBYTES[0].a/w2116 ) );
  XOR U718 ( .A(n165), .B(n163), .Z(n164) );
  IV U719 ( .A(\SUBBYTES[0].a/n99 ), .Z(n163) );
  AND U720 ( .A(n166), .B(\SUBBYTES[0].a/w2134 ), .Z(\SUBBYTES[0].a/w2111 ) );
  ANDN U721 ( .A(\SUBBYTES[0].a/w2135 ), .B(n167), .Z(\SUBBYTES[0].a/w2109 )
         );
  AND U722 ( .A(n168), .B(\SUBBYTES[0].a/w2138 ), .Z(\SUBBYTES[0].a/w2108 ) );
  AND U723 ( .A(\SUBBYTES[0].a/w2094 ), .B(\SUBBYTES[0].a/w2093 ), .Z(
        \SUBBYTES[0].a/w2095 ) );
  IV U724 ( .A(n165), .Z(\SUBBYTES[0].a/w2091 ) );
  NAND U725 ( .A(\SUBBYTES[0].a/w2070 ), .B(\SUBBYTES[0].a/w2085 ), .Z(n165)
         );
  AND U726 ( .A(\SUBBYTES[0].a/w2087 ), .B(\SUBBYTES[0].a/w2093 ), .Z(
        \SUBBYTES[0].a/w2088 ) );
  AND U727 ( .A(\SUBBYTES[0].a/w2072 ), .B(\SUBBYTES[0].a/w2070 ), .Z(
        \SUBBYTES[0].a/w2082 ) );
  AND U728 ( .A(\SUBBYTES[0].a/w2073 ), .B(\SUBBYTES[0].a/w2071 ), .Z(
        \SUBBYTES[0].a/w2080 ) );
  AND U729 ( .A(\SUBBYTES[0].a/w2087 ), .B(\SUBBYTES[0].a/w2094 ), .Z(
        \SUBBYTES[0].a/w2079 ) );
  AND U730 ( .A(\SUBBYTES[0].a/w2027 ), .B(\SUBBYTES[0].a/w2023 ), .Z(
        \SUBBYTES[0].a/w2064 ) );
  AND U731 ( .A(\SUBBYTES[0].a/w2028 ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2062 ) );
  AND U732 ( .A(\SUBBYTES[0].a/w2154 ), .B(n162), .Z(\SUBBYTES[0].a/w2061 ) );
  XNOR U733 ( .A(\w1[0][49] ), .B(n169), .Z(n162) );
  XOR U734 ( .A(g_input[49]), .B(state[49]), .Z(\w1[0][49] ) );
  AND U735 ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2029 ), .Z(
        \SUBBYTES[0].a/w2057 ) );
  XOR U736 ( .A(g_input[48]), .B(state[48]), .Z(\w1[0][48] ) );
  AND U737 ( .A(\SUBBYTES[0].a/w2030 ), .B(\SUBBYTES[0].a/w2026 ), .Z(
        \SUBBYTES[0].a/w2055 ) );
  AND U738 ( .A(\SUBBYTES[0].a/w2115 ), .B(\SUBBYTES[0].a/w2147 ), .Z(
        \SUBBYTES[0].a/w2054 ) );
  AND U739 ( .A(\SUBBYTES[0].a/w2136 ), .B(n166), .Z(\SUBBYTES[0].a/w2049 ) );
  XOR U740 ( .A(\w1[0][52] ), .B(\w1[0][55] ), .Z(n166) );
  ANDN U741 ( .A(\SUBBYTES[0].a/w2137 ), .B(n167), .Z(\SUBBYTES[0].a/w2047 )
         );
  XNOR U742 ( .A(\w1[0][50] ), .B(\w1[0][55] ), .Z(n167) );
  IV U743 ( .A(n169), .Z(\w1[0][55] ) );
  XNOR U744 ( .A(g_input[55]), .B(state[55]), .Z(n169) );
  AND U745 ( .A(\SUBBYTES[0].a/w2139 ), .B(n168), .Z(\SUBBYTES[0].a/w2046 ) );
  XOR U746 ( .A(\w1[0][50] ), .B(\w1[0][52] ), .Z(n168) );
  XOR U747 ( .A(g_input[52]), .B(state[52]), .Z(\w1[0][52] ) );
  XOR U748 ( .A(g_input[50]), .B(state[50]), .Z(\w1[0][50] ) );
  AND U749 ( .A(\SUBBYTES[0].a/w164 ), .B(\SUBBYTES[0].a/w160 ), .Z(
        \SUBBYTES[0].a/w201 ) );
  AND U750 ( .A(\SUBBYTES[0].a/w165 ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w199 ) );
  AND U751 ( .A(\SUBBYTES[0].a/w291 ), .B(n121), .Z(\SUBBYTES[0].a/w198 ) );
  XNOR U752 ( .A(\w1[0][121] ), .B(n170), .Z(n121) );
  XOR U753 ( .A(g_input[121]), .B(state[121]), .Z(\w1[0][121] ) );
  AND U754 ( .A(n171), .B(\SUBBYTES[0].a/w1816 ), .Z(\SUBBYTES[0].a/w1951 ) );
  AND U755 ( .A(n172), .B(\SUBBYTES[0].a/w1817 ), .Z(\SUBBYTES[0].a/w1949 ) );
  AND U756 ( .A(\SUBBYTES[0].a/w1947 ), .B(n173), .Z(\SUBBYTES[0].a/w1948 ) );
  ANDN U757 ( .A(\w1[0][56] ), .B(n174), .Z(\SUBBYTES[0].a/w1944 ) );
  AND U758 ( .A(n175), .B(\SUBBYTES[0].a/w1819 ), .Z(\SUBBYTES[0].a/w1942 ) );
  AND U759 ( .A(\SUBBYTES[0].a/w1940 ), .B(n176), .Z(\SUBBYTES[0].a/w1941 ) );
  XOR U760 ( .A(\SUBBYTES[0].a/w1884 ), .B(\SUBBYTES[0].a/n89 ), .Z(n176) );
  AND U761 ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w166 ), .Z(
        \SUBBYTES[0].a/w194 ) );
  XOR U762 ( .A(g_input[120]), .B(state[120]), .Z(\w1[0][120] ) );
  AND U763 ( .A(\SUBBYTES[0].a/w1927 ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/w1936 ) );
  AND U764 ( .A(\SUBBYTES[0].a/w1928 ), .B(\SUBBYTES[0].a/w1930 ), .Z(
        \SUBBYTES[0].a/w1934 ) );
  AND U765 ( .A(\SUBBYTES[0].a/w1931 ), .B(\SUBBYTES[0].a/w1932 ), .Z(
        \SUBBYTES[0].a/w1933 ) );
  AND U766 ( .A(\SUBBYTES[0].a/w167 ), .B(\SUBBYTES[0].a/w163 ), .Z(
        \SUBBYTES[0].a/w192 ) );
  AND U767 ( .A(\SUBBYTES[0].a/w1820 ), .B(n171), .Z(\SUBBYTES[0].a/w1919 ) );
  XOR U768 ( .A(\SUBBYTES[0].a/w1888 ), .B(n9), .Z(n171) );
  AND U769 ( .A(\SUBBYTES[0].a/w1821 ), .B(n172), .Z(\SUBBYTES[0].a/w1917 ) );
  XOR U770 ( .A(\SUBBYTES[0].a/n90 ), .B(\SUBBYTES[0].a/w1888 ), .Z(n172) );
  AND U771 ( .A(n177), .B(n173), .Z(\SUBBYTES[0].a/w1916 ) );
  XOR U772 ( .A(n9), .B(\SUBBYTES[0].a/n90 ), .Z(n173) );
  ANDN U773 ( .A(\SUBBYTES[0].a/w1822 ), .B(n174), .Z(\SUBBYTES[0].a/w1912 )
         );
  XNOR U774 ( .A(\SUBBYTES[0].a/w1881 ), .B(\SUBBYTES[0].a/w1884 ), .Z(n174)
         );
  AND U775 ( .A(\SUBBYTES[0].a/w1823 ), .B(n175), .Z(\SUBBYTES[0].a/w1910 ) );
  XNOR U776 ( .A(n178), .B(\SUBBYTES[0].a/w1881 ), .Z(n175) );
  AND U777 ( .A(\SUBBYTES[0].a/w252 ), .B(\SUBBYTES[0].a/w284 ), .Z(
        \SUBBYTES[0].a/w191 ) );
  AND U778 ( .A(\SUBBYTES[0].a/w1908 ), .B(n179), .Z(\SUBBYTES[0].a/w1909 ) );
  XOR U779 ( .A(n180), .B(n178), .Z(n179) );
  IV U780 ( .A(\SUBBYTES[0].a/n89 ), .Z(n178) );
  AND U781 ( .A(n181), .B(\SUBBYTES[0].a/w1927 ), .Z(\SUBBYTES[0].a/w1904 ) );
  ANDN U782 ( .A(\SUBBYTES[0].a/w1928 ), .B(n182), .Z(\SUBBYTES[0].a/w1902 )
         );
  AND U783 ( .A(n183), .B(\SUBBYTES[0].a/w1931 ), .Z(\SUBBYTES[0].a/w1901 ) );
  AND U784 ( .A(\SUBBYTES[0].a/w1887 ), .B(\SUBBYTES[0].a/w1886 ), .Z(
        \SUBBYTES[0].a/w1888 ) );
  IV U785 ( .A(n180), .Z(\SUBBYTES[0].a/w1884 ) );
  NAND U786 ( .A(\SUBBYTES[0].a/w1863 ), .B(\SUBBYTES[0].a/w1878 ), .Z(n180)
         );
  AND U787 ( .A(\SUBBYTES[0].a/w1880 ), .B(\SUBBYTES[0].a/w1886 ), .Z(
        \SUBBYTES[0].a/w1881 ) );
  AND U788 ( .A(\SUBBYTES[0].a/w1865 ), .B(\SUBBYTES[0].a/w1863 ), .Z(
        \SUBBYTES[0].a/w1875 ) );
  AND U789 ( .A(\SUBBYTES[0].a/w1866 ), .B(\SUBBYTES[0].a/w1864 ), .Z(
        \SUBBYTES[0].a/w1873 ) );
  AND U790 ( .A(\SUBBYTES[0].a/w1880 ), .B(\SUBBYTES[0].a/w1887 ), .Z(
        \SUBBYTES[0].a/w1872 ) );
  AND U791 ( .A(\SUBBYTES[0].a/w273 ), .B(n138), .Z(\SUBBYTES[0].a/w186 ) );
  XOR U792 ( .A(\w1[0][124] ), .B(\w1[0][127] ), .Z(n138) );
  AND U793 ( .A(\SUBBYTES[0].a/w1820 ), .B(\SUBBYTES[0].a/w1816 ), .Z(
        \SUBBYTES[0].a/w1857 ) );
  AND U794 ( .A(\SUBBYTES[0].a/w1821 ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1855 ) );
  AND U795 ( .A(\SUBBYTES[0].a/w1947 ), .B(n177), .Z(\SUBBYTES[0].a/w1854 ) );
  XNOR U796 ( .A(\w1[0][57] ), .B(n184), .Z(n177) );
  XOR U797 ( .A(g_input[57]), .B(state[57]), .Z(\w1[0][57] ) );
  AND U798 ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1822 ), .Z(
        \SUBBYTES[0].a/w1850 ) );
  XOR U799 ( .A(g_input[56]), .B(state[56]), .Z(\w1[0][56] ) );
  AND U800 ( .A(\SUBBYTES[0].a/w1823 ), .B(\SUBBYTES[0].a/w1819 ), .Z(
        \SUBBYTES[0].a/w1848 ) );
  AND U801 ( .A(\SUBBYTES[0].a/w1908 ), .B(\SUBBYTES[0].a/w1940 ), .Z(
        \SUBBYTES[0].a/w1847 ) );
  AND U802 ( .A(\SUBBYTES[0].a/w1929 ), .B(n181), .Z(\SUBBYTES[0].a/w1842 ) );
  XOR U803 ( .A(\w1[0][60] ), .B(\w1[0][63] ), .Z(n181) );
  ANDN U804 ( .A(\SUBBYTES[0].a/w1930 ), .B(n182), .Z(\SUBBYTES[0].a/w1840 )
         );
  XNOR U805 ( .A(\w1[0][58] ), .B(\w1[0][63] ), .Z(n182) );
  IV U806 ( .A(n184), .Z(\w1[0][63] ) );
  XNOR U807 ( .A(g_input[63]), .B(state[63]), .Z(n184) );
  ANDN U808 ( .A(\SUBBYTES[0].a/w274 ), .B(n140), .Z(\SUBBYTES[0].a/w184 ) );
  XNOR U809 ( .A(\w1[0][122] ), .B(\w1[0][127] ), .Z(n140) );
  IV U810 ( .A(n170), .Z(\w1[0][127] ) );
  XNOR U811 ( .A(g_input[127]), .B(state[127]), .Z(n170) );
  AND U812 ( .A(\SUBBYTES[0].a/w1932 ), .B(n183), .Z(\SUBBYTES[0].a/w1839 ) );
  XOR U813 ( .A(\w1[0][58] ), .B(\w1[0][60] ), .Z(n183) );
  XOR U814 ( .A(g_input[60]), .B(state[60]), .Z(\w1[0][60] ) );
  XOR U815 ( .A(g_input[58]), .B(state[58]), .Z(\w1[0][58] ) );
  AND U816 ( .A(\SUBBYTES[0].a/w276 ), .B(n141), .Z(\SUBBYTES[0].a/w183 ) );
  XOR U817 ( .A(\w1[0][122] ), .B(\w1[0][124] ), .Z(n141) );
  XOR U818 ( .A(g_input[124]), .B(state[124]), .Z(\w1[0][124] ) );
  XOR U819 ( .A(g_input[122]), .B(state[122]), .Z(\w1[0][122] ) );
  AND U820 ( .A(n185), .B(\SUBBYTES[0].a/w1609 ), .Z(\SUBBYTES[0].a/w1744 ) );
  AND U821 ( .A(n186), .B(\SUBBYTES[0].a/w1610 ), .Z(\SUBBYTES[0].a/w1742 ) );
  AND U822 ( .A(\SUBBYTES[0].a/w1740 ), .B(n187), .Z(\SUBBYTES[0].a/w1741 ) );
  ANDN U823 ( .A(\w1[0][64] ), .B(n188), .Z(\SUBBYTES[0].a/w1737 ) );
  AND U824 ( .A(n189), .B(\SUBBYTES[0].a/w1612 ), .Z(\SUBBYTES[0].a/w1735 ) );
  AND U825 ( .A(\SUBBYTES[0].a/w1733 ), .B(n190), .Z(\SUBBYTES[0].a/w1734 ) );
  XOR U826 ( .A(\SUBBYTES[0].a/w1677 ), .B(\SUBBYTES[0].a/n79 ), .Z(n190) );
  AND U827 ( .A(\SUBBYTES[0].a/w1720 ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/w1729 ) );
  AND U828 ( .A(\SUBBYTES[0].a/w1721 ), .B(\SUBBYTES[0].a/w1723 ), .Z(
        \SUBBYTES[0].a/w1727 ) );
  AND U829 ( .A(\SUBBYTES[0].a/w1724 ), .B(\SUBBYTES[0].a/w1725 ), .Z(
        \SUBBYTES[0].a/w1726 ) );
  AND U830 ( .A(\SUBBYTES[0].a/w1613 ), .B(n185), .Z(\SUBBYTES[0].a/w1712 ) );
  XOR U831 ( .A(\SUBBYTES[0].a/w1681 ), .B(n8), .Z(n185) );
  AND U832 ( .A(\SUBBYTES[0].a/w1614 ), .B(n186), .Z(\SUBBYTES[0].a/w1710 ) );
  XOR U833 ( .A(\SUBBYTES[0].a/n80 ), .B(\SUBBYTES[0].a/w1681 ), .Z(n186) );
  AND U834 ( .A(n191), .B(n187), .Z(\SUBBYTES[0].a/w1709 ) );
  XOR U835 ( .A(n8), .B(\SUBBYTES[0].a/n80 ), .Z(n187) );
  ANDN U836 ( .A(\SUBBYTES[0].a/w1615 ), .B(n188), .Z(\SUBBYTES[0].a/w1705 )
         );
  XNOR U837 ( .A(\SUBBYTES[0].a/w1674 ), .B(\SUBBYTES[0].a/w1677 ), .Z(n188)
         );
  AND U838 ( .A(\SUBBYTES[0].a/w1616 ), .B(n189), .Z(\SUBBYTES[0].a/w1703 ) );
  XNOR U839 ( .A(n192), .B(\SUBBYTES[0].a/w1674 ), .Z(n189) );
  AND U840 ( .A(\SUBBYTES[0].a/w1701 ), .B(n193), .Z(\SUBBYTES[0].a/w1702 ) );
  XOR U841 ( .A(n194), .B(n192), .Z(n193) );
  IV U842 ( .A(\SUBBYTES[0].a/n79 ), .Z(n192) );
  AND U843 ( .A(n195), .B(\SUBBYTES[0].a/w1720 ), .Z(\SUBBYTES[0].a/w1697 ) );
  ANDN U844 ( .A(\SUBBYTES[0].a/w1721 ), .B(n196), .Z(\SUBBYTES[0].a/w1695 )
         );
  AND U845 ( .A(n197), .B(\SUBBYTES[0].a/w1724 ), .Z(\SUBBYTES[0].a/w1694 ) );
  AND U846 ( .A(\SUBBYTES[0].a/w1680 ), .B(\SUBBYTES[0].a/w1679 ), .Z(
        \SUBBYTES[0].a/w1681 ) );
  IV U847 ( .A(n194), .Z(\SUBBYTES[0].a/w1677 ) );
  NAND U848 ( .A(\SUBBYTES[0].a/w1656 ), .B(\SUBBYTES[0].a/w1671 ), .Z(n194)
         );
  AND U849 ( .A(\SUBBYTES[0].a/w1673 ), .B(\SUBBYTES[0].a/w1679 ), .Z(
        \SUBBYTES[0].a/w1674 ) );
  AND U850 ( .A(\SUBBYTES[0].a/w1658 ), .B(\SUBBYTES[0].a/w1656 ), .Z(
        \SUBBYTES[0].a/w1668 ) );
  AND U851 ( .A(\SUBBYTES[0].a/w1659 ), .B(\SUBBYTES[0].a/w1657 ), .Z(
        \SUBBYTES[0].a/w1666 ) );
  AND U852 ( .A(\SUBBYTES[0].a/w1673 ), .B(\SUBBYTES[0].a/w1680 ), .Z(
        \SUBBYTES[0].a/w1665 ) );
  AND U853 ( .A(\SUBBYTES[0].a/w1613 ), .B(\SUBBYTES[0].a/w1609 ), .Z(
        \SUBBYTES[0].a/w1650 ) );
  AND U854 ( .A(\SUBBYTES[0].a/w1614 ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1648 ) );
  AND U855 ( .A(\SUBBYTES[0].a/w1740 ), .B(n191), .Z(\SUBBYTES[0].a/w1647 ) );
  XNOR U856 ( .A(\w1[0][65] ), .B(n198), .Z(n191) );
  XOR U857 ( .A(g_input[65]), .B(state[65]), .Z(\w1[0][65] ) );
  AND U858 ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1615 ), .Z(
        \SUBBYTES[0].a/w1643 ) );
  XOR U859 ( .A(g_input[64]), .B(state[64]), .Z(\w1[0][64] ) );
  AND U860 ( .A(\SUBBYTES[0].a/w1616 ), .B(\SUBBYTES[0].a/w1612 ), .Z(
        \SUBBYTES[0].a/w1641 ) );
  AND U861 ( .A(\SUBBYTES[0].a/w1701 ), .B(\SUBBYTES[0].a/w1733 ), .Z(
        \SUBBYTES[0].a/w1640 ) );
  AND U862 ( .A(\SUBBYTES[0].a/w1722 ), .B(n195), .Z(\SUBBYTES[0].a/w1635 ) );
  XOR U863 ( .A(\w1[0][68] ), .B(\w1[0][71] ), .Z(n195) );
  ANDN U864 ( .A(\SUBBYTES[0].a/w1723 ), .B(n196), .Z(\SUBBYTES[0].a/w1633 )
         );
  XNOR U865 ( .A(\w1[0][66] ), .B(\w1[0][71] ), .Z(n196) );
  IV U866 ( .A(n198), .Z(\w1[0][71] ) );
  XNOR U867 ( .A(g_input[71]), .B(state[71]), .Z(n198) );
  AND U868 ( .A(\SUBBYTES[0].a/w1725 ), .B(n197), .Z(\SUBBYTES[0].a/w1632 ) );
  XOR U869 ( .A(\w1[0][66] ), .B(\w1[0][68] ), .Z(n197) );
  XOR U870 ( .A(g_input[68]), .B(state[68]), .Z(\w1[0][68] ) );
  XOR U871 ( .A(g_input[66]), .B(state[66]), .Z(\w1[0][66] ) );
  AND U872 ( .A(n199), .B(\SUBBYTES[0].a/w1402 ), .Z(\SUBBYTES[0].a/w1537 ) );
  AND U873 ( .A(n200), .B(\SUBBYTES[0].a/w1403 ), .Z(\SUBBYTES[0].a/w1535 ) );
  AND U874 ( .A(\SUBBYTES[0].a/w1533 ), .B(n201), .Z(\SUBBYTES[0].a/w1534 ) );
  ANDN U875 ( .A(\w1[0][72] ), .B(n202), .Z(\SUBBYTES[0].a/w1530 ) );
  AND U876 ( .A(n203), .B(\SUBBYTES[0].a/w1405 ), .Z(\SUBBYTES[0].a/w1528 ) );
  AND U877 ( .A(\SUBBYTES[0].a/w1526 ), .B(n204), .Z(\SUBBYTES[0].a/w1527 ) );
  XOR U878 ( .A(\SUBBYTES[0].a/w1470 ), .B(\SUBBYTES[0].a/n69 ), .Z(n204) );
  AND U879 ( .A(\SUBBYTES[0].a/w1513 ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/w1522 ) );
  AND U880 ( .A(\SUBBYTES[0].a/w1514 ), .B(\SUBBYTES[0].a/w1516 ), .Z(
        \SUBBYTES[0].a/w1520 ) );
  AND U881 ( .A(\SUBBYTES[0].a/w1517 ), .B(\SUBBYTES[0].a/w1518 ), .Z(
        \SUBBYTES[0].a/w1519 ) );
  AND U882 ( .A(\SUBBYTES[0].a/w1406 ), .B(n199), .Z(\SUBBYTES[0].a/w1505 ) );
  XOR U883 ( .A(\SUBBYTES[0].a/w1474 ), .B(n7), .Z(n199) );
  AND U884 ( .A(\SUBBYTES[0].a/w1407 ), .B(n200), .Z(\SUBBYTES[0].a/w1503 ) );
  XOR U885 ( .A(\SUBBYTES[0].a/n70 ), .B(\SUBBYTES[0].a/w1474 ), .Z(n200) );
  AND U886 ( .A(n205), .B(n201), .Z(\SUBBYTES[0].a/w1502 ) );
  XOR U887 ( .A(n7), .B(\SUBBYTES[0].a/n70 ), .Z(n201) );
  ANDN U888 ( .A(\SUBBYTES[0].a/w1408 ), .B(n202), .Z(\SUBBYTES[0].a/w1498 )
         );
  XNOR U889 ( .A(\SUBBYTES[0].a/w1467 ), .B(\SUBBYTES[0].a/w1470 ), .Z(n202)
         );
  AND U890 ( .A(\SUBBYTES[0].a/w1409 ), .B(n203), .Z(\SUBBYTES[0].a/w1496 ) );
  XNOR U891 ( .A(n206), .B(\SUBBYTES[0].a/w1467 ), .Z(n203) );
  AND U892 ( .A(\SUBBYTES[0].a/w1494 ), .B(n207), .Z(\SUBBYTES[0].a/w1495 ) );
  XOR U893 ( .A(n208), .B(n206), .Z(n207) );
  IV U894 ( .A(\SUBBYTES[0].a/n69 ), .Z(n206) );
  AND U895 ( .A(n209), .B(\SUBBYTES[0].a/w1513 ), .Z(\SUBBYTES[0].a/w1490 ) );
  ANDN U896 ( .A(\SUBBYTES[0].a/w1514 ), .B(n210), .Z(\SUBBYTES[0].a/w1488 )
         );
  AND U897 ( .A(n211), .B(\SUBBYTES[0].a/w1517 ), .Z(\SUBBYTES[0].a/w1487 ) );
  AND U898 ( .A(\SUBBYTES[0].a/w1473 ), .B(\SUBBYTES[0].a/w1472 ), .Z(
        \SUBBYTES[0].a/w1474 ) );
  IV U899 ( .A(n208), .Z(\SUBBYTES[0].a/w1470 ) );
  NAND U900 ( .A(\SUBBYTES[0].a/w1449 ), .B(\SUBBYTES[0].a/w1464 ), .Z(n208)
         );
  AND U901 ( .A(\SUBBYTES[0].a/w1466 ), .B(\SUBBYTES[0].a/w1472 ), .Z(
        \SUBBYTES[0].a/w1467 ) );
  AND U902 ( .A(\SUBBYTES[0].a/w1451 ), .B(\SUBBYTES[0].a/w1449 ), .Z(
        \SUBBYTES[0].a/w1461 ) );
  AND U903 ( .A(\SUBBYTES[0].a/w1452 ), .B(\SUBBYTES[0].a/w1450 ), .Z(
        \SUBBYTES[0].a/w1459 ) );
  AND U904 ( .A(\SUBBYTES[0].a/w1466 ), .B(\SUBBYTES[0].a/w1473 ), .Z(
        \SUBBYTES[0].a/w1458 ) );
  AND U905 ( .A(\SUBBYTES[0].a/w1406 ), .B(\SUBBYTES[0].a/w1402 ), .Z(
        \SUBBYTES[0].a/w1443 ) );
  AND U906 ( .A(\SUBBYTES[0].a/w1407 ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1441 ) );
  AND U907 ( .A(\SUBBYTES[0].a/w1533 ), .B(n205), .Z(\SUBBYTES[0].a/w1440 ) );
  XNOR U908 ( .A(\w1[0][73] ), .B(n212), .Z(n205) );
  XOR U909 ( .A(g_input[73]), .B(state[73]), .Z(\w1[0][73] ) );
  AND U910 ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1408 ), .Z(
        \SUBBYTES[0].a/w1436 ) );
  XOR U911 ( .A(g_input[72]), .B(state[72]), .Z(\w1[0][72] ) );
  AND U912 ( .A(\SUBBYTES[0].a/w1409 ), .B(\SUBBYTES[0].a/w1405 ), .Z(
        \SUBBYTES[0].a/w1434 ) );
  AND U913 ( .A(\SUBBYTES[0].a/w1494 ), .B(\SUBBYTES[0].a/w1526 ), .Z(
        \SUBBYTES[0].a/w1433 ) );
  AND U914 ( .A(\SUBBYTES[0].a/w1515 ), .B(n209), .Z(\SUBBYTES[0].a/w1428 ) );
  XOR U915 ( .A(\w1[0][76] ), .B(\w1[0][79] ), .Z(n209) );
  ANDN U916 ( .A(\SUBBYTES[0].a/w1516 ), .B(n210), .Z(\SUBBYTES[0].a/w1426 )
         );
  XNOR U917 ( .A(\w1[0][74] ), .B(\w1[0][79] ), .Z(n210) );
  IV U918 ( .A(n212), .Z(\w1[0][79] ) );
  XNOR U919 ( .A(g_input[79]), .B(state[79]), .Z(n212) );
  AND U920 ( .A(\SUBBYTES[0].a/w1518 ), .B(n211), .Z(\SUBBYTES[0].a/w1425 ) );
  XOR U921 ( .A(\w1[0][74] ), .B(\w1[0][76] ), .Z(n211) );
  XOR U922 ( .A(g_input[76]), .B(state[76]), .Z(\w1[0][76] ) );
  XOR U923 ( .A(g_input[74]), .B(state[74]), .Z(\w1[0][74] ) );
  AND U924 ( .A(n213), .B(\SUBBYTES[0].a/w1195 ), .Z(\SUBBYTES[0].a/w1330 ) );
  AND U925 ( .A(n214), .B(\SUBBYTES[0].a/w1196 ), .Z(\SUBBYTES[0].a/w1328 ) );
  AND U926 ( .A(\SUBBYTES[0].a/w1326 ), .B(n215), .Z(\SUBBYTES[0].a/w1327 ) );
  ANDN U927 ( .A(\w1[0][80] ), .B(n216), .Z(\SUBBYTES[0].a/w1323 ) );
  AND U928 ( .A(n217), .B(\SUBBYTES[0].a/w1198 ), .Z(\SUBBYTES[0].a/w1321 ) );
  AND U929 ( .A(\SUBBYTES[0].a/w1319 ), .B(n218), .Z(\SUBBYTES[0].a/w1320 ) );
  XOR U930 ( .A(\SUBBYTES[0].a/w1263 ), .B(\SUBBYTES[0].a/n59 ), .Z(n218) );
  AND U931 ( .A(\SUBBYTES[0].a/w1306 ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/w1315 ) );
  AND U932 ( .A(\SUBBYTES[0].a/w1307 ), .B(\SUBBYTES[0].a/w1309 ), .Z(
        \SUBBYTES[0].a/w1313 ) );
  AND U933 ( .A(\SUBBYTES[0].a/w1310 ), .B(\SUBBYTES[0].a/w1311 ), .Z(
        \SUBBYTES[0].a/w1312 ) );
  AND U934 ( .A(\SUBBYTES[0].a/w1199 ), .B(n213), .Z(\SUBBYTES[0].a/w1298 ) );
  XOR U935 ( .A(\SUBBYTES[0].a/w1267 ), .B(n6), .Z(n213) );
  AND U936 ( .A(\SUBBYTES[0].a/w1200 ), .B(n214), .Z(\SUBBYTES[0].a/w1296 ) );
  XOR U937 ( .A(\SUBBYTES[0].a/n60 ), .B(\SUBBYTES[0].a/w1267 ), .Z(n214) );
  AND U938 ( .A(n219), .B(n215), .Z(\SUBBYTES[0].a/w1295 ) );
  XOR U939 ( .A(n6), .B(\SUBBYTES[0].a/n60 ), .Z(n215) );
  ANDN U940 ( .A(\SUBBYTES[0].a/w1201 ), .B(n216), .Z(\SUBBYTES[0].a/w1291 )
         );
  XNOR U941 ( .A(\SUBBYTES[0].a/w1260 ), .B(\SUBBYTES[0].a/w1263 ), .Z(n216)
         );
  AND U942 ( .A(\SUBBYTES[0].a/w1202 ), .B(n217), .Z(\SUBBYTES[0].a/w1289 ) );
  XNOR U943 ( .A(n220), .B(\SUBBYTES[0].a/w1260 ), .Z(n217) );
  AND U944 ( .A(\SUBBYTES[0].a/w1287 ), .B(n221), .Z(\SUBBYTES[0].a/w1288 ) );
  XOR U945 ( .A(n222), .B(n220), .Z(n221) );
  IV U946 ( .A(\SUBBYTES[0].a/n59 ), .Z(n220) );
  AND U947 ( .A(n223), .B(\SUBBYTES[0].a/w1306 ), .Z(\SUBBYTES[0].a/w1283 ) );
  ANDN U948 ( .A(\SUBBYTES[0].a/w1307 ), .B(n224), .Z(\SUBBYTES[0].a/w1281 )
         );
  AND U949 ( .A(n225), .B(\SUBBYTES[0].a/w1310 ), .Z(\SUBBYTES[0].a/w1280 ) );
  AND U950 ( .A(\SUBBYTES[0].a/w1266 ), .B(\SUBBYTES[0].a/w1265 ), .Z(
        \SUBBYTES[0].a/w1267 ) );
  IV U951 ( .A(n222), .Z(\SUBBYTES[0].a/w1263 ) );
  NAND U952 ( .A(\SUBBYTES[0].a/w1242 ), .B(\SUBBYTES[0].a/w1257 ), .Z(n222)
         );
  AND U953 ( .A(\SUBBYTES[0].a/w1259 ), .B(\SUBBYTES[0].a/w1265 ), .Z(
        \SUBBYTES[0].a/w1260 ) );
  AND U954 ( .A(\SUBBYTES[0].a/w1244 ), .B(\SUBBYTES[0].a/w1242 ), .Z(
        \SUBBYTES[0].a/w1254 ) );
  AND U955 ( .A(\SUBBYTES[0].a/w1245 ), .B(\SUBBYTES[0].a/w1243 ), .Z(
        \SUBBYTES[0].a/w1252 ) );
  AND U956 ( .A(\SUBBYTES[0].a/w1259 ), .B(\SUBBYTES[0].a/w1266 ), .Z(
        \SUBBYTES[0].a/w1251 ) );
  AND U957 ( .A(\SUBBYTES[0].a/w1199 ), .B(\SUBBYTES[0].a/w1195 ), .Z(
        \SUBBYTES[0].a/w1236 ) );
  AND U958 ( .A(\SUBBYTES[0].a/w1200 ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1234 ) );
  AND U959 ( .A(\SUBBYTES[0].a/w1326 ), .B(n219), .Z(\SUBBYTES[0].a/w1233 ) );
  XNOR U960 ( .A(\w1[0][81] ), .B(n226), .Z(n219) );
  XOR U961 ( .A(g_input[81]), .B(state[81]), .Z(\w1[0][81] ) );
  AND U962 ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1201 ), .Z(
        \SUBBYTES[0].a/w1229 ) );
  XOR U963 ( .A(g_input[80]), .B(state[80]), .Z(\w1[0][80] ) );
  AND U964 ( .A(\SUBBYTES[0].a/w1202 ), .B(\SUBBYTES[0].a/w1198 ), .Z(
        \SUBBYTES[0].a/w1227 ) );
  AND U965 ( .A(\SUBBYTES[0].a/w1287 ), .B(\SUBBYTES[0].a/w1319 ), .Z(
        \SUBBYTES[0].a/w1226 ) );
  AND U966 ( .A(\SUBBYTES[0].a/w1308 ), .B(n223), .Z(\SUBBYTES[0].a/w1221 ) );
  XOR U967 ( .A(\w1[0][84] ), .B(\w1[0][87] ), .Z(n223) );
  ANDN U968 ( .A(\SUBBYTES[0].a/w1309 ), .B(n224), .Z(\SUBBYTES[0].a/w1219 )
         );
  XNOR U969 ( .A(\w1[0][82] ), .B(\w1[0][87] ), .Z(n224) );
  IV U970 ( .A(n226), .Z(\w1[0][87] ) );
  XNOR U971 ( .A(g_input[87]), .B(state[87]), .Z(n226) );
  AND U972 ( .A(\SUBBYTES[0].a/w1311 ), .B(n225), .Z(\SUBBYTES[0].a/w1218 ) );
  XOR U973 ( .A(\w1[0][82] ), .B(\w1[0][84] ), .Z(n225) );
  XOR U974 ( .A(g_input[84]), .B(state[84]), .Z(\w1[0][84] ) );
  XOR U975 ( .A(g_input[82]), .B(state[82]), .Z(\w1[0][82] ) );
  AND U976 ( .A(n227), .B(\SUBBYTES[0].a/w988 ), .Z(\SUBBYTES[0].a/w1123 ) );
  AND U977 ( .A(n228), .B(\SUBBYTES[0].a/w989 ), .Z(\SUBBYTES[0].a/w1121 ) );
  AND U978 ( .A(\SUBBYTES[0].a/w1119 ), .B(n229), .Z(\SUBBYTES[0].a/w1120 ) );
  ANDN U979 ( .A(\w1[0][88] ), .B(n230), .Z(\SUBBYTES[0].a/w1116 ) );
  AND U980 ( .A(n231), .B(\SUBBYTES[0].a/w991 ), .Z(\SUBBYTES[0].a/w1114 ) );
  AND U981 ( .A(\SUBBYTES[0].a/w1112 ), .B(n232), .Z(\SUBBYTES[0].a/w1113 ) );
  XOR U982 ( .A(\SUBBYTES[0].a/w1056 ), .B(\SUBBYTES[0].a/n49 ), .Z(n232) );
  AND U983 ( .A(\SUBBYTES[0].a/w1099 ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/w1108 ) );
  AND U984 ( .A(\SUBBYTES[0].a/w1100 ), .B(\SUBBYTES[0].a/w1102 ), .Z(
        \SUBBYTES[0].a/w1106 ) );
  AND U985 ( .A(\SUBBYTES[0].a/w1103 ), .B(\SUBBYTES[0].a/w1104 ), .Z(
        \SUBBYTES[0].a/w1105 ) );
  AND U986 ( .A(\SUBBYTES[0].a/w992 ), .B(n227), .Z(\SUBBYTES[0].a/w1091 ) );
  XOR U987 ( .A(\SUBBYTES[0].a/w1060 ), .B(n5), .Z(n227) );
  AND U988 ( .A(\SUBBYTES[0].a/w993 ), .B(n228), .Z(\SUBBYTES[0].a/w1089 ) );
  XOR U989 ( .A(\SUBBYTES[0].a/n50 ), .B(\SUBBYTES[0].a/w1060 ), .Z(n228) );
  AND U990 ( .A(n233), .B(n229), .Z(\SUBBYTES[0].a/w1088 ) );
  XOR U991 ( .A(n5), .B(\SUBBYTES[0].a/n50 ), .Z(n229) );
  ANDN U992 ( .A(\SUBBYTES[0].a/w994 ), .B(n230), .Z(\SUBBYTES[0].a/w1084 ) );
  XNOR U993 ( .A(\SUBBYTES[0].a/w1053 ), .B(\SUBBYTES[0].a/w1056 ), .Z(n230)
         );
  AND U994 ( .A(\SUBBYTES[0].a/w995 ), .B(n231), .Z(\SUBBYTES[0].a/w1082 ) );
  XNOR U995 ( .A(n234), .B(\SUBBYTES[0].a/w1053 ), .Z(n231) );
  AND U996 ( .A(\SUBBYTES[0].a/w1080 ), .B(n235), .Z(\SUBBYTES[0].a/w1081 ) );
  XOR U997 ( .A(n236), .B(n234), .Z(n235) );
  IV U998 ( .A(\SUBBYTES[0].a/n49 ), .Z(n234) );
  AND U999 ( .A(n237), .B(\SUBBYTES[0].a/w1099 ), .Z(\SUBBYTES[0].a/w1076 ) );
  ANDN U1000 ( .A(\SUBBYTES[0].a/w1100 ), .B(n238), .Z(\SUBBYTES[0].a/w1074 )
         );
  AND U1001 ( .A(n239), .B(\SUBBYTES[0].a/w1103 ), .Z(\SUBBYTES[0].a/w1073 )
         );
  AND U1002 ( .A(\SUBBYTES[0].a/w1059 ), .B(\SUBBYTES[0].a/w1058 ), .Z(
        \SUBBYTES[0].a/w1060 ) );
  IV U1003 ( .A(n236), .Z(\SUBBYTES[0].a/w1056 ) );
  NAND U1004 ( .A(\SUBBYTES[0].a/w1035 ), .B(\SUBBYTES[0].a/w1050 ), .Z(n236)
         );
  AND U1005 ( .A(\SUBBYTES[0].a/w1052 ), .B(\SUBBYTES[0].a/w1058 ), .Z(
        \SUBBYTES[0].a/w1053 ) );
  AND U1006 ( .A(\SUBBYTES[0].a/w1037 ), .B(\SUBBYTES[0].a/w1035 ), .Z(
        \SUBBYTES[0].a/w1047 ) );
  AND U1007 ( .A(\SUBBYTES[0].a/w1038 ), .B(\SUBBYTES[0].a/w1036 ), .Z(
        \SUBBYTES[0].a/w1045 ) );
  AND U1008 ( .A(\SUBBYTES[0].a/w1052 ), .B(\SUBBYTES[0].a/w1059 ), .Z(
        \SUBBYTES[0].a/w1044 ) );
  AND U1009 ( .A(\SUBBYTES[0].a/w992 ), .B(\SUBBYTES[0].a/w988 ), .Z(
        \SUBBYTES[0].a/w1029 ) );
  AND U1010 ( .A(\SUBBYTES[0].a/w993 ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w1027 ) );
  AND U1011 ( .A(\SUBBYTES[0].a/w1119 ), .B(n233), .Z(\SUBBYTES[0].a/w1026 )
         );
  XNOR U1012 ( .A(\w1[0][89] ), .B(n240), .Z(n233) );
  XOR U1013 ( .A(g_input[89]), .B(state[89]), .Z(\w1[0][89] ) );
  AND U1014 ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w994 ), .Z(
        \SUBBYTES[0].a/w1022 ) );
  XOR U1015 ( .A(g_input[88]), .B(state[88]), .Z(\w1[0][88] ) );
  AND U1016 ( .A(\SUBBYTES[0].a/w995 ), .B(\SUBBYTES[0].a/w991 ), .Z(
        \SUBBYTES[0].a/w1020 ) );
  AND U1017 ( .A(\SUBBYTES[0].a/w1080 ), .B(\SUBBYTES[0].a/w1112 ), .Z(
        \SUBBYTES[0].a/w1019 ) );
  AND U1018 ( .A(\SUBBYTES[0].a/w1101 ), .B(n237), .Z(\SUBBYTES[0].a/w1014 )
         );
  XOR U1019 ( .A(\w1[0][92] ), .B(\w1[0][95] ), .Z(n237) );
  ANDN U1020 ( .A(\SUBBYTES[0].a/w1102 ), .B(n238), .Z(\SUBBYTES[0].a/w1012 )
         );
  XNOR U1021 ( .A(\w1[0][90] ), .B(\w1[0][95] ), .Z(n238) );
  IV U1022 ( .A(n240), .Z(\w1[0][95] ) );
  XNOR U1023 ( .A(g_input[95]), .B(state[95]), .Z(n240) );
  AND U1024 ( .A(\SUBBYTES[0].a/w1104 ), .B(n239), .Z(\SUBBYTES[0].a/w1011 )
         );
  XOR U1025 ( .A(\w1[0][90] ), .B(\w1[0][92] ), .Z(n239) );
  XOR U1026 ( .A(g_input[92]), .B(state[92]), .Z(\w1[0][92] ) );
  XOR U1027 ( .A(g_input[90]), .B(state[90]), .Z(\w1[0][90] ) );
  AND U1028 ( .A(\SUBBYTES[0].a/w2084 ), .B(\SUBBYTES[0].a/w2071 ), .Z(
        \SUBBYTES[0].a/n99 ) );
  AND U1029 ( .A(\SUBBYTES[0].a/w1877 ), .B(\SUBBYTES[0].a/w1866 ), .Z(
        \SUBBYTES[0].a/n90 ) );
  AND U1030 ( .A(\SUBBYTES[0].a/w221 ), .B(\SUBBYTES[0].a/w208 ), .Z(
        \SUBBYTES[0].a/n9 ) );
  AND U1031 ( .A(\SUBBYTES[0].a/w1877 ), .B(\SUBBYTES[0].a/w1864 ), .Z(
        \SUBBYTES[0].a/n89 ) );
  AND U1032 ( .A(\SUBBYTES[0].a/w1670 ), .B(\SUBBYTES[0].a/w1659 ), .Z(
        \SUBBYTES[0].a/n80 ) );
  AND U1033 ( .A(\SUBBYTES[0].a/w1670 ), .B(\SUBBYTES[0].a/w1657 ), .Z(
        \SUBBYTES[0].a/n79 ) );
  AND U1034 ( .A(\SUBBYTES[0].a/w1463 ), .B(\SUBBYTES[0].a/w1452 ), .Z(
        \SUBBYTES[0].a/n70 ) );
  AND U1035 ( .A(\SUBBYTES[0].a/w1463 ), .B(\SUBBYTES[0].a/w1450 ), .Z(
        \SUBBYTES[0].a/n69 ) );
  AND U1036 ( .A(\SUBBYTES[0].a/w1256 ), .B(\SUBBYTES[0].a/w1245 ), .Z(
        \SUBBYTES[0].a/n60 ) );
  AND U1037 ( .A(\SUBBYTES[0].a/w1256 ), .B(\SUBBYTES[0].a/w1243 ), .Z(
        \SUBBYTES[0].a/n59 ) );
  AND U1038 ( .A(\SUBBYTES[0].a/w1049 ), .B(\SUBBYTES[0].a/w1038 ), .Z(
        \SUBBYTES[0].a/n50 ) );
  AND U1039 ( .A(\SUBBYTES[0].a/w1049 ), .B(\SUBBYTES[0].a/w1036 ), .Z(
        \SUBBYTES[0].a/n49 ) );
  AND U1040 ( .A(\SUBBYTES[0].a/w842 ), .B(\SUBBYTES[0].a/w831 ), .Z(
        \SUBBYTES[0].a/n40 ) );
  AND U1041 ( .A(\SUBBYTES[0].a/w842 ), .B(\SUBBYTES[0].a/w829 ), .Z(
        \SUBBYTES[0].a/n39 ) );
  AND U1042 ( .A(\SUBBYTES[0].a/w635 ), .B(\SUBBYTES[0].a/w624 ), .Z(
        \SUBBYTES[0].a/n30 ) );
  AND U1043 ( .A(\SUBBYTES[0].a/w635 ), .B(\SUBBYTES[0].a/w622 ), .Z(
        \SUBBYTES[0].a/n29 ) );
  AND U1044 ( .A(\SUBBYTES[0].a/w428 ), .B(\SUBBYTES[0].a/w417 ), .Z(
        \SUBBYTES[0].a/n20 ) );
  AND U1045 ( .A(\SUBBYTES[0].a/w428 ), .B(\SUBBYTES[0].a/w415 ), .Z(
        \SUBBYTES[0].a/n19 ) );
  AND U1046 ( .A(\SUBBYTES[0].a/w3326 ), .B(\SUBBYTES[0].a/w3315 ), .Z(
        \SUBBYTES[0].a/n160 ) );
  AND U1047 ( .A(\SUBBYTES[0].a/w3326 ), .B(\SUBBYTES[0].a/w3313 ), .Z(
        \SUBBYTES[0].a/n159 ) );
  AND U1048 ( .A(\SUBBYTES[0].a/w3119 ), .B(\SUBBYTES[0].a/w3108 ), .Z(
        \SUBBYTES[0].a/n150 ) );
  AND U1049 ( .A(\SUBBYTES[0].a/w3119 ), .B(\SUBBYTES[0].a/w3106 ), .Z(
        \SUBBYTES[0].a/n149 ) );
  AND U1050 ( .A(\SUBBYTES[0].a/w2912 ), .B(\SUBBYTES[0].a/w2901 ), .Z(
        \SUBBYTES[0].a/n140 ) );
  AND U1051 ( .A(\SUBBYTES[0].a/w2912 ), .B(\SUBBYTES[0].a/w2899 ), .Z(
        \SUBBYTES[0].a/n139 ) );
  AND U1052 ( .A(\SUBBYTES[0].a/w2705 ), .B(\SUBBYTES[0].a/w2694 ), .Z(
        \SUBBYTES[0].a/n130 ) );
  AND U1053 ( .A(\SUBBYTES[0].a/w2705 ), .B(\SUBBYTES[0].a/w2692 ), .Z(
        \SUBBYTES[0].a/n129 ) );
  AND U1054 ( .A(\SUBBYTES[0].a/w2498 ), .B(\SUBBYTES[0].a/w2487 ), .Z(
        \SUBBYTES[0].a/n120 ) );
  AND U1055 ( .A(\SUBBYTES[0].a/w2498 ), .B(\SUBBYTES[0].a/w2485 ), .Z(
        \SUBBYTES[0].a/n119 ) );
  AND U1056 ( .A(\SUBBYTES[0].a/w2291 ), .B(\SUBBYTES[0].a/w2280 ), .Z(
        \SUBBYTES[0].a/n110 ) );
  AND U1057 ( .A(\SUBBYTES[0].a/w2291 ), .B(\SUBBYTES[0].a/w2278 ), .Z(
        \SUBBYTES[0].a/n109 ) );
  AND U1058 ( .A(\SUBBYTES[0].a/w2084 ), .B(\SUBBYTES[0].a/w2073 ), .Z(
        \SUBBYTES[0].a/n100 ) );
  AND U1059 ( .A(\SUBBYTES[0].a/w221 ), .B(\SUBBYTES[0].a/w210 ), .Z(
        \SUBBYTES[0].a/n10 ) );
endmodule

