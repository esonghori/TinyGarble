
module mult_N8_CC4 ( clk, rst, a, b, c );
  input [7:0] a;
  input [1:0] b;
  output [15:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94;
  wire   [15:0] sreg;

  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(sreg[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(sreg[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(sreg[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(sreg[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(sreg[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(sreg[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(sreg[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(sreg[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U5 ( .A(n72), .B(n70), .Z(n1) );
  XOR U6 ( .A(n72), .B(n70), .Z(n2) );
  NANDN U7 ( .A(n71), .B(n2), .Z(n3) );
  NAND U8 ( .A(n1), .B(n3), .Z(n79) );
  NAND U9 ( .A(n79), .B(n77), .Z(n4) );
  XOR U10 ( .A(n79), .B(n77), .Z(n5) );
  NANDN U11 ( .A(n78), .B(n5), .Z(n6) );
  NAND U12 ( .A(n4), .B(n6), .Z(n87) );
  NAND U13 ( .A(n65), .B(n63), .Z(n7) );
  XOR U14 ( .A(n65), .B(n63), .Z(n8) );
  NANDN U15 ( .A(n64), .B(n8), .Z(n9) );
  NAND U16 ( .A(n7), .B(n9), .Z(n72) );
  NAND U17 ( .A(n61), .B(n60), .Z(n10) );
  XOR U18 ( .A(n61), .B(n60), .Z(n11) );
  NANDN U19 ( .A(sreg[9]), .B(n11), .Z(n12) );
  NAND U20 ( .A(n10), .B(n12), .Z(n68) );
  NAND U21 ( .A(n81), .B(n80), .Z(n13) );
  XOR U22 ( .A(n81), .B(n80), .Z(n14) );
  NANDN U23 ( .A(sreg[12]), .B(n14), .Z(n15) );
  NAND U24 ( .A(n13), .B(n15), .Z(n84) );
  NAND U25 ( .A(n68), .B(n67), .Z(n16) );
  XOR U26 ( .A(n68), .B(n67), .Z(n17) );
  NANDN U27 ( .A(sreg[10]), .B(n17), .Z(n18) );
  NAND U28 ( .A(n16), .B(n18), .Z(n75) );
  NAND U29 ( .A(n84), .B(n83), .Z(n19) );
  XOR U30 ( .A(n84), .B(n83), .Z(n20) );
  NANDN U31 ( .A(sreg[13]), .B(n20), .Z(n21) );
  NAND U32 ( .A(n19), .B(n21), .Z(n93) );
  OR U33 ( .A(n56), .B(n58), .Z(n22) );
  NANDN U34 ( .A(n57), .B(n22), .Z(n23) );
  NANDN U35 ( .A(n58), .B(n57), .Z(n24) );
  NAND U36 ( .A(n55), .B(n24), .Z(n25) );
  NAND U37 ( .A(n23), .B(n25), .Z(n65) );
  NAND U38 ( .A(n75), .B(n74), .Z(n26) );
  XOR U39 ( .A(n75), .B(n74), .Z(n27) );
  NANDN U40 ( .A(sreg[11]), .B(n27), .Z(n28) );
  NAND U41 ( .A(n26), .B(n28), .Z(n81) );
  XOR U42 ( .A(n94), .B(n93), .Z(n29) );
  NANDN U43 ( .A(n92), .B(n29), .Z(n30) );
  NAND U44 ( .A(n93), .B(n94), .Z(n31) );
  AND U45 ( .A(n30), .B(n31), .Z(c[15]) );
  AND U46 ( .A(b[0]), .B(a[0]), .Z(n32) );
  XOR U47 ( .A(n32), .B(sreg[6]), .Z(c[6]) );
  AND U48 ( .A(b[0]), .B(a[1]), .Z(n56) );
  NAND U49 ( .A(b[1]), .B(a[0]), .Z(n44) );
  XOR U50 ( .A(n56), .B(n44), .Z(n39) );
  AND U51 ( .A(n32), .B(sreg[6]), .Z(n38) );
  IV U52 ( .A(n38), .Z(n37) );
  XNOR U53 ( .A(sreg[7]), .B(n37), .Z(n33) );
  XNOR U54 ( .A(n39), .B(n33), .Z(c[7]) );
  ANDN U55 ( .B(n56), .A(n44), .Z(n58) );
  AND U56 ( .A(a[2]), .B(b[0]), .Z(n35) );
  NAND U57 ( .A(a[1]), .B(b[1]), .Z(n34) );
  XNOR U58 ( .A(n35), .B(n34), .Z(n36) );
  XNOR U59 ( .A(n58), .B(n36), .Z(n50) );
  IV U60 ( .A(n50), .Z(n48) );
  NANDN U61 ( .A(sreg[7]), .B(n37), .Z(n42) );
  AND U62 ( .A(sreg[7]), .B(n38), .Z(n40) );
  NANDN U63 ( .A(n40), .B(n39), .Z(n41) );
  AND U64 ( .A(n42), .B(n41), .Z(n49) );
  XNOR U65 ( .A(n48), .B(n49), .Z(n43) );
  XNOR U66 ( .A(sreg[8]), .B(n43), .Z(c[8]) );
  AND U67 ( .A(b[0]), .B(a[3]), .Z(n55) );
  NAND U68 ( .A(b[1]), .B(a[2]), .Z(n57) );
  XNOR U69 ( .A(n56), .B(n57), .Z(n46) );
  NAND U70 ( .A(n56), .B(n44), .Z(n45) );
  NAND U71 ( .A(n46), .B(n45), .Z(n47) );
  XOR U72 ( .A(n55), .B(n47), .Z(n60) );
  NAND U73 ( .A(n48), .B(n49), .Z(n53) );
  ANDN U74 ( .B(n50), .A(n49), .Z(n51) );
  NANDN U75 ( .A(n51), .B(sreg[8]), .Z(n52) );
  AND U76 ( .A(n53), .B(n52), .Z(n61) );
  XNOR U77 ( .A(n61), .B(sreg[9]), .Z(n54) );
  XNOR U78 ( .A(n60), .B(n54), .Z(c[9]) );
  NAND U79 ( .A(b[0]), .B(a[4]), .Z(n64) );
  AND U80 ( .A(b[1]), .B(a[3]), .Z(n63) );
  XNOR U81 ( .A(n65), .B(n63), .Z(n59) );
  XNOR U82 ( .A(n64), .B(n59), .Z(n67) );
  XNOR U83 ( .A(n68), .B(sreg[10]), .Z(n62) );
  XNOR U84 ( .A(n67), .B(n62), .Z(c[10]) );
  NAND U85 ( .A(b[0]), .B(a[5]), .Z(n71) );
  AND U86 ( .A(b[1]), .B(a[4]), .Z(n70) );
  XNOR U87 ( .A(n72), .B(n70), .Z(n66) );
  XNOR U88 ( .A(n71), .B(n66), .Z(n74) );
  XNOR U89 ( .A(n75), .B(sreg[11]), .Z(n69) );
  XNOR U90 ( .A(n74), .B(n69), .Z(c[11]) );
  NAND U91 ( .A(a[6]), .B(b[0]), .Z(n78) );
  AND U92 ( .A(b[1]), .B(a[5]), .Z(n77) );
  XNOR U93 ( .A(n79), .B(n77), .Z(n73) );
  XNOR U94 ( .A(n78), .B(n73), .Z(n80) );
  XNOR U95 ( .A(n81), .B(sreg[12]), .Z(n76) );
  XNOR U96 ( .A(n80), .B(n76), .Z(c[12]) );
  AND U97 ( .A(b[1]), .B(a[6]), .Z(n85) );
  NAND U98 ( .A(b[0]), .B(a[7]), .Z(n86) );
  XNOR U99 ( .A(n85), .B(n86), .Z(n88) );
  XNOR U100 ( .A(n88), .B(n87), .Z(n83) );
  XNOR U101 ( .A(n84), .B(sreg[13]), .Z(n82) );
  XNOR U102 ( .A(n83), .B(n82), .Z(c[13]) );
  NANDN U103 ( .A(n86), .B(n85), .Z(n90) );
  NAND U104 ( .A(n88), .B(n87), .Z(n89) );
  AND U105 ( .A(n90), .B(n89), .Z(n94) );
  AND U106 ( .A(b[1]), .B(a[7]), .Z(n92) );
  XNOR U107 ( .A(n94), .B(n92), .Z(n91) );
  XNOR U108 ( .A(n93), .B(n91), .Z(c[14]) );
endmodule

