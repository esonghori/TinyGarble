
module mult_N64_CC4 ( clk, rst, a, b, c );
  input [63:0] a;
  input [15:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094;
  wire   [127:0] sreg;

  DFF \sreg_reg[111]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[110]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[109]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[108]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[107]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[106]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[105]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[104]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[103]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[102]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[101]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[100]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[99]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[98]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[97]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[96]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[95]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[55]) );
  DFF \sreg_reg[54]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[54]) );
  DFF \sreg_reg[53]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[53]) );
  DFF \sreg_reg[52]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[52]) );
  DFF \sreg_reg[51]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[51]) );
  DFF \sreg_reg[50]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[50]) );
  DFF \sreg_reg[49]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[49]) );
  DFF \sreg_reg[48]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[48]) );
  DFF \sreg_reg[47]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U19 ( .A(n4501), .B(n4500), .Z(n4509) );
  XOR U20 ( .A(n4138), .B(n4137), .Z(n4139) );
  XOR U21 ( .A(n4341), .B(n4340), .Z(n4342) );
  XOR U22 ( .A(n4616), .B(n4615), .Z(n4617) );
  NAND U23 ( .A(n4648), .B(n5012), .Z(n1) );
  NANDN U24 ( .A(n43), .B(n4701), .Z(n2) );
  AND U25 ( .A(n1), .B(n2), .Z(n4682) );
  NAND U26 ( .A(n4755), .B(n4707), .Z(n3) );
  NANDN U27 ( .A(n4756), .B(n4708), .Z(n4) );
  NAND U28 ( .A(n3), .B(n4), .Z(n4772) );
  NAND U29 ( .A(n4950), .B(n4745), .Z(n5) );
  NANDN U30 ( .A(n4815), .B(n4863), .Z(n6) );
  NAND U31 ( .A(n5), .B(n6), .Z(n4806) );
  XNOR U32 ( .A(n4273), .B(n4272), .Z(n4243) );
  XNOR U33 ( .A(n4373), .B(n4372), .Z(n4325) );
  XNOR U34 ( .A(n4442), .B(n4441), .Z(n4396) );
  XNOR U35 ( .A(n4512), .B(n4511), .Z(n4465) );
  XOR U36 ( .A(n4658), .B(n4657), .Z(n4611) );
  NAND U37 ( .A(n4862), .B(n4950), .Z(n7) );
  NANDN U38 ( .A(n4903), .B(n4863), .Z(n8) );
  NAND U39 ( .A(n7), .B(n8), .Z(n4906) );
  XNOR U40 ( .A(n4892), .B(n4891), .Z(n4912) );
  XOR U41 ( .A(n4955), .B(n4954), .Z(n4957) );
  XOR U42 ( .A(n4977), .B(n4976), .Z(n4970) );
  NAND U43 ( .A(n5012), .B(n4984), .Z(n9) );
  NANDN U44 ( .A(n5013), .B(n4985), .Z(n10) );
  NAND U45 ( .A(n9), .B(n10), .Z(n5000) );
  NANDN U46 ( .A(b[0]), .B(a[63]), .Z(n11) );
  AND U47 ( .A(b[1]), .B(n11), .Z(n4424) );
  XOR U48 ( .A(n4182), .B(n4181), .Z(n4183) );
  XOR U49 ( .A(n4188), .B(n4187), .Z(n4189) );
  XOR U50 ( .A(n4286), .B(n4285), .Z(n4287) );
  XOR U51 ( .A(n4292), .B(n4291), .Z(n4293) );
  XOR U52 ( .A(n4506), .B(n4505), .Z(n4510) );
  XOR U53 ( .A(n4568), .B(n4567), .Z(n4541) );
  XOR U54 ( .A(n4628), .B(n4627), .Z(n4630) );
  XOR U55 ( .A(n4618), .B(n4617), .Z(n4649) );
  XNOR U56 ( .A(n4695), .B(n4694), .Z(n4681) );
  XOR U57 ( .A(n4804), .B(n4803), .Z(n4805) );
  NANDN U58 ( .A(n4121), .B(n4120), .Z(n12) );
  NANDN U59 ( .A(n4118), .B(n4119), .Z(n13) );
  AND U60 ( .A(n12), .B(n13), .Z(n4167) );
  XOR U61 ( .A(n4448), .B(n4447), .Z(n4399) );
  XOR U62 ( .A(n4518), .B(n4517), .Z(n4468) );
  XOR U63 ( .A(n4792), .B(n4791), .Z(n4793) );
  XOR U64 ( .A(n4848), .B(n4847), .Z(n4850) );
  XNOR U65 ( .A(n4909), .B(n4908), .Z(n4914) );
  XOR U66 ( .A(n4933), .B(n4932), .Z(n4934) );
  XOR U67 ( .A(n4969), .B(n4968), .Z(n4971) );
  XOR U68 ( .A(n4304), .B(n4303), .Z(n4305) );
  XOR U69 ( .A(n4383), .B(n4382), .Z(n4384) );
  XOR U70 ( .A(n4604), .B(n4603), .Z(n4605) );
  XOR U71 ( .A(n5001), .B(n5000), .Z(n5003) );
  XOR U72 ( .A(n4424), .B(n4423), .Z(n4425) );
  XNOR U73 ( .A(n4140), .B(n4139), .Z(n4118) );
  XOR U74 ( .A(n4347), .B(n4346), .Z(n4348) );
  XOR U75 ( .A(n4412), .B(n4411), .Z(n4413) );
  XOR U76 ( .A(n4420), .B(n4419), .Z(n4439) );
  XOR U77 ( .A(n4494), .B(n4493), .Z(n4495) );
  NAND U78 ( .A(n4471), .B(n4435), .Z(n14) );
  NANDN U79 ( .A(n4472), .B(n33), .Z(n15) );
  NAND U80 ( .A(n14), .B(n15), .Z(n4501) );
  XOR U81 ( .A(n4578), .B(n4577), .Z(n4579) );
  XOR U82 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U83 ( .A(n36), .B(n4559), .Z(n16) );
  NANDN U84 ( .A(n4636), .B(n4560), .Z(n17) );
  NAND U85 ( .A(n16), .B(n17), .Z(n4628) );
  XOR U86 ( .A(n4760), .B(n4759), .Z(n4761) );
  XOR U87 ( .A(n4768), .B(n4767), .Z(n4773) );
  NAND U88 ( .A(n41), .B(n4809), .Z(n18) );
  NANDN U89 ( .A(n4867), .B(n4810), .Z(n19) );
  NAND U90 ( .A(n18), .B(n19), .Z(n4871) );
  XNOR U91 ( .A(n4184), .B(n4183), .Z(n4220) );
  XNOR U92 ( .A(n4217), .B(n4216), .Z(n4166) );
  XNOR U93 ( .A(n4288), .B(n4287), .Z(n4297) );
  XOR U94 ( .A(n4379), .B(n4378), .Z(n4327) );
  XOR U95 ( .A(n4610), .B(n4609), .Z(n4612) );
  XOR U96 ( .A(n4452), .B(n4451), .Z(n4453) );
  XOR U97 ( .A(n4522), .B(n4521), .Z(n4523) );
  XNOR U98 ( .A(n4538), .B(n4537), .Z(n4589) );
  XNOR U99 ( .A(n4678), .B(n4677), .Z(n4669) );
  XNOR U100 ( .A(n4736), .B(n4735), .Z(n4727) );
  XOR U101 ( .A(n4786), .B(n4785), .Z(n4787) );
  XOR U102 ( .A(n4844), .B(n4843), .Z(n4835) );
  XOR U103 ( .A(n4885), .B(n4884), .Z(n4886) );
  XOR U104 ( .A(n4927), .B(n4926), .Z(n4929) );
  XOR U105 ( .A(n4987), .B(n4986), .Z(n4988) );
  XOR U106 ( .A(n5020), .B(n5019), .Z(n5021) );
  NANDN U107 ( .A(n95), .B(n94), .Z(n20) );
  NANDN U108 ( .A(n92), .B(n93), .Z(n21) );
  AND U109 ( .A(n20), .B(n21), .Z(n126) );
  XOR U110 ( .A(n4320), .B(n4319), .Z(n4321) );
  XOR U111 ( .A(n4606), .B(n4605), .Z(n4597) );
  XOR U112 ( .A(n5034), .B(n5033), .Z(n5035) );
  XOR U113 ( .A(n5074), .B(n5075), .Z(n5077) );
  XOR U114 ( .A(n4194), .B(n4193), .Z(n4195) );
  XOR U115 ( .A(n4250), .B(n4249), .Z(n4251) );
  XOR U116 ( .A(n4353), .B(n4352), .Z(n4354) );
  XOR U117 ( .A(n4190), .B(n4189), .Z(n4214) );
  XOR U118 ( .A(n4294), .B(n4293), .Z(n4270) );
  XOR U119 ( .A(n4349), .B(n4348), .Z(n4370) );
  XOR U120 ( .A(n4418), .B(n4417), .Z(n4419) );
  XOR U121 ( .A(n4426), .B(n4425), .Z(n4440) );
  XOR U122 ( .A(n4542), .B(n4541), .Z(n4543) );
  XOR U123 ( .A(n4650), .B(n4649), .Z(n4652) );
  XOR U124 ( .A(n4693), .B(n4692), .Z(n4694) );
  XNOR U125 ( .A(n4689), .B(n4688), .Z(n4683) );
  XOR U126 ( .A(n4772), .B(n4771), .Z(n4774) );
  XOR U127 ( .A(n4871), .B(n4870), .Z(n4873) );
  NANDN U128 ( .A(n618), .B(n619), .Z(n22) );
  NANDN U129 ( .A(n617), .B(n616), .Z(n23) );
  NAND U130 ( .A(n22), .B(n23), .Z(n637) );
  XOR U131 ( .A(n4223), .B(n4222), .Z(n4168) );
  NAND U132 ( .A(n4096), .B(n4095), .Z(n24) );
  NANDN U133 ( .A(n4093), .B(n4094), .Z(n25) );
  AND U134 ( .A(n24), .B(n25), .Z(n4229) );
  XOR U135 ( .A(n4300), .B(n4299), .Z(n4246) );
  XNOR U136 ( .A(n4343), .B(n4342), .Z(n4376) );
  XNOR U137 ( .A(n4414), .B(n4413), .Z(n4445) );
  XNOR U138 ( .A(n4496), .B(n4495), .Z(n4515) );
  XOR U139 ( .A(n4584), .B(n4583), .Z(n4585) );
  XOR U140 ( .A(n4536), .B(n4535), .Z(n4537) );
  XOR U141 ( .A(n4656), .B(n4655), .Z(n4657) );
  XOR U142 ( .A(n4714), .B(n4713), .Z(n4715) );
  XNOR U143 ( .A(n4762), .B(n4761), .Z(n4740) );
  XNOR U144 ( .A(n4806), .B(n4805), .Z(n4798) );
  XOR U145 ( .A(n4842), .B(n4841), .Z(n4843) );
  XOR U146 ( .A(n4907), .B(n4906), .Z(n4908) );
  XOR U147 ( .A(n5007), .B(n5006), .Z(n5008) );
  XOR U148 ( .A(n4788), .B(n4787), .Z(n4779) );
  XOR U149 ( .A(n4989), .B(n4988), .Z(n4962) );
  XNOR U150 ( .A(n5022), .B(n5021), .Z(n4995) );
  XNOR U151 ( .A(n5036), .B(n5035), .Z(n5027) );
  XOR U152 ( .A(n82), .B(n80), .Z(n26) );
  NANDN U153 ( .A(n81), .B(n26), .Z(n27) );
  NAND U154 ( .A(n82), .B(n80), .Z(n28) );
  AND U155 ( .A(n27), .B(n28), .Z(n95) );
  XOR U156 ( .A(n4391), .B(n4390), .Z(n4392) );
  XOR U157 ( .A(n4322), .B(n4321), .Z(n4314) );
  XOR U158 ( .A(n4460), .B(n4459), .Z(n4461) );
  XOR U159 ( .A(n4530), .B(n4529), .Z(n4531) );
  XOR U160 ( .A(n4598), .B(n4597), .Z(n4599) );
  XOR U161 ( .A(n4664), .B(n4663), .Z(n4665) );
  XOR U162 ( .A(n4722), .B(n4721), .Z(n4723) );
  XOR U163 ( .A(n4830), .B(n4829), .Z(n4831) );
  XOR U164 ( .A(n4921), .B(n4920), .Z(n4922) );
  XNOR U165 ( .A(n5083), .B(n5082), .Z(n5076) );
  XNOR U166 ( .A(b[2]), .B(b[1]), .Z(n29) );
  NAND U167 ( .A(n135), .B(n35), .Z(n30) );
  NAND U168 ( .A(n594), .B(n5051), .Z(n31) );
  NAND U169 ( .A(n300), .B(n39), .Z(n32) );
  IV U170 ( .A(n29), .Z(n33) );
  IV U171 ( .A(n4471), .Z(n34) );
  IV U172 ( .A(n4560), .Z(n35) );
  IV U173 ( .A(n30), .Z(n36) );
  IV U174 ( .A(n4708), .Z(n37) );
  IV U175 ( .A(n4755), .Z(n38) );
  IV U176 ( .A(n4810), .Z(n39) );
  IV U177 ( .A(n4863), .Z(n40) );
  IV U178 ( .A(n32), .Z(n41) );
  IV U179 ( .A(n31), .Z(n42) );
  IV U180 ( .A(n4985), .Z(n43) );
  AND U181 ( .A(b[0]), .B(a[0]), .Z(n45) );
  XOR U182 ( .A(n45), .B(sreg[48]), .Z(c[48]) );
  AND U183 ( .A(b[0]), .B(a[1]), .Z(n52) );
  NAND U184 ( .A(a[0]), .B(b[1]), .Z(n44) );
  XOR U185 ( .A(n52), .B(n44), .Z(n46) );
  XNOR U186 ( .A(sreg[49]), .B(n46), .Z(n48) );
  AND U187 ( .A(n45), .B(sreg[48]), .Z(n47) );
  XOR U188 ( .A(n48), .B(n47), .Z(c[49]) );
  NANDN U189 ( .A(n46), .B(sreg[49]), .Z(n50) );
  NAND U190 ( .A(n48), .B(n47), .Z(n49) );
  AND U191 ( .A(n50), .B(n49), .Z(n70) );
  XNOR U192 ( .A(n70), .B(sreg[50]), .Z(n72) );
  NAND U193 ( .A(a[0]), .B(b[2]), .Z(n51) );
  XNOR U194 ( .A(b[1]), .B(n51), .Z(n54) );
  NANDN U195 ( .A(a[0]), .B(n52), .Z(n53) );
  NAND U196 ( .A(n54), .B(n53), .Z(n58) );
  AND U197 ( .A(b[0]), .B(a[2]), .Z(n55) );
  XOR U198 ( .A(b[1]), .B(n55), .Z(n57) );
  NANDN U199 ( .A(b[0]), .B(a[1]), .Z(n56) );
  AND U200 ( .A(n57), .B(n56), .Z(n59) );
  XNOR U201 ( .A(n58), .B(n59), .Z(n71) );
  XOR U202 ( .A(n72), .B(n71), .Z(c[50]) );
  ANDN U203 ( .B(n59), .A(n58), .Z(n82) );
  XOR U204 ( .A(b[3]), .B(b[2]), .Z(n83) );
  XOR U205 ( .A(b[3]), .B(a[0]), .Z(n60) );
  NAND U206 ( .A(n83), .B(n60), .Z(n61) );
  NANDN U207 ( .A(n61), .B(n29), .Z(n63) );
  XOR U208 ( .A(b[3]), .B(a[1]), .Z(n84) );
  NANDN U209 ( .A(n29), .B(n84), .Z(n62) );
  AND U210 ( .A(n63), .B(n62), .Z(n91) );
  NAND U211 ( .A(b[0]), .B(a[3]), .Z(n64) );
  XNOR U212 ( .A(b[1]), .B(n64), .Z(n66) );
  NANDN U213 ( .A(b[0]), .B(a[2]), .Z(n65) );
  NAND U214 ( .A(n66), .B(n65), .Z(n90) );
  XNOR U215 ( .A(n91), .B(n90), .Z(n81) );
  NAND U216 ( .A(n33), .B(a[0]), .Z(n68) );
  NANDN U217 ( .A(b[2]), .B(b[3]), .Z(n67) );
  NAND U218 ( .A(n33), .B(b[3]), .Z(n4474) );
  AND U219 ( .A(n67), .B(n4474), .Z(n4622) );
  IV U220 ( .A(n4622), .Z(n4564) );
  AND U221 ( .A(n68), .B(n4564), .Z(n80) );
  XOR U222 ( .A(n81), .B(n80), .Z(n69) );
  XOR U223 ( .A(n82), .B(n69), .Z(n75) );
  XNOR U224 ( .A(sreg[51]), .B(n75), .Z(n77) );
  NANDN U225 ( .A(n70), .B(sreg[50]), .Z(n74) );
  NAND U226 ( .A(n72), .B(n71), .Z(n73) );
  NAND U227 ( .A(n74), .B(n73), .Z(n76) );
  XOR U228 ( .A(n77), .B(n76), .Z(c[51]) );
  NANDN U229 ( .A(n75), .B(sreg[51]), .Z(n79) );
  NAND U230 ( .A(n77), .B(n76), .Z(n78) );
  AND U231 ( .A(n79), .B(n78), .Z(n113) );
  XNOR U232 ( .A(n113), .B(sreg[52]), .Z(n115) );
  AND U233 ( .A(n83), .B(n29), .Z(n4471) );
  NAND U234 ( .A(n4471), .B(n84), .Z(n86) );
  XOR U235 ( .A(b[3]), .B(a[2]), .Z(n96) );
  NAND U236 ( .A(n33), .B(n96), .Z(n85) );
  AND U237 ( .A(n86), .B(n85), .Z(n110) );
  XOR U238 ( .A(b[4]), .B(b[3]), .Z(n4560) );
  AND U239 ( .A(a[0]), .B(n4560), .Z(n107) );
  NAND U240 ( .A(b[0]), .B(a[4]), .Z(n87) );
  XNOR U241 ( .A(b[1]), .B(n87), .Z(n89) );
  NANDN U242 ( .A(b[0]), .B(a[3]), .Z(n88) );
  NAND U243 ( .A(n89), .B(n88), .Z(n108) );
  XNOR U244 ( .A(n107), .B(n108), .Z(n109) );
  XNOR U245 ( .A(n110), .B(n109), .Z(n93) );
  OR U246 ( .A(n91), .B(n90), .Z(n92) );
  XNOR U247 ( .A(n93), .B(n92), .Z(n94) );
  XNOR U248 ( .A(n95), .B(n94), .Z(n114) );
  XOR U249 ( .A(n115), .B(n114), .Z(c[52]) );
  NAND U250 ( .A(n4471), .B(n96), .Z(n98) );
  XOR U251 ( .A(b[3]), .B(a[3]), .Z(n129) );
  NAND U252 ( .A(n33), .B(n129), .Z(n97) );
  AND U253 ( .A(n98), .B(n97), .Z(n142) );
  NANDN U254 ( .A(b[4]), .B(b[5]), .Z(n99) );
  NAND U255 ( .A(n4560), .B(b[5]), .Z(n4638) );
  NAND U256 ( .A(n99), .B(n4638), .Z(n4766) );
  ANDN U257 ( .B(n4766), .A(n107), .Z(n141) );
  XNOR U258 ( .A(n142), .B(n141), .Z(n144) );
  NAND U259 ( .A(b[0]), .B(a[5]), .Z(n100) );
  XNOR U260 ( .A(b[1]), .B(n100), .Z(n102) );
  NANDN U261 ( .A(b[0]), .B(a[4]), .Z(n101) );
  NAND U262 ( .A(n102), .B(n101), .Z(n139) );
  XOR U263 ( .A(b[5]), .B(b[4]), .Z(n135) );
  XOR U264 ( .A(b[5]), .B(a[0]), .Z(n103) );
  NAND U265 ( .A(n135), .B(n103), .Z(n104) );
  NANDN U266 ( .A(n104), .B(n35), .Z(n106) );
  XOR U267 ( .A(b[5]), .B(a[1]), .Z(n136) );
  NANDN U268 ( .A(n35), .B(n136), .Z(n105) );
  NAND U269 ( .A(n106), .B(n105), .Z(n140) );
  XNOR U270 ( .A(n139), .B(n140), .Z(n143) );
  XOR U271 ( .A(n144), .B(n143), .Z(n124) );
  NANDN U272 ( .A(n108), .B(n107), .Z(n112) );
  NANDN U273 ( .A(n110), .B(n109), .Z(n111) );
  AND U274 ( .A(n112), .B(n111), .Z(n123) );
  XNOR U275 ( .A(n124), .B(n123), .Z(n125) );
  XOR U276 ( .A(n126), .B(n125), .Z(n118) );
  XNOR U277 ( .A(n118), .B(sreg[53]), .Z(n120) );
  NANDN U278 ( .A(n113), .B(sreg[52]), .Z(n117) );
  NAND U279 ( .A(n115), .B(n114), .Z(n116) );
  NAND U280 ( .A(n117), .B(n116), .Z(n119) );
  XOR U281 ( .A(n120), .B(n119), .Z(c[53]) );
  NANDN U282 ( .A(n118), .B(sreg[53]), .Z(n122) );
  NAND U283 ( .A(n120), .B(n119), .Z(n121) );
  AND U284 ( .A(n122), .B(n121), .Z(n179) );
  XNOR U285 ( .A(n179), .B(sreg[54]), .Z(n181) );
  NANDN U286 ( .A(n124), .B(n123), .Z(n128) );
  NAND U287 ( .A(n126), .B(n125), .Z(n127) );
  AND U288 ( .A(n128), .B(n127), .Z(n149) );
  NAND U289 ( .A(n4471), .B(n129), .Z(n131) );
  XOR U290 ( .A(b[3]), .B(a[4]), .Z(n170) );
  NAND U291 ( .A(n33), .B(n170), .Z(n130) );
  AND U292 ( .A(n131), .B(n130), .Z(n155) );
  XOR U293 ( .A(b[6]), .B(b[5]), .Z(n4708) );
  AND U294 ( .A(a[0]), .B(n4708), .Z(n166) );
  NAND U295 ( .A(b[0]), .B(a[6]), .Z(n132) );
  XNOR U296 ( .A(b[1]), .B(n132), .Z(n134) );
  NANDN U297 ( .A(b[0]), .B(a[5]), .Z(n133) );
  NAND U298 ( .A(n134), .B(n133), .Z(n153) );
  XNOR U299 ( .A(n166), .B(n153), .Z(n154) );
  XNOR U300 ( .A(n155), .B(n154), .Z(n176) );
  NAND U301 ( .A(n36), .B(n136), .Z(n138) );
  XOR U302 ( .A(b[5]), .B(a[2]), .Z(n162) );
  NAND U303 ( .A(n4560), .B(n162), .Z(n137) );
  AND U304 ( .A(n138), .B(n137), .Z(n174) );
  ANDN U305 ( .B(n140), .A(n139), .Z(n173) );
  XNOR U306 ( .A(n174), .B(n173), .Z(n175) );
  XOR U307 ( .A(n176), .B(n175), .Z(n148) );
  NANDN U308 ( .A(n142), .B(n141), .Z(n146) );
  NAND U309 ( .A(n144), .B(n143), .Z(n145) );
  AND U310 ( .A(n146), .B(n145), .Z(n147) );
  XOR U311 ( .A(n148), .B(n147), .Z(n150) );
  XNOR U312 ( .A(n149), .B(n150), .Z(n180) );
  XOR U313 ( .A(n181), .B(n180), .Z(c[54]) );
  NANDN U314 ( .A(n148), .B(n147), .Z(n152) );
  OR U315 ( .A(n150), .B(n149), .Z(n151) );
  AND U316 ( .A(n152), .B(n151), .Z(n191) );
  NANDN U317 ( .A(n153), .B(n166), .Z(n157) );
  NANDN U318 ( .A(n155), .B(n154), .Z(n156) );
  AND U319 ( .A(n157), .B(n156), .Z(n197) );
  XOR U320 ( .A(b[7]), .B(b[6]), .Z(n207) );
  XOR U321 ( .A(b[7]), .B(a[0]), .Z(n158) );
  NAND U322 ( .A(n207), .B(n158), .Z(n159) );
  NANDN U323 ( .A(n159), .B(n37), .Z(n161) );
  XOR U324 ( .A(b[7]), .B(a[1]), .Z(n208) );
  NANDN U325 ( .A(n37), .B(n208), .Z(n160) );
  AND U326 ( .A(n161), .B(n160), .Z(n215) );
  NAND U327 ( .A(n36), .B(n162), .Z(n164) );
  XOR U328 ( .A(b[5]), .B(a[3]), .Z(n219) );
  NAND U329 ( .A(n4560), .B(n219), .Z(n163) );
  AND U330 ( .A(n164), .B(n163), .Z(n214) );
  XOR U331 ( .A(n215), .B(n214), .Z(n204) );
  NANDN U332 ( .A(b[6]), .B(b[7]), .Z(n165) );
  NAND U333 ( .A(n4708), .B(b[7]), .Z(n4758) );
  AND U334 ( .A(n165), .B(n4758), .Z(n4854) );
  IV U335 ( .A(n4854), .Z(n4814) );
  ANDN U336 ( .B(n4814), .A(n166), .Z(n202) );
  NAND U337 ( .A(b[0]), .B(a[7]), .Z(n167) );
  XNOR U338 ( .A(b[1]), .B(n167), .Z(n169) );
  NANDN U339 ( .A(b[0]), .B(a[6]), .Z(n168) );
  NAND U340 ( .A(n169), .B(n168), .Z(n201) );
  XNOR U341 ( .A(n202), .B(n201), .Z(n203) );
  XNOR U342 ( .A(n204), .B(n203), .Z(n195) );
  NANDN U343 ( .A(n34), .B(n170), .Z(n172) );
  XNOR U344 ( .A(b[3]), .B(a[5]), .Z(n211) );
  OR U345 ( .A(n211), .B(n29), .Z(n171) );
  NAND U346 ( .A(n172), .B(n171), .Z(n196) );
  XOR U347 ( .A(n195), .B(n196), .Z(n198) );
  XNOR U348 ( .A(n197), .B(n198), .Z(n189) );
  NANDN U349 ( .A(n174), .B(n173), .Z(n178) );
  NAND U350 ( .A(n176), .B(n175), .Z(n177) );
  NAND U351 ( .A(n178), .B(n177), .Z(n190) );
  XOR U352 ( .A(n189), .B(n190), .Z(n192) );
  XOR U353 ( .A(n191), .B(n192), .Z(n184) );
  XNOR U354 ( .A(n184), .B(sreg[55]), .Z(n186) );
  NANDN U355 ( .A(n179), .B(sreg[54]), .Z(n183) );
  NAND U356 ( .A(n181), .B(n180), .Z(n182) );
  NAND U357 ( .A(n183), .B(n182), .Z(n185) );
  XOR U358 ( .A(n186), .B(n185), .Z(c[55]) );
  NANDN U359 ( .A(n184), .B(sreg[55]), .Z(n188) );
  NAND U360 ( .A(n186), .B(n185), .Z(n187) );
  AND U361 ( .A(n188), .B(n187), .Z(n263) );
  XNOR U362 ( .A(n263), .B(sreg[56]), .Z(n265) );
  NANDN U363 ( .A(n190), .B(n189), .Z(n194) );
  OR U364 ( .A(n192), .B(n191), .Z(n193) );
  AND U365 ( .A(n194), .B(n193), .Z(n259) );
  NANDN U366 ( .A(n196), .B(n195), .Z(n200) );
  NANDN U367 ( .A(n198), .B(n197), .Z(n199) );
  AND U368 ( .A(n200), .B(n199), .Z(n258) );
  NANDN U369 ( .A(n202), .B(n201), .Z(n206) );
  NANDN U370 ( .A(n204), .B(n203), .Z(n205) );
  AND U371 ( .A(n206), .B(n205), .Z(n225) );
  AND U372 ( .A(n207), .B(n37), .Z(n4755) );
  NAND U373 ( .A(n4755), .B(n208), .Z(n210) );
  XOR U374 ( .A(b[7]), .B(a[2]), .Z(n239) );
  NAND U375 ( .A(n4708), .B(n239), .Z(n209) );
  AND U376 ( .A(n210), .B(n209), .Z(n229) );
  OR U377 ( .A(n211), .B(n34), .Z(n213) );
  XOR U378 ( .A(b[3]), .B(a[6]), .Z(n254) );
  NAND U379 ( .A(n33), .B(n254), .Z(n212) );
  NAND U380 ( .A(n213), .B(n212), .Z(n228) );
  XNOR U381 ( .A(n229), .B(n228), .Z(n231) );
  NOR U382 ( .A(n215), .B(n214), .Z(n230) );
  XOR U383 ( .A(n231), .B(n230), .Z(n223) );
  NAND U384 ( .A(b[0]), .B(a[8]), .Z(n216) );
  XNOR U385 ( .A(b[1]), .B(n216), .Z(n218) );
  NANDN U386 ( .A(b[0]), .B(a[7]), .Z(n217) );
  NAND U387 ( .A(n218), .B(n217), .Z(n236) );
  XOR U388 ( .A(b[8]), .B(b[7]), .Z(n4810) );
  AND U389 ( .A(a[0]), .B(n4810), .Z(n247) );
  NAND U390 ( .A(n36), .B(n219), .Z(n221) );
  XOR U391 ( .A(b[5]), .B(a[4]), .Z(n248) );
  NAND U392 ( .A(n4560), .B(n248), .Z(n220) );
  AND U393 ( .A(n221), .B(n220), .Z(n234) );
  XOR U394 ( .A(n247), .B(n234), .Z(n235) );
  XNOR U395 ( .A(n236), .B(n235), .Z(n222) );
  XNOR U396 ( .A(n223), .B(n222), .Z(n224) );
  XNOR U397 ( .A(n225), .B(n224), .Z(n257) );
  XOR U398 ( .A(n258), .B(n257), .Z(n260) );
  XNOR U399 ( .A(n259), .B(n260), .Z(n264) );
  XOR U400 ( .A(n265), .B(n264), .Z(c[56]) );
  NANDN U401 ( .A(n223), .B(n222), .Z(n227) );
  NANDN U402 ( .A(n225), .B(n224), .Z(n226) );
  AND U403 ( .A(n227), .B(n226), .Z(n273) );
  NANDN U404 ( .A(n229), .B(n228), .Z(n233) );
  NAND U405 ( .A(n231), .B(n230), .Z(n232) );
  AND U406 ( .A(n233), .B(n232), .Z(n312) );
  NANDN U407 ( .A(n234), .B(n247), .Z(n238) );
  OR U408 ( .A(n236), .B(n235), .Z(n237) );
  AND U409 ( .A(n238), .B(n237), .Z(n310) );
  NAND U410 ( .A(n4755), .B(n239), .Z(n241) );
  XOR U411 ( .A(b[7]), .B(a[3]), .Z(n294) );
  NAND U412 ( .A(n4708), .B(n294), .Z(n240) );
  AND U413 ( .A(n241), .B(n240), .Z(n304) );
  XOR U414 ( .A(b[9]), .B(b[8]), .Z(n300) );
  XOR U415 ( .A(b[9]), .B(a[0]), .Z(n242) );
  NAND U416 ( .A(n300), .B(n242), .Z(n243) );
  NANDN U417 ( .A(n243), .B(n39), .Z(n245) );
  XOR U418 ( .A(b[9]), .B(a[1]), .Z(n301) );
  NANDN U419 ( .A(n39), .B(n301), .Z(n244) );
  NAND U420 ( .A(n245), .B(n244), .Z(n305) );
  XOR U421 ( .A(n304), .B(n305), .Z(n281) );
  NANDN U422 ( .A(b[8]), .B(b[9]), .Z(n246) );
  NAND U423 ( .A(n4810), .B(b[9]), .Z(n4869) );
  AND U424 ( .A(n246), .B(n4869), .Z(n4942) );
  IV U425 ( .A(n4942), .Z(n4901) );
  ANDN U426 ( .B(n4901), .A(n247), .Z(n280) );
  NAND U427 ( .A(n36), .B(n248), .Z(n250) );
  XOR U428 ( .A(b[5]), .B(a[5]), .Z(n297) );
  NAND U429 ( .A(n4560), .B(n297), .Z(n249) );
  AND U430 ( .A(n250), .B(n249), .Z(n279) );
  XOR U431 ( .A(n280), .B(n279), .Z(n282) );
  XOR U432 ( .A(n281), .B(n282), .Z(n288) );
  NAND U433 ( .A(b[0]), .B(a[9]), .Z(n251) );
  XNOR U434 ( .A(b[1]), .B(n251), .Z(n253) );
  NANDN U435 ( .A(b[0]), .B(a[8]), .Z(n252) );
  NAND U436 ( .A(n253), .B(n252), .Z(n286) );
  NAND U437 ( .A(n4471), .B(n254), .Z(n256) );
  XOR U438 ( .A(b[3]), .B(a[7]), .Z(n306) );
  NAND U439 ( .A(n33), .B(n306), .Z(n255) );
  NAND U440 ( .A(n256), .B(n255), .Z(n285) );
  XNOR U441 ( .A(n286), .B(n285), .Z(n287) );
  XOR U442 ( .A(n288), .B(n287), .Z(n309) );
  XNOR U443 ( .A(n310), .B(n309), .Z(n311) );
  XOR U444 ( .A(n312), .B(n311), .Z(n274) );
  XNOR U445 ( .A(n273), .B(n274), .Z(n275) );
  NANDN U446 ( .A(n258), .B(n257), .Z(n262) );
  OR U447 ( .A(n260), .B(n259), .Z(n261) );
  NAND U448 ( .A(n262), .B(n261), .Z(n276) );
  XOR U449 ( .A(n275), .B(n276), .Z(n268) );
  XNOR U450 ( .A(sreg[57]), .B(n268), .Z(n270) );
  NANDN U451 ( .A(n263), .B(sreg[56]), .Z(n267) );
  NAND U452 ( .A(n265), .B(n264), .Z(n266) );
  NAND U453 ( .A(n267), .B(n266), .Z(n269) );
  XOR U454 ( .A(n270), .B(n269), .Z(c[57]) );
  NANDN U455 ( .A(n268), .B(sreg[57]), .Z(n272) );
  NAND U456 ( .A(n270), .B(n269), .Z(n271) );
  AND U457 ( .A(n272), .B(n271), .Z(n365) );
  XNOR U458 ( .A(sreg[58]), .B(n365), .Z(n367) );
  NANDN U459 ( .A(n274), .B(n273), .Z(n278) );
  NANDN U460 ( .A(n276), .B(n275), .Z(n277) );
  AND U461 ( .A(n278), .B(n277), .Z(n317) );
  NANDN U462 ( .A(n280), .B(n279), .Z(n284) );
  NANDN U463 ( .A(n282), .B(n281), .Z(n283) );
  AND U464 ( .A(n284), .B(n283), .Z(n360) );
  NANDN U465 ( .A(n286), .B(n285), .Z(n290) );
  NAND U466 ( .A(n288), .B(n287), .Z(n289) );
  AND U467 ( .A(n290), .B(n289), .Z(n359) );
  XNOR U468 ( .A(n360), .B(n359), .Z(n361) );
  NAND U469 ( .A(b[0]), .B(a[10]), .Z(n291) );
  XNOR U470 ( .A(b[1]), .B(n291), .Z(n293) );
  NANDN U471 ( .A(b[0]), .B(a[9]), .Z(n292) );
  NAND U472 ( .A(n293), .B(n292), .Z(n329) );
  XOR U473 ( .A(b[10]), .B(b[9]), .Z(n4863) );
  AND U474 ( .A(a[0]), .B(n4863), .Z(n358) );
  NAND U475 ( .A(n4755), .B(n294), .Z(n296) );
  XOR U476 ( .A(b[7]), .B(a[4]), .Z(n354) );
  NAND U477 ( .A(n4708), .B(n354), .Z(n295) );
  AND U478 ( .A(n296), .B(n295), .Z(n327) );
  XOR U479 ( .A(n358), .B(n327), .Z(n328) );
  XOR U480 ( .A(n329), .B(n328), .Z(n324) );
  NAND U481 ( .A(n36), .B(n297), .Z(n299) );
  XOR U482 ( .A(b[5]), .B(a[6]), .Z(n348) );
  NAND U483 ( .A(n4560), .B(n348), .Z(n298) );
  AND U484 ( .A(n299), .B(n298), .Z(n333) );
  NAND U485 ( .A(n41), .B(n301), .Z(n303) );
  XOR U486 ( .A(b[9]), .B(a[2]), .Z(n342) );
  NAND U487 ( .A(n4810), .B(n342), .Z(n302) );
  NAND U488 ( .A(n303), .B(n302), .Z(n332) );
  XNOR U489 ( .A(n333), .B(n332), .Z(n335) );
  ANDN U490 ( .B(n305), .A(n304), .Z(n334) );
  XOR U491 ( .A(n335), .B(n334), .Z(n322) );
  NANDN U492 ( .A(n34), .B(n306), .Z(n308) );
  XNOR U493 ( .A(b[3]), .B(a[8]), .Z(n351) );
  OR U494 ( .A(n351), .B(n29), .Z(n307) );
  AND U495 ( .A(n308), .B(n307), .Z(n321) );
  XNOR U496 ( .A(n322), .B(n321), .Z(n323) );
  XOR U497 ( .A(n324), .B(n323), .Z(n362) );
  XNOR U498 ( .A(n361), .B(n362), .Z(n315) );
  NANDN U499 ( .A(n310), .B(n309), .Z(n314) );
  NANDN U500 ( .A(n312), .B(n311), .Z(n313) );
  NAND U501 ( .A(n314), .B(n313), .Z(n316) );
  XOR U502 ( .A(n315), .B(n316), .Z(n318) );
  XNOR U503 ( .A(n317), .B(n318), .Z(n366) );
  XNOR U504 ( .A(n367), .B(n366), .Z(c[58]) );
  NANDN U505 ( .A(n316), .B(n315), .Z(n320) );
  NANDN U506 ( .A(n318), .B(n317), .Z(n319) );
  AND U507 ( .A(n320), .B(n319), .Z(n377) );
  NANDN U508 ( .A(n322), .B(n321), .Z(n326) );
  NANDN U509 ( .A(n324), .B(n323), .Z(n325) );
  AND U510 ( .A(n326), .B(n325), .Z(n423) );
  NANDN U511 ( .A(n327), .B(n358), .Z(n331) );
  OR U512 ( .A(n329), .B(n328), .Z(n330) );
  AND U513 ( .A(n331), .B(n330), .Z(n421) );
  NANDN U514 ( .A(n333), .B(n332), .Z(n337) );
  NAND U515 ( .A(n335), .B(n334), .Z(n336) );
  AND U516 ( .A(n337), .B(n336), .Z(n417) );
  XOR U517 ( .A(b[11]), .B(b[10]), .Z(n392) );
  XOR U518 ( .A(b[11]), .B(a[0]), .Z(n338) );
  NAND U519 ( .A(n392), .B(n338), .Z(n339) );
  NANDN U520 ( .A(n339), .B(n40), .Z(n341) );
  XOR U521 ( .A(b[11]), .B(a[1]), .Z(n393) );
  NANDN U522 ( .A(n40), .B(n393), .Z(n340) );
  AND U523 ( .A(n341), .B(n340), .Z(n382) );
  NAND U524 ( .A(n41), .B(n342), .Z(n344) );
  XOR U525 ( .A(b[9]), .B(a[3]), .Z(n399) );
  NAND U526 ( .A(n4810), .B(n399), .Z(n343) );
  AND U527 ( .A(n344), .B(n343), .Z(n381) );
  XOR U528 ( .A(n382), .B(n381), .Z(n404) );
  NAND U529 ( .A(b[0]), .B(a[11]), .Z(n345) );
  XNOR U530 ( .A(b[1]), .B(n345), .Z(n347) );
  NANDN U531 ( .A(b[0]), .B(a[10]), .Z(n346) );
  NAND U532 ( .A(n347), .B(n346), .Z(n402) );
  NANDN U533 ( .A(n30), .B(n348), .Z(n350) );
  XNOR U534 ( .A(b[5]), .B(a[7]), .Z(n389) );
  OR U535 ( .A(n389), .B(n35), .Z(n349) );
  NAND U536 ( .A(n350), .B(n349), .Z(n403) );
  XOR U537 ( .A(n402), .B(n403), .Z(n405) );
  XOR U538 ( .A(n404), .B(n405), .Z(n415) );
  OR U539 ( .A(n351), .B(n34), .Z(n353) );
  XOR U540 ( .A(b[3]), .B(a[9]), .Z(n383) );
  NAND U541 ( .A(n33), .B(n383), .Z(n352) );
  AND U542 ( .A(n353), .B(n352), .Z(n411) );
  NAND U543 ( .A(n4755), .B(n354), .Z(n356) );
  XOR U544 ( .A(b[7]), .B(a[5]), .Z(n386) );
  NAND U545 ( .A(n4708), .B(n386), .Z(n355) );
  AND U546 ( .A(n356), .B(n355), .Z(n409) );
  NANDN U547 ( .A(b[10]), .B(b[11]), .Z(n357) );
  NAND U548 ( .A(n4863), .B(b[11]), .Z(n4953) );
  AND U549 ( .A(n357), .B(n4953), .Z(n5007) );
  NOR U550 ( .A(n5007), .B(n358), .Z(n408) );
  XNOR U551 ( .A(n409), .B(n408), .Z(n410) );
  XNOR U552 ( .A(n411), .B(n410), .Z(n414) );
  XNOR U553 ( .A(n415), .B(n414), .Z(n416) );
  XNOR U554 ( .A(n417), .B(n416), .Z(n420) );
  XNOR U555 ( .A(n421), .B(n420), .Z(n422) );
  XOR U556 ( .A(n423), .B(n422), .Z(n376) );
  NANDN U557 ( .A(n360), .B(n359), .Z(n364) );
  NANDN U558 ( .A(n362), .B(n361), .Z(n363) );
  NAND U559 ( .A(n364), .B(n363), .Z(n375) );
  XOR U560 ( .A(n376), .B(n375), .Z(n378) );
  XOR U561 ( .A(n377), .B(n378), .Z(n370) );
  XNOR U562 ( .A(n370), .B(sreg[59]), .Z(n372) );
  NANDN U563 ( .A(sreg[58]), .B(n365), .Z(n369) );
  NAND U564 ( .A(n367), .B(n366), .Z(n368) );
  AND U565 ( .A(n369), .B(n368), .Z(n371) );
  XOR U566 ( .A(n372), .B(n371), .Z(c[59]) );
  NANDN U567 ( .A(n370), .B(sreg[59]), .Z(n374) );
  NAND U568 ( .A(n372), .B(n371), .Z(n373) );
  AND U569 ( .A(n374), .B(n373), .Z(n485) );
  XNOR U570 ( .A(sreg[60]), .B(n485), .Z(n487) );
  NANDN U571 ( .A(n376), .B(n375), .Z(n380) );
  OR U572 ( .A(n378), .B(n377), .Z(n379) );
  AND U573 ( .A(n380), .B(n379), .Z(n429) );
  NOR U574 ( .A(n382), .B(n381), .Z(n475) );
  NANDN U575 ( .A(n34), .B(n383), .Z(n385) );
  XNOR U576 ( .A(b[3]), .B(a[10]), .Z(n457) );
  OR U577 ( .A(n457), .B(n29), .Z(n384) );
  AND U578 ( .A(n385), .B(n384), .Z(n473) );
  NANDN U579 ( .A(n38), .B(n386), .Z(n388) );
  XNOR U580 ( .A(b[7]), .B(a[6]), .Z(n447) );
  OR U581 ( .A(n447), .B(n37), .Z(n387) );
  NAND U582 ( .A(n388), .B(n387), .Z(n474) );
  XOR U583 ( .A(n473), .B(n474), .Z(n476) );
  XOR U584 ( .A(n475), .B(n476), .Z(n441) );
  OR U585 ( .A(n389), .B(n30), .Z(n391) );
  XOR U586 ( .A(b[5]), .B(a[8]), .Z(n464) );
  NAND U587 ( .A(n4560), .B(n464), .Z(n390) );
  AND U588 ( .A(n391), .B(n390), .Z(n439) );
  AND U589 ( .A(n392), .B(n40), .Z(n4950) );
  NAND U590 ( .A(n4950), .B(n393), .Z(n395) );
  XOR U591 ( .A(b[11]), .B(a[2]), .Z(n454) );
  NAND U592 ( .A(n4863), .B(n454), .Z(n394) );
  NAND U593 ( .A(n395), .B(n394), .Z(n438) );
  XNOR U594 ( .A(n439), .B(n438), .Z(n440) );
  XNOR U595 ( .A(n441), .B(n440), .Z(n435) );
  NAND U596 ( .A(b[0]), .B(a[12]), .Z(n396) );
  XNOR U597 ( .A(b[1]), .B(n396), .Z(n398) );
  NANDN U598 ( .A(b[0]), .B(a[11]), .Z(n397) );
  NAND U599 ( .A(n398), .B(n397), .Z(n470) );
  XOR U600 ( .A(b[12]), .B(b[11]), .Z(n4985) );
  AND U601 ( .A(a[0]), .B(n4985), .Z(n467) );
  NAND U602 ( .A(n41), .B(n399), .Z(n401) );
  XOR U603 ( .A(b[9]), .B(a[4]), .Z(n460) );
  NAND U604 ( .A(n4810), .B(n460), .Z(n400) );
  AND U605 ( .A(n401), .B(n400), .Z(n468) );
  XNOR U606 ( .A(n467), .B(n468), .Z(n469) );
  XNOR U607 ( .A(n470), .B(n469), .Z(n432) );
  NANDN U608 ( .A(n403), .B(n402), .Z(n407) );
  OR U609 ( .A(n405), .B(n404), .Z(n406) );
  NAND U610 ( .A(n407), .B(n406), .Z(n433) );
  XNOR U611 ( .A(n432), .B(n433), .Z(n434) );
  XOR U612 ( .A(n435), .B(n434), .Z(n482) );
  NANDN U613 ( .A(n409), .B(n408), .Z(n413) );
  NANDN U614 ( .A(n411), .B(n410), .Z(n412) );
  AND U615 ( .A(n413), .B(n412), .Z(n479) );
  NANDN U616 ( .A(n415), .B(n414), .Z(n419) );
  NANDN U617 ( .A(n417), .B(n416), .Z(n418) );
  NAND U618 ( .A(n419), .B(n418), .Z(n480) );
  XNOR U619 ( .A(n479), .B(n480), .Z(n481) );
  XNOR U620 ( .A(n482), .B(n481), .Z(n426) );
  NANDN U621 ( .A(n421), .B(n420), .Z(n425) );
  NAND U622 ( .A(n423), .B(n422), .Z(n424) );
  NAND U623 ( .A(n425), .B(n424), .Z(n427) );
  XNOR U624 ( .A(n426), .B(n427), .Z(n428) );
  XNOR U625 ( .A(n429), .B(n428), .Z(n486) );
  XNOR U626 ( .A(n487), .B(n486), .Z(c[60]) );
  NANDN U627 ( .A(n427), .B(n426), .Z(n431) );
  NANDN U628 ( .A(n429), .B(n428), .Z(n430) );
  AND U629 ( .A(n431), .B(n430), .Z(n498) );
  NANDN U630 ( .A(n433), .B(n432), .Z(n437) );
  NAND U631 ( .A(n435), .B(n434), .Z(n436) );
  AND U632 ( .A(n437), .B(n436), .Z(n551) );
  NANDN U633 ( .A(n439), .B(n438), .Z(n443) );
  NANDN U634 ( .A(n441), .B(n440), .Z(n442) );
  AND U635 ( .A(n443), .B(n442), .Z(n550) );
  NAND U636 ( .A(b[0]), .B(a[13]), .Z(n444) );
  XNOR U637 ( .A(b[1]), .B(n444), .Z(n446) );
  NANDN U638 ( .A(b[0]), .B(a[12]), .Z(n445) );
  NAND U639 ( .A(n446), .B(n445), .Z(n535) );
  OR U640 ( .A(n447), .B(n38), .Z(n449) );
  XOR U641 ( .A(b[7]), .B(a[7]), .Z(n528) );
  NAND U642 ( .A(n4708), .B(n528), .Z(n448) );
  NAND U643 ( .A(n449), .B(n448), .Z(n534) );
  XNOR U644 ( .A(n535), .B(n534), .Z(n537) );
  XOR U645 ( .A(b[13]), .B(b[12]), .Z(n540) );
  XOR U646 ( .A(b[13]), .B(a[0]), .Z(n450) );
  NAND U647 ( .A(n540), .B(n450), .Z(n451) );
  NANDN U648 ( .A(n451), .B(n43), .Z(n453) );
  XOR U649 ( .A(b[13]), .B(a[1]), .Z(n541) );
  NANDN U650 ( .A(n43), .B(n541), .Z(n452) );
  AND U651 ( .A(n453), .B(n452), .Z(n548) );
  NAND U652 ( .A(n4950), .B(n454), .Z(n456) );
  XOR U653 ( .A(b[11]), .B(a[3]), .Z(n519) );
  NAND U654 ( .A(n4863), .B(n519), .Z(n455) );
  NAND U655 ( .A(n456), .B(n455), .Z(n547) );
  XNOR U656 ( .A(n548), .B(n547), .Z(n536) );
  XOR U657 ( .A(n537), .B(n536), .Z(n509) );
  OR U658 ( .A(n457), .B(n34), .Z(n459) );
  XOR U659 ( .A(b[3]), .B(a[11]), .Z(n531) );
  NAND U660 ( .A(n33), .B(n531), .Z(n458) );
  AND U661 ( .A(n459), .B(n458), .Z(n514) );
  NAND U662 ( .A(n41), .B(n460), .Z(n462) );
  XOR U663 ( .A(b[9]), .B(a[5]), .Z(n544) );
  NAND U664 ( .A(n4810), .B(n544), .Z(n461) );
  NAND U665 ( .A(n462), .B(n461), .Z(n513) );
  XNOR U666 ( .A(n514), .B(n513), .Z(n516) );
  NANDN U667 ( .A(b[12]), .B(b[13]), .Z(n463) );
  NAND U668 ( .A(n4985), .B(b[13]), .Z(n5015) );
  NAND U669 ( .A(n463), .B(n5015), .Z(n5047) );
  IV U670 ( .A(n5047), .Z(n5055) );
  NOR U671 ( .A(n5055), .B(n467), .Z(n515) );
  XOR U672 ( .A(n516), .B(n515), .Z(n508) );
  NANDN U673 ( .A(n30), .B(n464), .Z(n466) );
  XNOR U674 ( .A(b[5]), .B(a[9]), .Z(n525) );
  OR U675 ( .A(n525), .B(n35), .Z(n465) );
  AND U676 ( .A(n466), .B(n465), .Z(n507) );
  XOR U677 ( .A(n508), .B(n507), .Z(n510) );
  XOR U678 ( .A(n509), .B(n510), .Z(n504) );
  NANDN U679 ( .A(n468), .B(n467), .Z(n472) );
  NANDN U680 ( .A(n470), .B(n469), .Z(n471) );
  AND U681 ( .A(n472), .B(n471), .Z(n502) );
  NANDN U682 ( .A(n474), .B(n473), .Z(n478) );
  OR U683 ( .A(n476), .B(n475), .Z(n477) );
  AND U684 ( .A(n478), .B(n477), .Z(n501) );
  XNOR U685 ( .A(n502), .B(n501), .Z(n503) );
  XNOR U686 ( .A(n504), .B(n503), .Z(n549) );
  XOR U687 ( .A(n550), .B(n549), .Z(n552) );
  XOR U688 ( .A(n551), .B(n552), .Z(n496) );
  NANDN U689 ( .A(n480), .B(n479), .Z(n484) );
  NANDN U690 ( .A(n482), .B(n481), .Z(n483) );
  NAND U691 ( .A(n484), .B(n483), .Z(n495) );
  XNOR U692 ( .A(n496), .B(n495), .Z(n497) );
  XNOR U693 ( .A(n498), .B(n497), .Z(n490) );
  XNOR U694 ( .A(sreg[61]), .B(n490), .Z(n492) );
  NANDN U695 ( .A(sreg[60]), .B(n485), .Z(n489) );
  NAND U696 ( .A(n487), .B(n486), .Z(n488) );
  NAND U697 ( .A(n489), .B(n488), .Z(n491) );
  XNOR U698 ( .A(n492), .B(n491), .Z(c[61]) );
  NANDN U699 ( .A(sreg[61]), .B(n490), .Z(n494) );
  NAND U700 ( .A(n492), .B(n491), .Z(n493) );
  NAND U701 ( .A(n494), .B(n493), .Z(n555) );
  XNOR U702 ( .A(sreg[62]), .B(n555), .Z(n557) );
  NANDN U703 ( .A(n496), .B(n495), .Z(n500) );
  NANDN U704 ( .A(n498), .B(n497), .Z(n499) );
  AND U705 ( .A(n500), .B(n499), .Z(n562) );
  NANDN U706 ( .A(n502), .B(n501), .Z(n506) );
  NANDN U707 ( .A(n504), .B(n503), .Z(n505) );
  AND U708 ( .A(n506), .B(n505), .Z(n622) );
  NANDN U709 ( .A(n508), .B(n507), .Z(n512) );
  OR U710 ( .A(n510), .B(n509), .Z(n511) );
  AND U711 ( .A(n512), .B(n511), .Z(n620) );
  NANDN U712 ( .A(n514), .B(n513), .Z(n518) );
  NAND U713 ( .A(n516), .B(n515), .Z(n517) );
  AND U714 ( .A(n518), .B(n517), .Z(n607) );
  XNOR U715 ( .A(b[13]), .B(b[14]), .Z(n5051) );
  IV U716 ( .A(n5051), .Z(n4981) );
  AND U717 ( .A(a[0]), .B(n4981), .Z(n610) );
  NAND U718 ( .A(n4950), .B(n519), .Z(n521) );
  XOR U719 ( .A(b[11]), .B(a[4]), .Z(n582) );
  NAND U720 ( .A(n4863), .B(n582), .Z(n520) );
  AND U721 ( .A(n521), .B(n520), .Z(n611) );
  XNOR U722 ( .A(n610), .B(n611), .Z(n612) );
  NAND U723 ( .A(b[0]), .B(a[14]), .Z(n522) );
  XNOR U724 ( .A(b[1]), .B(n522), .Z(n524) );
  NANDN U725 ( .A(b[0]), .B(a[13]), .Z(n523) );
  NAND U726 ( .A(n524), .B(n523), .Z(n613) );
  XNOR U727 ( .A(n612), .B(n613), .Z(n604) );
  OR U728 ( .A(n525), .B(n30), .Z(n527) );
  XOR U729 ( .A(b[5]), .B(a[10]), .Z(n576) );
  NAND U730 ( .A(n4560), .B(n576), .Z(n526) );
  AND U731 ( .A(n527), .B(n526), .Z(n588) );
  NAND U732 ( .A(n4755), .B(n528), .Z(n530) );
  XOR U733 ( .A(b[7]), .B(a[8]), .Z(n572) );
  NAND U734 ( .A(n4708), .B(n572), .Z(n529) );
  AND U735 ( .A(n530), .B(n529), .Z(n586) );
  NAND U736 ( .A(n4471), .B(n531), .Z(n533) );
  XOR U737 ( .A(b[3]), .B(a[12]), .Z(n579) );
  NAND U738 ( .A(n33), .B(n579), .Z(n532) );
  NAND U739 ( .A(n533), .B(n532), .Z(n585) );
  XNOR U740 ( .A(n586), .B(n585), .Z(n587) );
  XOR U741 ( .A(n588), .B(n587), .Z(n605) );
  XNOR U742 ( .A(n604), .B(n605), .Z(n606) );
  XNOR U743 ( .A(n607), .B(n606), .Z(n568) );
  NANDN U744 ( .A(n535), .B(n534), .Z(n539) );
  NAND U745 ( .A(n537), .B(n536), .Z(n538) );
  AND U746 ( .A(n539), .B(n538), .Z(n567) );
  AND U747 ( .A(n540), .B(n43), .Z(n5012) );
  NAND U748 ( .A(n5012), .B(n541), .Z(n543) );
  XOR U749 ( .A(b[13]), .B(a[2]), .Z(n591) );
  NAND U750 ( .A(n4985), .B(n591), .Z(n542) );
  AND U751 ( .A(n543), .B(n542), .Z(n617) );
  NAND U752 ( .A(n41), .B(n544), .Z(n546) );
  XOR U753 ( .A(b[9]), .B(a[6]), .Z(n601) );
  NAND U754 ( .A(n4810), .B(n601), .Z(n545) );
  NAND U755 ( .A(n546), .B(n545), .Z(n616) );
  XNOR U756 ( .A(n617), .B(n616), .Z(n619) );
  NANDN U757 ( .A(n548), .B(n547), .Z(n618) );
  XNOR U758 ( .A(n619), .B(n618), .Z(n566) );
  XOR U759 ( .A(n567), .B(n566), .Z(n569) );
  XOR U760 ( .A(n568), .B(n569), .Z(n621) );
  XOR U761 ( .A(n620), .B(n621), .Z(n623) );
  XOR U762 ( .A(n622), .B(n623), .Z(n561) );
  NANDN U763 ( .A(n550), .B(n549), .Z(n554) );
  OR U764 ( .A(n552), .B(n551), .Z(n553) );
  AND U765 ( .A(n554), .B(n553), .Z(n560) );
  XOR U766 ( .A(n561), .B(n560), .Z(n563) );
  XNOR U767 ( .A(n562), .B(n563), .Z(n556) );
  XOR U768 ( .A(n557), .B(n556), .Z(c[62]) );
  NANDN U769 ( .A(n555), .B(sreg[62]), .Z(n559) );
  NAND U770 ( .A(n557), .B(n556), .Z(n558) );
  AND U771 ( .A(n559), .B(n558), .Z(n628) );
  NANDN U772 ( .A(n561), .B(n560), .Z(n565) );
  OR U773 ( .A(n563), .B(n562), .Z(n564) );
  AND U774 ( .A(n565), .B(n564), .Z(n634) );
  NANDN U775 ( .A(n567), .B(n566), .Z(n571) );
  NANDN U776 ( .A(n569), .B(n568), .Z(n570) );
  AND U777 ( .A(n571), .B(n570), .Z(n694) );
  NAND U778 ( .A(n4755), .B(n572), .Z(n574) );
  XOR U779 ( .A(b[7]), .B(a[9]), .Z(n681) );
  NAND U780 ( .A(n4708), .B(n681), .Z(n573) );
  AND U781 ( .A(n574), .B(n573), .Z(n668) );
  NAND U782 ( .A(b[13]), .B(b[14]), .Z(n5089) );
  ANDN U783 ( .B(n5089), .A(n610), .Z(n575) );
  AND U784 ( .A(b[15]), .B(n575), .Z(n667) );
  XNOR U785 ( .A(n668), .B(n667), .Z(n670) );
  NAND U786 ( .A(n36), .B(n576), .Z(n578) );
  XOR U787 ( .A(b[5]), .B(a[11]), .Z(n690) );
  NAND U788 ( .A(n4560), .B(n690), .Z(n577) );
  AND U789 ( .A(n578), .B(n577), .Z(n664) );
  NAND U790 ( .A(n4471), .B(n579), .Z(n581) );
  XOR U791 ( .A(b[3]), .B(a[13]), .Z(n675) );
  NAND U792 ( .A(n33), .B(n675), .Z(n580) );
  AND U793 ( .A(n581), .B(n580), .Z(n662) );
  NAND U794 ( .A(n4950), .B(n582), .Z(n584) );
  XOR U795 ( .A(b[11]), .B(a[5]), .Z(n684) );
  NAND U796 ( .A(n4863), .B(n684), .Z(n583) );
  NAND U797 ( .A(n584), .B(n583), .Z(n661) );
  XNOR U798 ( .A(n662), .B(n661), .Z(n663) );
  XNOR U799 ( .A(n664), .B(n663), .Z(n669) );
  XOR U800 ( .A(n670), .B(n669), .Z(n645) );
  NANDN U801 ( .A(n586), .B(n585), .Z(n590) );
  NANDN U802 ( .A(n588), .B(n587), .Z(n589) );
  AND U803 ( .A(n590), .B(n589), .Z(n643) );
  NAND U804 ( .A(n5012), .B(n591), .Z(n593) );
  XOR U805 ( .A(b[13]), .B(a[3]), .Z(n658) );
  NAND U806 ( .A(n4985), .B(n658), .Z(n592) );
  AND U807 ( .A(n593), .B(n592), .Z(n674) );
  XOR U808 ( .A(b[14]), .B(b[15]), .Z(n594) );
  XOR U809 ( .A(a[0]), .B(b[15]), .Z(n595) );
  NAND U810 ( .A(n42), .B(n595), .Z(n597) );
  XOR U811 ( .A(b[15]), .B(a[1]), .Z(n687) );
  AND U812 ( .A(n687), .B(n4981), .Z(n596) );
  ANDN U813 ( .B(n597), .A(n596), .Z(n673) );
  XOR U814 ( .A(n674), .B(n673), .Z(n652) );
  NAND U815 ( .A(b[0]), .B(a[15]), .Z(n598) );
  XNOR U816 ( .A(b[1]), .B(n598), .Z(n600) );
  NANDN U817 ( .A(b[0]), .B(a[14]), .Z(n599) );
  NAND U818 ( .A(n600), .B(n599), .Z(n649) );
  NANDN U819 ( .A(n32), .B(n601), .Z(n603) );
  XNOR U820 ( .A(b[9]), .B(a[7]), .Z(n678) );
  OR U821 ( .A(n678), .B(n39), .Z(n602) );
  NAND U822 ( .A(n603), .B(n602), .Z(n650) );
  XNOR U823 ( .A(n649), .B(n650), .Z(n651) );
  XOR U824 ( .A(n652), .B(n651), .Z(n644) );
  XOR U825 ( .A(n643), .B(n644), .Z(n646) );
  XNOR U826 ( .A(n645), .B(n646), .Z(n693) );
  XNOR U827 ( .A(n694), .B(n693), .Z(n696) );
  NANDN U828 ( .A(n605), .B(n604), .Z(n609) );
  NANDN U829 ( .A(n607), .B(n606), .Z(n608) );
  AND U830 ( .A(n609), .B(n608), .Z(n640) );
  NANDN U831 ( .A(n611), .B(n610), .Z(n615) );
  NANDN U832 ( .A(n613), .B(n612), .Z(n614) );
  AND U833 ( .A(n615), .B(n614), .Z(n638) );
  XNOR U834 ( .A(n638), .B(n637), .Z(n639) );
  XNOR U835 ( .A(n640), .B(n639), .Z(n695) );
  XOR U836 ( .A(n696), .B(n695), .Z(n632) );
  NANDN U837 ( .A(n621), .B(n620), .Z(n625) );
  OR U838 ( .A(n623), .B(n622), .Z(n624) );
  AND U839 ( .A(n625), .B(n624), .Z(n631) );
  XNOR U840 ( .A(n632), .B(n631), .Z(n633) );
  XNOR U841 ( .A(n634), .B(n633), .Z(n626) );
  XNOR U842 ( .A(sreg[63]), .B(n626), .Z(n627) );
  XNOR U843 ( .A(n628), .B(n627), .Z(c[63]) );
  NANDN U844 ( .A(sreg[63]), .B(n626), .Z(n630) );
  NAND U845 ( .A(n628), .B(n627), .Z(n629) );
  NAND U846 ( .A(n630), .B(n629), .Z(n771) );
  XNOR U847 ( .A(sreg[64]), .B(n771), .Z(n773) );
  NANDN U848 ( .A(n632), .B(n631), .Z(n636) );
  NANDN U849 ( .A(n634), .B(n633), .Z(n635) );
  AND U850 ( .A(n636), .B(n635), .Z(n701) );
  NANDN U851 ( .A(n638), .B(n637), .Z(n642) );
  NANDN U852 ( .A(n640), .B(n639), .Z(n641) );
  AND U853 ( .A(n642), .B(n641), .Z(n767) );
  NANDN U854 ( .A(n644), .B(n643), .Z(n648) );
  OR U855 ( .A(n646), .B(n645), .Z(n647) );
  AND U856 ( .A(n648), .B(n647), .Z(n765) );
  NANDN U857 ( .A(n650), .B(n649), .Z(n654) );
  NANDN U858 ( .A(n652), .B(n651), .Z(n653) );
  AND U859 ( .A(n654), .B(n653), .Z(n760) );
  NAND U860 ( .A(b[0]), .B(a[16]), .Z(n655) );
  XNOR U861 ( .A(b[1]), .B(n655), .Z(n657) );
  NANDN U862 ( .A(b[0]), .B(a[15]), .Z(n656) );
  NAND U863 ( .A(n657), .B(n656), .Z(n729) );
  NAND U864 ( .A(n5012), .B(n658), .Z(n660) );
  XOR U865 ( .A(b[13]), .B(a[4]), .Z(n735) );
  NAND U866 ( .A(n4985), .B(n735), .Z(n659) );
  AND U867 ( .A(n660), .B(n659), .Z(n727) );
  AND U868 ( .A(b[15]), .B(a[0]), .Z(n726) );
  XOR U869 ( .A(n727), .B(n726), .Z(n728) );
  XNOR U870 ( .A(n729), .B(n728), .Z(n759) );
  XNOR U871 ( .A(n760), .B(n759), .Z(n762) );
  NANDN U872 ( .A(n662), .B(n661), .Z(n666) );
  NANDN U873 ( .A(n664), .B(n663), .Z(n665) );
  AND U874 ( .A(n666), .B(n665), .Z(n761) );
  XOR U875 ( .A(n762), .B(n761), .Z(n756) );
  NANDN U876 ( .A(n668), .B(n667), .Z(n672) );
  NAND U877 ( .A(n670), .B(n669), .Z(n671) );
  AND U878 ( .A(n672), .B(n671), .Z(n754) );
  NOR U879 ( .A(n674), .B(n673), .Z(n707) );
  NANDN U880 ( .A(n34), .B(n675), .Z(n677) );
  XNOR U881 ( .A(b[3]), .B(a[14]), .Z(n744) );
  OR U882 ( .A(n744), .B(n29), .Z(n676) );
  AND U883 ( .A(n677), .B(n676), .Z(n705) );
  OR U884 ( .A(n678), .B(n32), .Z(n680) );
  XNOR U885 ( .A(b[9]), .B(a[8]), .Z(n717) );
  OR U886 ( .A(n717), .B(n39), .Z(n679) );
  NAND U887 ( .A(n680), .B(n679), .Z(n706) );
  XOR U888 ( .A(n705), .B(n706), .Z(n708) );
  XOR U889 ( .A(n707), .B(n708), .Z(n750) );
  NAND U890 ( .A(n4755), .B(n681), .Z(n683) );
  XOR U891 ( .A(b[7]), .B(a[10]), .Z(n741) );
  NAND U892 ( .A(n4708), .B(n741), .Z(n682) );
  AND U893 ( .A(n683), .B(n682), .Z(n748) );
  NAND U894 ( .A(n4950), .B(n684), .Z(n686) );
  XOR U895 ( .A(b[11]), .B(a[6]), .Z(n711) );
  NAND U896 ( .A(n4863), .B(n711), .Z(n685) );
  AND U897 ( .A(n686), .B(n685), .Z(n723) );
  NAND U898 ( .A(n42), .B(n687), .Z(n689) );
  XOR U899 ( .A(b[15]), .B(a[2]), .Z(n714) );
  NAND U900 ( .A(n4981), .B(n714), .Z(n688) );
  AND U901 ( .A(n689), .B(n688), .Z(n721) );
  NAND U902 ( .A(n36), .B(n690), .Z(n692) );
  XOR U903 ( .A(b[5]), .B(a[12]), .Z(n738) );
  NAND U904 ( .A(n4560), .B(n738), .Z(n691) );
  NAND U905 ( .A(n692), .B(n691), .Z(n720) );
  XNOR U906 ( .A(n721), .B(n720), .Z(n722) );
  XNOR U907 ( .A(n723), .B(n722), .Z(n747) );
  XNOR U908 ( .A(n748), .B(n747), .Z(n749) );
  XNOR U909 ( .A(n750), .B(n749), .Z(n753) );
  XNOR U910 ( .A(n754), .B(n753), .Z(n755) );
  XOR U911 ( .A(n756), .B(n755), .Z(n766) );
  XOR U912 ( .A(n765), .B(n766), .Z(n768) );
  XOR U913 ( .A(n767), .B(n768), .Z(n700) );
  NANDN U914 ( .A(n694), .B(n693), .Z(n698) );
  NAND U915 ( .A(n696), .B(n695), .Z(n697) );
  AND U916 ( .A(n698), .B(n697), .Z(n699) );
  XOR U917 ( .A(n700), .B(n699), .Z(n702) );
  XNOR U918 ( .A(n701), .B(n702), .Z(n772) );
  XOR U919 ( .A(n773), .B(n772), .Z(c[64]) );
  NANDN U920 ( .A(n700), .B(n699), .Z(n704) );
  OR U921 ( .A(n702), .B(n701), .Z(n703) );
  AND U922 ( .A(n704), .B(n703), .Z(n783) );
  NANDN U923 ( .A(n706), .B(n705), .Z(n710) );
  OR U924 ( .A(n708), .B(n707), .Z(n709) );
  AND U925 ( .A(n710), .B(n709), .Z(n842) );
  NAND U926 ( .A(n4950), .B(n711), .Z(n713) );
  XOR U927 ( .A(b[11]), .B(a[7]), .Z(n820) );
  NAND U928 ( .A(n4863), .B(n820), .Z(n712) );
  AND U929 ( .A(n713), .B(n712), .Z(n831) );
  NAND U930 ( .A(n42), .B(n714), .Z(n716) );
  XOR U931 ( .A(b[15]), .B(a[3]), .Z(n823) );
  NAND U932 ( .A(n4981), .B(n823), .Z(n715) );
  AND U933 ( .A(n716), .B(n715), .Z(n830) );
  OR U934 ( .A(n717), .B(n32), .Z(n719) );
  XOR U935 ( .A(b[9]), .B(a[9]), .Z(n826) );
  NAND U936 ( .A(n4810), .B(n826), .Z(n718) );
  NAND U937 ( .A(n719), .B(n718), .Z(n829) );
  XOR U938 ( .A(n830), .B(n829), .Z(n832) );
  XNOR U939 ( .A(n831), .B(n832), .Z(n841) );
  XNOR U940 ( .A(n842), .B(n841), .Z(n843) );
  NANDN U941 ( .A(n721), .B(n720), .Z(n725) );
  NANDN U942 ( .A(n723), .B(n722), .Z(n724) );
  NAND U943 ( .A(n725), .B(n724), .Z(n844) );
  XNOR U944 ( .A(n843), .B(n844), .Z(n790) );
  NANDN U945 ( .A(n727), .B(n726), .Z(n731) );
  OR U946 ( .A(n729), .B(n728), .Z(n730) );
  AND U947 ( .A(n731), .B(n730), .Z(n816) );
  NAND U948 ( .A(b[0]), .B(a[17]), .Z(n732) );
  XNOR U949 ( .A(b[1]), .B(n732), .Z(n734) );
  NANDN U950 ( .A(b[0]), .B(a[16]), .Z(n733) );
  NAND U951 ( .A(n734), .B(n733), .Z(n796) );
  NAND U952 ( .A(n5012), .B(n735), .Z(n737) );
  XOR U953 ( .A(b[13]), .B(a[5]), .Z(n802) );
  NAND U954 ( .A(n4985), .B(n802), .Z(n736) );
  AND U955 ( .A(n737), .B(n736), .Z(n794) );
  AND U956 ( .A(b[15]), .B(a[1]), .Z(n793) );
  XNOR U957 ( .A(n794), .B(n793), .Z(n795) );
  XNOR U958 ( .A(n796), .B(n795), .Z(n814) );
  NAND U959 ( .A(n36), .B(n738), .Z(n740) );
  XOR U960 ( .A(b[5]), .B(a[13]), .Z(n805) );
  NAND U961 ( .A(n4560), .B(n805), .Z(n739) );
  AND U962 ( .A(n740), .B(n739), .Z(n838) );
  NAND U963 ( .A(n4755), .B(n741), .Z(n743) );
  XOR U964 ( .A(b[7]), .B(a[11]), .Z(n808) );
  NAND U965 ( .A(n4708), .B(n808), .Z(n742) );
  AND U966 ( .A(n743), .B(n742), .Z(n836) );
  OR U967 ( .A(n744), .B(n34), .Z(n746) );
  XOR U968 ( .A(b[3]), .B(a[15]), .Z(n811) );
  NAND U969 ( .A(n33), .B(n811), .Z(n745) );
  NAND U970 ( .A(n746), .B(n745), .Z(n835) );
  XNOR U971 ( .A(n836), .B(n835), .Z(n837) );
  XOR U972 ( .A(n838), .B(n837), .Z(n815) );
  XOR U973 ( .A(n814), .B(n815), .Z(n817) );
  XOR U974 ( .A(n816), .B(n817), .Z(n788) );
  NANDN U975 ( .A(n748), .B(n747), .Z(n752) );
  NANDN U976 ( .A(n750), .B(n749), .Z(n751) );
  AND U977 ( .A(n752), .B(n751), .Z(n787) );
  XNOR U978 ( .A(n788), .B(n787), .Z(n789) );
  XOR U979 ( .A(n790), .B(n789), .Z(n849) );
  NANDN U980 ( .A(n754), .B(n753), .Z(n758) );
  NANDN U981 ( .A(n756), .B(n755), .Z(n757) );
  AND U982 ( .A(n758), .B(n757), .Z(n848) );
  NANDN U983 ( .A(n760), .B(n759), .Z(n764) );
  NAND U984 ( .A(n762), .B(n761), .Z(n763) );
  AND U985 ( .A(n764), .B(n763), .Z(n847) );
  XOR U986 ( .A(n848), .B(n847), .Z(n850) );
  XOR U987 ( .A(n849), .B(n850), .Z(n782) );
  NANDN U988 ( .A(n766), .B(n765), .Z(n770) );
  OR U989 ( .A(n768), .B(n767), .Z(n769) );
  AND U990 ( .A(n770), .B(n769), .Z(n781) );
  XOR U991 ( .A(n782), .B(n781), .Z(n784) );
  XOR U992 ( .A(n783), .B(n784), .Z(n776) );
  XNOR U993 ( .A(n776), .B(sreg[65]), .Z(n778) );
  NANDN U994 ( .A(n771), .B(sreg[64]), .Z(n775) );
  NAND U995 ( .A(n773), .B(n772), .Z(n774) );
  NAND U996 ( .A(n775), .B(n774), .Z(n777) );
  XOR U997 ( .A(n778), .B(n777), .Z(c[65]) );
  NANDN U998 ( .A(n776), .B(sreg[65]), .Z(n780) );
  NAND U999 ( .A(n778), .B(n777), .Z(n779) );
  AND U1000 ( .A(n780), .B(n779), .Z(n927) );
  NANDN U1001 ( .A(n782), .B(n781), .Z(n786) );
  OR U1002 ( .A(n784), .B(n783), .Z(n785) );
  AND U1003 ( .A(n786), .B(n785), .Z(n856) );
  NANDN U1004 ( .A(n788), .B(n787), .Z(n792) );
  NAND U1005 ( .A(n790), .B(n789), .Z(n791) );
  AND U1006 ( .A(n792), .B(n791), .Z(n922) );
  NANDN U1007 ( .A(n794), .B(n793), .Z(n798) );
  NANDN U1008 ( .A(n796), .B(n795), .Z(n797) );
  AND U1009 ( .A(n798), .B(n797), .Z(n888) );
  NAND U1010 ( .A(b[0]), .B(a[18]), .Z(n799) );
  XNOR U1011 ( .A(b[1]), .B(n799), .Z(n801) );
  NANDN U1012 ( .A(b[0]), .B(a[17]), .Z(n800) );
  NAND U1013 ( .A(n801), .B(n800), .Z(n868) );
  NAND U1014 ( .A(n5012), .B(n802), .Z(n804) );
  XOR U1015 ( .A(b[13]), .B(a[6]), .Z(n874) );
  NAND U1016 ( .A(n4985), .B(n874), .Z(n803) );
  AND U1017 ( .A(n804), .B(n803), .Z(n866) );
  AND U1018 ( .A(b[15]), .B(a[2]), .Z(n865) );
  XNOR U1019 ( .A(n866), .B(n865), .Z(n867) );
  XNOR U1020 ( .A(n868), .B(n867), .Z(n886) );
  NAND U1021 ( .A(n36), .B(n805), .Z(n807) );
  XOR U1022 ( .A(b[5]), .B(a[14]), .Z(n877) );
  NAND U1023 ( .A(n4560), .B(n877), .Z(n806) );
  AND U1024 ( .A(n807), .B(n806), .Z(n910) );
  NAND U1025 ( .A(n4755), .B(n808), .Z(n810) );
  XOR U1026 ( .A(b[7]), .B(a[12]), .Z(n880) );
  NAND U1027 ( .A(n4708), .B(n880), .Z(n809) );
  AND U1028 ( .A(n810), .B(n809), .Z(n908) );
  NAND U1029 ( .A(n4471), .B(n811), .Z(n813) );
  XOR U1030 ( .A(b[3]), .B(a[16]), .Z(n883) );
  NAND U1031 ( .A(n33), .B(n883), .Z(n812) );
  NAND U1032 ( .A(n813), .B(n812), .Z(n907) );
  XNOR U1033 ( .A(n908), .B(n907), .Z(n909) );
  XOR U1034 ( .A(n910), .B(n909), .Z(n887) );
  XOR U1035 ( .A(n886), .B(n887), .Z(n889) );
  XOR U1036 ( .A(n888), .B(n889), .Z(n860) );
  NANDN U1037 ( .A(n815), .B(n814), .Z(n819) );
  OR U1038 ( .A(n817), .B(n816), .Z(n818) );
  AND U1039 ( .A(n819), .B(n818), .Z(n859) );
  XNOR U1040 ( .A(n860), .B(n859), .Z(n862) );
  NAND U1041 ( .A(n4950), .B(n820), .Z(n822) );
  XOR U1042 ( .A(b[11]), .B(a[8]), .Z(n892) );
  NAND U1043 ( .A(n4863), .B(n892), .Z(n821) );
  AND U1044 ( .A(n822), .B(n821), .Z(n903) );
  NAND U1045 ( .A(n42), .B(n823), .Z(n825) );
  XOR U1046 ( .A(b[15]), .B(a[4]), .Z(n895) );
  NAND U1047 ( .A(n4981), .B(n895), .Z(n824) );
  AND U1048 ( .A(n825), .B(n824), .Z(n902) );
  NAND U1049 ( .A(n41), .B(n826), .Z(n828) );
  XOR U1050 ( .A(b[9]), .B(a[10]), .Z(n898) );
  NAND U1051 ( .A(n4810), .B(n898), .Z(n827) );
  NAND U1052 ( .A(n828), .B(n827), .Z(n901) );
  XOR U1053 ( .A(n902), .B(n901), .Z(n904) );
  XOR U1054 ( .A(n903), .B(n904), .Z(n914) );
  NANDN U1055 ( .A(n830), .B(n829), .Z(n834) );
  OR U1056 ( .A(n832), .B(n831), .Z(n833) );
  AND U1057 ( .A(n834), .B(n833), .Z(n913) );
  XNOR U1058 ( .A(n914), .B(n913), .Z(n915) );
  NANDN U1059 ( .A(n836), .B(n835), .Z(n840) );
  NANDN U1060 ( .A(n838), .B(n837), .Z(n839) );
  NAND U1061 ( .A(n840), .B(n839), .Z(n916) );
  XNOR U1062 ( .A(n915), .B(n916), .Z(n861) );
  XOR U1063 ( .A(n862), .B(n861), .Z(n920) );
  NANDN U1064 ( .A(n842), .B(n841), .Z(n846) );
  NANDN U1065 ( .A(n844), .B(n843), .Z(n845) );
  AND U1066 ( .A(n846), .B(n845), .Z(n919) );
  XNOR U1067 ( .A(n920), .B(n919), .Z(n921) );
  XOR U1068 ( .A(n922), .B(n921), .Z(n854) );
  NANDN U1069 ( .A(n848), .B(n847), .Z(n852) );
  OR U1070 ( .A(n850), .B(n849), .Z(n851) );
  AND U1071 ( .A(n852), .B(n851), .Z(n853) );
  XNOR U1072 ( .A(n854), .B(n853), .Z(n855) );
  XNOR U1073 ( .A(n856), .B(n855), .Z(n925) );
  XNOR U1074 ( .A(sreg[66]), .B(n925), .Z(n926) );
  XNOR U1075 ( .A(n927), .B(n926), .Z(c[66]) );
  NANDN U1076 ( .A(n854), .B(n853), .Z(n858) );
  NANDN U1077 ( .A(n856), .B(n855), .Z(n857) );
  AND U1078 ( .A(n858), .B(n857), .Z(n933) );
  NANDN U1079 ( .A(n860), .B(n859), .Z(n864) );
  NAND U1080 ( .A(n862), .B(n861), .Z(n863) );
  AND U1081 ( .A(n864), .B(n863), .Z(n999) );
  NANDN U1082 ( .A(n866), .B(n865), .Z(n870) );
  NANDN U1083 ( .A(n868), .B(n867), .Z(n869) );
  AND U1084 ( .A(n870), .B(n869), .Z(n965) );
  NAND U1085 ( .A(b[0]), .B(a[19]), .Z(n871) );
  XNOR U1086 ( .A(b[1]), .B(n871), .Z(n873) );
  NANDN U1087 ( .A(b[0]), .B(a[18]), .Z(n872) );
  NAND U1088 ( .A(n873), .B(n872), .Z(n945) );
  NAND U1089 ( .A(n5012), .B(n874), .Z(n876) );
  XOR U1090 ( .A(b[13]), .B(a[7]), .Z(n951) );
  NAND U1091 ( .A(n4985), .B(n951), .Z(n875) );
  AND U1092 ( .A(n876), .B(n875), .Z(n943) );
  AND U1093 ( .A(b[15]), .B(a[3]), .Z(n942) );
  XNOR U1094 ( .A(n943), .B(n942), .Z(n944) );
  XNOR U1095 ( .A(n945), .B(n944), .Z(n963) );
  NAND U1096 ( .A(n36), .B(n877), .Z(n879) );
  XOR U1097 ( .A(b[5]), .B(a[15]), .Z(n954) );
  NAND U1098 ( .A(n4560), .B(n954), .Z(n878) );
  AND U1099 ( .A(n879), .B(n878), .Z(n987) );
  NAND U1100 ( .A(n4755), .B(n880), .Z(n882) );
  XOR U1101 ( .A(b[7]), .B(a[13]), .Z(n957) );
  NAND U1102 ( .A(n4708), .B(n957), .Z(n881) );
  AND U1103 ( .A(n882), .B(n881), .Z(n985) );
  NAND U1104 ( .A(n4471), .B(n883), .Z(n885) );
  XOR U1105 ( .A(b[3]), .B(a[17]), .Z(n960) );
  NAND U1106 ( .A(n33), .B(n960), .Z(n884) );
  NAND U1107 ( .A(n885), .B(n884), .Z(n984) );
  XNOR U1108 ( .A(n985), .B(n984), .Z(n986) );
  XOR U1109 ( .A(n987), .B(n986), .Z(n964) );
  XOR U1110 ( .A(n963), .B(n964), .Z(n966) );
  XOR U1111 ( .A(n965), .B(n966), .Z(n937) );
  NANDN U1112 ( .A(n887), .B(n886), .Z(n891) );
  OR U1113 ( .A(n889), .B(n888), .Z(n890) );
  AND U1114 ( .A(n891), .B(n890), .Z(n936) );
  XNOR U1115 ( .A(n937), .B(n936), .Z(n939) );
  NAND U1116 ( .A(n4950), .B(n892), .Z(n894) );
  XOR U1117 ( .A(b[11]), .B(a[9]), .Z(n969) );
  NAND U1118 ( .A(n4863), .B(n969), .Z(n893) );
  AND U1119 ( .A(n894), .B(n893), .Z(n980) );
  NAND U1120 ( .A(n42), .B(n895), .Z(n897) );
  XOR U1121 ( .A(b[15]), .B(a[5]), .Z(n972) );
  NAND U1122 ( .A(n4981), .B(n972), .Z(n896) );
  AND U1123 ( .A(n897), .B(n896), .Z(n979) );
  NAND U1124 ( .A(n41), .B(n898), .Z(n900) );
  XOR U1125 ( .A(b[9]), .B(a[11]), .Z(n975) );
  NAND U1126 ( .A(n4810), .B(n975), .Z(n899) );
  NAND U1127 ( .A(n900), .B(n899), .Z(n978) );
  XOR U1128 ( .A(n979), .B(n978), .Z(n981) );
  XOR U1129 ( .A(n980), .B(n981), .Z(n991) );
  NANDN U1130 ( .A(n902), .B(n901), .Z(n906) );
  OR U1131 ( .A(n904), .B(n903), .Z(n905) );
  AND U1132 ( .A(n906), .B(n905), .Z(n990) );
  XNOR U1133 ( .A(n991), .B(n990), .Z(n992) );
  NANDN U1134 ( .A(n908), .B(n907), .Z(n912) );
  NANDN U1135 ( .A(n910), .B(n909), .Z(n911) );
  NAND U1136 ( .A(n912), .B(n911), .Z(n993) );
  XNOR U1137 ( .A(n992), .B(n993), .Z(n938) );
  XOR U1138 ( .A(n939), .B(n938), .Z(n997) );
  NANDN U1139 ( .A(n914), .B(n913), .Z(n918) );
  NANDN U1140 ( .A(n916), .B(n915), .Z(n917) );
  AND U1141 ( .A(n918), .B(n917), .Z(n996) );
  XNOR U1142 ( .A(n997), .B(n996), .Z(n998) );
  XOR U1143 ( .A(n999), .B(n998), .Z(n931) );
  NANDN U1144 ( .A(n920), .B(n919), .Z(n924) );
  NAND U1145 ( .A(n922), .B(n921), .Z(n923) );
  AND U1146 ( .A(n924), .B(n923), .Z(n930) );
  XNOR U1147 ( .A(n931), .B(n930), .Z(n932) );
  XNOR U1148 ( .A(n933), .B(n932), .Z(n1002) );
  XNOR U1149 ( .A(sreg[67]), .B(n1002), .Z(n1004) );
  NANDN U1150 ( .A(sreg[66]), .B(n925), .Z(n929) );
  NAND U1151 ( .A(n927), .B(n926), .Z(n928) );
  NAND U1152 ( .A(n929), .B(n928), .Z(n1003) );
  XNOR U1153 ( .A(n1004), .B(n1003), .Z(c[67]) );
  NANDN U1154 ( .A(n931), .B(n930), .Z(n935) );
  NANDN U1155 ( .A(n933), .B(n932), .Z(n934) );
  AND U1156 ( .A(n935), .B(n934), .Z(n1014) );
  NANDN U1157 ( .A(n937), .B(n936), .Z(n941) );
  NAND U1158 ( .A(n939), .B(n938), .Z(n940) );
  AND U1159 ( .A(n941), .B(n940), .Z(n1081) );
  NANDN U1160 ( .A(n943), .B(n942), .Z(n947) );
  NANDN U1161 ( .A(n945), .B(n944), .Z(n946) );
  AND U1162 ( .A(n947), .B(n946), .Z(n1068) );
  NAND U1163 ( .A(b[0]), .B(a[20]), .Z(n948) );
  XNOR U1164 ( .A(b[1]), .B(n948), .Z(n950) );
  NANDN U1165 ( .A(b[0]), .B(a[19]), .Z(n949) );
  NAND U1166 ( .A(n950), .B(n949), .Z(n1048) );
  NAND U1167 ( .A(n5012), .B(n951), .Z(n953) );
  XOR U1168 ( .A(b[13]), .B(a[8]), .Z(n1054) );
  NAND U1169 ( .A(n4985), .B(n1054), .Z(n952) );
  AND U1170 ( .A(n953), .B(n952), .Z(n1046) );
  AND U1171 ( .A(b[15]), .B(a[4]), .Z(n1045) );
  XNOR U1172 ( .A(n1046), .B(n1045), .Z(n1047) );
  XNOR U1173 ( .A(n1048), .B(n1047), .Z(n1066) );
  NAND U1174 ( .A(n36), .B(n954), .Z(n956) );
  XOR U1175 ( .A(b[5]), .B(a[16]), .Z(n1057) );
  NAND U1176 ( .A(n4560), .B(n1057), .Z(n955) );
  AND U1177 ( .A(n956), .B(n955), .Z(n1042) );
  NAND U1178 ( .A(n4755), .B(n957), .Z(n959) );
  XOR U1179 ( .A(b[7]), .B(a[14]), .Z(n1060) );
  NAND U1180 ( .A(n4708), .B(n1060), .Z(n958) );
  AND U1181 ( .A(n959), .B(n958), .Z(n1040) );
  NAND U1182 ( .A(n4471), .B(n960), .Z(n962) );
  XOR U1183 ( .A(b[3]), .B(a[18]), .Z(n1063) );
  NAND U1184 ( .A(n33), .B(n1063), .Z(n961) );
  NAND U1185 ( .A(n962), .B(n961), .Z(n1039) );
  XNOR U1186 ( .A(n1040), .B(n1039), .Z(n1041) );
  XOR U1187 ( .A(n1042), .B(n1041), .Z(n1067) );
  XOR U1188 ( .A(n1066), .B(n1067), .Z(n1069) );
  XOR U1189 ( .A(n1068), .B(n1069), .Z(n1019) );
  NANDN U1190 ( .A(n964), .B(n963), .Z(n968) );
  OR U1191 ( .A(n966), .B(n965), .Z(n967) );
  AND U1192 ( .A(n968), .B(n967), .Z(n1018) );
  XNOR U1193 ( .A(n1019), .B(n1018), .Z(n1021) );
  NAND U1194 ( .A(n4950), .B(n969), .Z(n971) );
  XOR U1195 ( .A(b[11]), .B(a[10]), .Z(n1024) );
  NAND U1196 ( .A(n4863), .B(n1024), .Z(n970) );
  AND U1197 ( .A(n971), .B(n970), .Z(n1035) );
  NAND U1198 ( .A(n42), .B(n972), .Z(n974) );
  XOR U1199 ( .A(b[15]), .B(a[6]), .Z(n1027) );
  NAND U1200 ( .A(n4981), .B(n1027), .Z(n973) );
  AND U1201 ( .A(n974), .B(n973), .Z(n1034) );
  NAND U1202 ( .A(n41), .B(n975), .Z(n977) );
  XOR U1203 ( .A(b[9]), .B(a[12]), .Z(n1030) );
  NAND U1204 ( .A(n4810), .B(n1030), .Z(n976) );
  NAND U1205 ( .A(n977), .B(n976), .Z(n1033) );
  XOR U1206 ( .A(n1034), .B(n1033), .Z(n1036) );
  XOR U1207 ( .A(n1035), .B(n1036), .Z(n1073) );
  NANDN U1208 ( .A(n979), .B(n978), .Z(n983) );
  OR U1209 ( .A(n981), .B(n980), .Z(n982) );
  AND U1210 ( .A(n983), .B(n982), .Z(n1072) );
  XNOR U1211 ( .A(n1073), .B(n1072), .Z(n1074) );
  NANDN U1212 ( .A(n985), .B(n984), .Z(n989) );
  NANDN U1213 ( .A(n987), .B(n986), .Z(n988) );
  NAND U1214 ( .A(n989), .B(n988), .Z(n1075) );
  XNOR U1215 ( .A(n1074), .B(n1075), .Z(n1020) );
  XOR U1216 ( .A(n1021), .B(n1020), .Z(n1079) );
  NANDN U1217 ( .A(n991), .B(n990), .Z(n995) );
  NANDN U1218 ( .A(n993), .B(n992), .Z(n994) );
  AND U1219 ( .A(n995), .B(n994), .Z(n1078) );
  XNOR U1220 ( .A(n1079), .B(n1078), .Z(n1080) );
  XOR U1221 ( .A(n1081), .B(n1080), .Z(n1013) );
  NANDN U1222 ( .A(n997), .B(n996), .Z(n1001) );
  NAND U1223 ( .A(n999), .B(n998), .Z(n1000) );
  AND U1224 ( .A(n1001), .B(n1000), .Z(n1012) );
  XOR U1225 ( .A(n1013), .B(n1012), .Z(n1015) );
  XOR U1226 ( .A(n1014), .B(n1015), .Z(n1007) );
  XNOR U1227 ( .A(n1007), .B(sreg[68]), .Z(n1009) );
  NANDN U1228 ( .A(sreg[67]), .B(n1002), .Z(n1006) );
  NAND U1229 ( .A(n1004), .B(n1003), .Z(n1005) );
  AND U1230 ( .A(n1006), .B(n1005), .Z(n1008) );
  XOR U1231 ( .A(n1009), .B(n1008), .Z(c[68]) );
  NANDN U1232 ( .A(n1007), .B(sreg[68]), .Z(n1011) );
  NAND U1233 ( .A(n1009), .B(n1008), .Z(n1010) );
  AND U1234 ( .A(n1011), .B(n1010), .Z(n1158) );
  NANDN U1235 ( .A(n1013), .B(n1012), .Z(n1017) );
  OR U1236 ( .A(n1015), .B(n1014), .Z(n1016) );
  AND U1237 ( .A(n1017), .B(n1016), .Z(n1087) );
  NANDN U1238 ( .A(n1019), .B(n1018), .Z(n1023) );
  NAND U1239 ( .A(n1021), .B(n1020), .Z(n1022) );
  AND U1240 ( .A(n1023), .B(n1022), .Z(n1153) );
  NAND U1241 ( .A(n4950), .B(n1024), .Z(n1026) );
  XOR U1242 ( .A(b[11]), .B(a[11]), .Z(n1123) );
  NAND U1243 ( .A(n4863), .B(n1123), .Z(n1025) );
  AND U1244 ( .A(n1026), .B(n1025), .Z(n1134) );
  NAND U1245 ( .A(n42), .B(n1027), .Z(n1029) );
  XOR U1246 ( .A(b[15]), .B(a[7]), .Z(n1126) );
  NAND U1247 ( .A(n4981), .B(n1126), .Z(n1028) );
  AND U1248 ( .A(n1029), .B(n1028), .Z(n1133) );
  NAND U1249 ( .A(n41), .B(n1030), .Z(n1032) );
  XOR U1250 ( .A(b[9]), .B(a[13]), .Z(n1129) );
  NAND U1251 ( .A(n4810), .B(n1129), .Z(n1031) );
  NAND U1252 ( .A(n1032), .B(n1031), .Z(n1132) );
  XOR U1253 ( .A(n1133), .B(n1132), .Z(n1135) );
  XOR U1254 ( .A(n1134), .B(n1135), .Z(n1145) );
  NANDN U1255 ( .A(n1034), .B(n1033), .Z(n1038) );
  OR U1256 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1257 ( .A(n1038), .B(n1037), .Z(n1144) );
  XNOR U1258 ( .A(n1145), .B(n1144), .Z(n1146) );
  NANDN U1259 ( .A(n1040), .B(n1039), .Z(n1044) );
  NANDN U1260 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1261 ( .A(n1044), .B(n1043), .Z(n1147) );
  XNOR U1262 ( .A(n1146), .B(n1147), .Z(n1093) );
  NANDN U1263 ( .A(n1046), .B(n1045), .Z(n1050) );
  NANDN U1264 ( .A(n1048), .B(n1047), .Z(n1049) );
  AND U1265 ( .A(n1050), .B(n1049), .Z(n1119) );
  NAND U1266 ( .A(b[0]), .B(a[21]), .Z(n1051) );
  XNOR U1267 ( .A(b[1]), .B(n1051), .Z(n1053) );
  NANDN U1268 ( .A(b[0]), .B(a[20]), .Z(n1052) );
  NAND U1269 ( .A(n1053), .B(n1052), .Z(n1099) );
  NAND U1270 ( .A(n5012), .B(n1054), .Z(n1056) );
  XOR U1271 ( .A(b[13]), .B(a[9]), .Z(n1102) );
  NAND U1272 ( .A(n4985), .B(n1102), .Z(n1055) );
  AND U1273 ( .A(n1056), .B(n1055), .Z(n1097) );
  AND U1274 ( .A(b[15]), .B(a[5]), .Z(n1096) );
  XNOR U1275 ( .A(n1097), .B(n1096), .Z(n1098) );
  XNOR U1276 ( .A(n1099), .B(n1098), .Z(n1117) );
  NAND U1277 ( .A(n36), .B(n1057), .Z(n1059) );
  XOR U1278 ( .A(b[5]), .B(a[17]), .Z(n1108) );
  NAND U1279 ( .A(n4560), .B(n1108), .Z(n1058) );
  AND U1280 ( .A(n1059), .B(n1058), .Z(n1141) );
  NAND U1281 ( .A(n4755), .B(n1060), .Z(n1062) );
  XOR U1282 ( .A(b[7]), .B(a[15]), .Z(n1111) );
  NAND U1283 ( .A(n4708), .B(n1111), .Z(n1061) );
  AND U1284 ( .A(n1062), .B(n1061), .Z(n1139) );
  NAND U1285 ( .A(n4471), .B(n1063), .Z(n1065) );
  XOR U1286 ( .A(b[3]), .B(a[19]), .Z(n1114) );
  NAND U1287 ( .A(n33), .B(n1114), .Z(n1064) );
  NAND U1288 ( .A(n1065), .B(n1064), .Z(n1138) );
  XNOR U1289 ( .A(n1139), .B(n1138), .Z(n1140) );
  XOR U1290 ( .A(n1141), .B(n1140), .Z(n1118) );
  XOR U1291 ( .A(n1117), .B(n1118), .Z(n1120) );
  XOR U1292 ( .A(n1119), .B(n1120), .Z(n1091) );
  NANDN U1293 ( .A(n1067), .B(n1066), .Z(n1071) );
  OR U1294 ( .A(n1069), .B(n1068), .Z(n1070) );
  AND U1295 ( .A(n1071), .B(n1070), .Z(n1090) );
  XNOR U1296 ( .A(n1091), .B(n1090), .Z(n1092) );
  XOR U1297 ( .A(n1093), .B(n1092), .Z(n1151) );
  NANDN U1298 ( .A(n1073), .B(n1072), .Z(n1077) );
  NANDN U1299 ( .A(n1075), .B(n1074), .Z(n1076) );
  AND U1300 ( .A(n1077), .B(n1076), .Z(n1150) );
  XNOR U1301 ( .A(n1151), .B(n1150), .Z(n1152) );
  XOR U1302 ( .A(n1153), .B(n1152), .Z(n1085) );
  NANDN U1303 ( .A(n1079), .B(n1078), .Z(n1083) );
  NAND U1304 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1305 ( .A(n1083), .B(n1082), .Z(n1084) );
  XNOR U1306 ( .A(n1085), .B(n1084), .Z(n1086) );
  XNOR U1307 ( .A(n1087), .B(n1086), .Z(n1156) );
  XNOR U1308 ( .A(sreg[69]), .B(n1156), .Z(n1157) );
  XNOR U1309 ( .A(n1158), .B(n1157), .Z(c[69]) );
  NANDN U1310 ( .A(n1085), .B(n1084), .Z(n1089) );
  NANDN U1311 ( .A(n1087), .B(n1086), .Z(n1088) );
  AND U1312 ( .A(n1089), .B(n1088), .Z(n1164) );
  NANDN U1313 ( .A(n1091), .B(n1090), .Z(n1095) );
  NAND U1314 ( .A(n1093), .B(n1092), .Z(n1094) );
  AND U1315 ( .A(n1095), .B(n1094), .Z(n1230) );
  NANDN U1316 ( .A(n1097), .B(n1096), .Z(n1101) );
  NANDN U1317 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1318 ( .A(n1101), .B(n1100), .Z(n1196) );
  NAND U1319 ( .A(n5012), .B(n1102), .Z(n1104) );
  XOR U1320 ( .A(b[13]), .B(a[10]), .Z(n1182) );
  NAND U1321 ( .A(n4985), .B(n1182), .Z(n1103) );
  AND U1322 ( .A(n1104), .B(n1103), .Z(n1174) );
  AND U1323 ( .A(b[15]), .B(a[6]), .Z(n1173) );
  XNOR U1324 ( .A(n1174), .B(n1173), .Z(n1175) );
  NAND U1325 ( .A(b[0]), .B(a[22]), .Z(n1105) );
  XNOR U1326 ( .A(b[1]), .B(n1105), .Z(n1107) );
  NANDN U1327 ( .A(b[0]), .B(a[21]), .Z(n1106) );
  NAND U1328 ( .A(n1107), .B(n1106), .Z(n1176) );
  XNOR U1329 ( .A(n1175), .B(n1176), .Z(n1194) );
  NAND U1330 ( .A(n36), .B(n1108), .Z(n1110) );
  XOR U1331 ( .A(b[5]), .B(a[18]), .Z(n1185) );
  NAND U1332 ( .A(n4560), .B(n1185), .Z(n1109) );
  AND U1333 ( .A(n1110), .B(n1109), .Z(n1218) );
  NAND U1334 ( .A(n4755), .B(n1111), .Z(n1113) );
  XOR U1335 ( .A(b[7]), .B(a[16]), .Z(n1188) );
  NAND U1336 ( .A(n4708), .B(n1188), .Z(n1112) );
  AND U1337 ( .A(n1113), .B(n1112), .Z(n1216) );
  NAND U1338 ( .A(n4471), .B(n1114), .Z(n1116) );
  XOR U1339 ( .A(b[3]), .B(a[20]), .Z(n1191) );
  NAND U1340 ( .A(n33), .B(n1191), .Z(n1115) );
  NAND U1341 ( .A(n1116), .B(n1115), .Z(n1215) );
  XNOR U1342 ( .A(n1216), .B(n1215), .Z(n1217) );
  XOR U1343 ( .A(n1218), .B(n1217), .Z(n1195) );
  XOR U1344 ( .A(n1194), .B(n1195), .Z(n1197) );
  XOR U1345 ( .A(n1196), .B(n1197), .Z(n1168) );
  NANDN U1346 ( .A(n1118), .B(n1117), .Z(n1122) );
  OR U1347 ( .A(n1120), .B(n1119), .Z(n1121) );
  AND U1348 ( .A(n1122), .B(n1121), .Z(n1167) );
  XNOR U1349 ( .A(n1168), .B(n1167), .Z(n1170) );
  NAND U1350 ( .A(n4950), .B(n1123), .Z(n1125) );
  XOR U1351 ( .A(b[11]), .B(a[12]), .Z(n1200) );
  NAND U1352 ( .A(n4863), .B(n1200), .Z(n1124) );
  AND U1353 ( .A(n1125), .B(n1124), .Z(n1211) );
  NAND U1354 ( .A(n42), .B(n1126), .Z(n1128) );
  XOR U1355 ( .A(b[15]), .B(a[8]), .Z(n1203) );
  NAND U1356 ( .A(n4981), .B(n1203), .Z(n1127) );
  AND U1357 ( .A(n1128), .B(n1127), .Z(n1210) );
  NAND U1358 ( .A(n41), .B(n1129), .Z(n1131) );
  XOR U1359 ( .A(b[9]), .B(a[14]), .Z(n1206) );
  NAND U1360 ( .A(n4810), .B(n1206), .Z(n1130) );
  NAND U1361 ( .A(n1131), .B(n1130), .Z(n1209) );
  XOR U1362 ( .A(n1210), .B(n1209), .Z(n1212) );
  XOR U1363 ( .A(n1211), .B(n1212), .Z(n1222) );
  NANDN U1364 ( .A(n1133), .B(n1132), .Z(n1137) );
  OR U1365 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U1366 ( .A(n1137), .B(n1136), .Z(n1221) );
  XNOR U1367 ( .A(n1222), .B(n1221), .Z(n1223) );
  NANDN U1368 ( .A(n1139), .B(n1138), .Z(n1143) );
  NANDN U1369 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U1370 ( .A(n1143), .B(n1142), .Z(n1224) );
  XNOR U1371 ( .A(n1223), .B(n1224), .Z(n1169) );
  XOR U1372 ( .A(n1170), .B(n1169), .Z(n1228) );
  NANDN U1373 ( .A(n1145), .B(n1144), .Z(n1149) );
  NANDN U1374 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1375 ( .A(n1149), .B(n1148), .Z(n1227) );
  XNOR U1376 ( .A(n1228), .B(n1227), .Z(n1229) );
  XOR U1377 ( .A(n1230), .B(n1229), .Z(n1162) );
  NANDN U1378 ( .A(n1151), .B(n1150), .Z(n1155) );
  NAND U1379 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U1380 ( .A(n1155), .B(n1154), .Z(n1161) );
  XNOR U1381 ( .A(n1162), .B(n1161), .Z(n1163) );
  XNOR U1382 ( .A(n1164), .B(n1163), .Z(n1233) );
  XNOR U1383 ( .A(sreg[70]), .B(n1233), .Z(n1235) );
  NANDN U1384 ( .A(sreg[69]), .B(n1156), .Z(n1160) );
  NAND U1385 ( .A(n1158), .B(n1157), .Z(n1159) );
  NAND U1386 ( .A(n1160), .B(n1159), .Z(n1234) );
  XNOR U1387 ( .A(n1235), .B(n1234), .Z(c[70]) );
  NANDN U1388 ( .A(n1162), .B(n1161), .Z(n1166) );
  NANDN U1389 ( .A(n1164), .B(n1163), .Z(n1165) );
  AND U1390 ( .A(n1166), .B(n1165), .Z(n1245) );
  NANDN U1391 ( .A(n1168), .B(n1167), .Z(n1172) );
  NAND U1392 ( .A(n1170), .B(n1169), .Z(n1171) );
  AND U1393 ( .A(n1172), .B(n1171), .Z(n1312) );
  NANDN U1394 ( .A(n1174), .B(n1173), .Z(n1178) );
  NANDN U1395 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1396 ( .A(n1178), .B(n1177), .Z(n1278) );
  NAND U1397 ( .A(b[0]), .B(a[23]), .Z(n1179) );
  XNOR U1398 ( .A(b[1]), .B(n1179), .Z(n1181) );
  NANDN U1399 ( .A(b[0]), .B(a[22]), .Z(n1180) );
  NAND U1400 ( .A(n1181), .B(n1180), .Z(n1258) );
  NAND U1401 ( .A(n5012), .B(n1182), .Z(n1184) );
  XOR U1402 ( .A(b[13]), .B(a[11]), .Z(n1264) );
  NAND U1403 ( .A(n4985), .B(n1264), .Z(n1183) );
  AND U1404 ( .A(n1184), .B(n1183), .Z(n1256) );
  AND U1405 ( .A(b[15]), .B(a[7]), .Z(n1255) );
  XNOR U1406 ( .A(n1256), .B(n1255), .Z(n1257) );
  XNOR U1407 ( .A(n1258), .B(n1257), .Z(n1276) );
  NAND U1408 ( .A(n36), .B(n1185), .Z(n1187) );
  XOR U1409 ( .A(b[5]), .B(a[19]), .Z(n1267) );
  NAND U1410 ( .A(n4560), .B(n1267), .Z(n1186) );
  AND U1411 ( .A(n1187), .B(n1186), .Z(n1300) );
  NAND U1412 ( .A(n4755), .B(n1188), .Z(n1190) );
  XOR U1413 ( .A(b[7]), .B(a[17]), .Z(n1270) );
  NAND U1414 ( .A(n4708), .B(n1270), .Z(n1189) );
  AND U1415 ( .A(n1190), .B(n1189), .Z(n1298) );
  NAND U1416 ( .A(n4471), .B(n1191), .Z(n1193) );
  XOR U1417 ( .A(b[3]), .B(a[21]), .Z(n1273) );
  NAND U1418 ( .A(n33), .B(n1273), .Z(n1192) );
  NAND U1419 ( .A(n1193), .B(n1192), .Z(n1297) );
  XNOR U1420 ( .A(n1298), .B(n1297), .Z(n1299) );
  XOR U1421 ( .A(n1300), .B(n1299), .Z(n1277) );
  XOR U1422 ( .A(n1276), .B(n1277), .Z(n1279) );
  XOR U1423 ( .A(n1278), .B(n1279), .Z(n1250) );
  NANDN U1424 ( .A(n1195), .B(n1194), .Z(n1199) );
  OR U1425 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U1426 ( .A(n1199), .B(n1198), .Z(n1249) );
  XNOR U1427 ( .A(n1250), .B(n1249), .Z(n1252) );
  NAND U1428 ( .A(n4950), .B(n1200), .Z(n1202) );
  XOR U1429 ( .A(b[11]), .B(a[13]), .Z(n1282) );
  NAND U1430 ( .A(n4863), .B(n1282), .Z(n1201) );
  AND U1431 ( .A(n1202), .B(n1201), .Z(n1293) );
  NAND U1432 ( .A(n42), .B(n1203), .Z(n1205) );
  XOR U1433 ( .A(b[15]), .B(a[9]), .Z(n1285) );
  NAND U1434 ( .A(n4981), .B(n1285), .Z(n1204) );
  AND U1435 ( .A(n1205), .B(n1204), .Z(n1292) );
  NAND U1436 ( .A(n41), .B(n1206), .Z(n1208) );
  XOR U1437 ( .A(b[9]), .B(a[15]), .Z(n1288) );
  NAND U1438 ( .A(n4810), .B(n1288), .Z(n1207) );
  NAND U1439 ( .A(n1208), .B(n1207), .Z(n1291) );
  XOR U1440 ( .A(n1292), .B(n1291), .Z(n1294) );
  XOR U1441 ( .A(n1293), .B(n1294), .Z(n1304) );
  NANDN U1442 ( .A(n1210), .B(n1209), .Z(n1214) );
  OR U1443 ( .A(n1212), .B(n1211), .Z(n1213) );
  AND U1444 ( .A(n1214), .B(n1213), .Z(n1303) );
  XNOR U1445 ( .A(n1304), .B(n1303), .Z(n1305) );
  NANDN U1446 ( .A(n1216), .B(n1215), .Z(n1220) );
  NANDN U1447 ( .A(n1218), .B(n1217), .Z(n1219) );
  NAND U1448 ( .A(n1220), .B(n1219), .Z(n1306) );
  XNOR U1449 ( .A(n1305), .B(n1306), .Z(n1251) );
  XOR U1450 ( .A(n1252), .B(n1251), .Z(n1310) );
  NANDN U1451 ( .A(n1222), .B(n1221), .Z(n1226) );
  NANDN U1452 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1453 ( .A(n1226), .B(n1225), .Z(n1309) );
  XNOR U1454 ( .A(n1310), .B(n1309), .Z(n1311) );
  XOR U1455 ( .A(n1312), .B(n1311), .Z(n1244) );
  NANDN U1456 ( .A(n1228), .B(n1227), .Z(n1232) );
  NAND U1457 ( .A(n1230), .B(n1229), .Z(n1231) );
  AND U1458 ( .A(n1232), .B(n1231), .Z(n1243) );
  XOR U1459 ( .A(n1244), .B(n1243), .Z(n1246) );
  XOR U1460 ( .A(n1245), .B(n1246), .Z(n1238) );
  XNOR U1461 ( .A(n1238), .B(sreg[71]), .Z(n1240) );
  NANDN U1462 ( .A(sreg[70]), .B(n1233), .Z(n1237) );
  NAND U1463 ( .A(n1235), .B(n1234), .Z(n1236) );
  AND U1464 ( .A(n1237), .B(n1236), .Z(n1239) );
  XOR U1465 ( .A(n1240), .B(n1239), .Z(c[71]) );
  NANDN U1466 ( .A(n1238), .B(sreg[71]), .Z(n1242) );
  NAND U1467 ( .A(n1240), .B(n1239), .Z(n1241) );
  AND U1468 ( .A(n1242), .B(n1241), .Z(n1389) );
  NANDN U1469 ( .A(n1244), .B(n1243), .Z(n1248) );
  OR U1470 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U1471 ( .A(n1248), .B(n1247), .Z(n1318) );
  NANDN U1472 ( .A(n1250), .B(n1249), .Z(n1254) );
  NAND U1473 ( .A(n1252), .B(n1251), .Z(n1253) );
  AND U1474 ( .A(n1254), .B(n1253), .Z(n1384) );
  NANDN U1475 ( .A(n1256), .B(n1255), .Z(n1260) );
  NANDN U1476 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U1477 ( .A(n1260), .B(n1259), .Z(n1350) );
  NAND U1478 ( .A(b[0]), .B(a[24]), .Z(n1261) );
  XNOR U1479 ( .A(b[1]), .B(n1261), .Z(n1263) );
  NANDN U1480 ( .A(b[0]), .B(a[23]), .Z(n1262) );
  NAND U1481 ( .A(n1263), .B(n1262), .Z(n1330) );
  NAND U1482 ( .A(n5012), .B(n1264), .Z(n1266) );
  XOR U1483 ( .A(b[13]), .B(a[12]), .Z(n1336) );
  NAND U1484 ( .A(n4985), .B(n1336), .Z(n1265) );
  AND U1485 ( .A(n1266), .B(n1265), .Z(n1328) );
  AND U1486 ( .A(b[15]), .B(a[8]), .Z(n1327) );
  XNOR U1487 ( .A(n1328), .B(n1327), .Z(n1329) );
  XNOR U1488 ( .A(n1330), .B(n1329), .Z(n1348) );
  NAND U1489 ( .A(n36), .B(n1267), .Z(n1269) );
  XOR U1490 ( .A(b[5]), .B(a[20]), .Z(n1339) );
  NAND U1491 ( .A(n4560), .B(n1339), .Z(n1268) );
  AND U1492 ( .A(n1269), .B(n1268), .Z(n1372) );
  NAND U1493 ( .A(n4755), .B(n1270), .Z(n1272) );
  XOR U1494 ( .A(b[7]), .B(a[18]), .Z(n1342) );
  NAND U1495 ( .A(n4708), .B(n1342), .Z(n1271) );
  AND U1496 ( .A(n1272), .B(n1271), .Z(n1370) );
  NAND U1497 ( .A(n4471), .B(n1273), .Z(n1275) );
  XOR U1498 ( .A(b[3]), .B(a[22]), .Z(n1345) );
  NAND U1499 ( .A(n33), .B(n1345), .Z(n1274) );
  NAND U1500 ( .A(n1275), .B(n1274), .Z(n1369) );
  XNOR U1501 ( .A(n1370), .B(n1369), .Z(n1371) );
  XOR U1502 ( .A(n1372), .B(n1371), .Z(n1349) );
  XOR U1503 ( .A(n1348), .B(n1349), .Z(n1351) );
  XOR U1504 ( .A(n1350), .B(n1351), .Z(n1322) );
  NANDN U1505 ( .A(n1277), .B(n1276), .Z(n1281) );
  OR U1506 ( .A(n1279), .B(n1278), .Z(n1280) );
  AND U1507 ( .A(n1281), .B(n1280), .Z(n1321) );
  XNOR U1508 ( .A(n1322), .B(n1321), .Z(n1324) );
  NAND U1509 ( .A(n4950), .B(n1282), .Z(n1284) );
  XOR U1510 ( .A(b[11]), .B(a[14]), .Z(n1354) );
  NAND U1511 ( .A(n4863), .B(n1354), .Z(n1283) );
  AND U1512 ( .A(n1284), .B(n1283), .Z(n1365) );
  NAND U1513 ( .A(n42), .B(n1285), .Z(n1287) );
  XOR U1514 ( .A(b[15]), .B(a[10]), .Z(n1357) );
  NAND U1515 ( .A(n4981), .B(n1357), .Z(n1286) );
  AND U1516 ( .A(n1287), .B(n1286), .Z(n1364) );
  NAND U1517 ( .A(n41), .B(n1288), .Z(n1290) );
  XOR U1518 ( .A(b[9]), .B(a[16]), .Z(n1360) );
  NAND U1519 ( .A(n4810), .B(n1360), .Z(n1289) );
  NAND U1520 ( .A(n1290), .B(n1289), .Z(n1363) );
  XOR U1521 ( .A(n1364), .B(n1363), .Z(n1366) );
  XOR U1522 ( .A(n1365), .B(n1366), .Z(n1376) );
  NANDN U1523 ( .A(n1292), .B(n1291), .Z(n1296) );
  OR U1524 ( .A(n1294), .B(n1293), .Z(n1295) );
  AND U1525 ( .A(n1296), .B(n1295), .Z(n1375) );
  XNOR U1526 ( .A(n1376), .B(n1375), .Z(n1377) );
  NANDN U1527 ( .A(n1298), .B(n1297), .Z(n1302) );
  NANDN U1528 ( .A(n1300), .B(n1299), .Z(n1301) );
  NAND U1529 ( .A(n1302), .B(n1301), .Z(n1378) );
  XNOR U1530 ( .A(n1377), .B(n1378), .Z(n1323) );
  XOR U1531 ( .A(n1324), .B(n1323), .Z(n1382) );
  NANDN U1532 ( .A(n1304), .B(n1303), .Z(n1308) );
  NANDN U1533 ( .A(n1306), .B(n1305), .Z(n1307) );
  AND U1534 ( .A(n1308), .B(n1307), .Z(n1381) );
  XNOR U1535 ( .A(n1382), .B(n1381), .Z(n1383) );
  XOR U1536 ( .A(n1384), .B(n1383), .Z(n1316) );
  NANDN U1537 ( .A(n1310), .B(n1309), .Z(n1314) );
  NAND U1538 ( .A(n1312), .B(n1311), .Z(n1313) );
  AND U1539 ( .A(n1314), .B(n1313), .Z(n1315) );
  XNOR U1540 ( .A(n1316), .B(n1315), .Z(n1317) );
  XNOR U1541 ( .A(n1318), .B(n1317), .Z(n1387) );
  XNOR U1542 ( .A(sreg[72]), .B(n1387), .Z(n1388) );
  XNOR U1543 ( .A(n1389), .B(n1388), .Z(c[72]) );
  NANDN U1544 ( .A(n1316), .B(n1315), .Z(n1320) );
  NANDN U1545 ( .A(n1318), .B(n1317), .Z(n1319) );
  AND U1546 ( .A(n1320), .B(n1319), .Z(n1395) );
  NANDN U1547 ( .A(n1322), .B(n1321), .Z(n1326) );
  NAND U1548 ( .A(n1324), .B(n1323), .Z(n1325) );
  AND U1549 ( .A(n1326), .B(n1325), .Z(n1461) );
  NANDN U1550 ( .A(n1328), .B(n1327), .Z(n1332) );
  NANDN U1551 ( .A(n1330), .B(n1329), .Z(n1331) );
  AND U1552 ( .A(n1332), .B(n1331), .Z(n1448) );
  NAND U1553 ( .A(b[0]), .B(a[25]), .Z(n1333) );
  XNOR U1554 ( .A(b[1]), .B(n1333), .Z(n1335) );
  NANDN U1555 ( .A(b[0]), .B(a[24]), .Z(n1334) );
  NAND U1556 ( .A(n1335), .B(n1334), .Z(n1428) );
  NAND U1557 ( .A(n5012), .B(n1336), .Z(n1338) );
  XOR U1558 ( .A(b[13]), .B(a[13]), .Z(n1431) );
  NAND U1559 ( .A(n4985), .B(n1431), .Z(n1337) );
  AND U1560 ( .A(n1338), .B(n1337), .Z(n1426) );
  AND U1561 ( .A(b[15]), .B(a[9]), .Z(n1425) );
  XNOR U1562 ( .A(n1426), .B(n1425), .Z(n1427) );
  XNOR U1563 ( .A(n1428), .B(n1427), .Z(n1446) );
  NAND U1564 ( .A(n36), .B(n1339), .Z(n1341) );
  XOR U1565 ( .A(b[5]), .B(a[21]), .Z(n1437) );
  NAND U1566 ( .A(n4560), .B(n1437), .Z(n1340) );
  AND U1567 ( .A(n1341), .B(n1340), .Z(n1422) );
  NAND U1568 ( .A(n4755), .B(n1342), .Z(n1344) );
  XOR U1569 ( .A(b[7]), .B(a[19]), .Z(n1440) );
  NAND U1570 ( .A(n4708), .B(n1440), .Z(n1343) );
  AND U1571 ( .A(n1344), .B(n1343), .Z(n1420) );
  NAND U1572 ( .A(n4471), .B(n1345), .Z(n1347) );
  XOR U1573 ( .A(b[3]), .B(a[23]), .Z(n1443) );
  NAND U1574 ( .A(n33), .B(n1443), .Z(n1346) );
  NAND U1575 ( .A(n1347), .B(n1346), .Z(n1419) );
  XNOR U1576 ( .A(n1420), .B(n1419), .Z(n1421) );
  XOR U1577 ( .A(n1422), .B(n1421), .Z(n1447) );
  XOR U1578 ( .A(n1446), .B(n1447), .Z(n1449) );
  XOR U1579 ( .A(n1448), .B(n1449), .Z(n1399) );
  NANDN U1580 ( .A(n1349), .B(n1348), .Z(n1353) );
  OR U1581 ( .A(n1351), .B(n1350), .Z(n1352) );
  AND U1582 ( .A(n1353), .B(n1352), .Z(n1398) );
  XNOR U1583 ( .A(n1399), .B(n1398), .Z(n1401) );
  NAND U1584 ( .A(n4950), .B(n1354), .Z(n1356) );
  XOR U1585 ( .A(b[11]), .B(a[15]), .Z(n1404) );
  NAND U1586 ( .A(n4863), .B(n1404), .Z(n1355) );
  AND U1587 ( .A(n1356), .B(n1355), .Z(n1415) );
  NAND U1588 ( .A(n42), .B(n1357), .Z(n1359) );
  XOR U1589 ( .A(b[15]), .B(a[11]), .Z(n1407) );
  NAND U1590 ( .A(n4981), .B(n1407), .Z(n1358) );
  AND U1591 ( .A(n1359), .B(n1358), .Z(n1414) );
  NAND U1592 ( .A(n41), .B(n1360), .Z(n1362) );
  XOR U1593 ( .A(b[9]), .B(a[17]), .Z(n1410) );
  NAND U1594 ( .A(n4810), .B(n1410), .Z(n1361) );
  NAND U1595 ( .A(n1362), .B(n1361), .Z(n1413) );
  XOR U1596 ( .A(n1414), .B(n1413), .Z(n1416) );
  XOR U1597 ( .A(n1415), .B(n1416), .Z(n1453) );
  NANDN U1598 ( .A(n1364), .B(n1363), .Z(n1368) );
  OR U1599 ( .A(n1366), .B(n1365), .Z(n1367) );
  AND U1600 ( .A(n1368), .B(n1367), .Z(n1452) );
  XNOR U1601 ( .A(n1453), .B(n1452), .Z(n1454) );
  NANDN U1602 ( .A(n1370), .B(n1369), .Z(n1374) );
  NANDN U1603 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1604 ( .A(n1374), .B(n1373), .Z(n1455) );
  XNOR U1605 ( .A(n1454), .B(n1455), .Z(n1400) );
  XOR U1606 ( .A(n1401), .B(n1400), .Z(n1459) );
  NANDN U1607 ( .A(n1376), .B(n1375), .Z(n1380) );
  NANDN U1608 ( .A(n1378), .B(n1377), .Z(n1379) );
  AND U1609 ( .A(n1380), .B(n1379), .Z(n1458) );
  XNOR U1610 ( .A(n1459), .B(n1458), .Z(n1460) );
  XOR U1611 ( .A(n1461), .B(n1460), .Z(n1393) );
  NANDN U1612 ( .A(n1382), .B(n1381), .Z(n1386) );
  NAND U1613 ( .A(n1384), .B(n1383), .Z(n1385) );
  AND U1614 ( .A(n1386), .B(n1385), .Z(n1392) );
  XNOR U1615 ( .A(n1393), .B(n1392), .Z(n1394) );
  XNOR U1616 ( .A(n1395), .B(n1394), .Z(n1464) );
  XNOR U1617 ( .A(sreg[73]), .B(n1464), .Z(n1466) );
  NANDN U1618 ( .A(sreg[72]), .B(n1387), .Z(n1391) );
  NAND U1619 ( .A(n1389), .B(n1388), .Z(n1390) );
  NAND U1620 ( .A(n1391), .B(n1390), .Z(n1465) );
  XNOR U1621 ( .A(n1466), .B(n1465), .Z(c[73]) );
  NANDN U1622 ( .A(n1393), .B(n1392), .Z(n1397) );
  NANDN U1623 ( .A(n1395), .B(n1394), .Z(n1396) );
  AND U1624 ( .A(n1397), .B(n1396), .Z(n1472) );
  NANDN U1625 ( .A(n1399), .B(n1398), .Z(n1403) );
  NAND U1626 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1627 ( .A(n1403), .B(n1402), .Z(n1538) );
  NAND U1628 ( .A(n4950), .B(n1404), .Z(n1406) );
  XOR U1629 ( .A(b[11]), .B(a[16]), .Z(n1508) );
  NAND U1630 ( .A(n4863), .B(n1508), .Z(n1405) );
  AND U1631 ( .A(n1406), .B(n1405), .Z(n1519) );
  NAND U1632 ( .A(n42), .B(n1407), .Z(n1409) );
  XOR U1633 ( .A(b[15]), .B(a[12]), .Z(n1511) );
  NAND U1634 ( .A(n4981), .B(n1511), .Z(n1408) );
  AND U1635 ( .A(n1409), .B(n1408), .Z(n1518) );
  NAND U1636 ( .A(n41), .B(n1410), .Z(n1412) );
  XOR U1637 ( .A(b[9]), .B(a[18]), .Z(n1514) );
  NAND U1638 ( .A(n4810), .B(n1514), .Z(n1411) );
  NAND U1639 ( .A(n1412), .B(n1411), .Z(n1517) );
  XOR U1640 ( .A(n1518), .B(n1517), .Z(n1520) );
  XOR U1641 ( .A(n1519), .B(n1520), .Z(n1530) );
  NANDN U1642 ( .A(n1414), .B(n1413), .Z(n1418) );
  OR U1643 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1644 ( .A(n1418), .B(n1417), .Z(n1529) );
  XNOR U1645 ( .A(n1530), .B(n1529), .Z(n1531) );
  NANDN U1646 ( .A(n1420), .B(n1419), .Z(n1424) );
  NANDN U1647 ( .A(n1422), .B(n1421), .Z(n1423) );
  NAND U1648 ( .A(n1424), .B(n1423), .Z(n1532) );
  XNOR U1649 ( .A(n1531), .B(n1532), .Z(n1478) );
  NANDN U1650 ( .A(n1426), .B(n1425), .Z(n1430) );
  NANDN U1651 ( .A(n1428), .B(n1427), .Z(n1429) );
  AND U1652 ( .A(n1430), .B(n1429), .Z(n1504) );
  NAND U1653 ( .A(n5012), .B(n1431), .Z(n1433) );
  XOR U1654 ( .A(b[13]), .B(a[14]), .Z(n1487) );
  NAND U1655 ( .A(n4985), .B(n1487), .Z(n1432) );
  AND U1656 ( .A(n1433), .B(n1432), .Z(n1482) );
  AND U1657 ( .A(b[15]), .B(a[10]), .Z(n1481) );
  XNOR U1658 ( .A(n1482), .B(n1481), .Z(n1483) );
  NAND U1659 ( .A(b[0]), .B(a[26]), .Z(n1434) );
  XNOR U1660 ( .A(b[1]), .B(n1434), .Z(n1436) );
  NANDN U1661 ( .A(b[0]), .B(a[25]), .Z(n1435) );
  NAND U1662 ( .A(n1436), .B(n1435), .Z(n1484) );
  XNOR U1663 ( .A(n1483), .B(n1484), .Z(n1502) );
  NAND U1664 ( .A(n36), .B(n1437), .Z(n1439) );
  XOR U1665 ( .A(b[5]), .B(a[22]), .Z(n1493) );
  NAND U1666 ( .A(n4560), .B(n1493), .Z(n1438) );
  AND U1667 ( .A(n1439), .B(n1438), .Z(n1526) );
  NAND U1668 ( .A(n4755), .B(n1440), .Z(n1442) );
  XOR U1669 ( .A(b[7]), .B(a[20]), .Z(n1496) );
  NAND U1670 ( .A(n4708), .B(n1496), .Z(n1441) );
  AND U1671 ( .A(n1442), .B(n1441), .Z(n1524) );
  NAND U1672 ( .A(n4471), .B(n1443), .Z(n1445) );
  XOR U1673 ( .A(b[3]), .B(a[24]), .Z(n1499) );
  NAND U1674 ( .A(n33), .B(n1499), .Z(n1444) );
  NAND U1675 ( .A(n1445), .B(n1444), .Z(n1523) );
  XNOR U1676 ( .A(n1524), .B(n1523), .Z(n1525) );
  XOR U1677 ( .A(n1526), .B(n1525), .Z(n1503) );
  XOR U1678 ( .A(n1502), .B(n1503), .Z(n1505) );
  XOR U1679 ( .A(n1504), .B(n1505), .Z(n1476) );
  NANDN U1680 ( .A(n1447), .B(n1446), .Z(n1451) );
  OR U1681 ( .A(n1449), .B(n1448), .Z(n1450) );
  AND U1682 ( .A(n1451), .B(n1450), .Z(n1475) );
  XNOR U1683 ( .A(n1476), .B(n1475), .Z(n1477) );
  XOR U1684 ( .A(n1478), .B(n1477), .Z(n1536) );
  NANDN U1685 ( .A(n1453), .B(n1452), .Z(n1457) );
  NANDN U1686 ( .A(n1455), .B(n1454), .Z(n1456) );
  AND U1687 ( .A(n1457), .B(n1456), .Z(n1535) );
  XNOR U1688 ( .A(n1536), .B(n1535), .Z(n1537) );
  XOR U1689 ( .A(n1538), .B(n1537), .Z(n1470) );
  NANDN U1690 ( .A(n1459), .B(n1458), .Z(n1463) );
  NAND U1691 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1692 ( .A(n1463), .B(n1462), .Z(n1469) );
  XNOR U1693 ( .A(n1470), .B(n1469), .Z(n1471) );
  XNOR U1694 ( .A(n1472), .B(n1471), .Z(n1541) );
  XNOR U1695 ( .A(sreg[74]), .B(n1541), .Z(n1543) );
  NANDN U1696 ( .A(sreg[73]), .B(n1464), .Z(n1468) );
  NAND U1697 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1698 ( .A(n1468), .B(n1467), .Z(n1542) );
  XNOR U1699 ( .A(n1543), .B(n1542), .Z(c[74]) );
  NANDN U1700 ( .A(n1470), .B(n1469), .Z(n1474) );
  NANDN U1701 ( .A(n1472), .B(n1471), .Z(n1473) );
  AND U1702 ( .A(n1474), .B(n1473), .Z(n1549) );
  NANDN U1703 ( .A(n1476), .B(n1475), .Z(n1480) );
  NAND U1704 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U1705 ( .A(n1480), .B(n1479), .Z(n1615) );
  NANDN U1706 ( .A(n1482), .B(n1481), .Z(n1486) );
  NANDN U1707 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1708 ( .A(n1486), .B(n1485), .Z(n1581) );
  NAND U1709 ( .A(n5012), .B(n1487), .Z(n1489) );
  XOR U1710 ( .A(b[13]), .B(a[15]), .Z(n1567) );
  NAND U1711 ( .A(n4985), .B(n1567), .Z(n1488) );
  AND U1712 ( .A(n1489), .B(n1488), .Z(n1559) );
  AND U1713 ( .A(b[15]), .B(a[11]), .Z(n1558) );
  XNOR U1714 ( .A(n1559), .B(n1558), .Z(n1560) );
  NAND U1715 ( .A(b[0]), .B(a[27]), .Z(n1490) );
  XNOR U1716 ( .A(b[1]), .B(n1490), .Z(n1492) );
  NANDN U1717 ( .A(b[0]), .B(a[26]), .Z(n1491) );
  NAND U1718 ( .A(n1492), .B(n1491), .Z(n1561) );
  XNOR U1719 ( .A(n1560), .B(n1561), .Z(n1579) );
  NAND U1720 ( .A(n36), .B(n1493), .Z(n1495) );
  XOR U1721 ( .A(b[5]), .B(a[23]), .Z(n1570) );
  NAND U1722 ( .A(n4560), .B(n1570), .Z(n1494) );
  AND U1723 ( .A(n1495), .B(n1494), .Z(n1603) );
  NAND U1724 ( .A(n4755), .B(n1496), .Z(n1498) );
  XOR U1725 ( .A(b[7]), .B(a[21]), .Z(n1573) );
  NAND U1726 ( .A(n4708), .B(n1573), .Z(n1497) );
  AND U1727 ( .A(n1498), .B(n1497), .Z(n1601) );
  NAND U1728 ( .A(n4471), .B(n1499), .Z(n1501) );
  XOR U1729 ( .A(b[3]), .B(a[25]), .Z(n1576) );
  NAND U1730 ( .A(n33), .B(n1576), .Z(n1500) );
  NAND U1731 ( .A(n1501), .B(n1500), .Z(n1600) );
  XNOR U1732 ( .A(n1601), .B(n1600), .Z(n1602) );
  XOR U1733 ( .A(n1603), .B(n1602), .Z(n1580) );
  XOR U1734 ( .A(n1579), .B(n1580), .Z(n1582) );
  XOR U1735 ( .A(n1581), .B(n1582), .Z(n1553) );
  NANDN U1736 ( .A(n1503), .B(n1502), .Z(n1507) );
  OR U1737 ( .A(n1505), .B(n1504), .Z(n1506) );
  AND U1738 ( .A(n1507), .B(n1506), .Z(n1552) );
  XNOR U1739 ( .A(n1553), .B(n1552), .Z(n1555) );
  NAND U1740 ( .A(n4950), .B(n1508), .Z(n1510) );
  XOR U1741 ( .A(b[11]), .B(a[17]), .Z(n1585) );
  NAND U1742 ( .A(n4863), .B(n1585), .Z(n1509) );
  AND U1743 ( .A(n1510), .B(n1509), .Z(n1596) );
  NAND U1744 ( .A(n42), .B(n1511), .Z(n1513) );
  XOR U1745 ( .A(b[15]), .B(a[13]), .Z(n1588) );
  NAND U1746 ( .A(n4981), .B(n1588), .Z(n1512) );
  AND U1747 ( .A(n1513), .B(n1512), .Z(n1595) );
  NAND U1748 ( .A(n41), .B(n1514), .Z(n1516) );
  XOR U1749 ( .A(b[9]), .B(a[19]), .Z(n1591) );
  NAND U1750 ( .A(n4810), .B(n1591), .Z(n1515) );
  NAND U1751 ( .A(n1516), .B(n1515), .Z(n1594) );
  XOR U1752 ( .A(n1595), .B(n1594), .Z(n1597) );
  XOR U1753 ( .A(n1596), .B(n1597), .Z(n1607) );
  NANDN U1754 ( .A(n1518), .B(n1517), .Z(n1522) );
  OR U1755 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1756 ( .A(n1522), .B(n1521), .Z(n1606) );
  XNOR U1757 ( .A(n1607), .B(n1606), .Z(n1608) );
  NANDN U1758 ( .A(n1524), .B(n1523), .Z(n1528) );
  NANDN U1759 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1760 ( .A(n1528), .B(n1527), .Z(n1609) );
  XNOR U1761 ( .A(n1608), .B(n1609), .Z(n1554) );
  XOR U1762 ( .A(n1555), .B(n1554), .Z(n1613) );
  NANDN U1763 ( .A(n1530), .B(n1529), .Z(n1534) );
  NANDN U1764 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1765 ( .A(n1534), .B(n1533), .Z(n1612) );
  XNOR U1766 ( .A(n1613), .B(n1612), .Z(n1614) );
  XOR U1767 ( .A(n1615), .B(n1614), .Z(n1547) );
  NANDN U1768 ( .A(n1536), .B(n1535), .Z(n1540) );
  NAND U1769 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1770 ( .A(n1540), .B(n1539), .Z(n1546) );
  XNOR U1771 ( .A(n1547), .B(n1546), .Z(n1548) );
  XNOR U1772 ( .A(n1549), .B(n1548), .Z(n1618) );
  XNOR U1773 ( .A(sreg[75]), .B(n1618), .Z(n1620) );
  NANDN U1774 ( .A(sreg[74]), .B(n1541), .Z(n1545) );
  NAND U1775 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U1776 ( .A(n1545), .B(n1544), .Z(n1619) );
  XNOR U1777 ( .A(n1620), .B(n1619), .Z(c[75]) );
  NANDN U1778 ( .A(n1547), .B(n1546), .Z(n1551) );
  NANDN U1779 ( .A(n1549), .B(n1548), .Z(n1550) );
  AND U1780 ( .A(n1551), .B(n1550), .Z(n1626) );
  NANDN U1781 ( .A(n1553), .B(n1552), .Z(n1557) );
  NAND U1782 ( .A(n1555), .B(n1554), .Z(n1556) );
  AND U1783 ( .A(n1557), .B(n1556), .Z(n1692) );
  NANDN U1784 ( .A(n1559), .B(n1558), .Z(n1563) );
  NANDN U1785 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1786 ( .A(n1563), .B(n1562), .Z(n1658) );
  NAND U1787 ( .A(b[0]), .B(a[28]), .Z(n1564) );
  XNOR U1788 ( .A(b[1]), .B(n1564), .Z(n1566) );
  NANDN U1789 ( .A(b[0]), .B(a[27]), .Z(n1565) );
  NAND U1790 ( .A(n1566), .B(n1565), .Z(n1638) );
  NAND U1791 ( .A(n5012), .B(n1567), .Z(n1569) );
  XOR U1792 ( .A(b[13]), .B(a[16]), .Z(n1644) );
  NAND U1793 ( .A(n4985), .B(n1644), .Z(n1568) );
  AND U1794 ( .A(n1569), .B(n1568), .Z(n1636) );
  AND U1795 ( .A(b[15]), .B(a[12]), .Z(n1635) );
  XNOR U1796 ( .A(n1636), .B(n1635), .Z(n1637) );
  XNOR U1797 ( .A(n1638), .B(n1637), .Z(n1656) );
  NAND U1798 ( .A(n36), .B(n1570), .Z(n1572) );
  XOR U1799 ( .A(b[5]), .B(a[24]), .Z(n1647) );
  NAND U1800 ( .A(n4560), .B(n1647), .Z(n1571) );
  AND U1801 ( .A(n1572), .B(n1571), .Z(n1680) );
  NAND U1802 ( .A(n4755), .B(n1573), .Z(n1575) );
  XOR U1803 ( .A(b[7]), .B(a[22]), .Z(n1650) );
  NAND U1804 ( .A(n4708), .B(n1650), .Z(n1574) );
  AND U1805 ( .A(n1575), .B(n1574), .Z(n1678) );
  NAND U1806 ( .A(n4471), .B(n1576), .Z(n1578) );
  XOR U1807 ( .A(b[3]), .B(a[26]), .Z(n1653) );
  NAND U1808 ( .A(n33), .B(n1653), .Z(n1577) );
  NAND U1809 ( .A(n1578), .B(n1577), .Z(n1677) );
  XNOR U1810 ( .A(n1678), .B(n1677), .Z(n1679) );
  XOR U1811 ( .A(n1680), .B(n1679), .Z(n1657) );
  XOR U1812 ( .A(n1656), .B(n1657), .Z(n1659) );
  XOR U1813 ( .A(n1658), .B(n1659), .Z(n1630) );
  NANDN U1814 ( .A(n1580), .B(n1579), .Z(n1584) );
  OR U1815 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U1816 ( .A(n1584), .B(n1583), .Z(n1629) );
  XNOR U1817 ( .A(n1630), .B(n1629), .Z(n1632) );
  NAND U1818 ( .A(n4950), .B(n1585), .Z(n1587) );
  XOR U1819 ( .A(b[11]), .B(a[18]), .Z(n1662) );
  NAND U1820 ( .A(n4863), .B(n1662), .Z(n1586) );
  AND U1821 ( .A(n1587), .B(n1586), .Z(n1673) );
  NAND U1822 ( .A(n42), .B(n1588), .Z(n1590) );
  XOR U1823 ( .A(b[15]), .B(a[14]), .Z(n1665) );
  NAND U1824 ( .A(n4981), .B(n1665), .Z(n1589) );
  AND U1825 ( .A(n1590), .B(n1589), .Z(n1672) );
  NAND U1826 ( .A(n41), .B(n1591), .Z(n1593) );
  XOR U1827 ( .A(b[9]), .B(a[20]), .Z(n1668) );
  NAND U1828 ( .A(n4810), .B(n1668), .Z(n1592) );
  NAND U1829 ( .A(n1593), .B(n1592), .Z(n1671) );
  XOR U1830 ( .A(n1672), .B(n1671), .Z(n1674) );
  XOR U1831 ( .A(n1673), .B(n1674), .Z(n1684) );
  NANDN U1832 ( .A(n1595), .B(n1594), .Z(n1599) );
  OR U1833 ( .A(n1597), .B(n1596), .Z(n1598) );
  AND U1834 ( .A(n1599), .B(n1598), .Z(n1683) );
  XNOR U1835 ( .A(n1684), .B(n1683), .Z(n1685) );
  NANDN U1836 ( .A(n1601), .B(n1600), .Z(n1605) );
  NANDN U1837 ( .A(n1603), .B(n1602), .Z(n1604) );
  NAND U1838 ( .A(n1605), .B(n1604), .Z(n1686) );
  XNOR U1839 ( .A(n1685), .B(n1686), .Z(n1631) );
  XOR U1840 ( .A(n1632), .B(n1631), .Z(n1690) );
  NANDN U1841 ( .A(n1607), .B(n1606), .Z(n1611) );
  NANDN U1842 ( .A(n1609), .B(n1608), .Z(n1610) );
  AND U1843 ( .A(n1611), .B(n1610), .Z(n1689) );
  XNOR U1844 ( .A(n1690), .B(n1689), .Z(n1691) );
  XOR U1845 ( .A(n1692), .B(n1691), .Z(n1624) );
  NANDN U1846 ( .A(n1613), .B(n1612), .Z(n1617) );
  NAND U1847 ( .A(n1615), .B(n1614), .Z(n1616) );
  AND U1848 ( .A(n1617), .B(n1616), .Z(n1623) );
  XNOR U1849 ( .A(n1624), .B(n1623), .Z(n1625) );
  XNOR U1850 ( .A(n1626), .B(n1625), .Z(n1695) );
  XNOR U1851 ( .A(sreg[76]), .B(n1695), .Z(n1697) );
  NANDN U1852 ( .A(sreg[75]), .B(n1618), .Z(n1622) );
  NAND U1853 ( .A(n1620), .B(n1619), .Z(n1621) );
  NAND U1854 ( .A(n1622), .B(n1621), .Z(n1696) );
  XNOR U1855 ( .A(n1697), .B(n1696), .Z(c[76]) );
  NANDN U1856 ( .A(n1624), .B(n1623), .Z(n1628) );
  NANDN U1857 ( .A(n1626), .B(n1625), .Z(n1627) );
  AND U1858 ( .A(n1628), .B(n1627), .Z(n1703) );
  NANDN U1859 ( .A(n1630), .B(n1629), .Z(n1634) );
  NAND U1860 ( .A(n1632), .B(n1631), .Z(n1633) );
  AND U1861 ( .A(n1634), .B(n1633), .Z(n1769) );
  NANDN U1862 ( .A(n1636), .B(n1635), .Z(n1640) );
  NANDN U1863 ( .A(n1638), .B(n1637), .Z(n1639) );
  AND U1864 ( .A(n1640), .B(n1639), .Z(n1735) );
  NAND U1865 ( .A(b[0]), .B(a[29]), .Z(n1641) );
  XNOR U1866 ( .A(b[1]), .B(n1641), .Z(n1643) );
  NANDN U1867 ( .A(b[0]), .B(a[28]), .Z(n1642) );
  NAND U1868 ( .A(n1643), .B(n1642), .Z(n1715) );
  NAND U1869 ( .A(n5012), .B(n1644), .Z(n1646) );
  XOR U1870 ( .A(b[13]), .B(a[17]), .Z(n1721) );
  NAND U1871 ( .A(n4985), .B(n1721), .Z(n1645) );
  AND U1872 ( .A(n1646), .B(n1645), .Z(n1713) );
  AND U1873 ( .A(b[15]), .B(a[13]), .Z(n1712) );
  XNOR U1874 ( .A(n1713), .B(n1712), .Z(n1714) );
  XNOR U1875 ( .A(n1715), .B(n1714), .Z(n1733) );
  NAND U1876 ( .A(n36), .B(n1647), .Z(n1649) );
  XOR U1877 ( .A(b[5]), .B(a[25]), .Z(n1724) );
  NAND U1878 ( .A(n4560), .B(n1724), .Z(n1648) );
  AND U1879 ( .A(n1649), .B(n1648), .Z(n1757) );
  NAND U1880 ( .A(n4755), .B(n1650), .Z(n1652) );
  XOR U1881 ( .A(b[7]), .B(a[23]), .Z(n1727) );
  NAND U1882 ( .A(n4708), .B(n1727), .Z(n1651) );
  AND U1883 ( .A(n1652), .B(n1651), .Z(n1755) );
  NAND U1884 ( .A(n4471), .B(n1653), .Z(n1655) );
  XOR U1885 ( .A(b[3]), .B(a[27]), .Z(n1730) );
  NAND U1886 ( .A(n33), .B(n1730), .Z(n1654) );
  NAND U1887 ( .A(n1655), .B(n1654), .Z(n1754) );
  XNOR U1888 ( .A(n1755), .B(n1754), .Z(n1756) );
  XOR U1889 ( .A(n1757), .B(n1756), .Z(n1734) );
  XOR U1890 ( .A(n1733), .B(n1734), .Z(n1736) );
  XOR U1891 ( .A(n1735), .B(n1736), .Z(n1707) );
  NANDN U1892 ( .A(n1657), .B(n1656), .Z(n1661) );
  OR U1893 ( .A(n1659), .B(n1658), .Z(n1660) );
  AND U1894 ( .A(n1661), .B(n1660), .Z(n1706) );
  XNOR U1895 ( .A(n1707), .B(n1706), .Z(n1709) );
  NAND U1896 ( .A(n4950), .B(n1662), .Z(n1664) );
  XOR U1897 ( .A(b[11]), .B(a[19]), .Z(n1739) );
  NAND U1898 ( .A(n4863), .B(n1739), .Z(n1663) );
  AND U1899 ( .A(n1664), .B(n1663), .Z(n1750) );
  NAND U1900 ( .A(n42), .B(n1665), .Z(n1667) );
  XOR U1901 ( .A(b[15]), .B(a[15]), .Z(n1742) );
  NAND U1902 ( .A(n4981), .B(n1742), .Z(n1666) );
  AND U1903 ( .A(n1667), .B(n1666), .Z(n1749) );
  NAND U1904 ( .A(n41), .B(n1668), .Z(n1670) );
  XOR U1905 ( .A(b[9]), .B(a[21]), .Z(n1745) );
  NAND U1906 ( .A(n4810), .B(n1745), .Z(n1669) );
  NAND U1907 ( .A(n1670), .B(n1669), .Z(n1748) );
  XOR U1908 ( .A(n1749), .B(n1748), .Z(n1751) );
  XOR U1909 ( .A(n1750), .B(n1751), .Z(n1761) );
  NANDN U1910 ( .A(n1672), .B(n1671), .Z(n1676) );
  OR U1911 ( .A(n1674), .B(n1673), .Z(n1675) );
  AND U1912 ( .A(n1676), .B(n1675), .Z(n1760) );
  XNOR U1913 ( .A(n1761), .B(n1760), .Z(n1762) );
  NANDN U1914 ( .A(n1678), .B(n1677), .Z(n1682) );
  NANDN U1915 ( .A(n1680), .B(n1679), .Z(n1681) );
  NAND U1916 ( .A(n1682), .B(n1681), .Z(n1763) );
  XNOR U1917 ( .A(n1762), .B(n1763), .Z(n1708) );
  XOR U1918 ( .A(n1709), .B(n1708), .Z(n1767) );
  NANDN U1919 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U1920 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U1921 ( .A(n1688), .B(n1687), .Z(n1766) );
  XNOR U1922 ( .A(n1767), .B(n1766), .Z(n1768) );
  XOR U1923 ( .A(n1769), .B(n1768), .Z(n1701) );
  NANDN U1924 ( .A(n1690), .B(n1689), .Z(n1694) );
  NAND U1925 ( .A(n1692), .B(n1691), .Z(n1693) );
  AND U1926 ( .A(n1694), .B(n1693), .Z(n1700) );
  XNOR U1927 ( .A(n1701), .B(n1700), .Z(n1702) );
  XNOR U1928 ( .A(n1703), .B(n1702), .Z(n1772) );
  XNOR U1929 ( .A(sreg[77]), .B(n1772), .Z(n1774) );
  NANDN U1930 ( .A(sreg[76]), .B(n1695), .Z(n1699) );
  NAND U1931 ( .A(n1697), .B(n1696), .Z(n1698) );
  NAND U1932 ( .A(n1699), .B(n1698), .Z(n1773) );
  XNOR U1933 ( .A(n1774), .B(n1773), .Z(c[77]) );
  NANDN U1934 ( .A(n1701), .B(n1700), .Z(n1705) );
  NANDN U1935 ( .A(n1703), .B(n1702), .Z(n1704) );
  AND U1936 ( .A(n1705), .B(n1704), .Z(n1780) );
  NANDN U1937 ( .A(n1707), .B(n1706), .Z(n1711) );
  NAND U1938 ( .A(n1709), .B(n1708), .Z(n1710) );
  AND U1939 ( .A(n1711), .B(n1710), .Z(n1846) );
  NANDN U1940 ( .A(n1713), .B(n1712), .Z(n1717) );
  NANDN U1941 ( .A(n1715), .B(n1714), .Z(n1716) );
  AND U1942 ( .A(n1717), .B(n1716), .Z(n1812) );
  NAND U1943 ( .A(b[0]), .B(a[30]), .Z(n1718) );
  XNOR U1944 ( .A(b[1]), .B(n1718), .Z(n1720) );
  NANDN U1945 ( .A(b[0]), .B(a[29]), .Z(n1719) );
  NAND U1946 ( .A(n1720), .B(n1719), .Z(n1792) );
  NAND U1947 ( .A(n5012), .B(n1721), .Z(n1723) );
  XOR U1948 ( .A(b[13]), .B(a[18]), .Z(n1798) );
  NAND U1949 ( .A(n4985), .B(n1798), .Z(n1722) );
  AND U1950 ( .A(n1723), .B(n1722), .Z(n1790) );
  AND U1951 ( .A(b[15]), .B(a[14]), .Z(n1789) );
  XNOR U1952 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U1953 ( .A(n1792), .B(n1791), .Z(n1810) );
  NAND U1954 ( .A(n36), .B(n1724), .Z(n1726) );
  XOR U1955 ( .A(b[5]), .B(a[26]), .Z(n1801) );
  NAND U1956 ( .A(n4560), .B(n1801), .Z(n1725) );
  AND U1957 ( .A(n1726), .B(n1725), .Z(n1834) );
  NAND U1958 ( .A(n4755), .B(n1727), .Z(n1729) );
  XOR U1959 ( .A(b[7]), .B(a[24]), .Z(n1804) );
  NAND U1960 ( .A(n4708), .B(n1804), .Z(n1728) );
  AND U1961 ( .A(n1729), .B(n1728), .Z(n1832) );
  NAND U1962 ( .A(n4471), .B(n1730), .Z(n1732) );
  XOR U1963 ( .A(b[3]), .B(a[28]), .Z(n1807) );
  NAND U1964 ( .A(n33), .B(n1807), .Z(n1731) );
  NAND U1965 ( .A(n1732), .B(n1731), .Z(n1831) );
  XNOR U1966 ( .A(n1832), .B(n1831), .Z(n1833) );
  XOR U1967 ( .A(n1834), .B(n1833), .Z(n1811) );
  XOR U1968 ( .A(n1810), .B(n1811), .Z(n1813) );
  XOR U1969 ( .A(n1812), .B(n1813), .Z(n1784) );
  NANDN U1970 ( .A(n1734), .B(n1733), .Z(n1738) );
  OR U1971 ( .A(n1736), .B(n1735), .Z(n1737) );
  AND U1972 ( .A(n1738), .B(n1737), .Z(n1783) );
  XNOR U1973 ( .A(n1784), .B(n1783), .Z(n1786) );
  NAND U1974 ( .A(n4950), .B(n1739), .Z(n1741) );
  XOR U1975 ( .A(b[11]), .B(a[20]), .Z(n1816) );
  NAND U1976 ( .A(n4863), .B(n1816), .Z(n1740) );
  AND U1977 ( .A(n1741), .B(n1740), .Z(n1827) );
  NAND U1978 ( .A(n42), .B(n1742), .Z(n1744) );
  XOR U1979 ( .A(b[15]), .B(a[16]), .Z(n1819) );
  NAND U1980 ( .A(n4981), .B(n1819), .Z(n1743) );
  AND U1981 ( .A(n1744), .B(n1743), .Z(n1826) );
  NAND U1982 ( .A(n41), .B(n1745), .Z(n1747) );
  XOR U1983 ( .A(b[9]), .B(a[22]), .Z(n1822) );
  NAND U1984 ( .A(n4810), .B(n1822), .Z(n1746) );
  NAND U1985 ( .A(n1747), .B(n1746), .Z(n1825) );
  XOR U1986 ( .A(n1826), .B(n1825), .Z(n1828) );
  XOR U1987 ( .A(n1827), .B(n1828), .Z(n1838) );
  NANDN U1988 ( .A(n1749), .B(n1748), .Z(n1753) );
  OR U1989 ( .A(n1751), .B(n1750), .Z(n1752) );
  AND U1990 ( .A(n1753), .B(n1752), .Z(n1837) );
  XNOR U1991 ( .A(n1838), .B(n1837), .Z(n1839) );
  NANDN U1992 ( .A(n1755), .B(n1754), .Z(n1759) );
  NANDN U1993 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U1994 ( .A(n1759), .B(n1758), .Z(n1840) );
  XNOR U1995 ( .A(n1839), .B(n1840), .Z(n1785) );
  XOR U1996 ( .A(n1786), .B(n1785), .Z(n1844) );
  NANDN U1997 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U1998 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U1999 ( .A(n1765), .B(n1764), .Z(n1843) );
  XNOR U2000 ( .A(n1844), .B(n1843), .Z(n1845) );
  XOR U2001 ( .A(n1846), .B(n1845), .Z(n1778) );
  NANDN U2002 ( .A(n1767), .B(n1766), .Z(n1771) );
  NAND U2003 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U2004 ( .A(n1771), .B(n1770), .Z(n1777) );
  XNOR U2005 ( .A(n1778), .B(n1777), .Z(n1779) );
  XNOR U2006 ( .A(n1780), .B(n1779), .Z(n1849) );
  XNOR U2007 ( .A(sreg[78]), .B(n1849), .Z(n1851) );
  NANDN U2008 ( .A(sreg[77]), .B(n1772), .Z(n1776) );
  NAND U2009 ( .A(n1774), .B(n1773), .Z(n1775) );
  NAND U2010 ( .A(n1776), .B(n1775), .Z(n1850) );
  XNOR U2011 ( .A(n1851), .B(n1850), .Z(c[78]) );
  NANDN U2012 ( .A(n1778), .B(n1777), .Z(n1782) );
  NANDN U2013 ( .A(n1780), .B(n1779), .Z(n1781) );
  AND U2014 ( .A(n1782), .B(n1781), .Z(n1857) );
  NANDN U2015 ( .A(n1784), .B(n1783), .Z(n1788) );
  NAND U2016 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2017 ( .A(n1788), .B(n1787), .Z(n1923) );
  NANDN U2018 ( .A(n1790), .B(n1789), .Z(n1794) );
  NANDN U2019 ( .A(n1792), .B(n1791), .Z(n1793) );
  AND U2020 ( .A(n1794), .B(n1793), .Z(n1889) );
  NAND U2021 ( .A(b[0]), .B(a[31]), .Z(n1795) );
  XNOR U2022 ( .A(b[1]), .B(n1795), .Z(n1797) );
  NANDN U2023 ( .A(b[0]), .B(a[30]), .Z(n1796) );
  NAND U2024 ( .A(n1797), .B(n1796), .Z(n1869) );
  NAND U2025 ( .A(n5012), .B(n1798), .Z(n1800) );
  XOR U2026 ( .A(b[13]), .B(a[19]), .Z(n1872) );
  NAND U2027 ( .A(n4985), .B(n1872), .Z(n1799) );
  AND U2028 ( .A(n1800), .B(n1799), .Z(n1867) );
  AND U2029 ( .A(b[15]), .B(a[15]), .Z(n1866) );
  XNOR U2030 ( .A(n1867), .B(n1866), .Z(n1868) );
  XNOR U2031 ( .A(n1869), .B(n1868), .Z(n1887) );
  NAND U2032 ( .A(n36), .B(n1801), .Z(n1803) );
  XOR U2033 ( .A(b[5]), .B(a[27]), .Z(n1878) );
  NAND U2034 ( .A(n4560), .B(n1878), .Z(n1802) );
  AND U2035 ( .A(n1803), .B(n1802), .Z(n1911) );
  NAND U2036 ( .A(n4755), .B(n1804), .Z(n1806) );
  XOR U2037 ( .A(b[7]), .B(a[25]), .Z(n1881) );
  NAND U2038 ( .A(n4708), .B(n1881), .Z(n1805) );
  AND U2039 ( .A(n1806), .B(n1805), .Z(n1909) );
  NAND U2040 ( .A(n4471), .B(n1807), .Z(n1809) );
  XOR U2041 ( .A(b[3]), .B(a[29]), .Z(n1884) );
  NAND U2042 ( .A(n33), .B(n1884), .Z(n1808) );
  NAND U2043 ( .A(n1809), .B(n1808), .Z(n1908) );
  XNOR U2044 ( .A(n1909), .B(n1908), .Z(n1910) );
  XOR U2045 ( .A(n1911), .B(n1910), .Z(n1888) );
  XOR U2046 ( .A(n1887), .B(n1888), .Z(n1890) );
  XOR U2047 ( .A(n1889), .B(n1890), .Z(n1861) );
  NANDN U2048 ( .A(n1811), .B(n1810), .Z(n1815) );
  OR U2049 ( .A(n1813), .B(n1812), .Z(n1814) );
  AND U2050 ( .A(n1815), .B(n1814), .Z(n1860) );
  XNOR U2051 ( .A(n1861), .B(n1860), .Z(n1863) );
  NAND U2052 ( .A(n4950), .B(n1816), .Z(n1818) );
  XOR U2053 ( .A(b[11]), .B(a[21]), .Z(n1893) );
  NAND U2054 ( .A(n4863), .B(n1893), .Z(n1817) );
  AND U2055 ( .A(n1818), .B(n1817), .Z(n1904) );
  NAND U2056 ( .A(n42), .B(n1819), .Z(n1821) );
  XOR U2057 ( .A(b[15]), .B(a[17]), .Z(n1896) );
  NAND U2058 ( .A(n4981), .B(n1896), .Z(n1820) );
  AND U2059 ( .A(n1821), .B(n1820), .Z(n1903) );
  NAND U2060 ( .A(n41), .B(n1822), .Z(n1824) );
  XOR U2061 ( .A(b[9]), .B(a[23]), .Z(n1899) );
  NAND U2062 ( .A(n4810), .B(n1899), .Z(n1823) );
  NAND U2063 ( .A(n1824), .B(n1823), .Z(n1902) );
  XOR U2064 ( .A(n1903), .B(n1902), .Z(n1905) );
  XOR U2065 ( .A(n1904), .B(n1905), .Z(n1915) );
  NANDN U2066 ( .A(n1826), .B(n1825), .Z(n1830) );
  OR U2067 ( .A(n1828), .B(n1827), .Z(n1829) );
  AND U2068 ( .A(n1830), .B(n1829), .Z(n1914) );
  XNOR U2069 ( .A(n1915), .B(n1914), .Z(n1916) );
  NANDN U2070 ( .A(n1832), .B(n1831), .Z(n1836) );
  NANDN U2071 ( .A(n1834), .B(n1833), .Z(n1835) );
  NAND U2072 ( .A(n1836), .B(n1835), .Z(n1917) );
  XNOR U2073 ( .A(n1916), .B(n1917), .Z(n1862) );
  XOR U2074 ( .A(n1863), .B(n1862), .Z(n1921) );
  NANDN U2075 ( .A(n1838), .B(n1837), .Z(n1842) );
  NANDN U2076 ( .A(n1840), .B(n1839), .Z(n1841) );
  AND U2077 ( .A(n1842), .B(n1841), .Z(n1920) );
  XNOR U2078 ( .A(n1921), .B(n1920), .Z(n1922) );
  XOR U2079 ( .A(n1923), .B(n1922), .Z(n1855) );
  NANDN U2080 ( .A(n1844), .B(n1843), .Z(n1848) );
  NAND U2081 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U2082 ( .A(n1848), .B(n1847), .Z(n1854) );
  XNOR U2083 ( .A(n1855), .B(n1854), .Z(n1856) );
  XNOR U2084 ( .A(n1857), .B(n1856), .Z(n1926) );
  XNOR U2085 ( .A(sreg[79]), .B(n1926), .Z(n1928) );
  NANDN U2086 ( .A(sreg[78]), .B(n1849), .Z(n1853) );
  NAND U2087 ( .A(n1851), .B(n1850), .Z(n1852) );
  NAND U2088 ( .A(n1853), .B(n1852), .Z(n1927) );
  XNOR U2089 ( .A(n1928), .B(n1927), .Z(c[79]) );
  NANDN U2090 ( .A(n1855), .B(n1854), .Z(n1859) );
  NANDN U2091 ( .A(n1857), .B(n1856), .Z(n1858) );
  AND U2092 ( .A(n1859), .B(n1858), .Z(n1934) );
  NANDN U2093 ( .A(n1861), .B(n1860), .Z(n1865) );
  NAND U2094 ( .A(n1863), .B(n1862), .Z(n1864) );
  AND U2095 ( .A(n1865), .B(n1864), .Z(n2000) );
  NANDN U2096 ( .A(n1867), .B(n1866), .Z(n1871) );
  NANDN U2097 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2098 ( .A(n1871), .B(n1870), .Z(n1966) );
  NAND U2099 ( .A(n5012), .B(n1872), .Z(n1874) );
  XOR U2100 ( .A(b[13]), .B(a[20]), .Z(n1949) );
  NAND U2101 ( .A(n4985), .B(n1949), .Z(n1873) );
  AND U2102 ( .A(n1874), .B(n1873), .Z(n1944) );
  AND U2103 ( .A(b[15]), .B(a[16]), .Z(n1943) );
  XNOR U2104 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2105 ( .A(b[0]), .B(a[32]), .Z(n1875) );
  XNOR U2106 ( .A(b[1]), .B(n1875), .Z(n1877) );
  NANDN U2107 ( .A(b[0]), .B(a[31]), .Z(n1876) );
  NAND U2108 ( .A(n1877), .B(n1876), .Z(n1946) );
  XNOR U2109 ( .A(n1945), .B(n1946), .Z(n1964) );
  NAND U2110 ( .A(n36), .B(n1878), .Z(n1880) );
  XOR U2111 ( .A(b[5]), .B(a[28]), .Z(n1955) );
  NAND U2112 ( .A(n4560), .B(n1955), .Z(n1879) );
  AND U2113 ( .A(n1880), .B(n1879), .Z(n1988) );
  NAND U2114 ( .A(n4755), .B(n1881), .Z(n1883) );
  XOR U2115 ( .A(b[7]), .B(a[26]), .Z(n1958) );
  NAND U2116 ( .A(n4708), .B(n1958), .Z(n1882) );
  AND U2117 ( .A(n1883), .B(n1882), .Z(n1986) );
  NAND U2118 ( .A(n4471), .B(n1884), .Z(n1886) );
  XOR U2119 ( .A(b[3]), .B(a[30]), .Z(n1961) );
  NAND U2120 ( .A(n33), .B(n1961), .Z(n1885) );
  NAND U2121 ( .A(n1886), .B(n1885), .Z(n1985) );
  XNOR U2122 ( .A(n1986), .B(n1985), .Z(n1987) );
  XOR U2123 ( .A(n1988), .B(n1987), .Z(n1965) );
  XOR U2124 ( .A(n1964), .B(n1965), .Z(n1967) );
  XOR U2125 ( .A(n1966), .B(n1967), .Z(n1938) );
  NANDN U2126 ( .A(n1888), .B(n1887), .Z(n1892) );
  OR U2127 ( .A(n1890), .B(n1889), .Z(n1891) );
  AND U2128 ( .A(n1892), .B(n1891), .Z(n1937) );
  XNOR U2129 ( .A(n1938), .B(n1937), .Z(n1940) );
  NAND U2130 ( .A(n4950), .B(n1893), .Z(n1895) );
  XOR U2131 ( .A(b[11]), .B(a[22]), .Z(n1970) );
  NAND U2132 ( .A(n4863), .B(n1970), .Z(n1894) );
  AND U2133 ( .A(n1895), .B(n1894), .Z(n1981) );
  NAND U2134 ( .A(n42), .B(n1896), .Z(n1898) );
  XOR U2135 ( .A(b[15]), .B(a[18]), .Z(n1973) );
  NAND U2136 ( .A(n4981), .B(n1973), .Z(n1897) );
  AND U2137 ( .A(n1898), .B(n1897), .Z(n1980) );
  NAND U2138 ( .A(n41), .B(n1899), .Z(n1901) );
  XOR U2139 ( .A(b[9]), .B(a[24]), .Z(n1976) );
  NAND U2140 ( .A(n4810), .B(n1976), .Z(n1900) );
  NAND U2141 ( .A(n1901), .B(n1900), .Z(n1979) );
  XOR U2142 ( .A(n1980), .B(n1979), .Z(n1982) );
  XOR U2143 ( .A(n1981), .B(n1982), .Z(n1992) );
  NANDN U2144 ( .A(n1903), .B(n1902), .Z(n1907) );
  OR U2145 ( .A(n1905), .B(n1904), .Z(n1906) );
  AND U2146 ( .A(n1907), .B(n1906), .Z(n1991) );
  XNOR U2147 ( .A(n1992), .B(n1991), .Z(n1993) );
  NANDN U2148 ( .A(n1909), .B(n1908), .Z(n1913) );
  NANDN U2149 ( .A(n1911), .B(n1910), .Z(n1912) );
  NAND U2150 ( .A(n1913), .B(n1912), .Z(n1994) );
  XNOR U2151 ( .A(n1993), .B(n1994), .Z(n1939) );
  XOR U2152 ( .A(n1940), .B(n1939), .Z(n1998) );
  NANDN U2153 ( .A(n1915), .B(n1914), .Z(n1919) );
  NANDN U2154 ( .A(n1917), .B(n1916), .Z(n1918) );
  AND U2155 ( .A(n1919), .B(n1918), .Z(n1997) );
  XNOR U2156 ( .A(n1998), .B(n1997), .Z(n1999) );
  XOR U2157 ( .A(n2000), .B(n1999), .Z(n1932) );
  NANDN U2158 ( .A(n1921), .B(n1920), .Z(n1925) );
  NAND U2159 ( .A(n1923), .B(n1922), .Z(n1924) );
  AND U2160 ( .A(n1925), .B(n1924), .Z(n1931) );
  XNOR U2161 ( .A(n1932), .B(n1931), .Z(n1933) );
  XNOR U2162 ( .A(n1934), .B(n1933), .Z(n2003) );
  XNOR U2163 ( .A(sreg[80]), .B(n2003), .Z(n2005) );
  NANDN U2164 ( .A(sreg[79]), .B(n1926), .Z(n1930) );
  NAND U2165 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2166 ( .A(n1930), .B(n1929), .Z(n2004) );
  XNOR U2167 ( .A(n2005), .B(n2004), .Z(c[80]) );
  NANDN U2168 ( .A(n1932), .B(n1931), .Z(n1936) );
  NANDN U2169 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U2170 ( .A(n1936), .B(n1935), .Z(n2011) );
  NANDN U2171 ( .A(n1938), .B(n1937), .Z(n1942) );
  NAND U2172 ( .A(n1940), .B(n1939), .Z(n1941) );
  AND U2173 ( .A(n1942), .B(n1941), .Z(n2077) );
  NANDN U2174 ( .A(n1944), .B(n1943), .Z(n1948) );
  NANDN U2175 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2176 ( .A(n1948), .B(n1947), .Z(n2043) );
  NAND U2177 ( .A(n5012), .B(n1949), .Z(n1951) );
  XOR U2178 ( .A(b[13]), .B(a[21]), .Z(n2029) );
  NAND U2179 ( .A(n4985), .B(n2029), .Z(n1950) );
  AND U2180 ( .A(n1951), .B(n1950), .Z(n2021) );
  AND U2181 ( .A(b[15]), .B(a[17]), .Z(n2020) );
  XNOR U2182 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U2183 ( .A(b[0]), .B(a[33]), .Z(n1952) );
  XNOR U2184 ( .A(b[1]), .B(n1952), .Z(n1954) );
  NANDN U2185 ( .A(b[0]), .B(a[32]), .Z(n1953) );
  NAND U2186 ( .A(n1954), .B(n1953), .Z(n2023) );
  XNOR U2187 ( .A(n2022), .B(n2023), .Z(n2041) );
  NAND U2188 ( .A(n36), .B(n1955), .Z(n1957) );
  XOR U2189 ( .A(b[5]), .B(a[29]), .Z(n2032) );
  NAND U2190 ( .A(n4560), .B(n2032), .Z(n1956) );
  AND U2191 ( .A(n1957), .B(n1956), .Z(n2065) );
  NAND U2192 ( .A(n4755), .B(n1958), .Z(n1960) );
  XOR U2193 ( .A(b[7]), .B(a[27]), .Z(n2035) );
  NAND U2194 ( .A(n4708), .B(n2035), .Z(n1959) );
  AND U2195 ( .A(n1960), .B(n1959), .Z(n2063) );
  NAND U2196 ( .A(n4471), .B(n1961), .Z(n1963) );
  XOR U2197 ( .A(b[3]), .B(a[31]), .Z(n2038) );
  NAND U2198 ( .A(n33), .B(n2038), .Z(n1962) );
  NAND U2199 ( .A(n1963), .B(n1962), .Z(n2062) );
  XNOR U2200 ( .A(n2063), .B(n2062), .Z(n2064) );
  XOR U2201 ( .A(n2065), .B(n2064), .Z(n2042) );
  XOR U2202 ( .A(n2041), .B(n2042), .Z(n2044) );
  XOR U2203 ( .A(n2043), .B(n2044), .Z(n2015) );
  NANDN U2204 ( .A(n1965), .B(n1964), .Z(n1969) );
  OR U2205 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2206 ( .A(n1969), .B(n1968), .Z(n2014) );
  XNOR U2207 ( .A(n2015), .B(n2014), .Z(n2017) );
  NAND U2208 ( .A(n4950), .B(n1970), .Z(n1972) );
  XOR U2209 ( .A(b[11]), .B(a[23]), .Z(n2047) );
  NAND U2210 ( .A(n4863), .B(n2047), .Z(n1971) );
  AND U2211 ( .A(n1972), .B(n1971), .Z(n2058) );
  NAND U2212 ( .A(n42), .B(n1973), .Z(n1975) );
  XOR U2213 ( .A(b[15]), .B(a[19]), .Z(n2050) );
  NAND U2214 ( .A(n4981), .B(n2050), .Z(n1974) );
  AND U2215 ( .A(n1975), .B(n1974), .Z(n2057) );
  NAND U2216 ( .A(n41), .B(n1976), .Z(n1978) );
  XOR U2217 ( .A(b[9]), .B(a[25]), .Z(n2053) );
  NAND U2218 ( .A(n4810), .B(n2053), .Z(n1977) );
  NAND U2219 ( .A(n1978), .B(n1977), .Z(n2056) );
  XOR U2220 ( .A(n2057), .B(n2056), .Z(n2059) );
  XOR U2221 ( .A(n2058), .B(n2059), .Z(n2069) );
  NANDN U2222 ( .A(n1980), .B(n1979), .Z(n1984) );
  OR U2223 ( .A(n1982), .B(n1981), .Z(n1983) );
  AND U2224 ( .A(n1984), .B(n1983), .Z(n2068) );
  XNOR U2225 ( .A(n2069), .B(n2068), .Z(n2070) );
  NANDN U2226 ( .A(n1986), .B(n1985), .Z(n1990) );
  NANDN U2227 ( .A(n1988), .B(n1987), .Z(n1989) );
  NAND U2228 ( .A(n1990), .B(n1989), .Z(n2071) );
  XNOR U2229 ( .A(n2070), .B(n2071), .Z(n2016) );
  XOR U2230 ( .A(n2017), .B(n2016), .Z(n2075) );
  NANDN U2231 ( .A(n1992), .B(n1991), .Z(n1996) );
  NANDN U2232 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U2233 ( .A(n1996), .B(n1995), .Z(n2074) );
  XNOR U2234 ( .A(n2075), .B(n2074), .Z(n2076) );
  XOR U2235 ( .A(n2077), .B(n2076), .Z(n2009) );
  NANDN U2236 ( .A(n1998), .B(n1997), .Z(n2002) );
  NAND U2237 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2238 ( .A(n2002), .B(n2001), .Z(n2008) );
  XNOR U2239 ( .A(n2009), .B(n2008), .Z(n2010) );
  XNOR U2240 ( .A(n2011), .B(n2010), .Z(n2080) );
  XNOR U2241 ( .A(sreg[81]), .B(n2080), .Z(n2082) );
  NANDN U2242 ( .A(sreg[80]), .B(n2003), .Z(n2007) );
  NAND U2243 ( .A(n2005), .B(n2004), .Z(n2006) );
  NAND U2244 ( .A(n2007), .B(n2006), .Z(n2081) );
  XNOR U2245 ( .A(n2082), .B(n2081), .Z(c[81]) );
  NANDN U2246 ( .A(n2009), .B(n2008), .Z(n2013) );
  NANDN U2247 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2248 ( .A(n2013), .B(n2012), .Z(n2088) );
  NANDN U2249 ( .A(n2015), .B(n2014), .Z(n2019) );
  NAND U2250 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U2251 ( .A(n2019), .B(n2018), .Z(n2154) );
  NANDN U2252 ( .A(n2021), .B(n2020), .Z(n2025) );
  NANDN U2253 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2254 ( .A(n2025), .B(n2024), .Z(n2120) );
  NAND U2255 ( .A(b[0]), .B(a[34]), .Z(n2026) );
  XNOR U2256 ( .A(b[1]), .B(n2026), .Z(n2028) );
  NANDN U2257 ( .A(b[0]), .B(a[33]), .Z(n2027) );
  NAND U2258 ( .A(n2028), .B(n2027), .Z(n2100) );
  NAND U2259 ( .A(n5012), .B(n2029), .Z(n2031) );
  XOR U2260 ( .A(b[13]), .B(a[22]), .Z(n2106) );
  NAND U2261 ( .A(n4985), .B(n2106), .Z(n2030) );
  AND U2262 ( .A(n2031), .B(n2030), .Z(n2098) );
  AND U2263 ( .A(b[15]), .B(a[18]), .Z(n2097) );
  XNOR U2264 ( .A(n2098), .B(n2097), .Z(n2099) );
  XNOR U2265 ( .A(n2100), .B(n2099), .Z(n2118) );
  NAND U2266 ( .A(n36), .B(n2032), .Z(n2034) );
  XOR U2267 ( .A(b[5]), .B(a[30]), .Z(n2109) );
  NAND U2268 ( .A(n4560), .B(n2109), .Z(n2033) );
  AND U2269 ( .A(n2034), .B(n2033), .Z(n2142) );
  NAND U2270 ( .A(n4755), .B(n2035), .Z(n2037) );
  XOR U2271 ( .A(b[7]), .B(a[28]), .Z(n2112) );
  NAND U2272 ( .A(n4708), .B(n2112), .Z(n2036) );
  AND U2273 ( .A(n2037), .B(n2036), .Z(n2140) );
  NAND U2274 ( .A(n4471), .B(n2038), .Z(n2040) );
  XOR U2275 ( .A(b[3]), .B(a[32]), .Z(n2115) );
  NAND U2276 ( .A(n33), .B(n2115), .Z(n2039) );
  NAND U2277 ( .A(n2040), .B(n2039), .Z(n2139) );
  XNOR U2278 ( .A(n2140), .B(n2139), .Z(n2141) );
  XOR U2279 ( .A(n2142), .B(n2141), .Z(n2119) );
  XOR U2280 ( .A(n2118), .B(n2119), .Z(n2121) );
  XOR U2281 ( .A(n2120), .B(n2121), .Z(n2092) );
  NANDN U2282 ( .A(n2042), .B(n2041), .Z(n2046) );
  OR U2283 ( .A(n2044), .B(n2043), .Z(n2045) );
  AND U2284 ( .A(n2046), .B(n2045), .Z(n2091) );
  XNOR U2285 ( .A(n2092), .B(n2091), .Z(n2094) );
  NAND U2286 ( .A(n4950), .B(n2047), .Z(n2049) );
  XOR U2287 ( .A(b[11]), .B(a[24]), .Z(n2124) );
  NAND U2288 ( .A(n4863), .B(n2124), .Z(n2048) );
  AND U2289 ( .A(n2049), .B(n2048), .Z(n2135) );
  NAND U2290 ( .A(n42), .B(n2050), .Z(n2052) );
  XOR U2291 ( .A(b[15]), .B(a[20]), .Z(n2127) );
  NAND U2292 ( .A(n4981), .B(n2127), .Z(n2051) );
  AND U2293 ( .A(n2052), .B(n2051), .Z(n2134) );
  NAND U2294 ( .A(n41), .B(n2053), .Z(n2055) );
  XOR U2295 ( .A(b[9]), .B(a[26]), .Z(n2130) );
  NAND U2296 ( .A(n4810), .B(n2130), .Z(n2054) );
  NAND U2297 ( .A(n2055), .B(n2054), .Z(n2133) );
  XOR U2298 ( .A(n2134), .B(n2133), .Z(n2136) );
  XOR U2299 ( .A(n2135), .B(n2136), .Z(n2146) );
  NANDN U2300 ( .A(n2057), .B(n2056), .Z(n2061) );
  OR U2301 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2302 ( .A(n2061), .B(n2060), .Z(n2145) );
  XNOR U2303 ( .A(n2146), .B(n2145), .Z(n2147) );
  NANDN U2304 ( .A(n2063), .B(n2062), .Z(n2067) );
  NANDN U2305 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U2306 ( .A(n2067), .B(n2066), .Z(n2148) );
  XNOR U2307 ( .A(n2147), .B(n2148), .Z(n2093) );
  XOR U2308 ( .A(n2094), .B(n2093), .Z(n2152) );
  NANDN U2309 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U2310 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2311 ( .A(n2073), .B(n2072), .Z(n2151) );
  XNOR U2312 ( .A(n2152), .B(n2151), .Z(n2153) );
  XOR U2313 ( .A(n2154), .B(n2153), .Z(n2086) );
  NANDN U2314 ( .A(n2075), .B(n2074), .Z(n2079) );
  NAND U2315 ( .A(n2077), .B(n2076), .Z(n2078) );
  AND U2316 ( .A(n2079), .B(n2078), .Z(n2085) );
  XNOR U2317 ( .A(n2086), .B(n2085), .Z(n2087) );
  XNOR U2318 ( .A(n2088), .B(n2087), .Z(n2157) );
  XNOR U2319 ( .A(sreg[82]), .B(n2157), .Z(n2159) );
  NANDN U2320 ( .A(sreg[81]), .B(n2080), .Z(n2084) );
  NAND U2321 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2322 ( .A(n2084), .B(n2083), .Z(n2158) );
  XNOR U2323 ( .A(n2159), .B(n2158), .Z(c[82]) );
  NANDN U2324 ( .A(n2086), .B(n2085), .Z(n2090) );
  NANDN U2325 ( .A(n2088), .B(n2087), .Z(n2089) );
  AND U2326 ( .A(n2090), .B(n2089), .Z(n2165) );
  NANDN U2327 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U2328 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U2329 ( .A(n2096), .B(n2095), .Z(n2231) );
  NANDN U2330 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U2331 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2332 ( .A(n2102), .B(n2101), .Z(n2197) );
  NAND U2333 ( .A(b[0]), .B(a[35]), .Z(n2103) );
  XNOR U2334 ( .A(b[1]), .B(n2103), .Z(n2105) );
  NANDN U2335 ( .A(b[0]), .B(a[34]), .Z(n2104) );
  NAND U2336 ( .A(n2105), .B(n2104), .Z(n2177) );
  NAND U2337 ( .A(n5012), .B(n2106), .Z(n2108) );
  XOR U2338 ( .A(b[13]), .B(a[23]), .Z(n2183) );
  NAND U2339 ( .A(n4985), .B(n2183), .Z(n2107) );
  AND U2340 ( .A(n2108), .B(n2107), .Z(n2175) );
  AND U2341 ( .A(b[15]), .B(a[19]), .Z(n2174) );
  XNOR U2342 ( .A(n2175), .B(n2174), .Z(n2176) );
  XNOR U2343 ( .A(n2177), .B(n2176), .Z(n2195) );
  NAND U2344 ( .A(n36), .B(n2109), .Z(n2111) );
  XOR U2345 ( .A(b[5]), .B(a[31]), .Z(n2186) );
  NAND U2346 ( .A(n4560), .B(n2186), .Z(n2110) );
  AND U2347 ( .A(n2111), .B(n2110), .Z(n2219) );
  NAND U2348 ( .A(n4755), .B(n2112), .Z(n2114) );
  XOR U2349 ( .A(b[7]), .B(a[29]), .Z(n2189) );
  NAND U2350 ( .A(n4708), .B(n2189), .Z(n2113) );
  AND U2351 ( .A(n2114), .B(n2113), .Z(n2217) );
  NAND U2352 ( .A(n4471), .B(n2115), .Z(n2117) );
  XOR U2353 ( .A(b[3]), .B(a[33]), .Z(n2192) );
  NAND U2354 ( .A(n33), .B(n2192), .Z(n2116) );
  NAND U2355 ( .A(n2117), .B(n2116), .Z(n2216) );
  XNOR U2356 ( .A(n2217), .B(n2216), .Z(n2218) );
  XOR U2357 ( .A(n2219), .B(n2218), .Z(n2196) );
  XOR U2358 ( .A(n2195), .B(n2196), .Z(n2198) );
  XOR U2359 ( .A(n2197), .B(n2198), .Z(n2169) );
  NANDN U2360 ( .A(n2119), .B(n2118), .Z(n2123) );
  OR U2361 ( .A(n2121), .B(n2120), .Z(n2122) );
  AND U2362 ( .A(n2123), .B(n2122), .Z(n2168) );
  XNOR U2363 ( .A(n2169), .B(n2168), .Z(n2171) );
  NAND U2364 ( .A(n4950), .B(n2124), .Z(n2126) );
  XOR U2365 ( .A(b[11]), .B(a[25]), .Z(n2201) );
  NAND U2366 ( .A(n4863), .B(n2201), .Z(n2125) );
  AND U2367 ( .A(n2126), .B(n2125), .Z(n2212) );
  NAND U2368 ( .A(n42), .B(n2127), .Z(n2129) );
  XOR U2369 ( .A(b[15]), .B(a[21]), .Z(n2204) );
  NAND U2370 ( .A(n4981), .B(n2204), .Z(n2128) );
  AND U2371 ( .A(n2129), .B(n2128), .Z(n2211) );
  NAND U2372 ( .A(n41), .B(n2130), .Z(n2132) );
  XOR U2373 ( .A(b[9]), .B(a[27]), .Z(n2207) );
  NAND U2374 ( .A(n4810), .B(n2207), .Z(n2131) );
  NAND U2375 ( .A(n2132), .B(n2131), .Z(n2210) );
  XOR U2376 ( .A(n2211), .B(n2210), .Z(n2213) );
  XOR U2377 ( .A(n2212), .B(n2213), .Z(n2223) );
  NANDN U2378 ( .A(n2134), .B(n2133), .Z(n2138) );
  OR U2379 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U2380 ( .A(n2138), .B(n2137), .Z(n2222) );
  XNOR U2381 ( .A(n2223), .B(n2222), .Z(n2224) );
  NANDN U2382 ( .A(n2140), .B(n2139), .Z(n2144) );
  NANDN U2383 ( .A(n2142), .B(n2141), .Z(n2143) );
  NAND U2384 ( .A(n2144), .B(n2143), .Z(n2225) );
  XNOR U2385 ( .A(n2224), .B(n2225), .Z(n2170) );
  XOR U2386 ( .A(n2171), .B(n2170), .Z(n2229) );
  NANDN U2387 ( .A(n2146), .B(n2145), .Z(n2150) );
  NANDN U2388 ( .A(n2148), .B(n2147), .Z(n2149) );
  AND U2389 ( .A(n2150), .B(n2149), .Z(n2228) );
  XNOR U2390 ( .A(n2229), .B(n2228), .Z(n2230) );
  XOR U2391 ( .A(n2231), .B(n2230), .Z(n2163) );
  NANDN U2392 ( .A(n2152), .B(n2151), .Z(n2156) );
  NAND U2393 ( .A(n2154), .B(n2153), .Z(n2155) );
  AND U2394 ( .A(n2156), .B(n2155), .Z(n2162) );
  XNOR U2395 ( .A(n2163), .B(n2162), .Z(n2164) );
  XNOR U2396 ( .A(n2165), .B(n2164), .Z(n2234) );
  XNOR U2397 ( .A(sreg[83]), .B(n2234), .Z(n2236) );
  NANDN U2398 ( .A(sreg[82]), .B(n2157), .Z(n2161) );
  NAND U2399 ( .A(n2159), .B(n2158), .Z(n2160) );
  NAND U2400 ( .A(n2161), .B(n2160), .Z(n2235) );
  XNOR U2401 ( .A(n2236), .B(n2235), .Z(c[83]) );
  NANDN U2402 ( .A(n2163), .B(n2162), .Z(n2167) );
  NANDN U2403 ( .A(n2165), .B(n2164), .Z(n2166) );
  AND U2404 ( .A(n2167), .B(n2166), .Z(n2242) );
  NANDN U2405 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2406 ( .A(n2171), .B(n2170), .Z(n2172) );
  AND U2407 ( .A(n2173), .B(n2172), .Z(n2308) );
  NANDN U2408 ( .A(n2175), .B(n2174), .Z(n2179) );
  NANDN U2409 ( .A(n2177), .B(n2176), .Z(n2178) );
  AND U2410 ( .A(n2179), .B(n2178), .Z(n2274) );
  NAND U2411 ( .A(b[0]), .B(a[36]), .Z(n2180) );
  XNOR U2412 ( .A(b[1]), .B(n2180), .Z(n2182) );
  NANDN U2413 ( .A(b[0]), .B(a[35]), .Z(n2181) );
  NAND U2414 ( .A(n2182), .B(n2181), .Z(n2254) );
  NAND U2415 ( .A(n5012), .B(n2183), .Z(n2185) );
  XOR U2416 ( .A(b[13]), .B(a[24]), .Z(n2260) );
  NAND U2417 ( .A(n4985), .B(n2260), .Z(n2184) );
  AND U2418 ( .A(n2185), .B(n2184), .Z(n2252) );
  AND U2419 ( .A(b[15]), .B(a[20]), .Z(n2251) );
  XNOR U2420 ( .A(n2252), .B(n2251), .Z(n2253) );
  XNOR U2421 ( .A(n2254), .B(n2253), .Z(n2272) );
  NAND U2422 ( .A(n36), .B(n2186), .Z(n2188) );
  XOR U2423 ( .A(b[5]), .B(a[32]), .Z(n2263) );
  NAND U2424 ( .A(n4560), .B(n2263), .Z(n2187) );
  AND U2425 ( .A(n2188), .B(n2187), .Z(n2296) );
  NAND U2426 ( .A(n4755), .B(n2189), .Z(n2191) );
  XOR U2427 ( .A(b[7]), .B(a[30]), .Z(n2266) );
  NAND U2428 ( .A(n4708), .B(n2266), .Z(n2190) );
  AND U2429 ( .A(n2191), .B(n2190), .Z(n2294) );
  NAND U2430 ( .A(n4471), .B(n2192), .Z(n2194) );
  XOR U2431 ( .A(b[3]), .B(a[34]), .Z(n2269) );
  NAND U2432 ( .A(n33), .B(n2269), .Z(n2193) );
  NAND U2433 ( .A(n2194), .B(n2193), .Z(n2293) );
  XNOR U2434 ( .A(n2294), .B(n2293), .Z(n2295) );
  XOR U2435 ( .A(n2296), .B(n2295), .Z(n2273) );
  XOR U2436 ( .A(n2272), .B(n2273), .Z(n2275) );
  XOR U2437 ( .A(n2274), .B(n2275), .Z(n2246) );
  NANDN U2438 ( .A(n2196), .B(n2195), .Z(n2200) );
  OR U2439 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U2440 ( .A(n2200), .B(n2199), .Z(n2245) );
  XNOR U2441 ( .A(n2246), .B(n2245), .Z(n2248) );
  NAND U2442 ( .A(n4950), .B(n2201), .Z(n2203) );
  XOR U2443 ( .A(b[11]), .B(a[26]), .Z(n2278) );
  NAND U2444 ( .A(n4863), .B(n2278), .Z(n2202) );
  AND U2445 ( .A(n2203), .B(n2202), .Z(n2289) );
  NAND U2446 ( .A(n42), .B(n2204), .Z(n2206) );
  XOR U2447 ( .A(b[15]), .B(a[22]), .Z(n2281) );
  NAND U2448 ( .A(n4981), .B(n2281), .Z(n2205) );
  AND U2449 ( .A(n2206), .B(n2205), .Z(n2288) );
  NAND U2450 ( .A(n41), .B(n2207), .Z(n2209) );
  XOR U2451 ( .A(b[9]), .B(a[28]), .Z(n2284) );
  NAND U2452 ( .A(n4810), .B(n2284), .Z(n2208) );
  NAND U2453 ( .A(n2209), .B(n2208), .Z(n2287) );
  XOR U2454 ( .A(n2288), .B(n2287), .Z(n2290) );
  XOR U2455 ( .A(n2289), .B(n2290), .Z(n2300) );
  NANDN U2456 ( .A(n2211), .B(n2210), .Z(n2215) );
  OR U2457 ( .A(n2213), .B(n2212), .Z(n2214) );
  AND U2458 ( .A(n2215), .B(n2214), .Z(n2299) );
  XNOR U2459 ( .A(n2300), .B(n2299), .Z(n2301) );
  NANDN U2460 ( .A(n2217), .B(n2216), .Z(n2221) );
  NANDN U2461 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2462 ( .A(n2221), .B(n2220), .Z(n2302) );
  XNOR U2463 ( .A(n2301), .B(n2302), .Z(n2247) );
  XOR U2464 ( .A(n2248), .B(n2247), .Z(n2306) );
  NANDN U2465 ( .A(n2223), .B(n2222), .Z(n2227) );
  NANDN U2466 ( .A(n2225), .B(n2224), .Z(n2226) );
  AND U2467 ( .A(n2227), .B(n2226), .Z(n2305) );
  XNOR U2468 ( .A(n2306), .B(n2305), .Z(n2307) );
  XOR U2469 ( .A(n2308), .B(n2307), .Z(n2240) );
  NANDN U2470 ( .A(n2229), .B(n2228), .Z(n2233) );
  NAND U2471 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U2472 ( .A(n2233), .B(n2232), .Z(n2239) );
  XNOR U2473 ( .A(n2240), .B(n2239), .Z(n2241) );
  XNOR U2474 ( .A(n2242), .B(n2241), .Z(n2311) );
  XNOR U2475 ( .A(sreg[84]), .B(n2311), .Z(n2313) );
  NANDN U2476 ( .A(sreg[83]), .B(n2234), .Z(n2238) );
  NAND U2477 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2478 ( .A(n2238), .B(n2237), .Z(n2312) );
  XNOR U2479 ( .A(n2313), .B(n2312), .Z(c[84]) );
  NANDN U2480 ( .A(n2240), .B(n2239), .Z(n2244) );
  NANDN U2481 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2482 ( .A(n2244), .B(n2243), .Z(n2319) );
  NANDN U2483 ( .A(n2246), .B(n2245), .Z(n2250) );
  NAND U2484 ( .A(n2248), .B(n2247), .Z(n2249) );
  AND U2485 ( .A(n2250), .B(n2249), .Z(n2385) );
  NANDN U2486 ( .A(n2252), .B(n2251), .Z(n2256) );
  NANDN U2487 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2488 ( .A(n2256), .B(n2255), .Z(n2351) );
  NAND U2489 ( .A(b[0]), .B(a[37]), .Z(n2257) );
  XNOR U2490 ( .A(b[1]), .B(n2257), .Z(n2259) );
  NANDN U2491 ( .A(b[0]), .B(a[36]), .Z(n2258) );
  NAND U2492 ( .A(n2259), .B(n2258), .Z(n2331) );
  NAND U2493 ( .A(n5012), .B(n2260), .Z(n2262) );
  XOR U2494 ( .A(b[13]), .B(a[25]), .Z(n2334) );
  NAND U2495 ( .A(n4985), .B(n2334), .Z(n2261) );
  AND U2496 ( .A(n2262), .B(n2261), .Z(n2329) );
  AND U2497 ( .A(b[15]), .B(a[21]), .Z(n2328) );
  XNOR U2498 ( .A(n2329), .B(n2328), .Z(n2330) );
  XNOR U2499 ( .A(n2331), .B(n2330), .Z(n2349) );
  NAND U2500 ( .A(n36), .B(n2263), .Z(n2265) );
  XOR U2501 ( .A(b[5]), .B(a[33]), .Z(n2340) );
  NAND U2502 ( .A(n4560), .B(n2340), .Z(n2264) );
  AND U2503 ( .A(n2265), .B(n2264), .Z(n2373) );
  NAND U2504 ( .A(n4755), .B(n2266), .Z(n2268) );
  XOR U2505 ( .A(b[7]), .B(a[31]), .Z(n2343) );
  NAND U2506 ( .A(n4708), .B(n2343), .Z(n2267) );
  AND U2507 ( .A(n2268), .B(n2267), .Z(n2371) );
  NAND U2508 ( .A(n4471), .B(n2269), .Z(n2271) );
  XOR U2509 ( .A(b[3]), .B(a[35]), .Z(n2346) );
  NAND U2510 ( .A(n33), .B(n2346), .Z(n2270) );
  NAND U2511 ( .A(n2271), .B(n2270), .Z(n2370) );
  XNOR U2512 ( .A(n2371), .B(n2370), .Z(n2372) );
  XOR U2513 ( .A(n2373), .B(n2372), .Z(n2350) );
  XOR U2514 ( .A(n2349), .B(n2350), .Z(n2352) );
  XOR U2515 ( .A(n2351), .B(n2352), .Z(n2323) );
  NANDN U2516 ( .A(n2273), .B(n2272), .Z(n2277) );
  OR U2517 ( .A(n2275), .B(n2274), .Z(n2276) );
  AND U2518 ( .A(n2277), .B(n2276), .Z(n2322) );
  XNOR U2519 ( .A(n2323), .B(n2322), .Z(n2325) );
  NAND U2520 ( .A(n4950), .B(n2278), .Z(n2280) );
  XOR U2521 ( .A(b[11]), .B(a[27]), .Z(n2355) );
  NAND U2522 ( .A(n4863), .B(n2355), .Z(n2279) );
  AND U2523 ( .A(n2280), .B(n2279), .Z(n2366) );
  NAND U2524 ( .A(n42), .B(n2281), .Z(n2283) );
  XOR U2525 ( .A(b[15]), .B(a[23]), .Z(n2358) );
  NAND U2526 ( .A(n4981), .B(n2358), .Z(n2282) );
  AND U2527 ( .A(n2283), .B(n2282), .Z(n2365) );
  NAND U2528 ( .A(n41), .B(n2284), .Z(n2286) );
  XOR U2529 ( .A(b[9]), .B(a[29]), .Z(n2361) );
  NAND U2530 ( .A(n4810), .B(n2361), .Z(n2285) );
  NAND U2531 ( .A(n2286), .B(n2285), .Z(n2364) );
  XOR U2532 ( .A(n2365), .B(n2364), .Z(n2367) );
  XOR U2533 ( .A(n2366), .B(n2367), .Z(n2377) );
  NANDN U2534 ( .A(n2288), .B(n2287), .Z(n2292) );
  OR U2535 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U2536 ( .A(n2292), .B(n2291), .Z(n2376) );
  XNOR U2537 ( .A(n2377), .B(n2376), .Z(n2378) );
  NANDN U2538 ( .A(n2294), .B(n2293), .Z(n2298) );
  NANDN U2539 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2540 ( .A(n2298), .B(n2297), .Z(n2379) );
  XNOR U2541 ( .A(n2378), .B(n2379), .Z(n2324) );
  XOR U2542 ( .A(n2325), .B(n2324), .Z(n2383) );
  NANDN U2543 ( .A(n2300), .B(n2299), .Z(n2304) );
  NANDN U2544 ( .A(n2302), .B(n2301), .Z(n2303) );
  AND U2545 ( .A(n2304), .B(n2303), .Z(n2382) );
  XNOR U2546 ( .A(n2383), .B(n2382), .Z(n2384) );
  XOR U2547 ( .A(n2385), .B(n2384), .Z(n2317) );
  NANDN U2548 ( .A(n2306), .B(n2305), .Z(n2310) );
  NAND U2549 ( .A(n2308), .B(n2307), .Z(n2309) );
  AND U2550 ( .A(n2310), .B(n2309), .Z(n2316) );
  XNOR U2551 ( .A(n2317), .B(n2316), .Z(n2318) );
  XNOR U2552 ( .A(n2319), .B(n2318), .Z(n2388) );
  XNOR U2553 ( .A(sreg[85]), .B(n2388), .Z(n2390) );
  NANDN U2554 ( .A(sreg[84]), .B(n2311), .Z(n2315) );
  NAND U2555 ( .A(n2313), .B(n2312), .Z(n2314) );
  NAND U2556 ( .A(n2315), .B(n2314), .Z(n2389) );
  XNOR U2557 ( .A(n2390), .B(n2389), .Z(c[85]) );
  NANDN U2558 ( .A(n2317), .B(n2316), .Z(n2321) );
  NANDN U2559 ( .A(n2319), .B(n2318), .Z(n2320) );
  AND U2560 ( .A(n2321), .B(n2320), .Z(n2396) );
  NANDN U2561 ( .A(n2323), .B(n2322), .Z(n2327) );
  NAND U2562 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2563 ( .A(n2327), .B(n2326), .Z(n2462) );
  NANDN U2564 ( .A(n2329), .B(n2328), .Z(n2333) );
  NANDN U2565 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U2566 ( .A(n2333), .B(n2332), .Z(n2428) );
  NAND U2567 ( .A(n5012), .B(n2334), .Z(n2336) );
  XOR U2568 ( .A(b[13]), .B(a[26]), .Z(n2414) );
  NAND U2569 ( .A(n4985), .B(n2414), .Z(n2335) );
  AND U2570 ( .A(n2336), .B(n2335), .Z(n2406) );
  AND U2571 ( .A(b[15]), .B(a[22]), .Z(n2405) );
  XNOR U2572 ( .A(n2406), .B(n2405), .Z(n2407) );
  NAND U2573 ( .A(b[0]), .B(a[38]), .Z(n2337) );
  XNOR U2574 ( .A(b[1]), .B(n2337), .Z(n2339) );
  NANDN U2575 ( .A(b[0]), .B(a[37]), .Z(n2338) );
  NAND U2576 ( .A(n2339), .B(n2338), .Z(n2408) );
  XNOR U2577 ( .A(n2407), .B(n2408), .Z(n2426) );
  NAND U2578 ( .A(n36), .B(n2340), .Z(n2342) );
  XOR U2579 ( .A(b[5]), .B(a[34]), .Z(n2417) );
  NAND U2580 ( .A(n4560), .B(n2417), .Z(n2341) );
  AND U2581 ( .A(n2342), .B(n2341), .Z(n2450) );
  NAND U2582 ( .A(n4755), .B(n2343), .Z(n2345) );
  XOR U2583 ( .A(b[7]), .B(a[32]), .Z(n2420) );
  NAND U2584 ( .A(n4708), .B(n2420), .Z(n2344) );
  AND U2585 ( .A(n2345), .B(n2344), .Z(n2448) );
  NAND U2586 ( .A(n4471), .B(n2346), .Z(n2348) );
  XOR U2587 ( .A(b[3]), .B(a[36]), .Z(n2423) );
  NAND U2588 ( .A(n33), .B(n2423), .Z(n2347) );
  NAND U2589 ( .A(n2348), .B(n2347), .Z(n2447) );
  XNOR U2590 ( .A(n2448), .B(n2447), .Z(n2449) );
  XOR U2591 ( .A(n2450), .B(n2449), .Z(n2427) );
  XOR U2592 ( .A(n2426), .B(n2427), .Z(n2429) );
  XOR U2593 ( .A(n2428), .B(n2429), .Z(n2400) );
  NANDN U2594 ( .A(n2350), .B(n2349), .Z(n2354) );
  OR U2595 ( .A(n2352), .B(n2351), .Z(n2353) );
  AND U2596 ( .A(n2354), .B(n2353), .Z(n2399) );
  XNOR U2597 ( .A(n2400), .B(n2399), .Z(n2402) );
  NAND U2598 ( .A(n4950), .B(n2355), .Z(n2357) );
  XOR U2599 ( .A(b[11]), .B(a[28]), .Z(n2432) );
  NAND U2600 ( .A(n4863), .B(n2432), .Z(n2356) );
  AND U2601 ( .A(n2357), .B(n2356), .Z(n2443) );
  NAND U2602 ( .A(n42), .B(n2358), .Z(n2360) );
  XOR U2603 ( .A(b[15]), .B(a[24]), .Z(n2435) );
  NAND U2604 ( .A(n4981), .B(n2435), .Z(n2359) );
  AND U2605 ( .A(n2360), .B(n2359), .Z(n2442) );
  NAND U2606 ( .A(n41), .B(n2361), .Z(n2363) );
  XOR U2607 ( .A(b[9]), .B(a[30]), .Z(n2438) );
  NAND U2608 ( .A(n4810), .B(n2438), .Z(n2362) );
  NAND U2609 ( .A(n2363), .B(n2362), .Z(n2441) );
  XOR U2610 ( .A(n2442), .B(n2441), .Z(n2444) );
  XOR U2611 ( .A(n2443), .B(n2444), .Z(n2454) );
  NANDN U2612 ( .A(n2365), .B(n2364), .Z(n2369) );
  OR U2613 ( .A(n2367), .B(n2366), .Z(n2368) );
  AND U2614 ( .A(n2369), .B(n2368), .Z(n2453) );
  XNOR U2615 ( .A(n2454), .B(n2453), .Z(n2455) );
  NANDN U2616 ( .A(n2371), .B(n2370), .Z(n2375) );
  NANDN U2617 ( .A(n2373), .B(n2372), .Z(n2374) );
  NAND U2618 ( .A(n2375), .B(n2374), .Z(n2456) );
  XNOR U2619 ( .A(n2455), .B(n2456), .Z(n2401) );
  XOR U2620 ( .A(n2402), .B(n2401), .Z(n2460) );
  NANDN U2621 ( .A(n2377), .B(n2376), .Z(n2381) );
  NANDN U2622 ( .A(n2379), .B(n2378), .Z(n2380) );
  AND U2623 ( .A(n2381), .B(n2380), .Z(n2459) );
  XNOR U2624 ( .A(n2460), .B(n2459), .Z(n2461) );
  XOR U2625 ( .A(n2462), .B(n2461), .Z(n2394) );
  NANDN U2626 ( .A(n2383), .B(n2382), .Z(n2387) );
  NAND U2627 ( .A(n2385), .B(n2384), .Z(n2386) );
  AND U2628 ( .A(n2387), .B(n2386), .Z(n2393) );
  XNOR U2629 ( .A(n2394), .B(n2393), .Z(n2395) );
  XNOR U2630 ( .A(n2396), .B(n2395), .Z(n2465) );
  XNOR U2631 ( .A(sreg[86]), .B(n2465), .Z(n2467) );
  NANDN U2632 ( .A(sreg[85]), .B(n2388), .Z(n2392) );
  NAND U2633 ( .A(n2390), .B(n2389), .Z(n2391) );
  NAND U2634 ( .A(n2392), .B(n2391), .Z(n2466) );
  XNOR U2635 ( .A(n2467), .B(n2466), .Z(c[86]) );
  NANDN U2636 ( .A(n2394), .B(n2393), .Z(n2398) );
  NANDN U2637 ( .A(n2396), .B(n2395), .Z(n2397) );
  AND U2638 ( .A(n2398), .B(n2397), .Z(n2473) );
  NANDN U2639 ( .A(n2400), .B(n2399), .Z(n2404) );
  NAND U2640 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U2641 ( .A(n2404), .B(n2403), .Z(n2539) );
  NANDN U2642 ( .A(n2406), .B(n2405), .Z(n2410) );
  NANDN U2643 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U2644 ( .A(n2410), .B(n2409), .Z(n2505) );
  NAND U2645 ( .A(b[0]), .B(a[39]), .Z(n2411) );
  XNOR U2646 ( .A(b[1]), .B(n2411), .Z(n2413) );
  NANDN U2647 ( .A(b[0]), .B(a[38]), .Z(n2412) );
  NAND U2648 ( .A(n2413), .B(n2412), .Z(n2485) );
  NAND U2649 ( .A(n5012), .B(n2414), .Z(n2416) );
  XOR U2650 ( .A(b[13]), .B(a[27]), .Z(n2491) );
  NAND U2651 ( .A(n4985), .B(n2491), .Z(n2415) );
  AND U2652 ( .A(n2416), .B(n2415), .Z(n2483) );
  AND U2653 ( .A(b[15]), .B(a[23]), .Z(n2482) );
  XNOR U2654 ( .A(n2483), .B(n2482), .Z(n2484) );
  XNOR U2655 ( .A(n2485), .B(n2484), .Z(n2503) );
  NAND U2656 ( .A(n36), .B(n2417), .Z(n2419) );
  XOR U2657 ( .A(b[5]), .B(a[35]), .Z(n2494) );
  NAND U2658 ( .A(n4560), .B(n2494), .Z(n2418) );
  AND U2659 ( .A(n2419), .B(n2418), .Z(n2527) );
  NAND U2660 ( .A(n4755), .B(n2420), .Z(n2422) );
  XOR U2661 ( .A(b[7]), .B(a[33]), .Z(n2497) );
  NAND U2662 ( .A(n4708), .B(n2497), .Z(n2421) );
  AND U2663 ( .A(n2422), .B(n2421), .Z(n2525) );
  NAND U2664 ( .A(n4471), .B(n2423), .Z(n2425) );
  XOR U2665 ( .A(b[3]), .B(a[37]), .Z(n2500) );
  NAND U2666 ( .A(n33), .B(n2500), .Z(n2424) );
  NAND U2667 ( .A(n2425), .B(n2424), .Z(n2524) );
  XNOR U2668 ( .A(n2525), .B(n2524), .Z(n2526) );
  XOR U2669 ( .A(n2527), .B(n2526), .Z(n2504) );
  XOR U2670 ( .A(n2503), .B(n2504), .Z(n2506) );
  XOR U2671 ( .A(n2505), .B(n2506), .Z(n2477) );
  NANDN U2672 ( .A(n2427), .B(n2426), .Z(n2431) );
  OR U2673 ( .A(n2429), .B(n2428), .Z(n2430) );
  AND U2674 ( .A(n2431), .B(n2430), .Z(n2476) );
  XNOR U2675 ( .A(n2477), .B(n2476), .Z(n2479) );
  NAND U2676 ( .A(n4950), .B(n2432), .Z(n2434) );
  XOR U2677 ( .A(b[11]), .B(a[29]), .Z(n2509) );
  NAND U2678 ( .A(n4863), .B(n2509), .Z(n2433) );
  AND U2679 ( .A(n2434), .B(n2433), .Z(n2520) );
  NAND U2680 ( .A(n42), .B(n2435), .Z(n2437) );
  XOR U2681 ( .A(b[15]), .B(a[25]), .Z(n2512) );
  NAND U2682 ( .A(n4981), .B(n2512), .Z(n2436) );
  AND U2683 ( .A(n2437), .B(n2436), .Z(n2519) );
  NAND U2684 ( .A(n41), .B(n2438), .Z(n2440) );
  XOR U2685 ( .A(b[9]), .B(a[31]), .Z(n2515) );
  NAND U2686 ( .A(n4810), .B(n2515), .Z(n2439) );
  NAND U2687 ( .A(n2440), .B(n2439), .Z(n2518) );
  XOR U2688 ( .A(n2519), .B(n2518), .Z(n2521) );
  XOR U2689 ( .A(n2520), .B(n2521), .Z(n2531) );
  NANDN U2690 ( .A(n2442), .B(n2441), .Z(n2446) );
  OR U2691 ( .A(n2444), .B(n2443), .Z(n2445) );
  AND U2692 ( .A(n2446), .B(n2445), .Z(n2530) );
  XNOR U2693 ( .A(n2531), .B(n2530), .Z(n2532) );
  NANDN U2694 ( .A(n2448), .B(n2447), .Z(n2452) );
  NANDN U2695 ( .A(n2450), .B(n2449), .Z(n2451) );
  NAND U2696 ( .A(n2452), .B(n2451), .Z(n2533) );
  XNOR U2697 ( .A(n2532), .B(n2533), .Z(n2478) );
  XOR U2698 ( .A(n2479), .B(n2478), .Z(n2537) );
  NANDN U2699 ( .A(n2454), .B(n2453), .Z(n2458) );
  NANDN U2700 ( .A(n2456), .B(n2455), .Z(n2457) );
  AND U2701 ( .A(n2458), .B(n2457), .Z(n2536) );
  XNOR U2702 ( .A(n2537), .B(n2536), .Z(n2538) );
  XOR U2703 ( .A(n2539), .B(n2538), .Z(n2471) );
  NANDN U2704 ( .A(n2460), .B(n2459), .Z(n2464) );
  NAND U2705 ( .A(n2462), .B(n2461), .Z(n2463) );
  AND U2706 ( .A(n2464), .B(n2463), .Z(n2470) );
  XNOR U2707 ( .A(n2471), .B(n2470), .Z(n2472) );
  XNOR U2708 ( .A(n2473), .B(n2472), .Z(n2542) );
  XNOR U2709 ( .A(sreg[87]), .B(n2542), .Z(n2544) );
  NANDN U2710 ( .A(sreg[86]), .B(n2465), .Z(n2469) );
  NAND U2711 ( .A(n2467), .B(n2466), .Z(n2468) );
  NAND U2712 ( .A(n2469), .B(n2468), .Z(n2543) );
  XNOR U2713 ( .A(n2544), .B(n2543), .Z(c[87]) );
  NANDN U2714 ( .A(n2471), .B(n2470), .Z(n2475) );
  NANDN U2715 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U2716 ( .A(n2475), .B(n2474), .Z(n2550) );
  NANDN U2717 ( .A(n2477), .B(n2476), .Z(n2481) );
  NAND U2718 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2719 ( .A(n2481), .B(n2480), .Z(n2616) );
  NANDN U2720 ( .A(n2483), .B(n2482), .Z(n2487) );
  NANDN U2721 ( .A(n2485), .B(n2484), .Z(n2486) );
  AND U2722 ( .A(n2487), .B(n2486), .Z(n2582) );
  NAND U2723 ( .A(b[0]), .B(a[40]), .Z(n2488) );
  XNOR U2724 ( .A(b[1]), .B(n2488), .Z(n2490) );
  NANDN U2725 ( .A(b[0]), .B(a[39]), .Z(n2489) );
  NAND U2726 ( .A(n2490), .B(n2489), .Z(n2562) );
  NAND U2727 ( .A(n5012), .B(n2491), .Z(n2493) );
  XOR U2728 ( .A(b[13]), .B(a[28]), .Z(n2568) );
  NAND U2729 ( .A(n4985), .B(n2568), .Z(n2492) );
  AND U2730 ( .A(n2493), .B(n2492), .Z(n2560) );
  AND U2731 ( .A(b[15]), .B(a[24]), .Z(n2559) );
  XNOR U2732 ( .A(n2560), .B(n2559), .Z(n2561) );
  XNOR U2733 ( .A(n2562), .B(n2561), .Z(n2580) );
  NAND U2734 ( .A(n36), .B(n2494), .Z(n2496) );
  XOR U2735 ( .A(b[5]), .B(a[36]), .Z(n2571) );
  NAND U2736 ( .A(n4560), .B(n2571), .Z(n2495) );
  AND U2737 ( .A(n2496), .B(n2495), .Z(n2604) );
  NAND U2738 ( .A(n4755), .B(n2497), .Z(n2499) );
  XOR U2739 ( .A(b[7]), .B(a[34]), .Z(n2574) );
  NAND U2740 ( .A(n4708), .B(n2574), .Z(n2498) );
  AND U2741 ( .A(n2499), .B(n2498), .Z(n2602) );
  NAND U2742 ( .A(n4471), .B(n2500), .Z(n2502) );
  XOR U2743 ( .A(b[3]), .B(a[38]), .Z(n2577) );
  NAND U2744 ( .A(n33), .B(n2577), .Z(n2501) );
  NAND U2745 ( .A(n2502), .B(n2501), .Z(n2601) );
  XNOR U2746 ( .A(n2602), .B(n2601), .Z(n2603) );
  XOR U2747 ( .A(n2604), .B(n2603), .Z(n2581) );
  XOR U2748 ( .A(n2580), .B(n2581), .Z(n2583) );
  XOR U2749 ( .A(n2582), .B(n2583), .Z(n2554) );
  NANDN U2750 ( .A(n2504), .B(n2503), .Z(n2508) );
  OR U2751 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U2752 ( .A(n2508), .B(n2507), .Z(n2553) );
  XNOR U2753 ( .A(n2554), .B(n2553), .Z(n2556) );
  NAND U2754 ( .A(n4950), .B(n2509), .Z(n2511) );
  XOR U2755 ( .A(b[11]), .B(a[30]), .Z(n2586) );
  NAND U2756 ( .A(n4863), .B(n2586), .Z(n2510) );
  AND U2757 ( .A(n2511), .B(n2510), .Z(n2597) );
  NAND U2758 ( .A(n42), .B(n2512), .Z(n2514) );
  XOR U2759 ( .A(b[15]), .B(a[26]), .Z(n2589) );
  NAND U2760 ( .A(n4981), .B(n2589), .Z(n2513) );
  AND U2761 ( .A(n2514), .B(n2513), .Z(n2596) );
  NAND U2762 ( .A(n41), .B(n2515), .Z(n2517) );
  XOR U2763 ( .A(b[9]), .B(a[32]), .Z(n2592) );
  NAND U2764 ( .A(n4810), .B(n2592), .Z(n2516) );
  NAND U2765 ( .A(n2517), .B(n2516), .Z(n2595) );
  XOR U2766 ( .A(n2596), .B(n2595), .Z(n2598) );
  XOR U2767 ( .A(n2597), .B(n2598), .Z(n2608) );
  NANDN U2768 ( .A(n2519), .B(n2518), .Z(n2523) );
  OR U2769 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U2770 ( .A(n2523), .B(n2522), .Z(n2607) );
  XNOR U2771 ( .A(n2608), .B(n2607), .Z(n2609) );
  NANDN U2772 ( .A(n2525), .B(n2524), .Z(n2529) );
  NANDN U2773 ( .A(n2527), .B(n2526), .Z(n2528) );
  NAND U2774 ( .A(n2529), .B(n2528), .Z(n2610) );
  XNOR U2775 ( .A(n2609), .B(n2610), .Z(n2555) );
  XOR U2776 ( .A(n2556), .B(n2555), .Z(n2614) );
  NANDN U2777 ( .A(n2531), .B(n2530), .Z(n2535) );
  NANDN U2778 ( .A(n2533), .B(n2532), .Z(n2534) );
  AND U2779 ( .A(n2535), .B(n2534), .Z(n2613) );
  XNOR U2780 ( .A(n2614), .B(n2613), .Z(n2615) );
  XOR U2781 ( .A(n2616), .B(n2615), .Z(n2548) );
  NANDN U2782 ( .A(n2537), .B(n2536), .Z(n2541) );
  NAND U2783 ( .A(n2539), .B(n2538), .Z(n2540) );
  AND U2784 ( .A(n2541), .B(n2540), .Z(n2547) );
  XNOR U2785 ( .A(n2548), .B(n2547), .Z(n2549) );
  XNOR U2786 ( .A(n2550), .B(n2549), .Z(n2619) );
  XNOR U2787 ( .A(sreg[88]), .B(n2619), .Z(n2621) );
  NANDN U2788 ( .A(sreg[87]), .B(n2542), .Z(n2546) );
  NAND U2789 ( .A(n2544), .B(n2543), .Z(n2545) );
  NAND U2790 ( .A(n2546), .B(n2545), .Z(n2620) );
  XNOR U2791 ( .A(n2621), .B(n2620), .Z(c[88]) );
  NANDN U2792 ( .A(n2548), .B(n2547), .Z(n2552) );
  NANDN U2793 ( .A(n2550), .B(n2549), .Z(n2551) );
  AND U2794 ( .A(n2552), .B(n2551), .Z(n2627) );
  NANDN U2795 ( .A(n2554), .B(n2553), .Z(n2558) );
  NAND U2796 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U2797 ( .A(n2558), .B(n2557), .Z(n2693) );
  NANDN U2798 ( .A(n2560), .B(n2559), .Z(n2564) );
  NANDN U2799 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2800 ( .A(n2564), .B(n2563), .Z(n2680) );
  NAND U2801 ( .A(b[0]), .B(a[41]), .Z(n2565) );
  XNOR U2802 ( .A(b[1]), .B(n2565), .Z(n2567) );
  NANDN U2803 ( .A(b[0]), .B(a[40]), .Z(n2566) );
  NAND U2804 ( .A(n2567), .B(n2566), .Z(n2660) );
  NAND U2805 ( .A(n5012), .B(n2568), .Z(n2570) );
  XOR U2806 ( .A(b[13]), .B(a[29]), .Z(n2666) );
  NAND U2807 ( .A(n4985), .B(n2666), .Z(n2569) );
  AND U2808 ( .A(n2570), .B(n2569), .Z(n2658) );
  AND U2809 ( .A(b[15]), .B(a[25]), .Z(n2657) );
  XNOR U2810 ( .A(n2658), .B(n2657), .Z(n2659) );
  XNOR U2811 ( .A(n2660), .B(n2659), .Z(n2678) );
  NAND U2812 ( .A(n36), .B(n2571), .Z(n2573) );
  XOR U2813 ( .A(b[5]), .B(a[37]), .Z(n2669) );
  NAND U2814 ( .A(n4560), .B(n2669), .Z(n2572) );
  AND U2815 ( .A(n2573), .B(n2572), .Z(n2654) );
  NAND U2816 ( .A(n4755), .B(n2574), .Z(n2576) );
  XOR U2817 ( .A(b[7]), .B(a[35]), .Z(n2672) );
  NAND U2818 ( .A(n4708), .B(n2672), .Z(n2575) );
  AND U2819 ( .A(n2576), .B(n2575), .Z(n2652) );
  NAND U2820 ( .A(n4471), .B(n2577), .Z(n2579) );
  XOR U2821 ( .A(b[3]), .B(a[39]), .Z(n2675) );
  NAND U2822 ( .A(n33), .B(n2675), .Z(n2578) );
  NAND U2823 ( .A(n2579), .B(n2578), .Z(n2651) );
  XNOR U2824 ( .A(n2652), .B(n2651), .Z(n2653) );
  XOR U2825 ( .A(n2654), .B(n2653), .Z(n2679) );
  XOR U2826 ( .A(n2678), .B(n2679), .Z(n2681) );
  XOR U2827 ( .A(n2680), .B(n2681), .Z(n2631) );
  NANDN U2828 ( .A(n2581), .B(n2580), .Z(n2585) );
  OR U2829 ( .A(n2583), .B(n2582), .Z(n2584) );
  AND U2830 ( .A(n2585), .B(n2584), .Z(n2630) );
  XNOR U2831 ( .A(n2631), .B(n2630), .Z(n2633) );
  NAND U2832 ( .A(n4950), .B(n2586), .Z(n2588) );
  XOR U2833 ( .A(b[11]), .B(a[31]), .Z(n2636) );
  NAND U2834 ( .A(n4863), .B(n2636), .Z(n2587) );
  AND U2835 ( .A(n2588), .B(n2587), .Z(n2647) );
  NAND U2836 ( .A(n42), .B(n2589), .Z(n2591) );
  XOR U2837 ( .A(b[15]), .B(a[27]), .Z(n2639) );
  NAND U2838 ( .A(n4981), .B(n2639), .Z(n2590) );
  AND U2839 ( .A(n2591), .B(n2590), .Z(n2646) );
  NAND U2840 ( .A(n41), .B(n2592), .Z(n2594) );
  XOR U2841 ( .A(b[9]), .B(a[33]), .Z(n2642) );
  NAND U2842 ( .A(n4810), .B(n2642), .Z(n2593) );
  NAND U2843 ( .A(n2594), .B(n2593), .Z(n2645) );
  XOR U2844 ( .A(n2646), .B(n2645), .Z(n2648) );
  XOR U2845 ( .A(n2647), .B(n2648), .Z(n2685) );
  NANDN U2846 ( .A(n2596), .B(n2595), .Z(n2600) );
  OR U2847 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U2848 ( .A(n2600), .B(n2599), .Z(n2684) );
  XNOR U2849 ( .A(n2685), .B(n2684), .Z(n2686) );
  NANDN U2850 ( .A(n2602), .B(n2601), .Z(n2606) );
  NANDN U2851 ( .A(n2604), .B(n2603), .Z(n2605) );
  NAND U2852 ( .A(n2606), .B(n2605), .Z(n2687) );
  XNOR U2853 ( .A(n2686), .B(n2687), .Z(n2632) );
  XOR U2854 ( .A(n2633), .B(n2632), .Z(n2691) );
  NANDN U2855 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U2856 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U2857 ( .A(n2612), .B(n2611), .Z(n2690) );
  XNOR U2858 ( .A(n2691), .B(n2690), .Z(n2692) );
  XOR U2859 ( .A(n2693), .B(n2692), .Z(n2625) );
  NANDN U2860 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U2861 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U2862 ( .A(n2618), .B(n2617), .Z(n2624) );
  XNOR U2863 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U2864 ( .A(n2627), .B(n2626), .Z(n2696) );
  XNOR U2865 ( .A(sreg[89]), .B(n2696), .Z(n2698) );
  NANDN U2866 ( .A(sreg[88]), .B(n2619), .Z(n2623) );
  NAND U2867 ( .A(n2621), .B(n2620), .Z(n2622) );
  NAND U2868 ( .A(n2623), .B(n2622), .Z(n2697) );
  XNOR U2869 ( .A(n2698), .B(n2697), .Z(c[89]) );
  NANDN U2870 ( .A(n2625), .B(n2624), .Z(n2629) );
  NANDN U2871 ( .A(n2627), .B(n2626), .Z(n2628) );
  AND U2872 ( .A(n2629), .B(n2628), .Z(n2704) );
  NANDN U2873 ( .A(n2631), .B(n2630), .Z(n2635) );
  NAND U2874 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2875 ( .A(n2635), .B(n2634), .Z(n2770) );
  NAND U2876 ( .A(n4950), .B(n2636), .Z(n2638) );
  XOR U2877 ( .A(b[11]), .B(a[32]), .Z(n2713) );
  NAND U2878 ( .A(n4863), .B(n2713), .Z(n2637) );
  AND U2879 ( .A(n2638), .B(n2637), .Z(n2724) );
  NAND U2880 ( .A(n42), .B(n2639), .Z(n2641) );
  XOR U2881 ( .A(b[15]), .B(a[28]), .Z(n2716) );
  NAND U2882 ( .A(n4981), .B(n2716), .Z(n2640) );
  AND U2883 ( .A(n2641), .B(n2640), .Z(n2723) );
  NAND U2884 ( .A(n41), .B(n2642), .Z(n2644) );
  XOR U2885 ( .A(b[9]), .B(a[34]), .Z(n2719) );
  NAND U2886 ( .A(n4810), .B(n2719), .Z(n2643) );
  NAND U2887 ( .A(n2644), .B(n2643), .Z(n2722) );
  XOR U2888 ( .A(n2723), .B(n2722), .Z(n2725) );
  XOR U2889 ( .A(n2724), .B(n2725), .Z(n2762) );
  NANDN U2890 ( .A(n2646), .B(n2645), .Z(n2650) );
  OR U2891 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U2892 ( .A(n2650), .B(n2649), .Z(n2761) );
  XNOR U2893 ( .A(n2762), .B(n2761), .Z(n2763) );
  NANDN U2894 ( .A(n2652), .B(n2651), .Z(n2656) );
  NANDN U2895 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U2896 ( .A(n2656), .B(n2655), .Z(n2764) );
  XNOR U2897 ( .A(n2763), .B(n2764), .Z(n2710) );
  NANDN U2898 ( .A(n2658), .B(n2657), .Z(n2662) );
  NANDN U2899 ( .A(n2660), .B(n2659), .Z(n2661) );
  AND U2900 ( .A(n2662), .B(n2661), .Z(n2757) );
  NAND U2901 ( .A(b[0]), .B(a[42]), .Z(n2663) );
  XNOR U2902 ( .A(b[1]), .B(n2663), .Z(n2665) );
  NANDN U2903 ( .A(b[0]), .B(a[41]), .Z(n2664) );
  NAND U2904 ( .A(n2665), .B(n2664), .Z(n2737) );
  NAND U2905 ( .A(n5012), .B(n2666), .Z(n2668) );
  XOR U2906 ( .A(b[13]), .B(a[30]), .Z(n2743) );
  NAND U2907 ( .A(n4985), .B(n2743), .Z(n2667) );
  AND U2908 ( .A(n2668), .B(n2667), .Z(n2735) );
  AND U2909 ( .A(b[15]), .B(a[26]), .Z(n2734) );
  XNOR U2910 ( .A(n2735), .B(n2734), .Z(n2736) );
  XNOR U2911 ( .A(n2737), .B(n2736), .Z(n2755) );
  NAND U2912 ( .A(n36), .B(n2669), .Z(n2671) );
  XOR U2913 ( .A(b[5]), .B(a[38]), .Z(n2746) );
  NAND U2914 ( .A(n4560), .B(n2746), .Z(n2670) );
  AND U2915 ( .A(n2671), .B(n2670), .Z(n2731) );
  NAND U2916 ( .A(n4755), .B(n2672), .Z(n2674) );
  XOR U2917 ( .A(b[7]), .B(a[36]), .Z(n2749) );
  NAND U2918 ( .A(n4708), .B(n2749), .Z(n2673) );
  AND U2919 ( .A(n2674), .B(n2673), .Z(n2729) );
  NAND U2920 ( .A(n4471), .B(n2675), .Z(n2677) );
  XOR U2921 ( .A(b[3]), .B(a[40]), .Z(n2752) );
  NAND U2922 ( .A(n33), .B(n2752), .Z(n2676) );
  NAND U2923 ( .A(n2677), .B(n2676), .Z(n2728) );
  XNOR U2924 ( .A(n2729), .B(n2728), .Z(n2730) );
  XOR U2925 ( .A(n2731), .B(n2730), .Z(n2756) );
  XOR U2926 ( .A(n2755), .B(n2756), .Z(n2758) );
  XOR U2927 ( .A(n2757), .B(n2758), .Z(n2708) );
  NANDN U2928 ( .A(n2679), .B(n2678), .Z(n2683) );
  OR U2929 ( .A(n2681), .B(n2680), .Z(n2682) );
  AND U2930 ( .A(n2683), .B(n2682), .Z(n2707) );
  XNOR U2931 ( .A(n2708), .B(n2707), .Z(n2709) );
  XOR U2932 ( .A(n2710), .B(n2709), .Z(n2768) );
  NANDN U2933 ( .A(n2685), .B(n2684), .Z(n2689) );
  NANDN U2934 ( .A(n2687), .B(n2686), .Z(n2688) );
  AND U2935 ( .A(n2689), .B(n2688), .Z(n2767) );
  XNOR U2936 ( .A(n2768), .B(n2767), .Z(n2769) );
  XOR U2937 ( .A(n2770), .B(n2769), .Z(n2702) );
  NANDN U2938 ( .A(n2691), .B(n2690), .Z(n2695) );
  NAND U2939 ( .A(n2693), .B(n2692), .Z(n2694) );
  AND U2940 ( .A(n2695), .B(n2694), .Z(n2701) );
  XNOR U2941 ( .A(n2702), .B(n2701), .Z(n2703) );
  XNOR U2942 ( .A(n2704), .B(n2703), .Z(n2773) );
  XNOR U2943 ( .A(sreg[90]), .B(n2773), .Z(n2775) );
  NANDN U2944 ( .A(sreg[89]), .B(n2696), .Z(n2700) );
  NAND U2945 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U2946 ( .A(n2700), .B(n2699), .Z(n2774) );
  XNOR U2947 ( .A(n2775), .B(n2774), .Z(c[90]) );
  NANDN U2948 ( .A(n2702), .B(n2701), .Z(n2706) );
  NANDN U2949 ( .A(n2704), .B(n2703), .Z(n2705) );
  AND U2950 ( .A(n2706), .B(n2705), .Z(n2781) );
  NANDN U2951 ( .A(n2708), .B(n2707), .Z(n2712) );
  NAND U2952 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U2953 ( .A(n2712), .B(n2711), .Z(n2847) );
  NAND U2954 ( .A(n4950), .B(n2713), .Z(n2715) );
  XOR U2955 ( .A(b[11]), .B(a[33]), .Z(n2817) );
  NAND U2956 ( .A(n4863), .B(n2817), .Z(n2714) );
  AND U2957 ( .A(n2715), .B(n2714), .Z(n2828) );
  NAND U2958 ( .A(n42), .B(n2716), .Z(n2718) );
  XOR U2959 ( .A(b[15]), .B(a[29]), .Z(n2820) );
  NAND U2960 ( .A(n4981), .B(n2820), .Z(n2717) );
  AND U2961 ( .A(n2718), .B(n2717), .Z(n2827) );
  NAND U2962 ( .A(n41), .B(n2719), .Z(n2721) );
  XOR U2963 ( .A(b[9]), .B(a[35]), .Z(n2823) );
  NAND U2964 ( .A(n4810), .B(n2823), .Z(n2720) );
  NAND U2965 ( .A(n2721), .B(n2720), .Z(n2826) );
  XOR U2966 ( .A(n2827), .B(n2826), .Z(n2829) );
  XOR U2967 ( .A(n2828), .B(n2829), .Z(n2839) );
  NANDN U2968 ( .A(n2723), .B(n2722), .Z(n2727) );
  OR U2969 ( .A(n2725), .B(n2724), .Z(n2726) );
  AND U2970 ( .A(n2727), .B(n2726), .Z(n2838) );
  XNOR U2971 ( .A(n2839), .B(n2838), .Z(n2840) );
  NANDN U2972 ( .A(n2729), .B(n2728), .Z(n2733) );
  NANDN U2973 ( .A(n2731), .B(n2730), .Z(n2732) );
  NAND U2974 ( .A(n2733), .B(n2732), .Z(n2841) );
  XNOR U2975 ( .A(n2840), .B(n2841), .Z(n2787) );
  NANDN U2976 ( .A(n2735), .B(n2734), .Z(n2739) );
  NANDN U2977 ( .A(n2737), .B(n2736), .Z(n2738) );
  AND U2978 ( .A(n2739), .B(n2738), .Z(n2813) );
  NAND U2979 ( .A(b[0]), .B(a[43]), .Z(n2740) );
  XNOR U2980 ( .A(b[1]), .B(n2740), .Z(n2742) );
  NANDN U2981 ( .A(b[0]), .B(a[42]), .Z(n2741) );
  NAND U2982 ( .A(n2742), .B(n2741), .Z(n2793) );
  NAND U2983 ( .A(n5012), .B(n2743), .Z(n2745) );
  XOR U2984 ( .A(b[13]), .B(a[31]), .Z(n2799) );
  NAND U2985 ( .A(n4985), .B(n2799), .Z(n2744) );
  AND U2986 ( .A(n2745), .B(n2744), .Z(n2791) );
  AND U2987 ( .A(b[15]), .B(a[27]), .Z(n2790) );
  XNOR U2988 ( .A(n2791), .B(n2790), .Z(n2792) );
  XNOR U2989 ( .A(n2793), .B(n2792), .Z(n2811) );
  NAND U2990 ( .A(n36), .B(n2746), .Z(n2748) );
  XOR U2991 ( .A(b[5]), .B(a[39]), .Z(n2802) );
  NAND U2992 ( .A(n4560), .B(n2802), .Z(n2747) );
  AND U2993 ( .A(n2748), .B(n2747), .Z(n2835) );
  NAND U2994 ( .A(n4755), .B(n2749), .Z(n2751) );
  XOR U2995 ( .A(b[7]), .B(a[37]), .Z(n2805) );
  NAND U2996 ( .A(n4708), .B(n2805), .Z(n2750) );
  AND U2997 ( .A(n2751), .B(n2750), .Z(n2833) );
  NAND U2998 ( .A(n4471), .B(n2752), .Z(n2754) );
  XOR U2999 ( .A(b[3]), .B(a[41]), .Z(n2808) );
  NAND U3000 ( .A(n33), .B(n2808), .Z(n2753) );
  NAND U3001 ( .A(n2754), .B(n2753), .Z(n2832) );
  XNOR U3002 ( .A(n2833), .B(n2832), .Z(n2834) );
  XOR U3003 ( .A(n2835), .B(n2834), .Z(n2812) );
  XOR U3004 ( .A(n2811), .B(n2812), .Z(n2814) );
  XOR U3005 ( .A(n2813), .B(n2814), .Z(n2785) );
  NANDN U3006 ( .A(n2756), .B(n2755), .Z(n2760) );
  OR U3007 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U3008 ( .A(n2760), .B(n2759), .Z(n2784) );
  XNOR U3009 ( .A(n2785), .B(n2784), .Z(n2786) );
  XOR U3010 ( .A(n2787), .B(n2786), .Z(n2845) );
  NANDN U3011 ( .A(n2762), .B(n2761), .Z(n2766) );
  NANDN U3012 ( .A(n2764), .B(n2763), .Z(n2765) );
  AND U3013 ( .A(n2766), .B(n2765), .Z(n2844) );
  XNOR U3014 ( .A(n2845), .B(n2844), .Z(n2846) );
  XOR U3015 ( .A(n2847), .B(n2846), .Z(n2779) );
  NANDN U3016 ( .A(n2768), .B(n2767), .Z(n2772) );
  NAND U3017 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U3018 ( .A(n2772), .B(n2771), .Z(n2778) );
  XNOR U3019 ( .A(n2779), .B(n2778), .Z(n2780) );
  XNOR U3020 ( .A(n2781), .B(n2780), .Z(n2850) );
  XNOR U3021 ( .A(sreg[91]), .B(n2850), .Z(n2852) );
  NANDN U3022 ( .A(sreg[90]), .B(n2773), .Z(n2777) );
  NAND U3023 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3024 ( .A(n2777), .B(n2776), .Z(n2851) );
  XNOR U3025 ( .A(n2852), .B(n2851), .Z(c[91]) );
  NANDN U3026 ( .A(n2779), .B(n2778), .Z(n2783) );
  NANDN U3027 ( .A(n2781), .B(n2780), .Z(n2782) );
  AND U3028 ( .A(n2783), .B(n2782), .Z(n2858) );
  NANDN U3029 ( .A(n2785), .B(n2784), .Z(n2789) );
  NAND U3030 ( .A(n2787), .B(n2786), .Z(n2788) );
  AND U3031 ( .A(n2789), .B(n2788), .Z(n2924) );
  NANDN U3032 ( .A(n2791), .B(n2790), .Z(n2795) );
  NANDN U3033 ( .A(n2793), .B(n2792), .Z(n2794) );
  AND U3034 ( .A(n2795), .B(n2794), .Z(n2911) );
  NAND U3035 ( .A(b[0]), .B(a[44]), .Z(n2796) );
  XNOR U3036 ( .A(b[1]), .B(n2796), .Z(n2798) );
  NANDN U3037 ( .A(b[0]), .B(a[43]), .Z(n2797) );
  NAND U3038 ( .A(n2798), .B(n2797), .Z(n2891) );
  NAND U3039 ( .A(n5012), .B(n2799), .Z(n2801) );
  XOR U3040 ( .A(b[13]), .B(a[32]), .Z(n2897) );
  NAND U3041 ( .A(n4985), .B(n2897), .Z(n2800) );
  AND U3042 ( .A(n2801), .B(n2800), .Z(n2889) );
  AND U3043 ( .A(b[15]), .B(a[28]), .Z(n2888) );
  XNOR U3044 ( .A(n2889), .B(n2888), .Z(n2890) );
  XNOR U3045 ( .A(n2891), .B(n2890), .Z(n2909) );
  NAND U3046 ( .A(n36), .B(n2802), .Z(n2804) );
  XOR U3047 ( .A(b[5]), .B(a[40]), .Z(n2900) );
  NAND U3048 ( .A(n4560), .B(n2900), .Z(n2803) );
  AND U3049 ( .A(n2804), .B(n2803), .Z(n2885) );
  NAND U3050 ( .A(n4755), .B(n2805), .Z(n2807) );
  XOR U3051 ( .A(b[7]), .B(a[38]), .Z(n2903) );
  NAND U3052 ( .A(n4708), .B(n2903), .Z(n2806) );
  AND U3053 ( .A(n2807), .B(n2806), .Z(n2883) );
  NAND U3054 ( .A(n4471), .B(n2808), .Z(n2810) );
  XOR U3055 ( .A(b[3]), .B(a[42]), .Z(n2906) );
  NAND U3056 ( .A(n33), .B(n2906), .Z(n2809) );
  NAND U3057 ( .A(n2810), .B(n2809), .Z(n2882) );
  XNOR U3058 ( .A(n2883), .B(n2882), .Z(n2884) );
  XOR U3059 ( .A(n2885), .B(n2884), .Z(n2910) );
  XOR U3060 ( .A(n2909), .B(n2910), .Z(n2912) );
  XOR U3061 ( .A(n2911), .B(n2912), .Z(n2862) );
  NANDN U3062 ( .A(n2812), .B(n2811), .Z(n2816) );
  OR U3063 ( .A(n2814), .B(n2813), .Z(n2815) );
  AND U3064 ( .A(n2816), .B(n2815), .Z(n2861) );
  XNOR U3065 ( .A(n2862), .B(n2861), .Z(n2864) );
  NAND U3066 ( .A(n4950), .B(n2817), .Z(n2819) );
  XOR U3067 ( .A(b[11]), .B(a[34]), .Z(n2867) );
  NAND U3068 ( .A(n4863), .B(n2867), .Z(n2818) );
  AND U3069 ( .A(n2819), .B(n2818), .Z(n2878) );
  NAND U3070 ( .A(n42), .B(n2820), .Z(n2822) );
  XOR U3071 ( .A(b[15]), .B(a[30]), .Z(n2870) );
  NAND U3072 ( .A(n4981), .B(n2870), .Z(n2821) );
  AND U3073 ( .A(n2822), .B(n2821), .Z(n2877) );
  NAND U3074 ( .A(n41), .B(n2823), .Z(n2825) );
  XOR U3075 ( .A(b[9]), .B(a[36]), .Z(n2873) );
  NAND U3076 ( .A(n4810), .B(n2873), .Z(n2824) );
  NAND U3077 ( .A(n2825), .B(n2824), .Z(n2876) );
  XOR U3078 ( .A(n2877), .B(n2876), .Z(n2879) );
  XOR U3079 ( .A(n2878), .B(n2879), .Z(n2916) );
  NANDN U3080 ( .A(n2827), .B(n2826), .Z(n2831) );
  OR U3081 ( .A(n2829), .B(n2828), .Z(n2830) );
  AND U3082 ( .A(n2831), .B(n2830), .Z(n2915) );
  XNOR U3083 ( .A(n2916), .B(n2915), .Z(n2917) );
  NANDN U3084 ( .A(n2833), .B(n2832), .Z(n2837) );
  NANDN U3085 ( .A(n2835), .B(n2834), .Z(n2836) );
  NAND U3086 ( .A(n2837), .B(n2836), .Z(n2918) );
  XNOR U3087 ( .A(n2917), .B(n2918), .Z(n2863) );
  XOR U3088 ( .A(n2864), .B(n2863), .Z(n2922) );
  NANDN U3089 ( .A(n2839), .B(n2838), .Z(n2843) );
  NANDN U3090 ( .A(n2841), .B(n2840), .Z(n2842) );
  AND U3091 ( .A(n2843), .B(n2842), .Z(n2921) );
  XNOR U3092 ( .A(n2922), .B(n2921), .Z(n2923) );
  XOR U3093 ( .A(n2924), .B(n2923), .Z(n2856) );
  NANDN U3094 ( .A(n2845), .B(n2844), .Z(n2849) );
  NAND U3095 ( .A(n2847), .B(n2846), .Z(n2848) );
  AND U3096 ( .A(n2849), .B(n2848), .Z(n2855) );
  XNOR U3097 ( .A(n2856), .B(n2855), .Z(n2857) );
  XNOR U3098 ( .A(n2858), .B(n2857), .Z(n2927) );
  XNOR U3099 ( .A(sreg[92]), .B(n2927), .Z(n2929) );
  NANDN U3100 ( .A(sreg[91]), .B(n2850), .Z(n2854) );
  NAND U3101 ( .A(n2852), .B(n2851), .Z(n2853) );
  NAND U3102 ( .A(n2854), .B(n2853), .Z(n2928) );
  XNOR U3103 ( .A(n2929), .B(n2928), .Z(c[92]) );
  NANDN U3104 ( .A(n2856), .B(n2855), .Z(n2860) );
  NANDN U3105 ( .A(n2858), .B(n2857), .Z(n2859) );
  AND U3106 ( .A(n2860), .B(n2859), .Z(n2935) );
  NANDN U3107 ( .A(n2862), .B(n2861), .Z(n2866) );
  NAND U3108 ( .A(n2864), .B(n2863), .Z(n2865) );
  AND U3109 ( .A(n2866), .B(n2865), .Z(n3001) );
  NAND U3110 ( .A(n4950), .B(n2867), .Z(n2869) );
  XOR U3111 ( .A(b[11]), .B(a[35]), .Z(n2971) );
  NAND U3112 ( .A(n4863), .B(n2971), .Z(n2868) );
  AND U3113 ( .A(n2869), .B(n2868), .Z(n2982) );
  NAND U3114 ( .A(n42), .B(n2870), .Z(n2872) );
  XOR U3115 ( .A(b[15]), .B(a[31]), .Z(n2974) );
  NAND U3116 ( .A(n4981), .B(n2974), .Z(n2871) );
  AND U3117 ( .A(n2872), .B(n2871), .Z(n2981) );
  NAND U3118 ( .A(n41), .B(n2873), .Z(n2875) );
  XOR U3119 ( .A(b[9]), .B(a[37]), .Z(n2977) );
  NAND U3120 ( .A(n4810), .B(n2977), .Z(n2874) );
  NAND U3121 ( .A(n2875), .B(n2874), .Z(n2980) );
  XOR U3122 ( .A(n2981), .B(n2980), .Z(n2983) );
  XOR U3123 ( .A(n2982), .B(n2983), .Z(n2993) );
  NANDN U3124 ( .A(n2877), .B(n2876), .Z(n2881) );
  OR U3125 ( .A(n2879), .B(n2878), .Z(n2880) );
  AND U3126 ( .A(n2881), .B(n2880), .Z(n2992) );
  XNOR U3127 ( .A(n2993), .B(n2992), .Z(n2994) );
  NANDN U3128 ( .A(n2883), .B(n2882), .Z(n2887) );
  NANDN U3129 ( .A(n2885), .B(n2884), .Z(n2886) );
  NAND U3130 ( .A(n2887), .B(n2886), .Z(n2995) );
  XNOR U3131 ( .A(n2994), .B(n2995), .Z(n2941) );
  NANDN U3132 ( .A(n2889), .B(n2888), .Z(n2893) );
  NANDN U3133 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3134 ( .A(n2893), .B(n2892), .Z(n2967) );
  NAND U3135 ( .A(b[0]), .B(a[45]), .Z(n2894) );
  XNOR U3136 ( .A(b[1]), .B(n2894), .Z(n2896) );
  NANDN U3137 ( .A(b[0]), .B(a[44]), .Z(n2895) );
  NAND U3138 ( .A(n2896), .B(n2895), .Z(n2947) );
  NAND U3139 ( .A(n5012), .B(n2897), .Z(n2899) );
  XOR U3140 ( .A(b[13]), .B(a[33]), .Z(n2953) );
  NAND U3141 ( .A(n4985), .B(n2953), .Z(n2898) );
  AND U3142 ( .A(n2899), .B(n2898), .Z(n2945) );
  AND U3143 ( .A(b[15]), .B(a[29]), .Z(n2944) );
  XNOR U3144 ( .A(n2945), .B(n2944), .Z(n2946) );
  XNOR U3145 ( .A(n2947), .B(n2946), .Z(n2965) );
  NAND U3146 ( .A(n36), .B(n2900), .Z(n2902) );
  XOR U3147 ( .A(b[5]), .B(a[41]), .Z(n2956) );
  NAND U3148 ( .A(n4560), .B(n2956), .Z(n2901) );
  AND U3149 ( .A(n2902), .B(n2901), .Z(n2989) );
  NAND U3150 ( .A(n4755), .B(n2903), .Z(n2905) );
  XOR U3151 ( .A(b[7]), .B(a[39]), .Z(n2959) );
  NAND U3152 ( .A(n4708), .B(n2959), .Z(n2904) );
  AND U3153 ( .A(n2905), .B(n2904), .Z(n2987) );
  NAND U3154 ( .A(n4471), .B(n2906), .Z(n2908) );
  XOR U3155 ( .A(b[3]), .B(a[43]), .Z(n2962) );
  NAND U3156 ( .A(n33), .B(n2962), .Z(n2907) );
  NAND U3157 ( .A(n2908), .B(n2907), .Z(n2986) );
  XNOR U3158 ( .A(n2987), .B(n2986), .Z(n2988) );
  XOR U3159 ( .A(n2989), .B(n2988), .Z(n2966) );
  XOR U3160 ( .A(n2965), .B(n2966), .Z(n2968) );
  XOR U3161 ( .A(n2967), .B(n2968), .Z(n2939) );
  NANDN U3162 ( .A(n2910), .B(n2909), .Z(n2914) );
  OR U3163 ( .A(n2912), .B(n2911), .Z(n2913) );
  AND U3164 ( .A(n2914), .B(n2913), .Z(n2938) );
  XNOR U3165 ( .A(n2939), .B(n2938), .Z(n2940) );
  XOR U3166 ( .A(n2941), .B(n2940), .Z(n2999) );
  NANDN U3167 ( .A(n2916), .B(n2915), .Z(n2920) );
  NANDN U3168 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3169 ( .A(n2920), .B(n2919), .Z(n2998) );
  XNOR U3170 ( .A(n2999), .B(n2998), .Z(n3000) );
  XOR U3171 ( .A(n3001), .B(n3000), .Z(n2933) );
  NANDN U3172 ( .A(n2922), .B(n2921), .Z(n2926) );
  NAND U3173 ( .A(n2924), .B(n2923), .Z(n2925) );
  AND U3174 ( .A(n2926), .B(n2925), .Z(n2932) );
  XNOR U3175 ( .A(n2933), .B(n2932), .Z(n2934) );
  XNOR U3176 ( .A(n2935), .B(n2934), .Z(n3004) );
  XNOR U3177 ( .A(sreg[93]), .B(n3004), .Z(n3006) );
  NANDN U3178 ( .A(sreg[92]), .B(n2927), .Z(n2931) );
  NAND U3179 ( .A(n2929), .B(n2928), .Z(n2930) );
  NAND U3180 ( .A(n2931), .B(n2930), .Z(n3005) );
  XNOR U3181 ( .A(n3006), .B(n3005), .Z(c[93]) );
  NANDN U3182 ( .A(n2933), .B(n2932), .Z(n2937) );
  NANDN U3183 ( .A(n2935), .B(n2934), .Z(n2936) );
  AND U3184 ( .A(n2937), .B(n2936), .Z(n3012) );
  NANDN U3185 ( .A(n2939), .B(n2938), .Z(n2943) );
  NAND U3186 ( .A(n2941), .B(n2940), .Z(n2942) );
  AND U3187 ( .A(n2943), .B(n2942), .Z(n3078) );
  NANDN U3188 ( .A(n2945), .B(n2944), .Z(n2949) );
  NANDN U3189 ( .A(n2947), .B(n2946), .Z(n2948) );
  AND U3190 ( .A(n2949), .B(n2948), .Z(n3044) );
  NAND U3191 ( .A(b[0]), .B(a[46]), .Z(n2950) );
  XNOR U3192 ( .A(b[1]), .B(n2950), .Z(n2952) );
  NANDN U3193 ( .A(b[0]), .B(a[45]), .Z(n2951) );
  NAND U3194 ( .A(n2952), .B(n2951), .Z(n3024) );
  NAND U3195 ( .A(n5012), .B(n2953), .Z(n2955) );
  XOR U3196 ( .A(b[13]), .B(a[34]), .Z(n3030) );
  NAND U3197 ( .A(n4985), .B(n3030), .Z(n2954) );
  AND U3198 ( .A(n2955), .B(n2954), .Z(n3022) );
  AND U3199 ( .A(b[15]), .B(a[30]), .Z(n3021) );
  XNOR U3200 ( .A(n3022), .B(n3021), .Z(n3023) );
  XNOR U3201 ( .A(n3024), .B(n3023), .Z(n3042) );
  NAND U3202 ( .A(n36), .B(n2956), .Z(n2958) );
  XOR U3203 ( .A(b[5]), .B(a[42]), .Z(n3033) );
  NAND U3204 ( .A(n4560), .B(n3033), .Z(n2957) );
  AND U3205 ( .A(n2958), .B(n2957), .Z(n3066) );
  NAND U3206 ( .A(n4755), .B(n2959), .Z(n2961) );
  XOR U3207 ( .A(b[7]), .B(a[40]), .Z(n3036) );
  NAND U3208 ( .A(n4708), .B(n3036), .Z(n2960) );
  AND U3209 ( .A(n2961), .B(n2960), .Z(n3064) );
  NAND U3210 ( .A(n4471), .B(n2962), .Z(n2964) );
  XOR U3211 ( .A(b[3]), .B(a[44]), .Z(n3039) );
  NAND U3212 ( .A(n33), .B(n3039), .Z(n2963) );
  NAND U3213 ( .A(n2964), .B(n2963), .Z(n3063) );
  XNOR U3214 ( .A(n3064), .B(n3063), .Z(n3065) );
  XOR U3215 ( .A(n3066), .B(n3065), .Z(n3043) );
  XOR U3216 ( .A(n3042), .B(n3043), .Z(n3045) );
  XOR U3217 ( .A(n3044), .B(n3045), .Z(n3016) );
  NANDN U3218 ( .A(n2966), .B(n2965), .Z(n2970) );
  OR U3219 ( .A(n2968), .B(n2967), .Z(n2969) );
  AND U3220 ( .A(n2970), .B(n2969), .Z(n3015) );
  XNOR U3221 ( .A(n3016), .B(n3015), .Z(n3018) );
  NAND U3222 ( .A(n4950), .B(n2971), .Z(n2973) );
  XOR U3223 ( .A(b[11]), .B(a[36]), .Z(n3048) );
  NAND U3224 ( .A(n4863), .B(n3048), .Z(n2972) );
  AND U3225 ( .A(n2973), .B(n2972), .Z(n3059) );
  NAND U3226 ( .A(n42), .B(n2974), .Z(n2976) );
  XOR U3227 ( .A(b[15]), .B(a[32]), .Z(n3051) );
  NAND U3228 ( .A(n4981), .B(n3051), .Z(n2975) );
  AND U3229 ( .A(n2976), .B(n2975), .Z(n3058) );
  NAND U3230 ( .A(n41), .B(n2977), .Z(n2979) );
  XOR U3231 ( .A(b[9]), .B(a[38]), .Z(n3054) );
  NAND U3232 ( .A(n4810), .B(n3054), .Z(n2978) );
  NAND U3233 ( .A(n2979), .B(n2978), .Z(n3057) );
  XOR U3234 ( .A(n3058), .B(n3057), .Z(n3060) );
  XOR U3235 ( .A(n3059), .B(n3060), .Z(n3070) );
  NANDN U3236 ( .A(n2981), .B(n2980), .Z(n2985) );
  OR U3237 ( .A(n2983), .B(n2982), .Z(n2984) );
  AND U3238 ( .A(n2985), .B(n2984), .Z(n3069) );
  XNOR U3239 ( .A(n3070), .B(n3069), .Z(n3071) );
  NANDN U3240 ( .A(n2987), .B(n2986), .Z(n2991) );
  NANDN U3241 ( .A(n2989), .B(n2988), .Z(n2990) );
  NAND U3242 ( .A(n2991), .B(n2990), .Z(n3072) );
  XNOR U3243 ( .A(n3071), .B(n3072), .Z(n3017) );
  XOR U3244 ( .A(n3018), .B(n3017), .Z(n3076) );
  NANDN U3245 ( .A(n2993), .B(n2992), .Z(n2997) );
  NANDN U3246 ( .A(n2995), .B(n2994), .Z(n2996) );
  AND U3247 ( .A(n2997), .B(n2996), .Z(n3075) );
  XNOR U3248 ( .A(n3076), .B(n3075), .Z(n3077) );
  XOR U3249 ( .A(n3078), .B(n3077), .Z(n3010) );
  NANDN U3250 ( .A(n2999), .B(n2998), .Z(n3003) );
  NAND U3251 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3252 ( .A(n3003), .B(n3002), .Z(n3009) );
  XNOR U3253 ( .A(n3010), .B(n3009), .Z(n3011) );
  XNOR U3254 ( .A(n3012), .B(n3011), .Z(n3081) );
  XNOR U3255 ( .A(sreg[94]), .B(n3081), .Z(n3083) );
  NANDN U3256 ( .A(sreg[93]), .B(n3004), .Z(n3008) );
  NAND U3257 ( .A(n3006), .B(n3005), .Z(n3007) );
  NAND U3258 ( .A(n3008), .B(n3007), .Z(n3082) );
  XNOR U3259 ( .A(n3083), .B(n3082), .Z(c[94]) );
  NANDN U3260 ( .A(n3010), .B(n3009), .Z(n3014) );
  NANDN U3261 ( .A(n3012), .B(n3011), .Z(n3013) );
  AND U3262 ( .A(n3014), .B(n3013), .Z(n3089) );
  NANDN U3263 ( .A(n3016), .B(n3015), .Z(n3020) );
  NAND U3264 ( .A(n3018), .B(n3017), .Z(n3019) );
  AND U3265 ( .A(n3020), .B(n3019), .Z(n3155) );
  NANDN U3266 ( .A(n3022), .B(n3021), .Z(n3026) );
  NANDN U3267 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U3268 ( .A(n3026), .B(n3025), .Z(n3121) );
  NAND U3269 ( .A(b[0]), .B(a[47]), .Z(n3027) );
  XNOR U3270 ( .A(b[1]), .B(n3027), .Z(n3029) );
  NANDN U3271 ( .A(b[0]), .B(a[46]), .Z(n3028) );
  NAND U3272 ( .A(n3029), .B(n3028), .Z(n3101) );
  NAND U3273 ( .A(n5012), .B(n3030), .Z(n3032) );
  XOR U3274 ( .A(b[13]), .B(a[35]), .Z(n3104) );
  NAND U3275 ( .A(n4985), .B(n3104), .Z(n3031) );
  AND U3276 ( .A(n3032), .B(n3031), .Z(n3099) );
  AND U3277 ( .A(b[15]), .B(a[31]), .Z(n3098) );
  XNOR U3278 ( .A(n3099), .B(n3098), .Z(n3100) );
  XNOR U3279 ( .A(n3101), .B(n3100), .Z(n3119) );
  NAND U3280 ( .A(n36), .B(n3033), .Z(n3035) );
  XOR U3281 ( .A(b[5]), .B(a[43]), .Z(n3110) );
  NAND U3282 ( .A(n4560), .B(n3110), .Z(n3034) );
  AND U3283 ( .A(n3035), .B(n3034), .Z(n3143) );
  NAND U3284 ( .A(n4755), .B(n3036), .Z(n3038) );
  XOR U3285 ( .A(b[7]), .B(a[41]), .Z(n3113) );
  NAND U3286 ( .A(n4708), .B(n3113), .Z(n3037) );
  AND U3287 ( .A(n3038), .B(n3037), .Z(n3141) );
  NAND U3288 ( .A(n4471), .B(n3039), .Z(n3041) );
  XOR U3289 ( .A(b[3]), .B(a[45]), .Z(n3116) );
  NAND U3290 ( .A(n33), .B(n3116), .Z(n3040) );
  NAND U3291 ( .A(n3041), .B(n3040), .Z(n3140) );
  XNOR U3292 ( .A(n3141), .B(n3140), .Z(n3142) );
  XOR U3293 ( .A(n3143), .B(n3142), .Z(n3120) );
  XOR U3294 ( .A(n3119), .B(n3120), .Z(n3122) );
  XOR U3295 ( .A(n3121), .B(n3122), .Z(n3093) );
  NANDN U3296 ( .A(n3043), .B(n3042), .Z(n3047) );
  OR U3297 ( .A(n3045), .B(n3044), .Z(n3046) );
  AND U3298 ( .A(n3047), .B(n3046), .Z(n3092) );
  XNOR U3299 ( .A(n3093), .B(n3092), .Z(n3095) );
  NAND U3300 ( .A(n4950), .B(n3048), .Z(n3050) );
  XOR U3301 ( .A(b[11]), .B(a[37]), .Z(n3125) );
  NAND U3302 ( .A(n4863), .B(n3125), .Z(n3049) );
  AND U3303 ( .A(n3050), .B(n3049), .Z(n3136) );
  NAND U3304 ( .A(n42), .B(n3051), .Z(n3053) );
  XOR U3305 ( .A(b[15]), .B(a[33]), .Z(n3128) );
  NAND U3306 ( .A(n4981), .B(n3128), .Z(n3052) );
  AND U3307 ( .A(n3053), .B(n3052), .Z(n3135) );
  NAND U3308 ( .A(n41), .B(n3054), .Z(n3056) );
  XOR U3309 ( .A(b[9]), .B(a[39]), .Z(n3131) );
  NAND U3310 ( .A(n4810), .B(n3131), .Z(n3055) );
  NAND U3311 ( .A(n3056), .B(n3055), .Z(n3134) );
  XOR U3312 ( .A(n3135), .B(n3134), .Z(n3137) );
  XOR U3313 ( .A(n3136), .B(n3137), .Z(n3147) );
  NANDN U3314 ( .A(n3058), .B(n3057), .Z(n3062) );
  OR U3315 ( .A(n3060), .B(n3059), .Z(n3061) );
  AND U3316 ( .A(n3062), .B(n3061), .Z(n3146) );
  XNOR U3317 ( .A(n3147), .B(n3146), .Z(n3148) );
  NANDN U3318 ( .A(n3064), .B(n3063), .Z(n3068) );
  NANDN U3319 ( .A(n3066), .B(n3065), .Z(n3067) );
  NAND U3320 ( .A(n3068), .B(n3067), .Z(n3149) );
  XNOR U3321 ( .A(n3148), .B(n3149), .Z(n3094) );
  XOR U3322 ( .A(n3095), .B(n3094), .Z(n3153) );
  NANDN U3323 ( .A(n3070), .B(n3069), .Z(n3074) );
  NANDN U3324 ( .A(n3072), .B(n3071), .Z(n3073) );
  AND U3325 ( .A(n3074), .B(n3073), .Z(n3152) );
  XNOR U3326 ( .A(n3153), .B(n3152), .Z(n3154) );
  XOR U3327 ( .A(n3155), .B(n3154), .Z(n3087) );
  NANDN U3328 ( .A(n3076), .B(n3075), .Z(n3080) );
  NAND U3329 ( .A(n3078), .B(n3077), .Z(n3079) );
  AND U3330 ( .A(n3080), .B(n3079), .Z(n3086) );
  XNOR U3331 ( .A(n3087), .B(n3086), .Z(n3088) );
  XNOR U3332 ( .A(n3089), .B(n3088), .Z(n3158) );
  XNOR U3333 ( .A(sreg[95]), .B(n3158), .Z(n3160) );
  NANDN U3334 ( .A(sreg[94]), .B(n3081), .Z(n3085) );
  NAND U3335 ( .A(n3083), .B(n3082), .Z(n3084) );
  NAND U3336 ( .A(n3085), .B(n3084), .Z(n3159) );
  XNOR U3337 ( .A(n3160), .B(n3159), .Z(c[95]) );
  NANDN U3338 ( .A(n3087), .B(n3086), .Z(n3091) );
  NANDN U3339 ( .A(n3089), .B(n3088), .Z(n3090) );
  AND U3340 ( .A(n3091), .B(n3090), .Z(n3166) );
  NANDN U3341 ( .A(n3093), .B(n3092), .Z(n3097) );
  NAND U3342 ( .A(n3095), .B(n3094), .Z(n3096) );
  AND U3343 ( .A(n3097), .B(n3096), .Z(n3232) );
  NANDN U3344 ( .A(n3099), .B(n3098), .Z(n3103) );
  NANDN U3345 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3346 ( .A(n3103), .B(n3102), .Z(n3198) );
  NAND U3347 ( .A(n5012), .B(n3104), .Z(n3106) );
  XOR U3348 ( .A(b[13]), .B(a[36]), .Z(n3184) );
  NAND U3349 ( .A(n4985), .B(n3184), .Z(n3105) );
  AND U3350 ( .A(n3106), .B(n3105), .Z(n3176) );
  AND U3351 ( .A(b[15]), .B(a[32]), .Z(n3175) );
  XNOR U3352 ( .A(n3176), .B(n3175), .Z(n3177) );
  NAND U3353 ( .A(b[0]), .B(a[48]), .Z(n3107) );
  XNOR U3354 ( .A(b[1]), .B(n3107), .Z(n3109) );
  NANDN U3355 ( .A(b[0]), .B(a[47]), .Z(n3108) );
  NAND U3356 ( .A(n3109), .B(n3108), .Z(n3178) );
  XNOR U3357 ( .A(n3177), .B(n3178), .Z(n3196) );
  NAND U3358 ( .A(n36), .B(n3110), .Z(n3112) );
  XOR U3359 ( .A(b[5]), .B(a[44]), .Z(n3187) );
  NAND U3360 ( .A(n4560), .B(n3187), .Z(n3111) );
  AND U3361 ( .A(n3112), .B(n3111), .Z(n3220) );
  NAND U3362 ( .A(n4755), .B(n3113), .Z(n3115) );
  XOR U3363 ( .A(b[7]), .B(a[42]), .Z(n3190) );
  NAND U3364 ( .A(n4708), .B(n3190), .Z(n3114) );
  AND U3365 ( .A(n3115), .B(n3114), .Z(n3218) );
  NAND U3366 ( .A(n4471), .B(n3116), .Z(n3118) );
  XOR U3367 ( .A(b[3]), .B(a[46]), .Z(n3193) );
  NAND U3368 ( .A(n33), .B(n3193), .Z(n3117) );
  NAND U3369 ( .A(n3118), .B(n3117), .Z(n3217) );
  XNOR U3370 ( .A(n3218), .B(n3217), .Z(n3219) );
  XOR U3371 ( .A(n3220), .B(n3219), .Z(n3197) );
  XOR U3372 ( .A(n3196), .B(n3197), .Z(n3199) );
  XOR U3373 ( .A(n3198), .B(n3199), .Z(n3170) );
  NANDN U3374 ( .A(n3120), .B(n3119), .Z(n3124) );
  OR U3375 ( .A(n3122), .B(n3121), .Z(n3123) );
  AND U3376 ( .A(n3124), .B(n3123), .Z(n3169) );
  XNOR U3377 ( .A(n3170), .B(n3169), .Z(n3172) );
  NAND U3378 ( .A(n4950), .B(n3125), .Z(n3127) );
  XOR U3379 ( .A(b[11]), .B(a[38]), .Z(n3202) );
  NAND U3380 ( .A(n4863), .B(n3202), .Z(n3126) );
  AND U3381 ( .A(n3127), .B(n3126), .Z(n3213) );
  NAND U3382 ( .A(n42), .B(n3128), .Z(n3130) );
  XOR U3383 ( .A(b[15]), .B(a[34]), .Z(n3205) );
  NAND U3384 ( .A(n4981), .B(n3205), .Z(n3129) );
  AND U3385 ( .A(n3130), .B(n3129), .Z(n3212) );
  NAND U3386 ( .A(n41), .B(n3131), .Z(n3133) );
  XOR U3387 ( .A(b[9]), .B(a[40]), .Z(n3208) );
  NAND U3388 ( .A(n4810), .B(n3208), .Z(n3132) );
  NAND U3389 ( .A(n3133), .B(n3132), .Z(n3211) );
  XOR U3390 ( .A(n3212), .B(n3211), .Z(n3214) );
  XOR U3391 ( .A(n3213), .B(n3214), .Z(n3224) );
  NANDN U3392 ( .A(n3135), .B(n3134), .Z(n3139) );
  OR U3393 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3394 ( .A(n3139), .B(n3138), .Z(n3223) );
  XNOR U3395 ( .A(n3224), .B(n3223), .Z(n3225) );
  NANDN U3396 ( .A(n3141), .B(n3140), .Z(n3145) );
  NANDN U3397 ( .A(n3143), .B(n3142), .Z(n3144) );
  NAND U3398 ( .A(n3145), .B(n3144), .Z(n3226) );
  XNOR U3399 ( .A(n3225), .B(n3226), .Z(n3171) );
  XOR U3400 ( .A(n3172), .B(n3171), .Z(n3230) );
  NANDN U3401 ( .A(n3147), .B(n3146), .Z(n3151) );
  NANDN U3402 ( .A(n3149), .B(n3148), .Z(n3150) );
  AND U3403 ( .A(n3151), .B(n3150), .Z(n3229) );
  XNOR U3404 ( .A(n3230), .B(n3229), .Z(n3231) );
  XOR U3405 ( .A(n3232), .B(n3231), .Z(n3164) );
  NANDN U3406 ( .A(n3153), .B(n3152), .Z(n3157) );
  NAND U3407 ( .A(n3155), .B(n3154), .Z(n3156) );
  AND U3408 ( .A(n3157), .B(n3156), .Z(n3163) );
  XNOR U3409 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U3410 ( .A(n3166), .B(n3165), .Z(n3235) );
  XNOR U3411 ( .A(sreg[96]), .B(n3235), .Z(n3237) );
  NANDN U3412 ( .A(sreg[95]), .B(n3158), .Z(n3162) );
  NAND U3413 ( .A(n3160), .B(n3159), .Z(n3161) );
  NAND U3414 ( .A(n3162), .B(n3161), .Z(n3236) );
  XNOR U3415 ( .A(n3237), .B(n3236), .Z(c[96]) );
  NANDN U3416 ( .A(n3164), .B(n3163), .Z(n3168) );
  NANDN U3417 ( .A(n3166), .B(n3165), .Z(n3167) );
  AND U3418 ( .A(n3168), .B(n3167), .Z(n3243) );
  NANDN U3419 ( .A(n3170), .B(n3169), .Z(n3174) );
  NAND U3420 ( .A(n3172), .B(n3171), .Z(n3173) );
  AND U3421 ( .A(n3174), .B(n3173), .Z(n3309) );
  NANDN U3422 ( .A(n3176), .B(n3175), .Z(n3180) );
  NANDN U3423 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3424 ( .A(n3180), .B(n3179), .Z(n3275) );
  NAND U3425 ( .A(b[0]), .B(a[49]), .Z(n3181) );
  XNOR U3426 ( .A(b[1]), .B(n3181), .Z(n3183) );
  NANDN U3427 ( .A(b[0]), .B(a[48]), .Z(n3182) );
  NAND U3428 ( .A(n3183), .B(n3182), .Z(n3255) );
  NAND U3429 ( .A(n5012), .B(n3184), .Z(n3186) );
  XOR U3430 ( .A(b[13]), .B(a[37]), .Z(n3261) );
  NAND U3431 ( .A(n4985), .B(n3261), .Z(n3185) );
  AND U3432 ( .A(n3186), .B(n3185), .Z(n3253) );
  AND U3433 ( .A(b[15]), .B(a[33]), .Z(n3252) );
  XNOR U3434 ( .A(n3253), .B(n3252), .Z(n3254) );
  XNOR U3435 ( .A(n3255), .B(n3254), .Z(n3273) );
  NAND U3436 ( .A(n36), .B(n3187), .Z(n3189) );
  XOR U3437 ( .A(b[5]), .B(a[45]), .Z(n3264) );
  NAND U3438 ( .A(n4560), .B(n3264), .Z(n3188) );
  AND U3439 ( .A(n3189), .B(n3188), .Z(n3297) );
  NAND U3440 ( .A(n4755), .B(n3190), .Z(n3192) );
  XOR U3441 ( .A(b[7]), .B(a[43]), .Z(n3267) );
  NAND U3442 ( .A(n4708), .B(n3267), .Z(n3191) );
  AND U3443 ( .A(n3192), .B(n3191), .Z(n3295) );
  NAND U3444 ( .A(n4471), .B(n3193), .Z(n3195) );
  XOR U3445 ( .A(b[3]), .B(a[47]), .Z(n3270) );
  NAND U3446 ( .A(n33), .B(n3270), .Z(n3194) );
  NAND U3447 ( .A(n3195), .B(n3194), .Z(n3294) );
  XNOR U3448 ( .A(n3295), .B(n3294), .Z(n3296) );
  XOR U3449 ( .A(n3297), .B(n3296), .Z(n3274) );
  XOR U3450 ( .A(n3273), .B(n3274), .Z(n3276) );
  XOR U3451 ( .A(n3275), .B(n3276), .Z(n3247) );
  NANDN U3452 ( .A(n3197), .B(n3196), .Z(n3201) );
  OR U3453 ( .A(n3199), .B(n3198), .Z(n3200) );
  AND U3454 ( .A(n3201), .B(n3200), .Z(n3246) );
  XNOR U3455 ( .A(n3247), .B(n3246), .Z(n3249) );
  NAND U3456 ( .A(n4950), .B(n3202), .Z(n3204) );
  XOR U3457 ( .A(b[11]), .B(a[39]), .Z(n3279) );
  NAND U3458 ( .A(n4863), .B(n3279), .Z(n3203) );
  AND U3459 ( .A(n3204), .B(n3203), .Z(n3290) );
  NAND U3460 ( .A(n42), .B(n3205), .Z(n3207) );
  XOR U3461 ( .A(b[15]), .B(a[35]), .Z(n3282) );
  NAND U3462 ( .A(n4981), .B(n3282), .Z(n3206) );
  AND U3463 ( .A(n3207), .B(n3206), .Z(n3289) );
  NAND U3464 ( .A(n41), .B(n3208), .Z(n3210) );
  XOR U3465 ( .A(b[9]), .B(a[41]), .Z(n3285) );
  NAND U3466 ( .A(n4810), .B(n3285), .Z(n3209) );
  NAND U3467 ( .A(n3210), .B(n3209), .Z(n3288) );
  XOR U3468 ( .A(n3289), .B(n3288), .Z(n3291) );
  XOR U3469 ( .A(n3290), .B(n3291), .Z(n3301) );
  NANDN U3470 ( .A(n3212), .B(n3211), .Z(n3216) );
  OR U3471 ( .A(n3214), .B(n3213), .Z(n3215) );
  AND U3472 ( .A(n3216), .B(n3215), .Z(n3300) );
  XNOR U3473 ( .A(n3301), .B(n3300), .Z(n3302) );
  NANDN U3474 ( .A(n3218), .B(n3217), .Z(n3222) );
  NANDN U3475 ( .A(n3220), .B(n3219), .Z(n3221) );
  NAND U3476 ( .A(n3222), .B(n3221), .Z(n3303) );
  XNOR U3477 ( .A(n3302), .B(n3303), .Z(n3248) );
  XOR U3478 ( .A(n3249), .B(n3248), .Z(n3307) );
  NANDN U3479 ( .A(n3224), .B(n3223), .Z(n3228) );
  NANDN U3480 ( .A(n3226), .B(n3225), .Z(n3227) );
  AND U3481 ( .A(n3228), .B(n3227), .Z(n3306) );
  XNOR U3482 ( .A(n3307), .B(n3306), .Z(n3308) );
  XOR U3483 ( .A(n3309), .B(n3308), .Z(n3241) );
  NANDN U3484 ( .A(n3230), .B(n3229), .Z(n3234) );
  NAND U3485 ( .A(n3232), .B(n3231), .Z(n3233) );
  AND U3486 ( .A(n3234), .B(n3233), .Z(n3240) );
  XNOR U3487 ( .A(n3241), .B(n3240), .Z(n3242) );
  XNOR U3488 ( .A(n3243), .B(n3242), .Z(n3312) );
  XNOR U3489 ( .A(sreg[97]), .B(n3312), .Z(n3314) );
  NANDN U3490 ( .A(sreg[96]), .B(n3235), .Z(n3239) );
  NAND U3491 ( .A(n3237), .B(n3236), .Z(n3238) );
  NAND U3492 ( .A(n3239), .B(n3238), .Z(n3313) );
  XNOR U3493 ( .A(n3314), .B(n3313), .Z(c[97]) );
  NANDN U3494 ( .A(n3241), .B(n3240), .Z(n3245) );
  NANDN U3495 ( .A(n3243), .B(n3242), .Z(n3244) );
  AND U3496 ( .A(n3245), .B(n3244), .Z(n3320) );
  NANDN U3497 ( .A(n3247), .B(n3246), .Z(n3251) );
  NAND U3498 ( .A(n3249), .B(n3248), .Z(n3250) );
  AND U3499 ( .A(n3251), .B(n3250), .Z(n3386) );
  NANDN U3500 ( .A(n3253), .B(n3252), .Z(n3257) );
  NANDN U3501 ( .A(n3255), .B(n3254), .Z(n3256) );
  AND U3502 ( .A(n3257), .B(n3256), .Z(n3352) );
  NAND U3503 ( .A(b[0]), .B(a[50]), .Z(n3258) );
  XNOR U3504 ( .A(b[1]), .B(n3258), .Z(n3260) );
  NANDN U3505 ( .A(b[0]), .B(a[49]), .Z(n3259) );
  NAND U3506 ( .A(n3260), .B(n3259), .Z(n3332) );
  NAND U3507 ( .A(n5012), .B(n3261), .Z(n3263) );
  XOR U3508 ( .A(b[13]), .B(a[38]), .Z(n3338) );
  NAND U3509 ( .A(n4985), .B(n3338), .Z(n3262) );
  AND U3510 ( .A(n3263), .B(n3262), .Z(n3330) );
  AND U3511 ( .A(b[15]), .B(a[34]), .Z(n3329) );
  XNOR U3512 ( .A(n3330), .B(n3329), .Z(n3331) );
  XNOR U3513 ( .A(n3332), .B(n3331), .Z(n3350) );
  NAND U3514 ( .A(n36), .B(n3264), .Z(n3266) );
  XOR U3515 ( .A(b[5]), .B(a[46]), .Z(n3341) );
  NAND U3516 ( .A(n4560), .B(n3341), .Z(n3265) );
  AND U3517 ( .A(n3266), .B(n3265), .Z(n3374) );
  NAND U3518 ( .A(n4755), .B(n3267), .Z(n3269) );
  XOR U3519 ( .A(b[7]), .B(a[44]), .Z(n3344) );
  NAND U3520 ( .A(n4708), .B(n3344), .Z(n3268) );
  AND U3521 ( .A(n3269), .B(n3268), .Z(n3372) );
  NAND U3522 ( .A(n4471), .B(n3270), .Z(n3272) );
  XOR U3523 ( .A(b[3]), .B(a[48]), .Z(n3347) );
  NAND U3524 ( .A(n33), .B(n3347), .Z(n3271) );
  NAND U3525 ( .A(n3272), .B(n3271), .Z(n3371) );
  XNOR U3526 ( .A(n3372), .B(n3371), .Z(n3373) );
  XOR U3527 ( .A(n3374), .B(n3373), .Z(n3351) );
  XOR U3528 ( .A(n3350), .B(n3351), .Z(n3353) );
  XOR U3529 ( .A(n3352), .B(n3353), .Z(n3324) );
  NANDN U3530 ( .A(n3274), .B(n3273), .Z(n3278) );
  OR U3531 ( .A(n3276), .B(n3275), .Z(n3277) );
  AND U3532 ( .A(n3278), .B(n3277), .Z(n3323) );
  XNOR U3533 ( .A(n3324), .B(n3323), .Z(n3326) );
  NAND U3534 ( .A(n4950), .B(n3279), .Z(n3281) );
  XOR U3535 ( .A(b[11]), .B(a[40]), .Z(n3356) );
  NAND U3536 ( .A(n4863), .B(n3356), .Z(n3280) );
  AND U3537 ( .A(n3281), .B(n3280), .Z(n3367) );
  NAND U3538 ( .A(n42), .B(n3282), .Z(n3284) );
  XOR U3539 ( .A(b[15]), .B(a[36]), .Z(n3359) );
  NAND U3540 ( .A(n4981), .B(n3359), .Z(n3283) );
  AND U3541 ( .A(n3284), .B(n3283), .Z(n3366) );
  NAND U3542 ( .A(n41), .B(n3285), .Z(n3287) );
  XOR U3543 ( .A(b[9]), .B(a[42]), .Z(n3362) );
  NAND U3544 ( .A(n4810), .B(n3362), .Z(n3286) );
  NAND U3545 ( .A(n3287), .B(n3286), .Z(n3365) );
  XOR U3546 ( .A(n3366), .B(n3365), .Z(n3368) );
  XOR U3547 ( .A(n3367), .B(n3368), .Z(n3378) );
  NANDN U3548 ( .A(n3289), .B(n3288), .Z(n3293) );
  OR U3549 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3550 ( .A(n3293), .B(n3292), .Z(n3377) );
  XNOR U3551 ( .A(n3378), .B(n3377), .Z(n3379) );
  NANDN U3552 ( .A(n3295), .B(n3294), .Z(n3299) );
  NANDN U3553 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3554 ( .A(n3299), .B(n3298), .Z(n3380) );
  XNOR U3555 ( .A(n3379), .B(n3380), .Z(n3325) );
  XOR U3556 ( .A(n3326), .B(n3325), .Z(n3384) );
  NANDN U3557 ( .A(n3301), .B(n3300), .Z(n3305) );
  NANDN U3558 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U3559 ( .A(n3305), .B(n3304), .Z(n3383) );
  XNOR U3560 ( .A(n3384), .B(n3383), .Z(n3385) );
  XOR U3561 ( .A(n3386), .B(n3385), .Z(n3318) );
  NANDN U3562 ( .A(n3307), .B(n3306), .Z(n3311) );
  NAND U3563 ( .A(n3309), .B(n3308), .Z(n3310) );
  AND U3564 ( .A(n3311), .B(n3310), .Z(n3317) );
  XNOR U3565 ( .A(n3318), .B(n3317), .Z(n3319) );
  XNOR U3566 ( .A(n3320), .B(n3319), .Z(n3389) );
  XNOR U3567 ( .A(sreg[98]), .B(n3389), .Z(n3391) );
  NANDN U3568 ( .A(sreg[97]), .B(n3312), .Z(n3316) );
  NAND U3569 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U3570 ( .A(n3316), .B(n3315), .Z(n3390) );
  XNOR U3571 ( .A(n3391), .B(n3390), .Z(c[98]) );
  NANDN U3572 ( .A(n3318), .B(n3317), .Z(n3322) );
  NANDN U3573 ( .A(n3320), .B(n3319), .Z(n3321) );
  AND U3574 ( .A(n3322), .B(n3321), .Z(n3397) );
  NANDN U3575 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U3576 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U3577 ( .A(n3328), .B(n3327), .Z(n3463) );
  NANDN U3578 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U3579 ( .A(n3332), .B(n3331), .Z(n3333) );
  AND U3580 ( .A(n3334), .B(n3333), .Z(n3429) );
  NAND U3581 ( .A(b[0]), .B(a[51]), .Z(n3335) );
  XNOR U3582 ( .A(b[1]), .B(n3335), .Z(n3337) );
  NANDN U3583 ( .A(b[0]), .B(a[50]), .Z(n3336) );
  NAND U3584 ( .A(n3337), .B(n3336), .Z(n3409) );
  NAND U3585 ( .A(n5012), .B(n3338), .Z(n3340) );
  XOR U3586 ( .A(b[13]), .B(a[39]), .Z(n3415) );
  NAND U3587 ( .A(n4985), .B(n3415), .Z(n3339) );
  AND U3588 ( .A(n3340), .B(n3339), .Z(n3407) );
  AND U3589 ( .A(b[15]), .B(a[35]), .Z(n3406) );
  XNOR U3590 ( .A(n3407), .B(n3406), .Z(n3408) );
  XNOR U3591 ( .A(n3409), .B(n3408), .Z(n3427) );
  NAND U3592 ( .A(n36), .B(n3341), .Z(n3343) );
  XOR U3593 ( .A(b[5]), .B(a[47]), .Z(n3418) );
  NAND U3594 ( .A(n4560), .B(n3418), .Z(n3342) );
  AND U3595 ( .A(n3343), .B(n3342), .Z(n3451) );
  NAND U3596 ( .A(n4755), .B(n3344), .Z(n3346) );
  XOR U3597 ( .A(b[7]), .B(a[45]), .Z(n3421) );
  NAND U3598 ( .A(n4708), .B(n3421), .Z(n3345) );
  AND U3599 ( .A(n3346), .B(n3345), .Z(n3449) );
  NAND U3600 ( .A(n4471), .B(n3347), .Z(n3349) );
  XOR U3601 ( .A(b[3]), .B(a[49]), .Z(n3424) );
  NAND U3602 ( .A(n33), .B(n3424), .Z(n3348) );
  NAND U3603 ( .A(n3349), .B(n3348), .Z(n3448) );
  XNOR U3604 ( .A(n3449), .B(n3448), .Z(n3450) );
  XOR U3605 ( .A(n3451), .B(n3450), .Z(n3428) );
  XOR U3606 ( .A(n3427), .B(n3428), .Z(n3430) );
  XOR U3607 ( .A(n3429), .B(n3430), .Z(n3401) );
  NANDN U3608 ( .A(n3351), .B(n3350), .Z(n3355) );
  OR U3609 ( .A(n3353), .B(n3352), .Z(n3354) );
  AND U3610 ( .A(n3355), .B(n3354), .Z(n3400) );
  XNOR U3611 ( .A(n3401), .B(n3400), .Z(n3403) );
  NAND U3612 ( .A(n4950), .B(n3356), .Z(n3358) );
  XOR U3613 ( .A(b[11]), .B(a[41]), .Z(n3433) );
  NAND U3614 ( .A(n4863), .B(n3433), .Z(n3357) );
  AND U3615 ( .A(n3358), .B(n3357), .Z(n3444) );
  NAND U3616 ( .A(n42), .B(n3359), .Z(n3361) );
  XOR U3617 ( .A(b[15]), .B(a[37]), .Z(n3436) );
  NAND U3618 ( .A(n4981), .B(n3436), .Z(n3360) );
  AND U3619 ( .A(n3361), .B(n3360), .Z(n3443) );
  NAND U3620 ( .A(n41), .B(n3362), .Z(n3364) );
  XOR U3621 ( .A(b[9]), .B(a[43]), .Z(n3439) );
  NAND U3622 ( .A(n4810), .B(n3439), .Z(n3363) );
  NAND U3623 ( .A(n3364), .B(n3363), .Z(n3442) );
  XOR U3624 ( .A(n3443), .B(n3442), .Z(n3445) );
  XOR U3625 ( .A(n3444), .B(n3445), .Z(n3455) );
  NANDN U3626 ( .A(n3366), .B(n3365), .Z(n3370) );
  OR U3627 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3628 ( .A(n3370), .B(n3369), .Z(n3454) );
  XNOR U3629 ( .A(n3455), .B(n3454), .Z(n3456) );
  NANDN U3630 ( .A(n3372), .B(n3371), .Z(n3376) );
  NANDN U3631 ( .A(n3374), .B(n3373), .Z(n3375) );
  NAND U3632 ( .A(n3376), .B(n3375), .Z(n3457) );
  XNOR U3633 ( .A(n3456), .B(n3457), .Z(n3402) );
  XOR U3634 ( .A(n3403), .B(n3402), .Z(n3461) );
  NANDN U3635 ( .A(n3378), .B(n3377), .Z(n3382) );
  NANDN U3636 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U3637 ( .A(n3382), .B(n3381), .Z(n3460) );
  XNOR U3638 ( .A(n3461), .B(n3460), .Z(n3462) );
  XOR U3639 ( .A(n3463), .B(n3462), .Z(n3395) );
  NANDN U3640 ( .A(n3384), .B(n3383), .Z(n3388) );
  NAND U3641 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U3642 ( .A(n3388), .B(n3387), .Z(n3394) );
  XNOR U3643 ( .A(n3395), .B(n3394), .Z(n3396) );
  XNOR U3644 ( .A(n3397), .B(n3396), .Z(n3466) );
  XNOR U3645 ( .A(sreg[99]), .B(n3466), .Z(n3468) );
  NANDN U3646 ( .A(sreg[98]), .B(n3389), .Z(n3393) );
  NAND U3647 ( .A(n3391), .B(n3390), .Z(n3392) );
  NAND U3648 ( .A(n3393), .B(n3392), .Z(n3467) );
  XNOR U3649 ( .A(n3468), .B(n3467), .Z(c[99]) );
  NANDN U3650 ( .A(n3395), .B(n3394), .Z(n3399) );
  NANDN U3651 ( .A(n3397), .B(n3396), .Z(n3398) );
  AND U3652 ( .A(n3399), .B(n3398), .Z(n3474) );
  NANDN U3653 ( .A(n3401), .B(n3400), .Z(n3405) );
  NAND U3654 ( .A(n3403), .B(n3402), .Z(n3404) );
  AND U3655 ( .A(n3405), .B(n3404), .Z(n3540) );
  NANDN U3656 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U3657 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U3658 ( .A(n3411), .B(n3410), .Z(n3506) );
  NAND U3659 ( .A(b[0]), .B(a[52]), .Z(n3412) );
  XNOR U3660 ( .A(b[1]), .B(n3412), .Z(n3414) );
  NANDN U3661 ( .A(b[0]), .B(a[51]), .Z(n3413) );
  NAND U3662 ( .A(n3414), .B(n3413), .Z(n3486) );
  NAND U3663 ( .A(n5012), .B(n3415), .Z(n3417) );
  XOR U3664 ( .A(b[13]), .B(a[40]), .Z(n3492) );
  NAND U3665 ( .A(n4985), .B(n3492), .Z(n3416) );
  AND U3666 ( .A(n3417), .B(n3416), .Z(n3484) );
  AND U3667 ( .A(b[15]), .B(a[36]), .Z(n3483) );
  XNOR U3668 ( .A(n3484), .B(n3483), .Z(n3485) );
  XNOR U3669 ( .A(n3486), .B(n3485), .Z(n3504) );
  NAND U3670 ( .A(n36), .B(n3418), .Z(n3420) );
  XOR U3671 ( .A(b[5]), .B(a[48]), .Z(n3495) );
  NAND U3672 ( .A(n4560), .B(n3495), .Z(n3419) );
  AND U3673 ( .A(n3420), .B(n3419), .Z(n3528) );
  NAND U3674 ( .A(n4755), .B(n3421), .Z(n3423) );
  XOR U3675 ( .A(b[7]), .B(a[46]), .Z(n3498) );
  NAND U3676 ( .A(n4708), .B(n3498), .Z(n3422) );
  AND U3677 ( .A(n3423), .B(n3422), .Z(n3526) );
  NAND U3678 ( .A(n4471), .B(n3424), .Z(n3426) );
  XOR U3679 ( .A(b[3]), .B(a[50]), .Z(n3501) );
  NAND U3680 ( .A(n33), .B(n3501), .Z(n3425) );
  NAND U3681 ( .A(n3426), .B(n3425), .Z(n3525) );
  XNOR U3682 ( .A(n3526), .B(n3525), .Z(n3527) );
  XOR U3683 ( .A(n3528), .B(n3527), .Z(n3505) );
  XOR U3684 ( .A(n3504), .B(n3505), .Z(n3507) );
  XOR U3685 ( .A(n3506), .B(n3507), .Z(n3478) );
  NANDN U3686 ( .A(n3428), .B(n3427), .Z(n3432) );
  OR U3687 ( .A(n3430), .B(n3429), .Z(n3431) );
  AND U3688 ( .A(n3432), .B(n3431), .Z(n3477) );
  XNOR U3689 ( .A(n3478), .B(n3477), .Z(n3480) );
  NAND U3690 ( .A(n4950), .B(n3433), .Z(n3435) );
  XOR U3691 ( .A(b[11]), .B(a[42]), .Z(n3510) );
  NAND U3692 ( .A(n4863), .B(n3510), .Z(n3434) );
  AND U3693 ( .A(n3435), .B(n3434), .Z(n3521) );
  NAND U3694 ( .A(n42), .B(n3436), .Z(n3438) );
  XOR U3695 ( .A(b[15]), .B(a[38]), .Z(n3513) );
  NAND U3696 ( .A(n4981), .B(n3513), .Z(n3437) );
  AND U3697 ( .A(n3438), .B(n3437), .Z(n3520) );
  NAND U3698 ( .A(n41), .B(n3439), .Z(n3441) );
  XOR U3699 ( .A(b[9]), .B(a[44]), .Z(n3516) );
  NAND U3700 ( .A(n4810), .B(n3516), .Z(n3440) );
  NAND U3701 ( .A(n3441), .B(n3440), .Z(n3519) );
  XOR U3702 ( .A(n3520), .B(n3519), .Z(n3522) );
  XOR U3703 ( .A(n3521), .B(n3522), .Z(n3532) );
  NANDN U3704 ( .A(n3443), .B(n3442), .Z(n3447) );
  OR U3705 ( .A(n3445), .B(n3444), .Z(n3446) );
  AND U3706 ( .A(n3447), .B(n3446), .Z(n3531) );
  XNOR U3707 ( .A(n3532), .B(n3531), .Z(n3533) );
  NANDN U3708 ( .A(n3449), .B(n3448), .Z(n3453) );
  NANDN U3709 ( .A(n3451), .B(n3450), .Z(n3452) );
  NAND U3710 ( .A(n3453), .B(n3452), .Z(n3534) );
  XNOR U3711 ( .A(n3533), .B(n3534), .Z(n3479) );
  XOR U3712 ( .A(n3480), .B(n3479), .Z(n3538) );
  NANDN U3713 ( .A(n3455), .B(n3454), .Z(n3459) );
  NANDN U3714 ( .A(n3457), .B(n3456), .Z(n3458) );
  AND U3715 ( .A(n3459), .B(n3458), .Z(n3537) );
  XNOR U3716 ( .A(n3538), .B(n3537), .Z(n3539) );
  XOR U3717 ( .A(n3540), .B(n3539), .Z(n3472) );
  NANDN U3718 ( .A(n3461), .B(n3460), .Z(n3465) );
  NAND U3719 ( .A(n3463), .B(n3462), .Z(n3464) );
  AND U3720 ( .A(n3465), .B(n3464), .Z(n3471) );
  XNOR U3721 ( .A(n3472), .B(n3471), .Z(n3473) );
  XNOR U3722 ( .A(n3474), .B(n3473), .Z(n3543) );
  XNOR U3723 ( .A(sreg[100]), .B(n3543), .Z(n3545) );
  NANDN U3724 ( .A(sreg[99]), .B(n3466), .Z(n3470) );
  NAND U3725 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U3726 ( .A(n3470), .B(n3469), .Z(n3544) );
  XNOR U3727 ( .A(n3545), .B(n3544), .Z(c[100]) );
  NANDN U3728 ( .A(n3472), .B(n3471), .Z(n3476) );
  NANDN U3729 ( .A(n3474), .B(n3473), .Z(n3475) );
  AND U3730 ( .A(n3476), .B(n3475), .Z(n3551) );
  NANDN U3731 ( .A(n3478), .B(n3477), .Z(n3482) );
  NAND U3732 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U3733 ( .A(n3482), .B(n3481), .Z(n3617) );
  NANDN U3734 ( .A(n3484), .B(n3483), .Z(n3488) );
  NANDN U3735 ( .A(n3486), .B(n3485), .Z(n3487) );
  AND U3736 ( .A(n3488), .B(n3487), .Z(n3583) );
  NAND U3737 ( .A(b[0]), .B(a[53]), .Z(n3489) );
  XNOR U3738 ( .A(b[1]), .B(n3489), .Z(n3491) );
  NANDN U3739 ( .A(b[0]), .B(a[52]), .Z(n3490) );
  NAND U3740 ( .A(n3491), .B(n3490), .Z(n3563) );
  NAND U3741 ( .A(n5012), .B(n3492), .Z(n3494) );
  XOR U3742 ( .A(b[13]), .B(a[41]), .Z(n3569) );
  NAND U3743 ( .A(n4985), .B(n3569), .Z(n3493) );
  AND U3744 ( .A(n3494), .B(n3493), .Z(n3561) );
  AND U3745 ( .A(b[15]), .B(a[37]), .Z(n3560) );
  XNOR U3746 ( .A(n3561), .B(n3560), .Z(n3562) );
  XNOR U3747 ( .A(n3563), .B(n3562), .Z(n3581) );
  NAND U3748 ( .A(n36), .B(n3495), .Z(n3497) );
  XOR U3749 ( .A(b[5]), .B(a[49]), .Z(n3572) );
  NAND U3750 ( .A(n4560), .B(n3572), .Z(n3496) );
  AND U3751 ( .A(n3497), .B(n3496), .Z(n3605) );
  NAND U3752 ( .A(n4755), .B(n3498), .Z(n3500) );
  XOR U3753 ( .A(b[7]), .B(a[47]), .Z(n3575) );
  NAND U3754 ( .A(n4708), .B(n3575), .Z(n3499) );
  AND U3755 ( .A(n3500), .B(n3499), .Z(n3603) );
  NAND U3756 ( .A(n4471), .B(n3501), .Z(n3503) );
  XOR U3757 ( .A(b[3]), .B(a[51]), .Z(n3578) );
  NAND U3758 ( .A(n33), .B(n3578), .Z(n3502) );
  NAND U3759 ( .A(n3503), .B(n3502), .Z(n3602) );
  XNOR U3760 ( .A(n3603), .B(n3602), .Z(n3604) );
  XOR U3761 ( .A(n3605), .B(n3604), .Z(n3582) );
  XOR U3762 ( .A(n3581), .B(n3582), .Z(n3584) );
  XOR U3763 ( .A(n3583), .B(n3584), .Z(n3555) );
  NANDN U3764 ( .A(n3505), .B(n3504), .Z(n3509) );
  OR U3765 ( .A(n3507), .B(n3506), .Z(n3508) );
  AND U3766 ( .A(n3509), .B(n3508), .Z(n3554) );
  XNOR U3767 ( .A(n3555), .B(n3554), .Z(n3557) );
  NAND U3768 ( .A(n4950), .B(n3510), .Z(n3512) );
  XOR U3769 ( .A(b[11]), .B(a[43]), .Z(n3587) );
  NAND U3770 ( .A(n4863), .B(n3587), .Z(n3511) );
  AND U3771 ( .A(n3512), .B(n3511), .Z(n3598) );
  NAND U3772 ( .A(n42), .B(n3513), .Z(n3515) );
  XOR U3773 ( .A(b[15]), .B(a[39]), .Z(n3590) );
  NAND U3774 ( .A(n4981), .B(n3590), .Z(n3514) );
  AND U3775 ( .A(n3515), .B(n3514), .Z(n3597) );
  NAND U3776 ( .A(n41), .B(n3516), .Z(n3518) );
  XOR U3777 ( .A(b[9]), .B(a[45]), .Z(n3593) );
  NAND U3778 ( .A(n4810), .B(n3593), .Z(n3517) );
  NAND U3779 ( .A(n3518), .B(n3517), .Z(n3596) );
  XOR U3780 ( .A(n3597), .B(n3596), .Z(n3599) );
  XOR U3781 ( .A(n3598), .B(n3599), .Z(n3609) );
  NANDN U3782 ( .A(n3520), .B(n3519), .Z(n3524) );
  OR U3783 ( .A(n3522), .B(n3521), .Z(n3523) );
  AND U3784 ( .A(n3524), .B(n3523), .Z(n3608) );
  XNOR U3785 ( .A(n3609), .B(n3608), .Z(n3610) );
  NANDN U3786 ( .A(n3526), .B(n3525), .Z(n3530) );
  NANDN U3787 ( .A(n3528), .B(n3527), .Z(n3529) );
  NAND U3788 ( .A(n3530), .B(n3529), .Z(n3611) );
  XNOR U3789 ( .A(n3610), .B(n3611), .Z(n3556) );
  XOR U3790 ( .A(n3557), .B(n3556), .Z(n3615) );
  NANDN U3791 ( .A(n3532), .B(n3531), .Z(n3536) );
  NANDN U3792 ( .A(n3534), .B(n3533), .Z(n3535) );
  AND U3793 ( .A(n3536), .B(n3535), .Z(n3614) );
  XNOR U3794 ( .A(n3615), .B(n3614), .Z(n3616) );
  XOR U3795 ( .A(n3617), .B(n3616), .Z(n3549) );
  NANDN U3796 ( .A(n3538), .B(n3537), .Z(n3542) );
  NAND U3797 ( .A(n3540), .B(n3539), .Z(n3541) );
  AND U3798 ( .A(n3542), .B(n3541), .Z(n3548) );
  XNOR U3799 ( .A(n3549), .B(n3548), .Z(n3550) );
  XNOR U3800 ( .A(n3551), .B(n3550), .Z(n3620) );
  XNOR U3801 ( .A(sreg[101]), .B(n3620), .Z(n3622) );
  NANDN U3802 ( .A(sreg[100]), .B(n3543), .Z(n3547) );
  NAND U3803 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U3804 ( .A(n3547), .B(n3546), .Z(n3621) );
  XNOR U3805 ( .A(n3622), .B(n3621), .Z(c[101]) );
  NANDN U3806 ( .A(n3549), .B(n3548), .Z(n3553) );
  NANDN U3807 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U3808 ( .A(n3553), .B(n3552), .Z(n3628) );
  NANDN U3809 ( .A(n3555), .B(n3554), .Z(n3559) );
  NAND U3810 ( .A(n3557), .B(n3556), .Z(n3558) );
  AND U3811 ( .A(n3559), .B(n3558), .Z(n3694) );
  NANDN U3812 ( .A(n3561), .B(n3560), .Z(n3565) );
  NANDN U3813 ( .A(n3563), .B(n3562), .Z(n3564) );
  AND U3814 ( .A(n3565), .B(n3564), .Z(n3660) );
  NAND U3815 ( .A(b[0]), .B(a[54]), .Z(n3566) );
  XNOR U3816 ( .A(b[1]), .B(n3566), .Z(n3568) );
  NANDN U3817 ( .A(b[0]), .B(a[53]), .Z(n3567) );
  NAND U3818 ( .A(n3568), .B(n3567), .Z(n3640) );
  NAND U3819 ( .A(n5012), .B(n3569), .Z(n3571) );
  XOR U3820 ( .A(b[13]), .B(a[42]), .Z(n3646) );
  NAND U3821 ( .A(n4985), .B(n3646), .Z(n3570) );
  AND U3822 ( .A(n3571), .B(n3570), .Z(n3638) );
  AND U3823 ( .A(b[15]), .B(a[38]), .Z(n3637) );
  XNOR U3824 ( .A(n3638), .B(n3637), .Z(n3639) );
  XNOR U3825 ( .A(n3640), .B(n3639), .Z(n3658) );
  NAND U3826 ( .A(n36), .B(n3572), .Z(n3574) );
  XOR U3827 ( .A(b[5]), .B(a[50]), .Z(n3649) );
  NAND U3828 ( .A(n4560), .B(n3649), .Z(n3573) );
  AND U3829 ( .A(n3574), .B(n3573), .Z(n3682) );
  NAND U3830 ( .A(n4755), .B(n3575), .Z(n3577) );
  XOR U3831 ( .A(b[7]), .B(a[48]), .Z(n3652) );
  NAND U3832 ( .A(n4708), .B(n3652), .Z(n3576) );
  AND U3833 ( .A(n3577), .B(n3576), .Z(n3680) );
  NAND U3834 ( .A(n4471), .B(n3578), .Z(n3580) );
  XOR U3835 ( .A(a[52]), .B(b[3]), .Z(n3655) );
  NAND U3836 ( .A(n33), .B(n3655), .Z(n3579) );
  NAND U3837 ( .A(n3580), .B(n3579), .Z(n3679) );
  XNOR U3838 ( .A(n3680), .B(n3679), .Z(n3681) );
  XOR U3839 ( .A(n3682), .B(n3681), .Z(n3659) );
  XOR U3840 ( .A(n3658), .B(n3659), .Z(n3661) );
  XOR U3841 ( .A(n3660), .B(n3661), .Z(n3632) );
  NANDN U3842 ( .A(n3582), .B(n3581), .Z(n3586) );
  OR U3843 ( .A(n3584), .B(n3583), .Z(n3585) );
  AND U3844 ( .A(n3586), .B(n3585), .Z(n3631) );
  XNOR U3845 ( .A(n3632), .B(n3631), .Z(n3634) );
  NAND U3846 ( .A(n4950), .B(n3587), .Z(n3589) );
  XOR U3847 ( .A(b[11]), .B(a[44]), .Z(n3664) );
  NAND U3848 ( .A(n4863), .B(n3664), .Z(n3588) );
  AND U3849 ( .A(n3589), .B(n3588), .Z(n3675) );
  NAND U3850 ( .A(n42), .B(n3590), .Z(n3592) );
  XOR U3851 ( .A(b[15]), .B(a[40]), .Z(n3667) );
  NAND U3852 ( .A(n4981), .B(n3667), .Z(n3591) );
  AND U3853 ( .A(n3592), .B(n3591), .Z(n3674) );
  NAND U3854 ( .A(n41), .B(n3593), .Z(n3595) );
  XOR U3855 ( .A(b[9]), .B(a[46]), .Z(n3670) );
  NAND U3856 ( .A(n4810), .B(n3670), .Z(n3594) );
  NAND U3857 ( .A(n3595), .B(n3594), .Z(n3673) );
  XOR U3858 ( .A(n3674), .B(n3673), .Z(n3676) );
  XOR U3859 ( .A(n3675), .B(n3676), .Z(n3686) );
  NANDN U3860 ( .A(n3597), .B(n3596), .Z(n3601) );
  OR U3861 ( .A(n3599), .B(n3598), .Z(n3600) );
  AND U3862 ( .A(n3601), .B(n3600), .Z(n3685) );
  XNOR U3863 ( .A(n3686), .B(n3685), .Z(n3687) );
  NANDN U3864 ( .A(n3603), .B(n3602), .Z(n3607) );
  NANDN U3865 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U3866 ( .A(n3607), .B(n3606), .Z(n3688) );
  XNOR U3867 ( .A(n3687), .B(n3688), .Z(n3633) );
  XOR U3868 ( .A(n3634), .B(n3633), .Z(n3692) );
  NANDN U3869 ( .A(n3609), .B(n3608), .Z(n3613) );
  NANDN U3870 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U3871 ( .A(n3613), .B(n3612), .Z(n3691) );
  XNOR U3872 ( .A(n3692), .B(n3691), .Z(n3693) );
  XOR U3873 ( .A(n3694), .B(n3693), .Z(n3626) );
  NANDN U3874 ( .A(n3615), .B(n3614), .Z(n3619) );
  NAND U3875 ( .A(n3617), .B(n3616), .Z(n3618) );
  AND U3876 ( .A(n3619), .B(n3618), .Z(n3625) );
  XNOR U3877 ( .A(n3626), .B(n3625), .Z(n3627) );
  XNOR U3878 ( .A(n3628), .B(n3627), .Z(n3697) );
  XNOR U3879 ( .A(sreg[102]), .B(n3697), .Z(n3699) );
  NANDN U3880 ( .A(sreg[101]), .B(n3620), .Z(n3624) );
  NAND U3881 ( .A(n3622), .B(n3621), .Z(n3623) );
  NAND U3882 ( .A(n3624), .B(n3623), .Z(n3698) );
  XNOR U3883 ( .A(n3699), .B(n3698), .Z(c[102]) );
  NANDN U3884 ( .A(n3626), .B(n3625), .Z(n3630) );
  NANDN U3885 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U3886 ( .A(n3630), .B(n3629), .Z(n3705) );
  NANDN U3887 ( .A(n3632), .B(n3631), .Z(n3636) );
  NAND U3888 ( .A(n3634), .B(n3633), .Z(n3635) );
  AND U3889 ( .A(n3636), .B(n3635), .Z(n3771) );
  NANDN U3890 ( .A(n3638), .B(n3637), .Z(n3642) );
  NANDN U3891 ( .A(n3640), .B(n3639), .Z(n3641) );
  AND U3892 ( .A(n3642), .B(n3641), .Z(n3737) );
  NAND U3893 ( .A(b[0]), .B(a[55]), .Z(n3643) );
  XNOR U3894 ( .A(b[1]), .B(n3643), .Z(n3645) );
  NANDN U3895 ( .A(b[0]), .B(a[54]), .Z(n3644) );
  NAND U3896 ( .A(n3645), .B(n3644), .Z(n3717) );
  NAND U3897 ( .A(n5012), .B(n3646), .Z(n3648) );
  XOR U3898 ( .A(b[13]), .B(a[43]), .Z(n3723) );
  NAND U3899 ( .A(n4985), .B(n3723), .Z(n3647) );
  AND U3900 ( .A(n3648), .B(n3647), .Z(n3715) );
  AND U3901 ( .A(b[15]), .B(a[39]), .Z(n3714) );
  XNOR U3902 ( .A(n3715), .B(n3714), .Z(n3716) );
  XNOR U3903 ( .A(n3717), .B(n3716), .Z(n3735) );
  NAND U3904 ( .A(n36), .B(n3649), .Z(n3651) );
  XOR U3905 ( .A(b[5]), .B(a[51]), .Z(n3726) );
  NAND U3906 ( .A(n4560), .B(n3726), .Z(n3650) );
  AND U3907 ( .A(n3651), .B(n3650), .Z(n3759) );
  NAND U3908 ( .A(n4755), .B(n3652), .Z(n3654) );
  XOR U3909 ( .A(b[7]), .B(a[49]), .Z(n3729) );
  NAND U3910 ( .A(n4708), .B(n3729), .Z(n3653) );
  AND U3911 ( .A(n3654), .B(n3653), .Z(n3757) );
  NAND U3912 ( .A(n4471), .B(n3655), .Z(n3657) );
  XOR U3913 ( .A(b[3]), .B(a[53]), .Z(n3732) );
  NAND U3914 ( .A(n33), .B(n3732), .Z(n3656) );
  NAND U3915 ( .A(n3657), .B(n3656), .Z(n3756) );
  XNOR U3916 ( .A(n3757), .B(n3756), .Z(n3758) );
  XOR U3917 ( .A(n3759), .B(n3758), .Z(n3736) );
  XOR U3918 ( .A(n3735), .B(n3736), .Z(n3738) );
  XOR U3919 ( .A(n3737), .B(n3738), .Z(n3709) );
  NANDN U3920 ( .A(n3659), .B(n3658), .Z(n3663) );
  OR U3921 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U3922 ( .A(n3663), .B(n3662), .Z(n3708) );
  XNOR U3923 ( .A(n3709), .B(n3708), .Z(n3711) );
  NAND U3924 ( .A(n4950), .B(n3664), .Z(n3666) );
  XOR U3925 ( .A(b[11]), .B(a[45]), .Z(n3741) );
  NAND U3926 ( .A(n4863), .B(n3741), .Z(n3665) );
  AND U3927 ( .A(n3666), .B(n3665), .Z(n3752) );
  NAND U3928 ( .A(n42), .B(n3667), .Z(n3669) );
  XOR U3929 ( .A(b[15]), .B(a[41]), .Z(n3744) );
  NAND U3930 ( .A(n4981), .B(n3744), .Z(n3668) );
  AND U3931 ( .A(n3669), .B(n3668), .Z(n3751) );
  NAND U3932 ( .A(n41), .B(n3670), .Z(n3672) );
  XOR U3933 ( .A(b[9]), .B(a[47]), .Z(n3747) );
  NAND U3934 ( .A(n4810), .B(n3747), .Z(n3671) );
  NAND U3935 ( .A(n3672), .B(n3671), .Z(n3750) );
  XOR U3936 ( .A(n3751), .B(n3750), .Z(n3753) );
  XOR U3937 ( .A(n3752), .B(n3753), .Z(n3763) );
  NANDN U3938 ( .A(n3674), .B(n3673), .Z(n3678) );
  OR U3939 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U3940 ( .A(n3678), .B(n3677), .Z(n3762) );
  XNOR U3941 ( .A(n3763), .B(n3762), .Z(n3764) );
  NANDN U3942 ( .A(n3680), .B(n3679), .Z(n3684) );
  NANDN U3943 ( .A(n3682), .B(n3681), .Z(n3683) );
  NAND U3944 ( .A(n3684), .B(n3683), .Z(n3765) );
  XNOR U3945 ( .A(n3764), .B(n3765), .Z(n3710) );
  XOR U3946 ( .A(n3711), .B(n3710), .Z(n3769) );
  NANDN U3947 ( .A(n3686), .B(n3685), .Z(n3690) );
  NANDN U3948 ( .A(n3688), .B(n3687), .Z(n3689) );
  AND U3949 ( .A(n3690), .B(n3689), .Z(n3768) );
  XNOR U3950 ( .A(n3769), .B(n3768), .Z(n3770) );
  XOR U3951 ( .A(n3771), .B(n3770), .Z(n3703) );
  NANDN U3952 ( .A(n3692), .B(n3691), .Z(n3696) );
  NAND U3953 ( .A(n3694), .B(n3693), .Z(n3695) );
  AND U3954 ( .A(n3696), .B(n3695), .Z(n3702) );
  XNOR U3955 ( .A(n3703), .B(n3702), .Z(n3704) );
  XNOR U3956 ( .A(n3705), .B(n3704), .Z(n3774) );
  XNOR U3957 ( .A(sreg[103]), .B(n3774), .Z(n3776) );
  NANDN U3958 ( .A(sreg[102]), .B(n3697), .Z(n3701) );
  NAND U3959 ( .A(n3699), .B(n3698), .Z(n3700) );
  NAND U3960 ( .A(n3701), .B(n3700), .Z(n3775) );
  XNOR U3961 ( .A(n3776), .B(n3775), .Z(c[103]) );
  NANDN U3962 ( .A(n3703), .B(n3702), .Z(n3707) );
  NANDN U3963 ( .A(n3705), .B(n3704), .Z(n3706) );
  AND U3964 ( .A(n3707), .B(n3706), .Z(n3782) );
  NANDN U3965 ( .A(n3709), .B(n3708), .Z(n3713) );
  NAND U3966 ( .A(n3711), .B(n3710), .Z(n3712) );
  AND U3967 ( .A(n3713), .B(n3712), .Z(n3848) );
  NANDN U3968 ( .A(n3715), .B(n3714), .Z(n3719) );
  NANDN U3969 ( .A(n3717), .B(n3716), .Z(n3718) );
  AND U3970 ( .A(n3719), .B(n3718), .Z(n3835) );
  NAND U3971 ( .A(b[0]), .B(a[56]), .Z(n3720) );
  XNOR U3972 ( .A(b[1]), .B(n3720), .Z(n3722) );
  NANDN U3973 ( .A(b[0]), .B(a[55]), .Z(n3721) );
  NAND U3974 ( .A(n3722), .B(n3721), .Z(n3815) );
  NAND U3975 ( .A(n5012), .B(n3723), .Z(n3725) );
  XOR U3976 ( .A(b[13]), .B(a[44]), .Z(n3821) );
  NAND U3977 ( .A(n4985), .B(n3821), .Z(n3724) );
  AND U3978 ( .A(n3725), .B(n3724), .Z(n3813) );
  AND U3979 ( .A(b[15]), .B(a[40]), .Z(n3812) );
  XNOR U3980 ( .A(n3813), .B(n3812), .Z(n3814) );
  XNOR U3981 ( .A(n3815), .B(n3814), .Z(n3833) );
  NAND U3982 ( .A(n36), .B(n3726), .Z(n3728) );
  XOR U3983 ( .A(b[5]), .B(a[52]), .Z(n3824) );
  NAND U3984 ( .A(n4560), .B(n3824), .Z(n3727) );
  AND U3985 ( .A(n3728), .B(n3727), .Z(n3809) );
  NAND U3986 ( .A(n4755), .B(n3729), .Z(n3731) );
  XOR U3987 ( .A(b[7]), .B(a[50]), .Z(n3827) );
  NAND U3988 ( .A(n4708), .B(n3827), .Z(n3730) );
  AND U3989 ( .A(n3731), .B(n3730), .Z(n3807) );
  NAND U3990 ( .A(n4471), .B(n3732), .Z(n3734) );
  XOR U3991 ( .A(a[54]), .B(b[3]), .Z(n3830) );
  NAND U3992 ( .A(n33), .B(n3830), .Z(n3733) );
  NAND U3993 ( .A(n3734), .B(n3733), .Z(n3806) );
  XNOR U3994 ( .A(n3807), .B(n3806), .Z(n3808) );
  XOR U3995 ( .A(n3809), .B(n3808), .Z(n3834) );
  XOR U3996 ( .A(n3833), .B(n3834), .Z(n3836) );
  XOR U3997 ( .A(n3835), .B(n3836), .Z(n3786) );
  NANDN U3998 ( .A(n3736), .B(n3735), .Z(n3740) );
  OR U3999 ( .A(n3738), .B(n3737), .Z(n3739) );
  AND U4000 ( .A(n3740), .B(n3739), .Z(n3785) );
  XNOR U4001 ( .A(n3786), .B(n3785), .Z(n3788) );
  NAND U4002 ( .A(n4950), .B(n3741), .Z(n3743) );
  XOR U4003 ( .A(b[11]), .B(a[46]), .Z(n3791) );
  NAND U4004 ( .A(n4863), .B(n3791), .Z(n3742) );
  AND U4005 ( .A(n3743), .B(n3742), .Z(n3802) );
  NAND U4006 ( .A(n42), .B(n3744), .Z(n3746) );
  XOR U4007 ( .A(b[15]), .B(a[42]), .Z(n3794) );
  NAND U4008 ( .A(n4981), .B(n3794), .Z(n3745) );
  AND U4009 ( .A(n3746), .B(n3745), .Z(n3801) );
  NAND U4010 ( .A(n41), .B(n3747), .Z(n3749) );
  XOR U4011 ( .A(b[9]), .B(a[48]), .Z(n3797) );
  NAND U4012 ( .A(n4810), .B(n3797), .Z(n3748) );
  NAND U4013 ( .A(n3749), .B(n3748), .Z(n3800) );
  XOR U4014 ( .A(n3801), .B(n3800), .Z(n3803) );
  XOR U4015 ( .A(n3802), .B(n3803), .Z(n3840) );
  NANDN U4016 ( .A(n3751), .B(n3750), .Z(n3755) );
  OR U4017 ( .A(n3753), .B(n3752), .Z(n3754) );
  AND U4018 ( .A(n3755), .B(n3754), .Z(n3839) );
  XNOR U4019 ( .A(n3840), .B(n3839), .Z(n3841) );
  NANDN U4020 ( .A(n3757), .B(n3756), .Z(n3761) );
  NANDN U4021 ( .A(n3759), .B(n3758), .Z(n3760) );
  NAND U4022 ( .A(n3761), .B(n3760), .Z(n3842) );
  XNOR U4023 ( .A(n3841), .B(n3842), .Z(n3787) );
  XOR U4024 ( .A(n3788), .B(n3787), .Z(n3846) );
  NANDN U4025 ( .A(n3763), .B(n3762), .Z(n3767) );
  NANDN U4026 ( .A(n3765), .B(n3764), .Z(n3766) );
  AND U4027 ( .A(n3767), .B(n3766), .Z(n3845) );
  XNOR U4028 ( .A(n3846), .B(n3845), .Z(n3847) );
  XOR U4029 ( .A(n3848), .B(n3847), .Z(n3780) );
  NANDN U4030 ( .A(n3769), .B(n3768), .Z(n3773) );
  NAND U4031 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U4032 ( .A(n3773), .B(n3772), .Z(n3779) );
  XNOR U4033 ( .A(n3780), .B(n3779), .Z(n3781) );
  XNOR U4034 ( .A(n3782), .B(n3781), .Z(n3851) );
  XNOR U4035 ( .A(sreg[104]), .B(n3851), .Z(n3853) );
  NANDN U4036 ( .A(sreg[103]), .B(n3774), .Z(n3778) );
  NAND U4037 ( .A(n3776), .B(n3775), .Z(n3777) );
  NAND U4038 ( .A(n3778), .B(n3777), .Z(n3852) );
  XNOR U4039 ( .A(n3853), .B(n3852), .Z(c[104]) );
  NANDN U4040 ( .A(n3780), .B(n3779), .Z(n3784) );
  NANDN U4041 ( .A(n3782), .B(n3781), .Z(n3783) );
  AND U4042 ( .A(n3784), .B(n3783), .Z(n3859) );
  NANDN U4043 ( .A(n3786), .B(n3785), .Z(n3790) );
  NAND U4044 ( .A(n3788), .B(n3787), .Z(n3789) );
  AND U4045 ( .A(n3790), .B(n3789), .Z(n3925) );
  NAND U4046 ( .A(n4950), .B(n3791), .Z(n3793) );
  XOR U4047 ( .A(b[11]), .B(a[47]), .Z(n3868) );
  NAND U4048 ( .A(n4863), .B(n3868), .Z(n3792) );
  AND U4049 ( .A(n3793), .B(n3792), .Z(n3879) );
  NAND U4050 ( .A(n42), .B(n3794), .Z(n3796) );
  XOR U4051 ( .A(b[15]), .B(a[43]), .Z(n3871) );
  NAND U4052 ( .A(n4981), .B(n3871), .Z(n3795) );
  AND U4053 ( .A(n3796), .B(n3795), .Z(n3878) );
  NAND U4054 ( .A(n41), .B(n3797), .Z(n3799) );
  XOR U4055 ( .A(b[9]), .B(a[49]), .Z(n3874) );
  NAND U4056 ( .A(n4810), .B(n3874), .Z(n3798) );
  NAND U4057 ( .A(n3799), .B(n3798), .Z(n3877) );
  XOR U4058 ( .A(n3878), .B(n3877), .Z(n3880) );
  XOR U4059 ( .A(n3879), .B(n3880), .Z(n3917) );
  NANDN U4060 ( .A(n3801), .B(n3800), .Z(n3805) );
  OR U4061 ( .A(n3803), .B(n3802), .Z(n3804) );
  AND U4062 ( .A(n3805), .B(n3804), .Z(n3916) );
  XNOR U4063 ( .A(n3917), .B(n3916), .Z(n3918) );
  NANDN U4064 ( .A(n3807), .B(n3806), .Z(n3811) );
  NANDN U4065 ( .A(n3809), .B(n3808), .Z(n3810) );
  NAND U4066 ( .A(n3811), .B(n3810), .Z(n3919) );
  XNOR U4067 ( .A(n3918), .B(n3919), .Z(n3865) );
  NANDN U4068 ( .A(n3813), .B(n3812), .Z(n3817) );
  NANDN U4069 ( .A(n3815), .B(n3814), .Z(n3816) );
  AND U4070 ( .A(n3817), .B(n3816), .Z(n3912) );
  NAND U4071 ( .A(b[0]), .B(a[57]), .Z(n3818) );
  XNOR U4072 ( .A(b[1]), .B(n3818), .Z(n3820) );
  NANDN U4073 ( .A(b[0]), .B(a[56]), .Z(n3819) );
  NAND U4074 ( .A(n3820), .B(n3819), .Z(n3892) );
  NAND U4075 ( .A(n5012), .B(n3821), .Z(n3823) );
  XOR U4076 ( .A(b[13]), .B(a[45]), .Z(n3898) );
  NAND U4077 ( .A(n4985), .B(n3898), .Z(n3822) );
  AND U4078 ( .A(n3823), .B(n3822), .Z(n3890) );
  AND U4079 ( .A(b[15]), .B(a[41]), .Z(n3889) );
  XNOR U4080 ( .A(n3890), .B(n3889), .Z(n3891) );
  XNOR U4081 ( .A(n3892), .B(n3891), .Z(n3910) );
  NAND U4082 ( .A(n36), .B(n3824), .Z(n3826) );
  XOR U4083 ( .A(b[5]), .B(a[53]), .Z(n3901) );
  NAND U4084 ( .A(n4560), .B(n3901), .Z(n3825) );
  AND U4085 ( .A(n3826), .B(n3825), .Z(n3886) );
  NAND U4086 ( .A(n4755), .B(n3827), .Z(n3829) );
  XOR U4087 ( .A(b[7]), .B(a[51]), .Z(n3904) );
  NAND U4088 ( .A(n4708), .B(n3904), .Z(n3828) );
  AND U4089 ( .A(n3829), .B(n3828), .Z(n3884) );
  NAND U4090 ( .A(n4471), .B(n3830), .Z(n3832) );
  XOR U4091 ( .A(a[55]), .B(b[3]), .Z(n3907) );
  NAND U4092 ( .A(n33), .B(n3907), .Z(n3831) );
  NAND U4093 ( .A(n3832), .B(n3831), .Z(n3883) );
  XNOR U4094 ( .A(n3884), .B(n3883), .Z(n3885) );
  XOR U4095 ( .A(n3886), .B(n3885), .Z(n3911) );
  XOR U4096 ( .A(n3910), .B(n3911), .Z(n3913) );
  XOR U4097 ( .A(n3912), .B(n3913), .Z(n3863) );
  NANDN U4098 ( .A(n3834), .B(n3833), .Z(n3838) );
  OR U4099 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U4100 ( .A(n3838), .B(n3837), .Z(n3862) );
  XNOR U4101 ( .A(n3863), .B(n3862), .Z(n3864) );
  XOR U4102 ( .A(n3865), .B(n3864), .Z(n3923) );
  NANDN U4103 ( .A(n3840), .B(n3839), .Z(n3844) );
  NANDN U4104 ( .A(n3842), .B(n3841), .Z(n3843) );
  AND U4105 ( .A(n3844), .B(n3843), .Z(n3922) );
  XNOR U4106 ( .A(n3923), .B(n3922), .Z(n3924) );
  XOR U4107 ( .A(n3925), .B(n3924), .Z(n3857) );
  NANDN U4108 ( .A(n3846), .B(n3845), .Z(n3850) );
  NAND U4109 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4110 ( .A(n3850), .B(n3849), .Z(n3856) );
  XNOR U4111 ( .A(n3857), .B(n3856), .Z(n3858) );
  XNOR U4112 ( .A(n3859), .B(n3858), .Z(n3928) );
  XNOR U4113 ( .A(sreg[105]), .B(n3928), .Z(n3930) );
  NANDN U4114 ( .A(sreg[104]), .B(n3851), .Z(n3855) );
  NAND U4115 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4116 ( .A(n3855), .B(n3854), .Z(n3929) );
  XNOR U4117 ( .A(n3930), .B(n3929), .Z(c[105]) );
  NANDN U4118 ( .A(n3857), .B(n3856), .Z(n3861) );
  NANDN U4119 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U4120 ( .A(n3861), .B(n3860), .Z(n3936) );
  NANDN U4121 ( .A(n3863), .B(n3862), .Z(n3867) );
  NAND U4122 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4123 ( .A(n3867), .B(n3866), .Z(n4002) );
  NAND U4124 ( .A(n4950), .B(n3868), .Z(n3870) );
  XOR U4125 ( .A(b[11]), .B(a[48]), .Z(n3972) );
  NAND U4126 ( .A(n4863), .B(n3972), .Z(n3869) );
  AND U4127 ( .A(n3870), .B(n3869), .Z(n3983) );
  NAND U4128 ( .A(n42), .B(n3871), .Z(n3873) );
  XOR U4129 ( .A(b[15]), .B(a[44]), .Z(n3975) );
  NAND U4130 ( .A(n4981), .B(n3975), .Z(n3872) );
  AND U4131 ( .A(n3873), .B(n3872), .Z(n3982) );
  NAND U4132 ( .A(n41), .B(n3874), .Z(n3876) );
  XOR U4133 ( .A(b[9]), .B(a[50]), .Z(n3978) );
  NAND U4134 ( .A(n4810), .B(n3978), .Z(n3875) );
  NAND U4135 ( .A(n3876), .B(n3875), .Z(n3981) );
  XOR U4136 ( .A(n3982), .B(n3981), .Z(n3984) );
  XOR U4137 ( .A(n3983), .B(n3984), .Z(n3994) );
  NANDN U4138 ( .A(n3878), .B(n3877), .Z(n3882) );
  OR U4139 ( .A(n3880), .B(n3879), .Z(n3881) );
  AND U4140 ( .A(n3882), .B(n3881), .Z(n3993) );
  XNOR U4141 ( .A(n3994), .B(n3993), .Z(n3995) );
  NANDN U4142 ( .A(n3884), .B(n3883), .Z(n3888) );
  NANDN U4143 ( .A(n3886), .B(n3885), .Z(n3887) );
  NAND U4144 ( .A(n3888), .B(n3887), .Z(n3996) );
  XNOR U4145 ( .A(n3995), .B(n3996), .Z(n3942) );
  NANDN U4146 ( .A(n3890), .B(n3889), .Z(n3894) );
  NANDN U4147 ( .A(n3892), .B(n3891), .Z(n3893) );
  AND U4148 ( .A(n3894), .B(n3893), .Z(n3968) );
  NAND U4149 ( .A(b[0]), .B(a[58]), .Z(n3895) );
  XNOR U4150 ( .A(b[1]), .B(n3895), .Z(n3897) );
  NANDN U4151 ( .A(b[0]), .B(a[57]), .Z(n3896) );
  NAND U4152 ( .A(n3897), .B(n3896), .Z(n3948) );
  NAND U4153 ( .A(n5012), .B(n3898), .Z(n3900) );
  XOR U4154 ( .A(b[13]), .B(a[46]), .Z(n3951) );
  NAND U4155 ( .A(n4985), .B(n3951), .Z(n3899) );
  AND U4156 ( .A(n3900), .B(n3899), .Z(n3946) );
  AND U4157 ( .A(b[15]), .B(a[42]), .Z(n3945) );
  XNOR U4158 ( .A(n3946), .B(n3945), .Z(n3947) );
  XNOR U4159 ( .A(n3948), .B(n3947), .Z(n3966) );
  NAND U4160 ( .A(n36), .B(n3901), .Z(n3903) );
  XOR U4161 ( .A(b[5]), .B(a[54]), .Z(n3957) );
  NAND U4162 ( .A(n4560), .B(n3957), .Z(n3902) );
  AND U4163 ( .A(n3903), .B(n3902), .Z(n3990) );
  NAND U4164 ( .A(n4755), .B(n3904), .Z(n3906) );
  XOR U4165 ( .A(b[7]), .B(a[52]), .Z(n3960) );
  NAND U4166 ( .A(n4708), .B(n3960), .Z(n3905) );
  AND U4167 ( .A(n3906), .B(n3905), .Z(n3988) );
  NAND U4168 ( .A(n4471), .B(n3907), .Z(n3909) );
  XOR U4169 ( .A(a[56]), .B(b[3]), .Z(n3963) );
  NAND U4170 ( .A(n33), .B(n3963), .Z(n3908) );
  NAND U4171 ( .A(n3909), .B(n3908), .Z(n3987) );
  XNOR U4172 ( .A(n3988), .B(n3987), .Z(n3989) );
  XOR U4173 ( .A(n3990), .B(n3989), .Z(n3967) );
  XOR U4174 ( .A(n3966), .B(n3967), .Z(n3969) );
  XOR U4175 ( .A(n3968), .B(n3969), .Z(n3940) );
  NANDN U4176 ( .A(n3911), .B(n3910), .Z(n3915) );
  OR U4177 ( .A(n3913), .B(n3912), .Z(n3914) );
  AND U4178 ( .A(n3915), .B(n3914), .Z(n3939) );
  XNOR U4179 ( .A(n3940), .B(n3939), .Z(n3941) );
  XOR U4180 ( .A(n3942), .B(n3941), .Z(n4000) );
  NANDN U4181 ( .A(n3917), .B(n3916), .Z(n3921) );
  NANDN U4182 ( .A(n3919), .B(n3918), .Z(n3920) );
  AND U4183 ( .A(n3921), .B(n3920), .Z(n3999) );
  XNOR U4184 ( .A(n4000), .B(n3999), .Z(n4001) );
  XOR U4185 ( .A(n4002), .B(n4001), .Z(n3934) );
  NANDN U4186 ( .A(n3923), .B(n3922), .Z(n3927) );
  NAND U4187 ( .A(n3925), .B(n3924), .Z(n3926) );
  AND U4188 ( .A(n3927), .B(n3926), .Z(n3933) );
  XNOR U4189 ( .A(n3934), .B(n3933), .Z(n3935) );
  XNOR U4190 ( .A(n3936), .B(n3935), .Z(n4005) );
  XNOR U4191 ( .A(sreg[106]), .B(n4005), .Z(n4007) );
  NANDN U4192 ( .A(sreg[105]), .B(n3928), .Z(n3932) );
  NAND U4193 ( .A(n3930), .B(n3929), .Z(n3931) );
  NAND U4194 ( .A(n3932), .B(n3931), .Z(n4006) );
  XNOR U4195 ( .A(n4007), .B(n4006), .Z(c[106]) );
  NANDN U4196 ( .A(n3934), .B(n3933), .Z(n3938) );
  NANDN U4197 ( .A(n3936), .B(n3935), .Z(n3937) );
  AND U4198 ( .A(n3938), .B(n3937), .Z(n4013) );
  NANDN U4199 ( .A(n3940), .B(n3939), .Z(n3944) );
  NAND U4200 ( .A(n3942), .B(n3941), .Z(n3943) );
  AND U4201 ( .A(n3944), .B(n3943), .Z(n4079) );
  NANDN U4202 ( .A(n3946), .B(n3945), .Z(n3950) );
  NANDN U4203 ( .A(n3948), .B(n3947), .Z(n3949) );
  AND U4204 ( .A(n3950), .B(n3949), .Z(n4045) );
  NAND U4205 ( .A(n5012), .B(n3951), .Z(n3953) );
  XOR U4206 ( .A(b[13]), .B(a[47]), .Z(n4028) );
  NAND U4207 ( .A(n4985), .B(n4028), .Z(n3952) );
  AND U4208 ( .A(n3953), .B(n3952), .Z(n4023) );
  AND U4209 ( .A(b[15]), .B(a[43]), .Z(n4022) );
  XNOR U4210 ( .A(n4023), .B(n4022), .Z(n4024) );
  NAND U4211 ( .A(b[0]), .B(a[59]), .Z(n3954) );
  XNOR U4212 ( .A(b[1]), .B(n3954), .Z(n3956) );
  NANDN U4213 ( .A(b[0]), .B(a[58]), .Z(n3955) );
  NAND U4214 ( .A(n3956), .B(n3955), .Z(n4025) );
  XNOR U4215 ( .A(n4024), .B(n4025), .Z(n4043) );
  NAND U4216 ( .A(n36), .B(n3957), .Z(n3959) );
  XOR U4217 ( .A(a[55]), .B(b[5]), .Z(n4034) );
  NAND U4218 ( .A(n4560), .B(n4034), .Z(n3958) );
  AND U4219 ( .A(n3959), .B(n3958), .Z(n4067) );
  NAND U4220 ( .A(n4755), .B(n3960), .Z(n3962) );
  XOR U4221 ( .A(b[7]), .B(a[53]), .Z(n4037) );
  NAND U4222 ( .A(n4708), .B(n4037), .Z(n3961) );
  AND U4223 ( .A(n3962), .B(n3961), .Z(n4065) );
  NAND U4224 ( .A(n4471), .B(n3963), .Z(n3965) );
  XOR U4225 ( .A(a[57]), .B(b[3]), .Z(n4040) );
  NAND U4226 ( .A(n33), .B(n4040), .Z(n3964) );
  NAND U4227 ( .A(n3965), .B(n3964), .Z(n4064) );
  XNOR U4228 ( .A(n4065), .B(n4064), .Z(n4066) );
  XOR U4229 ( .A(n4067), .B(n4066), .Z(n4044) );
  XOR U4230 ( .A(n4043), .B(n4044), .Z(n4046) );
  XOR U4231 ( .A(n4045), .B(n4046), .Z(n4017) );
  NANDN U4232 ( .A(n3967), .B(n3966), .Z(n3971) );
  OR U4233 ( .A(n3969), .B(n3968), .Z(n3970) );
  AND U4234 ( .A(n3971), .B(n3970), .Z(n4016) );
  XNOR U4235 ( .A(n4017), .B(n4016), .Z(n4019) );
  NAND U4236 ( .A(n4950), .B(n3972), .Z(n3974) );
  XOR U4237 ( .A(b[11]), .B(a[49]), .Z(n4049) );
  NAND U4238 ( .A(n4863), .B(n4049), .Z(n3973) );
  AND U4239 ( .A(n3974), .B(n3973), .Z(n4060) );
  NAND U4240 ( .A(n42), .B(n3975), .Z(n3977) );
  XOR U4241 ( .A(b[15]), .B(a[45]), .Z(n4052) );
  NAND U4242 ( .A(n4981), .B(n4052), .Z(n3976) );
  AND U4243 ( .A(n3977), .B(n3976), .Z(n4059) );
  NAND U4244 ( .A(n41), .B(n3978), .Z(n3980) );
  XOR U4245 ( .A(b[9]), .B(a[51]), .Z(n4055) );
  NAND U4246 ( .A(n4810), .B(n4055), .Z(n3979) );
  NAND U4247 ( .A(n3980), .B(n3979), .Z(n4058) );
  XOR U4248 ( .A(n4059), .B(n4058), .Z(n4061) );
  XOR U4249 ( .A(n4060), .B(n4061), .Z(n4071) );
  NANDN U4250 ( .A(n3982), .B(n3981), .Z(n3986) );
  OR U4251 ( .A(n3984), .B(n3983), .Z(n3985) );
  AND U4252 ( .A(n3986), .B(n3985), .Z(n4070) );
  XNOR U4253 ( .A(n4071), .B(n4070), .Z(n4072) );
  NANDN U4254 ( .A(n3988), .B(n3987), .Z(n3992) );
  NANDN U4255 ( .A(n3990), .B(n3989), .Z(n3991) );
  NAND U4256 ( .A(n3992), .B(n3991), .Z(n4073) );
  XNOR U4257 ( .A(n4072), .B(n4073), .Z(n4018) );
  XOR U4258 ( .A(n4019), .B(n4018), .Z(n4077) );
  NANDN U4259 ( .A(n3994), .B(n3993), .Z(n3998) );
  NANDN U4260 ( .A(n3996), .B(n3995), .Z(n3997) );
  AND U4261 ( .A(n3998), .B(n3997), .Z(n4076) );
  XNOR U4262 ( .A(n4077), .B(n4076), .Z(n4078) );
  XOR U4263 ( .A(n4079), .B(n4078), .Z(n4011) );
  NANDN U4264 ( .A(n4000), .B(n3999), .Z(n4004) );
  NAND U4265 ( .A(n4002), .B(n4001), .Z(n4003) );
  AND U4266 ( .A(n4004), .B(n4003), .Z(n4010) );
  XNOR U4267 ( .A(n4011), .B(n4010), .Z(n4012) );
  XNOR U4268 ( .A(n4013), .B(n4012), .Z(n4082) );
  XNOR U4269 ( .A(sreg[107]), .B(n4082), .Z(n4084) );
  NANDN U4270 ( .A(sreg[106]), .B(n4005), .Z(n4009) );
  NAND U4271 ( .A(n4007), .B(n4006), .Z(n4008) );
  NAND U4272 ( .A(n4009), .B(n4008), .Z(n4083) );
  XNOR U4273 ( .A(n4084), .B(n4083), .Z(c[107]) );
  NANDN U4274 ( .A(n4011), .B(n4010), .Z(n4015) );
  NANDN U4275 ( .A(n4013), .B(n4012), .Z(n4014) );
  AND U4276 ( .A(n4015), .B(n4014), .Z(n4090) );
  NANDN U4277 ( .A(n4017), .B(n4016), .Z(n4021) );
  NAND U4278 ( .A(n4019), .B(n4018), .Z(n4020) );
  AND U4279 ( .A(n4021), .B(n4020), .Z(n4152) );
  NANDN U4280 ( .A(n4023), .B(n4022), .Z(n4027) );
  NANDN U4281 ( .A(n4025), .B(n4024), .Z(n4026) );
  AND U4282 ( .A(n4027), .B(n4026), .Z(n4121) );
  NAND U4283 ( .A(n5012), .B(n4028), .Z(n4030) );
  XOR U4284 ( .A(b[13]), .B(a[48]), .Z(n4103) );
  NAND U4285 ( .A(n4985), .B(n4103), .Z(n4029) );
  AND U4286 ( .A(n4030), .B(n4029), .Z(n4098) );
  AND U4287 ( .A(b[15]), .B(a[44]), .Z(n4097) );
  XNOR U4288 ( .A(n4098), .B(n4097), .Z(n4099) );
  NAND U4289 ( .A(b[0]), .B(a[60]), .Z(n4031) );
  XNOR U4290 ( .A(b[1]), .B(n4031), .Z(n4033) );
  NANDN U4291 ( .A(b[0]), .B(a[59]), .Z(n4032) );
  NAND U4292 ( .A(n4033), .B(n4032), .Z(n4100) );
  XNOR U4293 ( .A(n4099), .B(n4100), .Z(n4119) );
  NAND U4294 ( .A(n36), .B(n4034), .Z(n4036) );
  XOR U4295 ( .A(a[56]), .B(b[5]), .Z(n4109) );
  NAND U4296 ( .A(n4560), .B(n4109), .Z(n4035) );
  NAND U4297 ( .A(n4036), .B(n4035), .Z(n4140) );
  NAND U4298 ( .A(n4755), .B(n4037), .Z(n4039) );
  XOR U4299 ( .A(b[7]), .B(a[54]), .Z(n4112) );
  NAND U4300 ( .A(n4708), .B(n4112), .Z(n4038) );
  NAND U4301 ( .A(n4039), .B(n4038), .Z(n4138) );
  NAND U4302 ( .A(n4471), .B(n4040), .Z(n4042) );
  XOR U4303 ( .A(a[58]), .B(b[3]), .Z(n4115) );
  NAND U4304 ( .A(n33), .B(n4115), .Z(n4041) );
  NAND U4305 ( .A(n4042), .B(n4041), .Z(n4137) );
  XNOR U4306 ( .A(n4119), .B(n4118), .Z(n4120) );
  XNOR U4307 ( .A(n4121), .B(n4120), .Z(n4093) );
  NANDN U4308 ( .A(n4044), .B(n4043), .Z(n4048) );
  OR U4309 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U4310 ( .A(n4048), .B(n4047), .Z(n4094) );
  XNOR U4311 ( .A(n4093), .B(n4094), .Z(n4096) );
  NAND U4312 ( .A(n4950), .B(n4049), .Z(n4051) );
  XOR U4313 ( .A(b[11]), .B(a[50]), .Z(n4122) );
  NAND U4314 ( .A(n4863), .B(n4122), .Z(n4050) );
  AND U4315 ( .A(n4051), .B(n4050), .Z(n4134) );
  NAND U4316 ( .A(n42), .B(n4052), .Z(n4054) );
  XOR U4317 ( .A(b[15]), .B(a[46]), .Z(n4125) );
  NAND U4318 ( .A(n4981), .B(n4125), .Z(n4053) );
  AND U4319 ( .A(n4054), .B(n4053), .Z(n4132) );
  NAND U4320 ( .A(n41), .B(n4055), .Z(n4057) );
  XOR U4321 ( .A(b[9]), .B(a[52]), .Z(n4128) );
  NAND U4322 ( .A(n4810), .B(n4128), .Z(n4056) );
  NAND U4323 ( .A(n4057), .B(n4056), .Z(n4131) );
  XNOR U4324 ( .A(n4132), .B(n4131), .Z(n4133) );
  XOR U4325 ( .A(n4134), .B(n4133), .Z(n4144) );
  NANDN U4326 ( .A(n4059), .B(n4058), .Z(n4063) );
  OR U4327 ( .A(n4061), .B(n4060), .Z(n4062) );
  AND U4328 ( .A(n4063), .B(n4062), .Z(n4143) );
  XOR U4329 ( .A(n4144), .B(n4143), .Z(n4145) );
  NANDN U4330 ( .A(n4065), .B(n4064), .Z(n4069) );
  NANDN U4331 ( .A(n4067), .B(n4066), .Z(n4068) );
  NAND U4332 ( .A(n4069), .B(n4068), .Z(n4146) );
  XNOR U4333 ( .A(n4145), .B(n4146), .Z(n4095) );
  XOR U4334 ( .A(n4096), .B(n4095), .Z(n4150) );
  NANDN U4335 ( .A(n4071), .B(n4070), .Z(n4075) );
  NANDN U4336 ( .A(n4073), .B(n4072), .Z(n4074) );
  AND U4337 ( .A(n4075), .B(n4074), .Z(n4149) );
  XNOR U4338 ( .A(n4150), .B(n4149), .Z(n4151) );
  XOR U4339 ( .A(n4152), .B(n4151), .Z(n4088) );
  NANDN U4340 ( .A(n4077), .B(n4076), .Z(n4081) );
  NAND U4341 ( .A(n4079), .B(n4078), .Z(n4080) );
  AND U4342 ( .A(n4081), .B(n4080), .Z(n4087) );
  XNOR U4343 ( .A(n4088), .B(n4087), .Z(n4089) );
  XNOR U4344 ( .A(n4090), .B(n4089), .Z(n4155) );
  XNOR U4345 ( .A(sreg[108]), .B(n4155), .Z(n4157) );
  NANDN U4346 ( .A(sreg[107]), .B(n4082), .Z(n4086) );
  NAND U4347 ( .A(n4084), .B(n4083), .Z(n4085) );
  NAND U4348 ( .A(n4086), .B(n4085), .Z(n4156) );
  XNOR U4349 ( .A(n4157), .B(n4156), .Z(c[108]) );
  NANDN U4350 ( .A(n4088), .B(n4087), .Z(n4092) );
  NANDN U4351 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U4352 ( .A(n4092), .B(n4091), .Z(n4163) );
  NANDN U4353 ( .A(n4098), .B(n4097), .Z(n4102) );
  NANDN U4354 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND U4355 ( .A(n4102), .B(n4101), .Z(n4217) );
  NAND U4356 ( .A(n5012), .B(n4103), .Z(n4105) );
  XOR U4357 ( .A(b[13]), .B(a[49]), .Z(n4199) );
  NAND U4358 ( .A(n4985), .B(n4199), .Z(n4104) );
  NAND U4359 ( .A(n4105), .B(n4104), .Z(n4194) );
  AND U4360 ( .A(b[15]), .B(a[45]), .Z(n4193) );
  NAND U4361 ( .A(b[0]), .B(a[61]), .Z(n4106) );
  XNOR U4362 ( .A(b[1]), .B(n4106), .Z(n4108) );
  NANDN U4363 ( .A(b[0]), .B(a[60]), .Z(n4107) );
  NAND U4364 ( .A(n4108), .B(n4107), .Z(n4196) );
  XNOR U4365 ( .A(n4195), .B(n4196), .Z(n4215) );
  NAND U4366 ( .A(n36), .B(n4109), .Z(n4111) );
  XOR U4367 ( .A(a[57]), .B(b[5]), .Z(n4205) );
  NAND U4368 ( .A(n4560), .B(n4205), .Z(n4110) );
  NAND U4369 ( .A(n4111), .B(n4110), .Z(n4190) );
  NAND U4370 ( .A(n4755), .B(n4112), .Z(n4114) );
  XOR U4371 ( .A(b[7]), .B(a[55]), .Z(n4208) );
  NAND U4372 ( .A(n4708), .B(n4208), .Z(n4113) );
  NAND U4373 ( .A(n4114), .B(n4113), .Z(n4188) );
  NAND U4374 ( .A(n4471), .B(n4115), .Z(n4117) );
  XOR U4375 ( .A(a[59]), .B(b[3]), .Z(n4211) );
  NAND U4376 ( .A(n33), .B(n4211), .Z(n4116) );
  NAND U4377 ( .A(n4117), .B(n4116), .Z(n4187) );
  XOR U4378 ( .A(n4215), .B(n4214), .Z(n4216) );
  XOR U4379 ( .A(n4166), .B(n4167), .Z(n4169) );
  NAND U4380 ( .A(n4950), .B(n4122), .Z(n4124) );
  XOR U4381 ( .A(b[11]), .B(a[51]), .Z(n4172) );
  NAND U4382 ( .A(n4863), .B(n4172), .Z(n4123) );
  NAND U4383 ( .A(n4124), .B(n4123), .Z(n4184) );
  NAND U4384 ( .A(n42), .B(n4125), .Z(n4127) );
  XOR U4385 ( .A(b[15]), .B(a[47]), .Z(n4175) );
  NAND U4386 ( .A(n4981), .B(n4175), .Z(n4126) );
  NAND U4387 ( .A(n4127), .B(n4126), .Z(n4182) );
  NAND U4388 ( .A(n41), .B(n4128), .Z(n4130) );
  XOR U4389 ( .A(b[9]), .B(a[53]), .Z(n4178) );
  NAND U4390 ( .A(n4810), .B(n4178), .Z(n4129) );
  NAND U4391 ( .A(n4130), .B(n4129), .Z(n4181) );
  NANDN U4392 ( .A(n4132), .B(n4131), .Z(n4136) );
  NANDN U4393 ( .A(n4134), .B(n4133), .Z(n4135) );
  AND U4394 ( .A(n4136), .B(n4135), .Z(n4221) );
  XOR U4395 ( .A(n4220), .B(n4221), .Z(n4222) );
  NAND U4396 ( .A(n4138), .B(n4137), .Z(n4142) );
  NAND U4397 ( .A(n4140), .B(n4139), .Z(n4141) );
  AND U4398 ( .A(n4142), .B(n4141), .Z(n4223) );
  XOR U4399 ( .A(n4169), .B(n4168), .Z(n4227) );
  NAND U4400 ( .A(n4144), .B(n4143), .Z(n4148) );
  NANDN U4401 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U4402 ( .A(n4148), .B(n4147), .Z(n4226) );
  XNOR U4403 ( .A(n4227), .B(n4226), .Z(n4228) );
  XOR U4404 ( .A(n4229), .B(n4228), .Z(n4161) );
  NANDN U4405 ( .A(n4150), .B(n4149), .Z(n4154) );
  NAND U4406 ( .A(n4152), .B(n4151), .Z(n4153) );
  AND U4407 ( .A(n4154), .B(n4153), .Z(n4160) );
  XNOR U4408 ( .A(n4161), .B(n4160), .Z(n4162) );
  XNOR U4409 ( .A(n4163), .B(n4162), .Z(n4232) );
  XNOR U4410 ( .A(sreg[109]), .B(n4232), .Z(n4234) );
  NANDN U4411 ( .A(sreg[108]), .B(n4155), .Z(n4159) );
  NAND U4412 ( .A(n4157), .B(n4156), .Z(n4158) );
  NAND U4413 ( .A(n4159), .B(n4158), .Z(n4233) );
  XNOR U4414 ( .A(n4234), .B(n4233), .Z(c[109]) );
  NANDN U4415 ( .A(n4161), .B(n4160), .Z(n4165) );
  NANDN U4416 ( .A(n4163), .B(n4162), .Z(n4164) );
  AND U4417 ( .A(n4165), .B(n4164), .Z(n4240) );
  NAND U4418 ( .A(n4167), .B(n4166), .Z(n4171) );
  NAND U4419 ( .A(n4169), .B(n4168), .Z(n4170) );
  AND U4420 ( .A(n4171), .B(n4170), .Z(n4306) );
  NAND U4421 ( .A(n4950), .B(n4172), .Z(n4174) );
  XOR U4422 ( .A(b[11]), .B(a[52]), .Z(n4276) );
  NAND U4423 ( .A(n4863), .B(n4276), .Z(n4173) );
  NAND U4424 ( .A(n4174), .B(n4173), .Z(n4288) );
  NAND U4425 ( .A(n42), .B(n4175), .Z(n4177) );
  XOR U4426 ( .A(b[15]), .B(a[48]), .Z(n4279) );
  NAND U4427 ( .A(n4981), .B(n4279), .Z(n4176) );
  NAND U4428 ( .A(n4177), .B(n4176), .Z(n4286) );
  NAND U4429 ( .A(n41), .B(n4178), .Z(n4180) );
  XOR U4430 ( .A(b[9]), .B(a[54]), .Z(n4282) );
  NAND U4431 ( .A(n4810), .B(n4282), .Z(n4179) );
  NAND U4432 ( .A(n4180), .B(n4179), .Z(n4285) );
  NAND U4433 ( .A(n4182), .B(n4181), .Z(n4186) );
  NAND U4434 ( .A(n4184), .B(n4183), .Z(n4185) );
  AND U4435 ( .A(n4186), .B(n4185), .Z(n4298) );
  XOR U4436 ( .A(n4297), .B(n4298), .Z(n4299) );
  NAND U4437 ( .A(n4188), .B(n4187), .Z(n4192) );
  NAND U4438 ( .A(n4190), .B(n4189), .Z(n4191) );
  AND U4439 ( .A(n4192), .B(n4191), .Z(n4300) );
  NAND U4440 ( .A(n4194), .B(n4193), .Z(n4198) );
  NANDN U4441 ( .A(n4196), .B(n4195), .Z(n4197) );
  NAND U4442 ( .A(n4198), .B(n4197), .Z(n4273) );
  NAND U4443 ( .A(n5012), .B(n4199), .Z(n4201) );
  XOR U4444 ( .A(b[13]), .B(a[50]), .Z(n4255) );
  NAND U4445 ( .A(n4985), .B(n4255), .Z(n4200) );
  NAND U4446 ( .A(n4201), .B(n4200), .Z(n4250) );
  AND U4447 ( .A(b[15]), .B(a[46]), .Z(n4249) );
  NAND U4448 ( .A(b[0]), .B(a[62]), .Z(n4202) );
  XNOR U4449 ( .A(b[1]), .B(n4202), .Z(n4204) );
  NANDN U4450 ( .A(b[0]), .B(a[61]), .Z(n4203) );
  NAND U4451 ( .A(n4204), .B(n4203), .Z(n4252) );
  XNOR U4452 ( .A(n4251), .B(n4252), .Z(n4271) );
  NAND U4453 ( .A(n36), .B(n4205), .Z(n4207) );
  XOR U4454 ( .A(a[58]), .B(b[5]), .Z(n4261) );
  NAND U4455 ( .A(n4560), .B(n4261), .Z(n4206) );
  NAND U4456 ( .A(n4207), .B(n4206), .Z(n4294) );
  NAND U4457 ( .A(n4755), .B(n4208), .Z(n4210) );
  XOR U4458 ( .A(b[7]), .B(a[56]), .Z(n4264) );
  NAND U4459 ( .A(n4708), .B(n4264), .Z(n4209) );
  NAND U4460 ( .A(n4210), .B(n4209), .Z(n4292) );
  NAND U4461 ( .A(n4471), .B(n4211), .Z(n4213) );
  XOR U4462 ( .A(a[60]), .B(b[3]), .Z(n4267) );
  NAND U4463 ( .A(n33), .B(n4267), .Z(n4212) );
  NAND U4464 ( .A(n4213), .B(n4212), .Z(n4291) );
  XOR U4465 ( .A(n4271), .B(n4270), .Z(n4272) );
  NAND U4466 ( .A(n4215), .B(n4214), .Z(n4219) );
  NAND U4467 ( .A(n4217), .B(n4216), .Z(n4218) );
  AND U4468 ( .A(n4219), .B(n4218), .Z(n4244) );
  XOR U4469 ( .A(n4243), .B(n4244), .Z(n4245) );
  XNOR U4470 ( .A(n4246), .B(n4245), .Z(n4304) );
  NAND U4471 ( .A(n4221), .B(n4220), .Z(n4225) );
  NAND U4472 ( .A(n4223), .B(n4222), .Z(n4224) );
  AND U4473 ( .A(n4225), .B(n4224), .Z(n4303) );
  XOR U4474 ( .A(n4306), .B(n4305), .Z(n4238) );
  NANDN U4475 ( .A(n4227), .B(n4226), .Z(n4231) );
  NAND U4476 ( .A(n4229), .B(n4228), .Z(n4230) );
  AND U4477 ( .A(n4231), .B(n4230), .Z(n4237) );
  XNOR U4478 ( .A(n4238), .B(n4237), .Z(n4239) );
  XNOR U4479 ( .A(n4240), .B(n4239), .Z(n4309) );
  XNOR U4480 ( .A(sreg[110]), .B(n4309), .Z(n4311) );
  NANDN U4481 ( .A(sreg[109]), .B(n4232), .Z(n4236) );
  NAND U4482 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U4483 ( .A(n4236), .B(n4235), .Z(n4310) );
  XNOR U4484 ( .A(n4311), .B(n4310), .Z(c[110]) );
  NANDN U4485 ( .A(n4238), .B(n4237), .Z(n4242) );
  NANDN U4486 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U4487 ( .A(n4242), .B(n4241), .Z(n4322) );
  NAND U4488 ( .A(n4244), .B(n4243), .Z(n4248) );
  NAND U4489 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U4490 ( .A(n4248), .B(n4247), .Z(n4385) );
  NAND U4491 ( .A(n4250), .B(n4249), .Z(n4254) );
  NANDN U4492 ( .A(n4252), .B(n4251), .Z(n4253) );
  NAND U4493 ( .A(n4254), .B(n4253), .Z(n4373) );
  NAND U4494 ( .A(n5012), .B(n4255), .Z(n4257) );
  XOR U4495 ( .A(b[13]), .B(a[51]), .Z(n4358) );
  NAND U4496 ( .A(n4985), .B(n4358), .Z(n4256) );
  NAND U4497 ( .A(n4257), .B(n4256), .Z(n4353) );
  AND U4498 ( .A(b[15]), .B(a[47]), .Z(n4352) );
  NAND U4499 ( .A(b[0]), .B(a[63]), .Z(n4258) );
  XNOR U4500 ( .A(b[1]), .B(n4258), .Z(n4260) );
  NANDN U4501 ( .A(b[0]), .B(a[62]), .Z(n4259) );
  NAND U4502 ( .A(n4260), .B(n4259), .Z(n4355) );
  XNOR U4503 ( .A(n4354), .B(n4355), .Z(n4371) );
  NAND U4504 ( .A(n36), .B(n4261), .Z(n4263) );
  XOR U4505 ( .A(a[59]), .B(b[5]), .Z(n4361) );
  NAND U4506 ( .A(n4560), .B(n4361), .Z(n4262) );
  NAND U4507 ( .A(n4263), .B(n4262), .Z(n4349) );
  NAND U4508 ( .A(n4755), .B(n4264), .Z(n4266) );
  XOR U4509 ( .A(a[57]), .B(b[7]), .Z(n4364) );
  NAND U4510 ( .A(n4708), .B(n4364), .Z(n4265) );
  NAND U4511 ( .A(n4266), .B(n4265), .Z(n4347) );
  NAND U4512 ( .A(n4471), .B(n4267), .Z(n4269) );
  XOR U4513 ( .A(a[61]), .B(b[3]), .Z(n4367) );
  NAND U4514 ( .A(n33), .B(n4367), .Z(n4268) );
  NAND U4515 ( .A(n4269), .B(n4268), .Z(n4346) );
  XOR U4516 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U4517 ( .A(n4271), .B(n4270), .Z(n4275) );
  NAND U4518 ( .A(n4273), .B(n4272), .Z(n4274) );
  AND U4519 ( .A(n4275), .B(n4274), .Z(n4326) );
  XOR U4520 ( .A(n4325), .B(n4326), .Z(n4328) );
  NAND U4521 ( .A(n4950), .B(n4276), .Z(n4278) );
  XOR U4522 ( .A(b[11]), .B(a[53]), .Z(n4331) );
  NAND U4523 ( .A(n4863), .B(n4331), .Z(n4277) );
  NAND U4524 ( .A(n4278), .B(n4277), .Z(n4343) );
  NAND U4525 ( .A(n42), .B(n4279), .Z(n4281) );
  XOR U4526 ( .A(b[15]), .B(a[49]), .Z(n4334) );
  NAND U4527 ( .A(n4981), .B(n4334), .Z(n4280) );
  NAND U4528 ( .A(n4281), .B(n4280), .Z(n4341) );
  NAND U4529 ( .A(n41), .B(n4282), .Z(n4284) );
  XOR U4530 ( .A(b[9]), .B(a[55]), .Z(n4337) );
  NAND U4531 ( .A(n4810), .B(n4337), .Z(n4283) );
  NAND U4532 ( .A(n4284), .B(n4283), .Z(n4340) );
  NAND U4533 ( .A(n4286), .B(n4285), .Z(n4290) );
  NAND U4534 ( .A(n4288), .B(n4287), .Z(n4289) );
  AND U4535 ( .A(n4290), .B(n4289), .Z(n4377) );
  XOR U4536 ( .A(n4376), .B(n4377), .Z(n4378) );
  NAND U4537 ( .A(n4292), .B(n4291), .Z(n4296) );
  NAND U4538 ( .A(n4294), .B(n4293), .Z(n4295) );
  AND U4539 ( .A(n4296), .B(n4295), .Z(n4379) );
  XNOR U4540 ( .A(n4328), .B(n4327), .Z(n4383) );
  NAND U4541 ( .A(n4298), .B(n4297), .Z(n4302) );
  NAND U4542 ( .A(n4300), .B(n4299), .Z(n4301) );
  AND U4543 ( .A(n4302), .B(n4301), .Z(n4382) );
  XNOR U4544 ( .A(n4385), .B(n4384), .Z(n4320) );
  NAND U4545 ( .A(n4304), .B(n4303), .Z(n4308) );
  NAND U4546 ( .A(n4306), .B(n4305), .Z(n4307) );
  AND U4547 ( .A(n4308), .B(n4307), .Z(n4319) );
  XNOR U4548 ( .A(sreg[111]), .B(n4314), .Z(n4316) );
  NANDN U4549 ( .A(sreg[110]), .B(n4309), .Z(n4313) );
  NAND U4550 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND U4551 ( .A(n4313), .B(n4312), .Z(n4315) );
  XNOR U4552 ( .A(n4316), .B(n4315), .Z(c[111]) );
  NANDN U4553 ( .A(sreg[111]), .B(n4314), .Z(n4318) );
  NAND U4554 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U4555 ( .A(n4318), .B(n4317), .Z(n4389) );
  NAND U4556 ( .A(n4320), .B(n4319), .Z(n4324) );
  NAND U4557 ( .A(n4322), .B(n4321), .Z(n4323) );
  AND U4558 ( .A(n4324), .B(n4323), .Z(n4393) );
  NAND U4559 ( .A(n4326), .B(n4325), .Z(n4330) );
  NAND U4560 ( .A(n4328), .B(n4327), .Z(n4329) );
  AND U4561 ( .A(n4330), .B(n4329), .Z(n4454) );
  NAND U4562 ( .A(n4950), .B(n4331), .Z(n4333) );
  XOR U4563 ( .A(b[11]), .B(a[54]), .Z(n4405) );
  NAND U4564 ( .A(n4863), .B(n4405), .Z(n4332) );
  NAND U4565 ( .A(n4333), .B(n4332), .Z(n4414) );
  NAND U4566 ( .A(n42), .B(n4334), .Z(n4336) );
  XOR U4567 ( .A(b[15]), .B(a[50]), .Z(n4429) );
  NAND U4568 ( .A(n4981), .B(n4429), .Z(n4335) );
  NAND U4569 ( .A(n4336), .B(n4335), .Z(n4412) );
  NAND U4570 ( .A(n41), .B(n4337), .Z(n4339) );
  XOR U4571 ( .A(b[9]), .B(a[56]), .Z(n4402) );
  NAND U4572 ( .A(n4810), .B(n4402), .Z(n4338) );
  NAND U4573 ( .A(n4339), .B(n4338), .Z(n4411) );
  NAND U4574 ( .A(n4341), .B(n4340), .Z(n4345) );
  NAND U4575 ( .A(n4343), .B(n4342), .Z(n4344) );
  AND U4576 ( .A(n4345), .B(n4344), .Z(n4446) );
  XOR U4577 ( .A(n4445), .B(n4446), .Z(n4447) );
  NAND U4578 ( .A(n4347), .B(n4346), .Z(n4351) );
  NAND U4579 ( .A(n4349), .B(n4348), .Z(n4350) );
  AND U4580 ( .A(n4351), .B(n4350), .Z(n4448) );
  NAND U4581 ( .A(n4353), .B(n4352), .Z(n4357) );
  NANDN U4582 ( .A(n4355), .B(n4354), .Z(n4356) );
  NAND U4583 ( .A(n4357), .B(n4356), .Z(n4442) );
  NAND U4584 ( .A(n5012), .B(n4358), .Z(n4360) );
  XOR U4585 ( .A(b[13]), .B(a[52]), .Z(n4432) );
  NAND U4586 ( .A(n4985), .B(n4432), .Z(n4359) );
  NAND U4587 ( .A(n4360), .B(n4359), .Z(n4426) );
  AND U4588 ( .A(b[15]), .B(a[48]), .Z(n4423) );
  NAND U4589 ( .A(n36), .B(n4361), .Z(n4363) );
  XOR U4590 ( .A(a[60]), .B(b[5]), .Z(n4436) );
  NAND U4591 ( .A(n4560), .B(n4436), .Z(n4362) );
  NAND U4592 ( .A(n4363), .B(n4362), .Z(n4420) );
  NAND U4593 ( .A(n4755), .B(n4364), .Z(n4366) );
  XOR U4594 ( .A(a[58]), .B(b[7]), .Z(n4408) );
  NAND U4595 ( .A(n4708), .B(n4408), .Z(n4365) );
  NAND U4596 ( .A(n4366), .B(n4365), .Z(n4418) );
  NAND U4597 ( .A(n4471), .B(n4367), .Z(n4369) );
  XOR U4598 ( .A(a[62]), .B(b[3]), .Z(n4435) );
  NAND U4599 ( .A(n33), .B(n4435), .Z(n4368) );
  NAND U4600 ( .A(n4369), .B(n4368), .Z(n4417) );
  XOR U4601 ( .A(n4440), .B(n4439), .Z(n4441) );
  NAND U4602 ( .A(n4371), .B(n4370), .Z(n4375) );
  NAND U4603 ( .A(n4373), .B(n4372), .Z(n4374) );
  AND U4604 ( .A(n4375), .B(n4374), .Z(n4397) );
  XOR U4605 ( .A(n4396), .B(n4397), .Z(n4398) );
  XNOR U4606 ( .A(n4399), .B(n4398), .Z(n4452) );
  NAND U4607 ( .A(n4377), .B(n4376), .Z(n4381) );
  NAND U4608 ( .A(n4379), .B(n4378), .Z(n4380) );
  AND U4609 ( .A(n4381), .B(n4380), .Z(n4451) );
  XNOR U4610 ( .A(n4454), .B(n4453), .Z(n4391) );
  NAND U4611 ( .A(n4383), .B(n4382), .Z(n4387) );
  NAND U4612 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U4613 ( .A(n4387), .B(n4386), .Z(n4390) );
  XOR U4614 ( .A(n4393), .B(n4392), .Z(n4388) );
  XOR U4615 ( .A(n4389), .B(n4388), .Z(c[112]) );
  AND U4616 ( .A(n4389), .B(n4388), .Z(n4458) );
  NAND U4617 ( .A(n4391), .B(n4390), .Z(n4395) );
  NANDN U4618 ( .A(n4393), .B(n4392), .Z(n4394) );
  AND U4619 ( .A(n4395), .B(n4394), .Z(n4462) );
  NAND U4620 ( .A(n4397), .B(n4396), .Z(n4401) );
  NAND U4621 ( .A(n4399), .B(n4398), .Z(n4400) );
  AND U4622 ( .A(n4401), .B(n4400), .Z(n4524) );
  NAND U4623 ( .A(n41), .B(n4402), .Z(n4404) );
  XOR U4624 ( .A(b[9]), .B(a[57]), .Z(n4490) );
  NAND U4625 ( .A(n4810), .B(n4490), .Z(n4403) );
  NAND U4626 ( .A(n4404), .B(n4403), .Z(n4496) );
  NAND U4627 ( .A(n4950), .B(n4405), .Z(n4407) );
  XOR U4628 ( .A(b[11]), .B(a[55]), .Z(n4478) );
  NAND U4629 ( .A(n4863), .B(n4478), .Z(n4406) );
  NAND U4630 ( .A(n4407), .B(n4406), .Z(n4494) );
  NAND U4631 ( .A(n4755), .B(n4408), .Z(n4410) );
  XOR U4632 ( .A(a[59]), .B(b[7]), .Z(n4484) );
  NAND U4633 ( .A(n4708), .B(n4484), .Z(n4409) );
  NAND U4634 ( .A(n4410), .B(n4409), .Z(n4493) );
  NAND U4635 ( .A(n4412), .B(n4411), .Z(n4416) );
  NAND U4636 ( .A(n4414), .B(n4413), .Z(n4415) );
  AND U4637 ( .A(n4416), .B(n4415), .Z(n4516) );
  XOR U4638 ( .A(n4515), .B(n4516), .Z(n4517) );
  NAND U4639 ( .A(n4418), .B(n4417), .Z(n4422) );
  NAND U4640 ( .A(n4420), .B(n4419), .Z(n4421) );
  AND U4641 ( .A(n4422), .B(n4421), .Z(n4518) );
  NAND U4642 ( .A(n4424), .B(n4423), .Z(n4428) );
  NAND U4643 ( .A(n4426), .B(n4425), .Z(n4427) );
  NAND U4644 ( .A(n4428), .B(n4427), .Z(n4512) );
  NAND U4645 ( .A(n42), .B(n4429), .Z(n4431) );
  XOR U4646 ( .A(b[15]), .B(a[51]), .Z(n4475) );
  NAND U4647 ( .A(n4981), .B(n4475), .Z(n4430) );
  NAND U4648 ( .A(n4431), .B(n4430), .Z(n4506) );
  AND U4649 ( .A(b[15]), .B(a[49]), .Z(n4624) );
  NAND U4650 ( .A(n5012), .B(n4432), .Z(n4434) );
  XOR U4651 ( .A(b[13]), .B(a[53]), .Z(n4481) );
  NAND U4652 ( .A(n4985), .B(n4481), .Z(n4433) );
  NAND U4653 ( .A(n4434), .B(n4433), .Z(n4504) );
  XNOR U4654 ( .A(n4624), .B(n4504), .Z(n4505) );
  XNOR U4655 ( .A(a[63]), .B(b[3]), .Z(n4472) );
  NAND U4656 ( .A(n36), .B(n4436), .Z(n4438) );
  XOR U4657 ( .A(a[61]), .B(b[5]), .Z(n4487) );
  NAND U4658 ( .A(n4560), .B(n4487), .Z(n4437) );
  NAND U4659 ( .A(n4438), .B(n4437), .Z(n4499) );
  XNOR U4660 ( .A(b[1]), .B(n4499), .Z(n4500) );
  XOR U4661 ( .A(n4510), .B(n4509), .Z(n4511) );
  NAND U4662 ( .A(n4440), .B(n4439), .Z(n4444) );
  NAND U4663 ( .A(n4442), .B(n4441), .Z(n4443) );
  AND U4664 ( .A(n4444), .B(n4443), .Z(n4466) );
  XOR U4665 ( .A(n4465), .B(n4466), .Z(n4467) );
  XNOR U4666 ( .A(n4468), .B(n4467), .Z(n4522) );
  NAND U4667 ( .A(n4446), .B(n4445), .Z(n4450) );
  NAND U4668 ( .A(n4448), .B(n4447), .Z(n4449) );
  AND U4669 ( .A(n4450), .B(n4449), .Z(n4521) );
  XNOR U4670 ( .A(n4524), .B(n4523), .Z(n4460) );
  NAND U4671 ( .A(n4452), .B(n4451), .Z(n4456) );
  NAND U4672 ( .A(n4454), .B(n4453), .Z(n4455) );
  AND U4673 ( .A(n4456), .B(n4455), .Z(n4459) );
  XOR U4674 ( .A(n4462), .B(n4461), .Z(n4457) );
  XOR U4675 ( .A(n4458), .B(n4457), .Z(c[113]) );
  AND U4676 ( .A(n4458), .B(n4457), .Z(n4528) );
  NAND U4677 ( .A(n4460), .B(n4459), .Z(n4464) );
  NANDN U4678 ( .A(n4462), .B(n4461), .Z(n4463) );
  AND U4679 ( .A(n4464), .B(n4463), .Z(n4532) );
  NAND U4680 ( .A(n4466), .B(n4465), .Z(n4470) );
  NAND U4681 ( .A(n4468), .B(n4467), .Z(n4469) );
  AND U4682 ( .A(n4470), .B(n4469), .Z(n4592) );
  NANDN U4683 ( .A(n4472), .B(n4471), .Z(n4473) );
  AND U4684 ( .A(n4474), .B(n4473), .Z(n4572) );
  AND U4685 ( .A(b[15]), .B(a[50]), .Z(n4571) );
  XNOR U4686 ( .A(n4572), .B(n4571), .Z(n4573) );
  XNOR U4687 ( .A(n4624), .B(n4573), .Z(n4580) );
  NAND U4688 ( .A(n42), .B(n4475), .Z(n4477) );
  XOR U4689 ( .A(b[15]), .B(a[52]), .Z(n4547) );
  NAND U4690 ( .A(n4981), .B(n4547), .Z(n4476) );
  NAND U4691 ( .A(n4477), .B(n4476), .Z(n4578) );
  NAND U4692 ( .A(n4950), .B(n4478), .Z(n4480) );
  XOR U4693 ( .A(b[11]), .B(a[56]), .Z(n4561) );
  NAND U4694 ( .A(n4863), .B(n4561), .Z(n4479) );
  NAND U4695 ( .A(n4480), .B(n4479), .Z(n4577) );
  XOR U4696 ( .A(n4580), .B(n4579), .Z(n4544) );
  NAND U4697 ( .A(n5012), .B(n4481), .Z(n4483) );
  XOR U4698 ( .A(b[13]), .B(a[54]), .Z(n4556) );
  NAND U4699 ( .A(n4985), .B(n4556), .Z(n4482) );
  NAND U4700 ( .A(n4483), .B(n4482), .Z(n4542) );
  NAND U4701 ( .A(n4755), .B(n4484), .Z(n4486) );
  XOR U4702 ( .A(a[60]), .B(b[7]), .Z(n4553) );
  NAND U4703 ( .A(n4708), .B(n4553), .Z(n4485) );
  NAND U4704 ( .A(n4486), .B(n4485), .Z(n4568) );
  NAND U4705 ( .A(n36), .B(n4487), .Z(n4489) );
  XOR U4706 ( .A(a[62]), .B(b[5]), .Z(n4559) );
  NAND U4707 ( .A(n4560), .B(n4559), .Z(n4488) );
  NAND U4708 ( .A(n4489), .B(n4488), .Z(n4566) );
  NAND U4709 ( .A(n41), .B(n4490), .Z(n4492) );
  XOR U4710 ( .A(b[9]), .B(a[58]), .Z(n4550) );
  NAND U4711 ( .A(n4810), .B(n4550), .Z(n4491) );
  NAND U4712 ( .A(n4492), .B(n4491), .Z(n4565) );
  XOR U4713 ( .A(n4544), .B(n4543), .Z(n4586) );
  NAND U4714 ( .A(n4494), .B(n4493), .Z(n4498) );
  NAND U4715 ( .A(n4496), .B(n4495), .Z(n4497) );
  NAND U4716 ( .A(n4498), .B(n4497), .Z(n4584) );
  NANDN U4717 ( .A(b[1]), .B(n4499), .Z(n4503) );
  NAND U4718 ( .A(n4501), .B(n4500), .Z(n4502) );
  NAND U4719 ( .A(n4503), .B(n4502), .Z(n4583) );
  XNOR U4720 ( .A(n4586), .B(n4585), .Z(n4538) );
  IV U4721 ( .A(n4624), .Z(n4574) );
  NAND U4722 ( .A(n4574), .B(n4504), .Z(n4508) );
  NAND U4723 ( .A(n4506), .B(n4505), .Z(n4507) );
  AND U4724 ( .A(n4508), .B(n4507), .Z(n4535) );
  NAND U4725 ( .A(n4510), .B(n4509), .Z(n4514) );
  NAND U4726 ( .A(n4512), .B(n4511), .Z(n4513) );
  AND U4727 ( .A(n4514), .B(n4513), .Z(n4536) );
  NAND U4728 ( .A(n4516), .B(n4515), .Z(n4520) );
  NAND U4729 ( .A(n4518), .B(n4517), .Z(n4519) );
  AND U4730 ( .A(n4520), .B(n4519), .Z(n4590) );
  XOR U4731 ( .A(n4589), .B(n4590), .Z(n4591) );
  XNOR U4732 ( .A(n4592), .B(n4591), .Z(n4530) );
  NAND U4733 ( .A(n4522), .B(n4521), .Z(n4526) );
  NAND U4734 ( .A(n4524), .B(n4523), .Z(n4525) );
  AND U4735 ( .A(n4526), .B(n4525), .Z(n4529) );
  XOR U4736 ( .A(n4532), .B(n4531), .Z(n4527) );
  XOR U4737 ( .A(n4528), .B(n4527), .Z(c[114]) );
  AND U4738 ( .A(n4528), .B(n4527), .Z(n4596) );
  NAND U4739 ( .A(n4530), .B(n4529), .Z(n4534) );
  NANDN U4740 ( .A(n4532), .B(n4531), .Z(n4533) );
  AND U4741 ( .A(n4534), .B(n4533), .Z(n4600) );
  NAND U4742 ( .A(n4536), .B(n4535), .Z(n4540) );
  NAND U4743 ( .A(n4538), .B(n4537), .Z(n4539) );
  NAND U4744 ( .A(n4540), .B(n4539), .Z(n4606) );
  NAND U4745 ( .A(n4542), .B(n4541), .Z(n4546) );
  NAND U4746 ( .A(n4544), .B(n4543), .Z(n4545) );
  NAND U4747 ( .A(n4546), .B(n4545), .Z(n4610) );
  NAND U4748 ( .A(n42), .B(n4547), .Z(n4549) );
  XOR U4749 ( .A(b[15]), .B(a[53]), .Z(n4633) );
  NAND U4750 ( .A(n4981), .B(n4633), .Z(n4548) );
  NAND U4751 ( .A(n4549), .B(n4548), .Z(n4650) );
  NAND U4752 ( .A(n41), .B(n4550), .Z(n4552) );
  XOR U4753 ( .A(a[59]), .B(b[9]), .Z(n4639) );
  NAND U4754 ( .A(n4810), .B(n4639), .Z(n4551) );
  NAND U4755 ( .A(n4552), .B(n4551), .Z(n4618) );
  NAND U4756 ( .A(n4755), .B(n4553), .Z(n4555) );
  XOR U4757 ( .A(a[61]), .B(b[7]), .Z(n4642) );
  NAND U4758 ( .A(n4708), .B(n4642), .Z(n4554) );
  NAND U4759 ( .A(n4555), .B(n4554), .Z(n4616) );
  NAND U4760 ( .A(n5012), .B(n4556), .Z(n4558) );
  XOR U4761 ( .A(b[13]), .B(a[55]), .Z(n4648) );
  NAND U4762 ( .A(n4985), .B(n4648), .Z(n4557) );
  NAND U4763 ( .A(n4558), .B(n4557), .Z(n4615) );
  XNOR U4764 ( .A(a[63]), .B(b[5]), .Z(n4636) );
  NAND U4765 ( .A(n4950), .B(n4561), .Z(n4563) );
  XOR U4766 ( .A(b[11]), .B(a[57]), .Z(n4645) );
  NAND U4767 ( .A(n4863), .B(n4645), .Z(n4562) );
  NAND U4768 ( .A(n4563), .B(n4562), .Z(n4627) );
  AND U4769 ( .A(b[15]), .B(a[51]), .Z(n4621) );
  XNOR U4770 ( .A(n4621), .B(n4564), .Z(n4623) );
  XOR U4771 ( .A(n4624), .B(n4623), .Z(n4629) );
  XOR U4772 ( .A(n4630), .B(n4629), .Z(n4651) );
  XOR U4773 ( .A(n4652), .B(n4651), .Z(n4609) );
  NAND U4774 ( .A(n4566), .B(n4565), .Z(n4570) );
  NAND U4775 ( .A(n4568), .B(n4567), .Z(n4569) );
  NAND U4776 ( .A(n4570), .B(n4569), .Z(n4658) );
  NANDN U4777 ( .A(n4572), .B(n4571), .Z(n4576) );
  NAND U4778 ( .A(n4574), .B(n4573), .Z(n4575) );
  NAND U4779 ( .A(n4576), .B(n4575), .Z(n4656) );
  NAND U4780 ( .A(n4578), .B(n4577), .Z(n4582) );
  NAND U4781 ( .A(n4580), .B(n4579), .Z(n4581) );
  NAND U4782 ( .A(n4582), .B(n4581), .Z(n4655) );
  XNOR U4783 ( .A(n4612), .B(n4611), .Z(n4604) );
  NAND U4784 ( .A(n4584), .B(n4583), .Z(n4588) );
  NAND U4785 ( .A(n4586), .B(n4585), .Z(n4587) );
  AND U4786 ( .A(n4588), .B(n4587), .Z(n4603) );
  NAND U4787 ( .A(n4590), .B(n4589), .Z(n4594) );
  NAND U4788 ( .A(n4592), .B(n4591), .Z(n4593) );
  AND U4789 ( .A(n4594), .B(n4593), .Z(n4598) );
  XOR U4790 ( .A(n4600), .B(n4599), .Z(n4595) );
  XOR U4791 ( .A(n4596), .B(n4595), .Z(c[115]) );
  AND U4792 ( .A(n4596), .B(n4595), .Z(n4662) );
  NAND U4793 ( .A(n4598), .B(n4597), .Z(n4602) );
  NANDN U4794 ( .A(n4600), .B(n4599), .Z(n4601) );
  AND U4795 ( .A(n4602), .B(n4601), .Z(n4666) );
  NAND U4796 ( .A(n4604), .B(n4603), .Z(n4608) );
  NAND U4797 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U4798 ( .A(n4608), .B(n4607), .Z(n4664) );
  NAND U4799 ( .A(n4610), .B(n4609), .Z(n4614) );
  NAND U4800 ( .A(n4612), .B(n4611), .Z(n4613) );
  AND U4801 ( .A(n4614), .B(n4613), .Z(n4672) );
  NAND U4802 ( .A(n4616), .B(n4615), .Z(n4620) );
  NAND U4803 ( .A(n4618), .B(n4617), .Z(n4619) );
  AND U4804 ( .A(n4620), .B(n4619), .Z(n4716) );
  NAND U4805 ( .A(n4622), .B(n4621), .Z(n4626) );
  NAND U4806 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U4807 ( .A(n4626), .B(n4625), .Z(n4713) );
  NAND U4808 ( .A(n4628), .B(n4627), .Z(n4632) );
  NAND U4809 ( .A(n4630), .B(n4629), .Z(n4631) );
  AND U4810 ( .A(n4632), .B(n4631), .Z(n4714) );
  XNOR U4811 ( .A(n4716), .B(n4715), .Z(n4678) );
  NAND U4812 ( .A(n42), .B(n4633), .Z(n4635) );
  XOR U4813 ( .A(b[15]), .B(a[54]), .Z(n4704) );
  NAND U4814 ( .A(n4981), .B(n4704), .Z(n4634) );
  NAND U4815 ( .A(n4635), .B(n4634), .Z(n4689) );
  NANDN U4816 ( .A(n4636), .B(n36), .Z(n4637) );
  AND U4817 ( .A(n4638), .B(n4637), .Z(n4687) );
  AND U4818 ( .A(b[15]), .B(a[52]), .Z(n4712) );
  IV U4819 ( .A(n4712), .Z(n4765) );
  XNOR U4820 ( .A(n4687), .B(n4765), .Z(n4688) );
  NAND U4821 ( .A(n41), .B(n4639), .Z(n4641) );
  XOR U4822 ( .A(a[60]), .B(b[9]), .Z(n4698) );
  NAND U4823 ( .A(n4810), .B(n4698), .Z(n4640) );
  NAND U4824 ( .A(n4641), .B(n4640), .Z(n4695) );
  NAND U4825 ( .A(n4755), .B(n4642), .Z(n4644) );
  XOR U4826 ( .A(a[62]), .B(b[7]), .Z(n4707) );
  NAND U4827 ( .A(n4708), .B(n4707), .Z(n4643) );
  NAND U4828 ( .A(n4644), .B(n4643), .Z(n4693) );
  NAND U4829 ( .A(n4950), .B(n4645), .Z(n4647) );
  XOR U4830 ( .A(b[11]), .B(a[58]), .Z(n4709) );
  NAND U4831 ( .A(n4863), .B(n4709), .Z(n4646) );
  NAND U4832 ( .A(n4647), .B(n4646), .Z(n4692) );
  XOR U4833 ( .A(b[13]), .B(a[56]), .Z(n4701) );
  XOR U4834 ( .A(n4681), .B(n4682), .Z(n4684) );
  XNOR U4835 ( .A(n4683), .B(n4684), .Z(n4676) );
  NAND U4836 ( .A(n4650), .B(n4649), .Z(n4654) );
  NAND U4837 ( .A(n4652), .B(n4651), .Z(n4653) );
  NAND U4838 ( .A(n4654), .B(n4653), .Z(n4675) );
  XOR U4839 ( .A(n4676), .B(n4675), .Z(n4677) );
  NAND U4840 ( .A(n4656), .B(n4655), .Z(n4660) );
  NAND U4841 ( .A(n4658), .B(n4657), .Z(n4659) );
  AND U4842 ( .A(n4660), .B(n4659), .Z(n4670) );
  XOR U4843 ( .A(n4669), .B(n4670), .Z(n4671) );
  XOR U4844 ( .A(n4672), .B(n4671), .Z(n4663) );
  XOR U4845 ( .A(n4666), .B(n4665), .Z(n4661) );
  XOR U4846 ( .A(n4662), .B(n4661), .Z(c[116]) );
  AND U4847 ( .A(n4662), .B(n4661), .Z(n4720) );
  NAND U4848 ( .A(n4664), .B(n4663), .Z(n4668) );
  NANDN U4849 ( .A(n4666), .B(n4665), .Z(n4667) );
  AND U4850 ( .A(n4668), .B(n4667), .Z(n4724) );
  NAND U4851 ( .A(n4670), .B(n4669), .Z(n4674) );
  NAND U4852 ( .A(n4672), .B(n4671), .Z(n4673) );
  NAND U4853 ( .A(n4674), .B(n4673), .Z(n4722) );
  NAND U4854 ( .A(n4676), .B(n4675), .Z(n4680) );
  NAND U4855 ( .A(n4678), .B(n4677), .Z(n4679) );
  AND U4856 ( .A(n4680), .B(n4679), .Z(n4730) );
  NAND U4857 ( .A(n4682), .B(n4681), .Z(n4686) );
  NAND U4858 ( .A(n4684), .B(n4683), .Z(n4685) );
  NAND U4859 ( .A(n4686), .B(n4685), .Z(n4736) );
  NANDN U4860 ( .A(n4687), .B(n4765), .Z(n4691) );
  NAND U4861 ( .A(n4689), .B(n4688), .Z(n4690) );
  AND U4862 ( .A(n4691), .B(n4690), .Z(n4734) );
  NAND U4863 ( .A(n4693), .B(n4692), .Z(n4697) );
  NAND U4864 ( .A(n4695), .B(n4694), .Z(n4696) );
  AND U4865 ( .A(n4697), .B(n4696), .Z(n4742) );
  NAND U4866 ( .A(n41), .B(n4698), .Z(n4700) );
  XOR U4867 ( .A(a[61]), .B(b[9]), .Z(n4746) );
  NAND U4868 ( .A(n4810), .B(n4746), .Z(n4699) );
  NAND U4869 ( .A(n4700), .B(n4699), .Z(n4762) );
  NAND U4870 ( .A(n5012), .B(n4701), .Z(n4703) );
  XOR U4871 ( .A(b[13]), .B(a[57]), .Z(n4749) );
  NAND U4872 ( .A(n4985), .B(n4749), .Z(n4702) );
  NAND U4873 ( .A(n4703), .B(n4702), .Z(n4760) );
  NAND U4874 ( .A(n42), .B(n4704), .Z(n4706) );
  XOR U4875 ( .A(b[15]), .B(a[55]), .Z(n4752) );
  NAND U4876 ( .A(n4981), .B(n4752), .Z(n4705) );
  NAND U4877 ( .A(n4706), .B(n4705), .Z(n4759) );
  XNOR U4878 ( .A(a[63]), .B(b[7]), .Z(n4756) );
  NAND U4879 ( .A(n4950), .B(n4709), .Z(n4711) );
  XOR U4880 ( .A(b[11]), .B(a[59]), .Z(n4745) );
  NAND U4881 ( .A(n4863), .B(n4745), .Z(n4710) );
  NAND U4882 ( .A(n4711), .B(n4710), .Z(n4771) );
  XNOR U4883 ( .A(n4712), .B(n4766), .Z(n4767) );
  AND U4884 ( .A(b[15]), .B(a[53]), .Z(n4768) );
  XNOR U4885 ( .A(n4774), .B(n4773), .Z(n4739) );
  XOR U4886 ( .A(n4740), .B(n4739), .Z(n4741) );
  XOR U4887 ( .A(n4742), .B(n4741), .Z(n4733) );
  XOR U4888 ( .A(n4734), .B(n4733), .Z(n4735) );
  NAND U4889 ( .A(n4714), .B(n4713), .Z(n4718) );
  NAND U4890 ( .A(n4716), .B(n4715), .Z(n4717) );
  AND U4891 ( .A(n4718), .B(n4717), .Z(n4728) );
  XOR U4892 ( .A(n4727), .B(n4728), .Z(n4729) );
  XOR U4893 ( .A(n4730), .B(n4729), .Z(n4721) );
  XOR U4894 ( .A(n4724), .B(n4723), .Z(n4719) );
  XOR U4895 ( .A(n4720), .B(n4719), .Z(c[117]) );
  AND U4896 ( .A(n4720), .B(n4719), .Z(n4778) );
  NAND U4897 ( .A(n4722), .B(n4721), .Z(n4726) );
  NANDN U4898 ( .A(n4724), .B(n4723), .Z(n4725) );
  AND U4899 ( .A(n4726), .B(n4725), .Z(n4782) );
  NAND U4900 ( .A(n4728), .B(n4727), .Z(n4732) );
  NANDN U4901 ( .A(n4730), .B(n4729), .Z(n4731) );
  AND U4902 ( .A(n4732), .B(n4731), .Z(n4780) );
  NAND U4903 ( .A(n4734), .B(n4733), .Z(n4738) );
  NAND U4904 ( .A(n4736), .B(n4735), .Z(n4737) );
  NAND U4905 ( .A(n4738), .B(n4737), .Z(n4788) );
  NAND U4906 ( .A(n4740), .B(n4739), .Z(n4744) );
  NAND U4907 ( .A(n4742), .B(n4741), .Z(n4743) );
  NAND U4908 ( .A(n4744), .B(n4743), .Z(n4786) );
  XNOR U4909 ( .A(b[11]), .B(a[60]), .Z(n4815) );
  NAND U4910 ( .A(n41), .B(n4746), .Z(n4748) );
  XOR U4911 ( .A(a[62]), .B(b[9]), .Z(n4809) );
  NAND U4912 ( .A(n4810), .B(n4809), .Z(n4747) );
  NAND U4913 ( .A(n4748), .B(n4747), .Z(n4804) );
  NAND U4914 ( .A(n5012), .B(n4749), .Z(n4751) );
  XOR U4915 ( .A(b[13]), .B(a[58]), .Z(n4811) );
  NAND U4916 ( .A(n4985), .B(n4811), .Z(n4750) );
  NAND U4917 ( .A(n4751), .B(n4750), .Z(n4803) );
  NAND U4918 ( .A(n42), .B(n4752), .Z(n4754) );
  XOR U4919 ( .A(b[15]), .B(a[56]), .Z(n4818) );
  NAND U4920 ( .A(n4981), .B(n4818), .Z(n4753) );
  AND U4921 ( .A(n4754), .B(n4753), .Z(n4824) );
  NANDN U4922 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U4923 ( .A(n4758), .B(n4757), .Z(n4822) );
  AND U4924 ( .A(b[15]), .B(a[54]), .Z(n4856) );
  IV U4925 ( .A(n4856), .Z(n4821) );
  XNOR U4926 ( .A(n4822), .B(n4821), .Z(n4823) );
  XOR U4927 ( .A(n4824), .B(n4823), .Z(n4797) );
  XOR U4928 ( .A(n4798), .B(n4797), .Z(n4800) );
  NAND U4929 ( .A(n4760), .B(n4759), .Z(n4764) );
  NAND U4930 ( .A(n4762), .B(n4761), .Z(n4763) );
  AND U4931 ( .A(n4764), .B(n4763), .Z(n4799) );
  XOR U4932 ( .A(n4800), .B(n4799), .Z(n4794) );
  OR U4933 ( .A(n4766), .B(n4765), .Z(n4770) );
  NAND U4934 ( .A(n4768), .B(n4767), .Z(n4769) );
  NAND U4935 ( .A(n4770), .B(n4769), .Z(n4792) );
  NAND U4936 ( .A(n4772), .B(n4771), .Z(n4776) );
  NAND U4937 ( .A(n4774), .B(n4773), .Z(n4775) );
  NAND U4938 ( .A(n4776), .B(n4775), .Z(n4791) );
  XOR U4939 ( .A(n4794), .B(n4793), .Z(n4785) );
  XOR U4940 ( .A(n4780), .B(n4779), .Z(n4781) );
  XOR U4941 ( .A(n4782), .B(n4781), .Z(n4777) );
  XOR U4942 ( .A(n4778), .B(n4777), .Z(c[118]) );
  AND U4943 ( .A(n4778), .B(n4777), .Z(n4828) );
  NAND U4944 ( .A(n4780), .B(n4779), .Z(n4784) );
  NANDN U4945 ( .A(n4782), .B(n4781), .Z(n4783) );
  AND U4946 ( .A(n4784), .B(n4783), .Z(n4832) );
  NAND U4947 ( .A(n4786), .B(n4785), .Z(n4790) );
  NAND U4948 ( .A(n4788), .B(n4787), .Z(n4789) );
  NAND U4949 ( .A(n4790), .B(n4789), .Z(n4830) );
  NAND U4950 ( .A(n4792), .B(n4791), .Z(n4796) );
  NANDN U4951 ( .A(n4794), .B(n4793), .Z(n4795) );
  AND U4952 ( .A(n4796), .B(n4795), .Z(n4838) );
  NAND U4953 ( .A(n4798), .B(n4797), .Z(n4802) );
  NAND U4954 ( .A(n4800), .B(n4799), .Z(n4801) );
  AND U4955 ( .A(n4802), .B(n4801), .Z(n4836) );
  NAND U4956 ( .A(n4804), .B(n4803), .Z(n4808) );
  NAND U4957 ( .A(n4806), .B(n4805), .Z(n4807) );
  NAND U4958 ( .A(n4808), .B(n4807), .Z(n4844) );
  XNOR U4959 ( .A(a[63]), .B(b[9]), .Z(n4867) );
  NAND U4960 ( .A(n5012), .B(n4811), .Z(n4813) );
  XOR U4961 ( .A(b[13]), .B(a[59]), .Z(n4859) );
  NAND U4962 ( .A(n4985), .B(n4859), .Z(n4812) );
  NAND U4963 ( .A(n4813), .B(n4812), .Z(n4870) );
  AND U4964 ( .A(b[15]), .B(a[55]), .Z(n4853) );
  XNOR U4965 ( .A(n4853), .B(n4814), .Z(n4855) );
  XNOR U4966 ( .A(n4821), .B(n4855), .Z(n4872) );
  XNOR U4967 ( .A(n4873), .B(n4872), .Z(n4848) );
  NANDN U4968 ( .A(n4815), .B(n4950), .Z(n4817) );
  XOR U4969 ( .A(a[61]), .B(b[11]), .Z(n4862) );
  NANDN U4970 ( .A(n40), .B(n4862), .Z(n4816) );
  AND U4971 ( .A(n4817), .B(n4816), .Z(n4847) );
  NANDN U4972 ( .A(n31), .B(n4818), .Z(n4820) );
  XOR U4973 ( .A(b[15]), .B(a[57]), .Z(n4864) );
  NANDN U4974 ( .A(n5051), .B(n4864), .Z(n4819) );
  AND U4975 ( .A(n4820), .B(n4819), .Z(n4849) );
  XNOR U4976 ( .A(n4850), .B(n4849), .Z(n4842) );
  NANDN U4977 ( .A(n4822), .B(n4821), .Z(n4826) );
  NANDN U4978 ( .A(n4824), .B(n4823), .Z(n4825) );
  NAND U4979 ( .A(n4826), .B(n4825), .Z(n4841) );
  XOR U4980 ( .A(n4836), .B(n4835), .Z(n4837) );
  XOR U4981 ( .A(n4838), .B(n4837), .Z(n4829) );
  XOR U4982 ( .A(n4832), .B(n4831), .Z(n4827) );
  XOR U4983 ( .A(n4828), .B(n4827), .Z(c[119]) );
  AND U4984 ( .A(n4828), .B(n4827), .Z(n4877) );
  NAND U4985 ( .A(n4830), .B(n4829), .Z(n4834) );
  NANDN U4986 ( .A(n4832), .B(n4831), .Z(n4833) );
  AND U4987 ( .A(n4834), .B(n4833), .Z(n4881) );
  NAND U4988 ( .A(n4836), .B(n4835), .Z(n4840) );
  NANDN U4989 ( .A(n4838), .B(n4837), .Z(n4839) );
  AND U4990 ( .A(n4840), .B(n4839), .Z(n4879) );
  NAND U4991 ( .A(n4842), .B(n4841), .Z(n4846) );
  NAND U4992 ( .A(n4844), .B(n4843), .Z(n4845) );
  AND U4993 ( .A(n4846), .B(n4845), .Z(n4887) );
  NAND U4994 ( .A(n4848), .B(n4847), .Z(n4852) );
  NAND U4995 ( .A(n4850), .B(n4849), .Z(n4851) );
  NAND U4996 ( .A(n4852), .B(n4851), .Z(n4885) );
  NAND U4997 ( .A(n4854), .B(n4853), .Z(n4858) );
  NAND U4998 ( .A(n4856), .B(n4855), .Z(n4857) );
  NAND U4999 ( .A(n4858), .B(n4857), .Z(n4909) );
  NAND U5000 ( .A(n5012), .B(n4859), .Z(n4861) );
  XOR U5001 ( .A(b[13]), .B(a[60]), .Z(n4895) );
  NAND U5002 ( .A(n4985), .B(n4895), .Z(n4860) );
  NAND U5003 ( .A(n4861), .B(n4860), .Z(n4907) );
  XNOR U5004 ( .A(a[62]), .B(b[11]), .Z(n4903) );
  NAND U5005 ( .A(n42), .B(n4864), .Z(n4866) );
  XOR U5006 ( .A(b[15]), .B(a[58]), .Z(n4898) );
  NAND U5007 ( .A(n4981), .B(n4898), .Z(n4865) );
  NAND U5008 ( .A(n4866), .B(n4865), .Z(n4892) );
  NANDN U5009 ( .A(n4867), .B(n41), .Z(n4868) );
  AND U5010 ( .A(n4869), .B(n4868), .Z(n4890) );
  AND U5011 ( .A(b[15]), .B(a[56]), .Z(n4944) );
  IV U5012 ( .A(n4944), .Z(n4902) );
  XNOR U5013 ( .A(n4890), .B(n4902), .Z(n4891) );
  NAND U5014 ( .A(n4871), .B(n4870), .Z(n4875) );
  NAND U5015 ( .A(n4873), .B(n4872), .Z(n4874) );
  AND U5016 ( .A(n4875), .B(n4874), .Z(n4913) );
  XOR U5017 ( .A(n4912), .B(n4913), .Z(n4915) );
  XOR U5018 ( .A(n4914), .B(n4915), .Z(n4884) );
  XOR U5019 ( .A(n4887), .B(n4886), .Z(n4878) );
  XOR U5020 ( .A(n4879), .B(n4878), .Z(n4880) );
  XOR U5021 ( .A(n4881), .B(n4880), .Z(n4876) );
  XOR U5022 ( .A(n4877), .B(n4876), .Z(c[120]) );
  AND U5023 ( .A(n4877), .B(n4876), .Z(n4919) );
  NAND U5024 ( .A(n4879), .B(n4878), .Z(n4883) );
  NANDN U5025 ( .A(n4881), .B(n4880), .Z(n4882) );
  AND U5026 ( .A(n4883), .B(n4882), .Z(n4923) );
  NAND U5027 ( .A(n4885), .B(n4884), .Z(n4889) );
  NAND U5028 ( .A(n4887), .B(n4886), .Z(n4888) );
  NAND U5029 ( .A(n4889), .B(n4888), .Z(n4921) );
  NANDN U5030 ( .A(n4890), .B(n4902), .Z(n4894) );
  NAND U5031 ( .A(n4892), .B(n4891), .Z(n4893) );
  AND U5032 ( .A(n4894), .B(n4893), .Z(n4935) );
  NAND U5033 ( .A(n5012), .B(n4895), .Z(n4897) );
  XOR U5034 ( .A(b[13]), .B(a[61]), .Z(n4938) );
  NAND U5035 ( .A(n4985), .B(n4938), .Z(n4896) );
  NAND U5036 ( .A(n4897), .B(n4896), .Z(n4955) );
  NAND U5037 ( .A(n42), .B(n4898), .Z(n4900) );
  XOR U5038 ( .A(b[15]), .B(a[59]), .Z(n4947) );
  NAND U5039 ( .A(n4981), .B(n4947), .Z(n4899) );
  NAND U5040 ( .A(n4900), .B(n4899), .Z(n4954) );
  AND U5041 ( .A(b[15]), .B(a[57]), .Z(n4941) );
  XNOR U5042 ( .A(n4941), .B(n4901), .Z(n4943) );
  XNOR U5043 ( .A(n4902), .B(n4943), .Z(n4956) );
  XNOR U5044 ( .A(n4957), .B(n4956), .Z(n4933) );
  NANDN U5045 ( .A(n4903), .B(n4950), .Z(n4905) );
  XNOR U5046 ( .A(a[63]), .B(b[11]), .Z(n4951) );
  OR U5047 ( .A(n4951), .B(n40), .Z(n4904) );
  AND U5048 ( .A(n4905), .B(n4904), .Z(n4932) );
  XNOR U5049 ( .A(n4935), .B(n4934), .Z(n4927) );
  NAND U5050 ( .A(n4907), .B(n4906), .Z(n4911) );
  NAND U5051 ( .A(n4909), .B(n4908), .Z(n4910) );
  NAND U5052 ( .A(n4911), .B(n4910), .Z(n4926) );
  NAND U5053 ( .A(n4913), .B(n4912), .Z(n4917) );
  NAND U5054 ( .A(n4915), .B(n4914), .Z(n4916) );
  AND U5055 ( .A(n4917), .B(n4916), .Z(n4928) );
  XNOR U5056 ( .A(n4929), .B(n4928), .Z(n4920) );
  XOR U5057 ( .A(n4923), .B(n4922), .Z(n4918) );
  XOR U5058 ( .A(n4919), .B(n4918), .Z(c[121]) );
  AND U5059 ( .A(n4919), .B(n4918), .Z(n4961) );
  NAND U5060 ( .A(n4921), .B(n4920), .Z(n4925) );
  NANDN U5061 ( .A(n4923), .B(n4922), .Z(n4924) );
  AND U5062 ( .A(n4925), .B(n4924), .Z(n4965) );
  NAND U5063 ( .A(n4927), .B(n4926), .Z(n4931) );
  NAND U5064 ( .A(n4929), .B(n4928), .Z(n4930) );
  AND U5065 ( .A(n4931), .B(n4930), .Z(n4963) );
  NAND U5066 ( .A(n4933), .B(n4932), .Z(n4937) );
  NAND U5067 ( .A(n4935), .B(n4934), .Z(n4936) );
  NAND U5068 ( .A(n4937), .B(n4936), .Z(n4989) );
  NAND U5069 ( .A(n5012), .B(n4938), .Z(n4940) );
  XOR U5070 ( .A(a[62]), .B(b[13]), .Z(n4984) );
  NAND U5071 ( .A(n4985), .B(n4984), .Z(n4939) );
  NAND U5072 ( .A(n4940), .B(n4939), .Z(n4969) );
  NAND U5073 ( .A(n4942), .B(n4941), .Z(n4946) );
  NAND U5074 ( .A(n4944), .B(n4943), .Z(n4945) );
  NAND U5075 ( .A(n4946), .B(n4945), .Z(n4968) );
  NAND U5076 ( .A(n42), .B(n4947), .Z(n4949) );
  XOR U5077 ( .A(b[15]), .B(a[60]), .Z(n4980) );
  NAND U5078 ( .A(n4981), .B(n4980), .Z(n4948) );
  NAND U5079 ( .A(n4949), .B(n4948), .Z(n4977) );
  NANDN U5080 ( .A(n4951), .B(n4950), .Z(n4952) );
  AND U5081 ( .A(n4953), .B(n4952), .Z(n4975) );
  AND U5082 ( .A(b[15]), .B(a[58]), .Z(n5009) );
  IV U5083 ( .A(n5009), .Z(n4974) );
  XNOR U5084 ( .A(n4975), .B(n4974), .Z(n4976) );
  XNOR U5085 ( .A(n4971), .B(n4970), .Z(n4987) );
  NAND U5086 ( .A(n4955), .B(n4954), .Z(n4959) );
  NAND U5087 ( .A(n4957), .B(n4956), .Z(n4958) );
  AND U5088 ( .A(n4959), .B(n4958), .Z(n4986) );
  XOR U5089 ( .A(n4963), .B(n4962), .Z(n4964) );
  XOR U5090 ( .A(n4965), .B(n4964), .Z(n4960) );
  XOR U5091 ( .A(n4961), .B(n4960), .Z(c[122]) );
  AND U5092 ( .A(n4961), .B(n4960), .Z(n4993) );
  NAND U5093 ( .A(n4963), .B(n4962), .Z(n4967) );
  NANDN U5094 ( .A(n4965), .B(n4964), .Z(n4966) );
  AND U5095 ( .A(n4967), .B(n4966), .Z(n4997) );
  NAND U5096 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U5097 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U5098 ( .A(n4973), .B(n4972), .Z(n5022) );
  NANDN U5099 ( .A(n4975), .B(n4974), .Z(n4979) );
  NAND U5100 ( .A(n4977), .B(n4976), .Z(n4978) );
  NAND U5101 ( .A(n4979), .B(n4978), .Z(n5020) );
  NAND U5102 ( .A(n42), .B(n4980), .Z(n4983) );
  XOR U5103 ( .A(b[15]), .B(a[61]), .Z(n5016) );
  NAND U5104 ( .A(n4981), .B(n5016), .Z(n4982) );
  NAND U5105 ( .A(n4983), .B(n4982), .Z(n5001) );
  XNOR U5106 ( .A(a[63]), .B(b[13]), .Z(n5013) );
  AND U5107 ( .A(b[15]), .B(a[59]), .Z(n5006) );
  XOR U5108 ( .A(n5009), .B(n5008), .Z(n5002) );
  XOR U5109 ( .A(n5003), .B(n5002), .Z(n5019) );
  NAND U5110 ( .A(n4987), .B(n4986), .Z(n4991) );
  NAND U5111 ( .A(n4989), .B(n4988), .Z(n4990) );
  NAND U5112 ( .A(n4991), .B(n4990), .Z(n4994) );
  XOR U5113 ( .A(n4995), .B(n4994), .Z(n4996) );
  XOR U5114 ( .A(n4997), .B(n4996), .Z(n4992) );
  XOR U5115 ( .A(n4993), .B(n4992), .Z(c[123]) );
  AND U5116 ( .A(n4993), .B(n4992), .Z(n5026) );
  NAND U5117 ( .A(n4995), .B(n4994), .Z(n4999) );
  NANDN U5118 ( .A(n4997), .B(n4996), .Z(n4998) );
  AND U5119 ( .A(n4999), .B(n4998), .Z(n5030) );
  NAND U5120 ( .A(n5001), .B(n5000), .Z(n5005) );
  NAND U5121 ( .A(n5003), .B(n5002), .Z(n5004) );
  NAND U5122 ( .A(n5005), .B(n5004), .Z(n5036) );
  NAND U5123 ( .A(n5007), .B(n5006), .Z(n5011) );
  NAND U5124 ( .A(n5009), .B(n5008), .Z(n5010) );
  NAND U5125 ( .A(n5011), .B(n5010), .Z(n5034) );
  NANDN U5126 ( .A(n5013), .B(n5012), .Z(n5014) );
  AND U5127 ( .A(n5015), .B(n5014), .Z(n5039) );
  AND U5128 ( .A(b[15]), .B(a[60]), .Z(n5057) );
  XOR U5129 ( .A(n5039), .B(n5057), .Z(n5041) );
  NANDN U5130 ( .A(n31), .B(n5016), .Z(n5018) );
  XNOR U5131 ( .A(b[15]), .B(a[62]), .Z(n5044) );
  OR U5132 ( .A(n5044), .B(n5051), .Z(n5017) );
  NAND U5133 ( .A(n5018), .B(n5017), .Z(n5040) );
  XOR U5134 ( .A(n5041), .B(n5040), .Z(n5033) );
  NAND U5135 ( .A(n5020), .B(n5019), .Z(n5024) );
  NAND U5136 ( .A(n5022), .B(n5021), .Z(n5023) );
  AND U5137 ( .A(n5024), .B(n5023), .Z(n5028) );
  XOR U5138 ( .A(n5027), .B(n5028), .Z(n5029) );
  XOR U5139 ( .A(n5030), .B(n5029), .Z(n5025) );
  XOR U5140 ( .A(n5026), .B(n5025), .Z(c[124]) );
  AND U5141 ( .A(n5026), .B(n5025), .Z(n5049) );
  NAND U5142 ( .A(n5028), .B(n5027), .Z(n5032) );
  NANDN U5143 ( .A(n5030), .B(n5029), .Z(n5031) );
  AND U5144 ( .A(n5032), .B(n5031), .Z(n5063) );
  NAND U5145 ( .A(n5034), .B(n5033), .Z(n5038) );
  NAND U5146 ( .A(n5036), .B(n5035), .Z(n5037) );
  AND U5147 ( .A(n5038), .B(n5037), .Z(n5061) );
  OR U5148 ( .A(n5039), .B(n5057), .Z(n5043) );
  NAND U5149 ( .A(n5041), .B(n5040), .Z(n5042) );
  AND U5150 ( .A(n5043), .B(n5042), .Z(n5069) );
  OR U5151 ( .A(n5044), .B(n31), .Z(n5046) );
  XNOR U5152 ( .A(b[15]), .B(a[63]), .Z(n5050) );
  OR U5153 ( .A(n5050), .B(n5051), .Z(n5045) );
  AND U5154 ( .A(n5046), .B(n5045), .Z(n5067) );
  AND U5155 ( .A(b[15]), .B(a[61]), .Z(n5054) );
  XNOR U5156 ( .A(n5054), .B(n5047), .Z(n5056) );
  XNOR U5157 ( .A(n5057), .B(n5056), .Z(n5066) );
  XOR U5158 ( .A(n5067), .B(n5066), .Z(n5068) );
  XOR U5159 ( .A(n5069), .B(n5068), .Z(n5060) );
  XOR U5160 ( .A(n5061), .B(n5060), .Z(n5062) );
  XOR U5161 ( .A(n5063), .B(n5062), .Z(n5048) );
  XOR U5162 ( .A(n5049), .B(n5048), .Z(c[125]) );
  AND U5163 ( .A(n5049), .B(n5048), .Z(n5073) );
  NAND U5164 ( .A(b[15]), .B(a[62]), .Z(n5082) );
  OR U5165 ( .A(n5050), .B(n31), .Z(n5053) );
  NANDN U5166 ( .A(n5051), .B(b[15]), .Z(n5052) );
  NAND U5167 ( .A(n5053), .B(n5052), .Z(n5085) );
  NAND U5168 ( .A(n5055), .B(n5054), .Z(n5059) );
  NAND U5169 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U5170 ( .A(n5059), .B(n5058), .Z(n5084) );
  XOR U5171 ( .A(n5085), .B(n5084), .Z(n5083) );
  NAND U5172 ( .A(n5061), .B(n5060), .Z(n5065) );
  NANDN U5173 ( .A(n5063), .B(n5062), .Z(n5064) );
  NAND U5174 ( .A(n5065), .B(n5064), .Z(n5074) );
  NAND U5175 ( .A(n5067), .B(n5066), .Z(n5071) );
  NAND U5176 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U5177 ( .A(n5071), .B(n5070), .Z(n5075) );
  XNOR U5178 ( .A(n5076), .B(n5077), .Z(n5072) );
  XOR U5179 ( .A(n5073), .B(n5072), .Z(c[126]) );
  NAND U5180 ( .A(n5073), .B(n5072), .Z(n5081) );
  AND U5181 ( .A(n5075), .B(n5074), .Z(n5079) );
  AND U5182 ( .A(n5077), .B(n5076), .Z(n5078) );
  OR U5183 ( .A(n5079), .B(n5078), .Z(n5080) );
  AND U5184 ( .A(n5081), .B(n5080), .Z(n5094) );
  NAND U5185 ( .A(n5083), .B(n5082), .Z(n5087) );
  NAND U5186 ( .A(n5085), .B(n5084), .Z(n5086) );
  AND U5187 ( .A(n5087), .B(n5086), .Z(n5092) );
  XNOR U5188 ( .A(a[62]), .B(a[63]), .Z(n5088) );
  XNOR U5189 ( .A(n5089), .B(n5088), .Z(n5090) );
  NAND U5190 ( .A(b[15]), .B(n5090), .Z(n5091) );
  XNOR U5191 ( .A(n5092), .B(n5091), .Z(n5093) );
  XNOR U5192 ( .A(n5094), .B(n5093), .Z(c[127]) );
endmodule

